module xpb_first
(
    input [263:0] data_in0,
    input [263:0] data_in1,

    output [105:0] col_out_0,
    output [105:0] col_out_1,
    output [105:0] col_out_2,
    output [105:0] col_out_3,
    output [105:0] col_out_4,
    output [105:0] col_out_5,
    output [105:0] col_out_6,
    output [105:0] col_out_7,
    output [105:0] col_out_8,
    output [105:0] col_out_9,
    output [105:0] col_out_10,
    output [105:0] col_out_11,
    output [105:0] col_out_12,
    output [105:0] col_out_13,
    output [105:0] col_out_14,
    output [105:0] col_out_15,
    output [105:0] col_out_16,
    output [105:0] col_out_17,
    output [105:0] col_out_18,
    output [105:0] col_out_19,
    output [105:0] col_out_20,
    output [105:0] col_out_21,
    output [105:0] col_out_22,
    output [105:0] col_out_23,
    output [105:0] col_out_24,
    output [105:0] col_out_25,
    output [105:0] col_out_26,
    output [105:0] col_out_27,
    output [105:0] col_out_28,
    output [105:0] col_out_29,
    output [105:0] col_out_30,
    output [105:0] col_out_31,
    output [105:0] col_out_32,
    output [105:0] col_out_33,
    output [105:0] col_out_34,
    output [105:0] col_out_35,
    output [105:0] col_out_36,
    output [105:0] col_out_37,
    output [105:0] col_out_38,
    output [105:0] col_out_39,
    output [105:0] col_out_40,
    output [105:0] col_out_41,
    output [105:0] col_out_42,
    output [105:0] col_out_43,
    output [105:0] col_out_44,
    output [105:0] col_out_45,
    output [105:0] col_out_46,
    output [105:0] col_out_47,
    output [105:0] col_out_48,
    output [105:0] col_out_49,
    output [105:0] col_out_50,
    output [105:0] col_out_51,
    output [105:0] col_out_52,
    output [105:0] col_out_53,
    output [105:0] col_out_54,
    output [105:0] col_out_55,
    output [105:0] col_out_56,
    output [105:0] col_out_57,
    output [105:0] col_out_58,
    output [105:0] col_out_59,
    output [105:0] col_out_60,
    output [105:0] col_out_61,
    output [105:0] col_out_62,
    output [105:0] col_out_63,
    output [105:0] col_out_64,
    output [105:0] col_out_65,
    output [105:0] col_out_66,
    output [105:0] col_out_67,
    output [105:0] col_out_68,
    output [105:0] col_out_69,
    output [105:0] col_out_70,
    output [105:0] col_out_71,
    output [105:0] col_out_72,
    output [105:0] col_out_73,
    output [105:0] col_out_74,
    output [105:0] col_out_75,
    output [105:0] col_out_76,
    output [105:0] col_out_77,
    output [105:0] col_out_78,
    output [105:0] col_out_79,
    output [105:0] col_out_80,
    output [105:0] col_out_81,
    output [105:0] col_out_82,
    output [105:0] col_out_83,
    output [105:0] col_out_84,
    output [105:0] col_out_85,
    output [105:0] col_out_86,
    output [105:0] col_out_87,
    output [105:0] col_out_88,
    output [105:0] col_out_89,
    output [105:0] col_out_90,
    output [105:0] col_out_91,
    output [105:0] col_out_92,
    output [105:0] col_out_93,
    output [105:0] col_out_94,
    output [105:0] col_out_95,
    output [105:0] col_out_96,
    output [105:0] col_out_97,
    output [105:0] col_out_98,
    output [105:0] col_out_99,
    output [105:0] col_out_100,
    output [105:0] col_out_101,
    output [105:0] col_out_102,
    output [105:0] col_out_103,
    output [105:0] col_out_104,
    output [105:0] col_out_105,
    output [105:0] col_out_106,
    output [105:0] col_out_107,
    output [105:0] col_out_108,
    output [105:0] col_out_109,
    output [105:0] col_out_110,
    output [105:0] col_out_111,
    output [105:0] col_out_112,
    output [105:0] col_out_113,
    output [105:0] col_out_114,
    output [105:0] col_out_115,
    output [105:0] col_out_116,
    output [105:0] col_out_117,
    output [105:0] col_out_118,
    output [105:0] col_out_119,
    output [105:0] col_out_120,
    output [105:0] col_out_121,
    output [105:0] col_out_122,
    output [105:0] col_out_123,
    output [105:0] col_out_124,
    output [105:0] col_out_125,
    output [105:0] col_out_126,
    output [105:0] col_out_127,
    output [105:0] col_out_128,
    output [105:0] col_out_129,
    output [105:0] col_out_130,
    output [105:0] col_out_131,
    output [105:0] col_out_132,
    output [105:0] col_out_133,
    output [105:0] col_out_134,
    output [105:0] col_out_135,
    output [105:0] col_out_136,
    output [105:0] col_out_137,
    output [105:0] col_out_138,
    output [105:0] col_out_139,
    output [105:0] col_out_140,
    output [105:0] col_out_141,
    output [105:0] col_out_142,
    output [105:0] col_out_143,
    output [105:0] col_out_144,
    output [105:0] col_out_145,
    output [105:0] col_out_146,
    output [105:0] col_out_147,
    output [105:0] col_out_148,
    output [105:0] col_out_149,
    output [105:0] col_out_150,
    output [105:0] col_out_151,
    output [105:0] col_out_152,
    output [105:0] col_out_153,
    output [105:0] col_out_154,
    output [105:0] col_out_155,
    output [105:0] col_out_156,
    output [105:0] col_out_157,
    output [105:0] col_out_158,
    output [105:0] col_out_159,
    output [105:0] col_out_160,
    output [105:0] col_out_161,
    output [105:0] col_out_162,
    output [105:0] col_out_163,
    output [105:0] col_out_164,
    output [105:0] col_out_165,
    output [105:0] col_out_166,
    output [105:0] col_out_167,
    output [105:0] col_out_168,
    output [105:0] col_out_169,
    output [105:0] col_out_170,
    output [105:0] col_out_171,
    output [105:0] col_out_172,
    output [105:0] col_out_173,
    output [105:0] col_out_174,
    output [105:0] col_out_175,
    output [105:0] col_out_176,
    output [105:0] col_out_177,
    output [105:0] col_out_178,
    output [105:0] col_out_179,
    output [105:0] col_out_180,
    output [105:0] col_out_181,
    output [105:0] col_out_182,
    output [105:0] col_out_183,
    output [105:0] col_out_184,
    output [105:0] col_out_185,
    output [105:0] col_out_186,
    output [105:0] col_out_187,
    output [105:0] col_out_188,
    output [105:0] col_out_189,
    output [105:0] col_out_190,
    output [105:0] col_out_191,
    output [105:0] col_out_192,
    output [105:0] col_out_193,
    output [105:0] col_out_194,
    output [105:0] col_out_195,
    output [105:0] col_out_196,
    output [105:0] col_out_197,
    output [105:0] col_out_198,
    output [105:0] col_out_199,
    output [105:0] col_out_200,
    output [105:0] col_out_201,
    output [105:0] col_out_202,
    output [105:0] col_out_203,
    output [105:0] col_out_204,
    output [105:0] col_out_205,
    output [105:0] col_out_206,
    output [105:0] col_out_207,
    output [105:0] col_out_208,
    output [105:0] col_out_209,
    output [105:0] col_out_210,
    output [105:0] col_out_211,
    output [105:0] col_out_212,
    output [105:0] col_out_213,
    output [105:0] col_out_214,
    output [105:0] col_out_215,
    output [105:0] col_out_216,
    output [105:0] col_out_217,
    output [105:0] col_out_218,
    output [105:0] col_out_219,
    output [105:0] col_out_220,
    output [105:0] col_out_221,
    output [105:0] col_out_222,
    output [105:0] col_out_223,
    output [105:0] col_out_224,
    output [105:0] col_out_225,
    output [105:0] col_out_226,
    output [105:0] col_out_227,
    output [105:0] col_out_228,
    output [105:0] col_out_229,
    output [105:0] col_out_230,
    output [105:0] col_out_231,
    output [105:0] col_out_232,
    output [105:0] col_out_233,
    output [105:0] col_out_234,
    output [105:0] col_out_235,
    output [105:0] col_out_236,
    output [105:0] col_out_237,
    output [105:0] col_out_238,
    output [105:0] col_out_239,
    output [105:0] col_out_240,
    output [105:0] col_out_241,
    output [105:0] col_out_242,
    output [105:0] col_out_243,
    output [105:0] col_out_244,
    output [105:0] col_out_245,
    output [105:0] col_out_246,
    output [105:0] col_out_247,
    output [105:0] col_out_248,
    output [105:0] col_out_249,
    output [105:0] col_out_250,
    output [105:0] col_out_251,
    output [105:0] col_out_252,
    output [105:0] col_out_253,
    output [105:0] col_out_254,
    output [105:0] col_out_255,
    output [105:0] col_out_256,
    output [105:0] col_out_257,
    output [105:0] col_out_258,
    output [105:0] col_out_259,
    output [105:0] col_out_260,
    output [105:0] col_out_261,
    output [105:0] col_out_262,
    output [105:0] col_out_263,
    output [105:0] col_out_264,
    output [105:0] col_out_265,
    output [105:0] col_out_266,
    output [105:0] col_out_267,
    output [105:0] col_out_268,
    output [105:0] col_out_269,
    output [105:0] col_out_270,
    output [105:0] col_out_271,
    output [105:0] col_out_272,
    output [105:0] col_out_273,
    output [105:0] col_out_274,
    output [105:0] col_out_275,
    output [105:0] col_out_276,
    output [105:0] col_out_277,
    output [105:0] col_out_278,
    output [105:0] col_out_279,
    output [105:0] col_out_280,
    output [105:0] col_out_281,
    output [105:0] col_out_282,
    output [105:0] col_out_283,
    output [105:0] col_out_284,
    output [105:0] col_out_285,
    output [105:0] col_out_286,
    output [105:0] col_out_287,
    output [105:0] col_out_288,
    output [105:0] col_out_289,
    output [105:0] col_out_290,
    output [105:0] col_out_291,
    output [105:0] col_out_292,
    output [105:0] col_out_293,
    output [105:0] col_out_294,
    output [105:0] col_out_295,
    output [105:0] col_out_296,
    output [105:0] col_out_297,
    output [105:0] col_out_298,
    output [105:0] col_out_299,
    output [105:0] col_out_300,
    output [105:0] col_out_301,
    output [105:0] col_out_302,
    output [105:0] col_out_303,
    output [105:0] col_out_304,
    output [105:0] col_out_305,
    output [105:0] col_out_306,
    output [105:0] col_out_307,
    output [105:0] col_out_308,
    output [105:0] col_out_309,
    output [105:0] col_out_310,
    output [105:0] col_out_311,
    output [105:0] col_out_312,
    output [105:0] col_out_313,
    output [105:0] col_out_314,
    output [105:0] col_out_315,
    output [105:0] col_out_316,
    output [105:0] col_out_317,
    output [105:0] col_out_318,
    output [105:0] col_out_319,
    output [105:0] col_out_320,
    output [105:0] col_out_321,
    output [105:0] col_out_322,
    output [105:0] col_out_323,
    output [105:0] col_out_324,
    output [105:0] col_out_325,
    output [105:0] col_out_326,
    output [105:0] col_out_327,
    output [105:0] col_out_328,
    output [105:0] col_out_329,
    output [105:0] col_out_330,
    output [105:0] col_out_331,
    output [105:0] col_out_332,
    output [105:0] col_out_333,
    output [105:0] col_out_334,
    output [105:0] col_out_335,
    output [105:0] col_out_336,
    output [105:0] col_out_337,
    output [105:0] col_out_338,
    output [105:0] col_out_339,
    output [105:0] col_out_340,
    output [105:0] col_out_341,
    output [105:0] col_out_342,
    output [105:0] col_out_343,
    output [105:0] col_out_344,
    output [105:0] col_out_345,
    output [105:0] col_out_346,
    output [105:0] col_out_347,
    output [105:0] col_out_348,
    output [105:0] col_out_349,
    output [105:0] col_out_350,
    output [105:0] col_out_351,
    output [105:0] col_out_352,
    output [105:0] col_out_353,
    output [105:0] col_out_354,
    output [105:0] col_out_355,
    output [105:0] col_out_356,
    output [105:0] col_out_357,
    output [105:0] col_out_358,
    output [105:0] col_out_359,
    output [105:0] col_out_360,
    output [105:0] col_out_361,
    output [105:0] col_out_362,
    output [105:0] col_out_363,
    output [105:0] col_out_364,
    output [105:0] col_out_365,
    output [105:0] col_out_366,
    output [105:0] col_out_367,
    output [105:0] col_out_368,
    output [105:0] col_out_369,
    output [105:0] col_out_370,
    output [105:0] col_out_371,
    output [105:0] col_out_372,
    output [105:0] col_out_373,
    output [105:0] col_out_374,
    output [105:0] col_out_375,
    output [105:0] col_out_376,
    output [105:0] col_out_377,
    output [105:0] col_out_378,
    output [105:0] col_out_379,
    output [105:0] col_out_380,
    output [105:0] col_out_381,
    output [105:0] col_out_382,
    output [105:0] col_out_383,
    output [105:0] col_out_384,
    output [105:0] col_out_385,
    output [105:0] col_out_386,
    output [105:0] col_out_387,
    output [105:0] col_out_388,
    output [105:0] col_out_389,
    output [105:0] col_out_390,
    output [105:0] col_out_391,
    output [105:0] col_out_392,
    output [105:0] col_out_393,
    output [105:0] col_out_394,
    output [105:0] col_out_395,
    output [105:0] col_out_396,
    output [105:0] col_out_397,
    output [105:0] col_out_398,
    output [105:0] col_out_399,
    output [105:0] col_out_400,
    output [105:0] col_out_401,
    output [105:0] col_out_402,
    output [105:0] col_out_403,
    output [105:0] col_out_404,
    output [105:0] col_out_405,
    output [105:0] col_out_406,
    output [105:0] col_out_407,
    output [105:0] col_out_408,
    output [105:0] col_out_409,
    output [105:0] col_out_410,
    output [105:0] col_out_411,
    output [105:0] col_out_412,
    output [105:0] col_out_413,
    output [105:0] col_out_414,
    output [105:0] col_out_415,
    output [105:0] col_out_416,
    output [105:0] col_out_417,
    output [105:0] col_out_418,
    output [105:0] col_out_419,
    output [105:0] col_out_420,
    output [105:0] col_out_421,
    output [105:0] col_out_422,
    output [105:0] col_out_423,
    output [105:0] col_out_424,
    output [105:0] col_out_425,
    output [105:0] col_out_426,
    output [105:0] col_out_427,
    output [105:0] col_out_428,
    output [105:0] col_out_429,
    output [105:0] col_out_430,
    output [105:0] col_out_431,
    output [105:0] col_out_432,
    output [105:0] col_out_433,
    output [105:0] col_out_434,
    output [105:0] col_out_435,
    output [105:0] col_out_436,
    output [105:0] col_out_437,
    output [105:0] col_out_438,
    output [105:0] col_out_439,
    output [105:0] col_out_440,
    output [105:0] col_out_441,
    output [105:0] col_out_442,
    output [105:0] col_out_443,
    output [105:0] col_out_444,
    output [105:0] col_out_445,
    output [105:0] col_out_446,
    output [105:0] col_out_447,
    output [105:0] col_out_448,
    output [105:0] col_out_449,
    output [105:0] col_out_450,
    output [105:0] col_out_451,
    output [105:0] col_out_452,
    output [105:0] col_out_453,
    output [105:0] col_out_454,
    output [105:0] col_out_455,
    output [105:0] col_out_456,
    output [105:0] col_out_457,
    output [105:0] col_out_458,
    output [105:0] col_out_459,
    output [105:0] col_out_460,
    output [105:0] col_out_461,
    output [105:0] col_out_462,
    output [105:0] col_out_463,
    output [105:0] col_out_464,
    output [105:0] col_out_465,
    output [105:0] col_out_466,
    output [105:0] col_out_467,
    output [105:0] col_out_468,
    output [105:0] col_out_469,
    output [105:0] col_out_470,
    output [105:0] col_out_471,
    output [105:0] col_out_472,
    output [105:0] col_out_473,
    output [105:0] col_out_474,
    output [105:0] col_out_475,
    output [105:0] col_out_476,
    output [105:0] col_out_477,
    output [105:0] col_out_478,
    output [105:0] col_out_479,
    output [105:0] col_out_480,
    output [105:0] col_out_481,
    output [105:0] col_out_482,
    output [105:0] col_out_483,
    output [105:0] col_out_484,
    output [105:0] col_out_485,
    output [105:0] col_out_486,
    output [105:0] col_out_487,
    output [105:0] col_out_488,
    output [105:0] col_out_489,
    output [105:0] col_out_490,
    output [105:0] col_out_491,
    output [105:0] col_out_492,
    output [105:0] col_out_493,
    output [105:0] col_out_494,
    output [105:0] col_out_495,
    output [105:0] col_out_496,
    output [105:0] col_out_497,
    output [105:0] col_out_498,
    output [105:0] col_out_499,
    output [105:0] col_out_500,
    output [105:0] col_out_501,
    output [105:0] col_out_502,
    output [105:0] col_out_503,
    output [105:0] col_out_504,
    output [105:0] col_out_505,
    output [105:0] col_out_506,
    output [105:0] col_out_507,
    output [105:0] col_out_508,
    output [105:0] col_out_509,
    output [105:0] col_out_510,
    output [105:0] col_out_511,
    output [105:0] col_out_512,
    output [105:0] col_out_513,
    output [105:0] col_out_514,
    output [105:0] col_out_515,
    output [105:0] col_out_516,
    output [105:0] col_out_517,
    output [105:0] col_out_518,
    output [105:0] col_out_519,
    output [105:0] col_out_520,
    output [105:0] col_out_521,
    output [105:0] col_out_522,
    output [105:0] col_out_523,
    output [105:0] col_out_524,
    output [105:0] col_out_525,
    output [105:0] col_out_526,
    output [105:0] col_out_527,
    output [105:0] col_out_528,
    output [105:0] col_out_529,
    output [105:0] col_out_530,
    output [105:0] col_out_531,
    output [105:0] col_out_532,
    output [105:0] col_out_533,
    output [105:0] col_out_534,
    output [105:0] col_out_535,
    output [105:0] col_out_536,
    output [105:0] col_out_537,
    output [105:0] col_out_538,
    output [105:0] col_out_539,
    output [105:0] col_out_540,
    output [105:0] col_out_541,
    output [105:0] col_out_542,
    output [105:0] col_out_543,
    output [105:0] col_out_544,
    output [105:0] col_out_545,
    output [105:0] col_out_546,
    output [105:0] col_out_547,
    output [105:0] col_out_548,
    output [105:0] col_out_549,
    output [105:0] col_out_550,
    output [105:0] col_out_551,
    output [105:0] col_out_552,
    output [105:0] col_out_553,
    output [105:0] col_out_554,
    output [105:0] col_out_555,
    output [105:0] col_out_556,
    output [105:0] col_out_557,
    output [105:0] col_out_558,
    output [105:0] col_out_559,
    output [105:0] col_out_560,
    output [105:0] col_out_561,
    output [105:0] col_out_562,
    output [105:0] col_out_563,
    output [105:0] col_out_564,
    output [105:0] col_out_565,
    output [105:0] col_out_566,
    output [105:0] col_out_567,
    output [105:0] col_out_568,
    output [105:0] col_out_569,
    output [105:0] col_out_570,
    output [105:0] col_out_571,
    output [105:0] col_out_572,
    output [105:0] col_out_573,
    output [105:0] col_out_574,
    output [105:0] col_out_575,
    output [105:0] col_out_576,
    output [105:0] col_out_577,
    output [105:0] col_out_578,
    output [105:0] col_out_579,
    output [105:0] col_out_580,
    output [105:0] col_out_581,
    output [105:0] col_out_582,
    output [105:0] col_out_583,
    output [105:0] col_out_584,
    output [105:0] col_out_585,
    output [105:0] col_out_586,
    output [105:0] col_out_587,
    output [105:0] col_out_588,
    output [105:0] col_out_589,
    output [105:0] col_out_590,
    output [105:0] col_out_591,
    output [105:0] col_out_592,
    output [105:0] col_out_593,
    output [105:0] col_out_594,
    output [105:0] col_out_595,
    output [105:0] col_out_596,
    output [105:0] col_out_597,
    output [105:0] col_out_598,
    output [105:0] col_out_599,
    output [105:0] col_out_600,
    output [105:0] col_out_601,
    output [105:0] col_out_602,
    output [105:0] col_out_603,
    output [105:0] col_out_604,
    output [105:0] col_out_605,
    output [105:0] col_out_606,
    output [105:0] col_out_607,
    output [105:0] col_out_608,
    output [105:0] col_out_609,
    output [105:0] col_out_610,
    output [105:0] col_out_611,
    output [105:0] col_out_612,
    output [105:0] col_out_613,
    output [105:0] col_out_614,
    output [105:0] col_out_615,
    output [105:0] col_out_616,
    output [105:0] col_out_617,
    output [105:0] col_out_618,
    output [105:0] col_out_619,
    output [105:0] col_out_620,
    output [105:0] col_out_621,
    output [105:0] col_out_622,
    output [105:0] col_out_623,
    output [105:0] col_out_624,
    output [105:0] col_out_625,
    output [105:0] col_out_626,
    output [105:0] col_out_627,
    output [105:0] col_out_628,
    output [105:0] col_out_629,
    output [105:0] col_out_630,
    output [105:0] col_out_631,
    output [105:0] col_out_632,
    output [105:0] col_out_633,
    output [105:0] col_out_634,
    output [105:0] col_out_635,
    output [105:0] col_out_636,
    output [105:0] col_out_637,
    output [105:0] col_out_638,
    output [105:0] col_out_639,
    output [105:0] col_out_640,
    output [105:0] col_out_641,
    output [105:0] col_out_642,
    output [105:0] col_out_643,
    output [105:0] col_out_644,
    output [105:0] col_out_645,
    output [105:0] col_out_646,
    output [105:0] col_out_647,
    output [105:0] col_out_648,
    output [105:0] col_out_649,
    output [105:0] col_out_650,
    output [105:0] col_out_651,
    output [105:0] col_out_652,
    output [105:0] col_out_653,
    output [105:0] col_out_654,
    output [105:0] col_out_655,
    output [105:0] col_out_656,
    output [105:0] col_out_657,
    output [105:0] col_out_658,
    output [105:0] col_out_659,
    output [105:0] col_out_660,
    output [105:0] col_out_661,
    output [105:0] col_out_662,
    output [105:0] col_out_663,
    output [105:0] col_out_664,
    output [105:0] col_out_665,
    output [105:0] col_out_666,
    output [105:0] col_out_667,
    output [105:0] col_out_668,
    output [105:0] col_out_669,
    output [105:0] col_out_670,
    output [105:0] col_out_671,
    output [105:0] col_out_672,
    output [105:0] col_out_673,
    output [105:0] col_out_674,
    output [105:0] col_out_675,
    output [105:0] col_out_676,
    output [105:0] col_out_677,
    output [105:0] col_out_678,
    output [105:0] col_out_679,
    output [105:0] col_out_680,
    output [105:0] col_out_681,
    output [105:0] col_out_682,
    output [105:0] col_out_683,
    output [105:0] col_out_684,
    output [105:0] col_out_685,
    output [105:0] col_out_686,
    output [105:0] col_out_687,
    output [105:0] col_out_688,
    output [105:0] col_out_689,
    output [105:0] col_out_690,
    output [105:0] col_out_691,
    output [105:0] col_out_692,
    output [105:0] col_out_693,
    output [105:0] col_out_694,
    output [105:0] col_out_695,
    output [105:0] col_out_696,
    output [105:0] col_out_697,
    output [105:0] col_out_698,
    output [105:0] col_out_699,
    output [105:0] col_out_700,
    output [105:0] col_out_701,
    output [105:0] col_out_702,
    output [105:0] col_out_703,
    output [105:0] col_out_704,
    output [105:0] col_out_705,
    output [105:0] col_out_706,
    output [105:0] col_out_707,
    output [105:0] col_out_708,
    output [105:0] col_out_709,
    output [105:0] col_out_710,
    output [105:0] col_out_711,
    output [105:0] col_out_712,
    output [105:0] col_out_713,
    output [105:0] col_out_714,
    output [105:0] col_out_715,
    output [105:0] col_out_716,
    output [105:0] col_out_717,
    output [105:0] col_out_718,
    output [105:0] col_out_719,
    output [105:0] col_out_720,
    output [105:0] col_out_721,
    output [105:0] col_out_722,
    output [105:0] col_out_723,
    output [105:0] col_out_724,
    output [105:0] col_out_725,
    output [105:0] col_out_726,
    output [105:0] col_out_727,
    output [105:0] col_out_728,
    output [105:0] col_out_729,
    output [105:0] col_out_730,
    output [105:0] col_out_731,
    output [105:0] col_out_732,
    output [105:0] col_out_733,
    output [105:0] col_out_734,
    output [105:0] col_out_735,
    output [105:0] col_out_736,
    output [105:0] col_out_737,
    output [105:0] col_out_738,
    output [105:0] col_out_739,
    output [105:0] col_out_740,
    output [105:0] col_out_741,
    output [105:0] col_out_742,
    output [105:0] col_out_743,
    output [105:0] col_out_744,
    output [105:0] col_out_745,
    output [105:0] col_out_746,
    output [105:0] col_out_747,
    output [105:0] col_out_748,
    output [105:0] col_out_749,
    output [105:0] col_out_750,
    output [105:0] col_out_751,
    output [105:0] col_out_752,
    output [105:0] col_out_753,
    output [105:0] col_out_754,
    output [105:0] col_out_755,
    output [105:0] col_out_756,
    output [105:0] col_out_757,
    output [105:0] col_out_758,
    output [105:0] col_out_759,
    output [105:0] col_out_760,
    output [105:0] col_out_761,
    output [105:0] col_out_762,
    output [105:0] col_out_763,
    output [105:0] col_out_764,
    output [105:0] col_out_765,
    output [105:0] col_out_766,
    output [105:0] col_out_767,
    output [105:0] col_out_768,
    output [105:0] col_out_769,
    output [105:0] col_out_770,
    output [105:0] col_out_771,
    output [105:0] col_out_772,
    output [105:0] col_out_773,
    output [105:0] col_out_774,
    output [105:0] col_out_775,
    output [105:0] col_out_776,
    output [105:0] col_out_777,
    output [105:0] col_out_778,
    output [105:0] col_out_779,
    output [105:0] col_out_780,
    output [105:0] col_out_781,
    output [105:0] col_out_782,
    output [105:0] col_out_783,
    output [105:0] col_out_784,
    output [105:0] col_out_785,
    output [105:0] col_out_786,
    output [105:0] col_out_787,
    output [105:0] col_out_788,
    output [105:0] col_out_789,
    output [105:0] col_out_790,
    output [105:0] col_out_791,
    output [105:0] col_out_792,
    output [105:0] col_out_793,
    output [105:0] col_out_794,
    output [105:0] col_out_795,
    output [105:0] col_out_796,
    output [105:0] col_out_797,
    output [105:0] col_out_798,
    output [105:0] col_out_799,
    output [105:0] col_out_800,
    output [105:0] col_out_801,
    output [105:0] col_out_802,
    output [105:0] col_out_803,
    output [105:0] col_out_804,
    output [105:0] col_out_805,
    output [105:0] col_out_806,
    output [105:0] col_out_807,
    output [105:0] col_out_808,
    output [105:0] col_out_809,
    output [105:0] col_out_810,
    output [105:0] col_out_811,
    output [105:0] col_out_812,
    output [105:0] col_out_813,
    output [105:0] col_out_814,
    output [105:0] col_out_815,
    output [105:0] col_out_816,
    output [105:0] col_out_817,
    output [105:0] col_out_818,
    output [105:0] col_out_819,
    output [105:0] col_out_820,
    output [105:0] col_out_821,
    output [105:0] col_out_822,
    output [105:0] col_out_823,
    output [105:0] col_out_824,
    output [105:0] col_out_825,
    output [105:0] col_out_826,
    output [105:0] col_out_827,
    output [105:0] col_out_828,
    output [105:0] col_out_829,
    output [105:0] col_out_830,
    output [105:0] col_out_831,
    output [105:0] col_out_832,
    output [105:0] col_out_833,
    output [105:0] col_out_834,
    output [105:0] col_out_835,
    output [105:0] col_out_836,
    output [105:0] col_out_837,
    output [105:0] col_out_838,
    output [105:0] col_out_839,
    output [105:0] col_out_840,
    output [105:0] col_out_841,
    output [105:0] col_out_842,
    output [105:0] col_out_843,
    output [105:0] col_out_844,
    output [105:0] col_out_845,
    output [105:0] col_out_846,
    output [105:0] col_out_847,
    output [105:0] col_out_848,
    output [105:0] col_out_849,
    output [105:0] col_out_850,
    output [105:0] col_out_851,
    output [105:0] col_out_852,
    output [105:0] col_out_853,
    output [105:0] col_out_854,
    output [105:0] col_out_855,
    output [105:0] col_out_856,
    output [105:0] col_out_857,
    output [105:0] col_out_858,
    output [105:0] col_out_859,
    output [105:0] col_out_860,
    output [105:0] col_out_861,
    output [105:0] col_out_862,
    output [105:0] col_out_863,
    output [105:0] col_out_864,
    output [105:0] col_out_865,
    output [105:0] col_out_866,
    output [105:0] col_out_867,
    output [105:0] col_out_868,
    output [105:0] col_out_869,
    output [105:0] col_out_870,
    output [105:0] col_out_871,
    output [105:0] col_out_872,
    output [105:0] col_out_873,
    output [105:0] col_out_874,
    output [105:0] col_out_875,
    output [105:0] col_out_876,
    output [105:0] col_out_877,
    output [105:0] col_out_878,
    output [105:0] col_out_879,
    output [105:0] col_out_880,
    output [105:0] col_out_881,
    output [105:0] col_out_882,
    output [105:0] col_out_883,
    output [105:0] col_out_884,
    output [105:0] col_out_885,
    output [105:0] col_out_886,
    output [105:0] col_out_887,
    output [105:0] col_out_888,
    output [105:0] col_out_889,
    output [105:0] col_out_890,
    output [105:0] col_out_891,
    output [105:0] col_out_892,
    output [105:0] col_out_893,
    output [105:0] col_out_894,
    output [105:0] col_out_895,
    output [105:0] col_out_896,
    output [105:0] col_out_897,
    output [105:0] col_out_898,
    output [105:0] col_out_899,
    output [105:0] col_out_900,
    output [105:0] col_out_901,
    output [105:0] col_out_902,
    output [105:0] col_out_903,
    output [105:0] col_out_904,
    output [105:0] col_out_905,
    output [105:0] col_out_906,
    output [105:0] col_out_907,
    output [105:0] col_out_908,
    output [105:0] col_out_909,
    output [105:0] col_out_910,
    output [105:0] col_out_911,
    output [105:0] col_out_912,
    output [105:0] col_out_913,
    output [105:0] col_out_914,
    output [105:0] col_out_915,
    output [105:0] col_out_916,
    output [105:0] col_out_917,
    output [105:0] col_out_918,
    output [105:0] col_out_919,
    output [105:0] col_out_920,
    output [105:0] col_out_921,
    output [105:0] col_out_922,
    output [105:0] col_out_923,
    output [105:0] col_out_924,
    output [105:0] col_out_925,
    output [105:0] col_out_926,
    output [105:0] col_out_927,
    output [105:0] col_out_928,
    output [105:0] col_out_929,
    output [105:0] col_out_930,
    output [105:0] col_out_931,
    output [105:0] col_out_932,
    output [105:0] col_out_933,
    output [105:0] col_out_934,
    output [105:0] col_out_935,
    output [105:0] col_out_936,
    output [105:0] col_out_937,
    output [105:0] col_out_938,
    output [105:0] col_out_939,
    output [105:0] col_out_940,
    output [105:0] col_out_941,
    output [105:0] col_out_942,
    output [105:0] col_out_943,
    output [105:0] col_out_944,
    output [105:0] col_out_945,
    output [105:0] col_out_946,
    output [105:0] col_out_947,
    output [105:0] col_out_948,
    output [105:0] col_out_949,
    output [105:0] col_out_950,
    output [105:0] col_out_951,
    output [105:0] col_out_952,
    output [105:0] col_out_953,
    output [105:0] col_out_954,
    output [105:0] col_out_955,
    output [105:0] col_out_956,
    output [105:0] col_out_957,
    output [105:0] col_out_958,
    output [105:0] col_out_959,
    output [105:0] col_out_960,
    output [105:0] col_out_961,
    output [105:0] col_out_962,
    output [105:0] col_out_963,
    output [105:0] col_out_964,
    output [105:0] col_out_965,
    output [105:0] col_out_966,
    output [105:0] col_out_967,
    output [105:0] col_out_968,
    output [105:0] col_out_969,
    output [105:0] col_out_970,
    output [105:0] col_out_971,
    output [105:0] col_out_972,
    output [105:0] col_out_973,
    output [105:0] col_out_974,
    output [105:0] col_out_975,
    output [105:0] col_out_976,
    output [105:0] col_out_977,
    output [105:0] col_out_978,
    output [105:0] col_out_979,
    output [105:0] col_out_980,
    output [105:0] col_out_981,
    output [105:0] col_out_982,
    output [105:0] col_out_983,
    output [105:0] col_out_984,
    output [105:0] col_out_985,
    output [105:0] col_out_986,
    output [105:0] col_out_987,
    output [105:0] col_out_988,
    output [105:0] col_out_989,
    output [105:0] col_out_990,
    output [105:0] col_out_991,
    output [105:0] col_out_992,
    output [105:0] col_out_993,
    output [105:0] col_out_994,
    output [105:0] col_out_995,
    output [105:0] col_out_996,
    output [105:0] col_out_997,
    output [105:0] col_out_998,
    output [105:0] col_out_999,
    output [105:0] col_out_1000,
    output [105:0] col_out_1001,
    output [105:0] col_out_1002,
    output [105:0] col_out_1003,
    output [105:0] col_out_1004,
    output [105:0] col_out_1005,
    output [105:0] col_out_1006,
    output [105:0] col_out_1007,
    output [105:0] col_out_1008,
    output [105:0] col_out_1009,
    output [105:0] col_out_1010,
    output [105:0] col_out_1011,
    output [105:0] col_out_1012,
    output [105:0] col_out_1013,
    output [105:0] col_out_1014,
    output [105:0] col_out_1015,
    output [105:0] col_out_1016,
    output [105:0] col_out_1017,
    output [105:0] col_out_1018,
    output [105:0] col_out_1019,
    output [105:0] col_out_1020,
    output [105:0] col_out_1021,
    output [105:0] col_out_1022,
    output [105:0] col_out_1023
);


wire [1023:0] u_xpb_out[105:0];



xpb_264 u0_xpb_4_260(
    .data_in(data_in0), 

    .data_out_0(u_xpb_out[0]),
    .data_out_1(u_xpb_out[1]),
    .data_out_2(u_xpb_out[2]),
    .data_out_3(u_xpb_out[3]),
    .data_out_4(u_xpb_out[4]),
    .data_out_5(u_xpb_out[5]),
    .data_out_6(u_xpb_out[6]),
    .data_out_7(u_xpb_out[7]),
    .data_out_8(u_xpb_out[8]),
    .data_out_9(u_xpb_out[9]),
    .data_out_10(u_xpb_out[10]),
    .data_out_11(u_xpb_out[11]),
    .data_out_12(u_xpb_out[12]),
    .data_out_13(u_xpb_out[13]),
    .data_out_14(u_xpb_out[14]),
    .data_out_15(u_xpb_out[15]),
    .data_out_16(u_xpb_out[16]),
    .data_out_17(u_xpb_out[17]),
    .data_out_18(u_xpb_out[18]),
    .data_out_19(u_xpb_out[19]),
    .data_out_20(u_xpb_out[20]),
    .data_out_21(u_xpb_out[21]),
    .data_out_22(u_xpb_out[22]),
    .data_out_23(u_xpb_out[23]),
    .data_out_24(u_xpb_out[24]),
    .data_out_25(u_xpb_out[25]),
    .data_out_26(u_xpb_out[26]),
    .data_out_27(u_xpb_out[27]),
    .data_out_28(u_xpb_out[28]),
    .data_out_29(u_xpb_out[29]),
    .data_out_30(u_xpb_out[30]),
    .data_out_31(u_xpb_out[31]),
    .data_out_32(u_xpb_out[32]),
    .data_out_33(u_xpb_out[33]),
    .data_out_34(u_xpb_out[34]),
    .data_out_35(u_xpb_out[35]),
    .data_out_36(u_xpb_out[36]),
    .data_out_37(u_xpb_out[37]),
    .data_out_38(u_xpb_out[38]),
    .data_out_39(u_xpb_out[39]),
    .data_out_40(u_xpb_out[40]),
    .data_out_41(u_xpb_out[41]),
    .data_out_42(u_xpb_out[42]),
    .data_out_43(u_xpb_out[43]),
    .data_out_44(u_xpb_out[44]),
    .data_out_45(u_xpb_out[45]),
    .data_out_46(u_xpb_out[46]),
    .data_out_47(u_xpb_out[47]),
    .data_out_48(u_xpb_out[48]),
    .data_out_49(u_xpb_out[49]),
    .data_out_50(u_xpb_out[50]),
    .data_out_51(u_xpb_out[51]),
    .data_out_52(u_xpb_out[52])
);


xpb_264 u1_xpb_4_260(
    .data_in(data_in1), 

    .data_out_0(u_xpb_out[53]),
    .data_out_1(u_xpb_out[54]),
    .data_out_2(u_xpb_out[55]),
    .data_out_3(u_xpb_out[56]),
    .data_out_4(u_xpb_out[57]),
    .data_out_5(u_xpb_out[58]),
    .data_out_6(u_xpb_out[59]),
    .data_out_7(u_xpb_out[60]),
    .data_out_8(u_xpb_out[61]),
    .data_out_9(u_xpb_out[62]),
    .data_out_10(u_xpb_out[63]),
    .data_out_11(u_xpb_out[64]),
    .data_out_12(u_xpb_out[65]),
    .data_out_13(u_xpb_out[66]),
    .data_out_14(u_xpb_out[67]),
    .data_out_15(u_xpb_out[68]),
    .data_out_16(u_xpb_out[69]),
    .data_out_17(u_xpb_out[70]),
    .data_out_18(u_xpb_out[71]),
    .data_out_19(u_xpb_out[72]),
    .data_out_20(u_xpb_out[73]),
    .data_out_21(u_xpb_out[74]),
    .data_out_22(u_xpb_out[75]),
    .data_out_23(u_xpb_out[76]),
    .data_out_24(u_xpb_out[77]),
    .data_out_25(u_xpb_out[78]),
    .data_out_26(u_xpb_out[79]),
    .data_out_27(u_xpb_out[80]),
    .data_out_28(u_xpb_out[81]),
    .data_out_29(u_xpb_out[82]),
    .data_out_30(u_xpb_out[83]),
    .data_out_31(u_xpb_out[84]),
    .data_out_32(u_xpb_out[85]),
    .data_out_33(u_xpb_out[86]),
    .data_out_34(u_xpb_out[87]),
    .data_out_35(u_xpb_out[88]),
    .data_out_36(u_xpb_out[89]),
    .data_out_37(u_xpb_out[90]),
    .data_out_38(u_xpb_out[91]),
    .data_out_39(u_xpb_out[92]),
    .data_out_40(u_xpb_out[93]),
    .data_out_41(u_xpb_out[94]),
    .data_out_42(u_xpb_out[95]),
    .data_out_43(u_xpb_out[96]),
    .data_out_44(u_xpb_out[97]),
    .data_out_45(u_xpb_out[98]),
    .data_out_46(u_xpb_out[99]),
    .data_out_47(u_xpb_out[100]),
    .data_out_48(u_xpb_out[101]),
    .data_out_49(u_xpb_out[102]),
    .data_out_50(u_xpb_out[103]),
    .data_out_51(u_xpb_out[104]),
    .data_out_52(u_xpb_out[105])
);


assign col_out_0 = {u_xpb_out[0][0],u_xpb_out[1][0],u_xpb_out[2][0],u_xpb_out[3][0],u_xpb_out[4][0],u_xpb_out[5][0],u_xpb_out[6][0],u_xpb_out[7][0],u_xpb_out[8][0],u_xpb_out[9][0],u_xpb_out[10][0],u_xpb_out[11][0],u_xpb_out[12][0],u_xpb_out[13][0],u_xpb_out[14][0],u_xpb_out[15][0],u_xpb_out[16][0],u_xpb_out[17][0],u_xpb_out[18][0],u_xpb_out[19][0],u_xpb_out[20][0],u_xpb_out[21][0],u_xpb_out[22][0],u_xpb_out[23][0],u_xpb_out[24][0],u_xpb_out[25][0],u_xpb_out[26][0],u_xpb_out[27][0],u_xpb_out[28][0],u_xpb_out[29][0],u_xpb_out[30][0],u_xpb_out[31][0],u_xpb_out[32][0],u_xpb_out[33][0],u_xpb_out[34][0],u_xpb_out[35][0],u_xpb_out[36][0],u_xpb_out[37][0],u_xpb_out[38][0],u_xpb_out[39][0],u_xpb_out[40][0],u_xpb_out[41][0],u_xpb_out[42][0],u_xpb_out[43][0],u_xpb_out[44][0],u_xpb_out[45][0],u_xpb_out[46][0],u_xpb_out[47][0],u_xpb_out[48][0],u_xpb_out[49][0],u_xpb_out[50][0],u_xpb_out[51][0],u_xpb_out[52][0],u_xpb_out[53][0],u_xpb_out[54][0],u_xpb_out[55][0],u_xpb_out[56][0],u_xpb_out[57][0],u_xpb_out[58][0],u_xpb_out[59][0],u_xpb_out[60][0],u_xpb_out[61][0],u_xpb_out[62][0],u_xpb_out[63][0],u_xpb_out[64][0],u_xpb_out[65][0],u_xpb_out[66][0],u_xpb_out[67][0],u_xpb_out[68][0],u_xpb_out[69][0],u_xpb_out[70][0],u_xpb_out[71][0],u_xpb_out[72][0],u_xpb_out[73][0],u_xpb_out[74][0],u_xpb_out[75][0],u_xpb_out[76][0],u_xpb_out[77][0],u_xpb_out[78][0],u_xpb_out[79][0],u_xpb_out[80][0],u_xpb_out[81][0],u_xpb_out[82][0],u_xpb_out[83][0],u_xpb_out[84][0],u_xpb_out[85][0],u_xpb_out[86][0],u_xpb_out[87][0],u_xpb_out[88][0],u_xpb_out[89][0],u_xpb_out[90][0],u_xpb_out[91][0],u_xpb_out[92][0],u_xpb_out[93][0],u_xpb_out[94][0],u_xpb_out[95][0],u_xpb_out[96][0],u_xpb_out[97][0],u_xpb_out[98][0],u_xpb_out[99][0],u_xpb_out[100][0],u_xpb_out[101][0],u_xpb_out[102][0],u_xpb_out[103][0],u_xpb_out[104][0],u_xpb_out[105][0]};

assign col_out_1 = {u_xpb_out[0][1],u_xpb_out[1][1],u_xpb_out[2][1],u_xpb_out[3][1],u_xpb_out[4][1],u_xpb_out[5][1],u_xpb_out[6][1],u_xpb_out[7][1],u_xpb_out[8][1],u_xpb_out[9][1],u_xpb_out[10][1],u_xpb_out[11][1],u_xpb_out[12][1],u_xpb_out[13][1],u_xpb_out[14][1],u_xpb_out[15][1],u_xpb_out[16][1],u_xpb_out[17][1],u_xpb_out[18][1],u_xpb_out[19][1],u_xpb_out[20][1],u_xpb_out[21][1],u_xpb_out[22][1],u_xpb_out[23][1],u_xpb_out[24][1],u_xpb_out[25][1],u_xpb_out[26][1],u_xpb_out[27][1],u_xpb_out[28][1],u_xpb_out[29][1],u_xpb_out[30][1],u_xpb_out[31][1],u_xpb_out[32][1],u_xpb_out[33][1],u_xpb_out[34][1],u_xpb_out[35][1],u_xpb_out[36][1],u_xpb_out[37][1],u_xpb_out[38][1],u_xpb_out[39][1],u_xpb_out[40][1],u_xpb_out[41][1],u_xpb_out[42][1],u_xpb_out[43][1],u_xpb_out[44][1],u_xpb_out[45][1],u_xpb_out[46][1],u_xpb_out[47][1],u_xpb_out[48][1],u_xpb_out[49][1],u_xpb_out[50][1],u_xpb_out[51][1],u_xpb_out[52][1],u_xpb_out[53][1],u_xpb_out[54][1],u_xpb_out[55][1],u_xpb_out[56][1],u_xpb_out[57][1],u_xpb_out[58][1],u_xpb_out[59][1],u_xpb_out[60][1],u_xpb_out[61][1],u_xpb_out[62][1],u_xpb_out[63][1],u_xpb_out[64][1],u_xpb_out[65][1],u_xpb_out[66][1],u_xpb_out[67][1],u_xpb_out[68][1],u_xpb_out[69][1],u_xpb_out[70][1],u_xpb_out[71][1],u_xpb_out[72][1],u_xpb_out[73][1],u_xpb_out[74][1],u_xpb_out[75][1],u_xpb_out[76][1],u_xpb_out[77][1],u_xpb_out[78][1],u_xpb_out[79][1],u_xpb_out[80][1],u_xpb_out[81][1],u_xpb_out[82][1],u_xpb_out[83][1],u_xpb_out[84][1],u_xpb_out[85][1],u_xpb_out[86][1],u_xpb_out[87][1],u_xpb_out[88][1],u_xpb_out[89][1],u_xpb_out[90][1],u_xpb_out[91][1],u_xpb_out[92][1],u_xpb_out[93][1],u_xpb_out[94][1],u_xpb_out[95][1],u_xpb_out[96][1],u_xpb_out[97][1],u_xpb_out[98][1],u_xpb_out[99][1],u_xpb_out[100][1],u_xpb_out[101][1],u_xpb_out[102][1],u_xpb_out[103][1],u_xpb_out[104][1],u_xpb_out[105][1]};

assign col_out_2 = {u_xpb_out[0][2],u_xpb_out[1][2],u_xpb_out[2][2],u_xpb_out[3][2],u_xpb_out[4][2],u_xpb_out[5][2],u_xpb_out[6][2],u_xpb_out[7][2],u_xpb_out[8][2],u_xpb_out[9][2],u_xpb_out[10][2],u_xpb_out[11][2],u_xpb_out[12][2],u_xpb_out[13][2],u_xpb_out[14][2],u_xpb_out[15][2],u_xpb_out[16][2],u_xpb_out[17][2],u_xpb_out[18][2],u_xpb_out[19][2],u_xpb_out[20][2],u_xpb_out[21][2],u_xpb_out[22][2],u_xpb_out[23][2],u_xpb_out[24][2],u_xpb_out[25][2],u_xpb_out[26][2],u_xpb_out[27][2],u_xpb_out[28][2],u_xpb_out[29][2],u_xpb_out[30][2],u_xpb_out[31][2],u_xpb_out[32][2],u_xpb_out[33][2],u_xpb_out[34][2],u_xpb_out[35][2],u_xpb_out[36][2],u_xpb_out[37][2],u_xpb_out[38][2],u_xpb_out[39][2],u_xpb_out[40][2],u_xpb_out[41][2],u_xpb_out[42][2],u_xpb_out[43][2],u_xpb_out[44][2],u_xpb_out[45][2],u_xpb_out[46][2],u_xpb_out[47][2],u_xpb_out[48][2],u_xpb_out[49][2],u_xpb_out[50][2],u_xpb_out[51][2],u_xpb_out[52][2],u_xpb_out[53][2],u_xpb_out[54][2],u_xpb_out[55][2],u_xpb_out[56][2],u_xpb_out[57][2],u_xpb_out[58][2],u_xpb_out[59][2],u_xpb_out[60][2],u_xpb_out[61][2],u_xpb_out[62][2],u_xpb_out[63][2],u_xpb_out[64][2],u_xpb_out[65][2],u_xpb_out[66][2],u_xpb_out[67][2],u_xpb_out[68][2],u_xpb_out[69][2],u_xpb_out[70][2],u_xpb_out[71][2],u_xpb_out[72][2],u_xpb_out[73][2],u_xpb_out[74][2],u_xpb_out[75][2],u_xpb_out[76][2],u_xpb_out[77][2],u_xpb_out[78][2],u_xpb_out[79][2],u_xpb_out[80][2],u_xpb_out[81][2],u_xpb_out[82][2],u_xpb_out[83][2],u_xpb_out[84][2],u_xpb_out[85][2],u_xpb_out[86][2],u_xpb_out[87][2],u_xpb_out[88][2],u_xpb_out[89][2],u_xpb_out[90][2],u_xpb_out[91][2],u_xpb_out[92][2],u_xpb_out[93][2],u_xpb_out[94][2],u_xpb_out[95][2],u_xpb_out[96][2],u_xpb_out[97][2],u_xpb_out[98][2],u_xpb_out[99][2],u_xpb_out[100][2],u_xpb_out[101][2],u_xpb_out[102][2],u_xpb_out[103][2],u_xpb_out[104][2],u_xpb_out[105][2]};

assign col_out_3 = {u_xpb_out[0][3],u_xpb_out[1][3],u_xpb_out[2][3],u_xpb_out[3][3],u_xpb_out[4][3],u_xpb_out[5][3],u_xpb_out[6][3],u_xpb_out[7][3],u_xpb_out[8][3],u_xpb_out[9][3],u_xpb_out[10][3],u_xpb_out[11][3],u_xpb_out[12][3],u_xpb_out[13][3],u_xpb_out[14][3],u_xpb_out[15][3],u_xpb_out[16][3],u_xpb_out[17][3],u_xpb_out[18][3],u_xpb_out[19][3],u_xpb_out[20][3],u_xpb_out[21][3],u_xpb_out[22][3],u_xpb_out[23][3],u_xpb_out[24][3],u_xpb_out[25][3],u_xpb_out[26][3],u_xpb_out[27][3],u_xpb_out[28][3],u_xpb_out[29][3],u_xpb_out[30][3],u_xpb_out[31][3],u_xpb_out[32][3],u_xpb_out[33][3],u_xpb_out[34][3],u_xpb_out[35][3],u_xpb_out[36][3],u_xpb_out[37][3],u_xpb_out[38][3],u_xpb_out[39][3],u_xpb_out[40][3],u_xpb_out[41][3],u_xpb_out[42][3],u_xpb_out[43][3],u_xpb_out[44][3],u_xpb_out[45][3],u_xpb_out[46][3],u_xpb_out[47][3],u_xpb_out[48][3],u_xpb_out[49][3],u_xpb_out[50][3],u_xpb_out[51][3],u_xpb_out[52][3],u_xpb_out[53][3],u_xpb_out[54][3],u_xpb_out[55][3],u_xpb_out[56][3],u_xpb_out[57][3],u_xpb_out[58][3],u_xpb_out[59][3],u_xpb_out[60][3],u_xpb_out[61][3],u_xpb_out[62][3],u_xpb_out[63][3],u_xpb_out[64][3],u_xpb_out[65][3],u_xpb_out[66][3],u_xpb_out[67][3],u_xpb_out[68][3],u_xpb_out[69][3],u_xpb_out[70][3],u_xpb_out[71][3],u_xpb_out[72][3],u_xpb_out[73][3],u_xpb_out[74][3],u_xpb_out[75][3],u_xpb_out[76][3],u_xpb_out[77][3],u_xpb_out[78][3],u_xpb_out[79][3],u_xpb_out[80][3],u_xpb_out[81][3],u_xpb_out[82][3],u_xpb_out[83][3],u_xpb_out[84][3],u_xpb_out[85][3],u_xpb_out[86][3],u_xpb_out[87][3],u_xpb_out[88][3],u_xpb_out[89][3],u_xpb_out[90][3],u_xpb_out[91][3],u_xpb_out[92][3],u_xpb_out[93][3],u_xpb_out[94][3],u_xpb_out[95][3],u_xpb_out[96][3],u_xpb_out[97][3],u_xpb_out[98][3],u_xpb_out[99][3],u_xpb_out[100][3],u_xpb_out[101][3],u_xpb_out[102][3],u_xpb_out[103][3],u_xpb_out[104][3],u_xpb_out[105][3]};

assign col_out_4 = {u_xpb_out[0][4],u_xpb_out[1][4],u_xpb_out[2][4],u_xpb_out[3][4],u_xpb_out[4][4],u_xpb_out[5][4],u_xpb_out[6][4],u_xpb_out[7][4],u_xpb_out[8][4],u_xpb_out[9][4],u_xpb_out[10][4],u_xpb_out[11][4],u_xpb_out[12][4],u_xpb_out[13][4],u_xpb_out[14][4],u_xpb_out[15][4],u_xpb_out[16][4],u_xpb_out[17][4],u_xpb_out[18][4],u_xpb_out[19][4],u_xpb_out[20][4],u_xpb_out[21][4],u_xpb_out[22][4],u_xpb_out[23][4],u_xpb_out[24][4],u_xpb_out[25][4],u_xpb_out[26][4],u_xpb_out[27][4],u_xpb_out[28][4],u_xpb_out[29][4],u_xpb_out[30][4],u_xpb_out[31][4],u_xpb_out[32][4],u_xpb_out[33][4],u_xpb_out[34][4],u_xpb_out[35][4],u_xpb_out[36][4],u_xpb_out[37][4],u_xpb_out[38][4],u_xpb_out[39][4],u_xpb_out[40][4],u_xpb_out[41][4],u_xpb_out[42][4],u_xpb_out[43][4],u_xpb_out[44][4],u_xpb_out[45][4],u_xpb_out[46][4],u_xpb_out[47][4],u_xpb_out[48][4],u_xpb_out[49][4],u_xpb_out[50][4],u_xpb_out[51][4],u_xpb_out[52][4],u_xpb_out[53][4],u_xpb_out[54][4],u_xpb_out[55][4],u_xpb_out[56][4],u_xpb_out[57][4],u_xpb_out[58][4],u_xpb_out[59][4],u_xpb_out[60][4],u_xpb_out[61][4],u_xpb_out[62][4],u_xpb_out[63][4],u_xpb_out[64][4],u_xpb_out[65][4],u_xpb_out[66][4],u_xpb_out[67][4],u_xpb_out[68][4],u_xpb_out[69][4],u_xpb_out[70][4],u_xpb_out[71][4],u_xpb_out[72][4],u_xpb_out[73][4],u_xpb_out[74][4],u_xpb_out[75][4],u_xpb_out[76][4],u_xpb_out[77][4],u_xpb_out[78][4],u_xpb_out[79][4],u_xpb_out[80][4],u_xpb_out[81][4],u_xpb_out[82][4],u_xpb_out[83][4],u_xpb_out[84][4],u_xpb_out[85][4],u_xpb_out[86][4],u_xpb_out[87][4],u_xpb_out[88][4],u_xpb_out[89][4],u_xpb_out[90][4],u_xpb_out[91][4],u_xpb_out[92][4],u_xpb_out[93][4],u_xpb_out[94][4],u_xpb_out[95][4],u_xpb_out[96][4],u_xpb_out[97][4],u_xpb_out[98][4],u_xpb_out[99][4],u_xpb_out[100][4],u_xpb_out[101][4],u_xpb_out[102][4],u_xpb_out[103][4],u_xpb_out[104][4],u_xpb_out[105][4]};

assign col_out_5 = {u_xpb_out[0][5],u_xpb_out[1][5],u_xpb_out[2][5],u_xpb_out[3][5],u_xpb_out[4][5],u_xpb_out[5][5],u_xpb_out[6][5],u_xpb_out[7][5],u_xpb_out[8][5],u_xpb_out[9][5],u_xpb_out[10][5],u_xpb_out[11][5],u_xpb_out[12][5],u_xpb_out[13][5],u_xpb_out[14][5],u_xpb_out[15][5],u_xpb_out[16][5],u_xpb_out[17][5],u_xpb_out[18][5],u_xpb_out[19][5],u_xpb_out[20][5],u_xpb_out[21][5],u_xpb_out[22][5],u_xpb_out[23][5],u_xpb_out[24][5],u_xpb_out[25][5],u_xpb_out[26][5],u_xpb_out[27][5],u_xpb_out[28][5],u_xpb_out[29][5],u_xpb_out[30][5],u_xpb_out[31][5],u_xpb_out[32][5],u_xpb_out[33][5],u_xpb_out[34][5],u_xpb_out[35][5],u_xpb_out[36][5],u_xpb_out[37][5],u_xpb_out[38][5],u_xpb_out[39][5],u_xpb_out[40][5],u_xpb_out[41][5],u_xpb_out[42][5],u_xpb_out[43][5],u_xpb_out[44][5],u_xpb_out[45][5],u_xpb_out[46][5],u_xpb_out[47][5],u_xpb_out[48][5],u_xpb_out[49][5],u_xpb_out[50][5],u_xpb_out[51][5],u_xpb_out[52][5],u_xpb_out[53][5],u_xpb_out[54][5],u_xpb_out[55][5],u_xpb_out[56][5],u_xpb_out[57][5],u_xpb_out[58][5],u_xpb_out[59][5],u_xpb_out[60][5],u_xpb_out[61][5],u_xpb_out[62][5],u_xpb_out[63][5],u_xpb_out[64][5],u_xpb_out[65][5],u_xpb_out[66][5],u_xpb_out[67][5],u_xpb_out[68][5],u_xpb_out[69][5],u_xpb_out[70][5],u_xpb_out[71][5],u_xpb_out[72][5],u_xpb_out[73][5],u_xpb_out[74][5],u_xpb_out[75][5],u_xpb_out[76][5],u_xpb_out[77][5],u_xpb_out[78][5],u_xpb_out[79][5],u_xpb_out[80][5],u_xpb_out[81][5],u_xpb_out[82][5],u_xpb_out[83][5],u_xpb_out[84][5],u_xpb_out[85][5],u_xpb_out[86][5],u_xpb_out[87][5],u_xpb_out[88][5],u_xpb_out[89][5],u_xpb_out[90][5],u_xpb_out[91][5],u_xpb_out[92][5],u_xpb_out[93][5],u_xpb_out[94][5],u_xpb_out[95][5],u_xpb_out[96][5],u_xpb_out[97][5],u_xpb_out[98][5],u_xpb_out[99][5],u_xpb_out[100][5],u_xpb_out[101][5],u_xpb_out[102][5],u_xpb_out[103][5],u_xpb_out[104][5],u_xpb_out[105][5]};

assign col_out_6 = {u_xpb_out[0][6],u_xpb_out[1][6],u_xpb_out[2][6],u_xpb_out[3][6],u_xpb_out[4][6],u_xpb_out[5][6],u_xpb_out[6][6],u_xpb_out[7][6],u_xpb_out[8][6],u_xpb_out[9][6],u_xpb_out[10][6],u_xpb_out[11][6],u_xpb_out[12][6],u_xpb_out[13][6],u_xpb_out[14][6],u_xpb_out[15][6],u_xpb_out[16][6],u_xpb_out[17][6],u_xpb_out[18][6],u_xpb_out[19][6],u_xpb_out[20][6],u_xpb_out[21][6],u_xpb_out[22][6],u_xpb_out[23][6],u_xpb_out[24][6],u_xpb_out[25][6],u_xpb_out[26][6],u_xpb_out[27][6],u_xpb_out[28][6],u_xpb_out[29][6],u_xpb_out[30][6],u_xpb_out[31][6],u_xpb_out[32][6],u_xpb_out[33][6],u_xpb_out[34][6],u_xpb_out[35][6],u_xpb_out[36][6],u_xpb_out[37][6],u_xpb_out[38][6],u_xpb_out[39][6],u_xpb_out[40][6],u_xpb_out[41][6],u_xpb_out[42][6],u_xpb_out[43][6],u_xpb_out[44][6],u_xpb_out[45][6],u_xpb_out[46][6],u_xpb_out[47][6],u_xpb_out[48][6],u_xpb_out[49][6],u_xpb_out[50][6],u_xpb_out[51][6],u_xpb_out[52][6],u_xpb_out[53][6],u_xpb_out[54][6],u_xpb_out[55][6],u_xpb_out[56][6],u_xpb_out[57][6],u_xpb_out[58][6],u_xpb_out[59][6],u_xpb_out[60][6],u_xpb_out[61][6],u_xpb_out[62][6],u_xpb_out[63][6],u_xpb_out[64][6],u_xpb_out[65][6],u_xpb_out[66][6],u_xpb_out[67][6],u_xpb_out[68][6],u_xpb_out[69][6],u_xpb_out[70][6],u_xpb_out[71][6],u_xpb_out[72][6],u_xpb_out[73][6],u_xpb_out[74][6],u_xpb_out[75][6],u_xpb_out[76][6],u_xpb_out[77][6],u_xpb_out[78][6],u_xpb_out[79][6],u_xpb_out[80][6],u_xpb_out[81][6],u_xpb_out[82][6],u_xpb_out[83][6],u_xpb_out[84][6],u_xpb_out[85][6],u_xpb_out[86][6],u_xpb_out[87][6],u_xpb_out[88][6],u_xpb_out[89][6],u_xpb_out[90][6],u_xpb_out[91][6],u_xpb_out[92][6],u_xpb_out[93][6],u_xpb_out[94][6],u_xpb_out[95][6],u_xpb_out[96][6],u_xpb_out[97][6],u_xpb_out[98][6],u_xpb_out[99][6],u_xpb_out[100][6],u_xpb_out[101][6],u_xpb_out[102][6],u_xpb_out[103][6],u_xpb_out[104][6],u_xpb_out[105][6]};

assign col_out_7 = {u_xpb_out[0][7],u_xpb_out[1][7],u_xpb_out[2][7],u_xpb_out[3][7],u_xpb_out[4][7],u_xpb_out[5][7],u_xpb_out[6][7],u_xpb_out[7][7],u_xpb_out[8][7],u_xpb_out[9][7],u_xpb_out[10][7],u_xpb_out[11][7],u_xpb_out[12][7],u_xpb_out[13][7],u_xpb_out[14][7],u_xpb_out[15][7],u_xpb_out[16][7],u_xpb_out[17][7],u_xpb_out[18][7],u_xpb_out[19][7],u_xpb_out[20][7],u_xpb_out[21][7],u_xpb_out[22][7],u_xpb_out[23][7],u_xpb_out[24][7],u_xpb_out[25][7],u_xpb_out[26][7],u_xpb_out[27][7],u_xpb_out[28][7],u_xpb_out[29][7],u_xpb_out[30][7],u_xpb_out[31][7],u_xpb_out[32][7],u_xpb_out[33][7],u_xpb_out[34][7],u_xpb_out[35][7],u_xpb_out[36][7],u_xpb_out[37][7],u_xpb_out[38][7],u_xpb_out[39][7],u_xpb_out[40][7],u_xpb_out[41][7],u_xpb_out[42][7],u_xpb_out[43][7],u_xpb_out[44][7],u_xpb_out[45][7],u_xpb_out[46][7],u_xpb_out[47][7],u_xpb_out[48][7],u_xpb_out[49][7],u_xpb_out[50][7],u_xpb_out[51][7],u_xpb_out[52][7],u_xpb_out[53][7],u_xpb_out[54][7],u_xpb_out[55][7],u_xpb_out[56][7],u_xpb_out[57][7],u_xpb_out[58][7],u_xpb_out[59][7],u_xpb_out[60][7],u_xpb_out[61][7],u_xpb_out[62][7],u_xpb_out[63][7],u_xpb_out[64][7],u_xpb_out[65][7],u_xpb_out[66][7],u_xpb_out[67][7],u_xpb_out[68][7],u_xpb_out[69][7],u_xpb_out[70][7],u_xpb_out[71][7],u_xpb_out[72][7],u_xpb_out[73][7],u_xpb_out[74][7],u_xpb_out[75][7],u_xpb_out[76][7],u_xpb_out[77][7],u_xpb_out[78][7],u_xpb_out[79][7],u_xpb_out[80][7],u_xpb_out[81][7],u_xpb_out[82][7],u_xpb_out[83][7],u_xpb_out[84][7],u_xpb_out[85][7],u_xpb_out[86][7],u_xpb_out[87][7],u_xpb_out[88][7],u_xpb_out[89][7],u_xpb_out[90][7],u_xpb_out[91][7],u_xpb_out[92][7],u_xpb_out[93][7],u_xpb_out[94][7],u_xpb_out[95][7],u_xpb_out[96][7],u_xpb_out[97][7],u_xpb_out[98][7],u_xpb_out[99][7],u_xpb_out[100][7],u_xpb_out[101][7],u_xpb_out[102][7],u_xpb_out[103][7],u_xpb_out[104][7],u_xpb_out[105][7]};

assign col_out_8 = {u_xpb_out[0][8],u_xpb_out[1][8],u_xpb_out[2][8],u_xpb_out[3][8],u_xpb_out[4][8],u_xpb_out[5][8],u_xpb_out[6][8],u_xpb_out[7][8],u_xpb_out[8][8],u_xpb_out[9][8],u_xpb_out[10][8],u_xpb_out[11][8],u_xpb_out[12][8],u_xpb_out[13][8],u_xpb_out[14][8],u_xpb_out[15][8],u_xpb_out[16][8],u_xpb_out[17][8],u_xpb_out[18][8],u_xpb_out[19][8],u_xpb_out[20][8],u_xpb_out[21][8],u_xpb_out[22][8],u_xpb_out[23][8],u_xpb_out[24][8],u_xpb_out[25][8],u_xpb_out[26][8],u_xpb_out[27][8],u_xpb_out[28][8],u_xpb_out[29][8],u_xpb_out[30][8],u_xpb_out[31][8],u_xpb_out[32][8],u_xpb_out[33][8],u_xpb_out[34][8],u_xpb_out[35][8],u_xpb_out[36][8],u_xpb_out[37][8],u_xpb_out[38][8],u_xpb_out[39][8],u_xpb_out[40][8],u_xpb_out[41][8],u_xpb_out[42][8],u_xpb_out[43][8],u_xpb_out[44][8],u_xpb_out[45][8],u_xpb_out[46][8],u_xpb_out[47][8],u_xpb_out[48][8],u_xpb_out[49][8],u_xpb_out[50][8],u_xpb_out[51][8],u_xpb_out[52][8],u_xpb_out[53][8],u_xpb_out[54][8],u_xpb_out[55][8],u_xpb_out[56][8],u_xpb_out[57][8],u_xpb_out[58][8],u_xpb_out[59][8],u_xpb_out[60][8],u_xpb_out[61][8],u_xpb_out[62][8],u_xpb_out[63][8],u_xpb_out[64][8],u_xpb_out[65][8],u_xpb_out[66][8],u_xpb_out[67][8],u_xpb_out[68][8],u_xpb_out[69][8],u_xpb_out[70][8],u_xpb_out[71][8],u_xpb_out[72][8],u_xpb_out[73][8],u_xpb_out[74][8],u_xpb_out[75][8],u_xpb_out[76][8],u_xpb_out[77][8],u_xpb_out[78][8],u_xpb_out[79][8],u_xpb_out[80][8],u_xpb_out[81][8],u_xpb_out[82][8],u_xpb_out[83][8],u_xpb_out[84][8],u_xpb_out[85][8],u_xpb_out[86][8],u_xpb_out[87][8],u_xpb_out[88][8],u_xpb_out[89][8],u_xpb_out[90][8],u_xpb_out[91][8],u_xpb_out[92][8],u_xpb_out[93][8],u_xpb_out[94][8],u_xpb_out[95][8],u_xpb_out[96][8],u_xpb_out[97][8],u_xpb_out[98][8],u_xpb_out[99][8],u_xpb_out[100][8],u_xpb_out[101][8],u_xpb_out[102][8],u_xpb_out[103][8],u_xpb_out[104][8],u_xpb_out[105][8]};

assign col_out_9 = {u_xpb_out[0][9],u_xpb_out[1][9],u_xpb_out[2][9],u_xpb_out[3][9],u_xpb_out[4][9],u_xpb_out[5][9],u_xpb_out[6][9],u_xpb_out[7][9],u_xpb_out[8][9],u_xpb_out[9][9],u_xpb_out[10][9],u_xpb_out[11][9],u_xpb_out[12][9],u_xpb_out[13][9],u_xpb_out[14][9],u_xpb_out[15][9],u_xpb_out[16][9],u_xpb_out[17][9],u_xpb_out[18][9],u_xpb_out[19][9],u_xpb_out[20][9],u_xpb_out[21][9],u_xpb_out[22][9],u_xpb_out[23][9],u_xpb_out[24][9],u_xpb_out[25][9],u_xpb_out[26][9],u_xpb_out[27][9],u_xpb_out[28][9],u_xpb_out[29][9],u_xpb_out[30][9],u_xpb_out[31][9],u_xpb_out[32][9],u_xpb_out[33][9],u_xpb_out[34][9],u_xpb_out[35][9],u_xpb_out[36][9],u_xpb_out[37][9],u_xpb_out[38][9],u_xpb_out[39][9],u_xpb_out[40][9],u_xpb_out[41][9],u_xpb_out[42][9],u_xpb_out[43][9],u_xpb_out[44][9],u_xpb_out[45][9],u_xpb_out[46][9],u_xpb_out[47][9],u_xpb_out[48][9],u_xpb_out[49][9],u_xpb_out[50][9],u_xpb_out[51][9],u_xpb_out[52][9],u_xpb_out[53][9],u_xpb_out[54][9],u_xpb_out[55][9],u_xpb_out[56][9],u_xpb_out[57][9],u_xpb_out[58][9],u_xpb_out[59][9],u_xpb_out[60][9],u_xpb_out[61][9],u_xpb_out[62][9],u_xpb_out[63][9],u_xpb_out[64][9],u_xpb_out[65][9],u_xpb_out[66][9],u_xpb_out[67][9],u_xpb_out[68][9],u_xpb_out[69][9],u_xpb_out[70][9],u_xpb_out[71][9],u_xpb_out[72][9],u_xpb_out[73][9],u_xpb_out[74][9],u_xpb_out[75][9],u_xpb_out[76][9],u_xpb_out[77][9],u_xpb_out[78][9],u_xpb_out[79][9],u_xpb_out[80][9],u_xpb_out[81][9],u_xpb_out[82][9],u_xpb_out[83][9],u_xpb_out[84][9],u_xpb_out[85][9],u_xpb_out[86][9],u_xpb_out[87][9],u_xpb_out[88][9],u_xpb_out[89][9],u_xpb_out[90][9],u_xpb_out[91][9],u_xpb_out[92][9],u_xpb_out[93][9],u_xpb_out[94][9],u_xpb_out[95][9],u_xpb_out[96][9],u_xpb_out[97][9],u_xpb_out[98][9],u_xpb_out[99][9],u_xpb_out[100][9],u_xpb_out[101][9],u_xpb_out[102][9],u_xpb_out[103][9],u_xpb_out[104][9],u_xpb_out[105][9]};

assign col_out_10 = {u_xpb_out[0][10],u_xpb_out[1][10],u_xpb_out[2][10],u_xpb_out[3][10],u_xpb_out[4][10],u_xpb_out[5][10],u_xpb_out[6][10],u_xpb_out[7][10],u_xpb_out[8][10],u_xpb_out[9][10],u_xpb_out[10][10],u_xpb_out[11][10],u_xpb_out[12][10],u_xpb_out[13][10],u_xpb_out[14][10],u_xpb_out[15][10],u_xpb_out[16][10],u_xpb_out[17][10],u_xpb_out[18][10],u_xpb_out[19][10],u_xpb_out[20][10],u_xpb_out[21][10],u_xpb_out[22][10],u_xpb_out[23][10],u_xpb_out[24][10],u_xpb_out[25][10],u_xpb_out[26][10],u_xpb_out[27][10],u_xpb_out[28][10],u_xpb_out[29][10],u_xpb_out[30][10],u_xpb_out[31][10],u_xpb_out[32][10],u_xpb_out[33][10],u_xpb_out[34][10],u_xpb_out[35][10],u_xpb_out[36][10],u_xpb_out[37][10],u_xpb_out[38][10],u_xpb_out[39][10],u_xpb_out[40][10],u_xpb_out[41][10],u_xpb_out[42][10],u_xpb_out[43][10],u_xpb_out[44][10],u_xpb_out[45][10],u_xpb_out[46][10],u_xpb_out[47][10],u_xpb_out[48][10],u_xpb_out[49][10],u_xpb_out[50][10],u_xpb_out[51][10],u_xpb_out[52][10],u_xpb_out[53][10],u_xpb_out[54][10],u_xpb_out[55][10],u_xpb_out[56][10],u_xpb_out[57][10],u_xpb_out[58][10],u_xpb_out[59][10],u_xpb_out[60][10],u_xpb_out[61][10],u_xpb_out[62][10],u_xpb_out[63][10],u_xpb_out[64][10],u_xpb_out[65][10],u_xpb_out[66][10],u_xpb_out[67][10],u_xpb_out[68][10],u_xpb_out[69][10],u_xpb_out[70][10],u_xpb_out[71][10],u_xpb_out[72][10],u_xpb_out[73][10],u_xpb_out[74][10],u_xpb_out[75][10],u_xpb_out[76][10],u_xpb_out[77][10],u_xpb_out[78][10],u_xpb_out[79][10],u_xpb_out[80][10],u_xpb_out[81][10],u_xpb_out[82][10],u_xpb_out[83][10],u_xpb_out[84][10],u_xpb_out[85][10],u_xpb_out[86][10],u_xpb_out[87][10],u_xpb_out[88][10],u_xpb_out[89][10],u_xpb_out[90][10],u_xpb_out[91][10],u_xpb_out[92][10],u_xpb_out[93][10],u_xpb_out[94][10],u_xpb_out[95][10],u_xpb_out[96][10],u_xpb_out[97][10],u_xpb_out[98][10],u_xpb_out[99][10],u_xpb_out[100][10],u_xpb_out[101][10],u_xpb_out[102][10],u_xpb_out[103][10],u_xpb_out[104][10],u_xpb_out[105][10]};

assign col_out_11 = {u_xpb_out[0][11],u_xpb_out[1][11],u_xpb_out[2][11],u_xpb_out[3][11],u_xpb_out[4][11],u_xpb_out[5][11],u_xpb_out[6][11],u_xpb_out[7][11],u_xpb_out[8][11],u_xpb_out[9][11],u_xpb_out[10][11],u_xpb_out[11][11],u_xpb_out[12][11],u_xpb_out[13][11],u_xpb_out[14][11],u_xpb_out[15][11],u_xpb_out[16][11],u_xpb_out[17][11],u_xpb_out[18][11],u_xpb_out[19][11],u_xpb_out[20][11],u_xpb_out[21][11],u_xpb_out[22][11],u_xpb_out[23][11],u_xpb_out[24][11],u_xpb_out[25][11],u_xpb_out[26][11],u_xpb_out[27][11],u_xpb_out[28][11],u_xpb_out[29][11],u_xpb_out[30][11],u_xpb_out[31][11],u_xpb_out[32][11],u_xpb_out[33][11],u_xpb_out[34][11],u_xpb_out[35][11],u_xpb_out[36][11],u_xpb_out[37][11],u_xpb_out[38][11],u_xpb_out[39][11],u_xpb_out[40][11],u_xpb_out[41][11],u_xpb_out[42][11],u_xpb_out[43][11],u_xpb_out[44][11],u_xpb_out[45][11],u_xpb_out[46][11],u_xpb_out[47][11],u_xpb_out[48][11],u_xpb_out[49][11],u_xpb_out[50][11],u_xpb_out[51][11],u_xpb_out[52][11],u_xpb_out[53][11],u_xpb_out[54][11],u_xpb_out[55][11],u_xpb_out[56][11],u_xpb_out[57][11],u_xpb_out[58][11],u_xpb_out[59][11],u_xpb_out[60][11],u_xpb_out[61][11],u_xpb_out[62][11],u_xpb_out[63][11],u_xpb_out[64][11],u_xpb_out[65][11],u_xpb_out[66][11],u_xpb_out[67][11],u_xpb_out[68][11],u_xpb_out[69][11],u_xpb_out[70][11],u_xpb_out[71][11],u_xpb_out[72][11],u_xpb_out[73][11],u_xpb_out[74][11],u_xpb_out[75][11],u_xpb_out[76][11],u_xpb_out[77][11],u_xpb_out[78][11],u_xpb_out[79][11],u_xpb_out[80][11],u_xpb_out[81][11],u_xpb_out[82][11],u_xpb_out[83][11],u_xpb_out[84][11],u_xpb_out[85][11],u_xpb_out[86][11],u_xpb_out[87][11],u_xpb_out[88][11],u_xpb_out[89][11],u_xpb_out[90][11],u_xpb_out[91][11],u_xpb_out[92][11],u_xpb_out[93][11],u_xpb_out[94][11],u_xpb_out[95][11],u_xpb_out[96][11],u_xpb_out[97][11],u_xpb_out[98][11],u_xpb_out[99][11],u_xpb_out[100][11],u_xpb_out[101][11],u_xpb_out[102][11],u_xpb_out[103][11],u_xpb_out[104][11],u_xpb_out[105][11]};

assign col_out_12 = {u_xpb_out[0][12],u_xpb_out[1][12],u_xpb_out[2][12],u_xpb_out[3][12],u_xpb_out[4][12],u_xpb_out[5][12],u_xpb_out[6][12],u_xpb_out[7][12],u_xpb_out[8][12],u_xpb_out[9][12],u_xpb_out[10][12],u_xpb_out[11][12],u_xpb_out[12][12],u_xpb_out[13][12],u_xpb_out[14][12],u_xpb_out[15][12],u_xpb_out[16][12],u_xpb_out[17][12],u_xpb_out[18][12],u_xpb_out[19][12],u_xpb_out[20][12],u_xpb_out[21][12],u_xpb_out[22][12],u_xpb_out[23][12],u_xpb_out[24][12],u_xpb_out[25][12],u_xpb_out[26][12],u_xpb_out[27][12],u_xpb_out[28][12],u_xpb_out[29][12],u_xpb_out[30][12],u_xpb_out[31][12],u_xpb_out[32][12],u_xpb_out[33][12],u_xpb_out[34][12],u_xpb_out[35][12],u_xpb_out[36][12],u_xpb_out[37][12],u_xpb_out[38][12],u_xpb_out[39][12],u_xpb_out[40][12],u_xpb_out[41][12],u_xpb_out[42][12],u_xpb_out[43][12],u_xpb_out[44][12],u_xpb_out[45][12],u_xpb_out[46][12],u_xpb_out[47][12],u_xpb_out[48][12],u_xpb_out[49][12],u_xpb_out[50][12],u_xpb_out[51][12],u_xpb_out[52][12],u_xpb_out[53][12],u_xpb_out[54][12],u_xpb_out[55][12],u_xpb_out[56][12],u_xpb_out[57][12],u_xpb_out[58][12],u_xpb_out[59][12],u_xpb_out[60][12],u_xpb_out[61][12],u_xpb_out[62][12],u_xpb_out[63][12],u_xpb_out[64][12],u_xpb_out[65][12],u_xpb_out[66][12],u_xpb_out[67][12],u_xpb_out[68][12],u_xpb_out[69][12],u_xpb_out[70][12],u_xpb_out[71][12],u_xpb_out[72][12],u_xpb_out[73][12],u_xpb_out[74][12],u_xpb_out[75][12],u_xpb_out[76][12],u_xpb_out[77][12],u_xpb_out[78][12],u_xpb_out[79][12],u_xpb_out[80][12],u_xpb_out[81][12],u_xpb_out[82][12],u_xpb_out[83][12],u_xpb_out[84][12],u_xpb_out[85][12],u_xpb_out[86][12],u_xpb_out[87][12],u_xpb_out[88][12],u_xpb_out[89][12],u_xpb_out[90][12],u_xpb_out[91][12],u_xpb_out[92][12],u_xpb_out[93][12],u_xpb_out[94][12],u_xpb_out[95][12],u_xpb_out[96][12],u_xpb_out[97][12],u_xpb_out[98][12],u_xpb_out[99][12],u_xpb_out[100][12],u_xpb_out[101][12],u_xpb_out[102][12],u_xpb_out[103][12],u_xpb_out[104][12],u_xpb_out[105][12]};

assign col_out_13 = {u_xpb_out[0][13],u_xpb_out[1][13],u_xpb_out[2][13],u_xpb_out[3][13],u_xpb_out[4][13],u_xpb_out[5][13],u_xpb_out[6][13],u_xpb_out[7][13],u_xpb_out[8][13],u_xpb_out[9][13],u_xpb_out[10][13],u_xpb_out[11][13],u_xpb_out[12][13],u_xpb_out[13][13],u_xpb_out[14][13],u_xpb_out[15][13],u_xpb_out[16][13],u_xpb_out[17][13],u_xpb_out[18][13],u_xpb_out[19][13],u_xpb_out[20][13],u_xpb_out[21][13],u_xpb_out[22][13],u_xpb_out[23][13],u_xpb_out[24][13],u_xpb_out[25][13],u_xpb_out[26][13],u_xpb_out[27][13],u_xpb_out[28][13],u_xpb_out[29][13],u_xpb_out[30][13],u_xpb_out[31][13],u_xpb_out[32][13],u_xpb_out[33][13],u_xpb_out[34][13],u_xpb_out[35][13],u_xpb_out[36][13],u_xpb_out[37][13],u_xpb_out[38][13],u_xpb_out[39][13],u_xpb_out[40][13],u_xpb_out[41][13],u_xpb_out[42][13],u_xpb_out[43][13],u_xpb_out[44][13],u_xpb_out[45][13],u_xpb_out[46][13],u_xpb_out[47][13],u_xpb_out[48][13],u_xpb_out[49][13],u_xpb_out[50][13],u_xpb_out[51][13],u_xpb_out[52][13],u_xpb_out[53][13],u_xpb_out[54][13],u_xpb_out[55][13],u_xpb_out[56][13],u_xpb_out[57][13],u_xpb_out[58][13],u_xpb_out[59][13],u_xpb_out[60][13],u_xpb_out[61][13],u_xpb_out[62][13],u_xpb_out[63][13],u_xpb_out[64][13],u_xpb_out[65][13],u_xpb_out[66][13],u_xpb_out[67][13],u_xpb_out[68][13],u_xpb_out[69][13],u_xpb_out[70][13],u_xpb_out[71][13],u_xpb_out[72][13],u_xpb_out[73][13],u_xpb_out[74][13],u_xpb_out[75][13],u_xpb_out[76][13],u_xpb_out[77][13],u_xpb_out[78][13],u_xpb_out[79][13],u_xpb_out[80][13],u_xpb_out[81][13],u_xpb_out[82][13],u_xpb_out[83][13],u_xpb_out[84][13],u_xpb_out[85][13],u_xpb_out[86][13],u_xpb_out[87][13],u_xpb_out[88][13],u_xpb_out[89][13],u_xpb_out[90][13],u_xpb_out[91][13],u_xpb_out[92][13],u_xpb_out[93][13],u_xpb_out[94][13],u_xpb_out[95][13],u_xpb_out[96][13],u_xpb_out[97][13],u_xpb_out[98][13],u_xpb_out[99][13],u_xpb_out[100][13],u_xpb_out[101][13],u_xpb_out[102][13],u_xpb_out[103][13],u_xpb_out[104][13],u_xpb_out[105][13]};

assign col_out_14 = {u_xpb_out[0][14],u_xpb_out[1][14],u_xpb_out[2][14],u_xpb_out[3][14],u_xpb_out[4][14],u_xpb_out[5][14],u_xpb_out[6][14],u_xpb_out[7][14],u_xpb_out[8][14],u_xpb_out[9][14],u_xpb_out[10][14],u_xpb_out[11][14],u_xpb_out[12][14],u_xpb_out[13][14],u_xpb_out[14][14],u_xpb_out[15][14],u_xpb_out[16][14],u_xpb_out[17][14],u_xpb_out[18][14],u_xpb_out[19][14],u_xpb_out[20][14],u_xpb_out[21][14],u_xpb_out[22][14],u_xpb_out[23][14],u_xpb_out[24][14],u_xpb_out[25][14],u_xpb_out[26][14],u_xpb_out[27][14],u_xpb_out[28][14],u_xpb_out[29][14],u_xpb_out[30][14],u_xpb_out[31][14],u_xpb_out[32][14],u_xpb_out[33][14],u_xpb_out[34][14],u_xpb_out[35][14],u_xpb_out[36][14],u_xpb_out[37][14],u_xpb_out[38][14],u_xpb_out[39][14],u_xpb_out[40][14],u_xpb_out[41][14],u_xpb_out[42][14],u_xpb_out[43][14],u_xpb_out[44][14],u_xpb_out[45][14],u_xpb_out[46][14],u_xpb_out[47][14],u_xpb_out[48][14],u_xpb_out[49][14],u_xpb_out[50][14],u_xpb_out[51][14],u_xpb_out[52][14],u_xpb_out[53][14],u_xpb_out[54][14],u_xpb_out[55][14],u_xpb_out[56][14],u_xpb_out[57][14],u_xpb_out[58][14],u_xpb_out[59][14],u_xpb_out[60][14],u_xpb_out[61][14],u_xpb_out[62][14],u_xpb_out[63][14],u_xpb_out[64][14],u_xpb_out[65][14],u_xpb_out[66][14],u_xpb_out[67][14],u_xpb_out[68][14],u_xpb_out[69][14],u_xpb_out[70][14],u_xpb_out[71][14],u_xpb_out[72][14],u_xpb_out[73][14],u_xpb_out[74][14],u_xpb_out[75][14],u_xpb_out[76][14],u_xpb_out[77][14],u_xpb_out[78][14],u_xpb_out[79][14],u_xpb_out[80][14],u_xpb_out[81][14],u_xpb_out[82][14],u_xpb_out[83][14],u_xpb_out[84][14],u_xpb_out[85][14],u_xpb_out[86][14],u_xpb_out[87][14],u_xpb_out[88][14],u_xpb_out[89][14],u_xpb_out[90][14],u_xpb_out[91][14],u_xpb_out[92][14],u_xpb_out[93][14],u_xpb_out[94][14],u_xpb_out[95][14],u_xpb_out[96][14],u_xpb_out[97][14],u_xpb_out[98][14],u_xpb_out[99][14],u_xpb_out[100][14],u_xpb_out[101][14],u_xpb_out[102][14],u_xpb_out[103][14],u_xpb_out[104][14],u_xpb_out[105][14]};

assign col_out_15 = {u_xpb_out[0][15],u_xpb_out[1][15],u_xpb_out[2][15],u_xpb_out[3][15],u_xpb_out[4][15],u_xpb_out[5][15],u_xpb_out[6][15],u_xpb_out[7][15],u_xpb_out[8][15],u_xpb_out[9][15],u_xpb_out[10][15],u_xpb_out[11][15],u_xpb_out[12][15],u_xpb_out[13][15],u_xpb_out[14][15],u_xpb_out[15][15],u_xpb_out[16][15],u_xpb_out[17][15],u_xpb_out[18][15],u_xpb_out[19][15],u_xpb_out[20][15],u_xpb_out[21][15],u_xpb_out[22][15],u_xpb_out[23][15],u_xpb_out[24][15],u_xpb_out[25][15],u_xpb_out[26][15],u_xpb_out[27][15],u_xpb_out[28][15],u_xpb_out[29][15],u_xpb_out[30][15],u_xpb_out[31][15],u_xpb_out[32][15],u_xpb_out[33][15],u_xpb_out[34][15],u_xpb_out[35][15],u_xpb_out[36][15],u_xpb_out[37][15],u_xpb_out[38][15],u_xpb_out[39][15],u_xpb_out[40][15],u_xpb_out[41][15],u_xpb_out[42][15],u_xpb_out[43][15],u_xpb_out[44][15],u_xpb_out[45][15],u_xpb_out[46][15],u_xpb_out[47][15],u_xpb_out[48][15],u_xpb_out[49][15],u_xpb_out[50][15],u_xpb_out[51][15],u_xpb_out[52][15],u_xpb_out[53][15],u_xpb_out[54][15],u_xpb_out[55][15],u_xpb_out[56][15],u_xpb_out[57][15],u_xpb_out[58][15],u_xpb_out[59][15],u_xpb_out[60][15],u_xpb_out[61][15],u_xpb_out[62][15],u_xpb_out[63][15],u_xpb_out[64][15],u_xpb_out[65][15],u_xpb_out[66][15],u_xpb_out[67][15],u_xpb_out[68][15],u_xpb_out[69][15],u_xpb_out[70][15],u_xpb_out[71][15],u_xpb_out[72][15],u_xpb_out[73][15],u_xpb_out[74][15],u_xpb_out[75][15],u_xpb_out[76][15],u_xpb_out[77][15],u_xpb_out[78][15],u_xpb_out[79][15],u_xpb_out[80][15],u_xpb_out[81][15],u_xpb_out[82][15],u_xpb_out[83][15],u_xpb_out[84][15],u_xpb_out[85][15],u_xpb_out[86][15],u_xpb_out[87][15],u_xpb_out[88][15],u_xpb_out[89][15],u_xpb_out[90][15],u_xpb_out[91][15],u_xpb_out[92][15],u_xpb_out[93][15],u_xpb_out[94][15],u_xpb_out[95][15],u_xpb_out[96][15],u_xpb_out[97][15],u_xpb_out[98][15],u_xpb_out[99][15],u_xpb_out[100][15],u_xpb_out[101][15],u_xpb_out[102][15],u_xpb_out[103][15],u_xpb_out[104][15],u_xpb_out[105][15]};

assign col_out_16 = {u_xpb_out[0][16],u_xpb_out[1][16],u_xpb_out[2][16],u_xpb_out[3][16],u_xpb_out[4][16],u_xpb_out[5][16],u_xpb_out[6][16],u_xpb_out[7][16],u_xpb_out[8][16],u_xpb_out[9][16],u_xpb_out[10][16],u_xpb_out[11][16],u_xpb_out[12][16],u_xpb_out[13][16],u_xpb_out[14][16],u_xpb_out[15][16],u_xpb_out[16][16],u_xpb_out[17][16],u_xpb_out[18][16],u_xpb_out[19][16],u_xpb_out[20][16],u_xpb_out[21][16],u_xpb_out[22][16],u_xpb_out[23][16],u_xpb_out[24][16],u_xpb_out[25][16],u_xpb_out[26][16],u_xpb_out[27][16],u_xpb_out[28][16],u_xpb_out[29][16],u_xpb_out[30][16],u_xpb_out[31][16],u_xpb_out[32][16],u_xpb_out[33][16],u_xpb_out[34][16],u_xpb_out[35][16],u_xpb_out[36][16],u_xpb_out[37][16],u_xpb_out[38][16],u_xpb_out[39][16],u_xpb_out[40][16],u_xpb_out[41][16],u_xpb_out[42][16],u_xpb_out[43][16],u_xpb_out[44][16],u_xpb_out[45][16],u_xpb_out[46][16],u_xpb_out[47][16],u_xpb_out[48][16],u_xpb_out[49][16],u_xpb_out[50][16],u_xpb_out[51][16],u_xpb_out[52][16],u_xpb_out[53][16],u_xpb_out[54][16],u_xpb_out[55][16],u_xpb_out[56][16],u_xpb_out[57][16],u_xpb_out[58][16],u_xpb_out[59][16],u_xpb_out[60][16],u_xpb_out[61][16],u_xpb_out[62][16],u_xpb_out[63][16],u_xpb_out[64][16],u_xpb_out[65][16],u_xpb_out[66][16],u_xpb_out[67][16],u_xpb_out[68][16],u_xpb_out[69][16],u_xpb_out[70][16],u_xpb_out[71][16],u_xpb_out[72][16],u_xpb_out[73][16],u_xpb_out[74][16],u_xpb_out[75][16],u_xpb_out[76][16],u_xpb_out[77][16],u_xpb_out[78][16],u_xpb_out[79][16],u_xpb_out[80][16],u_xpb_out[81][16],u_xpb_out[82][16],u_xpb_out[83][16],u_xpb_out[84][16],u_xpb_out[85][16],u_xpb_out[86][16],u_xpb_out[87][16],u_xpb_out[88][16],u_xpb_out[89][16],u_xpb_out[90][16],u_xpb_out[91][16],u_xpb_out[92][16],u_xpb_out[93][16],u_xpb_out[94][16],u_xpb_out[95][16],u_xpb_out[96][16],u_xpb_out[97][16],u_xpb_out[98][16],u_xpb_out[99][16],u_xpb_out[100][16],u_xpb_out[101][16],u_xpb_out[102][16],u_xpb_out[103][16],u_xpb_out[104][16],u_xpb_out[105][16]};

assign col_out_17 = {u_xpb_out[0][17],u_xpb_out[1][17],u_xpb_out[2][17],u_xpb_out[3][17],u_xpb_out[4][17],u_xpb_out[5][17],u_xpb_out[6][17],u_xpb_out[7][17],u_xpb_out[8][17],u_xpb_out[9][17],u_xpb_out[10][17],u_xpb_out[11][17],u_xpb_out[12][17],u_xpb_out[13][17],u_xpb_out[14][17],u_xpb_out[15][17],u_xpb_out[16][17],u_xpb_out[17][17],u_xpb_out[18][17],u_xpb_out[19][17],u_xpb_out[20][17],u_xpb_out[21][17],u_xpb_out[22][17],u_xpb_out[23][17],u_xpb_out[24][17],u_xpb_out[25][17],u_xpb_out[26][17],u_xpb_out[27][17],u_xpb_out[28][17],u_xpb_out[29][17],u_xpb_out[30][17],u_xpb_out[31][17],u_xpb_out[32][17],u_xpb_out[33][17],u_xpb_out[34][17],u_xpb_out[35][17],u_xpb_out[36][17],u_xpb_out[37][17],u_xpb_out[38][17],u_xpb_out[39][17],u_xpb_out[40][17],u_xpb_out[41][17],u_xpb_out[42][17],u_xpb_out[43][17],u_xpb_out[44][17],u_xpb_out[45][17],u_xpb_out[46][17],u_xpb_out[47][17],u_xpb_out[48][17],u_xpb_out[49][17],u_xpb_out[50][17],u_xpb_out[51][17],u_xpb_out[52][17],u_xpb_out[53][17],u_xpb_out[54][17],u_xpb_out[55][17],u_xpb_out[56][17],u_xpb_out[57][17],u_xpb_out[58][17],u_xpb_out[59][17],u_xpb_out[60][17],u_xpb_out[61][17],u_xpb_out[62][17],u_xpb_out[63][17],u_xpb_out[64][17],u_xpb_out[65][17],u_xpb_out[66][17],u_xpb_out[67][17],u_xpb_out[68][17],u_xpb_out[69][17],u_xpb_out[70][17],u_xpb_out[71][17],u_xpb_out[72][17],u_xpb_out[73][17],u_xpb_out[74][17],u_xpb_out[75][17],u_xpb_out[76][17],u_xpb_out[77][17],u_xpb_out[78][17],u_xpb_out[79][17],u_xpb_out[80][17],u_xpb_out[81][17],u_xpb_out[82][17],u_xpb_out[83][17],u_xpb_out[84][17],u_xpb_out[85][17],u_xpb_out[86][17],u_xpb_out[87][17],u_xpb_out[88][17],u_xpb_out[89][17],u_xpb_out[90][17],u_xpb_out[91][17],u_xpb_out[92][17],u_xpb_out[93][17],u_xpb_out[94][17],u_xpb_out[95][17],u_xpb_out[96][17],u_xpb_out[97][17],u_xpb_out[98][17],u_xpb_out[99][17],u_xpb_out[100][17],u_xpb_out[101][17],u_xpb_out[102][17],u_xpb_out[103][17],u_xpb_out[104][17],u_xpb_out[105][17]};

assign col_out_18 = {u_xpb_out[0][18],u_xpb_out[1][18],u_xpb_out[2][18],u_xpb_out[3][18],u_xpb_out[4][18],u_xpb_out[5][18],u_xpb_out[6][18],u_xpb_out[7][18],u_xpb_out[8][18],u_xpb_out[9][18],u_xpb_out[10][18],u_xpb_out[11][18],u_xpb_out[12][18],u_xpb_out[13][18],u_xpb_out[14][18],u_xpb_out[15][18],u_xpb_out[16][18],u_xpb_out[17][18],u_xpb_out[18][18],u_xpb_out[19][18],u_xpb_out[20][18],u_xpb_out[21][18],u_xpb_out[22][18],u_xpb_out[23][18],u_xpb_out[24][18],u_xpb_out[25][18],u_xpb_out[26][18],u_xpb_out[27][18],u_xpb_out[28][18],u_xpb_out[29][18],u_xpb_out[30][18],u_xpb_out[31][18],u_xpb_out[32][18],u_xpb_out[33][18],u_xpb_out[34][18],u_xpb_out[35][18],u_xpb_out[36][18],u_xpb_out[37][18],u_xpb_out[38][18],u_xpb_out[39][18],u_xpb_out[40][18],u_xpb_out[41][18],u_xpb_out[42][18],u_xpb_out[43][18],u_xpb_out[44][18],u_xpb_out[45][18],u_xpb_out[46][18],u_xpb_out[47][18],u_xpb_out[48][18],u_xpb_out[49][18],u_xpb_out[50][18],u_xpb_out[51][18],u_xpb_out[52][18],u_xpb_out[53][18],u_xpb_out[54][18],u_xpb_out[55][18],u_xpb_out[56][18],u_xpb_out[57][18],u_xpb_out[58][18],u_xpb_out[59][18],u_xpb_out[60][18],u_xpb_out[61][18],u_xpb_out[62][18],u_xpb_out[63][18],u_xpb_out[64][18],u_xpb_out[65][18],u_xpb_out[66][18],u_xpb_out[67][18],u_xpb_out[68][18],u_xpb_out[69][18],u_xpb_out[70][18],u_xpb_out[71][18],u_xpb_out[72][18],u_xpb_out[73][18],u_xpb_out[74][18],u_xpb_out[75][18],u_xpb_out[76][18],u_xpb_out[77][18],u_xpb_out[78][18],u_xpb_out[79][18],u_xpb_out[80][18],u_xpb_out[81][18],u_xpb_out[82][18],u_xpb_out[83][18],u_xpb_out[84][18],u_xpb_out[85][18],u_xpb_out[86][18],u_xpb_out[87][18],u_xpb_out[88][18],u_xpb_out[89][18],u_xpb_out[90][18],u_xpb_out[91][18],u_xpb_out[92][18],u_xpb_out[93][18],u_xpb_out[94][18],u_xpb_out[95][18],u_xpb_out[96][18],u_xpb_out[97][18],u_xpb_out[98][18],u_xpb_out[99][18],u_xpb_out[100][18],u_xpb_out[101][18],u_xpb_out[102][18],u_xpb_out[103][18],u_xpb_out[104][18],u_xpb_out[105][18]};

assign col_out_19 = {u_xpb_out[0][19],u_xpb_out[1][19],u_xpb_out[2][19],u_xpb_out[3][19],u_xpb_out[4][19],u_xpb_out[5][19],u_xpb_out[6][19],u_xpb_out[7][19],u_xpb_out[8][19],u_xpb_out[9][19],u_xpb_out[10][19],u_xpb_out[11][19],u_xpb_out[12][19],u_xpb_out[13][19],u_xpb_out[14][19],u_xpb_out[15][19],u_xpb_out[16][19],u_xpb_out[17][19],u_xpb_out[18][19],u_xpb_out[19][19],u_xpb_out[20][19],u_xpb_out[21][19],u_xpb_out[22][19],u_xpb_out[23][19],u_xpb_out[24][19],u_xpb_out[25][19],u_xpb_out[26][19],u_xpb_out[27][19],u_xpb_out[28][19],u_xpb_out[29][19],u_xpb_out[30][19],u_xpb_out[31][19],u_xpb_out[32][19],u_xpb_out[33][19],u_xpb_out[34][19],u_xpb_out[35][19],u_xpb_out[36][19],u_xpb_out[37][19],u_xpb_out[38][19],u_xpb_out[39][19],u_xpb_out[40][19],u_xpb_out[41][19],u_xpb_out[42][19],u_xpb_out[43][19],u_xpb_out[44][19],u_xpb_out[45][19],u_xpb_out[46][19],u_xpb_out[47][19],u_xpb_out[48][19],u_xpb_out[49][19],u_xpb_out[50][19],u_xpb_out[51][19],u_xpb_out[52][19],u_xpb_out[53][19],u_xpb_out[54][19],u_xpb_out[55][19],u_xpb_out[56][19],u_xpb_out[57][19],u_xpb_out[58][19],u_xpb_out[59][19],u_xpb_out[60][19],u_xpb_out[61][19],u_xpb_out[62][19],u_xpb_out[63][19],u_xpb_out[64][19],u_xpb_out[65][19],u_xpb_out[66][19],u_xpb_out[67][19],u_xpb_out[68][19],u_xpb_out[69][19],u_xpb_out[70][19],u_xpb_out[71][19],u_xpb_out[72][19],u_xpb_out[73][19],u_xpb_out[74][19],u_xpb_out[75][19],u_xpb_out[76][19],u_xpb_out[77][19],u_xpb_out[78][19],u_xpb_out[79][19],u_xpb_out[80][19],u_xpb_out[81][19],u_xpb_out[82][19],u_xpb_out[83][19],u_xpb_out[84][19],u_xpb_out[85][19],u_xpb_out[86][19],u_xpb_out[87][19],u_xpb_out[88][19],u_xpb_out[89][19],u_xpb_out[90][19],u_xpb_out[91][19],u_xpb_out[92][19],u_xpb_out[93][19],u_xpb_out[94][19],u_xpb_out[95][19],u_xpb_out[96][19],u_xpb_out[97][19],u_xpb_out[98][19],u_xpb_out[99][19],u_xpb_out[100][19],u_xpb_out[101][19],u_xpb_out[102][19],u_xpb_out[103][19],u_xpb_out[104][19],u_xpb_out[105][19]};

assign col_out_20 = {u_xpb_out[0][20],u_xpb_out[1][20],u_xpb_out[2][20],u_xpb_out[3][20],u_xpb_out[4][20],u_xpb_out[5][20],u_xpb_out[6][20],u_xpb_out[7][20],u_xpb_out[8][20],u_xpb_out[9][20],u_xpb_out[10][20],u_xpb_out[11][20],u_xpb_out[12][20],u_xpb_out[13][20],u_xpb_out[14][20],u_xpb_out[15][20],u_xpb_out[16][20],u_xpb_out[17][20],u_xpb_out[18][20],u_xpb_out[19][20],u_xpb_out[20][20],u_xpb_out[21][20],u_xpb_out[22][20],u_xpb_out[23][20],u_xpb_out[24][20],u_xpb_out[25][20],u_xpb_out[26][20],u_xpb_out[27][20],u_xpb_out[28][20],u_xpb_out[29][20],u_xpb_out[30][20],u_xpb_out[31][20],u_xpb_out[32][20],u_xpb_out[33][20],u_xpb_out[34][20],u_xpb_out[35][20],u_xpb_out[36][20],u_xpb_out[37][20],u_xpb_out[38][20],u_xpb_out[39][20],u_xpb_out[40][20],u_xpb_out[41][20],u_xpb_out[42][20],u_xpb_out[43][20],u_xpb_out[44][20],u_xpb_out[45][20],u_xpb_out[46][20],u_xpb_out[47][20],u_xpb_out[48][20],u_xpb_out[49][20],u_xpb_out[50][20],u_xpb_out[51][20],u_xpb_out[52][20],u_xpb_out[53][20],u_xpb_out[54][20],u_xpb_out[55][20],u_xpb_out[56][20],u_xpb_out[57][20],u_xpb_out[58][20],u_xpb_out[59][20],u_xpb_out[60][20],u_xpb_out[61][20],u_xpb_out[62][20],u_xpb_out[63][20],u_xpb_out[64][20],u_xpb_out[65][20],u_xpb_out[66][20],u_xpb_out[67][20],u_xpb_out[68][20],u_xpb_out[69][20],u_xpb_out[70][20],u_xpb_out[71][20],u_xpb_out[72][20],u_xpb_out[73][20],u_xpb_out[74][20],u_xpb_out[75][20],u_xpb_out[76][20],u_xpb_out[77][20],u_xpb_out[78][20],u_xpb_out[79][20],u_xpb_out[80][20],u_xpb_out[81][20],u_xpb_out[82][20],u_xpb_out[83][20],u_xpb_out[84][20],u_xpb_out[85][20],u_xpb_out[86][20],u_xpb_out[87][20],u_xpb_out[88][20],u_xpb_out[89][20],u_xpb_out[90][20],u_xpb_out[91][20],u_xpb_out[92][20],u_xpb_out[93][20],u_xpb_out[94][20],u_xpb_out[95][20],u_xpb_out[96][20],u_xpb_out[97][20],u_xpb_out[98][20],u_xpb_out[99][20],u_xpb_out[100][20],u_xpb_out[101][20],u_xpb_out[102][20],u_xpb_out[103][20],u_xpb_out[104][20],u_xpb_out[105][20]};

assign col_out_21 = {u_xpb_out[0][21],u_xpb_out[1][21],u_xpb_out[2][21],u_xpb_out[3][21],u_xpb_out[4][21],u_xpb_out[5][21],u_xpb_out[6][21],u_xpb_out[7][21],u_xpb_out[8][21],u_xpb_out[9][21],u_xpb_out[10][21],u_xpb_out[11][21],u_xpb_out[12][21],u_xpb_out[13][21],u_xpb_out[14][21],u_xpb_out[15][21],u_xpb_out[16][21],u_xpb_out[17][21],u_xpb_out[18][21],u_xpb_out[19][21],u_xpb_out[20][21],u_xpb_out[21][21],u_xpb_out[22][21],u_xpb_out[23][21],u_xpb_out[24][21],u_xpb_out[25][21],u_xpb_out[26][21],u_xpb_out[27][21],u_xpb_out[28][21],u_xpb_out[29][21],u_xpb_out[30][21],u_xpb_out[31][21],u_xpb_out[32][21],u_xpb_out[33][21],u_xpb_out[34][21],u_xpb_out[35][21],u_xpb_out[36][21],u_xpb_out[37][21],u_xpb_out[38][21],u_xpb_out[39][21],u_xpb_out[40][21],u_xpb_out[41][21],u_xpb_out[42][21],u_xpb_out[43][21],u_xpb_out[44][21],u_xpb_out[45][21],u_xpb_out[46][21],u_xpb_out[47][21],u_xpb_out[48][21],u_xpb_out[49][21],u_xpb_out[50][21],u_xpb_out[51][21],u_xpb_out[52][21],u_xpb_out[53][21],u_xpb_out[54][21],u_xpb_out[55][21],u_xpb_out[56][21],u_xpb_out[57][21],u_xpb_out[58][21],u_xpb_out[59][21],u_xpb_out[60][21],u_xpb_out[61][21],u_xpb_out[62][21],u_xpb_out[63][21],u_xpb_out[64][21],u_xpb_out[65][21],u_xpb_out[66][21],u_xpb_out[67][21],u_xpb_out[68][21],u_xpb_out[69][21],u_xpb_out[70][21],u_xpb_out[71][21],u_xpb_out[72][21],u_xpb_out[73][21],u_xpb_out[74][21],u_xpb_out[75][21],u_xpb_out[76][21],u_xpb_out[77][21],u_xpb_out[78][21],u_xpb_out[79][21],u_xpb_out[80][21],u_xpb_out[81][21],u_xpb_out[82][21],u_xpb_out[83][21],u_xpb_out[84][21],u_xpb_out[85][21],u_xpb_out[86][21],u_xpb_out[87][21],u_xpb_out[88][21],u_xpb_out[89][21],u_xpb_out[90][21],u_xpb_out[91][21],u_xpb_out[92][21],u_xpb_out[93][21],u_xpb_out[94][21],u_xpb_out[95][21],u_xpb_out[96][21],u_xpb_out[97][21],u_xpb_out[98][21],u_xpb_out[99][21],u_xpb_out[100][21],u_xpb_out[101][21],u_xpb_out[102][21],u_xpb_out[103][21],u_xpb_out[104][21],u_xpb_out[105][21]};

assign col_out_22 = {u_xpb_out[0][22],u_xpb_out[1][22],u_xpb_out[2][22],u_xpb_out[3][22],u_xpb_out[4][22],u_xpb_out[5][22],u_xpb_out[6][22],u_xpb_out[7][22],u_xpb_out[8][22],u_xpb_out[9][22],u_xpb_out[10][22],u_xpb_out[11][22],u_xpb_out[12][22],u_xpb_out[13][22],u_xpb_out[14][22],u_xpb_out[15][22],u_xpb_out[16][22],u_xpb_out[17][22],u_xpb_out[18][22],u_xpb_out[19][22],u_xpb_out[20][22],u_xpb_out[21][22],u_xpb_out[22][22],u_xpb_out[23][22],u_xpb_out[24][22],u_xpb_out[25][22],u_xpb_out[26][22],u_xpb_out[27][22],u_xpb_out[28][22],u_xpb_out[29][22],u_xpb_out[30][22],u_xpb_out[31][22],u_xpb_out[32][22],u_xpb_out[33][22],u_xpb_out[34][22],u_xpb_out[35][22],u_xpb_out[36][22],u_xpb_out[37][22],u_xpb_out[38][22],u_xpb_out[39][22],u_xpb_out[40][22],u_xpb_out[41][22],u_xpb_out[42][22],u_xpb_out[43][22],u_xpb_out[44][22],u_xpb_out[45][22],u_xpb_out[46][22],u_xpb_out[47][22],u_xpb_out[48][22],u_xpb_out[49][22],u_xpb_out[50][22],u_xpb_out[51][22],u_xpb_out[52][22],u_xpb_out[53][22],u_xpb_out[54][22],u_xpb_out[55][22],u_xpb_out[56][22],u_xpb_out[57][22],u_xpb_out[58][22],u_xpb_out[59][22],u_xpb_out[60][22],u_xpb_out[61][22],u_xpb_out[62][22],u_xpb_out[63][22],u_xpb_out[64][22],u_xpb_out[65][22],u_xpb_out[66][22],u_xpb_out[67][22],u_xpb_out[68][22],u_xpb_out[69][22],u_xpb_out[70][22],u_xpb_out[71][22],u_xpb_out[72][22],u_xpb_out[73][22],u_xpb_out[74][22],u_xpb_out[75][22],u_xpb_out[76][22],u_xpb_out[77][22],u_xpb_out[78][22],u_xpb_out[79][22],u_xpb_out[80][22],u_xpb_out[81][22],u_xpb_out[82][22],u_xpb_out[83][22],u_xpb_out[84][22],u_xpb_out[85][22],u_xpb_out[86][22],u_xpb_out[87][22],u_xpb_out[88][22],u_xpb_out[89][22],u_xpb_out[90][22],u_xpb_out[91][22],u_xpb_out[92][22],u_xpb_out[93][22],u_xpb_out[94][22],u_xpb_out[95][22],u_xpb_out[96][22],u_xpb_out[97][22],u_xpb_out[98][22],u_xpb_out[99][22],u_xpb_out[100][22],u_xpb_out[101][22],u_xpb_out[102][22],u_xpb_out[103][22],u_xpb_out[104][22],u_xpb_out[105][22]};

assign col_out_23 = {u_xpb_out[0][23],u_xpb_out[1][23],u_xpb_out[2][23],u_xpb_out[3][23],u_xpb_out[4][23],u_xpb_out[5][23],u_xpb_out[6][23],u_xpb_out[7][23],u_xpb_out[8][23],u_xpb_out[9][23],u_xpb_out[10][23],u_xpb_out[11][23],u_xpb_out[12][23],u_xpb_out[13][23],u_xpb_out[14][23],u_xpb_out[15][23],u_xpb_out[16][23],u_xpb_out[17][23],u_xpb_out[18][23],u_xpb_out[19][23],u_xpb_out[20][23],u_xpb_out[21][23],u_xpb_out[22][23],u_xpb_out[23][23],u_xpb_out[24][23],u_xpb_out[25][23],u_xpb_out[26][23],u_xpb_out[27][23],u_xpb_out[28][23],u_xpb_out[29][23],u_xpb_out[30][23],u_xpb_out[31][23],u_xpb_out[32][23],u_xpb_out[33][23],u_xpb_out[34][23],u_xpb_out[35][23],u_xpb_out[36][23],u_xpb_out[37][23],u_xpb_out[38][23],u_xpb_out[39][23],u_xpb_out[40][23],u_xpb_out[41][23],u_xpb_out[42][23],u_xpb_out[43][23],u_xpb_out[44][23],u_xpb_out[45][23],u_xpb_out[46][23],u_xpb_out[47][23],u_xpb_out[48][23],u_xpb_out[49][23],u_xpb_out[50][23],u_xpb_out[51][23],u_xpb_out[52][23],u_xpb_out[53][23],u_xpb_out[54][23],u_xpb_out[55][23],u_xpb_out[56][23],u_xpb_out[57][23],u_xpb_out[58][23],u_xpb_out[59][23],u_xpb_out[60][23],u_xpb_out[61][23],u_xpb_out[62][23],u_xpb_out[63][23],u_xpb_out[64][23],u_xpb_out[65][23],u_xpb_out[66][23],u_xpb_out[67][23],u_xpb_out[68][23],u_xpb_out[69][23],u_xpb_out[70][23],u_xpb_out[71][23],u_xpb_out[72][23],u_xpb_out[73][23],u_xpb_out[74][23],u_xpb_out[75][23],u_xpb_out[76][23],u_xpb_out[77][23],u_xpb_out[78][23],u_xpb_out[79][23],u_xpb_out[80][23],u_xpb_out[81][23],u_xpb_out[82][23],u_xpb_out[83][23],u_xpb_out[84][23],u_xpb_out[85][23],u_xpb_out[86][23],u_xpb_out[87][23],u_xpb_out[88][23],u_xpb_out[89][23],u_xpb_out[90][23],u_xpb_out[91][23],u_xpb_out[92][23],u_xpb_out[93][23],u_xpb_out[94][23],u_xpb_out[95][23],u_xpb_out[96][23],u_xpb_out[97][23],u_xpb_out[98][23],u_xpb_out[99][23],u_xpb_out[100][23],u_xpb_out[101][23],u_xpb_out[102][23],u_xpb_out[103][23],u_xpb_out[104][23],u_xpb_out[105][23]};

assign col_out_24 = {u_xpb_out[0][24],u_xpb_out[1][24],u_xpb_out[2][24],u_xpb_out[3][24],u_xpb_out[4][24],u_xpb_out[5][24],u_xpb_out[6][24],u_xpb_out[7][24],u_xpb_out[8][24],u_xpb_out[9][24],u_xpb_out[10][24],u_xpb_out[11][24],u_xpb_out[12][24],u_xpb_out[13][24],u_xpb_out[14][24],u_xpb_out[15][24],u_xpb_out[16][24],u_xpb_out[17][24],u_xpb_out[18][24],u_xpb_out[19][24],u_xpb_out[20][24],u_xpb_out[21][24],u_xpb_out[22][24],u_xpb_out[23][24],u_xpb_out[24][24],u_xpb_out[25][24],u_xpb_out[26][24],u_xpb_out[27][24],u_xpb_out[28][24],u_xpb_out[29][24],u_xpb_out[30][24],u_xpb_out[31][24],u_xpb_out[32][24],u_xpb_out[33][24],u_xpb_out[34][24],u_xpb_out[35][24],u_xpb_out[36][24],u_xpb_out[37][24],u_xpb_out[38][24],u_xpb_out[39][24],u_xpb_out[40][24],u_xpb_out[41][24],u_xpb_out[42][24],u_xpb_out[43][24],u_xpb_out[44][24],u_xpb_out[45][24],u_xpb_out[46][24],u_xpb_out[47][24],u_xpb_out[48][24],u_xpb_out[49][24],u_xpb_out[50][24],u_xpb_out[51][24],u_xpb_out[52][24],u_xpb_out[53][24],u_xpb_out[54][24],u_xpb_out[55][24],u_xpb_out[56][24],u_xpb_out[57][24],u_xpb_out[58][24],u_xpb_out[59][24],u_xpb_out[60][24],u_xpb_out[61][24],u_xpb_out[62][24],u_xpb_out[63][24],u_xpb_out[64][24],u_xpb_out[65][24],u_xpb_out[66][24],u_xpb_out[67][24],u_xpb_out[68][24],u_xpb_out[69][24],u_xpb_out[70][24],u_xpb_out[71][24],u_xpb_out[72][24],u_xpb_out[73][24],u_xpb_out[74][24],u_xpb_out[75][24],u_xpb_out[76][24],u_xpb_out[77][24],u_xpb_out[78][24],u_xpb_out[79][24],u_xpb_out[80][24],u_xpb_out[81][24],u_xpb_out[82][24],u_xpb_out[83][24],u_xpb_out[84][24],u_xpb_out[85][24],u_xpb_out[86][24],u_xpb_out[87][24],u_xpb_out[88][24],u_xpb_out[89][24],u_xpb_out[90][24],u_xpb_out[91][24],u_xpb_out[92][24],u_xpb_out[93][24],u_xpb_out[94][24],u_xpb_out[95][24],u_xpb_out[96][24],u_xpb_out[97][24],u_xpb_out[98][24],u_xpb_out[99][24],u_xpb_out[100][24],u_xpb_out[101][24],u_xpb_out[102][24],u_xpb_out[103][24],u_xpb_out[104][24],u_xpb_out[105][24]};

assign col_out_25 = {u_xpb_out[0][25],u_xpb_out[1][25],u_xpb_out[2][25],u_xpb_out[3][25],u_xpb_out[4][25],u_xpb_out[5][25],u_xpb_out[6][25],u_xpb_out[7][25],u_xpb_out[8][25],u_xpb_out[9][25],u_xpb_out[10][25],u_xpb_out[11][25],u_xpb_out[12][25],u_xpb_out[13][25],u_xpb_out[14][25],u_xpb_out[15][25],u_xpb_out[16][25],u_xpb_out[17][25],u_xpb_out[18][25],u_xpb_out[19][25],u_xpb_out[20][25],u_xpb_out[21][25],u_xpb_out[22][25],u_xpb_out[23][25],u_xpb_out[24][25],u_xpb_out[25][25],u_xpb_out[26][25],u_xpb_out[27][25],u_xpb_out[28][25],u_xpb_out[29][25],u_xpb_out[30][25],u_xpb_out[31][25],u_xpb_out[32][25],u_xpb_out[33][25],u_xpb_out[34][25],u_xpb_out[35][25],u_xpb_out[36][25],u_xpb_out[37][25],u_xpb_out[38][25],u_xpb_out[39][25],u_xpb_out[40][25],u_xpb_out[41][25],u_xpb_out[42][25],u_xpb_out[43][25],u_xpb_out[44][25],u_xpb_out[45][25],u_xpb_out[46][25],u_xpb_out[47][25],u_xpb_out[48][25],u_xpb_out[49][25],u_xpb_out[50][25],u_xpb_out[51][25],u_xpb_out[52][25],u_xpb_out[53][25],u_xpb_out[54][25],u_xpb_out[55][25],u_xpb_out[56][25],u_xpb_out[57][25],u_xpb_out[58][25],u_xpb_out[59][25],u_xpb_out[60][25],u_xpb_out[61][25],u_xpb_out[62][25],u_xpb_out[63][25],u_xpb_out[64][25],u_xpb_out[65][25],u_xpb_out[66][25],u_xpb_out[67][25],u_xpb_out[68][25],u_xpb_out[69][25],u_xpb_out[70][25],u_xpb_out[71][25],u_xpb_out[72][25],u_xpb_out[73][25],u_xpb_out[74][25],u_xpb_out[75][25],u_xpb_out[76][25],u_xpb_out[77][25],u_xpb_out[78][25],u_xpb_out[79][25],u_xpb_out[80][25],u_xpb_out[81][25],u_xpb_out[82][25],u_xpb_out[83][25],u_xpb_out[84][25],u_xpb_out[85][25],u_xpb_out[86][25],u_xpb_out[87][25],u_xpb_out[88][25],u_xpb_out[89][25],u_xpb_out[90][25],u_xpb_out[91][25],u_xpb_out[92][25],u_xpb_out[93][25],u_xpb_out[94][25],u_xpb_out[95][25],u_xpb_out[96][25],u_xpb_out[97][25],u_xpb_out[98][25],u_xpb_out[99][25],u_xpb_out[100][25],u_xpb_out[101][25],u_xpb_out[102][25],u_xpb_out[103][25],u_xpb_out[104][25],u_xpb_out[105][25]};

assign col_out_26 = {u_xpb_out[0][26],u_xpb_out[1][26],u_xpb_out[2][26],u_xpb_out[3][26],u_xpb_out[4][26],u_xpb_out[5][26],u_xpb_out[6][26],u_xpb_out[7][26],u_xpb_out[8][26],u_xpb_out[9][26],u_xpb_out[10][26],u_xpb_out[11][26],u_xpb_out[12][26],u_xpb_out[13][26],u_xpb_out[14][26],u_xpb_out[15][26],u_xpb_out[16][26],u_xpb_out[17][26],u_xpb_out[18][26],u_xpb_out[19][26],u_xpb_out[20][26],u_xpb_out[21][26],u_xpb_out[22][26],u_xpb_out[23][26],u_xpb_out[24][26],u_xpb_out[25][26],u_xpb_out[26][26],u_xpb_out[27][26],u_xpb_out[28][26],u_xpb_out[29][26],u_xpb_out[30][26],u_xpb_out[31][26],u_xpb_out[32][26],u_xpb_out[33][26],u_xpb_out[34][26],u_xpb_out[35][26],u_xpb_out[36][26],u_xpb_out[37][26],u_xpb_out[38][26],u_xpb_out[39][26],u_xpb_out[40][26],u_xpb_out[41][26],u_xpb_out[42][26],u_xpb_out[43][26],u_xpb_out[44][26],u_xpb_out[45][26],u_xpb_out[46][26],u_xpb_out[47][26],u_xpb_out[48][26],u_xpb_out[49][26],u_xpb_out[50][26],u_xpb_out[51][26],u_xpb_out[52][26],u_xpb_out[53][26],u_xpb_out[54][26],u_xpb_out[55][26],u_xpb_out[56][26],u_xpb_out[57][26],u_xpb_out[58][26],u_xpb_out[59][26],u_xpb_out[60][26],u_xpb_out[61][26],u_xpb_out[62][26],u_xpb_out[63][26],u_xpb_out[64][26],u_xpb_out[65][26],u_xpb_out[66][26],u_xpb_out[67][26],u_xpb_out[68][26],u_xpb_out[69][26],u_xpb_out[70][26],u_xpb_out[71][26],u_xpb_out[72][26],u_xpb_out[73][26],u_xpb_out[74][26],u_xpb_out[75][26],u_xpb_out[76][26],u_xpb_out[77][26],u_xpb_out[78][26],u_xpb_out[79][26],u_xpb_out[80][26],u_xpb_out[81][26],u_xpb_out[82][26],u_xpb_out[83][26],u_xpb_out[84][26],u_xpb_out[85][26],u_xpb_out[86][26],u_xpb_out[87][26],u_xpb_out[88][26],u_xpb_out[89][26],u_xpb_out[90][26],u_xpb_out[91][26],u_xpb_out[92][26],u_xpb_out[93][26],u_xpb_out[94][26],u_xpb_out[95][26],u_xpb_out[96][26],u_xpb_out[97][26],u_xpb_out[98][26],u_xpb_out[99][26],u_xpb_out[100][26],u_xpb_out[101][26],u_xpb_out[102][26],u_xpb_out[103][26],u_xpb_out[104][26],u_xpb_out[105][26]};

assign col_out_27 = {u_xpb_out[0][27],u_xpb_out[1][27],u_xpb_out[2][27],u_xpb_out[3][27],u_xpb_out[4][27],u_xpb_out[5][27],u_xpb_out[6][27],u_xpb_out[7][27],u_xpb_out[8][27],u_xpb_out[9][27],u_xpb_out[10][27],u_xpb_out[11][27],u_xpb_out[12][27],u_xpb_out[13][27],u_xpb_out[14][27],u_xpb_out[15][27],u_xpb_out[16][27],u_xpb_out[17][27],u_xpb_out[18][27],u_xpb_out[19][27],u_xpb_out[20][27],u_xpb_out[21][27],u_xpb_out[22][27],u_xpb_out[23][27],u_xpb_out[24][27],u_xpb_out[25][27],u_xpb_out[26][27],u_xpb_out[27][27],u_xpb_out[28][27],u_xpb_out[29][27],u_xpb_out[30][27],u_xpb_out[31][27],u_xpb_out[32][27],u_xpb_out[33][27],u_xpb_out[34][27],u_xpb_out[35][27],u_xpb_out[36][27],u_xpb_out[37][27],u_xpb_out[38][27],u_xpb_out[39][27],u_xpb_out[40][27],u_xpb_out[41][27],u_xpb_out[42][27],u_xpb_out[43][27],u_xpb_out[44][27],u_xpb_out[45][27],u_xpb_out[46][27],u_xpb_out[47][27],u_xpb_out[48][27],u_xpb_out[49][27],u_xpb_out[50][27],u_xpb_out[51][27],u_xpb_out[52][27],u_xpb_out[53][27],u_xpb_out[54][27],u_xpb_out[55][27],u_xpb_out[56][27],u_xpb_out[57][27],u_xpb_out[58][27],u_xpb_out[59][27],u_xpb_out[60][27],u_xpb_out[61][27],u_xpb_out[62][27],u_xpb_out[63][27],u_xpb_out[64][27],u_xpb_out[65][27],u_xpb_out[66][27],u_xpb_out[67][27],u_xpb_out[68][27],u_xpb_out[69][27],u_xpb_out[70][27],u_xpb_out[71][27],u_xpb_out[72][27],u_xpb_out[73][27],u_xpb_out[74][27],u_xpb_out[75][27],u_xpb_out[76][27],u_xpb_out[77][27],u_xpb_out[78][27],u_xpb_out[79][27],u_xpb_out[80][27],u_xpb_out[81][27],u_xpb_out[82][27],u_xpb_out[83][27],u_xpb_out[84][27],u_xpb_out[85][27],u_xpb_out[86][27],u_xpb_out[87][27],u_xpb_out[88][27],u_xpb_out[89][27],u_xpb_out[90][27],u_xpb_out[91][27],u_xpb_out[92][27],u_xpb_out[93][27],u_xpb_out[94][27],u_xpb_out[95][27],u_xpb_out[96][27],u_xpb_out[97][27],u_xpb_out[98][27],u_xpb_out[99][27],u_xpb_out[100][27],u_xpb_out[101][27],u_xpb_out[102][27],u_xpb_out[103][27],u_xpb_out[104][27],u_xpb_out[105][27]};

assign col_out_28 = {u_xpb_out[0][28],u_xpb_out[1][28],u_xpb_out[2][28],u_xpb_out[3][28],u_xpb_out[4][28],u_xpb_out[5][28],u_xpb_out[6][28],u_xpb_out[7][28],u_xpb_out[8][28],u_xpb_out[9][28],u_xpb_out[10][28],u_xpb_out[11][28],u_xpb_out[12][28],u_xpb_out[13][28],u_xpb_out[14][28],u_xpb_out[15][28],u_xpb_out[16][28],u_xpb_out[17][28],u_xpb_out[18][28],u_xpb_out[19][28],u_xpb_out[20][28],u_xpb_out[21][28],u_xpb_out[22][28],u_xpb_out[23][28],u_xpb_out[24][28],u_xpb_out[25][28],u_xpb_out[26][28],u_xpb_out[27][28],u_xpb_out[28][28],u_xpb_out[29][28],u_xpb_out[30][28],u_xpb_out[31][28],u_xpb_out[32][28],u_xpb_out[33][28],u_xpb_out[34][28],u_xpb_out[35][28],u_xpb_out[36][28],u_xpb_out[37][28],u_xpb_out[38][28],u_xpb_out[39][28],u_xpb_out[40][28],u_xpb_out[41][28],u_xpb_out[42][28],u_xpb_out[43][28],u_xpb_out[44][28],u_xpb_out[45][28],u_xpb_out[46][28],u_xpb_out[47][28],u_xpb_out[48][28],u_xpb_out[49][28],u_xpb_out[50][28],u_xpb_out[51][28],u_xpb_out[52][28],u_xpb_out[53][28],u_xpb_out[54][28],u_xpb_out[55][28],u_xpb_out[56][28],u_xpb_out[57][28],u_xpb_out[58][28],u_xpb_out[59][28],u_xpb_out[60][28],u_xpb_out[61][28],u_xpb_out[62][28],u_xpb_out[63][28],u_xpb_out[64][28],u_xpb_out[65][28],u_xpb_out[66][28],u_xpb_out[67][28],u_xpb_out[68][28],u_xpb_out[69][28],u_xpb_out[70][28],u_xpb_out[71][28],u_xpb_out[72][28],u_xpb_out[73][28],u_xpb_out[74][28],u_xpb_out[75][28],u_xpb_out[76][28],u_xpb_out[77][28],u_xpb_out[78][28],u_xpb_out[79][28],u_xpb_out[80][28],u_xpb_out[81][28],u_xpb_out[82][28],u_xpb_out[83][28],u_xpb_out[84][28],u_xpb_out[85][28],u_xpb_out[86][28],u_xpb_out[87][28],u_xpb_out[88][28],u_xpb_out[89][28],u_xpb_out[90][28],u_xpb_out[91][28],u_xpb_out[92][28],u_xpb_out[93][28],u_xpb_out[94][28],u_xpb_out[95][28],u_xpb_out[96][28],u_xpb_out[97][28],u_xpb_out[98][28],u_xpb_out[99][28],u_xpb_out[100][28],u_xpb_out[101][28],u_xpb_out[102][28],u_xpb_out[103][28],u_xpb_out[104][28],u_xpb_out[105][28]};

assign col_out_29 = {u_xpb_out[0][29],u_xpb_out[1][29],u_xpb_out[2][29],u_xpb_out[3][29],u_xpb_out[4][29],u_xpb_out[5][29],u_xpb_out[6][29],u_xpb_out[7][29],u_xpb_out[8][29],u_xpb_out[9][29],u_xpb_out[10][29],u_xpb_out[11][29],u_xpb_out[12][29],u_xpb_out[13][29],u_xpb_out[14][29],u_xpb_out[15][29],u_xpb_out[16][29],u_xpb_out[17][29],u_xpb_out[18][29],u_xpb_out[19][29],u_xpb_out[20][29],u_xpb_out[21][29],u_xpb_out[22][29],u_xpb_out[23][29],u_xpb_out[24][29],u_xpb_out[25][29],u_xpb_out[26][29],u_xpb_out[27][29],u_xpb_out[28][29],u_xpb_out[29][29],u_xpb_out[30][29],u_xpb_out[31][29],u_xpb_out[32][29],u_xpb_out[33][29],u_xpb_out[34][29],u_xpb_out[35][29],u_xpb_out[36][29],u_xpb_out[37][29],u_xpb_out[38][29],u_xpb_out[39][29],u_xpb_out[40][29],u_xpb_out[41][29],u_xpb_out[42][29],u_xpb_out[43][29],u_xpb_out[44][29],u_xpb_out[45][29],u_xpb_out[46][29],u_xpb_out[47][29],u_xpb_out[48][29],u_xpb_out[49][29],u_xpb_out[50][29],u_xpb_out[51][29],u_xpb_out[52][29],u_xpb_out[53][29],u_xpb_out[54][29],u_xpb_out[55][29],u_xpb_out[56][29],u_xpb_out[57][29],u_xpb_out[58][29],u_xpb_out[59][29],u_xpb_out[60][29],u_xpb_out[61][29],u_xpb_out[62][29],u_xpb_out[63][29],u_xpb_out[64][29],u_xpb_out[65][29],u_xpb_out[66][29],u_xpb_out[67][29],u_xpb_out[68][29],u_xpb_out[69][29],u_xpb_out[70][29],u_xpb_out[71][29],u_xpb_out[72][29],u_xpb_out[73][29],u_xpb_out[74][29],u_xpb_out[75][29],u_xpb_out[76][29],u_xpb_out[77][29],u_xpb_out[78][29],u_xpb_out[79][29],u_xpb_out[80][29],u_xpb_out[81][29],u_xpb_out[82][29],u_xpb_out[83][29],u_xpb_out[84][29],u_xpb_out[85][29],u_xpb_out[86][29],u_xpb_out[87][29],u_xpb_out[88][29],u_xpb_out[89][29],u_xpb_out[90][29],u_xpb_out[91][29],u_xpb_out[92][29],u_xpb_out[93][29],u_xpb_out[94][29],u_xpb_out[95][29],u_xpb_out[96][29],u_xpb_out[97][29],u_xpb_out[98][29],u_xpb_out[99][29],u_xpb_out[100][29],u_xpb_out[101][29],u_xpb_out[102][29],u_xpb_out[103][29],u_xpb_out[104][29],u_xpb_out[105][29]};

assign col_out_30 = {u_xpb_out[0][30],u_xpb_out[1][30],u_xpb_out[2][30],u_xpb_out[3][30],u_xpb_out[4][30],u_xpb_out[5][30],u_xpb_out[6][30],u_xpb_out[7][30],u_xpb_out[8][30],u_xpb_out[9][30],u_xpb_out[10][30],u_xpb_out[11][30],u_xpb_out[12][30],u_xpb_out[13][30],u_xpb_out[14][30],u_xpb_out[15][30],u_xpb_out[16][30],u_xpb_out[17][30],u_xpb_out[18][30],u_xpb_out[19][30],u_xpb_out[20][30],u_xpb_out[21][30],u_xpb_out[22][30],u_xpb_out[23][30],u_xpb_out[24][30],u_xpb_out[25][30],u_xpb_out[26][30],u_xpb_out[27][30],u_xpb_out[28][30],u_xpb_out[29][30],u_xpb_out[30][30],u_xpb_out[31][30],u_xpb_out[32][30],u_xpb_out[33][30],u_xpb_out[34][30],u_xpb_out[35][30],u_xpb_out[36][30],u_xpb_out[37][30],u_xpb_out[38][30],u_xpb_out[39][30],u_xpb_out[40][30],u_xpb_out[41][30],u_xpb_out[42][30],u_xpb_out[43][30],u_xpb_out[44][30],u_xpb_out[45][30],u_xpb_out[46][30],u_xpb_out[47][30],u_xpb_out[48][30],u_xpb_out[49][30],u_xpb_out[50][30],u_xpb_out[51][30],u_xpb_out[52][30],u_xpb_out[53][30],u_xpb_out[54][30],u_xpb_out[55][30],u_xpb_out[56][30],u_xpb_out[57][30],u_xpb_out[58][30],u_xpb_out[59][30],u_xpb_out[60][30],u_xpb_out[61][30],u_xpb_out[62][30],u_xpb_out[63][30],u_xpb_out[64][30],u_xpb_out[65][30],u_xpb_out[66][30],u_xpb_out[67][30],u_xpb_out[68][30],u_xpb_out[69][30],u_xpb_out[70][30],u_xpb_out[71][30],u_xpb_out[72][30],u_xpb_out[73][30],u_xpb_out[74][30],u_xpb_out[75][30],u_xpb_out[76][30],u_xpb_out[77][30],u_xpb_out[78][30],u_xpb_out[79][30],u_xpb_out[80][30],u_xpb_out[81][30],u_xpb_out[82][30],u_xpb_out[83][30],u_xpb_out[84][30],u_xpb_out[85][30],u_xpb_out[86][30],u_xpb_out[87][30],u_xpb_out[88][30],u_xpb_out[89][30],u_xpb_out[90][30],u_xpb_out[91][30],u_xpb_out[92][30],u_xpb_out[93][30],u_xpb_out[94][30],u_xpb_out[95][30],u_xpb_out[96][30],u_xpb_out[97][30],u_xpb_out[98][30],u_xpb_out[99][30],u_xpb_out[100][30],u_xpb_out[101][30],u_xpb_out[102][30],u_xpb_out[103][30],u_xpb_out[104][30],u_xpb_out[105][30]};

assign col_out_31 = {u_xpb_out[0][31],u_xpb_out[1][31],u_xpb_out[2][31],u_xpb_out[3][31],u_xpb_out[4][31],u_xpb_out[5][31],u_xpb_out[6][31],u_xpb_out[7][31],u_xpb_out[8][31],u_xpb_out[9][31],u_xpb_out[10][31],u_xpb_out[11][31],u_xpb_out[12][31],u_xpb_out[13][31],u_xpb_out[14][31],u_xpb_out[15][31],u_xpb_out[16][31],u_xpb_out[17][31],u_xpb_out[18][31],u_xpb_out[19][31],u_xpb_out[20][31],u_xpb_out[21][31],u_xpb_out[22][31],u_xpb_out[23][31],u_xpb_out[24][31],u_xpb_out[25][31],u_xpb_out[26][31],u_xpb_out[27][31],u_xpb_out[28][31],u_xpb_out[29][31],u_xpb_out[30][31],u_xpb_out[31][31],u_xpb_out[32][31],u_xpb_out[33][31],u_xpb_out[34][31],u_xpb_out[35][31],u_xpb_out[36][31],u_xpb_out[37][31],u_xpb_out[38][31],u_xpb_out[39][31],u_xpb_out[40][31],u_xpb_out[41][31],u_xpb_out[42][31],u_xpb_out[43][31],u_xpb_out[44][31],u_xpb_out[45][31],u_xpb_out[46][31],u_xpb_out[47][31],u_xpb_out[48][31],u_xpb_out[49][31],u_xpb_out[50][31],u_xpb_out[51][31],u_xpb_out[52][31],u_xpb_out[53][31],u_xpb_out[54][31],u_xpb_out[55][31],u_xpb_out[56][31],u_xpb_out[57][31],u_xpb_out[58][31],u_xpb_out[59][31],u_xpb_out[60][31],u_xpb_out[61][31],u_xpb_out[62][31],u_xpb_out[63][31],u_xpb_out[64][31],u_xpb_out[65][31],u_xpb_out[66][31],u_xpb_out[67][31],u_xpb_out[68][31],u_xpb_out[69][31],u_xpb_out[70][31],u_xpb_out[71][31],u_xpb_out[72][31],u_xpb_out[73][31],u_xpb_out[74][31],u_xpb_out[75][31],u_xpb_out[76][31],u_xpb_out[77][31],u_xpb_out[78][31],u_xpb_out[79][31],u_xpb_out[80][31],u_xpb_out[81][31],u_xpb_out[82][31],u_xpb_out[83][31],u_xpb_out[84][31],u_xpb_out[85][31],u_xpb_out[86][31],u_xpb_out[87][31],u_xpb_out[88][31],u_xpb_out[89][31],u_xpb_out[90][31],u_xpb_out[91][31],u_xpb_out[92][31],u_xpb_out[93][31],u_xpb_out[94][31],u_xpb_out[95][31],u_xpb_out[96][31],u_xpb_out[97][31],u_xpb_out[98][31],u_xpb_out[99][31],u_xpb_out[100][31],u_xpb_out[101][31],u_xpb_out[102][31],u_xpb_out[103][31],u_xpb_out[104][31],u_xpb_out[105][31]};

assign col_out_32 = {u_xpb_out[0][32],u_xpb_out[1][32],u_xpb_out[2][32],u_xpb_out[3][32],u_xpb_out[4][32],u_xpb_out[5][32],u_xpb_out[6][32],u_xpb_out[7][32],u_xpb_out[8][32],u_xpb_out[9][32],u_xpb_out[10][32],u_xpb_out[11][32],u_xpb_out[12][32],u_xpb_out[13][32],u_xpb_out[14][32],u_xpb_out[15][32],u_xpb_out[16][32],u_xpb_out[17][32],u_xpb_out[18][32],u_xpb_out[19][32],u_xpb_out[20][32],u_xpb_out[21][32],u_xpb_out[22][32],u_xpb_out[23][32],u_xpb_out[24][32],u_xpb_out[25][32],u_xpb_out[26][32],u_xpb_out[27][32],u_xpb_out[28][32],u_xpb_out[29][32],u_xpb_out[30][32],u_xpb_out[31][32],u_xpb_out[32][32],u_xpb_out[33][32],u_xpb_out[34][32],u_xpb_out[35][32],u_xpb_out[36][32],u_xpb_out[37][32],u_xpb_out[38][32],u_xpb_out[39][32],u_xpb_out[40][32],u_xpb_out[41][32],u_xpb_out[42][32],u_xpb_out[43][32],u_xpb_out[44][32],u_xpb_out[45][32],u_xpb_out[46][32],u_xpb_out[47][32],u_xpb_out[48][32],u_xpb_out[49][32],u_xpb_out[50][32],u_xpb_out[51][32],u_xpb_out[52][32],u_xpb_out[53][32],u_xpb_out[54][32],u_xpb_out[55][32],u_xpb_out[56][32],u_xpb_out[57][32],u_xpb_out[58][32],u_xpb_out[59][32],u_xpb_out[60][32],u_xpb_out[61][32],u_xpb_out[62][32],u_xpb_out[63][32],u_xpb_out[64][32],u_xpb_out[65][32],u_xpb_out[66][32],u_xpb_out[67][32],u_xpb_out[68][32],u_xpb_out[69][32],u_xpb_out[70][32],u_xpb_out[71][32],u_xpb_out[72][32],u_xpb_out[73][32],u_xpb_out[74][32],u_xpb_out[75][32],u_xpb_out[76][32],u_xpb_out[77][32],u_xpb_out[78][32],u_xpb_out[79][32],u_xpb_out[80][32],u_xpb_out[81][32],u_xpb_out[82][32],u_xpb_out[83][32],u_xpb_out[84][32],u_xpb_out[85][32],u_xpb_out[86][32],u_xpb_out[87][32],u_xpb_out[88][32],u_xpb_out[89][32],u_xpb_out[90][32],u_xpb_out[91][32],u_xpb_out[92][32],u_xpb_out[93][32],u_xpb_out[94][32],u_xpb_out[95][32],u_xpb_out[96][32],u_xpb_out[97][32],u_xpb_out[98][32],u_xpb_out[99][32],u_xpb_out[100][32],u_xpb_out[101][32],u_xpb_out[102][32],u_xpb_out[103][32],u_xpb_out[104][32],u_xpb_out[105][32]};

assign col_out_33 = {u_xpb_out[0][33],u_xpb_out[1][33],u_xpb_out[2][33],u_xpb_out[3][33],u_xpb_out[4][33],u_xpb_out[5][33],u_xpb_out[6][33],u_xpb_out[7][33],u_xpb_out[8][33],u_xpb_out[9][33],u_xpb_out[10][33],u_xpb_out[11][33],u_xpb_out[12][33],u_xpb_out[13][33],u_xpb_out[14][33],u_xpb_out[15][33],u_xpb_out[16][33],u_xpb_out[17][33],u_xpb_out[18][33],u_xpb_out[19][33],u_xpb_out[20][33],u_xpb_out[21][33],u_xpb_out[22][33],u_xpb_out[23][33],u_xpb_out[24][33],u_xpb_out[25][33],u_xpb_out[26][33],u_xpb_out[27][33],u_xpb_out[28][33],u_xpb_out[29][33],u_xpb_out[30][33],u_xpb_out[31][33],u_xpb_out[32][33],u_xpb_out[33][33],u_xpb_out[34][33],u_xpb_out[35][33],u_xpb_out[36][33],u_xpb_out[37][33],u_xpb_out[38][33],u_xpb_out[39][33],u_xpb_out[40][33],u_xpb_out[41][33],u_xpb_out[42][33],u_xpb_out[43][33],u_xpb_out[44][33],u_xpb_out[45][33],u_xpb_out[46][33],u_xpb_out[47][33],u_xpb_out[48][33],u_xpb_out[49][33],u_xpb_out[50][33],u_xpb_out[51][33],u_xpb_out[52][33],u_xpb_out[53][33],u_xpb_out[54][33],u_xpb_out[55][33],u_xpb_out[56][33],u_xpb_out[57][33],u_xpb_out[58][33],u_xpb_out[59][33],u_xpb_out[60][33],u_xpb_out[61][33],u_xpb_out[62][33],u_xpb_out[63][33],u_xpb_out[64][33],u_xpb_out[65][33],u_xpb_out[66][33],u_xpb_out[67][33],u_xpb_out[68][33],u_xpb_out[69][33],u_xpb_out[70][33],u_xpb_out[71][33],u_xpb_out[72][33],u_xpb_out[73][33],u_xpb_out[74][33],u_xpb_out[75][33],u_xpb_out[76][33],u_xpb_out[77][33],u_xpb_out[78][33],u_xpb_out[79][33],u_xpb_out[80][33],u_xpb_out[81][33],u_xpb_out[82][33],u_xpb_out[83][33],u_xpb_out[84][33],u_xpb_out[85][33],u_xpb_out[86][33],u_xpb_out[87][33],u_xpb_out[88][33],u_xpb_out[89][33],u_xpb_out[90][33],u_xpb_out[91][33],u_xpb_out[92][33],u_xpb_out[93][33],u_xpb_out[94][33],u_xpb_out[95][33],u_xpb_out[96][33],u_xpb_out[97][33],u_xpb_out[98][33],u_xpb_out[99][33],u_xpb_out[100][33],u_xpb_out[101][33],u_xpb_out[102][33],u_xpb_out[103][33],u_xpb_out[104][33],u_xpb_out[105][33]};

assign col_out_34 = {u_xpb_out[0][34],u_xpb_out[1][34],u_xpb_out[2][34],u_xpb_out[3][34],u_xpb_out[4][34],u_xpb_out[5][34],u_xpb_out[6][34],u_xpb_out[7][34],u_xpb_out[8][34],u_xpb_out[9][34],u_xpb_out[10][34],u_xpb_out[11][34],u_xpb_out[12][34],u_xpb_out[13][34],u_xpb_out[14][34],u_xpb_out[15][34],u_xpb_out[16][34],u_xpb_out[17][34],u_xpb_out[18][34],u_xpb_out[19][34],u_xpb_out[20][34],u_xpb_out[21][34],u_xpb_out[22][34],u_xpb_out[23][34],u_xpb_out[24][34],u_xpb_out[25][34],u_xpb_out[26][34],u_xpb_out[27][34],u_xpb_out[28][34],u_xpb_out[29][34],u_xpb_out[30][34],u_xpb_out[31][34],u_xpb_out[32][34],u_xpb_out[33][34],u_xpb_out[34][34],u_xpb_out[35][34],u_xpb_out[36][34],u_xpb_out[37][34],u_xpb_out[38][34],u_xpb_out[39][34],u_xpb_out[40][34],u_xpb_out[41][34],u_xpb_out[42][34],u_xpb_out[43][34],u_xpb_out[44][34],u_xpb_out[45][34],u_xpb_out[46][34],u_xpb_out[47][34],u_xpb_out[48][34],u_xpb_out[49][34],u_xpb_out[50][34],u_xpb_out[51][34],u_xpb_out[52][34],u_xpb_out[53][34],u_xpb_out[54][34],u_xpb_out[55][34],u_xpb_out[56][34],u_xpb_out[57][34],u_xpb_out[58][34],u_xpb_out[59][34],u_xpb_out[60][34],u_xpb_out[61][34],u_xpb_out[62][34],u_xpb_out[63][34],u_xpb_out[64][34],u_xpb_out[65][34],u_xpb_out[66][34],u_xpb_out[67][34],u_xpb_out[68][34],u_xpb_out[69][34],u_xpb_out[70][34],u_xpb_out[71][34],u_xpb_out[72][34],u_xpb_out[73][34],u_xpb_out[74][34],u_xpb_out[75][34],u_xpb_out[76][34],u_xpb_out[77][34],u_xpb_out[78][34],u_xpb_out[79][34],u_xpb_out[80][34],u_xpb_out[81][34],u_xpb_out[82][34],u_xpb_out[83][34],u_xpb_out[84][34],u_xpb_out[85][34],u_xpb_out[86][34],u_xpb_out[87][34],u_xpb_out[88][34],u_xpb_out[89][34],u_xpb_out[90][34],u_xpb_out[91][34],u_xpb_out[92][34],u_xpb_out[93][34],u_xpb_out[94][34],u_xpb_out[95][34],u_xpb_out[96][34],u_xpb_out[97][34],u_xpb_out[98][34],u_xpb_out[99][34],u_xpb_out[100][34],u_xpb_out[101][34],u_xpb_out[102][34],u_xpb_out[103][34],u_xpb_out[104][34],u_xpb_out[105][34]};

assign col_out_35 = {u_xpb_out[0][35],u_xpb_out[1][35],u_xpb_out[2][35],u_xpb_out[3][35],u_xpb_out[4][35],u_xpb_out[5][35],u_xpb_out[6][35],u_xpb_out[7][35],u_xpb_out[8][35],u_xpb_out[9][35],u_xpb_out[10][35],u_xpb_out[11][35],u_xpb_out[12][35],u_xpb_out[13][35],u_xpb_out[14][35],u_xpb_out[15][35],u_xpb_out[16][35],u_xpb_out[17][35],u_xpb_out[18][35],u_xpb_out[19][35],u_xpb_out[20][35],u_xpb_out[21][35],u_xpb_out[22][35],u_xpb_out[23][35],u_xpb_out[24][35],u_xpb_out[25][35],u_xpb_out[26][35],u_xpb_out[27][35],u_xpb_out[28][35],u_xpb_out[29][35],u_xpb_out[30][35],u_xpb_out[31][35],u_xpb_out[32][35],u_xpb_out[33][35],u_xpb_out[34][35],u_xpb_out[35][35],u_xpb_out[36][35],u_xpb_out[37][35],u_xpb_out[38][35],u_xpb_out[39][35],u_xpb_out[40][35],u_xpb_out[41][35],u_xpb_out[42][35],u_xpb_out[43][35],u_xpb_out[44][35],u_xpb_out[45][35],u_xpb_out[46][35],u_xpb_out[47][35],u_xpb_out[48][35],u_xpb_out[49][35],u_xpb_out[50][35],u_xpb_out[51][35],u_xpb_out[52][35],u_xpb_out[53][35],u_xpb_out[54][35],u_xpb_out[55][35],u_xpb_out[56][35],u_xpb_out[57][35],u_xpb_out[58][35],u_xpb_out[59][35],u_xpb_out[60][35],u_xpb_out[61][35],u_xpb_out[62][35],u_xpb_out[63][35],u_xpb_out[64][35],u_xpb_out[65][35],u_xpb_out[66][35],u_xpb_out[67][35],u_xpb_out[68][35],u_xpb_out[69][35],u_xpb_out[70][35],u_xpb_out[71][35],u_xpb_out[72][35],u_xpb_out[73][35],u_xpb_out[74][35],u_xpb_out[75][35],u_xpb_out[76][35],u_xpb_out[77][35],u_xpb_out[78][35],u_xpb_out[79][35],u_xpb_out[80][35],u_xpb_out[81][35],u_xpb_out[82][35],u_xpb_out[83][35],u_xpb_out[84][35],u_xpb_out[85][35],u_xpb_out[86][35],u_xpb_out[87][35],u_xpb_out[88][35],u_xpb_out[89][35],u_xpb_out[90][35],u_xpb_out[91][35],u_xpb_out[92][35],u_xpb_out[93][35],u_xpb_out[94][35],u_xpb_out[95][35],u_xpb_out[96][35],u_xpb_out[97][35],u_xpb_out[98][35],u_xpb_out[99][35],u_xpb_out[100][35],u_xpb_out[101][35],u_xpb_out[102][35],u_xpb_out[103][35],u_xpb_out[104][35],u_xpb_out[105][35]};

assign col_out_36 = {u_xpb_out[0][36],u_xpb_out[1][36],u_xpb_out[2][36],u_xpb_out[3][36],u_xpb_out[4][36],u_xpb_out[5][36],u_xpb_out[6][36],u_xpb_out[7][36],u_xpb_out[8][36],u_xpb_out[9][36],u_xpb_out[10][36],u_xpb_out[11][36],u_xpb_out[12][36],u_xpb_out[13][36],u_xpb_out[14][36],u_xpb_out[15][36],u_xpb_out[16][36],u_xpb_out[17][36],u_xpb_out[18][36],u_xpb_out[19][36],u_xpb_out[20][36],u_xpb_out[21][36],u_xpb_out[22][36],u_xpb_out[23][36],u_xpb_out[24][36],u_xpb_out[25][36],u_xpb_out[26][36],u_xpb_out[27][36],u_xpb_out[28][36],u_xpb_out[29][36],u_xpb_out[30][36],u_xpb_out[31][36],u_xpb_out[32][36],u_xpb_out[33][36],u_xpb_out[34][36],u_xpb_out[35][36],u_xpb_out[36][36],u_xpb_out[37][36],u_xpb_out[38][36],u_xpb_out[39][36],u_xpb_out[40][36],u_xpb_out[41][36],u_xpb_out[42][36],u_xpb_out[43][36],u_xpb_out[44][36],u_xpb_out[45][36],u_xpb_out[46][36],u_xpb_out[47][36],u_xpb_out[48][36],u_xpb_out[49][36],u_xpb_out[50][36],u_xpb_out[51][36],u_xpb_out[52][36],u_xpb_out[53][36],u_xpb_out[54][36],u_xpb_out[55][36],u_xpb_out[56][36],u_xpb_out[57][36],u_xpb_out[58][36],u_xpb_out[59][36],u_xpb_out[60][36],u_xpb_out[61][36],u_xpb_out[62][36],u_xpb_out[63][36],u_xpb_out[64][36],u_xpb_out[65][36],u_xpb_out[66][36],u_xpb_out[67][36],u_xpb_out[68][36],u_xpb_out[69][36],u_xpb_out[70][36],u_xpb_out[71][36],u_xpb_out[72][36],u_xpb_out[73][36],u_xpb_out[74][36],u_xpb_out[75][36],u_xpb_out[76][36],u_xpb_out[77][36],u_xpb_out[78][36],u_xpb_out[79][36],u_xpb_out[80][36],u_xpb_out[81][36],u_xpb_out[82][36],u_xpb_out[83][36],u_xpb_out[84][36],u_xpb_out[85][36],u_xpb_out[86][36],u_xpb_out[87][36],u_xpb_out[88][36],u_xpb_out[89][36],u_xpb_out[90][36],u_xpb_out[91][36],u_xpb_out[92][36],u_xpb_out[93][36],u_xpb_out[94][36],u_xpb_out[95][36],u_xpb_out[96][36],u_xpb_out[97][36],u_xpb_out[98][36],u_xpb_out[99][36],u_xpb_out[100][36],u_xpb_out[101][36],u_xpb_out[102][36],u_xpb_out[103][36],u_xpb_out[104][36],u_xpb_out[105][36]};

assign col_out_37 = {u_xpb_out[0][37],u_xpb_out[1][37],u_xpb_out[2][37],u_xpb_out[3][37],u_xpb_out[4][37],u_xpb_out[5][37],u_xpb_out[6][37],u_xpb_out[7][37],u_xpb_out[8][37],u_xpb_out[9][37],u_xpb_out[10][37],u_xpb_out[11][37],u_xpb_out[12][37],u_xpb_out[13][37],u_xpb_out[14][37],u_xpb_out[15][37],u_xpb_out[16][37],u_xpb_out[17][37],u_xpb_out[18][37],u_xpb_out[19][37],u_xpb_out[20][37],u_xpb_out[21][37],u_xpb_out[22][37],u_xpb_out[23][37],u_xpb_out[24][37],u_xpb_out[25][37],u_xpb_out[26][37],u_xpb_out[27][37],u_xpb_out[28][37],u_xpb_out[29][37],u_xpb_out[30][37],u_xpb_out[31][37],u_xpb_out[32][37],u_xpb_out[33][37],u_xpb_out[34][37],u_xpb_out[35][37],u_xpb_out[36][37],u_xpb_out[37][37],u_xpb_out[38][37],u_xpb_out[39][37],u_xpb_out[40][37],u_xpb_out[41][37],u_xpb_out[42][37],u_xpb_out[43][37],u_xpb_out[44][37],u_xpb_out[45][37],u_xpb_out[46][37],u_xpb_out[47][37],u_xpb_out[48][37],u_xpb_out[49][37],u_xpb_out[50][37],u_xpb_out[51][37],u_xpb_out[52][37],u_xpb_out[53][37],u_xpb_out[54][37],u_xpb_out[55][37],u_xpb_out[56][37],u_xpb_out[57][37],u_xpb_out[58][37],u_xpb_out[59][37],u_xpb_out[60][37],u_xpb_out[61][37],u_xpb_out[62][37],u_xpb_out[63][37],u_xpb_out[64][37],u_xpb_out[65][37],u_xpb_out[66][37],u_xpb_out[67][37],u_xpb_out[68][37],u_xpb_out[69][37],u_xpb_out[70][37],u_xpb_out[71][37],u_xpb_out[72][37],u_xpb_out[73][37],u_xpb_out[74][37],u_xpb_out[75][37],u_xpb_out[76][37],u_xpb_out[77][37],u_xpb_out[78][37],u_xpb_out[79][37],u_xpb_out[80][37],u_xpb_out[81][37],u_xpb_out[82][37],u_xpb_out[83][37],u_xpb_out[84][37],u_xpb_out[85][37],u_xpb_out[86][37],u_xpb_out[87][37],u_xpb_out[88][37],u_xpb_out[89][37],u_xpb_out[90][37],u_xpb_out[91][37],u_xpb_out[92][37],u_xpb_out[93][37],u_xpb_out[94][37],u_xpb_out[95][37],u_xpb_out[96][37],u_xpb_out[97][37],u_xpb_out[98][37],u_xpb_out[99][37],u_xpb_out[100][37],u_xpb_out[101][37],u_xpb_out[102][37],u_xpb_out[103][37],u_xpb_out[104][37],u_xpb_out[105][37]};

assign col_out_38 = {u_xpb_out[0][38],u_xpb_out[1][38],u_xpb_out[2][38],u_xpb_out[3][38],u_xpb_out[4][38],u_xpb_out[5][38],u_xpb_out[6][38],u_xpb_out[7][38],u_xpb_out[8][38],u_xpb_out[9][38],u_xpb_out[10][38],u_xpb_out[11][38],u_xpb_out[12][38],u_xpb_out[13][38],u_xpb_out[14][38],u_xpb_out[15][38],u_xpb_out[16][38],u_xpb_out[17][38],u_xpb_out[18][38],u_xpb_out[19][38],u_xpb_out[20][38],u_xpb_out[21][38],u_xpb_out[22][38],u_xpb_out[23][38],u_xpb_out[24][38],u_xpb_out[25][38],u_xpb_out[26][38],u_xpb_out[27][38],u_xpb_out[28][38],u_xpb_out[29][38],u_xpb_out[30][38],u_xpb_out[31][38],u_xpb_out[32][38],u_xpb_out[33][38],u_xpb_out[34][38],u_xpb_out[35][38],u_xpb_out[36][38],u_xpb_out[37][38],u_xpb_out[38][38],u_xpb_out[39][38],u_xpb_out[40][38],u_xpb_out[41][38],u_xpb_out[42][38],u_xpb_out[43][38],u_xpb_out[44][38],u_xpb_out[45][38],u_xpb_out[46][38],u_xpb_out[47][38],u_xpb_out[48][38],u_xpb_out[49][38],u_xpb_out[50][38],u_xpb_out[51][38],u_xpb_out[52][38],u_xpb_out[53][38],u_xpb_out[54][38],u_xpb_out[55][38],u_xpb_out[56][38],u_xpb_out[57][38],u_xpb_out[58][38],u_xpb_out[59][38],u_xpb_out[60][38],u_xpb_out[61][38],u_xpb_out[62][38],u_xpb_out[63][38],u_xpb_out[64][38],u_xpb_out[65][38],u_xpb_out[66][38],u_xpb_out[67][38],u_xpb_out[68][38],u_xpb_out[69][38],u_xpb_out[70][38],u_xpb_out[71][38],u_xpb_out[72][38],u_xpb_out[73][38],u_xpb_out[74][38],u_xpb_out[75][38],u_xpb_out[76][38],u_xpb_out[77][38],u_xpb_out[78][38],u_xpb_out[79][38],u_xpb_out[80][38],u_xpb_out[81][38],u_xpb_out[82][38],u_xpb_out[83][38],u_xpb_out[84][38],u_xpb_out[85][38],u_xpb_out[86][38],u_xpb_out[87][38],u_xpb_out[88][38],u_xpb_out[89][38],u_xpb_out[90][38],u_xpb_out[91][38],u_xpb_out[92][38],u_xpb_out[93][38],u_xpb_out[94][38],u_xpb_out[95][38],u_xpb_out[96][38],u_xpb_out[97][38],u_xpb_out[98][38],u_xpb_out[99][38],u_xpb_out[100][38],u_xpb_out[101][38],u_xpb_out[102][38],u_xpb_out[103][38],u_xpb_out[104][38],u_xpb_out[105][38]};

assign col_out_39 = {u_xpb_out[0][39],u_xpb_out[1][39],u_xpb_out[2][39],u_xpb_out[3][39],u_xpb_out[4][39],u_xpb_out[5][39],u_xpb_out[6][39],u_xpb_out[7][39],u_xpb_out[8][39],u_xpb_out[9][39],u_xpb_out[10][39],u_xpb_out[11][39],u_xpb_out[12][39],u_xpb_out[13][39],u_xpb_out[14][39],u_xpb_out[15][39],u_xpb_out[16][39],u_xpb_out[17][39],u_xpb_out[18][39],u_xpb_out[19][39],u_xpb_out[20][39],u_xpb_out[21][39],u_xpb_out[22][39],u_xpb_out[23][39],u_xpb_out[24][39],u_xpb_out[25][39],u_xpb_out[26][39],u_xpb_out[27][39],u_xpb_out[28][39],u_xpb_out[29][39],u_xpb_out[30][39],u_xpb_out[31][39],u_xpb_out[32][39],u_xpb_out[33][39],u_xpb_out[34][39],u_xpb_out[35][39],u_xpb_out[36][39],u_xpb_out[37][39],u_xpb_out[38][39],u_xpb_out[39][39],u_xpb_out[40][39],u_xpb_out[41][39],u_xpb_out[42][39],u_xpb_out[43][39],u_xpb_out[44][39],u_xpb_out[45][39],u_xpb_out[46][39],u_xpb_out[47][39],u_xpb_out[48][39],u_xpb_out[49][39],u_xpb_out[50][39],u_xpb_out[51][39],u_xpb_out[52][39],u_xpb_out[53][39],u_xpb_out[54][39],u_xpb_out[55][39],u_xpb_out[56][39],u_xpb_out[57][39],u_xpb_out[58][39],u_xpb_out[59][39],u_xpb_out[60][39],u_xpb_out[61][39],u_xpb_out[62][39],u_xpb_out[63][39],u_xpb_out[64][39],u_xpb_out[65][39],u_xpb_out[66][39],u_xpb_out[67][39],u_xpb_out[68][39],u_xpb_out[69][39],u_xpb_out[70][39],u_xpb_out[71][39],u_xpb_out[72][39],u_xpb_out[73][39],u_xpb_out[74][39],u_xpb_out[75][39],u_xpb_out[76][39],u_xpb_out[77][39],u_xpb_out[78][39],u_xpb_out[79][39],u_xpb_out[80][39],u_xpb_out[81][39],u_xpb_out[82][39],u_xpb_out[83][39],u_xpb_out[84][39],u_xpb_out[85][39],u_xpb_out[86][39],u_xpb_out[87][39],u_xpb_out[88][39],u_xpb_out[89][39],u_xpb_out[90][39],u_xpb_out[91][39],u_xpb_out[92][39],u_xpb_out[93][39],u_xpb_out[94][39],u_xpb_out[95][39],u_xpb_out[96][39],u_xpb_out[97][39],u_xpb_out[98][39],u_xpb_out[99][39],u_xpb_out[100][39],u_xpb_out[101][39],u_xpb_out[102][39],u_xpb_out[103][39],u_xpb_out[104][39],u_xpb_out[105][39]};

assign col_out_40 = {u_xpb_out[0][40],u_xpb_out[1][40],u_xpb_out[2][40],u_xpb_out[3][40],u_xpb_out[4][40],u_xpb_out[5][40],u_xpb_out[6][40],u_xpb_out[7][40],u_xpb_out[8][40],u_xpb_out[9][40],u_xpb_out[10][40],u_xpb_out[11][40],u_xpb_out[12][40],u_xpb_out[13][40],u_xpb_out[14][40],u_xpb_out[15][40],u_xpb_out[16][40],u_xpb_out[17][40],u_xpb_out[18][40],u_xpb_out[19][40],u_xpb_out[20][40],u_xpb_out[21][40],u_xpb_out[22][40],u_xpb_out[23][40],u_xpb_out[24][40],u_xpb_out[25][40],u_xpb_out[26][40],u_xpb_out[27][40],u_xpb_out[28][40],u_xpb_out[29][40],u_xpb_out[30][40],u_xpb_out[31][40],u_xpb_out[32][40],u_xpb_out[33][40],u_xpb_out[34][40],u_xpb_out[35][40],u_xpb_out[36][40],u_xpb_out[37][40],u_xpb_out[38][40],u_xpb_out[39][40],u_xpb_out[40][40],u_xpb_out[41][40],u_xpb_out[42][40],u_xpb_out[43][40],u_xpb_out[44][40],u_xpb_out[45][40],u_xpb_out[46][40],u_xpb_out[47][40],u_xpb_out[48][40],u_xpb_out[49][40],u_xpb_out[50][40],u_xpb_out[51][40],u_xpb_out[52][40],u_xpb_out[53][40],u_xpb_out[54][40],u_xpb_out[55][40],u_xpb_out[56][40],u_xpb_out[57][40],u_xpb_out[58][40],u_xpb_out[59][40],u_xpb_out[60][40],u_xpb_out[61][40],u_xpb_out[62][40],u_xpb_out[63][40],u_xpb_out[64][40],u_xpb_out[65][40],u_xpb_out[66][40],u_xpb_out[67][40],u_xpb_out[68][40],u_xpb_out[69][40],u_xpb_out[70][40],u_xpb_out[71][40],u_xpb_out[72][40],u_xpb_out[73][40],u_xpb_out[74][40],u_xpb_out[75][40],u_xpb_out[76][40],u_xpb_out[77][40],u_xpb_out[78][40],u_xpb_out[79][40],u_xpb_out[80][40],u_xpb_out[81][40],u_xpb_out[82][40],u_xpb_out[83][40],u_xpb_out[84][40],u_xpb_out[85][40],u_xpb_out[86][40],u_xpb_out[87][40],u_xpb_out[88][40],u_xpb_out[89][40],u_xpb_out[90][40],u_xpb_out[91][40],u_xpb_out[92][40],u_xpb_out[93][40],u_xpb_out[94][40],u_xpb_out[95][40],u_xpb_out[96][40],u_xpb_out[97][40],u_xpb_out[98][40],u_xpb_out[99][40],u_xpb_out[100][40],u_xpb_out[101][40],u_xpb_out[102][40],u_xpb_out[103][40],u_xpb_out[104][40],u_xpb_out[105][40]};

assign col_out_41 = {u_xpb_out[0][41],u_xpb_out[1][41],u_xpb_out[2][41],u_xpb_out[3][41],u_xpb_out[4][41],u_xpb_out[5][41],u_xpb_out[6][41],u_xpb_out[7][41],u_xpb_out[8][41],u_xpb_out[9][41],u_xpb_out[10][41],u_xpb_out[11][41],u_xpb_out[12][41],u_xpb_out[13][41],u_xpb_out[14][41],u_xpb_out[15][41],u_xpb_out[16][41],u_xpb_out[17][41],u_xpb_out[18][41],u_xpb_out[19][41],u_xpb_out[20][41],u_xpb_out[21][41],u_xpb_out[22][41],u_xpb_out[23][41],u_xpb_out[24][41],u_xpb_out[25][41],u_xpb_out[26][41],u_xpb_out[27][41],u_xpb_out[28][41],u_xpb_out[29][41],u_xpb_out[30][41],u_xpb_out[31][41],u_xpb_out[32][41],u_xpb_out[33][41],u_xpb_out[34][41],u_xpb_out[35][41],u_xpb_out[36][41],u_xpb_out[37][41],u_xpb_out[38][41],u_xpb_out[39][41],u_xpb_out[40][41],u_xpb_out[41][41],u_xpb_out[42][41],u_xpb_out[43][41],u_xpb_out[44][41],u_xpb_out[45][41],u_xpb_out[46][41],u_xpb_out[47][41],u_xpb_out[48][41],u_xpb_out[49][41],u_xpb_out[50][41],u_xpb_out[51][41],u_xpb_out[52][41],u_xpb_out[53][41],u_xpb_out[54][41],u_xpb_out[55][41],u_xpb_out[56][41],u_xpb_out[57][41],u_xpb_out[58][41],u_xpb_out[59][41],u_xpb_out[60][41],u_xpb_out[61][41],u_xpb_out[62][41],u_xpb_out[63][41],u_xpb_out[64][41],u_xpb_out[65][41],u_xpb_out[66][41],u_xpb_out[67][41],u_xpb_out[68][41],u_xpb_out[69][41],u_xpb_out[70][41],u_xpb_out[71][41],u_xpb_out[72][41],u_xpb_out[73][41],u_xpb_out[74][41],u_xpb_out[75][41],u_xpb_out[76][41],u_xpb_out[77][41],u_xpb_out[78][41],u_xpb_out[79][41],u_xpb_out[80][41],u_xpb_out[81][41],u_xpb_out[82][41],u_xpb_out[83][41],u_xpb_out[84][41],u_xpb_out[85][41],u_xpb_out[86][41],u_xpb_out[87][41],u_xpb_out[88][41],u_xpb_out[89][41],u_xpb_out[90][41],u_xpb_out[91][41],u_xpb_out[92][41],u_xpb_out[93][41],u_xpb_out[94][41],u_xpb_out[95][41],u_xpb_out[96][41],u_xpb_out[97][41],u_xpb_out[98][41],u_xpb_out[99][41],u_xpb_out[100][41],u_xpb_out[101][41],u_xpb_out[102][41],u_xpb_out[103][41],u_xpb_out[104][41],u_xpb_out[105][41]};

assign col_out_42 = {u_xpb_out[0][42],u_xpb_out[1][42],u_xpb_out[2][42],u_xpb_out[3][42],u_xpb_out[4][42],u_xpb_out[5][42],u_xpb_out[6][42],u_xpb_out[7][42],u_xpb_out[8][42],u_xpb_out[9][42],u_xpb_out[10][42],u_xpb_out[11][42],u_xpb_out[12][42],u_xpb_out[13][42],u_xpb_out[14][42],u_xpb_out[15][42],u_xpb_out[16][42],u_xpb_out[17][42],u_xpb_out[18][42],u_xpb_out[19][42],u_xpb_out[20][42],u_xpb_out[21][42],u_xpb_out[22][42],u_xpb_out[23][42],u_xpb_out[24][42],u_xpb_out[25][42],u_xpb_out[26][42],u_xpb_out[27][42],u_xpb_out[28][42],u_xpb_out[29][42],u_xpb_out[30][42],u_xpb_out[31][42],u_xpb_out[32][42],u_xpb_out[33][42],u_xpb_out[34][42],u_xpb_out[35][42],u_xpb_out[36][42],u_xpb_out[37][42],u_xpb_out[38][42],u_xpb_out[39][42],u_xpb_out[40][42],u_xpb_out[41][42],u_xpb_out[42][42],u_xpb_out[43][42],u_xpb_out[44][42],u_xpb_out[45][42],u_xpb_out[46][42],u_xpb_out[47][42],u_xpb_out[48][42],u_xpb_out[49][42],u_xpb_out[50][42],u_xpb_out[51][42],u_xpb_out[52][42],u_xpb_out[53][42],u_xpb_out[54][42],u_xpb_out[55][42],u_xpb_out[56][42],u_xpb_out[57][42],u_xpb_out[58][42],u_xpb_out[59][42],u_xpb_out[60][42],u_xpb_out[61][42],u_xpb_out[62][42],u_xpb_out[63][42],u_xpb_out[64][42],u_xpb_out[65][42],u_xpb_out[66][42],u_xpb_out[67][42],u_xpb_out[68][42],u_xpb_out[69][42],u_xpb_out[70][42],u_xpb_out[71][42],u_xpb_out[72][42],u_xpb_out[73][42],u_xpb_out[74][42],u_xpb_out[75][42],u_xpb_out[76][42],u_xpb_out[77][42],u_xpb_out[78][42],u_xpb_out[79][42],u_xpb_out[80][42],u_xpb_out[81][42],u_xpb_out[82][42],u_xpb_out[83][42],u_xpb_out[84][42],u_xpb_out[85][42],u_xpb_out[86][42],u_xpb_out[87][42],u_xpb_out[88][42],u_xpb_out[89][42],u_xpb_out[90][42],u_xpb_out[91][42],u_xpb_out[92][42],u_xpb_out[93][42],u_xpb_out[94][42],u_xpb_out[95][42],u_xpb_out[96][42],u_xpb_out[97][42],u_xpb_out[98][42],u_xpb_out[99][42],u_xpb_out[100][42],u_xpb_out[101][42],u_xpb_out[102][42],u_xpb_out[103][42],u_xpb_out[104][42],u_xpb_out[105][42]};

assign col_out_43 = {u_xpb_out[0][43],u_xpb_out[1][43],u_xpb_out[2][43],u_xpb_out[3][43],u_xpb_out[4][43],u_xpb_out[5][43],u_xpb_out[6][43],u_xpb_out[7][43],u_xpb_out[8][43],u_xpb_out[9][43],u_xpb_out[10][43],u_xpb_out[11][43],u_xpb_out[12][43],u_xpb_out[13][43],u_xpb_out[14][43],u_xpb_out[15][43],u_xpb_out[16][43],u_xpb_out[17][43],u_xpb_out[18][43],u_xpb_out[19][43],u_xpb_out[20][43],u_xpb_out[21][43],u_xpb_out[22][43],u_xpb_out[23][43],u_xpb_out[24][43],u_xpb_out[25][43],u_xpb_out[26][43],u_xpb_out[27][43],u_xpb_out[28][43],u_xpb_out[29][43],u_xpb_out[30][43],u_xpb_out[31][43],u_xpb_out[32][43],u_xpb_out[33][43],u_xpb_out[34][43],u_xpb_out[35][43],u_xpb_out[36][43],u_xpb_out[37][43],u_xpb_out[38][43],u_xpb_out[39][43],u_xpb_out[40][43],u_xpb_out[41][43],u_xpb_out[42][43],u_xpb_out[43][43],u_xpb_out[44][43],u_xpb_out[45][43],u_xpb_out[46][43],u_xpb_out[47][43],u_xpb_out[48][43],u_xpb_out[49][43],u_xpb_out[50][43],u_xpb_out[51][43],u_xpb_out[52][43],u_xpb_out[53][43],u_xpb_out[54][43],u_xpb_out[55][43],u_xpb_out[56][43],u_xpb_out[57][43],u_xpb_out[58][43],u_xpb_out[59][43],u_xpb_out[60][43],u_xpb_out[61][43],u_xpb_out[62][43],u_xpb_out[63][43],u_xpb_out[64][43],u_xpb_out[65][43],u_xpb_out[66][43],u_xpb_out[67][43],u_xpb_out[68][43],u_xpb_out[69][43],u_xpb_out[70][43],u_xpb_out[71][43],u_xpb_out[72][43],u_xpb_out[73][43],u_xpb_out[74][43],u_xpb_out[75][43],u_xpb_out[76][43],u_xpb_out[77][43],u_xpb_out[78][43],u_xpb_out[79][43],u_xpb_out[80][43],u_xpb_out[81][43],u_xpb_out[82][43],u_xpb_out[83][43],u_xpb_out[84][43],u_xpb_out[85][43],u_xpb_out[86][43],u_xpb_out[87][43],u_xpb_out[88][43],u_xpb_out[89][43],u_xpb_out[90][43],u_xpb_out[91][43],u_xpb_out[92][43],u_xpb_out[93][43],u_xpb_out[94][43],u_xpb_out[95][43],u_xpb_out[96][43],u_xpb_out[97][43],u_xpb_out[98][43],u_xpb_out[99][43],u_xpb_out[100][43],u_xpb_out[101][43],u_xpb_out[102][43],u_xpb_out[103][43],u_xpb_out[104][43],u_xpb_out[105][43]};

assign col_out_44 = {u_xpb_out[0][44],u_xpb_out[1][44],u_xpb_out[2][44],u_xpb_out[3][44],u_xpb_out[4][44],u_xpb_out[5][44],u_xpb_out[6][44],u_xpb_out[7][44],u_xpb_out[8][44],u_xpb_out[9][44],u_xpb_out[10][44],u_xpb_out[11][44],u_xpb_out[12][44],u_xpb_out[13][44],u_xpb_out[14][44],u_xpb_out[15][44],u_xpb_out[16][44],u_xpb_out[17][44],u_xpb_out[18][44],u_xpb_out[19][44],u_xpb_out[20][44],u_xpb_out[21][44],u_xpb_out[22][44],u_xpb_out[23][44],u_xpb_out[24][44],u_xpb_out[25][44],u_xpb_out[26][44],u_xpb_out[27][44],u_xpb_out[28][44],u_xpb_out[29][44],u_xpb_out[30][44],u_xpb_out[31][44],u_xpb_out[32][44],u_xpb_out[33][44],u_xpb_out[34][44],u_xpb_out[35][44],u_xpb_out[36][44],u_xpb_out[37][44],u_xpb_out[38][44],u_xpb_out[39][44],u_xpb_out[40][44],u_xpb_out[41][44],u_xpb_out[42][44],u_xpb_out[43][44],u_xpb_out[44][44],u_xpb_out[45][44],u_xpb_out[46][44],u_xpb_out[47][44],u_xpb_out[48][44],u_xpb_out[49][44],u_xpb_out[50][44],u_xpb_out[51][44],u_xpb_out[52][44],u_xpb_out[53][44],u_xpb_out[54][44],u_xpb_out[55][44],u_xpb_out[56][44],u_xpb_out[57][44],u_xpb_out[58][44],u_xpb_out[59][44],u_xpb_out[60][44],u_xpb_out[61][44],u_xpb_out[62][44],u_xpb_out[63][44],u_xpb_out[64][44],u_xpb_out[65][44],u_xpb_out[66][44],u_xpb_out[67][44],u_xpb_out[68][44],u_xpb_out[69][44],u_xpb_out[70][44],u_xpb_out[71][44],u_xpb_out[72][44],u_xpb_out[73][44],u_xpb_out[74][44],u_xpb_out[75][44],u_xpb_out[76][44],u_xpb_out[77][44],u_xpb_out[78][44],u_xpb_out[79][44],u_xpb_out[80][44],u_xpb_out[81][44],u_xpb_out[82][44],u_xpb_out[83][44],u_xpb_out[84][44],u_xpb_out[85][44],u_xpb_out[86][44],u_xpb_out[87][44],u_xpb_out[88][44],u_xpb_out[89][44],u_xpb_out[90][44],u_xpb_out[91][44],u_xpb_out[92][44],u_xpb_out[93][44],u_xpb_out[94][44],u_xpb_out[95][44],u_xpb_out[96][44],u_xpb_out[97][44],u_xpb_out[98][44],u_xpb_out[99][44],u_xpb_out[100][44],u_xpb_out[101][44],u_xpb_out[102][44],u_xpb_out[103][44],u_xpb_out[104][44],u_xpb_out[105][44]};

assign col_out_45 = {u_xpb_out[0][45],u_xpb_out[1][45],u_xpb_out[2][45],u_xpb_out[3][45],u_xpb_out[4][45],u_xpb_out[5][45],u_xpb_out[6][45],u_xpb_out[7][45],u_xpb_out[8][45],u_xpb_out[9][45],u_xpb_out[10][45],u_xpb_out[11][45],u_xpb_out[12][45],u_xpb_out[13][45],u_xpb_out[14][45],u_xpb_out[15][45],u_xpb_out[16][45],u_xpb_out[17][45],u_xpb_out[18][45],u_xpb_out[19][45],u_xpb_out[20][45],u_xpb_out[21][45],u_xpb_out[22][45],u_xpb_out[23][45],u_xpb_out[24][45],u_xpb_out[25][45],u_xpb_out[26][45],u_xpb_out[27][45],u_xpb_out[28][45],u_xpb_out[29][45],u_xpb_out[30][45],u_xpb_out[31][45],u_xpb_out[32][45],u_xpb_out[33][45],u_xpb_out[34][45],u_xpb_out[35][45],u_xpb_out[36][45],u_xpb_out[37][45],u_xpb_out[38][45],u_xpb_out[39][45],u_xpb_out[40][45],u_xpb_out[41][45],u_xpb_out[42][45],u_xpb_out[43][45],u_xpb_out[44][45],u_xpb_out[45][45],u_xpb_out[46][45],u_xpb_out[47][45],u_xpb_out[48][45],u_xpb_out[49][45],u_xpb_out[50][45],u_xpb_out[51][45],u_xpb_out[52][45],u_xpb_out[53][45],u_xpb_out[54][45],u_xpb_out[55][45],u_xpb_out[56][45],u_xpb_out[57][45],u_xpb_out[58][45],u_xpb_out[59][45],u_xpb_out[60][45],u_xpb_out[61][45],u_xpb_out[62][45],u_xpb_out[63][45],u_xpb_out[64][45],u_xpb_out[65][45],u_xpb_out[66][45],u_xpb_out[67][45],u_xpb_out[68][45],u_xpb_out[69][45],u_xpb_out[70][45],u_xpb_out[71][45],u_xpb_out[72][45],u_xpb_out[73][45],u_xpb_out[74][45],u_xpb_out[75][45],u_xpb_out[76][45],u_xpb_out[77][45],u_xpb_out[78][45],u_xpb_out[79][45],u_xpb_out[80][45],u_xpb_out[81][45],u_xpb_out[82][45],u_xpb_out[83][45],u_xpb_out[84][45],u_xpb_out[85][45],u_xpb_out[86][45],u_xpb_out[87][45],u_xpb_out[88][45],u_xpb_out[89][45],u_xpb_out[90][45],u_xpb_out[91][45],u_xpb_out[92][45],u_xpb_out[93][45],u_xpb_out[94][45],u_xpb_out[95][45],u_xpb_out[96][45],u_xpb_out[97][45],u_xpb_out[98][45],u_xpb_out[99][45],u_xpb_out[100][45],u_xpb_out[101][45],u_xpb_out[102][45],u_xpb_out[103][45],u_xpb_out[104][45],u_xpb_out[105][45]};

assign col_out_46 = {u_xpb_out[0][46],u_xpb_out[1][46],u_xpb_out[2][46],u_xpb_out[3][46],u_xpb_out[4][46],u_xpb_out[5][46],u_xpb_out[6][46],u_xpb_out[7][46],u_xpb_out[8][46],u_xpb_out[9][46],u_xpb_out[10][46],u_xpb_out[11][46],u_xpb_out[12][46],u_xpb_out[13][46],u_xpb_out[14][46],u_xpb_out[15][46],u_xpb_out[16][46],u_xpb_out[17][46],u_xpb_out[18][46],u_xpb_out[19][46],u_xpb_out[20][46],u_xpb_out[21][46],u_xpb_out[22][46],u_xpb_out[23][46],u_xpb_out[24][46],u_xpb_out[25][46],u_xpb_out[26][46],u_xpb_out[27][46],u_xpb_out[28][46],u_xpb_out[29][46],u_xpb_out[30][46],u_xpb_out[31][46],u_xpb_out[32][46],u_xpb_out[33][46],u_xpb_out[34][46],u_xpb_out[35][46],u_xpb_out[36][46],u_xpb_out[37][46],u_xpb_out[38][46],u_xpb_out[39][46],u_xpb_out[40][46],u_xpb_out[41][46],u_xpb_out[42][46],u_xpb_out[43][46],u_xpb_out[44][46],u_xpb_out[45][46],u_xpb_out[46][46],u_xpb_out[47][46],u_xpb_out[48][46],u_xpb_out[49][46],u_xpb_out[50][46],u_xpb_out[51][46],u_xpb_out[52][46],u_xpb_out[53][46],u_xpb_out[54][46],u_xpb_out[55][46],u_xpb_out[56][46],u_xpb_out[57][46],u_xpb_out[58][46],u_xpb_out[59][46],u_xpb_out[60][46],u_xpb_out[61][46],u_xpb_out[62][46],u_xpb_out[63][46],u_xpb_out[64][46],u_xpb_out[65][46],u_xpb_out[66][46],u_xpb_out[67][46],u_xpb_out[68][46],u_xpb_out[69][46],u_xpb_out[70][46],u_xpb_out[71][46],u_xpb_out[72][46],u_xpb_out[73][46],u_xpb_out[74][46],u_xpb_out[75][46],u_xpb_out[76][46],u_xpb_out[77][46],u_xpb_out[78][46],u_xpb_out[79][46],u_xpb_out[80][46],u_xpb_out[81][46],u_xpb_out[82][46],u_xpb_out[83][46],u_xpb_out[84][46],u_xpb_out[85][46],u_xpb_out[86][46],u_xpb_out[87][46],u_xpb_out[88][46],u_xpb_out[89][46],u_xpb_out[90][46],u_xpb_out[91][46],u_xpb_out[92][46],u_xpb_out[93][46],u_xpb_out[94][46],u_xpb_out[95][46],u_xpb_out[96][46],u_xpb_out[97][46],u_xpb_out[98][46],u_xpb_out[99][46],u_xpb_out[100][46],u_xpb_out[101][46],u_xpb_out[102][46],u_xpb_out[103][46],u_xpb_out[104][46],u_xpb_out[105][46]};

assign col_out_47 = {u_xpb_out[0][47],u_xpb_out[1][47],u_xpb_out[2][47],u_xpb_out[3][47],u_xpb_out[4][47],u_xpb_out[5][47],u_xpb_out[6][47],u_xpb_out[7][47],u_xpb_out[8][47],u_xpb_out[9][47],u_xpb_out[10][47],u_xpb_out[11][47],u_xpb_out[12][47],u_xpb_out[13][47],u_xpb_out[14][47],u_xpb_out[15][47],u_xpb_out[16][47],u_xpb_out[17][47],u_xpb_out[18][47],u_xpb_out[19][47],u_xpb_out[20][47],u_xpb_out[21][47],u_xpb_out[22][47],u_xpb_out[23][47],u_xpb_out[24][47],u_xpb_out[25][47],u_xpb_out[26][47],u_xpb_out[27][47],u_xpb_out[28][47],u_xpb_out[29][47],u_xpb_out[30][47],u_xpb_out[31][47],u_xpb_out[32][47],u_xpb_out[33][47],u_xpb_out[34][47],u_xpb_out[35][47],u_xpb_out[36][47],u_xpb_out[37][47],u_xpb_out[38][47],u_xpb_out[39][47],u_xpb_out[40][47],u_xpb_out[41][47],u_xpb_out[42][47],u_xpb_out[43][47],u_xpb_out[44][47],u_xpb_out[45][47],u_xpb_out[46][47],u_xpb_out[47][47],u_xpb_out[48][47],u_xpb_out[49][47],u_xpb_out[50][47],u_xpb_out[51][47],u_xpb_out[52][47],u_xpb_out[53][47],u_xpb_out[54][47],u_xpb_out[55][47],u_xpb_out[56][47],u_xpb_out[57][47],u_xpb_out[58][47],u_xpb_out[59][47],u_xpb_out[60][47],u_xpb_out[61][47],u_xpb_out[62][47],u_xpb_out[63][47],u_xpb_out[64][47],u_xpb_out[65][47],u_xpb_out[66][47],u_xpb_out[67][47],u_xpb_out[68][47],u_xpb_out[69][47],u_xpb_out[70][47],u_xpb_out[71][47],u_xpb_out[72][47],u_xpb_out[73][47],u_xpb_out[74][47],u_xpb_out[75][47],u_xpb_out[76][47],u_xpb_out[77][47],u_xpb_out[78][47],u_xpb_out[79][47],u_xpb_out[80][47],u_xpb_out[81][47],u_xpb_out[82][47],u_xpb_out[83][47],u_xpb_out[84][47],u_xpb_out[85][47],u_xpb_out[86][47],u_xpb_out[87][47],u_xpb_out[88][47],u_xpb_out[89][47],u_xpb_out[90][47],u_xpb_out[91][47],u_xpb_out[92][47],u_xpb_out[93][47],u_xpb_out[94][47],u_xpb_out[95][47],u_xpb_out[96][47],u_xpb_out[97][47],u_xpb_out[98][47],u_xpb_out[99][47],u_xpb_out[100][47],u_xpb_out[101][47],u_xpb_out[102][47],u_xpb_out[103][47],u_xpb_out[104][47],u_xpb_out[105][47]};

assign col_out_48 = {u_xpb_out[0][48],u_xpb_out[1][48],u_xpb_out[2][48],u_xpb_out[3][48],u_xpb_out[4][48],u_xpb_out[5][48],u_xpb_out[6][48],u_xpb_out[7][48],u_xpb_out[8][48],u_xpb_out[9][48],u_xpb_out[10][48],u_xpb_out[11][48],u_xpb_out[12][48],u_xpb_out[13][48],u_xpb_out[14][48],u_xpb_out[15][48],u_xpb_out[16][48],u_xpb_out[17][48],u_xpb_out[18][48],u_xpb_out[19][48],u_xpb_out[20][48],u_xpb_out[21][48],u_xpb_out[22][48],u_xpb_out[23][48],u_xpb_out[24][48],u_xpb_out[25][48],u_xpb_out[26][48],u_xpb_out[27][48],u_xpb_out[28][48],u_xpb_out[29][48],u_xpb_out[30][48],u_xpb_out[31][48],u_xpb_out[32][48],u_xpb_out[33][48],u_xpb_out[34][48],u_xpb_out[35][48],u_xpb_out[36][48],u_xpb_out[37][48],u_xpb_out[38][48],u_xpb_out[39][48],u_xpb_out[40][48],u_xpb_out[41][48],u_xpb_out[42][48],u_xpb_out[43][48],u_xpb_out[44][48],u_xpb_out[45][48],u_xpb_out[46][48],u_xpb_out[47][48],u_xpb_out[48][48],u_xpb_out[49][48],u_xpb_out[50][48],u_xpb_out[51][48],u_xpb_out[52][48],u_xpb_out[53][48],u_xpb_out[54][48],u_xpb_out[55][48],u_xpb_out[56][48],u_xpb_out[57][48],u_xpb_out[58][48],u_xpb_out[59][48],u_xpb_out[60][48],u_xpb_out[61][48],u_xpb_out[62][48],u_xpb_out[63][48],u_xpb_out[64][48],u_xpb_out[65][48],u_xpb_out[66][48],u_xpb_out[67][48],u_xpb_out[68][48],u_xpb_out[69][48],u_xpb_out[70][48],u_xpb_out[71][48],u_xpb_out[72][48],u_xpb_out[73][48],u_xpb_out[74][48],u_xpb_out[75][48],u_xpb_out[76][48],u_xpb_out[77][48],u_xpb_out[78][48],u_xpb_out[79][48],u_xpb_out[80][48],u_xpb_out[81][48],u_xpb_out[82][48],u_xpb_out[83][48],u_xpb_out[84][48],u_xpb_out[85][48],u_xpb_out[86][48],u_xpb_out[87][48],u_xpb_out[88][48],u_xpb_out[89][48],u_xpb_out[90][48],u_xpb_out[91][48],u_xpb_out[92][48],u_xpb_out[93][48],u_xpb_out[94][48],u_xpb_out[95][48],u_xpb_out[96][48],u_xpb_out[97][48],u_xpb_out[98][48],u_xpb_out[99][48],u_xpb_out[100][48],u_xpb_out[101][48],u_xpb_out[102][48],u_xpb_out[103][48],u_xpb_out[104][48],u_xpb_out[105][48]};

assign col_out_49 = {u_xpb_out[0][49],u_xpb_out[1][49],u_xpb_out[2][49],u_xpb_out[3][49],u_xpb_out[4][49],u_xpb_out[5][49],u_xpb_out[6][49],u_xpb_out[7][49],u_xpb_out[8][49],u_xpb_out[9][49],u_xpb_out[10][49],u_xpb_out[11][49],u_xpb_out[12][49],u_xpb_out[13][49],u_xpb_out[14][49],u_xpb_out[15][49],u_xpb_out[16][49],u_xpb_out[17][49],u_xpb_out[18][49],u_xpb_out[19][49],u_xpb_out[20][49],u_xpb_out[21][49],u_xpb_out[22][49],u_xpb_out[23][49],u_xpb_out[24][49],u_xpb_out[25][49],u_xpb_out[26][49],u_xpb_out[27][49],u_xpb_out[28][49],u_xpb_out[29][49],u_xpb_out[30][49],u_xpb_out[31][49],u_xpb_out[32][49],u_xpb_out[33][49],u_xpb_out[34][49],u_xpb_out[35][49],u_xpb_out[36][49],u_xpb_out[37][49],u_xpb_out[38][49],u_xpb_out[39][49],u_xpb_out[40][49],u_xpb_out[41][49],u_xpb_out[42][49],u_xpb_out[43][49],u_xpb_out[44][49],u_xpb_out[45][49],u_xpb_out[46][49],u_xpb_out[47][49],u_xpb_out[48][49],u_xpb_out[49][49],u_xpb_out[50][49],u_xpb_out[51][49],u_xpb_out[52][49],u_xpb_out[53][49],u_xpb_out[54][49],u_xpb_out[55][49],u_xpb_out[56][49],u_xpb_out[57][49],u_xpb_out[58][49],u_xpb_out[59][49],u_xpb_out[60][49],u_xpb_out[61][49],u_xpb_out[62][49],u_xpb_out[63][49],u_xpb_out[64][49],u_xpb_out[65][49],u_xpb_out[66][49],u_xpb_out[67][49],u_xpb_out[68][49],u_xpb_out[69][49],u_xpb_out[70][49],u_xpb_out[71][49],u_xpb_out[72][49],u_xpb_out[73][49],u_xpb_out[74][49],u_xpb_out[75][49],u_xpb_out[76][49],u_xpb_out[77][49],u_xpb_out[78][49],u_xpb_out[79][49],u_xpb_out[80][49],u_xpb_out[81][49],u_xpb_out[82][49],u_xpb_out[83][49],u_xpb_out[84][49],u_xpb_out[85][49],u_xpb_out[86][49],u_xpb_out[87][49],u_xpb_out[88][49],u_xpb_out[89][49],u_xpb_out[90][49],u_xpb_out[91][49],u_xpb_out[92][49],u_xpb_out[93][49],u_xpb_out[94][49],u_xpb_out[95][49],u_xpb_out[96][49],u_xpb_out[97][49],u_xpb_out[98][49],u_xpb_out[99][49],u_xpb_out[100][49],u_xpb_out[101][49],u_xpb_out[102][49],u_xpb_out[103][49],u_xpb_out[104][49],u_xpb_out[105][49]};

assign col_out_50 = {u_xpb_out[0][50],u_xpb_out[1][50],u_xpb_out[2][50],u_xpb_out[3][50],u_xpb_out[4][50],u_xpb_out[5][50],u_xpb_out[6][50],u_xpb_out[7][50],u_xpb_out[8][50],u_xpb_out[9][50],u_xpb_out[10][50],u_xpb_out[11][50],u_xpb_out[12][50],u_xpb_out[13][50],u_xpb_out[14][50],u_xpb_out[15][50],u_xpb_out[16][50],u_xpb_out[17][50],u_xpb_out[18][50],u_xpb_out[19][50],u_xpb_out[20][50],u_xpb_out[21][50],u_xpb_out[22][50],u_xpb_out[23][50],u_xpb_out[24][50],u_xpb_out[25][50],u_xpb_out[26][50],u_xpb_out[27][50],u_xpb_out[28][50],u_xpb_out[29][50],u_xpb_out[30][50],u_xpb_out[31][50],u_xpb_out[32][50],u_xpb_out[33][50],u_xpb_out[34][50],u_xpb_out[35][50],u_xpb_out[36][50],u_xpb_out[37][50],u_xpb_out[38][50],u_xpb_out[39][50],u_xpb_out[40][50],u_xpb_out[41][50],u_xpb_out[42][50],u_xpb_out[43][50],u_xpb_out[44][50],u_xpb_out[45][50],u_xpb_out[46][50],u_xpb_out[47][50],u_xpb_out[48][50],u_xpb_out[49][50],u_xpb_out[50][50],u_xpb_out[51][50],u_xpb_out[52][50],u_xpb_out[53][50],u_xpb_out[54][50],u_xpb_out[55][50],u_xpb_out[56][50],u_xpb_out[57][50],u_xpb_out[58][50],u_xpb_out[59][50],u_xpb_out[60][50],u_xpb_out[61][50],u_xpb_out[62][50],u_xpb_out[63][50],u_xpb_out[64][50],u_xpb_out[65][50],u_xpb_out[66][50],u_xpb_out[67][50],u_xpb_out[68][50],u_xpb_out[69][50],u_xpb_out[70][50],u_xpb_out[71][50],u_xpb_out[72][50],u_xpb_out[73][50],u_xpb_out[74][50],u_xpb_out[75][50],u_xpb_out[76][50],u_xpb_out[77][50],u_xpb_out[78][50],u_xpb_out[79][50],u_xpb_out[80][50],u_xpb_out[81][50],u_xpb_out[82][50],u_xpb_out[83][50],u_xpb_out[84][50],u_xpb_out[85][50],u_xpb_out[86][50],u_xpb_out[87][50],u_xpb_out[88][50],u_xpb_out[89][50],u_xpb_out[90][50],u_xpb_out[91][50],u_xpb_out[92][50],u_xpb_out[93][50],u_xpb_out[94][50],u_xpb_out[95][50],u_xpb_out[96][50],u_xpb_out[97][50],u_xpb_out[98][50],u_xpb_out[99][50],u_xpb_out[100][50],u_xpb_out[101][50],u_xpb_out[102][50],u_xpb_out[103][50],u_xpb_out[104][50],u_xpb_out[105][50]};

assign col_out_51 = {u_xpb_out[0][51],u_xpb_out[1][51],u_xpb_out[2][51],u_xpb_out[3][51],u_xpb_out[4][51],u_xpb_out[5][51],u_xpb_out[6][51],u_xpb_out[7][51],u_xpb_out[8][51],u_xpb_out[9][51],u_xpb_out[10][51],u_xpb_out[11][51],u_xpb_out[12][51],u_xpb_out[13][51],u_xpb_out[14][51],u_xpb_out[15][51],u_xpb_out[16][51],u_xpb_out[17][51],u_xpb_out[18][51],u_xpb_out[19][51],u_xpb_out[20][51],u_xpb_out[21][51],u_xpb_out[22][51],u_xpb_out[23][51],u_xpb_out[24][51],u_xpb_out[25][51],u_xpb_out[26][51],u_xpb_out[27][51],u_xpb_out[28][51],u_xpb_out[29][51],u_xpb_out[30][51],u_xpb_out[31][51],u_xpb_out[32][51],u_xpb_out[33][51],u_xpb_out[34][51],u_xpb_out[35][51],u_xpb_out[36][51],u_xpb_out[37][51],u_xpb_out[38][51],u_xpb_out[39][51],u_xpb_out[40][51],u_xpb_out[41][51],u_xpb_out[42][51],u_xpb_out[43][51],u_xpb_out[44][51],u_xpb_out[45][51],u_xpb_out[46][51],u_xpb_out[47][51],u_xpb_out[48][51],u_xpb_out[49][51],u_xpb_out[50][51],u_xpb_out[51][51],u_xpb_out[52][51],u_xpb_out[53][51],u_xpb_out[54][51],u_xpb_out[55][51],u_xpb_out[56][51],u_xpb_out[57][51],u_xpb_out[58][51],u_xpb_out[59][51],u_xpb_out[60][51],u_xpb_out[61][51],u_xpb_out[62][51],u_xpb_out[63][51],u_xpb_out[64][51],u_xpb_out[65][51],u_xpb_out[66][51],u_xpb_out[67][51],u_xpb_out[68][51],u_xpb_out[69][51],u_xpb_out[70][51],u_xpb_out[71][51],u_xpb_out[72][51],u_xpb_out[73][51],u_xpb_out[74][51],u_xpb_out[75][51],u_xpb_out[76][51],u_xpb_out[77][51],u_xpb_out[78][51],u_xpb_out[79][51],u_xpb_out[80][51],u_xpb_out[81][51],u_xpb_out[82][51],u_xpb_out[83][51],u_xpb_out[84][51],u_xpb_out[85][51],u_xpb_out[86][51],u_xpb_out[87][51],u_xpb_out[88][51],u_xpb_out[89][51],u_xpb_out[90][51],u_xpb_out[91][51],u_xpb_out[92][51],u_xpb_out[93][51],u_xpb_out[94][51],u_xpb_out[95][51],u_xpb_out[96][51],u_xpb_out[97][51],u_xpb_out[98][51],u_xpb_out[99][51],u_xpb_out[100][51],u_xpb_out[101][51],u_xpb_out[102][51],u_xpb_out[103][51],u_xpb_out[104][51],u_xpb_out[105][51]};

assign col_out_52 = {u_xpb_out[0][52],u_xpb_out[1][52],u_xpb_out[2][52],u_xpb_out[3][52],u_xpb_out[4][52],u_xpb_out[5][52],u_xpb_out[6][52],u_xpb_out[7][52],u_xpb_out[8][52],u_xpb_out[9][52],u_xpb_out[10][52],u_xpb_out[11][52],u_xpb_out[12][52],u_xpb_out[13][52],u_xpb_out[14][52],u_xpb_out[15][52],u_xpb_out[16][52],u_xpb_out[17][52],u_xpb_out[18][52],u_xpb_out[19][52],u_xpb_out[20][52],u_xpb_out[21][52],u_xpb_out[22][52],u_xpb_out[23][52],u_xpb_out[24][52],u_xpb_out[25][52],u_xpb_out[26][52],u_xpb_out[27][52],u_xpb_out[28][52],u_xpb_out[29][52],u_xpb_out[30][52],u_xpb_out[31][52],u_xpb_out[32][52],u_xpb_out[33][52],u_xpb_out[34][52],u_xpb_out[35][52],u_xpb_out[36][52],u_xpb_out[37][52],u_xpb_out[38][52],u_xpb_out[39][52],u_xpb_out[40][52],u_xpb_out[41][52],u_xpb_out[42][52],u_xpb_out[43][52],u_xpb_out[44][52],u_xpb_out[45][52],u_xpb_out[46][52],u_xpb_out[47][52],u_xpb_out[48][52],u_xpb_out[49][52],u_xpb_out[50][52],u_xpb_out[51][52],u_xpb_out[52][52],u_xpb_out[53][52],u_xpb_out[54][52],u_xpb_out[55][52],u_xpb_out[56][52],u_xpb_out[57][52],u_xpb_out[58][52],u_xpb_out[59][52],u_xpb_out[60][52],u_xpb_out[61][52],u_xpb_out[62][52],u_xpb_out[63][52],u_xpb_out[64][52],u_xpb_out[65][52],u_xpb_out[66][52],u_xpb_out[67][52],u_xpb_out[68][52],u_xpb_out[69][52],u_xpb_out[70][52],u_xpb_out[71][52],u_xpb_out[72][52],u_xpb_out[73][52],u_xpb_out[74][52],u_xpb_out[75][52],u_xpb_out[76][52],u_xpb_out[77][52],u_xpb_out[78][52],u_xpb_out[79][52],u_xpb_out[80][52],u_xpb_out[81][52],u_xpb_out[82][52],u_xpb_out[83][52],u_xpb_out[84][52],u_xpb_out[85][52],u_xpb_out[86][52],u_xpb_out[87][52],u_xpb_out[88][52],u_xpb_out[89][52],u_xpb_out[90][52],u_xpb_out[91][52],u_xpb_out[92][52],u_xpb_out[93][52],u_xpb_out[94][52],u_xpb_out[95][52],u_xpb_out[96][52],u_xpb_out[97][52],u_xpb_out[98][52],u_xpb_out[99][52],u_xpb_out[100][52],u_xpb_out[101][52],u_xpb_out[102][52],u_xpb_out[103][52],u_xpb_out[104][52],u_xpb_out[105][52]};

assign col_out_53 = {u_xpb_out[0][53],u_xpb_out[1][53],u_xpb_out[2][53],u_xpb_out[3][53],u_xpb_out[4][53],u_xpb_out[5][53],u_xpb_out[6][53],u_xpb_out[7][53],u_xpb_out[8][53],u_xpb_out[9][53],u_xpb_out[10][53],u_xpb_out[11][53],u_xpb_out[12][53],u_xpb_out[13][53],u_xpb_out[14][53],u_xpb_out[15][53],u_xpb_out[16][53],u_xpb_out[17][53],u_xpb_out[18][53],u_xpb_out[19][53],u_xpb_out[20][53],u_xpb_out[21][53],u_xpb_out[22][53],u_xpb_out[23][53],u_xpb_out[24][53],u_xpb_out[25][53],u_xpb_out[26][53],u_xpb_out[27][53],u_xpb_out[28][53],u_xpb_out[29][53],u_xpb_out[30][53],u_xpb_out[31][53],u_xpb_out[32][53],u_xpb_out[33][53],u_xpb_out[34][53],u_xpb_out[35][53],u_xpb_out[36][53],u_xpb_out[37][53],u_xpb_out[38][53],u_xpb_out[39][53],u_xpb_out[40][53],u_xpb_out[41][53],u_xpb_out[42][53],u_xpb_out[43][53],u_xpb_out[44][53],u_xpb_out[45][53],u_xpb_out[46][53],u_xpb_out[47][53],u_xpb_out[48][53],u_xpb_out[49][53],u_xpb_out[50][53],u_xpb_out[51][53],u_xpb_out[52][53],u_xpb_out[53][53],u_xpb_out[54][53],u_xpb_out[55][53],u_xpb_out[56][53],u_xpb_out[57][53],u_xpb_out[58][53],u_xpb_out[59][53],u_xpb_out[60][53],u_xpb_out[61][53],u_xpb_out[62][53],u_xpb_out[63][53],u_xpb_out[64][53],u_xpb_out[65][53],u_xpb_out[66][53],u_xpb_out[67][53],u_xpb_out[68][53],u_xpb_out[69][53],u_xpb_out[70][53],u_xpb_out[71][53],u_xpb_out[72][53],u_xpb_out[73][53],u_xpb_out[74][53],u_xpb_out[75][53],u_xpb_out[76][53],u_xpb_out[77][53],u_xpb_out[78][53],u_xpb_out[79][53],u_xpb_out[80][53],u_xpb_out[81][53],u_xpb_out[82][53],u_xpb_out[83][53],u_xpb_out[84][53],u_xpb_out[85][53],u_xpb_out[86][53],u_xpb_out[87][53],u_xpb_out[88][53],u_xpb_out[89][53],u_xpb_out[90][53],u_xpb_out[91][53],u_xpb_out[92][53],u_xpb_out[93][53],u_xpb_out[94][53],u_xpb_out[95][53],u_xpb_out[96][53],u_xpb_out[97][53],u_xpb_out[98][53],u_xpb_out[99][53],u_xpb_out[100][53],u_xpb_out[101][53],u_xpb_out[102][53],u_xpb_out[103][53],u_xpb_out[104][53],u_xpb_out[105][53]};

assign col_out_54 = {u_xpb_out[0][54],u_xpb_out[1][54],u_xpb_out[2][54],u_xpb_out[3][54],u_xpb_out[4][54],u_xpb_out[5][54],u_xpb_out[6][54],u_xpb_out[7][54],u_xpb_out[8][54],u_xpb_out[9][54],u_xpb_out[10][54],u_xpb_out[11][54],u_xpb_out[12][54],u_xpb_out[13][54],u_xpb_out[14][54],u_xpb_out[15][54],u_xpb_out[16][54],u_xpb_out[17][54],u_xpb_out[18][54],u_xpb_out[19][54],u_xpb_out[20][54],u_xpb_out[21][54],u_xpb_out[22][54],u_xpb_out[23][54],u_xpb_out[24][54],u_xpb_out[25][54],u_xpb_out[26][54],u_xpb_out[27][54],u_xpb_out[28][54],u_xpb_out[29][54],u_xpb_out[30][54],u_xpb_out[31][54],u_xpb_out[32][54],u_xpb_out[33][54],u_xpb_out[34][54],u_xpb_out[35][54],u_xpb_out[36][54],u_xpb_out[37][54],u_xpb_out[38][54],u_xpb_out[39][54],u_xpb_out[40][54],u_xpb_out[41][54],u_xpb_out[42][54],u_xpb_out[43][54],u_xpb_out[44][54],u_xpb_out[45][54],u_xpb_out[46][54],u_xpb_out[47][54],u_xpb_out[48][54],u_xpb_out[49][54],u_xpb_out[50][54],u_xpb_out[51][54],u_xpb_out[52][54],u_xpb_out[53][54],u_xpb_out[54][54],u_xpb_out[55][54],u_xpb_out[56][54],u_xpb_out[57][54],u_xpb_out[58][54],u_xpb_out[59][54],u_xpb_out[60][54],u_xpb_out[61][54],u_xpb_out[62][54],u_xpb_out[63][54],u_xpb_out[64][54],u_xpb_out[65][54],u_xpb_out[66][54],u_xpb_out[67][54],u_xpb_out[68][54],u_xpb_out[69][54],u_xpb_out[70][54],u_xpb_out[71][54],u_xpb_out[72][54],u_xpb_out[73][54],u_xpb_out[74][54],u_xpb_out[75][54],u_xpb_out[76][54],u_xpb_out[77][54],u_xpb_out[78][54],u_xpb_out[79][54],u_xpb_out[80][54],u_xpb_out[81][54],u_xpb_out[82][54],u_xpb_out[83][54],u_xpb_out[84][54],u_xpb_out[85][54],u_xpb_out[86][54],u_xpb_out[87][54],u_xpb_out[88][54],u_xpb_out[89][54],u_xpb_out[90][54],u_xpb_out[91][54],u_xpb_out[92][54],u_xpb_out[93][54],u_xpb_out[94][54],u_xpb_out[95][54],u_xpb_out[96][54],u_xpb_out[97][54],u_xpb_out[98][54],u_xpb_out[99][54],u_xpb_out[100][54],u_xpb_out[101][54],u_xpb_out[102][54],u_xpb_out[103][54],u_xpb_out[104][54],u_xpb_out[105][54]};

assign col_out_55 = {u_xpb_out[0][55],u_xpb_out[1][55],u_xpb_out[2][55],u_xpb_out[3][55],u_xpb_out[4][55],u_xpb_out[5][55],u_xpb_out[6][55],u_xpb_out[7][55],u_xpb_out[8][55],u_xpb_out[9][55],u_xpb_out[10][55],u_xpb_out[11][55],u_xpb_out[12][55],u_xpb_out[13][55],u_xpb_out[14][55],u_xpb_out[15][55],u_xpb_out[16][55],u_xpb_out[17][55],u_xpb_out[18][55],u_xpb_out[19][55],u_xpb_out[20][55],u_xpb_out[21][55],u_xpb_out[22][55],u_xpb_out[23][55],u_xpb_out[24][55],u_xpb_out[25][55],u_xpb_out[26][55],u_xpb_out[27][55],u_xpb_out[28][55],u_xpb_out[29][55],u_xpb_out[30][55],u_xpb_out[31][55],u_xpb_out[32][55],u_xpb_out[33][55],u_xpb_out[34][55],u_xpb_out[35][55],u_xpb_out[36][55],u_xpb_out[37][55],u_xpb_out[38][55],u_xpb_out[39][55],u_xpb_out[40][55],u_xpb_out[41][55],u_xpb_out[42][55],u_xpb_out[43][55],u_xpb_out[44][55],u_xpb_out[45][55],u_xpb_out[46][55],u_xpb_out[47][55],u_xpb_out[48][55],u_xpb_out[49][55],u_xpb_out[50][55],u_xpb_out[51][55],u_xpb_out[52][55],u_xpb_out[53][55],u_xpb_out[54][55],u_xpb_out[55][55],u_xpb_out[56][55],u_xpb_out[57][55],u_xpb_out[58][55],u_xpb_out[59][55],u_xpb_out[60][55],u_xpb_out[61][55],u_xpb_out[62][55],u_xpb_out[63][55],u_xpb_out[64][55],u_xpb_out[65][55],u_xpb_out[66][55],u_xpb_out[67][55],u_xpb_out[68][55],u_xpb_out[69][55],u_xpb_out[70][55],u_xpb_out[71][55],u_xpb_out[72][55],u_xpb_out[73][55],u_xpb_out[74][55],u_xpb_out[75][55],u_xpb_out[76][55],u_xpb_out[77][55],u_xpb_out[78][55],u_xpb_out[79][55],u_xpb_out[80][55],u_xpb_out[81][55],u_xpb_out[82][55],u_xpb_out[83][55],u_xpb_out[84][55],u_xpb_out[85][55],u_xpb_out[86][55],u_xpb_out[87][55],u_xpb_out[88][55],u_xpb_out[89][55],u_xpb_out[90][55],u_xpb_out[91][55],u_xpb_out[92][55],u_xpb_out[93][55],u_xpb_out[94][55],u_xpb_out[95][55],u_xpb_out[96][55],u_xpb_out[97][55],u_xpb_out[98][55],u_xpb_out[99][55],u_xpb_out[100][55],u_xpb_out[101][55],u_xpb_out[102][55],u_xpb_out[103][55],u_xpb_out[104][55],u_xpb_out[105][55]};

assign col_out_56 = {u_xpb_out[0][56],u_xpb_out[1][56],u_xpb_out[2][56],u_xpb_out[3][56],u_xpb_out[4][56],u_xpb_out[5][56],u_xpb_out[6][56],u_xpb_out[7][56],u_xpb_out[8][56],u_xpb_out[9][56],u_xpb_out[10][56],u_xpb_out[11][56],u_xpb_out[12][56],u_xpb_out[13][56],u_xpb_out[14][56],u_xpb_out[15][56],u_xpb_out[16][56],u_xpb_out[17][56],u_xpb_out[18][56],u_xpb_out[19][56],u_xpb_out[20][56],u_xpb_out[21][56],u_xpb_out[22][56],u_xpb_out[23][56],u_xpb_out[24][56],u_xpb_out[25][56],u_xpb_out[26][56],u_xpb_out[27][56],u_xpb_out[28][56],u_xpb_out[29][56],u_xpb_out[30][56],u_xpb_out[31][56],u_xpb_out[32][56],u_xpb_out[33][56],u_xpb_out[34][56],u_xpb_out[35][56],u_xpb_out[36][56],u_xpb_out[37][56],u_xpb_out[38][56],u_xpb_out[39][56],u_xpb_out[40][56],u_xpb_out[41][56],u_xpb_out[42][56],u_xpb_out[43][56],u_xpb_out[44][56],u_xpb_out[45][56],u_xpb_out[46][56],u_xpb_out[47][56],u_xpb_out[48][56],u_xpb_out[49][56],u_xpb_out[50][56],u_xpb_out[51][56],u_xpb_out[52][56],u_xpb_out[53][56],u_xpb_out[54][56],u_xpb_out[55][56],u_xpb_out[56][56],u_xpb_out[57][56],u_xpb_out[58][56],u_xpb_out[59][56],u_xpb_out[60][56],u_xpb_out[61][56],u_xpb_out[62][56],u_xpb_out[63][56],u_xpb_out[64][56],u_xpb_out[65][56],u_xpb_out[66][56],u_xpb_out[67][56],u_xpb_out[68][56],u_xpb_out[69][56],u_xpb_out[70][56],u_xpb_out[71][56],u_xpb_out[72][56],u_xpb_out[73][56],u_xpb_out[74][56],u_xpb_out[75][56],u_xpb_out[76][56],u_xpb_out[77][56],u_xpb_out[78][56],u_xpb_out[79][56],u_xpb_out[80][56],u_xpb_out[81][56],u_xpb_out[82][56],u_xpb_out[83][56],u_xpb_out[84][56],u_xpb_out[85][56],u_xpb_out[86][56],u_xpb_out[87][56],u_xpb_out[88][56],u_xpb_out[89][56],u_xpb_out[90][56],u_xpb_out[91][56],u_xpb_out[92][56],u_xpb_out[93][56],u_xpb_out[94][56],u_xpb_out[95][56],u_xpb_out[96][56],u_xpb_out[97][56],u_xpb_out[98][56],u_xpb_out[99][56],u_xpb_out[100][56],u_xpb_out[101][56],u_xpb_out[102][56],u_xpb_out[103][56],u_xpb_out[104][56],u_xpb_out[105][56]};

assign col_out_57 = {u_xpb_out[0][57],u_xpb_out[1][57],u_xpb_out[2][57],u_xpb_out[3][57],u_xpb_out[4][57],u_xpb_out[5][57],u_xpb_out[6][57],u_xpb_out[7][57],u_xpb_out[8][57],u_xpb_out[9][57],u_xpb_out[10][57],u_xpb_out[11][57],u_xpb_out[12][57],u_xpb_out[13][57],u_xpb_out[14][57],u_xpb_out[15][57],u_xpb_out[16][57],u_xpb_out[17][57],u_xpb_out[18][57],u_xpb_out[19][57],u_xpb_out[20][57],u_xpb_out[21][57],u_xpb_out[22][57],u_xpb_out[23][57],u_xpb_out[24][57],u_xpb_out[25][57],u_xpb_out[26][57],u_xpb_out[27][57],u_xpb_out[28][57],u_xpb_out[29][57],u_xpb_out[30][57],u_xpb_out[31][57],u_xpb_out[32][57],u_xpb_out[33][57],u_xpb_out[34][57],u_xpb_out[35][57],u_xpb_out[36][57],u_xpb_out[37][57],u_xpb_out[38][57],u_xpb_out[39][57],u_xpb_out[40][57],u_xpb_out[41][57],u_xpb_out[42][57],u_xpb_out[43][57],u_xpb_out[44][57],u_xpb_out[45][57],u_xpb_out[46][57],u_xpb_out[47][57],u_xpb_out[48][57],u_xpb_out[49][57],u_xpb_out[50][57],u_xpb_out[51][57],u_xpb_out[52][57],u_xpb_out[53][57],u_xpb_out[54][57],u_xpb_out[55][57],u_xpb_out[56][57],u_xpb_out[57][57],u_xpb_out[58][57],u_xpb_out[59][57],u_xpb_out[60][57],u_xpb_out[61][57],u_xpb_out[62][57],u_xpb_out[63][57],u_xpb_out[64][57],u_xpb_out[65][57],u_xpb_out[66][57],u_xpb_out[67][57],u_xpb_out[68][57],u_xpb_out[69][57],u_xpb_out[70][57],u_xpb_out[71][57],u_xpb_out[72][57],u_xpb_out[73][57],u_xpb_out[74][57],u_xpb_out[75][57],u_xpb_out[76][57],u_xpb_out[77][57],u_xpb_out[78][57],u_xpb_out[79][57],u_xpb_out[80][57],u_xpb_out[81][57],u_xpb_out[82][57],u_xpb_out[83][57],u_xpb_out[84][57],u_xpb_out[85][57],u_xpb_out[86][57],u_xpb_out[87][57],u_xpb_out[88][57],u_xpb_out[89][57],u_xpb_out[90][57],u_xpb_out[91][57],u_xpb_out[92][57],u_xpb_out[93][57],u_xpb_out[94][57],u_xpb_out[95][57],u_xpb_out[96][57],u_xpb_out[97][57],u_xpb_out[98][57],u_xpb_out[99][57],u_xpb_out[100][57],u_xpb_out[101][57],u_xpb_out[102][57],u_xpb_out[103][57],u_xpb_out[104][57],u_xpb_out[105][57]};

assign col_out_58 = {u_xpb_out[0][58],u_xpb_out[1][58],u_xpb_out[2][58],u_xpb_out[3][58],u_xpb_out[4][58],u_xpb_out[5][58],u_xpb_out[6][58],u_xpb_out[7][58],u_xpb_out[8][58],u_xpb_out[9][58],u_xpb_out[10][58],u_xpb_out[11][58],u_xpb_out[12][58],u_xpb_out[13][58],u_xpb_out[14][58],u_xpb_out[15][58],u_xpb_out[16][58],u_xpb_out[17][58],u_xpb_out[18][58],u_xpb_out[19][58],u_xpb_out[20][58],u_xpb_out[21][58],u_xpb_out[22][58],u_xpb_out[23][58],u_xpb_out[24][58],u_xpb_out[25][58],u_xpb_out[26][58],u_xpb_out[27][58],u_xpb_out[28][58],u_xpb_out[29][58],u_xpb_out[30][58],u_xpb_out[31][58],u_xpb_out[32][58],u_xpb_out[33][58],u_xpb_out[34][58],u_xpb_out[35][58],u_xpb_out[36][58],u_xpb_out[37][58],u_xpb_out[38][58],u_xpb_out[39][58],u_xpb_out[40][58],u_xpb_out[41][58],u_xpb_out[42][58],u_xpb_out[43][58],u_xpb_out[44][58],u_xpb_out[45][58],u_xpb_out[46][58],u_xpb_out[47][58],u_xpb_out[48][58],u_xpb_out[49][58],u_xpb_out[50][58],u_xpb_out[51][58],u_xpb_out[52][58],u_xpb_out[53][58],u_xpb_out[54][58],u_xpb_out[55][58],u_xpb_out[56][58],u_xpb_out[57][58],u_xpb_out[58][58],u_xpb_out[59][58],u_xpb_out[60][58],u_xpb_out[61][58],u_xpb_out[62][58],u_xpb_out[63][58],u_xpb_out[64][58],u_xpb_out[65][58],u_xpb_out[66][58],u_xpb_out[67][58],u_xpb_out[68][58],u_xpb_out[69][58],u_xpb_out[70][58],u_xpb_out[71][58],u_xpb_out[72][58],u_xpb_out[73][58],u_xpb_out[74][58],u_xpb_out[75][58],u_xpb_out[76][58],u_xpb_out[77][58],u_xpb_out[78][58],u_xpb_out[79][58],u_xpb_out[80][58],u_xpb_out[81][58],u_xpb_out[82][58],u_xpb_out[83][58],u_xpb_out[84][58],u_xpb_out[85][58],u_xpb_out[86][58],u_xpb_out[87][58],u_xpb_out[88][58],u_xpb_out[89][58],u_xpb_out[90][58],u_xpb_out[91][58],u_xpb_out[92][58],u_xpb_out[93][58],u_xpb_out[94][58],u_xpb_out[95][58],u_xpb_out[96][58],u_xpb_out[97][58],u_xpb_out[98][58],u_xpb_out[99][58],u_xpb_out[100][58],u_xpb_out[101][58],u_xpb_out[102][58],u_xpb_out[103][58],u_xpb_out[104][58],u_xpb_out[105][58]};

assign col_out_59 = {u_xpb_out[0][59],u_xpb_out[1][59],u_xpb_out[2][59],u_xpb_out[3][59],u_xpb_out[4][59],u_xpb_out[5][59],u_xpb_out[6][59],u_xpb_out[7][59],u_xpb_out[8][59],u_xpb_out[9][59],u_xpb_out[10][59],u_xpb_out[11][59],u_xpb_out[12][59],u_xpb_out[13][59],u_xpb_out[14][59],u_xpb_out[15][59],u_xpb_out[16][59],u_xpb_out[17][59],u_xpb_out[18][59],u_xpb_out[19][59],u_xpb_out[20][59],u_xpb_out[21][59],u_xpb_out[22][59],u_xpb_out[23][59],u_xpb_out[24][59],u_xpb_out[25][59],u_xpb_out[26][59],u_xpb_out[27][59],u_xpb_out[28][59],u_xpb_out[29][59],u_xpb_out[30][59],u_xpb_out[31][59],u_xpb_out[32][59],u_xpb_out[33][59],u_xpb_out[34][59],u_xpb_out[35][59],u_xpb_out[36][59],u_xpb_out[37][59],u_xpb_out[38][59],u_xpb_out[39][59],u_xpb_out[40][59],u_xpb_out[41][59],u_xpb_out[42][59],u_xpb_out[43][59],u_xpb_out[44][59],u_xpb_out[45][59],u_xpb_out[46][59],u_xpb_out[47][59],u_xpb_out[48][59],u_xpb_out[49][59],u_xpb_out[50][59],u_xpb_out[51][59],u_xpb_out[52][59],u_xpb_out[53][59],u_xpb_out[54][59],u_xpb_out[55][59],u_xpb_out[56][59],u_xpb_out[57][59],u_xpb_out[58][59],u_xpb_out[59][59],u_xpb_out[60][59],u_xpb_out[61][59],u_xpb_out[62][59],u_xpb_out[63][59],u_xpb_out[64][59],u_xpb_out[65][59],u_xpb_out[66][59],u_xpb_out[67][59],u_xpb_out[68][59],u_xpb_out[69][59],u_xpb_out[70][59],u_xpb_out[71][59],u_xpb_out[72][59],u_xpb_out[73][59],u_xpb_out[74][59],u_xpb_out[75][59],u_xpb_out[76][59],u_xpb_out[77][59],u_xpb_out[78][59],u_xpb_out[79][59],u_xpb_out[80][59],u_xpb_out[81][59],u_xpb_out[82][59],u_xpb_out[83][59],u_xpb_out[84][59],u_xpb_out[85][59],u_xpb_out[86][59],u_xpb_out[87][59],u_xpb_out[88][59],u_xpb_out[89][59],u_xpb_out[90][59],u_xpb_out[91][59],u_xpb_out[92][59],u_xpb_out[93][59],u_xpb_out[94][59],u_xpb_out[95][59],u_xpb_out[96][59],u_xpb_out[97][59],u_xpb_out[98][59],u_xpb_out[99][59],u_xpb_out[100][59],u_xpb_out[101][59],u_xpb_out[102][59],u_xpb_out[103][59],u_xpb_out[104][59],u_xpb_out[105][59]};

assign col_out_60 = {u_xpb_out[0][60],u_xpb_out[1][60],u_xpb_out[2][60],u_xpb_out[3][60],u_xpb_out[4][60],u_xpb_out[5][60],u_xpb_out[6][60],u_xpb_out[7][60],u_xpb_out[8][60],u_xpb_out[9][60],u_xpb_out[10][60],u_xpb_out[11][60],u_xpb_out[12][60],u_xpb_out[13][60],u_xpb_out[14][60],u_xpb_out[15][60],u_xpb_out[16][60],u_xpb_out[17][60],u_xpb_out[18][60],u_xpb_out[19][60],u_xpb_out[20][60],u_xpb_out[21][60],u_xpb_out[22][60],u_xpb_out[23][60],u_xpb_out[24][60],u_xpb_out[25][60],u_xpb_out[26][60],u_xpb_out[27][60],u_xpb_out[28][60],u_xpb_out[29][60],u_xpb_out[30][60],u_xpb_out[31][60],u_xpb_out[32][60],u_xpb_out[33][60],u_xpb_out[34][60],u_xpb_out[35][60],u_xpb_out[36][60],u_xpb_out[37][60],u_xpb_out[38][60],u_xpb_out[39][60],u_xpb_out[40][60],u_xpb_out[41][60],u_xpb_out[42][60],u_xpb_out[43][60],u_xpb_out[44][60],u_xpb_out[45][60],u_xpb_out[46][60],u_xpb_out[47][60],u_xpb_out[48][60],u_xpb_out[49][60],u_xpb_out[50][60],u_xpb_out[51][60],u_xpb_out[52][60],u_xpb_out[53][60],u_xpb_out[54][60],u_xpb_out[55][60],u_xpb_out[56][60],u_xpb_out[57][60],u_xpb_out[58][60],u_xpb_out[59][60],u_xpb_out[60][60],u_xpb_out[61][60],u_xpb_out[62][60],u_xpb_out[63][60],u_xpb_out[64][60],u_xpb_out[65][60],u_xpb_out[66][60],u_xpb_out[67][60],u_xpb_out[68][60],u_xpb_out[69][60],u_xpb_out[70][60],u_xpb_out[71][60],u_xpb_out[72][60],u_xpb_out[73][60],u_xpb_out[74][60],u_xpb_out[75][60],u_xpb_out[76][60],u_xpb_out[77][60],u_xpb_out[78][60],u_xpb_out[79][60],u_xpb_out[80][60],u_xpb_out[81][60],u_xpb_out[82][60],u_xpb_out[83][60],u_xpb_out[84][60],u_xpb_out[85][60],u_xpb_out[86][60],u_xpb_out[87][60],u_xpb_out[88][60],u_xpb_out[89][60],u_xpb_out[90][60],u_xpb_out[91][60],u_xpb_out[92][60],u_xpb_out[93][60],u_xpb_out[94][60],u_xpb_out[95][60],u_xpb_out[96][60],u_xpb_out[97][60],u_xpb_out[98][60],u_xpb_out[99][60],u_xpb_out[100][60],u_xpb_out[101][60],u_xpb_out[102][60],u_xpb_out[103][60],u_xpb_out[104][60],u_xpb_out[105][60]};

assign col_out_61 = {u_xpb_out[0][61],u_xpb_out[1][61],u_xpb_out[2][61],u_xpb_out[3][61],u_xpb_out[4][61],u_xpb_out[5][61],u_xpb_out[6][61],u_xpb_out[7][61],u_xpb_out[8][61],u_xpb_out[9][61],u_xpb_out[10][61],u_xpb_out[11][61],u_xpb_out[12][61],u_xpb_out[13][61],u_xpb_out[14][61],u_xpb_out[15][61],u_xpb_out[16][61],u_xpb_out[17][61],u_xpb_out[18][61],u_xpb_out[19][61],u_xpb_out[20][61],u_xpb_out[21][61],u_xpb_out[22][61],u_xpb_out[23][61],u_xpb_out[24][61],u_xpb_out[25][61],u_xpb_out[26][61],u_xpb_out[27][61],u_xpb_out[28][61],u_xpb_out[29][61],u_xpb_out[30][61],u_xpb_out[31][61],u_xpb_out[32][61],u_xpb_out[33][61],u_xpb_out[34][61],u_xpb_out[35][61],u_xpb_out[36][61],u_xpb_out[37][61],u_xpb_out[38][61],u_xpb_out[39][61],u_xpb_out[40][61],u_xpb_out[41][61],u_xpb_out[42][61],u_xpb_out[43][61],u_xpb_out[44][61],u_xpb_out[45][61],u_xpb_out[46][61],u_xpb_out[47][61],u_xpb_out[48][61],u_xpb_out[49][61],u_xpb_out[50][61],u_xpb_out[51][61],u_xpb_out[52][61],u_xpb_out[53][61],u_xpb_out[54][61],u_xpb_out[55][61],u_xpb_out[56][61],u_xpb_out[57][61],u_xpb_out[58][61],u_xpb_out[59][61],u_xpb_out[60][61],u_xpb_out[61][61],u_xpb_out[62][61],u_xpb_out[63][61],u_xpb_out[64][61],u_xpb_out[65][61],u_xpb_out[66][61],u_xpb_out[67][61],u_xpb_out[68][61],u_xpb_out[69][61],u_xpb_out[70][61],u_xpb_out[71][61],u_xpb_out[72][61],u_xpb_out[73][61],u_xpb_out[74][61],u_xpb_out[75][61],u_xpb_out[76][61],u_xpb_out[77][61],u_xpb_out[78][61],u_xpb_out[79][61],u_xpb_out[80][61],u_xpb_out[81][61],u_xpb_out[82][61],u_xpb_out[83][61],u_xpb_out[84][61],u_xpb_out[85][61],u_xpb_out[86][61],u_xpb_out[87][61],u_xpb_out[88][61],u_xpb_out[89][61],u_xpb_out[90][61],u_xpb_out[91][61],u_xpb_out[92][61],u_xpb_out[93][61],u_xpb_out[94][61],u_xpb_out[95][61],u_xpb_out[96][61],u_xpb_out[97][61],u_xpb_out[98][61],u_xpb_out[99][61],u_xpb_out[100][61],u_xpb_out[101][61],u_xpb_out[102][61],u_xpb_out[103][61],u_xpb_out[104][61],u_xpb_out[105][61]};

assign col_out_62 = {u_xpb_out[0][62],u_xpb_out[1][62],u_xpb_out[2][62],u_xpb_out[3][62],u_xpb_out[4][62],u_xpb_out[5][62],u_xpb_out[6][62],u_xpb_out[7][62],u_xpb_out[8][62],u_xpb_out[9][62],u_xpb_out[10][62],u_xpb_out[11][62],u_xpb_out[12][62],u_xpb_out[13][62],u_xpb_out[14][62],u_xpb_out[15][62],u_xpb_out[16][62],u_xpb_out[17][62],u_xpb_out[18][62],u_xpb_out[19][62],u_xpb_out[20][62],u_xpb_out[21][62],u_xpb_out[22][62],u_xpb_out[23][62],u_xpb_out[24][62],u_xpb_out[25][62],u_xpb_out[26][62],u_xpb_out[27][62],u_xpb_out[28][62],u_xpb_out[29][62],u_xpb_out[30][62],u_xpb_out[31][62],u_xpb_out[32][62],u_xpb_out[33][62],u_xpb_out[34][62],u_xpb_out[35][62],u_xpb_out[36][62],u_xpb_out[37][62],u_xpb_out[38][62],u_xpb_out[39][62],u_xpb_out[40][62],u_xpb_out[41][62],u_xpb_out[42][62],u_xpb_out[43][62],u_xpb_out[44][62],u_xpb_out[45][62],u_xpb_out[46][62],u_xpb_out[47][62],u_xpb_out[48][62],u_xpb_out[49][62],u_xpb_out[50][62],u_xpb_out[51][62],u_xpb_out[52][62],u_xpb_out[53][62],u_xpb_out[54][62],u_xpb_out[55][62],u_xpb_out[56][62],u_xpb_out[57][62],u_xpb_out[58][62],u_xpb_out[59][62],u_xpb_out[60][62],u_xpb_out[61][62],u_xpb_out[62][62],u_xpb_out[63][62],u_xpb_out[64][62],u_xpb_out[65][62],u_xpb_out[66][62],u_xpb_out[67][62],u_xpb_out[68][62],u_xpb_out[69][62],u_xpb_out[70][62],u_xpb_out[71][62],u_xpb_out[72][62],u_xpb_out[73][62],u_xpb_out[74][62],u_xpb_out[75][62],u_xpb_out[76][62],u_xpb_out[77][62],u_xpb_out[78][62],u_xpb_out[79][62],u_xpb_out[80][62],u_xpb_out[81][62],u_xpb_out[82][62],u_xpb_out[83][62],u_xpb_out[84][62],u_xpb_out[85][62],u_xpb_out[86][62],u_xpb_out[87][62],u_xpb_out[88][62],u_xpb_out[89][62],u_xpb_out[90][62],u_xpb_out[91][62],u_xpb_out[92][62],u_xpb_out[93][62],u_xpb_out[94][62],u_xpb_out[95][62],u_xpb_out[96][62],u_xpb_out[97][62],u_xpb_out[98][62],u_xpb_out[99][62],u_xpb_out[100][62],u_xpb_out[101][62],u_xpb_out[102][62],u_xpb_out[103][62],u_xpb_out[104][62],u_xpb_out[105][62]};

assign col_out_63 = {u_xpb_out[0][63],u_xpb_out[1][63],u_xpb_out[2][63],u_xpb_out[3][63],u_xpb_out[4][63],u_xpb_out[5][63],u_xpb_out[6][63],u_xpb_out[7][63],u_xpb_out[8][63],u_xpb_out[9][63],u_xpb_out[10][63],u_xpb_out[11][63],u_xpb_out[12][63],u_xpb_out[13][63],u_xpb_out[14][63],u_xpb_out[15][63],u_xpb_out[16][63],u_xpb_out[17][63],u_xpb_out[18][63],u_xpb_out[19][63],u_xpb_out[20][63],u_xpb_out[21][63],u_xpb_out[22][63],u_xpb_out[23][63],u_xpb_out[24][63],u_xpb_out[25][63],u_xpb_out[26][63],u_xpb_out[27][63],u_xpb_out[28][63],u_xpb_out[29][63],u_xpb_out[30][63],u_xpb_out[31][63],u_xpb_out[32][63],u_xpb_out[33][63],u_xpb_out[34][63],u_xpb_out[35][63],u_xpb_out[36][63],u_xpb_out[37][63],u_xpb_out[38][63],u_xpb_out[39][63],u_xpb_out[40][63],u_xpb_out[41][63],u_xpb_out[42][63],u_xpb_out[43][63],u_xpb_out[44][63],u_xpb_out[45][63],u_xpb_out[46][63],u_xpb_out[47][63],u_xpb_out[48][63],u_xpb_out[49][63],u_xpb_out[50][63],u_xpb_out[51][63],u_xpb_out[52][63],u_xpb_out[53][63],u_xpb_out[54][63],u_xpb_out[55][63],u_xpb_out[56][63],u_xpb_out[57][63],u_xpb_out[58][63],u_xpb_out[59][63],u_xpb_out[60][63],u_xpb_out[61][63],u_xpb_out[62][63],u_xpb_out[63][63],u_xpb_out[64][63],u_xpb_out[65][63],u_xpb_out[66][63],u_xpb_out[67][63],u_xpb_out[68][63],u_xpb_out[69][63],u_xpb_out[70][63],u_xpb_out[71][63],u_xpb_out[72][63],u_xpb_out[73][63],u_xpb_out[74][63],u_xpb_out[75][63],u_xpb_out[76][63],u_xpb_out[77][63],u_xpb_out[78][63],u_xpb_out[79][63],u_xpb_out[80][63],u_xpb_out[81][63],u_xpb_out[82][63],u_xpb_out[83][63],u_xpb_out[84][63],u_xpb_out[85][63],u_xpb_out[86][63],u_xpb_out[87][63],u_xpb_out[88][63],u_xpb_out[89][63],u_xpb_out[90][63],u_xpb_out[91][63],u_xpb_out[92][63],u_xpb_out[93][63],u_xpb_out[94][63],u_xpb_out[95][63],u_xpb_out[96][63],u_xpb_out[97][63],u_xpb_out[98][63],u_xpb_out[99][63],u_xpb_out[100][63],u_xpb_out[101][63],u_xpb_out[102][63],u_xpb_out[103][63],u_xpb_out[104][63],u_xpb_out[105][63]};

assign col_out_64 = {u_xpb_out[0][64],u_xpb_out[1][64],u_xpb_out[2][64],u_xpb_out[3][64],u_xpb_out[4][64],u_xpb_out[5][64],u_xpb_out[6][64],u_xpb_out[7][64],u_xpb_out[8][64],u_xpb_out[9][64],u_xpb_out[10][64],u_xpb_out[11][64],u_xpb_out[12][64],u_xpb_out[13][64],u_xpb_out[14][64],u_xpb_out[15][64],u_xpb_out[16][64],u_xpb_out[17][64],u_xpb_out[18][64],u_xpb_out[19][64],u_xpb_out[20][64],u_xpb_out[21][64],u_xpb_out[22][64],u_xpb_out[23][64],u_xpb_out[24][64],u_xpb_out[25][64],u_xpb_out[26][64],u_xpb_out[27][64],u_xpb_out[28][64],u_xpb_out[29][64],u_xpb_out[30][64],u_xpb_out[31][64],u_xpb_out[32][64],u_xpb_out[33][64],u_xpb_out[34][64],u_xpb_out[35][64],u_xpb_out[36][64],u_xpb_out[37][64],u_xpb_out[38][64],u_xpb_out[39][64],u_xpb_out[40][64],u_xpb_out[41][64],u_xpb_out[42][64],u_xpb_out[43][64],u_xpb_out[44][64],u_xpb_out[45][64],u_xpb_out[46][64],u_xpb_out[47][64],u_xpb_out[48][64],u_xpb_out[49][64],u_xpb_out[50][64],u_xpb_out[51][64],u_xpb_out[52][64],u_xpb_out[53][64],u_xpb_out[54][64],u_xpb_out[55][64],u_xpb_out[56][64],u_xpb_out[57][64],u_xpb_out[58][64],u_xpb_out[59][64],u_xpb_out[60][64],u_xpb_out[61][64],u_xpb_out[62][64],u_xpb_out[63][64],u_xpb_out[64][64],u_xpb_out[65][64],u_xpb_out[66][64],u_xpb_out[67][64],u_xpb_out[68][64],u_xpb_out[69][64],u_xpb_out[70][64],u_xpb_out[71][64],u_xpb_out[72][64],u_xpb_out[73][64],u_xpb_out[74][64],u_xpb_out[75][64],u_xpb_out[76][64],u_xpb_out[77][64],u_xpb_out[78][64],u_xpb_out[79][64],u_xpb_out[80][64],u_xpb_out[81][64],u_xpb_out[82][64],u_xpb_out[83][64],u_xpb_out[84][64],u_xpb_out[85][64],u_xpb_out[86][64],u_xpb_out[87][64],u_xpb_out[88][64],u_xpb_out[89][64],u_xpb_out[90][64],u_xpb_out[91][64],u_xpb_out[92][64],u_xpb_out[93][64],u_xpb_out[94][64],u_xpb_out[95][64],u_xpb_out[96][64],u_xpb_out[97][64],u_xpb_out[98][64],u_xpb_out[99][64],u_xpb_out[100][64],u_xpb_out[101][64],u_xpb_out[102][64],u_xpb_out[103][64],u_xpb_out[104][64],u_xpb_out[105][64]};

assign col_out_65 = {u_xpb_out[0][65],u_xpb_out[1][65],u_xpb_out[2][65],u_xpb_out[3][65],u_xpb_out[4][65],u_xpb_out[5][65],u_xpb_out[6][65],u_xpb_out[7][65],u_xpb_out[8][65],u_xpb_out[9][65],u_xpb_out[10][65],u_xpb_out[11][65],u_xpb_out[12][65],u_xpb_out[13][65],u_xpb_out[14][65],u_xpb_out[15][65],u_xpb_out[16][65],u_xpb_out[17][65],u_xpb_out[18][65],u_xpb_out[19][65],u_xpb_out[20][65],u_xpb_out[21][65],u_xpb_out[22][65],u_xpb_out[23][65],u_xpb_out[24][65],u_xpb_out[25][65],u_xpb_out[26][65],u_xpb_out[27][65],u_xpb_out[28][65],u_xpb_out[29][65],u_xpb_out[30][65],u_xpb_out[31][65],u_xpb_out[32][65],u_xpb_out[33][65],u_xpb_out[34][65],u_xpb_out[35][65],u_xpb_out[36][65],u_xpb_out[37][65],u_xpb_out[38][65],u_xpb_out[39][65],u_xpb_out[40][65],u_xpb_out[41][65],u_xpb_out[42][65],u_xpb_out[43][65],u_xpb_out[44][65],u_xpb_out[45][65],u_xpb_out[46][65],u_xpb_out[47][65],u_xpb_out[48][65],u_xpb_out[49][65],u_xpb_out[50][65],u_xpb_out[51][65],u_xpb_out[52][65],u_xpb_out[53][65],u_xpb_out[54][65],u_xpb_out[55][65],u_xpb_out[56][65],u_xpb_out[57][65],u_xpb_out[58][65],u_xpb_out[59][65],u_xpb_out[60][65],u_xpb_out[61][65],u_xpb_out[62][65],u_xpb_out[63][65],u_xpb_out[64][65],u_xpb_out[65][65],u_xpb_out[66][65],u_xpb_out[67][65],u_xpb_out[68][65],u_xpb_out[69][65],u_xpb_out[70][65],u_xpb_out[71][65],u_xpb_out[72][65],u_xpb_out[73][65],u_xpb_out[74][65],u_xpb_out[75][65],u_xpb_out[76][65],u_xpb_out[77][65],u_xpb_out[78][65],u_xpb_out[79][65],u_xpb_out[80][65],u_xpb_out[81][65],u_xpb_out[82][65],u_xpb_out[83][65],u_xpb_out[84][65],u_xpb_out[85][65],u_xpb_out[86][65],u_xpb_out[87][65],u_xpb_out[88][65],u_xpb_out[89][65],u_xpb_out[90][65],u_xpb_out[91][65],u_xpb_out[92][65],u_xpb_out[93][65],u_xpb_out[94][65],u_xpb_out[95][65],u_xpb_out[96][65],u_xpb_out[97][65],u_xpb_out[98][65],u_xpb_out[99][65],u_xpb_out[100][65],u_xpb_out[101][65],u_xpb_out[102][65],u_xpb_out[103][65],u_xpb_out[104][65],u_xpb_out[105][65]};

assign col_out_66 = {u_xpb_out[0][66],u_xpb_out[1][66],u_xpb_out[2][66],u_xpb_out[3][66],u_xpb_out[4][66],u_xpb_out[5][66],u_xpb_out[6][66],u_xpb_out[7][66],u_xpb_out[8][66],u_xpb_out[9][66],u_xpb_out[10][66],u_xpb_out[11][66],u_xpb_out[12][66],u_xpb_out[13][66],u_xpb_out[14][66],u_xpb_out[15][66],u_xpb_out[16][66],u_xpb_out[17][66],u_xpb_out[18][66],u_xpb_out[19][66],u_xpb_out[20][66],u_xpb_out[21][66],u_xpb_out[22][66],u_xpb_out[23][66],u_xpb_out[24][66],u_xpb_out[25][66],u_xpb_out[26][66],u_xpb_out[27][66],u_xpb_out[28][66],u_xpb_out[29][66],u_xpb_out[30][66],u_xpb_out[31][66],u_xpb_out[32][66],u_xpb_out[33][66],u_xpb_out[34][66],u_xpb_out[35][66],u_xpb_out[36][66],u_xpb_out[37][66],u_xpb_out[38][66],u_xpb_out[39][66],u_xpb_out[40][66],u_xpb_out[41][66],u_xpb_out[42][66],u_xpb_out[43][66],u_xpb_out[44][66],u_xpb_out[45][66],u_xpb_out[46][66],u_xpb_out[47][66],u_xpb_out[48][66],u_xpb_out[49][66],u_xpb_out[50][66],u_xpb_out[51][66],u_xpb_out[52][66],u_xpb_out[53][66],u_xpb_out[54][66],u_xpb_out[55][66],u_xpb_out[56][66],u_xpb_out[57][66],u_xpb_out[58][66],u_xpb_out[59][66],u_xpb_out[60][66],u_xpb_out[61][66],u_xpb_out[62][66],u_xpb_out[63][66],u_xpb_out[64][66],u_xpb_out[65][66],u_xpb_out[66][66],u_xpb_out[67][66],u_xpb_out[68][66],u_xpb_out[69][66],u_xpb_out[70][66],u_xpb_out[71][66],u_xpb_out[72][66],u_xpb_out[73][66],u_xpb_out[74][66],u_xpb_out[75][66],u_xpb_out[76][66],u_xpb_out[77][66],u_xpb_out[78][66],u_xpb_out[79][66],u_xpb_out[80][66],u_xpb_out[81][66],u_xpb_out[82][66],u_xpb_out[83][66],u_xpb_out[84][66],u_xpb_out[85][66],u_xpb_out[86][66],u_xpb_out[87][66],u_xpb_out[88][66],u_xpb_out[89][66],u_xpb_out[90][66],u_xpb_out[91][66],u_xpb_out[92][66],u_xpb_out[93][66],u_xpb_out[94][66],u_xpb_out[95][66],u_xpb_out[96][66],u_xpb_out[97][66],u_xpb_out[98][66],u_xpb_out[99][66],u_xpb_out[100][66],u_xpb_out[101][66],u_xpb_out[102][66],u_xpb_out[103][66],u_xpb_out[104][66],u_xpb_out[105][66]};

assign col_out_67 = {u_xpb_out[0][67],u_xpb_out[1][67],u_xpb_out[2][67],u_xpb_out[3][67],u_xpb_out[4][67],u_xpb_out[5][67],u_xpb_out[6][67],u_xpb_out[7][67],u_xpb_out[8][67],u_xpb_out[9][67],u_xpb_out[10][67],u_xpb_out[11][67],u_xpb_out[12][67],u_xpb_out[13][67],u_xpb_out[14][67],u_xpb_out[15][67],u_xpb_out[16][67],u_xpb_out[17][67],u_xpb_out[18][67],u_xpb_out[19][67],u_xpb_out[20][67],u_xpb_out[21][67],u_xpb_out[22][67],u_xpb_out[23][67],u_xpb_out[24][67],u_xpb_out[25][67],u_xpb_out[26][67],u_xpb_out[27][67],u_xpb_out[28][67],u_xpb_out[29][67],u_xpb_out[30][67],u_xpb_out[31][67],u_xpb_out[32][67],u_xpb_out[33][67],u_xpb_out[34][67],u_xpb_out[35][67],u_xpb_out[36][67],u_xpb_out[37][67],u_xpb_out[38][67],u_xpb_out[39][67],u_xpb_out[40][67],u_xpb_out[41][67],u_xpb_out[42][67],u_xpb_out[43][67],u_xpb_out[44][67],u_xpb_out[45][67],u_xpb_out[46][67],u_xpb_out[47][67],u_xpb_out[48][67],u_xpb_out[49][67],u_xpb_out[50][67],u_xpb_out[51][67],u_xpb_out[52][67],u_xpb_out[53][67],u_xpb_out[54][67],u_xpb_out[55][67],u_xpb_out[56][67],u_xpb_out[57][67],u_xpb_out[58][67],u_xpb_out[59][67],u_xpb_out[60][67],u_xpb_out[61][67],u_xpb_out[62][67],u_xpb_out[63][67],u_xpb_out[64][67],u_xpb_out[65][67],u_xpb_out[66][67],u_xpb_out[67][67],u_xpb_out[68][67],u_xpb_out[69][67],u_xpb_out[70][67],u_xpb_out[71][67],u_xpb_out[72][67],u_xpb_out[73][67],u_xpb_out[74][67],u_xpb_out[75][67],u_xpb_out[76][67],u_xpb_out[77][67],u_xpb_out[78][67],u_xpb_out[79][67],u_xpb_out[80][67],u_xpb_out[81][67],u_xpb_out[82][67],u_xpb_out[83][67],u_xpb_out[84][67],u_xpb_out[85][67],u_xpb_out[86][67],u_xpb_out[87][67],u_xpb_out[88][67],u_xpb_out[89][67],u_xpb_out[90][67],u_xpb_out[91][67],u_xpb_out[92][67],u_xpb_out[93][67],u_xpb_out[94][67],u_xpb_out[95][67],u_xpb_out[96][67],u_xpb_out[97][67],u_xpb_out[98][67],u_xpb_out[99][67],u_xpb_out[100][67],u_xpb_out[101][67],u_xpb_out[102][67],u_xpb_out[103][67],u_xpb_out[104][67],u_xpb_out[105][67]};

assign col_out_68 = {u_xpb_out[0][68],u_xpb_out[1][68],u_xpb_out[2][68],u_xpb_out[3][68],u_xpb_out[4][68],u_xpb_out[5][68],u_xpb_out[6][68],u_xpb_out[7][68],u_xpb_out[8][68],u_xpb_out[9][68],u_xpb_out[10][68],u_xpb_out[11][68],u_xpb_out[12][68],u_xpb_out[13][68],u_xpb_out[14][68],u_xpb_out[15][68],u_xpb_out[16][68],u_xpb_out[17][68],u_xpb_out[18][68],u_xpb_out[19][68],u_xpb_out[20][68],u_xpb_out[21][68],u_xpb_out[22][68],u_xpb_out[23][68],u_xpb_out[24][68],u_xpb_out[25][68],u_xpb_out[26][68],u_xpb_out[27][68],u_xpb_out[28][68],u_xpb_out[29][68],u_xpb_out[30][68],u_xpb_out[31][68],u_xpb_out[32][68],u_xpb_out[33][68],u_xpb_out[34][68],u_xpb_out[35][68],u_xpb_out[36][68],u_xpb_out[37][68],u_xpb_out[38][68],u_xpb_out[39][68],u_xpb_out[40][68],u_xpb_out[41][68],u_xpb_out[42][68],u_xpb_out[43][68],u_xpb_out[44][68],u_xpb_out[45][68],u_xpb_out[46][68],u_xpb_out[47][68],u_xpb_out[48][68],u_xpb_out[49][68],u_xpb_out[50][68],u_xpb_out[51][68],u_xpb_out[52][68],u_xpb_out[53][68],u_xpb_out[54][68],u_xpb_out[55][68],u_xpb_out[56][68],u_xpb_out[57][68],u_xpb_out[58][68],u_xpb_out[59][68],u_xpb_out[60][68],u_xpb_out[61][68],u_xpb_out[62][68],u_xpb_out[63][68],u_xpb_out[64][68],u_xpb_out[65][68],u_xpb_out[66][68],u_xpb_out[67][68],u_xpb_out[68][68],u_xpb_out[69][68],u_xpb_out[70][68],u_xpb_out[71][68],u_xpb_out[72][68],u_xpb_out[73][68],u_xpb_out[74][68],u_xpb_out[75][68],u_xpb_out[76][68],u_xpb_out[77][68],u_xpb_out[78][68],u_xpb_out[79][68],u_xpb_out[80][68],u_xpb_out[81][68],u_xpb_out[82][68],u_xpb_out[83][68],u_xpb_out[84][68],u_xpb_out[85][68],u_xpb_out[86][68],u_xpb_out[87][68],u_xpb_out[88][68],u_xpb_out[89][68],u_xpb_out[90][68],u_xpb_out[91][68],u_xpb_out[92][68],u_xpb_out[93][68],u_xpb_out[94][68],u_xpb_out[95][68],u_xpb_out[96][68],u_xpb_out[97][68],u_xpb_out[98][68],u_xpb_out[99][68],u_xpb_out[100][68],u_xpb_out[101][68],u_xpb_out[102][68],u_xpb_out[103][68],u_xpb_out[104][68],u_xpb_out[105][68]};

assign col_out_69 = {u_xpb_out[0][69],u_xpb_out[1][69],u_xpb_out[2][69],u_xpb_out[3][69],u_xpb_out[4][69],u_xpb_out[5][69],u_xpb_out[6][69],u_xpb_out[7][69],u_xpb_out[8][69],u_xpb_out[9][69],u_xpb_out[10][69],u_xpb_out[11][69],u_xpb_out[12][69],u_xpb_out[13][69],u_xpb_out[14][69],u_xpb_out[15][69],u_xpb_out[16][69],u_xpb_out[17][69],u_xpb_out[18][69],u_xpb_out[19][69],u_xpb_out[20][69],u_xpb_out[21][69],u_xpb_out[22][69],u_xpb_out[23][69],u_xpb_out[24][69],u_xpb_out[25][69],u_xpb_out[26][69],u_xpb_out[27][69],u_xpb_out[28][69],u_xpb_out[29][69],u_xpb_out[30][69],u_xpb_out[31][69],u_xpb_out[32][69],u_xpb_out[33][69],u_xpb_out[34][69],u_xpb_out[35][69],u_xpb_out[36][69],u_xpb_out[37][69],u_xpb_out[38][69],u_xpb_out[39][69],u_xpb_out[40][69],u_xpb_out[41][69],u_xpb_out[42][69],u_xpb_out[43][69],u_xpb_out[44][69],u_xpb_out[45][69],u_xpb_out[46][69],u_xpb_out[47][69],u_xpb_out[48][69],u_xpb_out[49][69],u_xpb_out[50][69],u_xpb_out[51][69],u_xpb_out[52][69],u_xpb_out[53][69],u_xpb_out[54][69],u_xpb_out[55][69],u_xpb_out[56][69],u_xpb_out[57][69],u_xpb_out[58][69],u_xpb_out[59][69],u_xpb_out[60][69],u_xpb_out[61][69],u_xpb_out[62][69],u_xpb_out[63][69],u_xpb_out[64][69],u_xpb_out[65][69],u_xpb_out[66][69],u_xpb_out[67][69],u_xpb_out[68][69],u_xpb_out[69][69],u_xpb_out[70][69],u_xpb_out[71][69],u_xpb_out[72][69],u_xpb_out[73][69],u_xpb_out[74][69],u_xpb_out[75][69],u_xpb_out[76][69],u_xpb_out[77][69],u_xpb_out[78][69],u_xpb_out[79][69],u_xpb_out[80][69],u_xpb_out[81][69],u_xpb_out[82][69],u_xpb_out[83][69],u_xpb_out[84][69],u_xpb_out[85][69],u_xpb_out[86][69],u_xpb_out[87][69],u_xpb_out[88][69],u_xpb_out[89][69],u_xpb_out[90][69],u_xpb_out[91][69],u_xpb_out[92][69],u_xpb_out[93][69],u_xpb_out[94][69],u_xpb_out[95][69],u_xpb_out[96][69],u_xpb_out[97][69],u_xpb_out[98][69],u_xpb_out[99][69],u_xpb_out[100][69],u_xpb_out[101][69],u_xpb_out[102][69],u_xpb_out[103][69],u_xpb_out[104][69],u_xpb_out[105][69]};

assign col_out_70 = {u_xpb_out[0][70],u_xpb_out[1][70],u_xpb_out[2][70],u_xpb_out[3][70],u_xpb_out[4][70],u_xpb_out[5][70],u_xpb_out[6][70],u_xpb_out[7][70],u_xpb_out[8][70],u_xpb_out[9][70],u_xpb_out[10][70],u_xpb_out[11][70],u_xpb_out[12][70],u_xpb_out[13][70],u_xpb_out[14][70],u_xpb_out[15][70],u_xpb_out[16][70],u_xpb_out[17][70],u_xpb_out[18][70],u_xpb_out[19][70],u_xpb_out[20][70],u_xpb_out[21][70],u_xpb_out[22][70],u_xpb_out[23][70],u_xpb_out[24][70],u_xpb_out[25][70],u_xpb_out[26][70],u_xpb_out[27][70],u_xpb_out[28][70],u_xpb_out[29][70],u_xpb_out[30][70],u_xpb_out[31][70],u_xpb_out[32][70],u_xpb_out[33][70],u_xpb_out[34][70],u_xpb_out[35][70],u_xpb_out[36][70],u_xpb_out[37][70],u_xpb_out[38][70],u_xpb_out[39][70],u_xpb_out[40][70],u_xpb_out[41][70],u_xpb_out[42][70],u_xpb_out[43][70],u_xpb_out[44][70],u_xpb_out[45][70],u_xpb_out[46][70],u_xpb_out[47][70],u_xpb_out[48][70],u_xpb_out[49][70],u_xpb_out[50][70],u_xpb_out[51][70],u_xpb_out[52][70],u_xpb_out[53][70],u_xpb_out[54][70],u_xpb_out[55][70],u_xpb_out[56][70],u_xpb_out[57][70],u_xpb_out[58][70],u_xpb_out[59][70],u_xpb_out[60][70],u_xpb_out[61][70],u_xpb_out[62][70],u_xpb_out[63][70],u_xpb_out[64][70],u_xpb_out[65][70],u_xpb_out[66][70],u_xpb_out[67][70],u_xpb_out[68][70],u_xpb_out[69][70],u_xpb_out[70][70],u_xpb_out[71][70],u_xpb_out[72][70],u_xpb_out[73][70],u_xpb_out[74][70],u_xpb_out[75][70],u_xpb_out[76][70],u_xpb_out[77][70],u_xpb_out[78][70],u_xpb_out[79][70],u_xpb_out[80][70],u_xpb_out[81][70],u_xpb_out[82][70],u_xpb_out[83][70],u_xpb_out[84][70],u_xpb_out[85][70],u_xpb_out[86][70],u_xpb_out[87][70],u_xpb_out[88][70],u_xpb_out[89][70],u_xpb_out[90][70],u_xpb_out[91][70],u_xpb_out[92][70],u_xpb_out[93][70],u_xpb_out[94][70],u_xpb_out[95][70],u_xpb_out[96][70],u_xpb_out[97][70],u_xpb_out[98][70],u_xpb_out[99][70],u_xpb_out[100][70],u_xpb_out[101][70],u_xpb_out[102][70],u_xpb_out[103][70],u_xpb_out[104][70],u_xpb_out[105][70]};

assign col_out_71 = {u_xpb_out[0][71],u_xpb_out[1][71],u_xpb_out[2][71],u_xpb_out[3][71],u_xpb_out[4][71],u_xpb_out[5][71],u_xpb_out[6][71],u_xpb_out[7][71],u_xpb_out[8][71],u_xpb_out[9][71],u_xpb_out[10][71],u_xpb_out[11][71],u_xpb_out[12][71],u_xpb_out[13][71],u_xpb_out[14][71],u_xpb_out[15][71],u_xpb_out[16][71],u_xpb_out[17][71],u_xpb_out[18][71],u_xpb_out[19][71],u_xpb_out[20][71],u_xpb_out[21][71],u_xpb_out[22][71],u_xpb_out[23][71],u_xpb_out[24][71],u_xpb_out[25][71],u_xpb_out[26][71],u_xpb_out[27][71],u_xpb_out[28][71],u_xpb_out[29][71],u_xpb_out[30][71],u_xpb_out[31][71],u_xpb_out[32][71],u_xpb_out[33][71],u_xpb_out[34][71],u_xpb_out[35][71],u_xpb_out[36][71],u_xpb_out[37][71],u_xpb_out[38][71],u_xpb_out[39][71],u_xpb_out[40][71],u_xpb_out[41][71],u_xpb_out[42][71],u_xpb_out[43][71],u_xpb_out[44][71],u_xpb_out[45][71],u_xpb_out[46][71],u_xpb_out[47][71],u_xpb_out[48][71],u_xpb_out[49][71],u_xpb_out[50][71],u_xpb_out[51][71],u_xpb_out[52][71],u_xpb_out[53][71],u_xpb_out[54][71],u_xpb_out[55][71],u_xpb_out[56][71],u_xpb_out[57][71],u_xpb_out[58][71],u_xpb_out[59][71],u_xpb_out[60][71],u_xpb_out[61][71],u_xpb_out[62][71],u_xpb_out[63][71],u_xpb_out[64][71],u_xpb_out[65][71],u_xpb_out[66][71],u_xpb_out[67][71],u_xpb_out[68][71],u_xpb_out[69][71],u_xpb_out[70][71],u_xpb_out[71][71],u_xpb_out[72][71],u_xpb_out[73][71],u_xpb_out[74][71],u_xpb_out[75][71],u_xpb_out[76][71],u_xpb_out[77][71],u_xpb_out[78][71],u_xpb_out[79][71],u_xpb_out[80][71],u_xpb_out[81][71],u_xpb_out[82][71],u_xpb_out[83][71],u_xpb_out[84][71],u_xpb_out[85][71],u_xpb_out[86][71],u_xpb_out[87][71],u_xpb_out[88][71],u_xpb_out[89][71],u_xpb_out[90][71],u_xpb_out[91][71],u_xpb_out[92][71],u_xpb_out[93][71],u_xpb_out[94][71],u_xpb_out[95][71],u_xpb_out[96][71],u_xpb_out[97][71],u_xpb_out[98][71],u_xpb_out[99][71],u_xpb_out[100][71],u_xpb_out[101][71],u_xpb_out[102][71],u_xpb_out[103][71],u_xpb_out[104][71],u_xpb_out[105][71]};

assign col_out_72 = {u_xpb_out[0][72],u_xpb_out[1][72],u_xpb_out[2][72],u_xpb_out[3][72],u_xpb_out[4][72],u_xpb_out[5][72],u_xpb_out[6][72],u_xpb_out[7][72],u_xpb_out[8][72],u_xpb_out[9][72],u_xpb_out[10][72],u_xpb_out[11][72],u_xpb_out[12][72],u_xpb_out[13][72],u_xpb_out[14][72],u_xpb_out[15][72],u_xpb_out[16][72],u_xpb_out[17][72],u_xpb_out[18][72],u_xpb_out[19][72],u_xpb_out[20][72],u_xpb_out[21][72],u_xpb_out[22][72],u_xpb_out[23][72],u_xpb_out[24][72],u_xpb_out[25][72],u_xpb_out[26][72],u_xpb_out[27][72],u_xpb_out[28][72],u_xpb_out[29][72],u_xpb_out[30][72],u_xpb_out[31][72],u_xpb_out[32][72],u_xpb_out[33][72],u_xpb_out[34][72],u_xpb_out[35][72],u_xpb_out[36][72],u_xpb_out[37][72],u_xpb_out[38][72],u_xpb_out[39][72],u_xpb_out[40][72],u_xpb_out[41][72],u_xpb_out[42][72],u_xpb_out[43][72],u_xpb_out[44][72],u_xpb_out[45][72],u_xpb_out[46][72],u_xpb_out[47][72],u_xpb_out[48][72],u_xpb_out[49][72],u_xpb_out[50][72],u_xpb_out[51][72],u_xpb_out[52][72],u_xpb_out[53][72],u_xpb_out[54][72],u_xpb_out[55][72],u_xpb_out[56][72],u_xpb_out[57][72],u_xpb_out[58][72],u_xpb_out[59][72],u_xpb_out[60][72],u_xpb_out[61][72],u_xpb_out[62][72],u_xpb_out[63][72],u_xpb_out[64][72],u_xpb_out[65][72],u_xpb_out[66][72],u_xpb_out[67][72],u_xpb_out[68][72],u_xpb_out[69][72],u_xpb_out[70][72],u_xpb_out[71][72],u_xpb_out[72][72],u_xpb_out[73][72],u_xpb_out[74][72],u_xpb_out[75][72],u_xpb_out[76][72],u_xpb_out[77][72],u_xpb_out[78][72],u_xpb_out[79][72],u_xpb_out[80][72],u_xpb_out[81][72],u_xpb_out[82][72],u_xpb_out[83][72],u_xpb_out[84][72],u_xpb_out[85][72],u_xpb_out[86][72],u_xpb_out[87][72],u_xpb_out[88][72],u_xpb_out[89][72],u_xpb_out[90][72],u_xpb_out[91][72],u_xpb_out[92][72],u_xpb_out[93][72],u_xpb_out[94][72],u_xpb_out[95][72],u_xpb_out[96][72],u_xpb_out[97][72],u_xpb_out[98][72],u_xpb_out[99][72],u_xpb_out[100][72],u_xpb_out[101][72],u_xpb_out[102][72],u_xpb_out[103][72],u_xpb_out[104][72],u_xpb_out[105][72]};

assign col_out_73 = {u_xpb_out[0][73],u_xpb_out[1][73],u_xpb_out[2][73],u_xpb_out[3][73],u_xpb_out[4][73],u_xpb_out[5][73],u_xpb_out[6][73],u_xpb_out[7][73],u_xpb_out[8][73],u_xpb_out[9][73],u_xpb_out[10][73],u_xpb_out[11][73],u_xpb_out[12][73],u_xpb_out[13][73],u_xpb_out[14][73],u_xpb_out[15][73],u_xpb_out[16][73],u_xpb_out[17][73],u_xpb_out[18][73],u_xpb_out[19][73],u_xpb_out[20][73],u_xpb_out[21][73],u_xpb_out[22][73],u_xpb_out[23][73],u_xpb_out[24][73],u_xpb_out[25][73],u_xpb_out[26][73],u_xpb_out[27][73],u_xpb_out[28][73],u_xpb_out[29][73],u_xpb_out[30][73],u_xpb_out[31][73],u_xpb_out[32][73],u_xpb_out[33][73],u_xpb_out[34][73],u_xpb_out[35][73],u_xpb_out[36][73],u_xpb_out[37][73],u_xpb_out[38][73],u_xpb_out[39][73],u_xpb_out[40][73],u_xpb_out[41][73],u_xpb_out[42][73],u_xpb_out[43][73],u_xpb_out[44][73],u_xpb_out[45][73],u_xpb_out[46][73],u_xpb_out[47][73],u_xpb_out[48][73],u_xpb_out[49][73],u_xpb_out[50][73],u_xpb_out[51][73],u_xpb_out[52][73],u_xpb_out[53][73],u_xpb_out[54][73],u_xpb_out[55][73],u_xpb_out[56][73],u_xpb_out[57][73],u_xpb_out[58][73],u_xpb_out[59][73],u_xpb_out[60][73],u_xpb_out[61][73],u_xpb_out[62][73],u_xpb_out[63][73],u_xpb_out[64][73],u_xpb_out[65][73],u_xpb_out[66][73],u_xpb_out[67][73],u_xpb_out[68][73],u_xpb_out[69][73],u_xpb_out[70][73],u_xpb_out[71][73],u_xpb_out[72][73],u_xpb_out[73][73],u_xpb_out[74][73],u_xpb_out[75][73],u_xpb_out[76][73],u_xpb_out[77][73],u_xpb_out[78][73],u_xpb_out[79][73],u_xpb_out[80][73],u_xpb_out[81][73],u_xpb_out[82][73],u_xpb_out[83][73],u_xpb_out[84][73],u_xpb_out[85][73],u_xpb_out[86][73],u_xpb_out[87][73],u_xpb_out[88][73],u_xpb_out[89][73],u_xpb_out[90][73],u_xpb_out[91][73],u_xpb_out[92][73],u_xpb_out[93][73],u_xpb_out[94][73],u_xpb_out[95][73],u_xpb_out[96][73],u_xpb_out[97][73],u_xpb_out[98][73],u_xpb_out[99][73],u_xpb_out[100][73],u_xpb_out[101][73],u_xpb_out[102][73],u_xpb_out[103][73],u_xpb_out[104][73],u_xpb_out[105][73]};

assign col_out_74 = {u_xpb_out[0][74],u_xpb_out[1][74],u_xpb_out[2][74],u_xpb_out[3][74],u_xpb_out[4][74],u_xpb_out[5][74],u_xpb_out[6][74],u_xpb_out[7][74],u_xpb_out[8][74],u_xpb_out[9][74],u_xpb_out[10][74],u_xpb_out[11][74],u_xpb_out[12][74],u_xpb_out[13][74],u_xpb_out[14][74],u_xpb_out[15][74],u_xpb_out[16][74],u_xpb_out[17][74],u_xpb_out[18][74],u_xpb_out[19][74],u_xpb_out[20][74],u_xpb_out[21][74],u_xpb_out[22][74],u_xpb_out[23][74],u_xpb_out[24][74],u_xpb_out[25][74],u_xpb_out[26][74],u_xpb_out[27][74],u_xpb_out[28][74],u_xpb_out[29][74],u_xpb_out[30][74],u_xpb_out[31][74],u_xpb_out[32][74],u_xpb_out[33][74],u_xpb_out[34][74],u_xpb_out[35][74],u_xpb_out[36][74],u_xpb_out[37][74],u_xpb_out[38][74],u_xpb_out[39][74],u_xpb_out[40][74],u_xpb_out[41][74],u_xpb_out[42][74],u_xpb_out[43][74],u_xpb_out[44][74],u_xpb_out[45][74],u_xpb_out[46][74],u_xpb_out[47][74],u_xpb_out[48][74],u_xpb_out[49][74],u_xpb_out[50][74],u_xpb_out[51][74],u_xpb_out[52][74],u_xpb_out[53][74],u_xpb_out[54][74],u_xpb_out[55][74],u_xpb_out[56][74],u_xpb_out[57][74],u_xpb_out[58][74],u_xpb_out[59][74],u_xpb_out[60][74],u_xpb_out[61][74],u_xpb_out[62][74],u_xpb_out[63][74],u_xpb_out[64][74],u_xpb_out[65][74],u_xpb_out[66][74],u_xpb_out[67][74],u_xpb_out[68][74],u_xpb_out[69][74],u_xpb_out[70][74],u_xpb_out[71][74],u_xpb_out[72][74],u_xpb_out[73][74],u_xpb_out[74][74],u_xpb_out[75][74],u_xpb_out[76][74],u_xpb_out[77][74],u_xpb_out[78][74],u_xpb_out[79][74],u_xpb_out[80][74],u_xpb_out[81][74],u_xpb_out[82][74],u_xpb_out[83][74],u_xpb_out[84][74],u_xpb_out[85][74],u_xpb_out[86][74],u_xpb_out[87][74],u_xpb_out[88][74],u_xpb_out[89][74],u_xpb_out[90][74],u_xpb_out[91][74],u_xpb_out[92][74],u_xpb_out[93][74],u_xpb_out[94][74],u_xpb_out[95][74],u_xpb_out[96][74],u_xpb_out[97][74],u_xpb_out[98][74],u_xpb_out[99][74],u_xpb_out[100][74],u_xpb_out[101][74],u_xpb_out[102][74],u_xpb_out[103][74],u_xpb_out[104][74],u_xpb_out[105][74]};

assign col_out_75 = {u_xpb_out[0][75],u_xpb_out[1][75],u_xpb_out[2][75],u_xpb_out[3][75],u_xpb_out[4][75],u_xpb_out[5][75],u_xpb_out[6][75],u_xpb_out[7][75],u_xpb_out[8][75],u_xpb_out[9][75],u_xpb_out[10][75],u_xpb_out[11][75],u_xpb_out[12][75],u_xpb_out[13][75],u_xpb_out[14][75],u_xpb_out[15][75],u_xpb_out[16][75],u_xpb_out[17][75],u_xpb_out[18][75],u_xpb_out[19][75],u_xpb_out[20][75],u_xpb_out[21][75],u_xpb_out[22][75],u_xpb_out[23][75],u_xpb_out[24][75],u_xpb_out[25][75],u_xpb_out[26][75],u_xpb_out[27][75],u_xpb_out[28][75],u_xpb_out[29][75],u_xpb_out[30][75],u_xpb_out[31][75],u_xpb_out[32][75],u_xpb_out[33][75],u_xpb_out[34][75],u_xpb_out[35][75],u_xpb_out[36][75],u_xpb_out[37][75],u_xpb_out[38][75],u_xpb_out[39][75],u_xpb_out[40][75],u_xpb_out[41][75],u_xpb_out[42][75],u_xpb_out[43][75],u_xpb_out[44][75],u_xpb_out[45][75],u_xpb_out[46][75],u_xpb_out[47][75],u_xpb_out[48][75],u_xpb_out[49][75],u_xpb_out[50][75],u_xpb_out[51][75],u_xpb_out[52][75],u_xpb_out[53][75],u_xpb_out[54][75],u_xpb_out[55][75],u_xpb_out[56][75],u_xpb_out[57][75],u_xpb_out[58][75],u_xpb_out[59][75],u_xpb_out[60][75],u_xpb_out[61][75],u_xpb_out[62][75],u_xpb_out[63][75],u_xpb_out[64][75],u_xpb_out[65][75],u_xpb_out[66][75],u_xpb_out[67][75],u_xpb_out[68][75],u_xpb_out[69][75],u_xpb_out[70][75],u_xpb_out[71][75],u_xpb_out[72][75],u_xpb_out[73][75],u_xpb_out[74][75],u_xpb_out[75][75],u_xpb_out[76][75],u_xpb_out[77][75],u_xpb_out[78][75],u_xpb_out[79][75],u_xpb_out[80][75],u_xpb_out[81][75],u_xpb_out[82][75],u_xpb_out[83][75],u_xpb_out[84][75],u_xpb_out[85][75],u_xpb_out[86][75],u_xpb_out[87][75],u_xpb_out[88][75],u_xpb_out[89][75],u_xpb_out[90][75],u_xpb_out[91][75],u_xpb_out[92][75],u_xpb_out[93][75],u_xpb_out[94][75],u_xpb_out[95][75],u_xpb_out[96][75],u_xpb_out[97][75],u_xpb_out[98][75],u_xpb_out[99][75],u_xpb_out[100][75],u_xpb_out[101][75],u_xpb_out[102][75],u_xpb_out[103][75],u_xpb_out[104][75],u_xpb_out[105][75]};

assign col_out_76 = {u_xpb_out[0][76],u_xpb_out[1][76],u_xpb_out[2][76],u_xpb_out[3][76],u_xpb_out[4][76],u_xpb_out[5][76],u_xpb_out[6][76],u_xpb_out[7][76],u_xpb_out[8][76],u_xpb_out[9][76],u_xpb_out[10][76],u_xpb_out[11][76],u_xpb_out[12][76],u_xpb_out[13][76],u_xpb_out[14][76],u_xpb_out[15][76],u_xpb_out[16][76],u_xpb_out[17][76],u_xpb_out[18][76],u_xpb_out[19][76],u_xpb_out[20][76],u_xpb_out[21][76],u_xpb_out[22][76],u_xpb_out[23][76],u_xpb_out[24][76],u_xpb_out[25][76],u_xpb_out[26][76],u_xpb_out[27][76],u_xpb_out[28][76],u_xpb_out[29][76],u_xpb_out[30][76],u_xpb_out[31][76],u_xpb_out[32][76],u_xpb_out[33][76],u_xpb_out[34][76],u_xpb_out[35][76],u_xpb_out[36][76],u_xpb_out[37][76],u_xpb_out[38][76],u_xpb_out[39][76],u_xpb_out[40][76],u_xpb_out[41][76],u_xpb_out[42][76],u_xpb_out[43][76],u_xpb_out[44][76],u_xpb_out[45][76],u_xpb_out[46][76],u_xpb_out[47][76],u_xpb_out[48][76],u_xpb_out[49][76],u_xpb_out[50][76],u_xpb_out[51][76],u_xpb_out[52][76],u_xpb_out[53][76],u_xpb_out[54][76],u_xpb_out[55][76],u_xpb_out[56][76],u_xpb_out[57][76],u_xpb_out[58][76],u_xpb_out[59][76],u_xpb_out[60][76],u_xpb_out[61][76],u_xpb_out[62][76],u_xpb_out[63][76],u_xpb_out[64][76],u_xpb_out[65][76],u_xpb_out[66][76],u_xpb_out[67][76],u_xpb_out[68][76],u_xpb_out[69][76],u_xpb_out[70][76],u_xpb_out[71][76],u_xpb_out[72][76],u_xpb_out[73][76],u_xpb_out[74][76],u_xpb_out[75][76],u_xpb_out[76][76],u_xpb_out[77][76],u_xpb_out[78][76],u_xpb_out[79][76],u_xpb_out[80][76],u_xpb_out[81][76],u_xpb_out[82][76],u_xpb_out[83][76],u_xpb_out[84][76],u_xpb_out[85][76],u_xpb_out[86][76],u_xpb_out[87][76],u_xpb_out[88][76],u_xpb_out[89][76],u_xpb_out[90][76],u_xpb_out[91][76],u_xpb_out[92][76],u_xpb_out[93][76],u_xpb_out[94][76],u_xpb_out[95][76],u_xpb_out[96][76],u_xpb_out[97][76],u_xpb_out[98][76],u_xpb_out[99][76],u_xpb_out[100][76],u_xpb_out[101][76],u_xpb_out[102][76],u_xpb_out[103][76],u_xpb_out[104][76],u_xpb_out[105][76]};

assign col_out_77 = {u_xpb_out[0][77],u_xpb_out[1][77],u_xpb_out[2][77],u_xpb_out[3][77],u_xpb_out[4][77],u_xpb_out[5][77],u_xpb_out[6][77],u_xpb_out[7][77],u_xpb_out[8][77],u_xpb_out[9][77],u_xpb_out[10][77],u_xpb_out[11][77],u_xpb_out[12][77],u_xpb_out[13][77],u_xpb_out[14][77],u_xpb_out[15][77],u_xpb_out[16][77],u_xpb_out[17][77],u_xpb_out[18][77],u_xpb_out[19][77],u_xpb_out[20][77],u_xpb_out[21][77],u_xpb_out[22][77],u_xpb_out[23][77],u_xpb_out[24][77],u_xpb_out[25][77],u_xpb_out[26][77],u_xpb_out[27][77],u_xpb_out[28][77],u_xpb_out[29][77],u_xpb_out[30][77],u_xpb_out[31][77],u_xpb_out[32][77],u_xpb_out[33][77],u_xpb_out[34][77],u_xpb_out[35][77],u_xpb_out[36][77],u_xpb_out[37][77],u_xpb_out[38][77],u_xpb_out[39][77],u_xpb_out[40][77],u_xpb_out[41][77],u_xpb_out[42][77],u_xpb_out[43][77],u_xpb_out[44][77],u_xpb_out[45][77],u_xpb_out[46][77],u_xpb_out[47][77],u_xpb_out[48][77],u_xpb_out[49][77],u_xpb_out[50][77],u_xpb_out[51][77],u_xpb_out[52][77],u_xpb_out[53][77],u_xpb_out[54][77],u_xpb_out[55][77],u_xpb_out[56][77],u_xpb_out[57][77],u_xpb_out[58][77],u_xpb_out[59][77],u_xpb_out[60][77],u_xpb_out[61][77],u_xpb_out[62][77],u_xpb_out[63][77],u_xpb_out[64][77],u_xpb_out[65][77],u_xpb_out[66][77],u_xpb_out[67][77],u_xpb_out[68][77],u_xpb_out[69][77],u_xpb_out[70][77],u_xpb_out[71][77],u_xpb_out[72][77],u_xpb_out[73][77],u_xpb_out[74][77],u_xpb_out[75][77],u_xpb_out[76][77],u_xpb_out[77][77],u_xpb_out[78][77],u_xpb_out[79][77],u_xpb_out[80][77],u_xpb_out[81][77],u_xpb_out[82][77],u_xpb_out[83][77],u_xpb_out[84][77],u_xpb_out[85][77],u_xpb_out[86][77],u_xpb_out[87][77],u_xpb_out[88][77],u_xpb_out[89][77],u_xpb_out[90][77],u_xpb_out[91][77],u_xpb_out[92][77],u_xpb_out[93][77],u_xpb_out[94][77],u_xpb_out[95][77],u_xpb_out[96][77],u_xpb_out[97][77],u_xpb_out[98][77],u_xpb_out[99][77],u_xpb_out[100][77],u_xpb_out[101][77],u_xpb_out[102][77],u_xpb_out[103][77],u_xpb_out[104][77],u_xpb_out[105][77]};

assign col_out_78 = {u_xpb_out[0][78],u_xpb_out[1][78],u_xpb_out[2][78],u_xpb_out[3][78],u_xpb_out[4][78],u_xpb_out[5][78],u_xpb_out[6][78],u_xpb_out[7][78],u_xpb_out[8][78],u_xpb_out[9][78],u_xpb_out[10][78],u_xpb_out[11][78],u_xpb_out[12][78],u_xpb_out[13][78],u_xpb_out[14][78],u_xpb_out[15][78],u_xpb_out[16][78],u_xpb_out[17][78],u_xpb_out[18][78],u_xpb_out[19][78],u_xpb_out[20][78],u_xpb_out[21][78],u_xpb_out[22][78],u_xpb_out[23][78],u_xpb_out[24][78],u_xpb_out[25][78],u_xpb_out[26][78],u_xpb_out[27][78],u_xpb_out[28][78],u_xpb_out[29][78],u_xpb_out[30][78],u_xpb_out[31][78],u_xpb_out[32][78],u_xpb_out[33][78],u_xpb_out[34][78],u_xpb_out[35][78],u_xpb_out[36][78],u_xpb_out[37][78],u_xpb_out[38][78],u_xpb_out[39][78],u_xpb_out[40][78],u_xpb_out[41][78],u_xpb_out[42][78],u_xpb_out[43][78],u_xpb_out[44][78],u_xpb_out[45][78],u_xpb_out[46][78],u_xpb_out[47][78],u_xpb_out[48][78],u_xpb_out[49][78],u_xpb_out[50][78],u_xpb_out[51][78],u_xpb_out[52][78],u_xpb_out[53][78],u_xpb_out[54][78],u_xpb_out[55][78],u_xpb_out[56][78],u_xpb_out[57][78],u_xpb_out[58][78],u_xpb_out[59][78],u_xpb_out[60][78],u_xpb_out[61][78],u_xpb_out[62][78],u_xpb_out[63][78],u_xpb_out[64][78],u_xpb_out[65][78],u_xpb_out[66][78],u_xpb_out[67][78],u_xpb_out[68][78],u_xpb_out[69][78],u_xpb_out[70][78],u_xpb_out[71][78],u_xpb_out[72][78],u_xpb_out[73][78],u_xpb_out[74][78],u_xpb_out[75][78],u_xpb_out[76][78],u_xpb_out[77][78],u_xpb_out[78][78],u_xpb_out[79][78],u_xpb_out[80][78],u_xpb_out[81][78],u_xpb_out[82][78],u_xpb_out[83][78],u_xpb_out[84][78],u_xpb_out[85][78],u_xpb_out[86][78],u_xpb_out[87][78],u_xpb_out[88][78],u_xpb_out[89][78],u_xpb_out[90][78],u_xpb_out[91][78],u_xpb_out[92][78],u_xpb_out[93][78],u_xpb_out[94][78],u_xpb_out[95][78],u_xpb_out[96][78],u_xpb_out[97][78],u_xpb_out[98][78],u_xpb_out[99][78],u_xpb_out[100][78],u_xpb_out[101][78],u_xpb_out[102][78],u_xpb_out[103][78],u_xpb_out[104][78],u_xpb_out[105][78]};

assign col_out_79 = {u_xpb_out[0][79],u_xpb_out[1][79],u_xpb_out[2][79],u_xpb_out[3][79],u_xpb_out[4][79],u_xpb_out[5][79],u_xpb_out[6][79],u_xpb_out[7][79],u_xpb_out[8][79],u_xpb_out[9][79],u_xpb_out[10][79],u_xpb_out[11][79],u_xpb_out[12][79],u_xpb_out[13][79],u_xpb_out[14][79],u_xpb_out[15][79],u_xpb_out[16][79],u_xpb_out[17][79],u_xpb_out[18][79],u_xpb_out[19][79],u_xpb_out[20][79],u_xpb_out[21][79],u_xpb_out[22][79],u_xpb_out[23][79],u_xpb_out[24][79],u_xpb_out[25][79],u_xpb_out[26][79],u_xpb_out[27][79],u_xpb_out[28][79],u_xpb_out[29][79],u_xpb_out[30][79],u_xpb_out[31][79],u_xpb_out[32][79],u_xpb_out[33][79],u_xpb_out[34][79],u_xpb_out[35][79],u_xpb_out[36][79],u_xpb_out[37][79],u_xpb_out[38][79],u_xpb_out[39][79],u_xpb_out[40][79],u_xpb_out[41][79],u_xpb_out[42][79],u_xpb_out[43][79],u_xpb_out[44][79],u_xpb_out[45][79],u_xpb_out[46][79],u_xpb_out[47][79],u_xpb_out[48][79],u_xpb_out[49][79],u_xpb_out[50][79],u_xpb_out[51][79],u_xpb_out[52][79],u_xpb_out[53][79],u_xpb_out[54][79],u_xpb_out[55][79],u_xpb_out[56][79],u_xpb_out[57][79],u_xpb_out[58][79],u_xpb_out[59][79],u_xpb_out[60][79],u_xpb_out[61][79],u_xpb_out[62][79],u_xpb_out[63][79],u_xpb_out[64][79],u_xpb_out[65][79],u_xpb_out[66][79],u_xpb_out[67][79],u_xpb_out[68][79],u_xpb_out[69][79],u_xpb_out[70][79],u_xpb_out[71][79],u_xpb_out[72][79],u_xpb_out[73][79],u_xpb_out[74][79],u_xpb_out[75][79],u_xpb_out[76][79],u_xpb_out[77][79],u_xpb_out[78][79],u_xpb_out[79][79],u_xpb_out[80][79],u_xpb_out[81][79],u_xpb_out[82][79],u_xpb_out[83][79],u_xpb_out[84][79],u_xpb_out[85][79],u_xpb_out[86][79],u_xpb_out[87][79],u_xpb_out[88][79],u_xpb_out[89][79],u_xpb_out[90][79],u_xpb_out[91][79],u_xpb_out[92][79],u_xpb_out[93][79],u_xpb_out[94][79],u_xpb_out[95][79],u_xpb_out[96][79],u_xpb_out[97][79],u_xpb_out[98][79],u_xpb_out[99][79],u_xpb_out[100][79],u_xpb_out[101][79],u_xpb_out[102][79],u_xpb_out[103][79],u_xpb_out[104][79],u_xpb_out[105][79]};

assign col_out_80 = {u_xpb_out[0][80],u_xpb_out[1][80],u_xpb_out[2][80],u_xpb_out[3][80],u_xpb_out[4][80],u_xpb_out[5][80],u_xpb_out[6][80],u_xpb_out[7][80],u_xpb_out[8][80],u_xpb_out[9][80],u_xpb_out[10][80],u_xpb_out[11][80],u_xpb_out[12][80],u_xpb_out[13][80],u_xpb_out[14][80],u_xpb_out[15][80],u_xpb_out[16][80],u_xpb_out[17][80],u_xpb_out[18][80],u_xpb_out[19][80],u_xpb_out[20][80],u_xpb_out[21][80],u_xpb_out[22][80],u_xpb_out[23][80],u_xpb_out[24][80],u_xpb_out[25][80],u_xpb_out[26][80],u_xpb_out[27][80],u_xpb_out[28][80],u_xpb_out[29][80],u_xpb_out[30][80],u_xpb_out[31][80],u_xpb_out[32][80],u_xpb_out[33][80],u_xpb_out[34][80],u_xpb_out[35][80],u_xpb_out[36][80],u_xpb_out[37][80],u_xpb_out[38][80],u_xpb_out[39][80],u_xpb_out[40][80],u_xpb_out[41][80],u_xpb_out[42][80],u_xpb_out[43][80],u_xpb_out[44][80],u_xpb_out[45][80],u_xpb_out[46][80],u_xpb_out[47][80],u_xpb_out[48][80],u_xpb_out[49][80],u_xpb_out[50][80],u_xpb_out[51][80],u_xpb_out[52][80],u_xpb_out[53][80],u_xpb_out[54][80],u_xpb_out[55][80],u_xpb_out[56][80],u_xpb_out[57][80],u_xpb_out[58][80],u_xpb_out[59][80],u_xpb_out[60][80],u_xpb_out[61][80],u_xpb_out[62][80],u_xpb_out[63][80],u_xpb_out[64][80],u_xpb_out[65][80],u_xpb_out[66][80],u_xpb_out[67][80],u_xpb_out[68][80],u_xpb_out[69][80],u_xpb_out[70][80],u_xpb_out[71][80],u_xpb_out[72][80],u_xpb_out[73][80],u_xpb_out[74][80],u_xpb_out[75][80],u_xpb_out[76][80],u_xpb_out[77][80],u_xpb_out[78][80],u_xpb_out[79][80],u_xpb_out[80][80],u_xpb_out[81][80],u_xpb_out[82][80],u_xpb_out[83][80],u_xpb_out[84][80],u_xpb_out[85][80],u_xpb_out[86][80],u_xpb_out[87][80],u_xpb_out[88][80],u_xpb_out[89][80],u_xpb_out[90][80],u_xpb_out[91][80],u_xpb_out[92][80],u_xpb_out[93][80],u_xpb_out[94][80],u_xpb_out[95][80],u_xpb_out[96][80],u_xpb_out[97][80],u_xpb_out[98][80],u_xpb_out[99][80],u_xpb_out[100][80],u_xpb_out[101][80],u_xpb_out[102][80],u_xpb_out[103][80],u_xpb_out[104][80],u_xpb_out[105][80]};

assign col_out_81 = {u_xpb_out[0][81],u_xpb_out[1][81],u_xpb_out[2][81],u_xpb_out[3][81],u_xpb_out[4][81],u_xpb_out[5][81],u_xpb_out[6][81],u_xpb_out[7][81],u_xpb_out[8][81],u_xpb_out[9][81],u_xpb_out[10][81],u_xpb_out[11][81],u_xpb_out[12][81],u_xpb_out[13][81],u_xpb_out[14][81],u_xpb_out[15][81],u_xpb_out[16][81],u_xpb_out[17][81],u_xpb_out[18][81],u_xpb_out[19][81],u_xpb_out[20][81],u_xpb_out[21][81],u_xpb_out[22][81],u_xpb_out[23][81],u_xpb_out[24][81],u_xpb_out[25][81],u_xpb_out[26][81],u_xpb_out[27][81],u_xpb_out[28][81],u_xpb_out[29][81],u_xpb_out[30][81],u_xpb_out[31][81],u_xpb_out[32][81],u_xpb_out[33][81],u_xpb_out[34][81],u_xpb_out[35][81],u_xpb_out[36][81],u_xpb_out[37][81],u_xpb_out[38][81],u_xpb_out[39][81],u_xpb_out[40][81],u_xpb_out[41][81],u_xpb_out[42][81],u_xpb_out[43][81],u_xpb_out[44][81],u_xpb_out[45][81],u_xpb_out[46][81],u_xpb_out[47][81],u_xpb_out[48][81],u_xpb_out[49][81],u_xpb_out[50][81],u_xpb_out[51][81],u_xpb_out[52][81],u_xpb_out[53][81],u_xpb_out[54][81],u_xpb_out[55][81],u_xpb_out[56][81],u_xpb_out[57][81],u_xpb_out[58][81],u_xpb_out[59][81],u_xpb_out[60][81],u_xpb_out[61][81],u_xpb_out[62][81],u_xpb_out[63][81],u_xpb_out[64][81],u_xpb_out[65][81],u_xpb_out[66][81],u_xpb_out[67][81],u_xpb_out[68][81],u_xpb_out[69][81],u_xpb_out[70][81],u_xpb_out[71][81],u_xpb_out[72][81],u_xpb_out[73][81],u_xpb_out[74][81],u_xpb_out[75][81],u_xpb_out[76][81],u_xpb_out[77][81],u_xpb_out[78][81],u_xpb_out[79][81],u_xpb_out[80][81],u_xpb_out[81][81],u_xpb_out[82][81],u_xpb_out[83][81],u_xpb_out[84][81],u_xpb_out[85][81],u_xpb_out[86][81],u_xpb_out[87][81],u_xpb_out[88][81],u_xpb_out[89][81],u_xpb_out[90][81],u_xpb_out[91][81],u_xpb_out[92][81],u_xpb_out[93][81],u_xpb_out[94][81],u_xpb_out[95][81],u_xpb_out[96][81],u_xpb_out[97][81],u_xpb_out[98][81],u_xpb_out[99][81],u_xpb_out[100][81],u_xpb_out[101][81],u_xpb_out[102][81],u_xpb_out[103][81],u_xpb_out[104][81],u_xpb_out[105][81]};

assign col_out_82 = {u_xpb_out[0][82],u_xpb_out[1][82],u_xpb_out[2][82],u_xpb_out[3][82],u_xpb_out[4][82],u_xpb_out[5][82],u_xpb_out[6][82],u_xpb_out[7][82],u_xpb_out[8][82],u_xpb_out[9][82],u_xpb_out[10][82],u_xpb_out[11][82],u_xpb_out[12][82],u_xpb_out[13][82],u_xpb_out[14][82],u_xpb_out[15][82],u_xpb_out[16][82],u_xpb_out[17][82],u_xpb_out[18][82],u_xpb_out[19][82],u_xpb_out[20][82],u_xpb_out[21][82],u_xpb_out[22][82],u_xpb_out[23][82],u_xpb_out[24][82],u_xpb_out[25][82],u_xpb_out[26][82],u_xpb_out[27][82],u_xpb_out[28][82],u_xpb_out[29][82],u_xpb_out[30][82],u_xpb_out[31][82],u_xpb_out[32][82],u_xpb_out[33][82],u_xpb_out[34][82],u_xpb_out[35][82],u_xpb_out[36][82],u_xpb_out[37][82],u_xpb_out[38][82],u_xpb_out[39][82],u_xpb_out[40][82],u_xpb_out[41][82],u_xpb_out[42][82],u_xpb_out[43][82],u_xpb_out[44][82],u_xpb_out[45][82],u_xpb_out[46][82],u_xpb_out[47][82],u_xpb_out[48][82],u_xpb_out[49][82],u_xpb_out[50][82],u_xpb_out[51][82],u_xpb_out[52][82],u_xpb_out[53][82],u_xpb_out[54][82],u_xpb_out[55][82],u_xpb_out[56][82],u_xpb_out[57][82],u_xpb_out[58][82],u_xpb_out[59][82],u_xpb_out[60][82],u_xpb_out[61][82],u_xpb_out[62][82],u_xpb_out[63][82],u_xpb_out[64][82],u_xpb_out[65][82],u_xpb_out[66][82],u_xpb_out[67][82],u_xpb_out[68][82],u_xpb_out[69][82],u_xpb_out[70][82],u_xpb_out[71][82],u_xpb_out[72][82],u_xpb_out[73][82],u_xpb_out[74][82],u_xpb_out[75][82],u_xpb_out[76][82],u_xpb_out[77][82],u_xpb_out[78][82],u_xpb_out[79][82],u_xpb_out[80][82],u_xpb_out[81][82],u_xpb_out[82][82],u_xpb_out[83][82],u_xpb_out[84][82],u_xpb_out[85][82],u_xpb_out[86][82],u_xpb_out[87][82],u_xpb_out[88][82],u_xpb_out[89][82],u_xpb_out[90][82],u_xpb_out[91][82],u_xpb_out[92][82],u_xpb_out[93][82],u_xpb_out[94][82],u_xpb_out[95][82],u_xpb_out[96][82],u_xpb_out[97][82],u_xpb_out[98][82],u_xpb_out[99][82],u_xpb_out[100][82],u_xpb_out[101][82],u_xpb_out[102][82],u_xpb_out[103][82],u_xpb_out[104][82],u_xpb_out[105][82]};

assign col_out_83 = {u_xpb_out[0][83],u_xpb_out[1][83],u_xpb_out[2][83],u_xpb_out[3][83],u_xpb_out[4][83],u_xpb_out[5][83],u_xpb_out[6][83],u_xpb_out[7][83],u_xpb_out[8][83],u_xpb_out[9][83],u_xpb_out[10][83],u_xpb_out[11][83],u_xpb_out[12][83],u_xpb_out[13][83],u_xpb_out[14][83],u_xpb_out[15][83],u_xpb_out[16][83],u_xpb_out[17][83],u_xpb_out[18][83],u_xpb_out[19][83],u_xpb_out[20][83],u_xpb_out[21][83],u_xpb_out[22][83],u_xpb_out[23][83],u_xpb_out[24][83],u_xpb_out[25][83],u_xpb_out[26][83],u_xpb_out[27][83],u_xpb_out[28][83],u_xpb_out[29][83],u_xpb_out[30][83],u_xpb_out[31][83],u_xpb_out[32][83],u_xpb_out[33][83],u_xpb_out[34][83],u_xpb_out[35][83],u_xpb_out[36][83],u_xpb_out[37][83],u_xpb_out[38][83],u_xpb_out[39][83],u_xpb_out[40][83],u_xpb_out[41][83],u_xpb_out[42][83],u_xpb_out[43][83],u_xpb_out[44][83],u_xpb_out[45][83],u_xpb_out[46][83],u_xpb_out[47][83],u_xpb_out[48][83],u_xpb_out[49][83],u_xpb_out[50][83],u_xpb_out[51][83],u_xpb_out[52][83],u_xpb_out[53][83],u_xpb_out[54][83],u_xpb_out[55][83],u_xpb_out[56][83],u_xpb_out[57][83],u_xpb_out[58][83],u_xpb_out[59][83],u_xpb_out[60][83],u_xpb_out[61][83],u_xpb_out[62][83],u_xpb_out[63][83],u_xpb_out[64][83],u_xpb_out[65][83],u_xpb_out[66][83],u_xpb_out[67][83],u_xpb_out[68][83],u_xpb_out[69][83],u_xpb_out[70][83],u_xpb_out[71][83],u_xpb_out[72][83],u_xpb_out[73][83],u_xpb_out[74][83],u_xpb_out[75][83],u_xpb_out[76][83],u_xpb_out[77][83],u_xpb_out[78][83],u_xpb_out[79][83],u_xpb_out[80][83],u_xpb_out[81][83],u_xpb_out[82][83],u_xpb_out[83][83],u_xpb_out[84][83],u_xpb_out[85][83],u_xpb_out[86][83],u_xpb_out[87][83],u_xpb_out[88][83],u_xpb_out[89][83],u_xpb_out[90][83],u_xpb_out[91][83],u_xpb_out[92][83],u_xpb_out[93][83],u_xpb_out[94][83],u_xpb_out[95][83],u_xpb_out[96][83],u_xpb_out[97][83],u_xpb_out[98][83],u_xpb_out[99][83],u_xpb_out[100][83],u_xpb_out[101][83],u_xpb_out[102][83],u_xpb_out[103][83],u_xpb_out[104][83],u_xpb_out[105][83]};

assign col_out_84 = {u_xpb_out[0][84],u_xpb_out[1][84],u_xpb_out[2][84],u_xpb_out[3][84],u_xpb_out[4][84],u_xpb_out[5][84],u_xpb_out[6][84],u_xpb_out[7][84],u_xpb_out[8][84],u_xpb_out[9][84],u_xpb_out[10][84],u_xpb_out[11][84],u_xpb_out[12][84],u_xpb_out[13][84],u_xpb_out[14][84],u_xpb_out[15][84],u_xpb_out[16][84],u_xpb_out[17][84],u_xpb_out[18][84],u_xpb_out[19][84],u_xpb_out[20][84],u_xpb_out[21][84],u_xpb_out[22][84],u_xpb_out[23][84],u_xpb_out[24][84],u_xpb_out[25][84],u_xpb_out[26][84],u_xpb_out[27][84],u_xpb_out[28][84],u_xpb_out[29][84],u_xpb_out[30][84],u_xpb_out[31][84],u_xpb_out[32][84],u_xpb_out[33][84],u_xpb_out[34][84],u_xpb_out[35][84],u_xpb_out[36][84],u_xpb_out[37][84],u_xpb_out[38][84],u_xpb_out[39][84],u_xpb_out[40][84],u_xpb_out[41][84],u_xpb_out[42][84],u_xpb_out[43][84],u_xpb_out[44][84],u_xpb_out[45][84],u_xpb_out[46][84],u_xpb_out[47][84],u_xpb_out[48][84],u_xpb_out[49][84],u_xpb_out[50][84],u_xpb_out[51][84],u_xpb_out[52][84],u_xpb_out[53][84],u_xpb_out[54][84],u_xpb_out[55][84],u_xpb_out[56][84],u_xpb_out[57][84],u_xpb_out[58][84],u_xpb_out[59][84],u_xpb_out[60][84],u_xpb_out[61][84],u_xpb_out[62][84],u_xpb_out[63][84],u_xpb_out[64][84],u_xpb_out[65][84],u_xpb_out[66][84],u_xpb_out[67][84],u_xpb_out[68][84],u_xpb_out[69][84],u_xpb_out[70][84],u_xpb_out[71][84],u_xpb_out[72][84],u_xpb_out[73][84],u_xpb_out[74][84],u_xpb_out[75][84],u_xpb_out[76][84],u_xpb_out[77][84],u_xpb_out[78][84],u_xpb_out[79][84],u_xpb_out[80][84],u_xpb_out[81][84],u_xpb_out[82][84],u_xpb_out[83][84],u_xpb_out[84][84],u_xpb_out[85][84],u_xpb_out[86][84],u_xpb_out[87][84],u_xpb_out[88][84],u_xpb_out[89][84],u_xpb_out[90][84],u_xpb_out[91][84],u_xpb_out[92][84],u_xpb_out[93][84],u_xpb_out[94][84],u_xpb_out[95][84],u_xpb_out[96][84],u_xpb_out[97][84],u_xpb_out[98][84],u_xpb_out[99][84],u_xpb_out[100][84],u_xpb_out[101][84],u_xpb_out[102][84],u_xpb_out[103][84],u_xpb_out[104][84],u_xpb_out[105][84]};

assign col_out_85 = {u_xpb_out[0][85],u_xpb_out[1][85],u_xpb_out[2][85],u_xpb_out[3][85],u_xpb_out[4][85],u_xpb_out[5][85],u_xpb_out[6][85],u_xpb_out[7][85],u_xpb_out[8][85],u_xpb_out[9][85],u_xpb_out[10][85],u_xpb_out[11][85],u_xpb_out[12][85],u_xpb_out[13][85],u_xpb_out[14][85],u_xpb_out[15][85],u_xpb_out[16][85],u_xpb_out[17][85],u_xpb_out[18][85],u_xpb_out[19][85],u_xpb_out[20][85],u_xpb_out[21][85],u_xpb_out[22][85],u_xpb_out[23][85],u_xpb_out[24][85],u_xpb_out[25][85],u_xpb_out[26][85],u_xpb_out[27][85],u_xpb_out[28][85],u_xpb_out[29][85],u_xpb_out[30][85],u_xpb_out[31][85],u_xpb_out[32][85],u_xpb_out[33][85],u_xpb_out[34][85],u_xpb_out[35][85],u_xpb_out[36][85],u_xpb_out[37][85],u_xpb_out[38][85],u_xpb_out[39][85],u_xpb_out[40][85],u_xpb_out[41][85],u_xpb_out[42][85],u_xpb_out[43][85],u_xpb_out[44][85],u_xpb_out[45][85],u_xpb_out[46][85],u_xpb_out[47][85],u_xpb_out[48][85],u_xpb_out[49][85],u_xpb_out[50][85],u_xpb_out[51][85],u_xpb_out[52][85],u_xpb_out[53][85],u_xpb_out[54][85],u_xpb_out[55][85],u_xpb_out[56][85],u_xpb_out[57][85],u_xpb_out[58][85],u_xpb_out[59][85],u_xpb_out[60][85],u_xpb_out[61][85],u_xpb_out[62][85],u_xpb_out[63][85],u_xpb_out[64][85],u_xpb_out[65][85],u_xpb_out[66][85],u_xpb_out[67][85],u_xpb_out[68][85],u_xpb_out[69][85],u_xpb_out[70][85],u_xpb_out[71][85],u_xpb_out[72][85],u_xpb_out[73][85],u_xpb_out[74][85],u_xpb_out[75][85],u_xpb_out[76][85],u_xpb_out[77][85],u_xpb_out[78][85],u_xpb_out[79][85],u_xpb_out[80][85],u_xpb_out[81][85],u_xpb_out[82][85],u_xpb_out[83][85],u_xpb_out[84][85],u_xpb_out[85][85],u_xpb_out[86][85],u_xpb_out[87][85],u_xpb_out[88][85],u_xpb_out[89][85],u_xpb_out[90][85],u_xpb_out[91][85],u_xpb_out[92][85],u_xpb_out[93][85],u_xpb_out[94][85],u_xpb_out[95][85],u_xpb_out[96][85],u_xpb_out[97][85],u_xpb_out[98][85],u_xpb_out[99][85],u_xpb_out[100][85],u_xpb_out[101][85],u_xpb_out[102][85],u_xpb_out[103][85],u_xpb_out[104][85],u_xpb_out[105][85]};

assign col_out_86 = {u_xpb_out[0][86],u_xpb_out[1][86],u_xpb_out[2][86],u_xpb_out[3][86],u_xpb_out[4][86],u_xpb_out[5][86],u_xpb_out[6][86],u_xpb_out[7][86],u_xpb_out[8][86],u_xpb_out[9][86],u_xpb_out[10][86],u_xpb_out[11][86],u_xpb_out[12][86],u_xpb_out[13][86],u_xpb_out[14][86],u_xpb_out[15][86],u_xpb_out[16][86],u_xpb_out[17][86],u_xpb_out[18][86],u_xpb_out[19][86],u_xpb_out[20][86],u_xpb_out[21][86],u_xpb_out[22][86],u_xpb_out[23][86],u_xpb_out[24][86],u_xpb_out[25][86],u_xpb_out[26][86],u_xpb_out[27][86],u_xpb_out[28][86],u_xpb_out[29][86],u_xpb_out[30][86],u_xpb_out[31][86],u_xpb_out[32][86],u_xpb_out[33][86],u_xpb_out[34][86],u_xpb_out[35][86],u_xpb_out[36][86],u_xpb_out[37][86],u_xpb_out[38][86],u_xpb_out[39][86],u_xpb_out[40][86],u_xpb_out[41][86],u_xpb_out[42][86],u_xpb_out[43][86],u_xpb_out[44][86],u_xpb_out[45][86],u_xpb_out[46][86],u_xpb_out[47][86],u_xpb_out[48][86],u_xpb_out[49][86],u_xpb_out[50][86],u_xpb_out[51][86],u_xpb_out[52][86],u_xpb_out[53][86],u_xpb_out[54][86],u_xpb_out[55][86],u_xpb_out[56][86],u_xpb_out[57][86],u_xpb_out[58][86],u_xpb_out[59][86],u_xpb_out[60][86],u_xpb_out[61][86],u_xpb_out[62][86],u_xpb_out[63][86],u_xpb_out[64][86],u_xpb_out[65][86],u_xpb_out[66][86],u_xpb_out[67][86],u_xpb_out[68][86],u_xpb_out[69][86],u_xpb_out[70][86],u_xpb_out[71][86],u_xpb_out[72][86],u_xpb_out[73][86],u_xpb_out[74][86],u_xpb_out[75][86],u_xpb_out[76][86],u_xpb_out[77][86],u_xpb_out[78][86],u_xpb_out[79][86],u_xpb_out[80][86],u_xpb_out[81][86],u_xpb_out[82][86],u_xpb_out[83][86],u_xpb_out[84][86],u_xpb_out[85][86],u_xpb_out[86][86],u_xpb_out[87][86],u_xpb_out[88][86],u_xpb_out[89][86],u_xpb_out[90][86],u_xpb_out[91][86],u_xpb_out[92][86],u_xpb_out[93][86],u_xpb_out[94][86],u_xpb_out[95][86],u_xpb_out[96][86],u_xpb_out[97][86],u_xpb_out[98][86],u_xpb_out[99][86],u_xpb_out[100][86],u_xpb_out[101][86],u_xpb_out[102][86],u_xpb_out[103][86],u_xpb_out[104][86],u_xpb_out[105][86]};

assign col_out_87 = {u_xpb_out[0][87],u_xpb_out[1][87],u_xpb_out[2][87],u_xpb_out[3][87],u_xpb_out[4][87],u_xpb_out[5][87],u_xpb_out[6][87],u_xpb_out[7][87],u_xpb_out[8][87],u_xpb_out[9][87],u_xpb_out[10][87],u_xpb_out[11][87],u_xpb_out[12][87],u_xpb_out[13][87],u_xpb_out[14][87],u_xpb_out[15][87],u_xpb_out[16][87],u_xpb_out[17][87],u_xpb_out[18][87],u_xpb_out[19][87],u_xpb_out[20][87],u_xpb_out[21][87],u_xpb_out[22][87],u_xpb_out[23][87],u_xpb_out[24][87],u_xpb_out[25][87],u_xpb_out[26][87],u_xpb_out[27][87],u_xpb_out[28][87],u_xpb_out[29][87],u_xpb_out[30][87],u_xpb_out[31][87],u_xpb_out[32][87],u_xpb_out[33][87],u_xpb_out[34][87],u_xpb_out[35][87],u_xpb_out[36][87],u_xpb_out[37][87],u_xpb_out[38][87],u_xpb_out[39][87],u_xpb_out[40][87],u_xpb_out[41][87],u_xpb_out[42][87],u_xpb_out[43][87],u_xpb_out[44][87],u_xpb_out[45][87],u_xpb_out[46][87],u_xpb_out[47][87],u_xpb_out[48][87],u_xpb_out[49][87],u_xpb_out[50][87],u_xpb_out[51][87],u_xpb_out[52][87],u_xpb_out[53][87],u_xpb_out[54][87],u_xpb_out[55][87],u_xpb_out[56][87],u_xpb_out[57][87],u_xpb_out[58][87],u_xpb_out[59][87],u_xpb_out[60][87],u_xpb_out[61][87],u_xpb_out[62][87],u_xpb_out[63][87],u_xpb_out[64][87],u_xpb_out[65][87],u_xpb_out[66][87],u_xpb_out[67][87],u_xpb_out[68][87],u_xpb_out[69][87],u_xpb_out[70][87],u_xpb_out[71][87],u_xpb_out[72][87],u_xpb_out[73][87],u_xpb_out[74][87],u_xpb_out[75][87],u_xpb_out[76][87],u_xpb_out[77][87],u_xpb_out[78][87],u_xpb_out[79][87],u_xpb_out[80][87],u_xpb_out[81][87],u_xpb_out[82][87],u_xpb_out[83][87],u_xpb_out[84][87],u_xpb_out[85][87],u_xpb_out[86][87],u_xpb_out[87][87],u_xpb_out[88][87],u_xpb_out[89][87],u_xpb_out[90][87],u_xpb_out[91][87],u_xpb_out[92][87],u_xpb_out[93][87],u_xpb_out[94][87],u_xpb_out[95][87],u_xpb_out[96][87],u_xpb_out[97][87],u_xpb_out[98][87],u_xpb_out[99][87],u_xpb_out[100][87],u_xpb_out[101][87],u_xpb_out[102][87],u_xpb_out[103][87],u_xpb_out[104][87],u_xpb_out[105][87]};

assign col_out_88 = {u_xpb_out[0][88],u_xpb_out[1][88],u_xpb_out[2][88],u_xpb_out[3][88],u_xpb_out[4][88],u_xpb_out[5][88],u_xpb_out[6][88],u_xpb_out[7][88],u_xpb_out[8][88],u_xpb_out[9][88],u_xpb_out[10][88],u_xpb_out[11][88],u_xpb_out[12][88],u_xpb_out[13][88],u_xpb_out[14][88],u_xpb_out[15][88],u_xpb_out[16][88],u_xpb_out[17][88],u_xpb_out[18][88],u_xpb_out[19][88],u_xpb_out[20][88],u_xpb_out[21][88],u_xpb_out[22][88],u_xpb_out[23][88],u_xpb_out[24][88],u_xpb_out[25][88],u_xpb_out[26][88],u_xpb_out[27][88],u_xpb_out[28][88],u_xpb_out[29][88],u_xpb_out[30][88],u_xpb_out[31][88],u_xpb_out[32][88],u_xpb_out[33][88],u_xpb_out[34][88],u_xpb_out[35][88],u_xpb_out[36][88],u_xpb_out[37][88],u_xpb_out[38][88],u_xpb_out[39][88],u_xpb_out[40][88],u_xpb_out[41][88],u_xpb_out[42][88],u_xpb_out[43][88],u_xpb_out[44][88],u_xpb_out[45][88],u_xpb_out[46][88],u_xpb_out[47][88],u_xpb_out[48][88],u_xpb_out[49][88],u_xpb_out[50][88],u_xpb_out[51][88],u_xpb_out[52][88],u_xpb_out[53][88],u_xpb_out[54][88],u_xpb_out[55][88],u_xpb_out[56][88],u_xpb_out[57][88],u_xpb_out[58][88],u_xpb_out[59][88],u_xpb_out[60][88],u_xpb_out[61][88],u_xpb_out[62][88],u_xpb_out[63][88],u_xpb_out[64][88],u_xpb_out[65][88],u_xpb_out[66][88],u_xpb_out[67][88],u_xpb_out[68][88],u_xpb_out[69][88],u_xpb_out[70][88],u_xpb_out[71][88],u_xpb_out[72][88],u_xpb_out[73][88],u_xpb_out[74][88],u_xpb_out[75][88],u_xpb_out[76][88],u_xpb_out[77][88],u_xpb_out[78][88],u_xpb_out[79][88],u_xpb_out[80][88],u_xpb_out[81][88],u_xpb_out[82][88],u_xpb_out[83][88],u_xpb_out[84][88],u_xpb_out[85][88],u_xpb_out[86][88],u_xpb_out[87][88],u_xpb_out[88][88],u_xpb_out[89][88],u_xpb_out[90][88],u_xpb_out[91][88],u_xpb_out[92][88],u_xpb_out[93][88],u_xpb_out[94][88],u_xpb_out[95][88],u_xpb_out[96][88],u_xpb_out[97][88],u_xpb_out[98][88],u_xpb_out[99][88],u_xpb_out[100][88],u_xpb_out[101][88],u_xpb_out[102][88],u_xpb_out[103][88],u_xpb_out[104][88],u_xpb_out[105][88]};

assign col_out_89 = {u_xpb_out[0][89],u_xpb_out[1][89],u_xpb_out[2][89],u_xpb_out[3][89],u_xpb_out[4][89],u_xpb_out[5][89],u_xpb_out[6][89],u_xpb_out[7][89],u_xpb_out[8][89],u_xpb_out[9][89],u_xpb_out[10][89],u_xpb_out[11][89],u_xpb_out[12][89],u_xpb_out[13][89],u_xpb_out[14][89],u_xpb_out[15][89],u_xpb_out[16][89],u_xpb_out[17][89],u_xpb_out[18][89],u_xpb_out[19][89],u_xpb_out[20][89],u_xpb_out[21][89],u_xpb_out[22][89],u_xpb_out[23][89],u_xpb_out[24][89],u_xpb_out[25][89],u_xpb_out[26][89],u_xpb_out[27][89],u_xpb_out[28][89],u_xpb_out[29][89],u_xpb_out[30][89],u_xpb_out[31][89],u_xpb_out[32][89],u_xpb_out[33][89],u_xpb_out[34][89],u_xpb_out[35][89],u_xpb_out[36][89],u_xpb_out[37][89],u_xpb_out[38][89],u_xpb_out[39][89],u_xpb_out[40][89],u_xpb_out[41][89],u_xpb_out[42][89],u_xpb_out[43][89],u_xpb_out[44][89],u_xpb_out[45][89],u_xpb_out[46][89],u_xpb_out[47][89],u_xpb_out[48][89],u_xpb_out[49][89],u_xpb_out[50][89],u_xpb_out[51][89],u_xpb_out[52][89],u_xpb_out[53][89],u_xpb_out[54][89],u_xpb_out[55][89],u_xpb_out[56][89],u_xpb_out[57][89],u_xpb_out[58][89],u_xpb_out[59][89],u_xpb_out[60][89],u_xpb_out[61][89],u_xpb_out[62][89],u_xpb_out[63][89],u_xpb_out[64][89],u_xpb_out[65][89],u_xpb_out[66][89],u_xpb_out[67][89],u_xpb_out[68][89],u_xpb_out[69][89],u_xpb_out[70][89],u_xpb_out[71][89],u_xpb_out[72][89],u_xpb_out[73][89],u_xpb_out[74][89],u_xpb_out[75][89],u_xpb_out[76][89],u_xpb_out[77][89],u_xpb_out[78][89],u_xpb_out[79][89],u_xpb_out[80][89],u_xpb_out[81][89],u_xpb_out[82][89],u_xpb_out[83][89],u_xpb_out[84][89],u_xpb_out[85][89],u_xpb_out[86][89],u_xpb_out[87][89],u_xpb_out[88][89],u_xpb_out[89][89],u_xpb_out[90][89],u_xpb_out[91][89],u_xpb_out[92][89],u_xpb_out[93][89],u_xpb_out[94][89],u_xpb_out[95][89],u_xpb_out[96][89],u_xpb_out[97][89],u_xpb_out[98][89],u_xpb_out[99][89],u_xpb_out[100][89],u_xpb_out[101][89],u_xpb_out[102][89],u_xpb_out[103][89],u_xpb_out[104][89],u_xpb_out[105][89]};

assign col_out_90 = {u_xpb_out[0][90],u_xpb_out[1][90],u_xpb_out[2][90],u_xpb_out[3][90],u_xpb_out[4][90],u_xpb_out[5][90],u_xpb_out[6][90],u_xpb_out[7][90],u_xpb_out[8][90],u_xpb_out[9][90],u_xpb_out[10][90],u_xpb_out[11][90],u_xpb_out[12][90],u_xpb_out[13][90],u_xpb_out[14][90],u_xpb_out[15][90],u_xpb_out[16][90],u_xpb_out[17][90],u_xpb_out[18][90],u_xpb_out[19][90],u_xpb_out[20][90],u_xpb_out[21][90],u_xpb_out[22][90],u_xpb_out[23][90],u_xpb_out[24][90],u_xpb_out[25][90],u_xpb_out[26][90],u_xpb_out[27][90],u_xpb_out[28][90],u_xpb_out[29][90],u_xpb_out[30][90],u_xpb_out[31][90],u_xpb_out[32][90],u_xpb_out[33][90],u_xpb_out[34][90],u_xpb_out[35][90],u_xpb_out[36][90],u_xpb_out[37][90],u_xpb_out[38][90],u_xpb_out[39][90],u_xpb_out[40][90],u_xpb_out[41][90],u_xpb_out[42][90],u_xpb_out[43][90],u_xpb_out[44][90],u_xpb_out[45][90],u_xpb_out[46][90],u_xpb_out[47][90],u_xpb_out[48][90],u_xpb_out[49][90],u_xpb_out[50][90],u_xpb_out[51][90],u_xpb_out[52][90],u_xpb_out[53][90],u_xpb_out[54][90],u_xpb_out[55][90],u_xpb_out[56][90],u_xpb_out[57][90],u_xpb_out[58][90],u_xpb_out[59][90],u_xpb_out[60][90],u_xpb_out[61][90],u_xpb_out[62][90],u_xpb_out[63][90],u_xpb_out[64][90],u_xpb_out[65][90],u_xpb_out[66][90],u_xpb_out[67][90],u_xpb_out[68][90],u_xpb_out[69][90],u_xpb_out[70][90],u_xpb_out[71][90],u_xpb_out[72][90],u_xpb_out[73][90],u_xpb_out[74][90],u_xpb_out[75][90],u_xpb_out[76][90],u_xpb_out[77][90],u_xpb_out[78][90],u_xpb_out[79][90],u_xpb_out[80][90],u_xpb_out[81][90],u_xpb_out[82][90],u_xpb_out[83][90],u_xpb_out[84][90],u_xpb_out[85][90],u_xpb_out[86][90],u_xpb_out[87][90],u_xpb_out[88][90],u_xpb_out[89][90],u_xpb_out[90][90],u_xpb_out[91][90],u_xpb_out[92][90],u_xpb_out[93][90],u_xpb_out[94][90],u_xpb_out[95][90],u_xpb_out[96][90],u_xpb_out[97][90],u_xpb_out[98][90],u_xpb_out[99][90],u_xpb_out[100][90],u_xpb_out[101][90],u_xpb_out[102][90],u_xpb_out[103][90],u_xpb_out[104][90],u_xpb_out[105][90]};

assign col_out_91 = {u_xpb_out[0][91],u_xpb_out[1][91],u_xpb_out[2][91],u_xpb_out[3][91],u_xpb_out[4][91],u_xpb_out[5][91],u_xpb_out[6][91],u_xpb_out[7][91],u_xpb_out[8][91],u_xpb_out[9][91],u_xpb_out[10][91],u_xpb_out[11][91],u_xpb_out[12][91],u_xpb_out[13][91],u_xpb_out[14][91],u_xpb_out[15][91],u_xpb_out[16][91],u_xpb_out[17][91],u_xpb_out[18][91],u_xpb_out[19][91],u_xpb_out[20][91],u_xpb_out[21][91],u_xpb_out[22][91],u_xpb_out[23][91],u_xpb_out[24][91],u_xpb_out[25][91],u_xpb_out[26][91],u_xpb_out[27][91],u_xpb_out[28][91],u_xpb_out[29][91],u_xpb_out[30][91],u_xpb_out[31][91],u_xpb_out[32][91],u_xpb_out[33][91],u_xpb_out[34][91],u_xpb_out[35][91],u_xpb_out[36][91],u_xpb_out[37][91],u_xpb_out[38][91],u_xpb_out[39][91],u_xpb_out[40][91],u_xpb_out[41][91],u_xpb_out[42][91],u_xpb_out[43][91],u_xpb_out[44][91],u_xpb_out[45][91],u_xpb_out[46][91],u_xpb_out[47][91],u_xpb_out[48][91],u_xpb_out[49][91],u_xpb_out[50][91],u_xpb_out[51][91],u_xpb_out[52][91],u_xpb_out[53][91],u_xpb_out[54][91],u_xpb_out[55][91],u_xpb_out[56][91],u_xpb_out[57][91],u_xpb_out[58][91],u_xpb_out[59][91],u_xpb_out[60][91],u_xpb_out[61][91],u_xpb_out[62][91],u_xpb_out[63][91],u_xpb_out[64][91],u_xpb_out[65][91],u_xpb_out[66][91],u_xpb_out[67][91],u_xpb_out[68][91],u_xpb_out[69][91],u_xpb_out[70][91],u_xpb_out[71][91],u_xpb_out[72][91],u_xpb_out[73][91],u_xpb_out[74][91],u_xpb_out[75][91],u_xpb_out[76][91],u_xpb_out[77][91],u_xpb_out[78][91],u_xpb_out[79][91],u_xpb_out[80][91],u_xpb_out[81][91],u_xpb_out[82][91],u_xpb_out[83][91],u_xpb_out[84][91],u_xpb_out[85][91],u_xpb_out[86][91],u_xpb_out[87][91],u_xpb_out[88][91],u_xpb_out[89][91],u_xpb_out[90][91],u_xpb_out[91][91],u_xpb_out[92][91],u_xpb_out[93][91],u_xpb_out[94][91],u_xpb_out[95][91],u_xpb_out[96][91],u_xpb_out[97][91],u_xpb_out[98][91],u_xpb_out[99][91],u_xpb_out[100][91],u_xpb_out[101][91],u_xpb_out[102][91],u_xpb_out[103][91],u_xpb_out[104][91],u_xpb_out[105][91]};

assign col_out_92 = {u_xpb_out[0][92],u_xpb_out[1][92],u_xpb_out[2][92],u_xpb_out[3][92],u_xpb_out[4][92],u_xpb_out[5][92],u_xpb_out[6][92],u_xpb_out[7][92],u_xpb_out[8][92],u_xpb_out[9][92],u_xpb_out[10][92],u_xpb_out[11][92],u_xpb_out[12][92],u_xpb_out[13][92],u_xpb_out[14][92],u_xpb_out[15][92],u_xpb_out[16][92],u_xpb_out[17][92],u_xpb_out[18][92],u_xpb_out[19][92],u_xpb_out[20][92],u_xpb_out[21][92],u_xpb_out[22][92],u_xpb_out[23][92],u_xpb_out[24][92],u_xpb_out[25][92],u_xpb_out[26][92],u_xpb_out[27][92],u_xpb_out[28][92],u_xpb_out[29][92],u_xpb_out[30][92],u_xpb_out[31][92],u_xpb_out[32][92],u_xpb_out[33][92],u_xpb_out[34][92],u_xpb_out[35][92],u_xpb_out[36][92],u_xpb_out[37][92],u_xpb_out[38][92],u_xpb_out[39][92],u_xpb_out[40][92],u_xpb_out[41][92],u_xpb_out[42][92],u_xpb_out[43][92],u_xpb_out[44][92],u_xpb_out[45][92],u_xpb_out[46][92],u_xpb_out[47][92],u_xpb_out[48][92],u_xpb_out[49][92],u_xpb_out[50][92],u_xpb_out[51][92],u_xpb_out[52][92],u_xpb_out[53][92],u_xpb_out[54][92],u_xpb_out[55][92],u_xpb_out[56][92],u_xpb_out[57][92],u_xpb_out[58][92],u_xpb_out[59][92],u_xpb_out[60][92],u_xpb_out[61][92],u_xpb_out[62][92],u_xpb_out[63][92],u_xpb_out[64][92],u_xpb_out[65][92],u_xpb_out[66][92],u_xpb_out[67][92],u_xpb_out[68][92],u_xpb_out[69][92],u_xpb_out[70][92],u_xpb_out[71][92],u_xpb_out[72][92],u_xpb_out[73][92],u_xpb_out[74][92],u_xpb_out[75][92],u_xpb_out[76][92],u_xpb_out[77][92],u_xpb_out[78][92],u_xpb_out[79][92],u_xpb_out[80][92],u_xpb_out[81][92],u_xpb_out[82][92],u_xpb_out[83][92],u_xpb_out[84][92],u_xpb_out[85][92],u_xpb_out[86][92],u_xpb_out[87][92],u_xpb_out[88][92],u_xpb_out[89][92],u_xpb_out[90][92],u_xpb_out[91][92],u_xpb_out[92][92],u_xpb_out[93][92],u_xpb_out[94][92],u_xpb_out[95][92],u_xpb_out[96][92],u_xpb_out[97][92],u_xpb_out[98][92],u_xpb_out[99][92],u_xpb_out[100][92],u_xpb_out[101][92],u_xpb_out[102][92],u_xpb_out[103][92],u_xpb_out[104][92],u_xpb_out[105][92]};

assign col_out_93 = {u_xpb_out[0][93],u_xpb_out[1][93],u_xpb_out[2][93],u_xpb_out[3][93],u_xpb_out[4][93],u_xpb_out[5][93],u_xpb_out[6][93],u_xpb_out[7][93],u_xpb_out[8][93],u_xpb_out[9][93],u_xpb_out[10][93],u_xpb_out[11][93],u_xpb_out[12][93],u_xpb_out[13][93],u_xpb_out[14][93],u_xpb_out[15][93],u_xpb_out[16][93],u_xpb_out[17][93],u_xpb_out[18][93],u_xpb_out[19][93],u_xpb_out[20][93],u_xpb_out[21][93],u_xpb_out[22][93],u_xpb_out[23][93],u_xpb_out[24][93],u_xpb_out[25][93],u_xpb_out[26][93],u_xpb_out[27][93],u_xpb_out[28][93],u_xpb_out[29][93],u_xpb_out[30][93],u_xpb_out[31][93],u_xpb_out[32][93],u_xpb_out[33][93],u_xpb_out[34][93],u_xpb_out[35][93],u_xpb_out[36][93],u_xpb_out[37][93],u_xpb_out[38][93],u_xpb_out[39][93],u_xpb_out[40][93],u_xpb_out[41][93],u_xpb_out[42][93],u_xpb_out[43][93],u_xpb_out[44][93],u_xpb_out[45][93],u_xpb_out[46][93],u_xpb_out[47][93],u_xpb_out[48][93],u_xpb_out[49][93],u_xpb_out[50][93],u_xpb_out[51][93],u_xpb_out[52][93],u_xpb_out[53][93],u_xpb_out[54][93],u_xpb_out[55][93],u_xpb_out[56][93],u_xpb_out[57][93],u_xpb_out[58][93],u_xpb_out[59][93],u_xpb_out[60][93],u_xpb_out[61][93],u_xpb_out[62][93],u_xpb_out[63][93],u_xpb_out[64][93],u_xpb_out[65][93],u_xpb_out[66][93],u_xpb_out[67][93],u_xpb_out[68][93],u_xpb_out[69][93],u_xpb_out[70][93],u_xpb_out[71][93],u_xpb_out[72][93],u_xpb_out[73][93],u_xpb_out[74][93],u_xpb_out[75][93],u_xpb_out[76][93],u_xpb_out[77][93],u_xpb_out[78][93],u_xpb_out[79][93],u_xpb_out[80][93],u_xpb_out[81][93],u_xpb_out[82][93],u_xpb_out[83][93],u_xpb_out[84][93],u_xpb_out[85][93],u_xpb_out[86][93],u_xpb_out[87][93],u_xpb_out[88][93],u_xpb_out[89][93],u_xpb_out[90][93],u_xpb_out[91][93],u_xpb_out[92][93],u_xpb_out[93][93],u_xpb_out[94][93],u_xpb_out[95][93],u_xpb_out[96][93],u_xpb_out[97][93],u_xpb_out[98][93],u_xpb_out[99][93],u_xpb_out[100][93],u_xpb_out[101][93],u_xpb_out[102][93],u_xpb_out[103][93],u_xpb_out[104][93],u_xpb_out[105][93]};

assign col_out_94 = {u_xpb_out[0][94],u_xpb_out[1][94],u_xpb_out[2][94],u_xpb_out[3][94],u_xpb_out[4][94],u_xpb_out[5][94],u_xpb_out[6][94],u_xpb_out[7][94],u_xpb_out[8][94],u_xpb_out[9][94],u_xpb_out[10][94],u_xpb_out[11][94],u_xpb_out[12][94],u_xpb_out[13][94],u_xpb_out[14][94],u_xpb_out[15][94],u_xpb_out[16][94],u_xpb_out[17][94],u_xpb_out[18][94],u_xpb_out[19][94],u_xpb_out[20][94],u_xpb_out[21][94],u_xpb_out[22][94],u_xpb_out[23][94],u_xpb_out[24][94],u_xpb_out[25][94],u_xpb_out[26][94],u_xpb_out[27][94],u_xpb_out[28][94],u_xpb_out[29][94],u_xpb_out[30][94],u_xpb_out[31][94],u_xpb_out[32][94],u_xpb_out[33][94],u_xpb_out[34][94],u_xpb_out[35][94],u_xpb_out[36][94],u_xpb_out[37][94],u_xpb_out[38][94],u_xpb_out[39][94],u_xpb_out[40][94],u_xpb_out[41][94],u_xpb_out[42][94],u_xpb_out[43][94],u_xpb_out[44][94],u_xpb_out[45][94],u_xpb_out[46][94],u_xpb_out[47][94],u_xpb_out[48][94],u_xpb_out[49][94],u_xpb_out[50][94],u_xpb_out[51][94],u_xpb_out[52][94],u_xpb_out[53][94],u_xpb_out[54][94],u_xpb_out[55][94],u_xpb_out[56][94],u_xpb_out[57][94],u_xpb_out[58][94],u_xpb_out[59][94],u_xpb_out[60][94],u_xpb_out[61][94],u_xpb_out[62][94],u_xpb_out[63][94],u_xpb_out[64][94],u_xpb_out[65][94],u_xpb_out[66][94],u_xpb_out[67][94],u_xpb_out[68][94],u_xpb_out[69][94],u_xpb_out[70][94],u_xpb_out[71][94],u_xpb_out[72][94],u_xpb_out[73][94],u_xpb_out[74][94],u_xpb_out[75][94],u_xpb_out[76][94],u_xpb_out[77][94],u_xpb_out[78][94],u_xpb_out[79][94],u_xpb_out[80][94],u_xpb_out[81][94],u_xpb_out[82][94],u_xpb_out[83][94],u_xpb_out[84][94],u_xpb_out[85][94],u_xpb_out[86][94],u_xpb_out[87][94],u_xpb_out[88][94],u_xpb_out[89][94],u_xpb_out[90][94],u_xpb_out[91][94],u_xpb_out[92][94],u_xpb_out[93][94],u_xpb_out[94][94],u_xpb_out[95][94],u_xpb_out[96][94],u_xpb_out[97][94],u_xpb_out[98][94],u_xpb_out[99][94],u_xpb_out[100][94],u_xpb_out[101][94],u_xpb_out[102][94],u_xpb_out[103][94],u_xpb_out[104][94],u_xpb_out[105][94]};

assign col_out_95 = {u_xpb_out[0][95],u_xpb_out[1][95],u_xpb_out[2][95],u_xpb_out[3][95],u_xpb_out[4][95],u_xpb_out[5][95],u_xpb_out[6][95],u_xpb_out[7][95],u_xpb_out[8][95],u_xpb_out[9][95],u_xpb_out[10][95],u_xpb_out[11][95],u_xpb_out[12][95],u_xpb_out[13][95],u_xpb_out[14][95],u_xpb_out[15][95],u_xpb_out[16][95],u_xpb_out[17][95],u_xpb_out[18][95],u_xpb_out[19][95],u_xpb_out[20][95],u_xpb_out[21][95],u_xpb_out[22][95],u_xpb_out[23][95],u_xpb_out[24][95],u_xpb_out[25][95],u_xpb_out[26][95],u_xpb_out[27][95],u_xpb_out[28][95],u_xpb_out[29][95],u_xpb_out[30][95],u_xpb_out[31][95],u_xpb_out[32][95],u_xpb_out[33][95],u_xpb_out[34][95],u_xpb_out[35][95],u_xpb_out[36][95],u_xpb_out[37][95],u_xpb_out[38][95],u_xpb_out[39][95],u_xpb_out[40][95],u_xpb_out[41][95],u_xpb_out[42][95],u_xpb_out[43][95],u_xpb_out[44][95],u_xpb_out[45][95],u_xpb_out[46][95],u_xpb_out[47][95],u_xpb_out[48][95],u_xpb_out[49][95],u_xpb_out[50][95],u_xpb_out[51][95],u_xpb_out[52][95],u_xpb_out[53][95],u_xpb_out[54][95],u_xpb_out[55][95],u_xpb_out[56][95],u_xpb_out[57][95],u_xpb_out[58][95],u_xpb_out[59][95],u_xpb_out[60][95],u_xpb_out[61][95],u_xpb_out[62][95],u_xpb_out[63][95],u_xpb_out[64][95],u_xpb_out[65][95],u_xpb_out[66][95],u_xpb_out[67][95],u_xpb_out[68][95],u_xpb_out[69][95],u_xpb_out[70][95],u_xpb_out[71][95],u_xpb_out[72][95],u_xpb_out[73][95],u_xpb_out[74][95],u_xpb_out[75][95],u_xpb_out[76][95],u_xpb_out[77][95],u_xpb_out[78][95],u_xpb_out[79][95],u_xpb_out[80][95],u_xpb_out[81][95],u_xpb_out[82][95],u_xpb_out[83][95],u_xpb_out[84][95],u_xpb_out[85][95],u_xpb_out[86][95],u_xpb_out[87][95],u_xpb_out[88][95],u_xpb_out[89][95],u_xpb_out[90][95],u_xpb_out[91][95],u_xpb_out[92][95],u_xpb_out[93][95],u_xpb_out[94][95],u_xpb_out[95][95],u_xpb_out[96][95],u_xpb_out[97][95],u_xpb_out[98][95],u_xpb_out[99][95],u_xpb_out[100][95],u_xpb_out[101][95],u_xpb_out[102][95],u_xpb_out[103][95],u_xpb_out[104][95],u_xpb_out[105][95]};

assign col_out_96 = {u_xpb_out[0][96],u_xpb_out[1][96],u_xpb_out[2][96],u_xpb_out[3][96],u_xpb_out[4][96],u_xpb_out[5][96],u_xpb_out[6][96],u_xpb_out[7][96],u_xpb_out[8][96],u_xpb_out[9][96],u_xpb_out[10][96],u_xpb_out[11][96],u_xpb_out[12][96],u_xpb_out[13][96],u_xpb_out[14][96],u_xpb_out[15][96],u_xpb_out[16][96],u_xpb_out[17][96],u_xpb_out[18][96],u_xpb_out[19][96],u_xpb_out[20][96],u_xpb_out[21][96],u_xpb_out[22][96],u_xpb_out[23][96],u_xpb_out[24][96],u_xpb_out[25][96],u_xpb_out[26][96],u_xpb_out[27][96],u_xpb_out[28][96],u_xpb_out[29][96],u_xpb_out[30][96],u_xpb_out[31][96],u_xpb_out[32][96],u_xpb_out[33][96],u_xpb_out[34][96],u_xpb_out[35][96],u_xpb_out[36][96],u_xpb_out[37][96],u_xpb_out[38][96],u_xpb_out[39][96],u_xpb_out[40][96],u_xpb_out[41][96],u_xpb_out[42][96],u_xpb_out[43][96],u_xpb_out[44][96],u_xpb_out[45][96],u_xpb_out[46][96],u_xpb_out[47][96],u_xpb_out[48][96],u_xpb_out[49][96],u_xpb_out[50][96],u_xpb_out[51][96],u_xpb_out[52][96],u_xpb_out[53][96],u_xpb_out[54][96],u_xpb_out[55][96],u_xpb_out[56][96],u_xpb_out[57][96],u_xpb_out[58][96],u_xpb_out[59][96],u_xpb_out[60][96],u_xpb_out[61][96],u_xpb_out[62][96],u_xpb_out[63][96],u_xpb_out[64][96],u_xpb_out[65][96],u_xpb_out[66][96],u_xpb_out[67][96],u_xpb_out[68][96],u_xpb_out[69][96],u_xpb_out[70][96],u_xpb_out[71][96],u_xpb_out[72][96],u_xpb_out[73][96],u_xpb_out[74][96],u_xpb_out[75][96],u_xpb_out[76][96],u_xpb_out[77][96],u_xpb_out[78][96],u_xpb_out[79][96],u_xpb_out[80][96],u_xpb_out[81][96],u_xpb_out[82][96],u_xpb_out[83][96],u_xpb_out[84][96],u_xpb_out[85][96],u_xpb_out[86][96],u_xpb_out[87][96],u_xpb_out[88][96],u_xpb_out[89][96],u_xpb_out[90][96],u_xpb_out[91][96],u_xpb_out[92][96],u_xpb_out[93][96],u_xpb_out[94][96],u_xpb_out[95][96],u_xpb_out[96][96],u_xpb_out[97][96],u_xpb_out[98][96],u_xpb_out[99][96],u_xpb_out[100][96],u_xpb_out[101][96],u_xpb_out[102][96],u_xpb_out[103][96],u_xpb_out[104][96],u_xpb_out[105][96]};

assign col_out_97 = {u_xpb_out[0][97],u_xpb_out[1][97],u_xpb_out[2][97],u_xpb_out[3][97],u_xpb_out[4][97],u_xpb_out[5][97],u_xpb_out[6][97],u_xpb_out[7][97],u_xpb_out[8][97],u_xpb_out[9][97],u_xpb_out[10][97],u_xpb_out[11][97],u_xpb_out[12][97],u_xpb_out[13][97],u_xpb_out[14][97],u_xpb_out[15][97],u_xpb_out[16][97],u_xpb_out[17][97],u_xpb_out[18][97],u_xpb_out[19][97],u_xpb_out[20][97],u_xpb_out[21][97],u_xpb_out[22][97],u_xpb_out[23][97],u_xpb_out[24][97],u_xpb_out[25][97],u_xpb_out[26][97],u_xpb_out[27][97],u_xpb_out[28][97],u_xpb_out[29][97],u_xpb_out[30][97],u_xpb_out[31][97],u_xpb_out[32][97],u_xpb_out[33][97],u_xpb_out[34][97],u_xpb_out[35][97],u_xpb_out[36][97],u_xpb_out[37][97],u_xpb_out[38][97],u_xpb_out[39][97],u_xpb_out[40][97],u_xpb_out[41][97],u_xpb_out[42][97],u_xpb_out[43][97],u_xpb_out[44][97],u_xpb_out[45][97],u_xpb_out[46][97],u_xpb_out[47][97],u_xpb_out[48][97],u_xpb_out[49][97],u_xpb_out[50][97],u_xpb_out[51][97],u_xpb_out[52][97],u_xpb_out[53][97],u_xpb_out[54][97],u_xpb_out[55][97],u_xpb_out[56][97],u_xpb_out[57][97],u_xpb_out[58][97],u_xpb_out[59][97],u_xpb_out[60][97],u_xpb_out[61][97],u_xpb_out[62][97],u_xpb_out[63][97],u_xpb_out[64][97],u_xpb_out[65][97],u_xpb_out[66][97],u_xpb_out[67][97],u_xpb_out[68][97],u_xpb_out[69][97],u_xpb_out[70][97],u_xpb_out[71][97],u_xpb_out[72][97],u_xpb_out[73][97],u_xpb_out[74][97],u_xpb_out[75][97],u_xpb_out[76][97],u_xpb_out[77][97],u_xpb_out[78][97],u_xpb_out[79][97],u_xpb_out[80][97],u_xpb_out[81][97],u_xpb_out[82][97],u_xpb_out[83][97],u_xpb_out[84][97],u_xpb_out[85][97],u_xpb_out[86][97],u_xpb_out[87][97],u_xpb_out[88][97],u_xpb_out[89][97],u_xpb_out[90][97],u_xpb_out[91][97],u_xpb_out[92][97],u_xpb_out[93][97],u_xpb_out[94][97],u_xpb_out[95][97],u_xpb_out[96][97],u_xpb_out[97][97],u_xpb_out[98][97],u_xpb_out[99][97],u_xpb_out[100][97],u_xpb_out[101][97],u_xpb_out[102][97],u_xpb_out[103][97],u_xpb_out[104][97],u_xpb_out[105][97]};

assign col_out_98 = {u_xpb_out[0][98],u_xpb_out[1][98],u_xpb_out[2][98],u_xpb_out[3][98],u_xpb_out[4][98],u_xpb_out[5][98],u_xpb_out[6][98],u_xpb_out[7][98],u_xpb_out[8][98],u_xpb_out[9][98],u_xpb_out[10][98],u_xpb_out[11][98],u_xpb_out[12][98],u_xpb_out[13][98],u_xpb_out[14][98],u_xpb_out[15][98],u_xpb_out[16][98],u_xpb_out[17][98],u_xpb_out[18][98],u_xpb_out[19][98],u_xpb_out[20][98],u_xpb_out[21][98],u_xpb_out[22][98],u_xpb_out[23][98],u_xpb_out[24][98],u_xpb_out[25][98],u_xpb_out[26][98],u_xpb_out[27][98],u_xpb_out[28][98],u_xpb_out[29][98],u_xpb_out[30][98],u_xpb_out[31][98],u_xpb_out[32][98],u_xpb_out[33][98],u_xpb_out[34][98],u_xpb_out[35][98],u_xpb_out[36][98],u_xpb_out[37][98],u_xpb_out[38][98],u_xpb_out[39][98],u_xpb_out[40][98],u_xpb_out[41][98],u_xpb_out[42][98],u_xpb_out[43][98],u_xpb_out[44][98],u_xpb_out[45][98],u_xpb_out[46][98],u_xpb_out[47][98],u_xpb_out[48][98],u_xpb_out[49][98],u_xpb_out[50][98],u_xpb_out[51][98],u_xpb_out[52][98],u_xpb_out[53][98],u_xpb_out[54][98],u_xpb_out[55][98],u_xpb_out[56][98],u_xpb_out[57][98],u_xpb_out[58][98],u_xpb_out[59][98],u_xpb_out[60][98],u_xpb_out[61][98],u_xpb_out[62][98],u_xpb_out[63][98],u_xpb_out[64][98],u_xpb_out[65][98],u_xpb_out[66][98],u_xpb_out[67][98],u_xpb_out[68][98],u_xpb_out[69][98],u_xpb_out[70][98],u_xpb_out[71][98],u_xpb_out[72][98],u_xpb_out[73][98],u_xpb_out[74][98],u_xpb_out[75][98],u_xpb_out[76][98],u_xpb_out[77][98],u_xpb_out[78][98],u_xpb_out[79][98],u_xpb_out[80][98],u_xpb_out[81][98],u_xpb_out[82][98],u_xpb_out[83][98],u_xpb_out[84][98],u_xpb_out[85][98],u_xpb_out[86][98],u_xpb_out[87][98],u_xpb_out[88][98],u_xpb_out[89][98],u_xpb_out[90][98],u_xpb_out[91][98],u_xpb_out[92][98],u_xpb_out[93][98],u_xpb_out[94][98],u_xpb_out[95][98],u_xpb_out[96][98],u_xpb_out[97][98],u_xpb_out[98][98],u_xpb_out[99][98],u_xpb_out[100][98],u_xpb_out[101][98],u_xpb_out[102][98],u_xpb_out[103][98],u_xpb_out[104][98],u_xpb_out[105][98]};

assign col_out_99 = {u_xpb_out[0][99],u_xpb_out[1][99],u_xpb_out[2][99],u_xpb_out[3][99],u_xpb_out[4][99],u_xpb_out[5][99],u_xpb_out[6][99],u_xpb_out[7][99],u_xpb_out[8][99],u_xpb_out[9][99],u_xpb_out[10][99],u_xpb_out[11][99],u_xpb_out[12][99],u_xpb_out[13][99],u_xpb_out[14][99],u_xpb_out[15][99],u_xpb_out[16][99],u_xpb_out[17][99],u_xpb_out[18][99],u_xpb_out[19][99],u_xpb_out[20][99],u_xpb_out[21][99],u_xpb_out[22][99],u_xpb_out[23][99],u_xpb_out[24][99],u_xpb_out[25][99],u_xpb_out[26][99],u_xpb_out[27][99],u_xpb_out[28][99],u_xpb_out[29][99],u_xpb_out[30][99],u_xpb_out[31][99],u_xpb_out[32][99],u_xpb_out[33][99],u_xpb_out[34][99],u_xpb_out[35][99],u_xpb_out[36][99],u_xpb_out[37][99],u_xpb_out[38][99],u_xpb_out[39][99],u_xpb_out[40][99],u_xpb_out[41][99],u_xpb_out[42][99],u_xpb_out[43][99],u_xpb_out[44][99],u_xpb_out[45][99],u_xpb_out[46][99],u_xpb_out[47][99],u_xpb_out[48][99],u_xpb_out[49][99],u_xpb_out[50][99],u_xpb_out[51][99],u_xpb_out[52][99],u_xpb_out[53][99],u_xpb_out[54][99],u_xpb_out[55][99],u_xpb_out[56][99],u_xpb_out[57][99],u_xpb_out[58][99],u_xpb_out[59][99],u_xpb_out[60][99],u_xpb_out[61][99],u_xpb_out[62][99],u_xpb_out[63][99],u_xpb_out[64][99],u_xpb_out[65][99],u_xpb_out[66][99],u_xpb_out[67][99],u_xpb_out[68][99],u_xpb_out[69][99],u_xpb_out[70][99],u_xpb_out[71][99],u_xpb_out[72][99],u_xpb_out[73][99],u_xpb_out[74][99],u_xpb_out[75][99],u_xpb_out[76][99],u_xpb_out[77][99],u_xpb_out[78][99],u_xpb_out[79][99],u_xpb_out[80][99],u_xpb_out[81][99],u_xpb_out[82][99],u_xpb_out[83][99],u_xpb_out[84][99],u_xpb_out[85][99],u_xpb_out[86][99],u_xpb_out[87][99],u_xpb_out[88][99],u_xpb_out[89][99],u_xpb_out[90][99],u_xpb_out[91][99],u_xpb_out[92][99],u_xpb_out[93][99],u_xpb_out[94][99],u_xpb_out[95][99],u_xpb_out[96][99],u_xpb_out[97][99],u_xpb_out[98][99],u_xpb_out[99][99],u_xpb_out[100][99],u_xpb_out[101][99],u_xpb_out[102][99],u_xpb_out[103][99],u_xpb_out[104][99],u_xpb_out[105][99]};

assign col_out_100 = {u_xpb_out[0][100],u_xpb_out[1][100],u_xpb_out[2][100],u_xpb_out[3][100],u_xpb_out[4][100],u_xpb_out[5][100],u_xpb_out[6][100],u_xpb_out[7][100],u_xpb_out[8][100],u_xpb_out[9][100],u_xpb_out[10][100],u_xpb_out[11][100],u_xpb_out[12][100],u_xpb_out[13][100],u_xpb_out[14][100],u_xpb_out[15][100],u_xpb_out[16][100],u_xpb_out[17][100],u_xpb_out[18][100],u_xpb_out[19][100],u_xpb_out[20][100],u_xpb_out[21][100],u_xpb_out[22][100],u_xpb_out[23][100],u_xpb_out[24][100],u_xpb_out[25][100],u_xpb_out[26][100],u_xpb_out[27][100],u_xpb_out[28][100],u_xpb_out[29][100],u_xpb_out[30][100],u_xpb_out[31][100],u_xpb_out[32][100],u_xpb_out[33][100],u_xpb_out[34][100],u_xpb_out[35][100],u_xpb_out[36][100],u_xpb_out[37][100],u_xpb_out[38][100],u_xpb_out[39][100],u_xpb_out[40][100],u_xpb_out[41][100],u_xpb_out[42][100],u_xpb_out[43][100],u_xpb_out[44][100],u_xpb_out[45][100],u_xpb_out[46][100],u_xpb_out[47][100],u_xpb_out[48][100],u_xpb_out[49][100],u_xpb_out[50][100],u_xpb_out[51][100],u_xpb_out[52][100],u_xpb_out[53][100],u_xpb_out[54][100],u_xpb_out[55][100],u_xpb_out[56][100],u_xpb_out[57][100],u_xpb_out[58][100],u_xpb_out[59][100],u_xpb_out[60][100],u_xpb_out[61][100],u_xpb_out[62][100],u_xpb_out[63][100],u_xpb_out[64][100],u_xpb_out[65][100],u_xpb_out[66][100],u_xpb_out[67][100],u_xpb_out[68][100],u_xpb_out[69][100],u_xpb_out[70][100],u_xpb_out[71][100],u_xpb_out[72][100],u_xpb_out[73][100],u_xpb_out[74][100],u_xpb_out[75][100],u_xpb_out[76][100],u_xpb_out[77][100],u_xpb_out[78][100],u_xpb_out[79][100],u_xpb_out[80][100],u_xpb_out[81][100],u_xpb_out[82][100],u_xpb_out[83][100],u_xpb_out[84][100],u_xpb_out[85][100],u_xpb_out[86][100],u_xpb_out[87][100],u_xpb_out[88][100],u_xpb_out[89][100],u_xpb_out[90][100],u_xpb_out[91][100],u_xpb_out[92][100],u_xpb_out[93][100],u_xpb_out[94][100],u_xpb_out[95][100],u_xpb_out[96][100],u_xpb_out[97][100],u_xpb_out[98][100],u_xpb_out[99][100],u_xpb_out[100][100],u_xpb_out[101][100],u_xpb_out[102][100],u_xpb_out[103][100],u_xpb_out[104][100],u_xpb_out[105][100]};

assign col_out_101 = {u_xpb_out[0][101],u_xpb_out[1][101],u_xpb_out[2][101],u_xpb_out[3][101],u_xpb_out[4][101],u_xpb_out[5][101],u_xpb_out[6][101],u_xpb_out[7][101],u_xpb_out[8][101],u_xpb_out[9][101],u_xpb_out[10][101],u_xpb_out[11][101],u_xpb_out[12][101],u_xpb_out[13][101],u_xpb_out[14][101],u_xpb_out[15][101],u_xpb_out[16][101],u_xpb_out[17][101],u_xpb_out[18][101],u_xpb_out[19][101],u_xpb_out[20][101],u_xpb_out[21][101],u_xpb_out[22][101],u_xpb_out[23][101],u_xpb_out[24][101],u_xpb_out[25][101],u_xpb_out[26][101],u_xpb_out[27][101],u_xpb_out[28][101],u_xpb_out[29][101],u_xpb_out[30][101],u_xpb_out[31][101],u_xpb_out[32][101],u_xpb_out[33][101],u_xpb_out[34][101],u_xpb_out[35][101],u_xpb_out[36][101],u_xpb_out[37][101],u_xpb_out[38][101],u_xpb_out[39][101],u_xpb_out[40][101],u_xpb_out[41][101],u_xpb_out[42][101],u_xpb_out[43][101],u_xpb_out[44][101],u_xpb_out[45][101],u_xpb_out[46][101],u_xpb_out[47][101],u_xpb_out[48][101],u_xpb_out[49][101],u_xpb_out[50][101],u_xpb_out[51][101],u_xpb_out[52][101],u_xpb_out[53][101],u_xpb_out[54][101],u_xpb_out[55][101],u_xpb_out[56][101],u_xpb_out[57][101],u_xpb_out[58][101],u_xpb_out[59][101],u_xpb_out[60][101],u_xpb_out[61][101],u_xpb_out[62][101],u_xpb_out[63][101],u_xpb_out[64][101],u_xpb_out[65][101],u_xpb_out[66][101],u_xpb_out[67][101],u_xpb_out[68][101],u_xpb_out[69][101],u_xpb_out[70][101],u_xpb_out[71][101],u_xpb_out[72][101],u_xpb_out[73][101],u_xpb_out[74][101],u_xpb_out[75][101],u_xpb_out[76][101],u_xpb_out[77][101],u_xpb_out[78][101],u_xpb_out[79][101],u_xpb_out[80][101],u_xpb_out[81][101],u_xpb_out[82][101],u_xpb_out[83][101],u_xpb_out[84][101],u_xpb_out[85][101],u_xpb_out[86][101],u_xpb_out[87][101],u_xpb_out[88][101],u_xpb_out[89][101],u_xpb_out[90][101],u_xpb_out[91][101],u_xpb_out[92][101],u_xpb_out[93][101],u_xpb_out[94][101],u_xpb_out[95][101],u_xpb_out[96][101],u_xpb_out[97][101],u_xpb_out[98][101],u_xpb_out[99][101],u_xpb_out[100][101],u_xpb_out[101][101],u_xpb_out[102][101],u_xpb_out[103][101],u_xpb_out[104][101],u_xpb_out[105][101]};

assign col_out_102 = {u_xpb_out[0][102],u_xpb_out[1][102],u_xpb_out[2][102],u_xpb_out[3][102],u_xpb_out[4][102],u_xpb_out[5][102],u_xpb_out[6][102],u_xpb_out[7][102],u_xpb_out[8][102],u_xpb_out[9][102],u_xpb_out[10][102],u_xpb_out[11][102],u_xpb_out[12][102],u_xpb_out[13][102],u_xpb_out[14][102],u_xpb_out[15][102],u_xpb_out[16][102],u_xpb_out[17][102],u_xpb_out[18][102],u_xpb_out[19][102],u_xpb_out[20][102],u_xpb_out[21][102],u_xpb_out[22][102],u_xpb_out[23][102],u_xpb_out[24][102],u_xpb_out[25][102],u_xpb_out[26][102],u_xpb_out[27][102],u_xpb_out[28][102],u_xpb_out[29][102],u_xpb_out[30][102],u_xpb_out[31][102],u_xpb_out[32][102],u_xpb_out[33][102],u_xpb_out[34][102],u_xpb_out[35][102],u_xpb_out[36][102],u_xpb_out[37][102],u_xpb_out[38][102],u_xpb_out[39][102],u_xpb_out[40][102],u_xpb_out[41][102],u_xpb_out[42][102],u_xpb_out[43][102],u_xpb_out[44][102],u_xpb_out[45][102],u_xpb_out[46][102],u_xpb_out[47][102],u_xpb_out[48][102],u_xpb_out[49][102],u_xpb_out[50][102],u_xpb_out[51][102],u_xpb_out[52][102],u_xpb_out[53][102],u_xpb_out[54][102],u_xpb_out[55][102],u_xpb_out[56][102],u_xpb_out[57][102],u_xpb_out[58][102],u_xpb_out[59][102],u_xpb_out[60][102],u_xpb_out[61][102],u_xpb_out[62][102],u_xpb_out[63][102],u_xpb_out[64][102],u_xpb_out[65][102],u_xpb_out[66][102],u_xpb_out[67][102],u_xpb_out[68][102],u_xpb_out[69][102],u_xpb_out[70][102],u_xpb_out[71][102],u_xpb_out[72][102],u_xpb_out[73][102],u_xpb_out[74][102],u_xpb_out[75][102],u_xpb_out[76][102],u_xpb_out[77][102],u_xpb_out[78][102],u_xpb_out[79][102],u_xpb_out[80][102],u_xpb_out[81][102],u_xpb_out[82][102],u_xpb_out[83][102],u_xpb_out[84][102],u_xpb_out[85][102],u_xpb_out[86][102],u_xpb_out[87][102],u_xpb_out[88][102],u_xpb_out[89][102],u_xpb_out[90][102],u_xpb_out[91][102],u_xpb_out[92][102],u_xpb_out[93][102],u_xpb_out[94][102],u_xpb_out[95][102],u_xpb_out[96][102],u_xpb_out[97][102],u_xpb_out[98][102],u_xpb_out[99][102],u_xpb_out[100][102],u_xpb_out[101][102],u_xpb_out[102][102],u_xpb_out[103][102],u_xpb_out[104][102],u_xpb_out[105][102]};

assign col_out_103 = {u_xpb_out[0][103],u_xpb_out[1][103],u_xpb_out[2][103],u_xpb_out[3][103],u_xpb_out[4][103],u_xpb_out[5][103],u_xpb_out[6][103],u_xpb_out[7][103],u_xpb_out[8][103],u_xpb_out[9][103],u_xpb_out[10][103],u_xpb_out[11][103],u_xpb_out[12][103],u_xpb_out[13][103],u_xpb_out[14][103],u_xpb_out[15][103],u_xpb_out[16][103],u_xpb_out[17][103],u_xpb_out[18][103],u_xpb_out[19][103],u_xpb_out[20][103],u_xpb_out[21][103],u_xpb_out[22][103],u_xpb_out[23][103],u_xpb_out[24][103],u_xpb_out[25][103],u_xpb_out[26][103],u_xpb_out[27][103],u_xpb_out[28][103],u_xpb_out[29][103],u_xpb_out[30][103],u_xpb_out[31][103],u_xpb_out[32][103],u_xpb_out[33][103],u_xpb_out[34][103],u_xpb_out[35][103],u_xpb_out[36][103],u_xpb_out[37][103],u_xpb_out[38][103],u_xpb_out[39][103],u_xpb_out[40][103],u_xpb_out[41][103],u_xpb_out[42][103],u_xpb_out[43][103],u_xpb_out[44][103],u_xpb_out[45][103],u_xpb_out[46][103],u_xpb_out[47][103],u_xpb_out[48][103],u_xpb_out[49][103],u_xpb_out[50][103],u_xpb_out[51][103],u_xpb_out[52][103],u_xpb_out[53][103],u_xpb_out[54][103],u_xpb_out[55][103],u_xpb_out[56][103],u_xpb_out[57][103],u_xpb_out[58][103],u_xpb_out[59][103],u_xpb_out[60][103],u_xpb_out[61][103],u_xpb_out[62][103],u_xpb_out[63][103],u_xpb_out[64][103],u_xpb_out[65][103],u_xpb_out[66][103],u_xpb_out[67][103],u_xpb_out[68][103],u_xpb_out[69][103],u_xpb_out[70][103],u_xpb_out[71][103],u_xpb_out[72][103],u_xpb_out[73][103],u_xpb_out[74][103],u_xpb_out[75][103],u_xpb_out[76][103],u_xpb_out[77][103],u_xpb_out[78][103],u_xpb_out[79][103],u_xpb_out[80][103],u_xpb_out[81][103],u_xpb_out[82][103],u_xpb_out[83][103],u_xpb_out[84][103],u_xpb_out[85][103],u_xpb_out[86][103],u_xpb_out[87][103],u_xpb_out[88][103],u_xpb_out[89][103],u_xpb_out[90][103],u_xpb_out[91][103],u_xpb_out[92][103],u_xpb_out[93][103],u_xpb_out[94][103],u_xpb_out[95][103],u_xpb_out[96][103],u_xpb_out[97][103],u_xpb_out[98][103],u_xpb_out[99][103],u_xpb_out[100][103],u_xpb_out[101][103],u_xpb_out[102][103],u_xpb_out[103][103],u_xpb_out[104][103],u_xpb_out[105][103]};

assign col_out_104 = {u_xpb_out[0][104],u_xpb_out[1][104],u_xpb_out[2][104],u_xpb_out[3][104],u_xpb_out[4][104],u_xpb_out[5][104],u_xpb_out[6][104],u_xpb_out[7][104],u_xpb_out[8][104],u_xpb_out[9][104],u_xpb_out[10][104],u_xpb_out[11][104],u_xpb_out[12][104],u_xpb_out[13][104],u_xpb_out[14][104],u_xpb_out[15][104],u_xpb_out[16][104],u_xpb_out[17][104],u_xpb_out[18][104],u_xpb_out[19][104],u_xpb_out[20][104],u_xpb_out[21][104],u_xpb_out[22][104],u_xpb_out[23][104],u_xpb_out[24][104],u_xpb_out[25][104],u_xpb_out[26][104],u_xpb_out[27][104],u_xpb_out[28][104],u_xpb_out[29][104],u_xpb_out[30][104],u_xpb_out[31][104],u_xpb_out[32][104],u_xpb_out[33][104],u_xpb_out[34][104],u_xpb_out[35][104],u_xpb_out[36][104],u_xpb_out[37][104],u_xpb_out[38][104],u_xpb_out[39][104],u_xpb_out[40][104],u_xpb_out[41][104],u_xpb_out[42][104],u_xpb_out[43][104],u_xpb_out[44][104],u_xpb_out[45][104],u_xpb_out[46][104],u_xpb_out[47][104],u_xpb_out[48][104],u_xpb_out[49][104],u_xpb_out[50][104],u_xpb_out[51][104],u_xpb_out[52][104],u_xpb_out[53][104],u_xpb_out[54][104],u_xpb_out[55][104],u_xpb_out[56][104],u_xpb_out[57][104],u_xpb_out[58][104],u_xpb_out[59][104],u_xpb_out[60][104],u_xpb_out[61][104],u_xpb_out[62][104],u_xpb_out[63][104],u_xpb_out[64][104],u_xpb_out[65][104],u_xpb_out[66][104],u_xpb_out[67][104],u_xpb_out[68][104],u_xpb_out[69][104],u_xpb_out[70][104],u_xpb_out[71][104],u_xpb_out[72][104],u_xpb_out[73][104],u_xpb_out[74][104],u_xpb_out[75][104],u_xpb_out[76][104],u_xpb_out[77][104],u_xpb_out[78][104],u_xpb_out[79][104],u_xpb_out[80][104],u_xpb_out[81][104],u_xpb_out[82][104],u_xpb_out[83][104],u_xpb_out[84][104],u_xpb_out[85][104],u_xpb_out[86][104],u_xpb_out[87][104],u_xpb_out[88][104],u_xpb_out[89][104],u_xpb_out[90][104],u_xpb_out[91][104],u_xpb_out[92][104],u_xpb_out[93][104],u_xpb_out[94][104],u_xpb_out[95][104],u_xpb_out[96][104],u_xpb_out[97][104],u_xpb_out[98][104],u_xpb_out[99][104],u_xpb_out[100][104],u_xpb_out[101][104],u_xpb_out[102][104],u_xpb_out[103][104],u_xpb_out[104][104],u_xpb_out[105][104]};

assign col_out_105 = {u_xpb_out[0][105],u_xpb_out[1][105],u_xpb_out[2][105],u_xpb_out[3][105],u_xpb_out[4][105],u_xpb_out[5][105],u_xpb_out[6][105],u_xpb_out[7][105],u_xpb_out[8][105],u_xpb_out[9][105],u_xpb_out[10][105],u_xpb_out[11][105],u_xpb_out[12][105],u_xpb_out[13][105],u_xpb_out[14][105],u_xpb_out[15][105],u_xpb_out[16][105],u_xpb_out[17][105],u_xpb_out[18][105],u_xpb_out[19][105],u_xpb_out[20][105],u_xpb_out[21][105],u_xpb_out[22][105],u_xpb_out[23][105],u_xpb_out[24][105],u_xpb_out[25][105],u_xpb_out[26][105],u_xpb_out[27][105],u_xpb_out[28][105],u_xpb_out[29][105],u_xpb_out[30][105],u_xpb_out[31][105],u_xpb_out[32][105],u_xpb_out[33][105],u_xpb_out[34][105],u_xpb_out[35][105],u_xpb_out[36][105],u_xpb_out[37][105],u_xpb_out[38][105],u_xpb_out[39][105],u_xpb_out[40][105],u_xpb_out[41][105],u_xpb_out[42][105],u_xpb_out[43][105],u_xpb_out[44][105],u_xpb_out[45][105],u_xpb_out[46][105],u_xpb_out[47][105],u_xpb_out[48][105],u_xpb_out[49][105],u_xpb_out[50][105],u_xpb_out[51][105],u_xpb_out[52][105],u_xpb_out[53][105],u_xpb_out[54][105],u_xpb_out[55][105],u_xpb_out[56][105],u_xpb_out[57][105],u_xpb_out[58][105],u_xpb_out[59][105],u_xpb_out[60][105],u_xpb_out[61][105],u_xpb_out[62][105],u_xpb_out[63][105],u_xpb_out[64][105],u_xpb_out[65][105],u_xpb_out[66][105],u_xpb_out[67][105],u_xpb_out[68][105],u_xpb_out[69][105],u_xpb_out[70][105],u_xpb_out[71][105],u_xpb_out[72][105],u_xpb_out[73][105],u_xpb_out[74][105],u_xpb_out[75][105],u_xpb_out[76][105],u_xpb_out[77][105],u_xpb_out[78][105],u_xpb_out[79][105],u_xpb_out[80][105],u_xpb_out[81][105],u_xpb_out[82][105],u_xpb_out[83][105],u_xpb_out[84][105],u_xpb_out[85][105],u_xpb_out[86][105],u_xpb_out[87][105],u_xpb_out[88][105],u_xpb_out[89][105],u_xpb_out[90][105],u_xpb_out[91][105],u_xpb_out[92][105],u_xpb_out[93][105],u_xpb_out[94][105],u_xpb_out[95][105],u_xpb_out[96][105],u_xpb_out[97][105],u_xpb_out[98][105],u_xpb_out[99][105],u_xpb_out[100][105],u_xpb_out[101][105],u_xpb_out[102][105],u_xpb_out[103][105],u_xpb_out[104][105],u_xpb_out[105][105]};

assign col_out_106 = {u_xpb_out[0][106],u_xpb_out[1][106],u_xpb_out[2][106],u_xpb_out[3][106],u_xpb_out[4][106],u_xpb_out[5][106],u_xpb_out[6][106],u_xpb_out[7][106],u_xpb_out[8][106],u_xpb_out[9][106],u_xpb_out[10][106],u_xpb_out[11][106],u_xpb_out[12][106],u_xpb_out[13][106],u_xpb_out[14][106],u_xpb_out[15][106],u_xpb_out[16][106],u_xpb_out[17][106],u_xpb_out[18][106],u_xpb_out[19][106],u_xpb_out[20][106],u_xpb_out[21][106],u_xpb_out[22][106],u_xpb_out[23][106],u_xpb_out[24][106],u_xpb_out[25][106],u_xpb_out[26][106],u_xpb_out[27][106],u_xpb_out[28][106],u_xpb_out[29][106],u_xpb_out[30][106],u_xpb_out[31][106],u_xpb_out[32][106],u_xpb_out[33][106],u_xpb_out[34][106],u_xpb_out[35][106],u_xpb_out[36][106],u_xpb_out[37][106],u_xpb_out[38][106],u_xpb_out[39][106],u_xpb_out[40][106],u_xpb_out[41][106],u_xpb_out[42][106],u_xpb_out[43][106],u_xpb_out[44][106],u_xpb_out[45][106],u_xpb_out[46][106],u_xpb_out[47][106],u_xpb_out[48][106],u_xpb_out[49][106],u_xpb_out[50][106],u_xpb_out[51][106],u_xpb_out[52][106],u_xpb_out[53][106],u_xpb_out[54][106],u_xpb_out[55][106],u_xpb_out[56][106],u_xpb_out[57][106],u_xpb_out[58][106],u_xpb_out[59][106],u_xpb_out[60][106],u_xpb_out[61][106],u_xpb_out[62][106],u_xpb_out[63][106],u_xpb_out[64][106],u_xpb_out[65][106],u_xpb_out[66][106],u_xpb_out[67][106],u_xpb_out[68][106],u_xpb_out[69][106],u_xpb_out[70][106],u_xpb_out[71][106],u_xpb_out[72][106],u_xpb_out[73][106],u_xpb_out[74][106],u_xpb_out[75][106],u_xpb_out[76][106],u_xpb_out[77][106],u_xpb_out[78][106],u_xpb_out[79][106],u_xpb_out[80][106],u_xpb_out[81][106],u_xpb_out[82][106],u_xpb_out[83][106],u_xpb_out[84][106],u_xpb_out[85][106],u_xpb_out[86][106],u_xpb_out[87][106],u_xpb_out[88][106],u_xpb_out[89][106],u_xpb_out[90][106],u_xpb_out[91][106],u_xpb_out[92][106],u_xpb_out[93][106],u_xpb_out[94][106],u_xpb_out[95][106],u_xpb_out[96][106],u_xpb_out[97][106],u_xpb_out[98][106],u_xpb_out[99][106],u_xpb_out[100][106],u_xpb_out[101][106],u_xpb_out[102][106],u_xpb_out[103][106],u_xpb_out[104][106],u_xpb_out[105][106]};

assign col_out_107 = {u_xpb_out[0][107],u_xpb_out[1][107],u_xpb_out[2][107],u_xpb_out[3][107],u_xpb_out[4][107],u_xpb_out[5][107],u_xpb_out[6][107],u_xpb_out[7][107],u_xpb_out[8][107],u_xpb_out[9][107],u_xpb_out[10][107],u_xpb_out[11][107],u_xpb_out[12][107],u_xpb_out[13][107],u_xpb_out[14][107],u_xpb_out[15][107],u_xpb_out[16][107],u_xpb_out[17][107],u_xpb_out[18][107],u_xpb_out[19][107],u_xpb_out[20][107],u_xpb_out[21][107],u_xpb_out[22][107],u_xpb_out[23][107],u_xpb_out[24][107],u_xpb_out[25][107],u_xpb_out[26][107],u_xpb_out[27][107],u_xpb_out[28][107],u_xpb_out[29][107],u_xpb_out[30][107],u_xpb_out[31][107],u_xpb_out[32][107],u_xpb_out[33][107],u_xpb_out[34][107],u_xpb_out[35][107],u_xpb_out[36][107],u_xpb_out[37][107],u_xpb_out[38][107],u_xpb_out[39][107],u_xpb_out[40][107],u_xpb_out[41][107],u_xpb_out[42][107],u_xpb_out[43][107],u_xpb_out[44][107],u_xpb_out[45][107],u_xpb_out[46][107],u_xpb_out[47][107],u_xpb_out[48][107],u_xpb_out[49][107],u_xpb_out[50][107],u_xpb_out[51][107],u_xpb_out[52][107],u_xpb_out[53][107],u_xpb_out[54][107],u_xpb_out[55][107],u_xpb_out[56][107],u_xpb_out[57][107],u_xpb_out[58][107],u_xpb_out[59][107],u_xpb_out[60][107],u_xpb_out[61][107],u_xpb_out[62][107],u_xpb_out[63][107],u_xpb_out[64][107],u_xpb_out[65][107],u_xpb_out[66][107],u_xpb_out[67][107],u_xpb_out[68][107],u_xpb_out[69][107],u_xpb_out[70][107],u_xpb_out[71][107],u_xpb_out[72][107],u_xpb_out[73][107],u_xpb_out[74][107],u_xpb_out[75][107],u_xpb_out[76][107],u_xpb_out[77][107],u_xpb_out[78][107],u_xpb_out[79][107],u_xpb_out[80][107],u_xpb_out[81][107],u_xpb_out[82][107],u_xpb_out[83][107],u_xpb_out[84][107],u_xpb_out[85][107],u_xpb_out[86][107],u_xpb_out[87][107],u_xpb_out[88][107],u_xpb_out[89][107],u_xpb_out[90][107],u_xpb_out[91][107],u_xpb_out[92][107],u_xpb_out[93][107],u_xpb_out[94][107],u_xpb_out[95][107],u_xpb_out[96][107],u_xpb_out[97][107],u_xpb_out[98][107],u_xpb_out[99][107],u_xpb_out[100][107],u_xpb_out[101][107],u_xpb_out[102][107],u_xpb_out[103][107],u_xpb_out[104][107],u_xpb_out[105][107]};

assign col_out_108 = {u_xpb_out[0][108],u_xpb_out[1][108],u_xpb_out[2][108],u_xpb_out[3][108],u_xpb_out[4][108],u_xpb_out[5][108],u_xpb_out[6][108],u_xpb_out[7][108],u_xpb_out[8][108],u_xpb_out[9][108],u_xpb_out[10][108],u_xpb_out[11][108],u_xpb_out[12][108],u_xpb_out[13][108],u_xpb_out[14][108],u_xpb_out[15][108],u_xpb_out[16][108],u_xpb_out[17][108],u_xpb_out[18][108],u_xpb_out[19][108],u_xpb_out[20][108],u_xpb_out[21][108],u_xpb_out[22][108],u_xpb_out[23][108],u_xpb_out[24][108],u_xpb_out[25][108],u_xpb_out[26][108],u_xpb_out[27][108],u_xpb_out[28][108],u_xpb_out[29][108],u_xpb_out[30][108],u_xpb_out[31][108],u_xpb_out[32][108],u_xpb_out[33][108],u_xpb_out[34][108],u_xpb_out[35][108],u_xpb_out[36][108],u_xpb_out[37][108],u_xpb_out[38][108],u_xpb_out[39][108],u_xpb_out[40][108],u_xpb_out[41][108],u_xpb_out[42][108],u_xpb_out[43][108],u_xpb_out[44][108],u_xpb_out[45][108],u_xpb_out[46][108],u_xpb_out[47][108],u_xpb_out[48][108],u_xpb_out[49][108],u_xpb_out[50][108],u_xpb_out[51][108],u_xpb_out[52][108],u_xpb_out[53][108],u_xpb_out[54][108],u_xpb_out[55][108],u_xpb_out[56][108],u_xpb_out[57][108],u_xpb_out[58][108],u_xpb_out[59][108],u_xpb_out[60][108],u_xpb_out[61][108],u_xpb_out[62][108],u_xpb_out[63][108],u_xpb_out[64][108],u_xpb_out[65][108],u_xpb_out[66][108],u_xpb_out[67][108],u_xpb_out[68][108],u_xpb_out[69][108],u_xpb_out[70][108],u_xpb_out[71][108],u_xpb_out[72][108],u_xpb_out[73][108],u_xpb_out[74][108],u_xpb_out[75][108],u_xpb_out[76][108],u_xpb_out[77][108],u_xpb_out[78][108],u_xpb_out[79][108],u_xpb_out[80][108],u_xpb_out[81][108],u_xpb_out[82][108],u_xpb_out[83][108],u_xpb_out[84][108],u_xpb_out[85][108],u_xpb_out[86][108],u_xpb_out[87][108],u_xpb_out[88][108],u_xpb_out[89][108],u_xpb_out[90][108],u_xpb_out[91][108],u_xpb_out[92][108],u_xpb_out[93][108],u_xpb_out[94][108],u_xpb_out[95][108],u_xpb_out[96][108],u_xpb_out[97][108],u_xpb_out[98][108],u_xpb_out[99][108],u_xpb_out[100][108],u_xpb_out[101][108],u_xpb_out[102][108],u_xpb_out[103][108],u_xpb_out[104][108],u_xpb_out[105][108]};

assign col_out_109 = {u_xpb_out[0][109],u_xpb_out[1][109],u_xpb_out[2][109],u_xpb_out[3][109],u_xpb_out[4][109],u_xpb_out[5][109],u_xpb_out[6][109],u_xpb_out[7][109],u_xpb_out[8][109],u_xpb_out[9][109],u_xpb_out[10][109],u_xpb_out[11][109],u_xpb_out[12][109],u_xpb_out[13][109],u_xpb_out[14][109],u_xpb_out[15][109],u_xpb_out[16][109],u_xpb_out[17][109],u_xpb_out[18][109],u_xpb_out[19][109],u_xpb_out[20][109],u_xpb_out[21][109],u_xpb_out[22][109],u_xpb_out[23][109],u_xpb_out[24][109],u_xpb_out[25][109],u_xpb_out[26][109],u_xpb_out[27][109],u_xpb_out[28][109],u_xpb_out[29][109],u_xpb_out[30][109],u_xpb_out[31][109],u_xpb_out[32][109],u_xpb_out[33][109],u_xpb_out[34][109],u_xpb_out[35][109],u_xpb_out[36][109],u_xpb_out[37][109],u_xpb_out[38][109],u_xpb_out[39][109],u_xpb_out[40][109],u_xpb_out[41][109],u_xpb_out[42][109],u_xpb_out[43][109],u_xpb_out[44][109],u_xpb_out[45][109],u_xpb_out[46][109],u_xpb_out[47][109],u_xpb_out[48][109],u_xpb_out[49][109],u_xpb_out[50][109],u_xpb_out[51][109],u_xpb_out[52][109],u_xpb_out[53][109],u_xpb_out[54][109],u_xpb_out[55][109],u_xpb_out[56][109],u_xpb_out[57][109],u_xpb_out[58][109],u_xpb_out[59][109],u_xpb_out[60][109],u_xpb_out[61][109],u_xpb_out[62][109],u_xpb_out[63][109],u_xpb_out[64][109],u_xpb_out[65][109],u_xpb_out[66][109],u_xpb_out[67][109],u_xpb_out[68][109],u_xpb_out[69][109],u_xpb_out[70][109],u_xpb_out[71][109],u_xpb_out[72][109],u_xpb_out[73][109],u_xpb_out[74][109],u_xpb_out[75][109],u_xpb_out[76][109],u_xpb_out[77][109],u_xpb_out[78][109],u_xpb_out[79][109],u_xpb_out[80][109],u_xpb_out[81][109],u_xpb_out[82][109],u_xpb_out[83][109],u_xpb_out[84][109],u_xpb_out[85][109],u_xpb_out[86][109],u_xpb_out[87][109],u_xpb_out[88][109],u_xpb_out[89][109],u_xpb_out[90][109],u_xpb_out[91][109],u_xpb_out[92][109],u_xpb_out[93][109],u_xpb_out[94][109],u_xpb_out[95][109],u_xpb_out[96][109],u_xpb_out[97][109],u_xpb_out[98][109],u_xpb_out[99][109],u_xpb_out[100][109],u_xpb_out[101][109],u_xpb_out[102][109],u_xpb_out[103][109],u_xpb_out[104][109],u_xpb_out[105][109]};

assign col_out_110 = {u_xpb_out[0][110],u_xpb_out[1][110],u_xpb_out[2][110],u_xpb_out[3][110],u_xpb_out[4][110],u_xpb_out[5][110],u_xpb_out[6][110],u_xpb_out[7][110],u_xpb_out[8][110],u_xpb_out[9][110],u_xpb_out[10][110],u_xpb_out[11][110],u_xpb_out[12][110],u_xpb_out[13][110],u_xpb_out[14][110],u_xpb_out[15][110],u_xpb_out[16][110],u_xpb_out[17][110],u_xpb_out[18][110],u_xpb_out[19][110],u_xpb_out[20][110],u_xpb_out[21][110],u_xpb_out[22][110],u_xpb_out[23][110],u_xpb_out[24][110],u_xpb_out[25][110],u_xpb_out[26][110],u_xpb_out[27][110],u_xpb_out[28][110],u_xpb_out[29][110],u_xpb_out[30][110],u_xpb_out[31][110],u_xpb_out[32][110],u_xpb_out[33][110],u_xpb_out[34][110],u_xpb_out[35][110],u_xpb_out[36][110],u_xpb_out[37][110],u_xpb_out[38][110],u_xpb_out[39][110],u_xpb_out[40][110],u_xpb_out[41][110],u_xpb_out[42][110],u_xpb_out[43][110],u_xpb_out[44][110],u_xpb_out[45][110],u_xpb_out[46][110],u_xpb_out[47][110],u_xpb_out[48][110],u_xpb_out[49][110],u_xpb_out[50][110],u_xpb_out[51][110],u_xpb_out[52][110],u_xpb_out[53][110],u_xpb_out[54][110],u_xpb_out[55][110],u_xpb_out[56][110],u_xpb_out[57][110],u_xpb_out[58][110],u_xpb_out[59][110],u_xpb_out[60][110],u_xpb_out[61][110],u_xpb_out[62][110],u_xpb_out[63][110],u_xpb_out[64][110],u_xpb_out[65][110],u_xpb_out[66][110],u_xpb_out[67][110],u_xpb_out[68][110],u_xpb_out[69][110],u_xpb_out[70][110],u_xpb_out[71][110],u_xpb_out[72][110],u_xpb_out[73][110],u_xpb_out[74][110],u_xpb_out[75][110],u_xpb_out[76][110],u_xpb_out[77][110],u_xpb_out[78][110],u_xpb_out[79][110],u_xpb_out[80][110],u_xpb_out[81][110],u_xpb_out[82][110],u_xpb_out[83][110],u_xpb_out[84][110],u_xpb_out[85][110],u_xpb_out[86][110],u_xpb_out[87][110],u_xpb_out[88][110],u_xpb_out[89][110],u_xpb_out[90][110],u_xpb_out[91][110],u_xpb_out[92][110],u_xpb_out[93][110],u_xpb_out[94][110],u_xpb_out[95][110],u_xpb_out[96][110],u_xpb_out[97][110],u_xpb_out[98][110],u_xpb_out[99][110],u_xpb_out[100][110],u_xpb_out[101][110],u_xpb_out[102][110],u_xpb_out[103][110],u_xpb_out[104][110],u_xpb_out[105][110]};

assign col_out_111 = {u_xpb_out[0][111],u_xpb_out[1][111],u_xpb_out[2][111],u_xpb_out[3][111],u_xpb_out[4][111],u_xpb_out[5][111],u_xpb_out[6][111],u_xpb_out[7][111],u_xpb_out[8][111],u_xpb_out[9][111],u_xpb_out[10][111],u_xpb_out[11][111],u_xpb_out[12][111],u_xpb_out[13][111],u_xpb_out[14][111],u_xpb_out[15][111],u_xpb_out[16][111],u_xpb_out[17][111],u_xpb_out[18][111],u_xpb_out[19][111],u_xpb_out[20][111],u_xpb_out[21][111],u_xpb_out[22][111],u_xpb_out[23][111],u_xpb_out[24][111],u_xpb_out[25][111],u_xpb_out[26][111],u_xpb_out[27][111],u_xpb_out[28][111],u_xpb_out[29][111],u_xpb_out[30][111],u_xpb_out[31][111],u_xpb_out[32][111],u_xpb_out[33][111],u_xpb_out[34][111],u_xpb_out[35][111],u_xpb_out[36][111],u_xpb_out[37][111],u_xpb_out[38][111],u_xpb_out[39][111],u_xpb_out[40][111],u_xpb_out[41][111],u_xpb_out[42][111],u_xpb_out[43][111],u_xpb_out[44][111],u_xpb_out[45][111],u_xpb_out[46][111],u_xpb_out[47][111],u_xpb_out[48][111],u_xpb_out[49][111],u_xpb_out[50][111],u_xpb_out[51][111],u_xpb_out[52][111],u_xpb_out[53][111],u_xpb_out[54][111],u_xpb_out[55][111],u_xpb_out[56][111],u_xpb_out[57][111],u_xpb_out[58][111],u_xpb_out[59][111],u_xpb_out[60][111],u_xpb_out[61][111],u_xpb_out[62][111],u_xpb_out[63][111],u_xpb_out[64][111],u_xpb_out[65][111],u_xpb_out[66][111],u_xpb_out[67][111],u_xpb_out[68][111],u_xpb_out[69][111],u_xpb_out[70][111],u_xpb_out[71][111],u_xpb_out[72][111],u_xpb_out[73][111],u_xpb_out[74][111],u_xpb_out[75][111],u_xpb_out[76][111],u_xpb_out[77][111],u_xpb_out[78][111],u_xpb_out[79][111],u_xpb_out[80][111],u_xpb_out[81][111],u_xpb_out[82][111],u_xpb_out[83][111],u_xpb_out[84][111],u_xpb_out[85][111],u_xpb_out[86][111],u_xpb_out[87][111],u_xpb_out[88][111],u_xpb_out[89][111],u_xpb_out[90][111],u_xpb_out[91][111],u_xpb_out[92][111],u_xpb_out[93][111],u_xpb_out[94][111],u_xpb_out[95][111],u_xpb_out[96][111],u_xpb_out[97][111],u_xpb_out[98][111],u_xpb_out[99][111],u_xpb_out[100][111],u_xpb_out[101][111],u_xpb_out[102][111],u_xpb_out[103][111],u_xpb_out[104][111],u_xpb_out[105][111]};

assign col_out_112 = {u_xpb_out[0][112],u_xpb_out[1][112],u_xpb_out[2][112],u_xpb_out[3][112],u_xpb_out[4][112],u_xpb_out[5][112],u_xpb_out[6][112],u_xpb_out[7][112],u_xpb_out[8][112],u_xpb_out[9][112],u_xpb_out[10][112],u_xpb_out[11][112],u_xpb_out[12][112],u_xpb_out[13][112],u_xpb_out[14][112],u_xpb_out[15][112],u_xpb_out[16][112],u_xpb_out[17][112],u_xpb_out[18][112],u_xpb_out[19][112],u_xpb_out[20][112],u_xpb_out[21][112],u_xpb_out[22][112],u_xpb_out[23][112],u_xpb_out[24][112],u_xpb_out[25][112],u_xpb_out[26][112],u_xpb_out[27][112],u_xpb_out[28][112],u_xpb_out[29][112],u_xpb_out[30][112],u_xpb_out[31][112],u_xpb_out[32][112],u_xpb_out[33][112],u_xpb_out[34][112],u_xpb_out[35][112],u_xpb_out[36][112],u_xpb_out[37][112],u_xpb_out[38][112],u_xpb_out[39][112],u_xpb_out[40][112],u_xpb_out[41][112],u_xpb_out[42][112],u_xpb_out[43][112],u_xpb_out[44][112],u_xpb_out[45][112],u_xpb_out[46][112],u_xpb_out[47][112],u_xpb_out[48][112],u_xpb_out[49][112],u_xpb_out[50][112],u_xpb_out[51][112],u_xpb_out[52][112],u_xpb_out[53][112],u_xpb_out[54][112],u_xpb_out[55][112],u_xpb_out[56][112],u_xpb_out[57][112],u_xpb_out[58][112],u_xpb_out[59][112],u_xpb_out[60][112],u_xpb_out[61][112],u_xpb_out[62][112],u_xpb_out[63][112],u_xpb_out[64][112],u_xpb_out[65][112],u_xpb_out[66][112],u_xpb_out[67][112],u_xpb_out[68][112],u_xpb_out[69][112],u_xpb_out[70][112],u_xpb_out[71][112],u_xpb_out[72][112],u_xpb_out[73][112],u_xpb_out[74][112],u_xpb_out[75][112],u_xpb_out[76][112],u_xpb_out[77][112],u_xpb_out[78][112],u_xpb_out[79][112],u_xpb_out[80][112],u_xpb_out[81][112],u_xpb_out[82][112],u_xpb_out[83][112],u_xpb_out[84][112],u_xpb_out[85][112],u_xpb_out[86][112],u_xpb_out[87][112],u_xpb_out[88][112],u_xpb_out[89][112],u_xpb_out[90][112],u_xpb_out[91][112],u_xpb_out[92][112],u_xpb_out[93][112],u_xpb_out[94][112],u_xpb_out[95][112],u_xpb_out[96][112],u_xpb_out[97][112],u_xpb_out[98][112],u_xpb_out[99][112],u_xpb_out[100][112],u_xpb_out[101][112],u_xpb_out[102][112],u_xpb_out[103][112],u_xpb_out[104][112],u_xpb_out[105][112]};

assign col_out_113 = {u_xpb_out[0][113],u_xpb_out[1][113],u_xpb_out[2][113],u_xpb_out[3][113],u_xpb_out[4][113],u_xpb_out[5][113],u_xpb_out[6][113],u_xpb_out[7][113],u_xpb_out[8][113],u_xpb_out[9][113],u_xpb_out[10][113],u_xpb_out[11][113],u_xpb_out[12][113],u_xpb_out[13][113],u_xpb_out[14][113],u_xpb_out[15][113],u_xpb_out[16][113],u_xpb_out[17][113],u_xpb_out[18][113],u_xpb_out[19][113],u_xpb_out[20][113],u_xpb_out[21][113],u_xpb_out[22][113],u_xpb_out[23][113],u_xpb_out[24][113],u_xpb_out[25][113],u_xpb_out[26][113],u_xpb_out[27][113],u_xpb_out[28][113],u_xpb_out[29][113],u_xpb_out[30][113],u_xpb_out[31][113],u_xpb_out[32][113],u_xpb_out[33][113],u_xpb_out[34][113],u_xpb_out[35][113],u_xpb_out[36][113],u_xpb_out[37][113],u_xpb_out[38][113],u_xpb_out[39][113],u_xpb_out[40][113],u_xpb_out[41][113],u_xpb_out[42][113],u_xpb_out[43][113],u_xpb_out[44][113],u_xpb_out[45][113],u_xpb_out[46][113],u_xpb_out[47][113],u_xpb_out[48][113],u_xpb_out[49][113],u_xpb_out[50][113],u_xpb_out[51][113],u_xpb_out[52][113],u_xpb_out[53][113],u_xpb_out[54][113],u_xpb_out[55][113],u_xpb_out[56][113],u_xpb_out[57][113],u_xpb_out[58][113],u_xpb_out[59][113],u_xpb_out[60][113],u_xpb_out[61][113],u_xpb_out[62][113],u_xpb_out[63][113],u_xpb_out[64][113],u_xpb_out[65][113],u_xpb_out[66][113],u_xpb_out[67][113],u_xpb_out[68][113],u_xpb_out[69][113],u_xpb_out[70][113],u_xpb_out[71][113],u_xpb_out[72][113],u_xpb_out[73][113],u_xpb_out[74][113],u_xpb_out[75][113],u_xpb_out[76][113],u_xpb_out[77][113],u_xpb_out[78][113],u_xpb_out[79][113],u_xpb_out[80][113],u_xpb_out[81][113],u_xpb_out[82][113],u_xpb_out[83][113],u_xpb_out[84][113],u_xpb_out[85][113],u_xpb_out[86][113],u_xpb_out[87][113],u_xpb_out[88][113],u_xpb_out[89][113],u_xpb_out[90][113],u_xpb_out[91][113],u_xpb_out[92][113],u_xpb_out[93][113],u_xpb_out[94][113],u_xpb_out[95][113],u_xpb_out[96][113],u_xpb_out[97][113],u_xpb_out[98][113],u_xpb_out[99][113],u_xpb_out[100][113],u_xpb_out[101][113],u_xpb_out[102][113],u_xpb_out[103][113],u_xpb_out[104][113],u_xpb_out[105][113]};

assign col_out_114 = {u_xpb_out[0][114],u_xpb_out[1][114],u_xpb_out[2][114],u_xpb_out[3][114],u_xpb_out[4][114],u_xpb_out[5][114],u_xpb_out[6][114],u_xpb_out[7][114],u_xpb_out[8][114],u_xpb_out[9][114],u_xpb_out[10][114],u_xpb_out[11][114],u_xpb_out[12][114],u_xpb_out[13][114],u_xpb_out[14][114],u_xpb_out[15][114],u_xpb_out[16][114],u_xpb_out[17][114],u_xpb_out[18][114],u_xpb_out[19][114],u_xpb_out[20][114],u_xpb_out[21][114],u_xpb_out[22][114],u_xpb_out[23][114],u_xpb_out[24][114],u_xpb_out[25][114],u_xpb_out[26][114],u_xpb_out[27][114],u_xpb_out[28][114],u_xpb_out[29][114],u_xpb_out[30][114],u_xpb_out[31][114],u_xpb_out[32][114],u_xpb_out[33][114],u_xpb_out[34][114],u_xpb_out[35][114],u_xpb_out[36][114],u_xpb_out[37][114],u_xpb_out[38][114],u_xpb_out[39][114],u_xpb_out[40][114],u_xpb_out[41][114],u_xpb_out[42][114],u_xpb_out[43][114],u_xpb_out[44][114],u_xpb_out[45][114],u_xpb_out[46][114],u_xpb_out[47][114],u_xpb_out[48][114],u_xpb_out[49][114],u_xpb_out[50][114],u_xpb_out[51][114],u_xpb_out[52][114],u_xpb_out[53][114],u_xpb_out[54][114],u_xpb_out[55][114],u_xpb_out[56][114],u_xpb_out[57][114],u_xpb_out[58][114],u_xpb_out[59][114],u_xpb_out[60][114],u_xpb_out[61][114],u_xpb_out[62][114],u_xpb_out[63][114],u_xpb_out[64][114],u_xpb_out[65][114],u_xpb_out[66][114],u_xpb_out[67][114],u_xpb_out[68][114],u_xpb_out[69][114],u_xpb_out[70][114],u_xpb_out[71][114],u_xpb_out[72][114],u_xpb_out[73][114],u_xpb_out[74][114],u_xpb_out[75][114],u_xpb_out[76][114],u_xpb_out[77][114],u_xpb_out[78][114],u_xpb_out[79][114],u_xpb_out[80][114],u_xpb_out[81][114],u_xpb_out[82][114],u_xpb_out[83][114],u_xpb_out[84][114],u_xpb_out[85][114],u_xpb_out[86][114],u_xpb_out[87][114],u_xpb_out[88][114],u_xpb_out[89][114],u_xpb_out[90][114],u_xpb_out[91][114],u_xpb_out[92][114],u_xpb_out[93][114],u_xpb_out[94][114],u_xpb_out[95][114],u_xpb_out[96][114],u_xpb_out[97][114],u_xpb_out[98][114],u_xpb_out[99][114],u_xpb_out[100][114],u_xpb_out[101][114],u_xpb_out[102][114],u_xpb_out[103][114],u_xpb_out[104][114],u_xpb_out[105][114]};

assign col_out_115 = {u_xpb_out[0][115],u_xpb_out[1][115],u_xpb_out[2][115],u_xpb_out[3][115],u_xpb_out[4][115],u_xpb_out[5][115],u_xpb_out[6][115],u_xpb_out[7][115],u_xpb_out[8][115],u_xpb_out[9][115],u_xpb_out[10][115],u_xpb_out[11][115],u_xpb_out[12][115],u_xpb_out[13][115],u_xpb_out[14][115],u_xpb_out[15][115],u_xpb_out[16][115],u_xpb_out[17][115],u_xpb_out[18][115],u_xpb_out[19][115],u_xpb_out[20][115],u_xpb_out[21][115],u_xpb_out[22][115],u_xpb_out[23][115],u_xpb_out[24][115],u_xpb_out[25][115],u_xpb_out[26][115],u_xpb_out[27][115],u_xpb_out[28][115],u_xpb_out[29][115],u_xpb_out[30][115],u_xpb_out[31][115],u_xpb_out[32][115],u_xpb_out[33][115],u_xpb_out[34][115],u_xpb_out[35][115],u_xpb_out[36][115],u_xpb_out[37][115],u_xpb_out[38][115],u_xpb_out[39][115],u_xpb_out[40][115],u_xpb_out[41][115],u_xpb_out[42][115],u_xpb_out[43][115],u_xpb_out[44][115],u_xpb_out[45][115],u_xpb_out[46][115],u_xpb_out[47][115],u_xpb_out[48][115],u_xpb_out[49][115],u_xpb_out[50][115],u_xpb_out[51][115],u_xpb_out[52][115],u_xpb_out[53][115],u_xpb_out[54][115],u_xpb_out[55][115],u_xpb_out[56][115],u_xpb_out[57][115],u_xpb_out[58][115],u_xpb_out[59][115],u_xpb_out[60][115],u_xpb_out[61][115],u_xpb_out[62][115],u_xpb_out[63][115],u_xpb_out[64][115],u_xpb_out[65][115],u_xpb_out[66][115],u_xpb_out[67][115],u_xpb_out[68][115],u_xpb_out[69][115],u_xpb_out[70][115],u_xpb_out[71][115],u_xpb_out[72][115],u_xpb_out[73][115],u_xpb_out[74][115],u_xpb_out[75][115],u_xpb_out[76][115],u_xpb_out[77][115],u_xpb_out[78][115],u_xpb_out[79][115],u_xpb_out[80][115],u_xpb_out[81][115],u_xpb_out[82][115],u_xpb_out[83][115],u_xpb_out[84][115],u_xpb_out[85][115],u_xpb_out[86][115],u_xpb_out[87][115],u_xpb_out[88][115],u_xpb_out[89][115],u_xpb_out[90][115],u_xpb_out[91][115],u_xpb_out[92][115],u_xpb_out[93][115],u_xpb_out[94][115],u_xpb_out[95][115],u_xpb_out[96][115],u_xpb_out[97][115],u_xpb_out[98][115],u_xpb_out[99][115],u_xpb_out[100][115],u_xpb_out[101][115],u_xpb_out[102][115],u_xpb_out[103][115],u_xpb_out[104][115],u_xpb_out[105][115]};

assign col_out_116 = {u_xpb_out[0][116],u_xpb_out[1][116],u_xpb_out[2][116],u_xpb_out[3][116],u_xpb_out[4][116],u_xpb_out[5][116],u_xpb_out[6][116],u_xpb_out[7][116],u_xpb_out[8][116],u_xpb_out[9][116],u_xpb_out[10][116],u_xpb_out[11][116],u_xpb_out[12][116],u_xpb_out[13][116],u_xpb_out[14][116],u_xpb_out[15][116],u_xpb_out[16][116],u_xpb_out[17][116],u_xpb_out[18][116],u_xpb_out[19][116],u_xpb_out[20][116],u_xpb_out[21][116],u_xpb_out[22][116],u_xpb_out[23][116],u_xpb_out[24][116],u_xpb_out[25][116],u_xpb_out[26][116],u_xpb_out[27][116],u_xpb_out[28][116],u_xpb_out[29][116],u_xpb_out[30][116],u_xpb_out[31][116],u_xpb_out[32][116],u_xpb_out[33][116],u_xpb_out[34][116],u_xpb_out[35][116],u_xpb_out[36][116],u_xpb_out[37][116],u_xpb_out[38][116],u_xpb_out[39][116],u_xpb_out[40][116],u_xpb_out[41][116],u_xpb_out[42][116],u_xpb_out[43][116],u_xpb_out[44][116],u_xpb_out[45][116],u_xpb_out[46][116],u_xpb_out[47][116],u_xpb_out[48][116],u_xpb_out[49][116],u_xpb_out[50][116],u_xpb_out[51][116],u_xpb_out[52][116],u_xpb_out[53][116],u_xpb_out[54][116],u_xpb_out[55][116],u_xpb_out[56][116],u_xpb_out[57][116],u_xpb_out[58][116],u_xpb_out[59][116],u_xpb_out[60][116],u_xpb_out[61][116],u_xpb_out[62][116],u_xpb_out[63][116],u_xpb_out[64][116],u_xpb_out[65][116],u_xpb_out[66][116],u_xpb_out[67][116],u_xpb_out[68][116],u_xpb_out[69][116],u_xpb_out[70][116],u_xpb_out[71][116],u_xpb_out[72][116],u_xpb_out[73][116],u_xpb_out[74][116],u_xpb_out[75][116],u_xpb_out[76][116],u_xpb_out[77][116],u_xpb_out[78][116],u_xpb_out[79][116],u_xpb_out[80][116],u_xpb_out[81][116],u_xpb_out[82][116],u_xpb_out[83][116],u_xpb_out[84][116],u_xpb_out[85][116],u_xpb_out[86][116],u_xpb_out[87][116],u_xpb_out[88][116],u_xpb_out[89][116],u_xpb_out[90][116],u_xpb_out[91][116],u_xpb_out[92][116],u_xpb_out[93][116],u_xpb_out[94][116],u_xpb_out[95][116],u_xpb_out[96][116],u_xpb_out[97][116],u_xpb_out[98][116],u_xpb_out[99][116],u_xpb_out[100][116],u_xpb_out[101][116],u_xpb_out[102][116],u_xpb_out[103][116],u_xpb_out[104][116],u_xpb_out[105][116]};

assign col_out_117 = {u_xpb_out[0][117],u_xpb_out[1][117],u_xpb_out[2][117],u_xpb_out[3][117],u_xpb_out[4][117],u_xpb_out[5][117],u_xpb_out[6][117],u_xpb_out[7][117],u_xpb_out[8][117],u_xpb_out[9][117],u_xpb_out[10][117],u_xpb_out[11][117],u_xpb_out[12][117],u_xpb_out[13][117],u_xpb_out[14][117],u_xpb_out[15][117],u_xpb_out[16][117],u_xpb_out[17][117],u_xpb_out[18][117],u_xpb_out[19][117],u_xpb_out[20][117],u_xpb_out[21][117],u_xpb_out[22][117],u_xpb_out[23][117],u_xpb_out[24][117],u_xpb_out[25][117],u_xpb_out[26][117],u_xpb_out[27][117],u_xpb_out[28][117],u_xpb_out[29][117],u_xpb_out[30][117],u_xpb_out[31][117],u_xpb_out[32][117],u_xpb_out[33][117],u_xpb_out[34][117],u_xpb_out[35][117],u_xpb_out[36][117],u_xpb_out[37][117],u_xpb_out[38][117],u_xpb_out[39][117],u_xpb_out[40][117],u_xpb_out[41][117],u_xpb_out[42][117],u_xpb_out[43][117],u_xpb_out[44][117],u_xpb_out[45][117],u_xpb_out[46][117],u_xpb_out[47][117],u_xpb_out[48][117],u_xpb_out[49][117],u_xpb_out[50][117],u_xpb_out[51][117],u_xpb_out[52][117],u_xpb_out[53][117],u_xpb_out[54][117],u_xpb_out[55][117],u_xpb_out[56][117],u_xpb_out[57][117],u_xpb_out[58][117],u_xpb_out[59][117],u_xpb_out[60][117],u_xpb_out[61][117],u_xpb_out[62][117],u_xpb_out[63][117],u_xpb_out[64][117],u_xpb_out[65][117],u_xpb_out[66][117],u_xpb_out[67][117],u_xpb_out[68][117],u_xpb_out[69][117],u_xpb_out[70][117],u_xpb_out[71][117],u_xpb_out[72][117],u_xpb_out[73][117],u_xpb_out[74][117],u_xpb_out[75][117],u_xpb_out[76][117],u_xpb_out[77][117],u_xpb_out[78][117],u_xpb_out[79][117],u_xpb_out[80][117],u_xpb_out[81][117],u_xpb_out[82][117],u_xpb_out[83][117],u_xpb_out[84][117],u_xpb_out[85][117],u_xpb_out[86][117],u_xpb_out[87][117],u_xpb_out[88][117],u_xpb_out[89][117],u_xpb_out[90][117],u_xpb_out[91][117],u_xpb_out[92][117],u_xpb_out[93][117],u_xpb_out[94][117],u_xpb_out[95][117],u_xpb_out[96][117],u_xpb_out[97][117],u_xpb_out[98][117],u_xpb_out[99][117],u_xpb_out[100][117],u_xpb_out[101][117],u_xpb_out[102][117],u_xpb_out[103][117],u_xpb_out[104][117],u_xpb_out[105][117]};

assign col_out_118 = {u_xpb_out[0][118],u_xpb_out[1][118],u_xpb_out[2][118],u_xpb_out[3][118],u_xpb_out[4][118],u_xpb_out[5][118],u_xpb_out[6][118],u_xpb_out[7][118],u_xpb_out[8][118],u_xpb_out[9][118],u_xpb_out[10][118],u_xpb_out[11][118],u_xpb_out[12][118],u_xpb_out[13][118],u_xpb_out[14][118],u_xpb_out[15][118],u_xpb_out[16][118],u_xpb_out[17][118],u_xpb_out[18][118],u_xpb_out[19][118],u_xpb_out[20][118],u_xpb_out[21][118],u_xpb_out[22][118],u_xpb_out[23][118],u_xpb_out[24][118],u_xpb_out[25][118],u_xpb_out[26][118],u_xpb_out[27][118],u_xpb_out[28][118],u_xpb_out[29][118],u_xpb_out[30][118],u_xpb_out[31][118],u_xpb_out[32][118],u_xpb_out[33][118],u_xpb_out[34][118],u_xpb_out[35][118],u_xpb_out[36][118],u_xpb_out[37][118],u_xpb_out[38][118],u_xpb_out[39][118],u_xpb_out[40][118],u_xpb_out[41][118],u_xpb_out[42][118],u_xpb_out[43][118],u_xpb_out[44][118],u_xpb_out[45][118],u_xpb_out[46][118],u_xpb_out[47][118],u_xpb_out[48][118],u_xpb_out[49][118],u_xpb_out[50][118],u_xpb_out[51][118],u_xpb_out[52][118],u_xpb_out[53][118],u_xpb_out[54][118],u_xpb_out[55][118],u_xpb_out[56][118],u_xpb_out[57][118],u_xpb_out[58][118],u_xpb_out[59][118],u_xpb_out[60][118],u_xpb_out[61][118],u_xpb_out[62][118],u_xpb_out[63][118],u_xpb_out[64][118],u_xpb_out[65][118],u_xpb_out[66][118],u_xpb_out[67][118],u_xpb_out[68][118],u_xpb_out[69][118],u_xpb_out[70][118],u_xpb_out[71][118],u_xpb_out[72][118],u_xpb_out[73][118],u_xpb_out[74][118],u_xpb_out[75][118],u_xpb_out[76][118],u_xpb_out[77][118],u_xpb_out[78][118],u_xpb_out[79][118],u_xpb_out[80][118],u_xpb_out[81][118],u_xpb_out[82][118],u_xpb_out[83][118],u_xpb_out[84][118],u_xpb_out[85][118],u_xpb_out[86][118],u_xpb_out[87][118],u_xpb_out[88][118],u_xpb_out[89][118],u_xpb_out[90][118],u_xpb_out[91][118],u_xpb_out[92][118],u_xpb_out[93][118],u_xpb_out[94][118],u_xpb_out[95][118],u_xpb_out[96][118],u_xpb_out[97][118],u_xpb_out[98][118],u_xpb_out[99][118],u_xpb_out[100][118],u_xpb_out[101][118],u_xpb_out[102][118],u_xpb_out[103][118],u_xpb_out[104][118],u_xpb_out[105][118]};

assign col_out_119 = {u_xpb_out[0][119],u_xpb_out[1][119],u_xpb_out[2][119],u_xpb_out[3][119],u_xpb_out[4][119],u_xpb_out[5][119],u_xpb_out[6][119],u_xpb_out[7][119],u_xpb_out[8][119],u_xpb_out[9][119],u_xpb_out[10][119],u_xpb_out[11][119],u_xpb_out[12][119],u_xpb_out[13][119],u_xpb_out[14][119],u_xpb_out[15][119],u_xpb_out[16][119],u_xpb_out[17][119],u_xpb_out[18][119],u_xpb_out[19][119],u_xpb_out[20][119],u_xpb_out[21][119],u_xpb_out[22][119],u_xpb_out[23][119],u_xpb_out[24][119],u_xpb_out[25][119],u_xpb_out[26][119],u_xpb_out[27][119],u_xpb_out[28][119],u_xpb_out[29][119],u_xpb_out[30][119],u_xpb_out[31][119],u_xpb_out[32][119],u_xpb_out[33][119],u_xpb_out[34][119],u_xpb_out[35][119],u_xpb_out[36][119],u_xpb_out[37][119],u_xpb_out[38][119],u_xpb_out[39][119],u_xpb_out[40][119],u_xpb_out[41][119],u_xpb_out[42][119],u_xpb_out[43][119],u_xpb_out[44][119],u_xpb_out[45][119],u_xpb_out[46][119],u_xpb_out[47][119],u_xpb_out[48][119],u_xpb_out[49][119],u_xpb_out[50][119],u_xpb_out[51][119],u_xpb_out[52][119],u_xpb_out[53][119],u_xpb_out[54][119],u_xpb_out[55][119],u_xpb_out[56][119],u_xpb_out[57][119],u_xpb_out[58][119],u_xpb_out[59][119],u_xpb_out[60][119],u_xpb_out[61][119],u_xpb_out[62][119],u_xpb_out[63][119],u_xpb_out[64][119],u_xpb_out[65][119],u_xpb_out[66][119],u_xpb_out[67][119],u_xpb_out[68][119],u_xpb_out[69][119],u_xpb_out[70][119],u_xpb_out[71][119],u_xpb_out[72][119],u_xpb_out[73][119],u_xpb_out[74][119],u_xpb_out[75][119],u_xpb_out[76][119],u_xpb_out[77][119],u_xpb_out[78][119],u_xpb_out[79][119],u_xpb_out[80][119],u_xpb_out[81][119],u_xpb_out[82][119],u_xpb_out[83][119],u_xpb_out[84][119],u_xpb_out[85][119],u_xpb_out[86][119],u_xpb_out[87][119],u_xpb_out[88][119],u_xpb_out[89][119],u_xpb_out[90][119],u_xpb_out[91][119],u_xpb_out[92][119],u_xpb_out[93][119],u_xpb_out[94][119],u_xpb_out[95][119],u_xpb_out[96][119],u_xpb_out[97][119],u_xpb_out[98][119],u_xpb_out[99][119],u_xpb_out[100][119],u_xpb_out[101][119],u_xpb_out[102][119],u_xpb_out[103][119],u_xpb_out[104][119],u_xpb_out[105][119]};

assign col_out_120 = {u_xpb_out[0][120],u_xpb_out[1][120],u_xpb_out[2][120],u_xpb_out[3][120],u_xpb_out[4][120],u_xpb_out[5][120],u_xpb_out[6][120],u_xpb_out[7][120],u_xpb_out[8][120],u_xpb_out[9][120],u_xpb_out[10][120],u_xpb_out[11][120],u_xpb_out[12][120],u_xpb_out[13][120],u_xpb_out[14][120],u_xpb_out[15][120],u_xpb_out[16][120],u_xpb_out[17][120],u_xpb_out[18][120],u_xpb_out[19][120],u_xpb_out[20][120],u_xpb_out[21][120],u_xpb_out[22][120],u_xpb_out[23][120],u_xpb_out[24][120],u_xpb_out[25][120],u_xpb_out[26][120],u_xpb_out[27][120],u_xpb_out[28][120],u_xpb_out[29][120],u_xpb_out[30][120],u_xpb_out[31][120],u_xpb_out[32][120],u_xpb_out[33][120],u_xpb_out[34][120],u_xpb_out[35][120],u_xpb_out[36][120],u_xpb_out[37][120],u_xpb_out[38][120],u_xpb_out[39][120],u_xpb_out[40][120],u_xpb_out[41][120],u_xpb_out[42][120],u_xpb_out[43][120],u_xpb_out[44][120],u_xpb_out[45][120],u_xpb_out[46][120],u_xpb_out[47][120],u_xpb_out[48][120],u_xpb_out[49][120],u_xpb_out[50][120],u_xpb_out[51][120],u_xpb_out[52][120],u_xpb_out[53][120],u_xpb_out[54][120],u_xpb_out[55][120],u_xpb_out[56][120],u_xpb_out[57][120],u_xpb_out[58][120],u_xpb_out[59][120],u_xpb_out[60][120],u_xpb_out[61][120],u_xpb_out[62][120],u_xpb_out[63][120],u_xpb_out[64][120],u_xpb_out[65][120],u_xpb_out[66][120],u_xpb_out[67][120],u_xpb_out[68][120],u_xpb_out[69][120],u_xpb_out[70][120],u_xpb_out[71][120],u_xpb_out[72][120],u_xpb_out[73][120],u_xpb_out[74][120],u_xpb_out[75][120],u_xpb_out[76][120],u_xpb_out[77][120],u_xpb_out[78][120],u_xpb_out[79][120],u_xpb_out[80][120],u_xpb_out[81][120],u_xpb_out[82][120],u_xpb_out[83][120],u_xpb_out[84][120],u_xpb_out[85][120],u_xpb_out[86][120],u_xpb_out[87][120],u_xpb_out[88][120],u_xpb_out[89][120],u_xpb_out[90][120],u_xpb_out[91][120],u_xpb_out[92][120],u_xpb_out[93][120],u_xpb_out[94][120],u_xpb_out[95][120],u_xpb_out[96][120],u_xpb_out[97][120],u_xpb_out[98][120],u_xpb_out[99][120],u_xpb_out[100][120],u_xpb_out[101][120],u_xpb_out[102][120],u_xpb_out[103][120],u_xpb_out[104][120],u_xpb_out[105][120]};

assign col_out_121 = {u_xpb_out[0][121],u_xpb_out[1][121],u_xpb_out[2][121],u_xpb_out[3][121],u_xpb_out[4][121],u_xpb_out[5][121],u_xpb_out[6][121],u_xpb_out[7][121],u_xpb_out[8][121],u_xpb_out[9][121],u_xpb_out[10][121],u_xpb_out[11][121],u_xpb_out[12][121],u_xpb_out[13][121],u_xpb_out[14][121],u_xpb_out[15][121],u_xpb_out[16][121],u_xpb_out[17][121],u_xpb_out[18][121],u_xpb_out[19][121],u_xpb_out[20][121],u_xpb_out[21][121],u_xpb_out[22][121],u_xpb_out[23][121],u_xpb_out[24][121],u_xpb_out[25][121],u_xpb_out[26][121],u_xpb_out[27][121],u_xpb_out[28][121],u_xpb_out[29][121],u_xpb_out[30][121],u_xpb_out[31][121],u_xpb_out[32][121],u_xpb_out[33][121],u_xpb_out[34][121],u_xpb_out[35][121],u_xpb_out[36][121],u_xpb_out[37][121],u_xpb_out[38][121],u_xpb_out[39][121],u_xpb_out[40][121],u_xpb_out[41][121],u_xpb_out[42][121],u_xpb_out[43][121],u_xpb_out[44][121],u_xpb_out[45][121],u_xpb_out[46][121],u_xpb_out[47][121],u_xpb_out[48][121],u_xpb_out[49][121],u_xpb_out[50][121],u_xpb_out[51][121],u_xpb_out[52][121],u_xpb_out[53][121],u_xpb_out[54][121],u_xpb_out[55][121],u_xpb_out[56][121],u_xpb_out[57][121],u_xpb_out[58][121],u_xpb_out[59][121],u_xpb_out[60][121],u_xpb_out[61][121],u_xpb_out[62][121],u_xpb_out[63][121],u_xpb_out[64][121],u_xpb_out[65][121],u_xpb_out[66][121],u_xpb_out[67][121],u_xpb_out[68][121],u_xpb_out[69][121],u_xpb_out[70][121],u_xpb_out[71][121],u_xpb_out[72][121],u_xpb_out[73][121],u_xpb_out[74][121],u_xpb_out[75][121],u_xpb_out[76][121],u_xpb_out[77][121],u_xpb_out[78][121],u_xpb_out[79][121],u_xpb_out[80][121],u_xpb_out[81][121],u_xpb_out[82][121],u_xpb_out[83][121],u_xpb_out[84][121],u_xpb_out[85][121],u_xpb_out[86][121],u_xpb_out[87][121],u_xpb_out[88][121],u_xpb_out[89][121],u_xpb_out[90][121],u_xpb_out[91][121],u_xpb_out[92][121],u_xpb_out[93][121],u_xpb_out[94][121],u_xpb_out[95][121],u_xpb_out[96][121],u_xpb_out[97][121],u_xpb_out[98][121],u_xpb_out[99][121],u_xpb_out[100][121],u_xpb_out[101][121],u_xpb_out[102][121],u_xpb_out[103][121],u_xpb_out[104][121],u_xpb_out[105][121]};

assign col_out_122 = {u_xpb_out[0][122],u_xpb_out[1][122],u_xpb_out[2][122],u_xpb_out[3][122],u_xpb_out[4][122],u_xpb_out[5][122],u_xpb_out[6][122],u_xpb_out[7][122],u_xpb_out[8][122],u_xpb_out[9][122],u_xpb_out[10][122],u_xpb_out[11][122],u_xpb_out[12][122],u_xpb_out[13][122],u_xpb_out[14][122],u_xpb_out[15][122],u_xpb_out[16][122],u_xpb_out[17][122],u_xpb_out[18][122],u_xpb_out[19][122],u_xpb_out[20][122],u_xpb_out[21][122],u_xpb_out[22][122],u_xpb_out[23][122],u_xpb_out[24][122],u_xpb_out[25][122],u_xpb_out[26][122],u_xpb_out[27][122],u_xpb_out[28][122],u_xpb_out[29][122],u_xpb_out[30][122],u_xpb_out[31][122],u_xpb_out[32][122],u_xpb_out[33][122],u_xpb_out[34][122],u_xpb_out[35][122],u_xpb_out[36][122],u_xpb_out[37][122],u_xpb_out[38][122],u_xpb_out[39][122],u_xpb_out[40][122],u_xpb_out[41][122],u_xpb_out[42][122],u_xpb_out[43][122],u_xpb_out[44][122],u_xpb_out[45][122],u_xpb_out[46][122],u_xpb_out[47][122],u_xpb_out[48][122],u_xpb_out[49][122],u_xpb_out[50][122],u_xpb_out[51][122],u_xpb_out[52][122],u_xpb_out[53][122],u_xpb_out[54][122],u_xpb_out[55][122],u_xpb_out[56][122],u_xpb_out[57][122],u_xpb_out[58][122],u_xpb_out[59][122],u_xpb_out[60][122],u_xpb_out[61][122],u_xpb_out[62][122],u_xpb_out[63][122],u_xpb_out[64][122],u_xpb_out[65][122],u_xpb_out[66][122],u_xpb_out[67][122],u_xpb_out[68][122],u_xpb_out[69][122],u_xpb_out[70][122],u_xpb_out[71][122],u_xpb_out[72][122],u_xpb_out[73][122],u_xpb_out[74][122],u_xpb_out[75][122],u_xpb_out[76][122],u_xpb_out[77][122],u_xpb_out[78][122],u_xpb_out[79][122],u_xpb_out[80][122],u_xpb_out[81][122],u_xpb_out[82][122],u_xpb_out[83][122],u_xpb_out[84][122],u_xpb_out[85][122],u_xpb_out[86][122],u_xpb_out[87][122],u_xpb_out[88][122],u_xpb_out[89][122],u_xpb_out[90][122],u_xpb_out[91][122],u_xpb_out[92][122],u_xpb_out[93][122],u_xpb_out[94][122],u_xpb_out[95][122],u_xpb_out[96][122],u_xpb_out[97][122],u_xpb_out[98][122],u_xpb_out[99][122],u_xpb_out[100][122],u_xpb_out[101][122],u_xpb_out[102][122],u_xpb_out[103][122],u_xpb_out[104][122],u_xpb_out[105][122]};

assign col_out_123 = {u_xpb_out[0][123],u_xpb_out[1][123],u_xpb_out[2][123],u_xpb_out[3][123],u_xpb_out[4][123],u_xpb_out[5][123],u_xpb_out[6][123],u_xpb_out[7][123],u_xpb_out[8][123],u_xpb_out[9][123],u_xpb_out[10][123],u_xpb_out[11][123],u_xpb_out[12][123],u_xpb_out[13][123],u_xpb_out[14][123],u_xpb_out[15][123],u_xpb_out[16][123],u_xpb_out[17][123],u_xpb_out[18][123],u_xpb_out[19][123],u_xpb_out[20][123],u_xpb_out[21][123],u_xpb_out[22][123],u_xpb_out[23][123],u_xpb_out[24][123],u_xpb_out[25][123],u_xpb_out[26][123],u_xpb_out[27][123],u_xpb_out[28][123],u_xpb_out[29][123],u_xpb_out[30][123],u_xpb_out[31][123],u_xpb_out[32][123],u_xpb_out[33][123],u_xpb_out[34][123],u_xpb_out[35][123],u_xpb_out[36][123],u_xpb_out[37][123],u_xpb_out[38][123],u_xpb_out[39][123],u_xpb_out[40][123],u_xpb_out[41][123],u_xpb_out[42][123],u_xpb_out[43][123],u_xpb_out[44][123],u_xpb_out[45][123],u_xpb_out[46][123],u_xpb_out[47][123],u_xpb_out[48][123],u_xpb_out[49][123],u_xpb_out[50][123],u_xpb_out[51][123],u_xpb_out[52][123],u_xpb_out[53][123],u_xpb_out[54][123],u_xpb_out[55][123],u_xpb_out[56][123],u_xpb_out[57][123],u_xpb_out[58][123],u_xpb_out[59][123],u_xpb_out[60][123],u_xpb_out[61][123],u_xpb_out[62][123],u_xpb_out[63][123],u_xpb_out[64][123],u_xpb_out[65][123],u_xpb_out[66][123],u_xpb_out[67][123],u_xpb_out[68][123],u_xpb_out[69][123],u_xpb_out[70][123],u_xpb_out[71][123],u_xpb_out[72][123],u_xpb_out[73][123],u_xpb_out[74][123],u_xpb_out[75][123],u_xpb_out[76][123],u_xpb_out[77][123],u_xpb_out[78][123],u_xpb_out[79][123],u_xpb_out[80][123],u_xpb_out[81][123],u_xpb_out[82][123],u_xpb_out[83][123],u_xpb_out[84][123],u_xpb_out[85][123],u_xpb_out[86][123],u_xpb_out[87][123],u_xpb_out[88][123],u_xpb_out[89][123],u_xpb_out[90][123],u_xpb_out[91][123],u_xpb_out[92][123],u_xpb_out[93][123],u_xpb_out[94][123],u_xpb_out[95][123],u_xpb_out[96][123],u_xpb_out[97][123],u_xpb_out[98][123],u_xpb_out[99][123],u_xpb_out[100][123],u_xpb_out[101][123],u_xpb_out[102][123],u_xpb_out[103][123],u_xpb_out[104][123],u_xpb_out[105][123]};

assign col_out_124 = {u_xpb_out[0][124],u_xpb_out[1][124],u_xpb_out[2][124],u_xpb_out[3][124],u_xpb_out[4][124],u_xpb_out[5][124],u_xpb_out[6][124],u_xpb_out[7][124],u_xpb_out[8][124],u_xpb_out[9][124],u_xpb_out[10][124],u_xpb_out[11][124],u_xpb_out[12][124],u_xpb_out[13][124],u_xpb_out[14][124],u_xpb_out[15][124],u_xpb_out[16][124],u_xpb_out[17][124],u_xpb_out[18][124],u_xpb_out[19][124],u_xpb_out[20][124],u_xpb_out[21][124],u_xpb_out[22][124],u_xpb_out[23][124],u_xpb_out[24][124],u_xpb_out[25][124],u_xpb_out[26][124],u_xpb_out[27][124],u_xpb_out[28][124],u_xpb_out[29][124],u_xpb_out[30][124],u_xpb_out[31][124],u_xpb_out[32][124],u_xpb_out[33][124],u_xpb_out[34][124],u_xpb_out[35][124],u_xpb_out[36][124],u_xpb_out[37][124],u_xpb_out[38][124],u_xpb_out[39][124],u_xpb_out[40][124],u_xpb_out[41][124],u_xpb_out[42][124],u_xpb_out[43][124],u_xpb_out[44][124],u_xpb_out[45][124],u_xpb_out[46][124],u_xpb_out[47][124],u_xpb_out[48][124],u_xpb_out[49][124],u_xpb_out[50][124],u_xpb_out[51][124],u_xpb_out[52][124],u_xpb_out[53][124],u_xpb_out[54][124],u_xpb_out[55][124],u_xpb_out[56][124],u_xpb_out[57][124],u_xpb_out[58][124],u_xpb_out[59][124],u_xpb_out[60][124],u_xpb_out[61][124],u_xpb_out[62][124],u_xpb_out[63][124],u_xpb_out[64][124],u_xpb_out[65][124],u_xpb_out[66][124],u_xpb_out[67][124],u_xpb_out[68][124],u_xpb_out[69][124],u_xpb_out[70][124],u_xpb_out[71][124],u_xpb_out[72][124],u_xpb_out[73][124],u_xpb_out[74][124],u_xpb_out[75][124],u_xpb_out[76][124],u_xpb_out[77][124],u_xpb_out[78][124],u_xpb_out[79][124],u_xpb_out[80][124],u_xpb_out[81][124],u_xpb_out[82][124],u_xpb_out[83][124],u_xpb_out[84][124],u_xpb_out[85][124],u_xpb_out[86][124],u_xpb_out[87][124],u_xpb_out[88][124],u_xpb_out[89][124],u_xpb_out[90][124],u_xpb_out[91][124],u_xpb_out[92][124],u_xpb_out[93][124],u_xpb_out[94][124],u_xpb_out[95][124],u_xpb_out[96][124],u_xpb_out[97][124],u_xpb_out[98][124],u_xpb_out[99][124],u_xpb_out[100][124],u_xpb_out[101][124],u_xpb_out[102][124],u_xpb_out[103][124],u_xpb_out[104][124],u_xpb_out[105][124]};

assign col_out_125 = {u_xpb_out[0][125],u_xpb_out[1][125],u_xpb_out[2][125],u_xpb_out[3][125],u_xpb_out[4][125],u_xpb_out[5][125],u_xpb_out[6][125],u_xpb_out[7][125],u_xpb_out[8][125],u_xpb_out[9][125],u_xpb_out[10][125],u_xpb_out[11][125],u_xpb_out[12][125],u_xpb_out[13][125],u_xpb_out[14][125],u_xpb_out[15][125],u_xpb_out[16][125],u_xpb_out[17][125],u_xpb_out[18][125],u_xpb_out[19][125],u_xpb_out[20][125],u_xpb_out[21][125],u_xpb_out[22][125],u_xpb_out[23][125],u_xpb_out[24][125],u_xpb_out[25][125],u_xpb_out[26][125],u_xpb_out[27][125],u_xpb_out[28][125],u_xpb_out[29][125],u_xpb_out[30][125],u_xpb_out[31][125],u_xpb_out[32][125],u_xpb_out[33][125],u_xpb_out[34][125],u_xpb_out[35][125],u_xpb_out[36][125],u_xpb_out[37][125],u_xpb_out[38][125],u_xpb_out[39][125],u_xpb_out[40][125],u_xpb_out[41][125],u_xpb_out[42][125],u_xpb_out[43][125],u_xpb_out[44][125],u_xpb_out[45][125],u_xpb_out[46][125],u_xpb_out[47][125],u_xpb_out[48][125],u_xpb_out[49][125],u_xpb_out[50][125],u_xpb_out[51][125],u_xpb_out[52][125],u_xpb_out[53][125],u_xpb_out[54][125],u_xpb_out[55][125],u_xpb_out[56][125],u_xpb_out[57][125],u_xpb_out[58][125],u_xpb_out[59][125],u_xpb_out[60][125],u_xpb_out[61][125],u_xpb_out[62][125],u_xpb_out[63][125],u_xpb_out[64][125],u_xpb_out[65][125],u_xpb_out[66][125],u_xpb_out[67][125],u_xpb_out[68][125],u_xpb_out[69][125],u_xpb_out[70][125],u_xpb_out[71][125],u_xpb_out[72][125],u_xpb_out[73][125],u_xpb_out[74][125],u_xpb_out[75][125],u_xpb_out[76][125],u_xpb_out[77][125],u_xpb_out[78][125],u_xpb_out[79][125],u_xpb_out[80][125],u_xpb_out[81][125],u_xpb_out[82][125],u_xpb_out[83][125],u_xpb_out[84][125],u_xpb_out[85][125],u_xpb_out[86][125],u_xpb_out[87][125],u_xpb_out[88][125],u_xpb_out[89][125],u_xpb_out[90][125],u_xpb_out[91][125],u_xpb_out[92][125],u_xpb_out[93][125],u_xpb_out[94][125],u_xpb_out[95][125],u_xpb_out[96][125],u_xpb_out[97][125],u_xpb_out[98][125],u_xpb_out[99][125],u_xpb_out[100][125],u_xpb_out[101][125],u_xpb_out[102][125],u_xpb_out[103][125],u_xpb_out[104][125],u_xpb_out[105][125]};

assign col_out_126 = {u_xpb_out[0][126],u_xpb_out[1][126],u_xpb_out[2][126],u_xpb_out[3][126],u_xpb_out[4][126],u_xpb_out[5][126],u_xpb_out[6][126],u_xpb_out[7][126],u_xpb_out[8][126],u_xpb_out[9][126],u_xpb_out[10][126],u_xpb_out[11][126],u_xpb_out[12][126],u_xpb_out[13][126],u_xpb_out[14][126],u_xpb_out[15][126],u_xpb_out[16][126],u_xpb_out[17][126],u_xpb_out[18][126],u_xpb_out[19][126],u_xpb_out[20][126],u_xpb_out[21][126],u_xpb_out[22][126],u_xpb_out[23][126],u_xpb_out[24][126],u_xpb_out[25][126],u_xpb_out[26][126],u_xpb_out[27][126],u_xpb_out[28][126],u_xpb_out[29][126],u_xpb_out[30][126],u_xpb_out[31][126],u_xpb_out[32][126],u_xpb_out[33][126],u_xpb_out[34][126],u_xpb_out[35][126],u_xpb_out[36][126],u_xpb_out[37][126],u_xpb_out[38][126],u_xpb_out[39][126],u_xpb_out[40][126],u_xpb_out[41][126],u_xpb_out[42][126],u_xpb_out[43][126],u_xpb_out[44][126],u_xpb_out[45][126],u_xpb_out[46][126],u_xpb_out[47][126],u_xpb_out[48][126],u_xpb_out[49][126],u_xpb_out[50][126],u_xpb_out[51][126],u_xpb_out[52][126],u_xpb_out[53][126],u_xpb_out[54][126],u_xpb_out[55][126],u_xpb_out[56][126],u_xpb_out[57][126],u_xpb_out[58][126],u_xpb_out[59][126],u_xpb_out[60][126],u_xpb_out[61][126],u_xpb_out[62][126],u_xpb_out[63][126],u_xpb_out[64][126],u_xpb_out[65][126],u_xpb_out[66][126],u_xpb_out[67][126],u_xpb_out[68][126],u_xpb_out[69][126],u_xpb_out[70][126],u_xpb_out[71][126],u_xpb_out[72][126],u_xpb_out[73][126],u_xpb_out[74][126],u_xpb_out[75][126],u_xpb_out[76][126],u_xpb_out[77][126],u_xpb_out[78][126],u_xpb_out[79][126],u_xpb_out[80][126],u_xpb_out[81][126],u_xpb_out[82][126],u_xpb_out[83][126],u_xpb_out[84][126],u_xpb_out[85][126],u_xpb_out[86][126],u_xpb_out[87][126],u_xpb_out[88][126],u_xpb_out[89][126],u_xpb_out[90][126],u_xpb_out[91][126],u_xpb_out[92][126],u_xpb_out[93][126],u_xpb_out[94][126],u_xpb_out[95][126],u_xpb_out[96][126],u_xpb_out[97][126],u_xpb_out[98][126],u_xpb_out[99][126],u_xpb_out[100][126],u_xpb_out[101][126],u_xpb_out[102][126],u_xpb_out[103][126],u_xpb_out[104][126],u_xpb_out[105][126]};

assign col_out_127 = {u_xpb_out[0][127],u_xpb_out[1][127],u_xpb_out[2][127],u_xpb_out[3][127],u_xpb_out[4][127],u_xpb_out[5][127],u_xpb_out[6][127],u_xpb_out[7][127],u_xpb_out[8][127],u_xpb_out[9][127],u_xpb_out[10][127],u_xpb_out[11][127],u_xpb_out[12][127],u_xpb_out[13][127],u_xpb_out[14][127],u_xpb_out[15][127],u_xpb_out[16][127],u_xpb_out[17][127],u_xpb_out[18][127],u_xpb_out[19][127],u_xpb_out[20][127],u_xpb_out[21][127],u_xpb_out[22][127],u_xpb_out[23][127],u_xpb_out[24][127],u_xpb_out[25][127],u_xpb_out[26][127],u_xpb_out[27][127],u_xpb_out[28][127],u_xpb_out[29][127],u_xpb_out[30][127],u_xpb_out[31][127],u_xpb_out[32][127],u_xpb_out[33][127],u_xpb_out[34][127],u_xpb_out[35][127],u_xpb_out[36][127],u_xpb_out[37][127],u_xpb_out[38][127],u_xpb_out[39][127],u_xpb_out[40][127],u_xpb_out[41][127],u_xpb_out[42][127],u_xpb_out[43][127],u_xpb_out[44][127],u_xpb_out[45][127],u_xpb_out[46][127],u_xpb_out[47][127],u_xpb_out[48][127],u_xpb_out[49][127],u_xpb_out[50][127],u_xpb_out[51][127],u_xpb_out[52][127],u_xpb_out[53][127],u_xpb_out[54][127],u_xpb_out[55][127],u_xpb_out[56][127],u_xpb_out[57][127],u_xpb_out[58][127],u_xpb_out[59][127],u_xpb_out[60][127],u_xpb_out[61][127],u_xpb_out[62][127],u_xpb_out[63][127],u_xpb_out[64][127],u_xpb_out[65][127],u_xpb_out[66][127],u_xpb_out[67][127],u_xpb_out[68][127],u_xpb_out[69][127],u_xpb_out[70][127],u_xpb_out[71][127],u_xpb_out[72][127],u_xpb_out[73][127],u_xpb_out[74][127],u_xpb_out[75][127],u_xpb_out[76][127],u_xpb_out[77][127],u_xpb_out[78][127],u_xpb_out[79][127],u_xpb_out[80][127],u_xpb_out[81][127],u_xpb_out[82][127],u_xpb_out[83][127],u_xpb_out[84][127],u_xpb_out[85][127],u_xpb_out[86][127],u_xpb_out[87][127],u_xpb_out[88][127],u_xpb_out[89][127],u_xpb_out[90][127],u_xpb_out[91][127],u_xpb_out[92][127],u_xpb_out[93][127],u_xpb_out[94][127],u_xpb_out[95][127],u_xpb_out[96][127],u_xpb_out[97][127],u_xpb_out[98][127],u_xpb_out[99][127],u_xpb_out[100][127],u_xpb_out[101][127],u_xpb_out[102][127],u_xpb_out[103][127],u_xpb_out[104][127],u_xpb_out[105][127]};

assign col_out_128 = {u_xpb_out[0][128],u_xpb_out[1][128],u_xpb_out[2][128],u_xpb_out[3][128],u_xpb_out[4][128],u_xpb_out[5][128],u_xpb_out[6][128],u_xpb_out[7][128],u_xpb_out[8][128],u_xpb_out[9][128],u_xpb_out[10][128],u_xpb_out[11][128],u_xpb_out[12][128],u_xpb_out[13][128],u_xpb_out[14][128],u_xpb_out[15][128],u_xpb_out[16][128],u_xpb_out[17][128],u_xpb_out[18][128],u_xpb_out[19][128],u_xpb_out[20][128],u_xpb_out[21][128],u_xpb_out[22][128],u_xpb_out[23][128],u_xpb_out[24][128],u_xpb_out[25][128],u_xpb_out[26][128],u_xpb_out[27][128],u_xpb_out[28][128],u_xpb_out[29][128],u_xpb_out[30][128],u_xpb_out[31][128],u_xpb_out[32][128],u_xpb_out[33][128],u_xpb_out[34][128],u_xpb_out[35][128],u_xpb_out[36][128],u_xpb_out[37][128],u_xpb_out[38][128],u_xpb_out[39][128],u_xpb_out[40][128],u_xpb_out[41][128],u_xpb_out[42][128],u_xpb_out[43][128],u_xpb_out[44][128],u_xpb_out[45][128],u_xpb_out[46][128],u_xpb_out[47][128],u_xpb_out[48][128],u_xpb_out[49][128],u_xpb_out[50][128],u_xpb_out[51][128],u_xpb_out[52][128],u_xpb_out[53][128],u_xpb_out[54][128],u_xpb_out[55][128],u_xpb_out[56][128],u_xpb_out[57][128],u_xpb_out[58][128],u_xpb_out[59][128],u_xpb_out[60][128],u_xpb_out[61][128],u_xpb_out[62][128],u_xpb_out[63][128],u_xpb_out[64][128],u_xpb_out[65][128],u_xpb_out[66][128],u_xpb_out[67][128],u_xpb_out[68][128],u_xpb_out[69][128],u_xpb_out[70][128],u_xpb_out[71][128],u_xpb_out[72][128],u_xpb_out[73][128],u_xpb_out[74][128],u_xpb_out[75][128],u_xpb_out[76][128],u_xpb_out[77][128],u_xpb_out[78][128],u_xpb_out[79][128],u_xpb_out[80][128],u_xpb_out[81][128],u_xpb_out[82][128],u_xpb_out[83][128],u_xpb_out[84][128],u_xpb_out[85][128],u_xpb_out[86][128],u_xpb_out[87][128],u_xpb_out[88][128],u_xpb_out[89][128],u_xpb_out[90][128],u_xpb_out[91][128],u_xpb_out[92][128],u_xpb_out[93][128],u_xpb_out[94][128],u_xpb_out[95][128],u_xpb_out[96][128],u_xpb_out[97][128],u_xpb_out[98][128],u_xpb_out[99][128],u_xpb_out[100][128],u_xpb_out[101][128],u_xpb_out[102][128],u_xpb_out[103][128],u_xpb_out[104][128],u_xpb_out[105][128]};

assign col_out_129 = {u_xpb_out[0][129],u_xpb_out[1][129],u_xpb_out[2][129],u_xpb_out[3][129],u_xpb_out[4][129],u_xpb_out[5][129],u_xpb_out[6][129],u_xpb_out[7][129],u_xpb_out[8][129],u_xpb_out[9][129],u_xpb_out[10][129],u_xpb_out[11][129],u_xpb_out[12][129],u_xpb_out[13][129],u_xpb_out[14][129],u_xpb_out[15][129],u_xpb_out[16][129],u_xpb_out[17][129],u_xpb_out[18][129],u_xpb_out[19][129],u_xpb_out[20][129],u_xpb_out[21][129],u_xpb_out[22][129],u_xpb_out[23][129],u_xpb_out[24][129],u_xpb_out[25][129],u_xpb_out[26][129],u_xpb_out[27][129],u_xpb_out[28][129],u_xpb_out[29][129],u_xpb_out[30][129],u_xpb_out[31][129],u_xpb_out[32][129],u_xpb_out[33][129],u_xpb_out[34][129],u_xpb_out[35][129],u_xpb_out[36][129],u_xpb_out[37][129],u_xpb_out[38][129],u_xpb_out[39][129],u_xpb_out[40][129],u_xpb_out[41][129],u_xpb_out[42][129],u_xpb_out[43][129],u_xpb_out[44][129],u_xpb_out[45][129],u_xpb_out[46][129],u_xpb_out[47][129],u_xpb_out[48][129],u_xpb_out[49][129],u_xpb_out[50][129],u_xpb_out[51][129],u_xpb_out[52][129],u_xpb_out[53][129],u_xpb_out[54][129],u_xpb_out[55][129],u_xpb_out[56][129],u_xpb_out[57][129],u_xpb_out[58][129],u_xpb_out[59][129],u_xpb_out[60][129],u_xpb_out[61][129],u_xpb_out[62][129],u_xpb_out[63][129],u_xpb_out[64][129],u_xpb_out[65][129],u_xpb_out[66][129],u_xpb_out[67][129],u_xpb_out[68][129],u_xpb_out[69][129],u_xpb_out[70][129],u_xpb_out[71][129],u_xpb_out[72][129],u_xpb_out[73][129],u_xpb_out[74][129],u_xpb_out[75][129],u_xpb_out[76][129],u_xpb_out[77][129],u_xpb_out[78][129],u_xpb_out[79][129],u_xpb_out[80][129],u_xpb_out[81][129],u_xpb_out[82][129],u_xpb_out[83][129],u_xpb_out[84][129],u_xpb_out[85][129],u_xpb_out[86][129],u_xpb_out[87][129],u_xpb_out[88][129],u_xpb_out[89][129],u_xpb_out[90][129],u_xpb_out[91][129],u_xpb_out[92][129],u_xpb_out[93][129],u_xpb_out[94][129],u_xpb_out[95][129],u_xpb_out[96][129],u_xpb_out[97][129],u_xpb_out[98][129],u_xpb_out[99][129],u_xpb_out[100][129],u_xpb_out[101][129],u_xpb_out[102][129],u_xpb_out[103][129],u_xpb_out[104][129],u_xpb_out[105][129]};

assign col_out_130 = {u_xpb_out[0][130],u_xpb_out[1][130],u_xpb_out[2][130],u_xpb_out[3][130],u_xpb_out[4][130],u_xpb_out[5][130],u_xpb_out[6][130],u_xpb_out[7][130],u_xpb_out[8][130],u_xpb_out[9][130],u_xpb_out[10][130],u_xpb_out[11][130],u_xpb_out[12][130],u_xpb_out[13][130],u_xpb_out[14][130],u_xpb_out[15][130],u_xpb_out[16][130],u_xpb_out[17][130],u_xpb_out[18][130],u_xpb_out[19][130],u_xpb_out[20][130],u_xpb_out[21][130],u_xpb_out[22][130],u_xpb_out[23][130],u_xpb_out[24][130],u_xpb_out[25][130],u_xpb_out[26][130],u_xpb_out[27][130],u_xpb_out[28][130],u_xpb_out[29][130],u_xpb_out[30][130],u_xpb_out[31][130],u_xpb_out[32][130],u_xpb_out[33][130],u_xpb_out[34][130],u_xpb_out[35][130],u_xpb_out[36][130],u_xpb_out[37][130],u_xpb_out[38][130],u_xpb_out[39][130],u_xpb_out[40][130],u_xpb_out[41][130],u_xpb_out[42][130],u_xpb_out[43][130],u_xpb_out[44][130],u_xpb_out[45][130],u_xpb_out[46][130],u_xpb_out[47][130],u_xpb_out[48][130],u_xpb_out[49][130],u_xpb_out[50][130],u_xpb_out[51][130],u_xpb_out[52][130],u_xpb_out[53][130],u_xpb_out[54][130],u_xpb_out[55][130],u_xpb_out[56][130],u_xpb_out[57][130],u_xpb_out[58][130],u_xpb_out[59][130],u_xpb_out[60][130],u_xpb_out[61][130],u_xpb_out[62][130],u_xpb_out[63][130],u_xpb_out[64][130],u_xpb_out[65][130],u_xpb_out[66][130],u_xpb_out[67][130],u_xpb_out[68][130],u_xpb_out[69][130],u_xpb_out[70][130],u_xpb_out[71][130],u_xpb_out[72][130],u_xpb_out[73][130],u_xpb_out[74][130],u_xpb_out[75][130],u_xpb_out[76][130],u_xpb_out[77][130],u_xpb_out[78][130],u_xpb_out[79][130],u_xpb_out[80][130],u_xpb_out[81][130],u_xpb_out[82][130],u_xpb_out[83][130],u_xpb_out[84][130],u_xpb_out[85][130],u_xpb_out[86][130],u_xpb_out[87][130],u_xpb_out[88][130],u_xpb_out[89][130],u_xpb_out[90][130],u_xpb_out[91][130],u_xpb_out[92][130],u_xpb_out[93][130],u_xpb_out[94][130],u_xpb_out[95][130],u_xpb_out[96][130],u_xpb_out[97][130],u_xpb_out[98][130],u_xpb_out[99][130],u_xpb_out[100][130],u_xpb_out[101][130],u_xpb_out[102][130],u_xpb_out[103][130],u_xpb_out[104][130],u_xpb_out[105][130]};

assign col_out_131 = {u_xpb_out[0][131],u_xpb_out[1][131],u_xpb_out[2][131],u_xpb_out[3][131],u_xpb_out[4][131],u_xpb_out[5][131],u_xpb_out[6][131],u_xpb_out[7][131],u_xpb_out[8][131],u_xpb_out[9][131],u_xpb_out[10][131],u_xpb_out[11][131],u_xpb_out[12][131],u_xpb_out[13][131],u_xpb_out[14][131],u_xpb_out[15][131],u_xpb_out[16][131],u_xpb_out[17][131],u_xpb_out[18][131],u_xpb_out[19][131],u_xpb_out[20][131],u_xpb_out[21][131],u_xpb_out[22][131],u_xpb_out[23][131],u_xpb_out[24][131],u_xpb_out[25][131],u_xpb_out[26][131],u_xpb_out[27][131],u_xpb_out[28][131],u_xpb_out[29][131],u_xpb_out[30][131],u_xpb_out[31][131],u_xpb_out[32][131],u_xpb_out[33][131],u_xpb_out[34][131],u_xpb_out[35][131],u_xpb_out[36][131],u_xpb_out[37][131],u_xpb_out[38][131],u_xpb_out[39][131],u_xpb_out[40][131],u_xpb_out[41][131],u_xpb_out[42][131],u_xpb_out[43][131],u_xpb_out[44][131],u_xpb_out[45][131],u_xpb_out[46][131],u_xpb_out[47][131],u_xpb_out[48][131],u_xpb_out[49][131],u_xpb_out[50][131],u_xpb_out[51][131],u_xpb_out[52][131],u_xpb_out[53][131],u_xpb_out[54][131],u_xpb_out[55][131],u_xpb_out[56][131],u_xpb_out[57][131],u_xpb_out[58][131],u_xpb_out[59][131],u_xpb_out[60][131],u_xpb_out[61][131],u_xpb_out[62][131],u_xpb_out[63][131],u_xpb_out[64][131],u_xpb_out[65][131],u_xpb_out[66][131],u_xpb_out[67][131],u_xpb_out[68][131],u_xpb_out[69][131],u_xpb_out[70][131],u_xpb_out[71][131],u_xpb_out[72][131],u_xpb_out[73][131],u_xpb_out[74][131],u_xpb_out[75][131],u_xpb_out[76][131],u_xpb_out[77][131],u_xpb_out[78][131],u_xpb_out[79][131],u_xpb_out[80][131],u_xpb_out[81][131],u_xpb_out[82][131],u_xpb_out[83][131],u_xpb_out[84][131],u_xpb_out[85][131],u_xpb_out[86][131],u_xpb_out[87][131],u_xpb_out[88][131],u_xpb_out[89][131],u_xpb_out[90][131],u_xpb_out[91][131],u_xpb_out[92][131],u_xpb_out[93][131],u_xpb_out[94][131],u_xpb_out[95][131],u_xpb_out[96][131],u_xpb_out[97][131],u_xpb_out[98][131],u_xpb_out[99][131],u_xpb_out[100][131],u_xpb_out[101][131],u_xpb_out[102][131],u_xpb_out[103][131],u_xpb_out[104][131],u_xpb_out[105][131]};

assign col_out_132 = {u_xpb_out[0][132],u_xpb_out[1][132],u_xpb_out[2][132],u_xpb_out[3][132],u_xpb_out[4][132],u_xpb_out[5][132],u_xpb_out[6][132],u_xpb_out[7][132],u_xpb_out[8][132],u_xpb_out[9][132],u_xpb_out[10][132],u_xpb_out[11][132],u_xpb_out[12][132],u_xpb_out[13][132],u_xpb_out[14][132],u_xpb_out[15][132],u_xpb_out[16][132],u_xpb_out[17][132],u_xpb_out[18][132],u_xpb_out[19][132],u_xpb_out[20][132],u_xpb_out[21][132],u_xpb_out[22][132],u_xpb_out[23][132],u_xpb_out[24][132],u_xpb_out[25][132],u_xpb_out[26][132],u_xpb_out[27][132],u_xpb_out[28][132],u_xpb_out[29][132],u_xpb_out[30][132],u_xpb_out[31][132],u_xpb_out[32][132],u_xpb_out[33][132],u_xpb_out[34][132],u_xpb_out[35][132],u_xpb_out[36][132],u_xpb_out[37][132],u_xpb_out[38][132],u_xpb_out[39][132],u_xpb_out[40][132],u_xpb_out[41][132],u_xpb_out[42][132],u_xpb_out[43][132],u_xpb_out[44][132],u_xpb_out[45][132],u_xpb_out[46][132],u_xpb_out[47][132],u_xpb_out[48][132],u_xpb_out[49][132],u_xpb_out[50][132],u_xpb_out[51][132],u_xpb_out[52][132],u_xpb_out[53][132],u_xpb_out[54][132],u_xpb_out[55][132],u_xpb_out[56][132],u_xpb_out[57][132],u_xpb_out[58][132],u_xpb_out[59][132],u_xpb_out[60][132],u_xpb_out[61][132],u_xpb_out[62][132],u_xpb_out[63][132],u_xpb_out[64][132],u_xpb_out[65][132],u_xpb_out[66][132],u_xpb_out[67][132],u_xpb_out[68][132],u_xpb_out[69][132],u_xpb_out[70][132],u_xpb_out[71][132],u_xpb_out[72][132],u_xpb_out[73][132],u_xpb_out[74][132],u_xpb_out[75][132],u_xpb_out[76][132],u_xpb_out[77][132],u_xpb_out[78][132],u_xpb_out[79][132],u_xpb_out[80][132],u_xpb_out[81][132],u_xpb_out[82][132],u_xpb_out[83][132],u_xpb_out[84][132],u_xpb_out[85][132],u_xpb_out[86][132],u_xpb_out[87][132],u_xpb_out[88][132],u_xpb_out[89][132],u_xpb_out[90][132],u_xpb_out[91][132],u_xpb_out[92][132],u_xpb_out[93][132],u_xpb_out[94][132],u_xpb_out[95][132],u_xpb_out[96][132],u_xpb_out[97][132],u_xpb_out[98][132],u_xpb_out[99][132],u_xpb_out[100][132],u_xpb_out[101][132],u_xpb_out[102][132],u_xpb_out[103][132],u_xpb_out[104][132],u_xpb_out[105][132]};

assign col_out_133 = {u_xpb_out[0][133],u_xpb_out[1][133],u_xpb_out[2][133],u_xpb_out[3][133],u_xpb_out[4][133],u_xpb_out[5][133],u_xpb_out[6][133],u_xpb_out[7][133],u_xpb_out[8][133],u_xpb_out[9][133],u_xpb_out[10][133],u_xpb_out[11][133],u_xpb_out[12][133],u_xpb_out[13][133],u_xpb_out[14][133],u_xpb_out[15][133],u_xpb_out[16][133],u_xpb_out[17][133],u_xpb_out[18][133],u_xpb_out[19][133],u_xpb_out[20][133],u_xpb_out[21][133],u_xpb_out[22][133],u_xpb_out[23][133],u_xpb_out[24][133],u_xpb_out[25][133],u_xpb_out[26][133],u_xpb_out[27][133],u_xpb_out[28][133],u_xpb_out[29][133],u_xpb_out[30][133],u_xpb_out[31][133],u_xpb_out[32][133],u_xpb_out[33][133],u_xpb_out[34][133],u_xpb_out[35][133],u_xpb_out[36][133],u_xpb_out[37][133],u_xpb_out[38][133],u_xpb_out[39][133],u_xpb_out[40][133],u_xpb_out[41][133],u_xpb_out[42][133],u_xpb_out[43][133],u_xpb_out[44][133],u_xpb_out[45][133],u_xpb_out[46][133],u_xpb_out[47][133],u_xpb_out[48][133],u_xpb_out[49][133],u_xpb_out[50][133],u_xpb_out[51][133],u_xpb_out[52][133],u_xpb_out[53][133],u_xpb_out[54][133],u_xpb_out[55][133],u_xpb_out[56][133],u_xpb_out[57][133],u_xpb_out[58][133],u_xpb_out[59][133],u_xpb_out[60][133],u_xpb_out[61][133],u_xpb_out[62][133],u_xpb_out[63][133],u_xpb_out[64][133],u_xpb_out[65][133],u_xpb_out[66][133],u_xpb_out[67][133],u_xpb_out[68][133],u_xpb_out[69][133],u_xpb_out[70][133],u_xpb_out[71][133],u_xpb_out[72][133],u_xpb_out[73][133],u_xpb_out[74][133],u_xpb_out[75][133],u_xpb_out[76][133],u_xpb_out[77][133],u_xpb_out[78][133],u_xpb_out[79][133],u_xpb_out[80][133],u_xpb_out[81][133],u_xpb_out[82][133],u_xpb_out[83][133],u_xpb_out[84][133],u_xpb_out[85][133],u_xpb_out[86][133],u_xpb_out[87][133],u_xpb_out[88][133],u_xpb_out[89][133],u_xpb_out[90][133],u_xpb_out[91][133],u_xpb_out[92][133],u_xpb_out[93][133],u_xpb_out[94][133],u_xpb_out[95][133],u_xpb_out[96][133],u_xpb_out[97][133],u_xpb_out[98][133],u_xpb_out[99][133],u_xpb_out[100][133],u_xpb_out[101][133],u_xpb_out[102][133],u_xpb_out[103][133],u_xpb_out[104][133],u_xpb_out[105][133]};

assign col_out_134 = {u_xpb_out[0][134],u_xpb_out[1][134],u_xpb_out[2][134],u_xpb_out[3][134],u_xpb_out[4][134],u_xpb_out[5][134],u_xpb_out[6][134],u_xpb_out[7][134],u_xpb_out[8][134],u_xpb_out[9][134],u_xpb_out[10][134],u_xpb_out[11][134],u_xpb_out[12][134],u_xpb_out[13][134],u_xpb_out[14][134],u_xpb_out[15][134],u_xpb_out[16][134],u_xpb_out[17][134],u_xpb_out[18][134],u_xpb_out[19][134],u_xpb_out[20][134],u_xpb_out[21][134],u_xpb_out[22][134],u_xpb_out[23][134],u_xpb_out[24][134],u_xpb_out[25][134],u_xpb_out[26][134],u_xpb_out[27][134],u_xpb_out[28][134],u_xpb_out[29][134],u_xpb_out[30][134],u_xpb_out[31][134],u_xpb_out[32][134],u_xpb_out[33][134],u_xpb_out[34][134],u_xpb_out[35][134],u_xpb_out[36][134],u_xpb_out[37][134],u_xpb_out[38][134],u_xpb_out[39][134],u_xpb_out[40][134],u_xpb_out[41][134],u_xpb_out[42][134],u_xpb_out[43][134],u_xpb_out[44][134],u_xpb_out[45][134],u_xpb_out[46][134],u_xpb_out[47][134],u_xpb_out[48][134],u_xpb_out[49][134],u_xpb_out[50][134],u_xpb_out[51][134],u_xpb_out[52][134],u_xpb_out[53][134],u_xpb_out[54][134],u_xpb_out[55][134],u_xpb_out[56][134],u_xpb_out[57][134],u_xpb_out[58][134],u_xpb_out[59][134],u_xpb_out[60][134],u_xpb_out[61][134],u_xpb_out[62][134],u_xpb_out[63][134],u_xpb_out[64][134],u_xpb_out[65][134],u_xpb_out[66][134],u_xpb_out[67][134],u_xpb_out[68][134],u_xpb_out[69][134],u_xpb_out[70][134],u_xpb_out[71][134],u_xpb_out[72][134],u_xpb_out[73][134],u_xpb_out[74][134],u_xpb_out[75][134],u_xpb_out[76][134],u_xpb_out[77][134],u_xpb_out[78][134],u_xpb_out[79][134],u_xpb_out[80][134],u_xpb_out[81][134],u_xpb_out[82][134],u_xpb_out[83][134],u_xpb_out[84][134],u_xpb_out[85][134],u_xpb_out[86][134],u_xpb_out[87][134],u_xpb_out[88][134],u_xpb_out[89][134],u_xpb_out[90][134],u_xpb_out[91][134],u_xpb_out[92][134],u_xpb_out[93][134],u_xpb_out[94][134],u_xpb_out[95][134],u_xpb_out[96][134],u_xpb_out[97][134],u_xpb_out[98][134],u_xpb_out[99][134],u_xpb_out[100][134],u_xpb_out[101][134],u_xpb_out[102][134],u_xpb_out[103][134],u_xpb_out[104][134],u_xpb_out[105][134]};

assign col_out_135 = {u_xpb_out[0][135],u_xpb_out[1][135],u_xpb_out[2][135],u_xpb_out[3][135],u_xpb_out[4][135],u_xpb_out[5][135],u_xpb_out[6][135],u_xpb_out[7][135],u_xpb_out[8][135],u_xpb_out[9][135],u_xpb_out[10][135],u_xpb_out[11][135],u_xpb_out[12][135],u_xpb_out[13][135],u_xpb_out[14][135],u_xpb_out[15][135],u_xpb_out[16][135],u_xpb_out[17][135],u_xpb_out[18][135],u_xpb_out[19][135],u_xpb_out[20][135],u_xpb_out[21][135],u_xpb_out[22][135],u_xpb_out[23][135],u_xpb_out[24][135],u_xpb_out[25][135],u_xpb_out[26][135],u_xpb_out[27][135],u_xpb_out[28][135],u_xpb_out[29][135],u_xpb_out[30][135],u_xpb_out[31][135],u_xpb_out[32][135],u_xpb_out[33][135],u_xpb_out[34][135],u_xpb_out[35][135],u_xpb_out[36][135],u_xpb_out[37][135],u_xpb_out[38][135],u_xpb_out[39][135],u_xpb_out[40][135],u_xpb_out[41][135],u_xpb_out[42][135],u_xpb_out[43][135],u_xpb_out[44][135],u_xpb_out[45][135],u_xpb_out[46][135],u_xpb_out[47][135],u_xpb_out[48][135],u_xpb_out[49][135],u_xpb_out[50][135],u_xpb_out[51][135],u_xpb_out[52][135],u_xpb_out[53][135],u_xpb_out[54][135],u_xpb_out[55][135],u_xpb_out[56][135],u_xpb_out[57][135],u_xpb_out[58][135],u_xpb_out[59][135],u_xpb_out[60][135],u_xpb_out[61][135],u_xpb_out[62][135],u_xpb_out[63][135],u_xpb_out[64][135],u_xpb_out[65][135],u_xpb_out[66][135],u_xpb_out[67][135],u_xpb_out[68][135],u_xpb_out[69][135],u_xpb_out[70][135],u_xpb_out[71][135],u_xpb_out[72][135],u_xpb_out[73][135],u_xpb_out[74][135],u_xpb_out[75][135],u_xpb_out[76][135],u_xpb_out[77][135],u_xpb_out[78][135],u_xpb_out[79][135],u_xpb_out[80][135],u_xpb_out[81][135],u_xpb_out[82][135],u_xpb_out[83][135],u_xpb_out[84][135],u_xpb_out[85][135],u_xpb_out[86][135],u_xpb_out[87][135],u_xpb_out[88][135],u_xpb_out[89][135],u_xpb_out[90][135],u_xpb_out[91][135],u_xpb_out[92][135],u_xpb_out[93][135],u_xpb_out[94][135],u_xpb_out[95][135],u_xpb_out[96][135],u_xpb_out[97][135],u_xpb_out[98][135],u_xpb_out[99][135],u_xpb_out[100][135],u_xpb_out[101][135],u_xpb_out[102][135],u_xpb_out[103][135],u_xpb_out[104][135],u_xpb_out[105][135]};

assign col_out_136 = {u_xpb_out[0][136],u_xpb_out[1][136],u_xpb_out[2][136],u_xpb_out[3][136],u_xpb_out[4][136],u_xpb_out[5][136],u_xpb_out[6][136],u_xpb_out[7][136],u_xpb_out[8][136],u_xpb_out[9][136],u_xpb_out[10][136],u_xpb_out[11][136],u_xpb_out[12][136],u_xpb_out[13][136],u_xpb_out[14][136],u_xpb_out[15][136],u_xpb_out[16][136],u_xpb_out[17][136],u_xpb_out[18][136],u_xpb_out[19][136],u_xpb_out[20][136],u_xpb_out[21][136],u_xpb_out[22][136],u_xpb_out[23][136],u_xpb_out[24][136],u_xpb_out[25][136],u_xpb_out[26][136],u_xpb_out[27][136],u_xpb_out[28][136],u_xpb_out[29][136],u_xpb_out[30][136],u_xpb_out[31][136],u_xpb_out[32][136],u_xpb_out[33][136],u_xpb_out[34][136],u_xpb_out[35][136],u_xpb_out[36][136],u_xpb_out[37][136],u_xpb_out[38][136],u_xpb_out[39][136],u_xpb_out[40][136],u_xpb_out[41][136],u_xpb_out[42][136],u_xpb_out[43][136],u_xpb_out[44][136],u_xpb_out[45][136],u_xpb_out[46][136],u_xpb_out[47][136],u_xpb_out[48][136],u_xpb_out[49][136],u_xpb_out[50][136],u_xpb_out[51][136],u_xpb_out[52][136],u_xpb_out[53][136],u_xpb_out[54][136],u_xpb_out[55][136],u_xpb_out[56][136],u_xpb_out[57][136],u_xpb_out[58][136],u_xpb_out[59][136],u_xpb_out[60][136],u_xpb_out[61][136],u_xpb_out[62][136],u_xpb_out[63][136],u_xpb_out[64][136],u_xpb_out[65][136],u_xpb_out[66][136],u_xpb_out[67][136],u_xpb_out[68][136],u_xpb_out[69][136],u_xpb_out[70][136],u_xpb_out[71][136],u_xpb_out[72][136],u_xpb_out[73][136],u_xpb_out[74][136],u_xpb_out[75][136],u_xpb_out[76][136],u_xpb_out[77][136],u_xpb_out[78][136],u_xpb_out[79][136],u_xpb_out[80][136],u_xpb_out[81][136],u_xpb_out[82][136],u_xpb_out[83][136],u_xpb_out[84][136],u_xpb_out[85][136],u_xpb_out[86][136],u_xpb_out[87][136],u_xpb_out[88][136],u_xpb_out[89][136],u_xpb_out[90][136],u_xpb_out[91][136],u_xpb_out[92][136],u_xpb_out[93][136],u_xpb_out[94][136],u_xpb_out[95][136],u_xpb_out[96][136],u_xpb_out[97][136],u_xpb_out[98][136],u_xpb_out[99][136],u_xpb_out[100][136],u_xpb_out[101][136],u_xpb_out[102][136],u_xpb_out[103][136],u_xpb_out[104][136],u_xpb_out[105][136]};

assign col_out_137 = {u_xpb_out[0][137],u_xpb_out[1][137],u_xpb_out[2][137],u_xpb_out[3][137],u_xpb_out[4][137],u_xpb_out[5][137],u_xpb_out[6][137],u_xpb_out[7][137],u_xpb_out[8][137],u_xpb_out[9][137],u_xpb_out[10][137],u_xpb_out[11][137],u_xpb_out[12][137],u_xpb_out[13][137],u_xpb_out[14][137],u_xpb_out[15][137],u_xpb_out[16][137],u_xpb_out[17][137],u_xpb_out[18][137],u_xpb_out[19][137],u_xpb_out[20][137],u_xpb_out[21][137],u_xpb_out[22][137],u_xpb_out[23][137],u_xpb_out[24][137],u_xpb_out[25][137],u_xpb_out[26][137],u_xpb_out[27][137],u_xpb_out[28][137],u_xpb_out[29][137],u_xpb_out[30][137],u_xpb_out[31][137],u_xpb_out[32][137],u_xpb_out[33][137],u_xpb_out[34][137],u_xpb_out[35][137],u_xpb_out[36][137],u_xpb_out[37][137],u_xpb_out[38][137],u_xpb_out[39][137],u_xpb_out[40][137],u_xpb_out[41][137],u_xpb_out[42][137],u_xpb_out[43][137],u_xpb_out[44][137],u_xpb_out[45][137],u_xpb_out[46][137],u_xpb_out[47][137],u_xpb_out[48][137],u_xpb_out[49][137],u_xpb_out[50][137],u_xpb_out[51][137],u_xpb_out[52][137],u_xpb_out[53][137],u_xpb_out[54][137],u_xpb_out[55][137],u_xpb_out[56][137],u_xpb_out[57][137],u_xpb_out[58][137],u_xpb_out[59][137],u_xpb_out[60][137],u_xpb_out[61][137],u_xpb_out[62][137],u_xpb_out[63][137],u_xpb_out[64][137],u_xpb_out[65][137],u_xpb_out[66][137],u_xpb_out[67][137],u_xpb_out[68][137],u_xpb_out[69][137],u_xpb_out[70][137],u_xpb_out[71][137],u_xpb_out[72][137],u_xpb_out[73][137],u_xpb_out[74][137],u_xpb_out[75][137],u_xpb_out[76][137],u_xpb_out[77][137],u_xpb_out[78][137],u_xpb_out[79][137],u_xpb_out[80][137],u_xpb_out[81][137],u_xpb_out[82][137],u_xpb_out[83][137],u_xpb_out[84][137],u_xpb_out[85][137],u_xpb_out[86][137],u_xpb_out[87][137],u_xpb_out[88][137],u_xpb_out[89][137],u_xpb_out[90][137],u_xpb_out[91][137],u_xpb_out[92][137],u_xpb_out[93][137],u_xpb_out[94][137],u_xpb_out[95][137],u_xpb_out[96][137],u_xpb_out[97][137],u_xpb_out[98][137],u_xpb_out[99][137],u_xpb_out[100][137],u_xpb_out[101][137],u_xpb_out[102][137],u_xpb_out[103][137],u_xpb_out[104][137],u_xpb_out[105][137]};

assign col_out_138 = {u_xpb_out[0][138],u_xpb_out[1][138],u_xpb_out[2][138],u_xpb_out[3][138],u_xpb_out[4][138],u_xpb_out[5][138],u_xpb_out[6][138],u_xpb_out[7][138],u_xpb_out[8][138],u_xpb_out[9][138],u_xpb_out[10][138],u_xpb_out[11][138],u_xpb_out[12][138],u_xpb_out[13][138],u_xpb_out[14][138],u_xpb_out[15][138],u_xpb_out[16][138],u_xpb_out[17][138],u_xpb_out[18][138],u_xpb_out[19][138],u_xpb_out[20][138],u_xpb_out[21][138],u_xpb_out[22][138],u_xpb_out[23][138],u_xpb_out[24][138],u_xpb_out[25][138],u_xpb_out[26][138],u_xpb_out[27][138],u_xpb_out[28][138],u_xpb_out[29][138],u_xpb_out[30][138],u_xpb_out[31][138],u_xpb_out[32][138],u_xpb_out[33][138],u_xpb_out[34][138],u_xpb_out[35][138],u_xpb_out[36][138],u_xpb_out[37][138],u_xpb_out[38][138],u_xpb_out[39][138],u_xpb_out[40][138],u_xpb_out[41][138],u_xpb_out[42][138],u_xpb_out[43][138],u_xpb_out[44][138],u_xpb_out[45][138],u_xpb_out[46][138],u_xpb_out[47][138],u_xpb_out[48][138],u_xpb_out[49][138],u_xpb_out[50][138],u_xpb_out[51][138],u_xpb_out[52][138],u_xpb_out[53][138],u_xpb_out[54][138],u_xpb_out[55][138],u_xpb_out[56][138],u_xpb_out[57][138],u_xpb_out[58][138],u_xpb_out[59][138],u_xpb_out[60][138],u_xpb_out[61][138],u_xpb_out[62][138],u_xpb_out[63][138],u_xpb_out[64][138],u_xpb_out[65][138],u_xpb_out[66][138],u_xpb_out[67][138],u_xpb_out[68][138],u_xpb_out[69][138],u_xpb_out[70][138],u_xpb_out[71][138],u_xpb_out[72][138],u_xpb_out[73][138],u_xpb_out[74][138],u_xpb_out[75][138],u_xpb_out[76][138],u_xpb_out[77][138],u_xpb_out[78][138],u_xpb_out[79][138],u_xpb_out[80][138],u_xpb_out[81][138],u_xpb_out[82][138],u_xpb_out[83][138],u_xpb_out[84][138],u_xpb_out[85][138],u_xpb_out[86][138],u_xpb_out[87][138],u_xpb_out[88][138],u_xpb_out[89][138],u_xpb_out[90][138],u_xpb_out[91][138],u_xpb_out[92][138],u_xpb_out[93][138],u_xpb_out[94][138],u_xpb_out[95][138],u_xpb_out[96][138],u_xpb_out[97][138],u_xpb_out[98][138],u_xpb_out[99][138],u_xpb_out[100][138],u_xpb_out[101][138],u_xpb_out[102][138],u_xpb_out[103][138],u_xpb_out[104][138],u_xpb_out[105][138]};

assign col_out_139 = {u_xpb_out[0][139],u_xpb_out[1][139],u_xpb_out[2][139],u_xpb_out[3][139],u_xpb_out[4][139],u_xpb_out[5][139],u_xpb_out[6][139],u_xpb_out[7][139],u_xpb_out[8][139],u_xpb_out[9][139],u_xpb_out[10][139],u_xpb_out[11][139],u_xpb_out[12][139],u_xpb_out[13][139],u_xpb_out[14][139],u_xpb_out[15][139],u_xpb_out[16][139],u_xpb_out[17][139],u_xpb_out[18][139],u_xpb_out[19][139],u_xpb_out[20][139],u_xpb_out[21][139],u_xpb_out[22][139],u_xpb_out[23][139],u_xpb_out[24][139],u_xpb_out[25][139],u_xpb_out[26][139],u_xpb_out[27][139],u_xpb_out[28][139],u_xpb_out[29][139],u_xpb_out[30][139],u_xpb_out[31][139],u_xpb_out[32][139],u_xpb_out[33][139],u_xpb_out[34][139],u_xpb_out[35][139],u_xpb_out[36][139],u_xpb_out[37][139],u_xpb_out[38][139],u_xpb_out[39][139],u_xpb_out[40][139],u_xpb_out[41][139],u_xpb_out[42][139],u_xpb_out[43][139],u_xpb_out[44][139],u_xpb_out[45][139],u_xpb_out[46][139],u_xpb_out[47][139],u_xpb_out[48][139],u_xpb_out[49][139],u_xpb_out[50][139],u_xpb_out[51][139],u_xpb_out[52][139],u_xpb_out[53][139],u_xpb_out[54][139],u_xpb_out[55][139],u_xpb_out[56][139],u_xpb_out[57][139],u_xpb_out[58][139],u_xpb_out[59][139],u_xpb_out[60][139],u_xpb_out[61][139],u_xpb_out[62][139],u_xpb_out[63][139],u_xpb_out[64][139],u_xpb_out[65][139],u_xpb_out[66][139],u_xpb_out[67][139],u_xpb_out[68][139],u_xpb_out[69][139],u_xpb_out[70][139],u_xpb_out[71][139],u_xpb_out[72][139],u_xpb_out[73][139],u_xpb_out[74][139],u_xpb_out[75][139],u_xpb_out[76][139],u_xpb_out[77][139],u_xpb_out[78][139],u_xpb_out[79][139],u_xpb_out[80][139],u_xpb_out[81][139],u_xpb_out[82][139],u_xpb_out[83][139],u_xpb_out[84][139],u_xpb_out[85][139],u_xpb_out[86][139],u_xpb_out[87][139],u_xpb_out[88][139],u_xpb_out[89][139],u_xpb_out[90][139],u_xpb_out[91][139],u_xpb_out[92][139],u_xpb_out[93][139],u_xpb_out[94][139],u_xpb_out[95][139],u_xpb_out[96][139],u_xpb_out[97][139],u_xpb_out[98][139],u_xpb_out[99][139],u_xpb_out[100][139],u_xpb_out[101][139],u_xpb_out[102][139],u_xpb_out[103][139],u_xpb_out[104][139],u_xpb_out[105][139]};

assign col_out_140 = {u_xpb_out[0][140],u_xpb_out[1][140],u_xpb_out[2][140],u_xpb_out[3][140],u_xpb_out[4][140],u_xpb_out[5][140],u_xpb_out[6][140],u_xpb_out[7][140],u_xpb_out[8][140],u_xpb_out[9][140],u_xpb_out[10][140],u_xpb_out[11][140],u_xpb_out[12][140],u_xpb_out[13][140],u_xpb_out[14][140],u_xpb_out[15][140],u_xpb_out[16][140],u_xpb_out[17][140],u_xpb_out[18][140],u_xpb_out[19][140],u_xpb_out[20][140],u_xpb_out[21][140],u_xpb_out[22][140],u_xpb_out[23][140],u_xpb_out[24][140],u_xpb_out[25][140],u_xpb_out[26][140],u_xpb_out[27][140],u_xpb_out[28][140],u_xpb_out[29][140],u_xpb_out[30][140],u_xpb_out[31][140],u_xpb_out[32][140],u_xpb_out[33][140],u_xpb_out[34][140],u_xpb_out[35][140],u_xpb_out[36][140],u_xpb_out[37][140],u_xpb_out[38][140],u_xpb_out[39][140],u_xpb_out[40][140],u_xpb_out[41][140],u_xpb_out[42][140],u_xpb_out[43][140],u_xpb_out[44][140],u_xpb_out[45][140],u_xpb_out[46][140],u_xpb_out[47][140],u_xpb_out[48][140],u_xpb_out[49][140],u_xpb_out[50][140],u_xpb_out[51][140],u_xpb_out[52][140],u_xpb_out[53][140],u_xpb_out[54][140],u_xpb_out[55][140],u_xpb_out[56][140],u_xpb_out[57][140],u_xpb_out[58][140],u_xpb_out[59][140],u_xpb_out[60][140],u_xpb_out[61][140],u_xpb_out[62][140],u_xpb_out[63][140],u_xpb_out[64][140],u_xpb_out[65][140],u_xpb_out[66][140],u_xpb_out[67][140],u_xpb_out[68][140],u_xpb_out[69][140],u_xpb_out[70][140],u_xpb_out[71][140],u_xpb_out[72][140],u_xpb_out[73][140],u_xpb_out[74][140],u_xpb_out[75][140],u_xpb_out[76][140],u_xpb_out[77][140],u_xpb_out[78][140],u_xpb_out[79][140],u_xpb_out[80][140],u_xpb_out[81][140],u_xpb_out[82][140],u_xpb_out[83][140],u_xpb_out[84][140],u_xpb_out[85][140],u_xpb_out[86][140],u_xpb_out[87][140],u_xpb_out[88][140],u_xpb_out[89][140],u_xpb_out[90][140],u_xpb_out[91][140],u_xpb_out[92][140],u_xpb_out[93][140],u_xpb_out[94][140],u_xpb_out[95][140],u_xpb_out[96][140],u_xpb_out[97][140],u_xpb_out[98][140],u_xpb_out[99][140],u_xpb_out[100][140],u_xpb_out[101][140],u_xpb_out[102][140],u_xpb_out[103][140],u_xpb_out[104][140],u_xpb_out[105][140]};

assign col_out_141 = {u_xpb_out[0][141],u_xpb_out[1][141],u_xpb_out[2][141],u_xpb_out[3][141],u_xpb_out[4][141],u_xpb_out[5][141],u_xpb_out[6][141],u_xpb_out[7][141],u_xpb_out[8][141],u_xpb_out[9][141],u_xpb_out[10][141],u_xpb_out[11][141],u_xpb_out[12][141],u_xpb_out[13][141],u_xpb_out[14][141],u_xpb_out[15][141],u_xpb_out[16][141],u_xpb_out[17][141],u_xpb_out[18][141],u_xpb_out[19][141],u_xpb_out[20][141],u_xpb_out[21][141],u_xpb_out[22][141],u_xpb_out[23][141],u_xpb_out[24][141],u_xpb_out[25][141],u_xpb_out[26][141],u_xpb_out[27][141],u_xpb_out[28][141],u_xpb_out[29][141],u_xpb_out[30][141],u_xpb_out[31][141],u_xpb_out[32][141],u_xpb_out[33][141],u_xpb_out[34][141],u_xpb_out[35][141],u_xpb_out[36][141],u_xpb_out[37][141],u_xpb_out[38][141],u_xpb_out[39][141],u_xpb_out[40][141],u_xpb_out[41][141],u_xpb_out[42][141],u_xpb_out[43][141],u_xpb_out[44][141],u_xpb_out[45][141],u_xpb_out[46][141],u_xpb_out[47][141],u_xpb_out[48][141],u_xpb_out[49][141],u_xpb_out[50][141],u_xpb_out[51][141],u_xpb_out[52][141],u_xpb_out[53][141],u_xpb_out[54][141],u_xpb_out[55][141],u_xpb_out[56][141],u_xpb_out[57][141],u_xpb_out[58][141],u_xpb_out[59][141],u_xpb_out[60][141],u_xpb_out[61][141],u_xpb_out[62][141],u_xpb_out[63][141],u_xpb_out[64][141],u_xpb_out[65][141],u_xpb_out[66][141],u_xpb_out[67][141],u_xpb_out[68][141],u_xpb_out[69][141],u_xpb_out[70][141],u_xpb_out[71][141],u_xpb_out[72][141],u_xpb_out[73][141],u_xpb_out[74][141],u_xpb_out[75][141],u_xpb_out[76][141],u_xpb_out[77][141],u_xpb_out[78][141],u_xpb_out[79][141],u_xpb_out[80][141],u_xpb_out[81][141],u_xpb_out[82][141],u_xpb_out[83][141],u_xpb_out[84][141],u_xpb_out[85][141],u_xpb_out[86][141],u_xpb_out[87][141],u_xpb_out[88][141],u_xpb_out[89][141],u_xpb_out[90][141],u_xpb_out[91][141],u_xpb_out[92][141],u_xpb_out[93][141],u_xpb_out[94][141],u_xpb_out[95][141],u_xpb_out[96][141],u_xpb_out[97][141],u_xpb_out[98][141],u_xpb_out[99][141],u_xpb_out[100][141],u_xpb_out[101][141],u_xpb_out[102][141],u_xpb_out[103][141],u_xpb_out[104][141],u_xpb_out[105][141]};

assign col_out_142 = {u_xpb_out[0][142],u_xpb_out[1][142],u_xpb_out[2][142],u_xpb_out[3][142],u_xpb_out[4][142],u_xpb_out[5][142],u_xpb_out[6][142],u_xpb_out[7][142],u_xpb_out[8][142],u_xpb_out[9][142],u_xpb_out[10][142],u_xpb_out[11][142],u_xpb_out[12][142],u_xpb_out[13][142],u_xpb_out[14][142],u_xpb_out[15][142],u_xpb_out[16][142],u_xpb_out[17][142],u_xpb_out[18][142],u_xpb_out[19][142],u_xpb_out[20][142],u_xpb_out[21][142],u_xpb_out[22][142],u_xpb_out[23][142],u_xpb_out[24][142],u_xpb_out[25][142],u_xpb_out[26][142],u_xpb_out[27][142],u_xpb_out[28][142],u_xpb_out[29][142],u_xpb_out[30][142],u_xpb_out[31][142],u_xpb_out[32][142],u_xpb_out[33][142],u_xpb_out[34][142],u_xpb_out[35][142],u_xpb_out[36][142],u_xpb_out[37][142],u_xpb_out[38][142],u_xpb_out[39][142],u_xpb_out[40][142],u_xpb_out[41][142],u_xpb_out[42][142],u_xpb_out[43][142],u_xpb_out[44][142],u_xpb_out[45][142],u_xpb_out[46][142],u_xpb_out[47][142],u_xpb_out[48][142],u_xpb_out[49][142],u_xpb_out[50][142],u_xpb_out[51][142],u_xpb_out[52][142],u_xpb_out[53][142],u_xpb_out[54][142],u_xpb_out[55][142],u_xpb_out[56][142],u_xpb_out[57][142],u_xpb_out[58][142],u_xpb_out[59][142],u_xpb_out[60][142],u_xpb_out[61][142],u_xpb_out[62][142],u_xpb_out[63][142],u_xpb_out[64][142],u_xpb_out[65][142],u_xpb_out[66][142],u_xpb_out[67][142],u_xpb_out[68][142],u_xpb_out[69][142],u_xpb_out[70][142],u_xpb_out[71][142],u_xpb_out[72][142],u_xpb_out[73][142],u_xpb_out[74][142],u_xpb_out[75][142],u_xpb_out[76][142],u_xpb_out[77][142],u_xpb_out[78][142],u_xpb_out[79][142],u_xpb_out[80][142],u_xpb_out[81][142],u_xpb_out[82][142],u_xpb_out[83][142],u_xpb_out[84][142],u_xpb_out[85][142],u_xpb_out[86][142],u_xpb_out[87][142],u_xpb_out[88][142],u_xpb_out[89][142],u_xpb_out[90][142],u_xpb_out[91][142],u_xpb_out[92][142],u_xpb_out[93][142],u_xpb_out[94][142],u_xpb_out[95][142],u_xpb_out[96][142],u_xpb_out[97][142],u_xpb_out[98][142],u_xpb_out[99][142],u_xpb_out[100][142],u_xpb_out[101][142],u_xpb_out[102][142],u_xpb_out[103][142],u_xpb_out[104][142],u_xpb_out[105][142]};

assign col_out_143 = {u_xpb_out[0][143],u_xpb_out[1][143],u_xpb_out[2][143],u_xpb_out[3][143],u_xpb_out[4][143],u_xpb_out[5][143],u_xpb_out[6][143],u_xpb_out[7][143],u_xpb_out[8][143],u_xpb_out[9][143],u_xpb_out[10][143],u_xpb_out[11][143],u_xpb_out[12][143],u_xpb_out[13][143],u_xpb_out[14][143],u_xpb_out[15][143],u_xpb_out[16][143],u_xpb_out[17][143],u_xpb_out[18][143],u_xpb_out[19][143],u_xpb_out[20][143],u_xpb_out[21][143],u_xpb_out[22][143],u_xpb_out[23][143],u_xpb_out[24][143],u_xpb_out[25][143],u_xpb_out[26][143],u_xpb_out[27][143],u_xpb_out[28][143],u_xpb_out[29][143],u_xpb_out[30][143],u_xpb_out[31][143],u_xpb_out[32][143],u_xpb_out[33][143],u_xpb_out[34][143],u_xpb_out[35][143],u_xpb_out[36][143],u_xpb_out[37][143],u_xpb_out[38][143],u_xpb_out[39][143],u_xpb_out[40][143],u_xpb_out[41][143],u_xpb_out[42][143],u_xpb_out[43][143],u_xpb_out[44][143],u_xpb_out[45][143],u_xpb_out[46][143],u_xpb_out[47][143],u_xpb_out[48][143],u_xpb_out[49][143],u_xpb_out[50][143],u_xpb_out[51][143],u_xpb_out[52][143],u_xpb_out[53][143],u_xpb_out[54][143],u_xpb_out[55][143],u_xpb_out[56][143],u_xpb_out[57][143],u_xpb_out[58][143],u_xpb_out[59][143],u_xpb_out[60][143],u_xpb_out[61][143],u_xpb_out[62][143],u_xpb_out[63][143],u_xpb_out[64][143],u_xpb_out[65][143],u_xpb_out[66][143],u_xpb_out[67][143],u_xpb_out[68][143],u_xpb_out[69][143],u_xpb_out[70][143],u_xpb_out[71][143],u_xpb_out[72][143],u_xpb_out[73][143],u_xpb_out[74][143],u_xpb_out[75][143],u_xpb_out[76][143],u_xpb_out[77][143],u_xpb_out[78][143],u_xpb_out[79][143],u_xpb_out[80][143],u_xpb_out[81][143],u_xpb_out[82][143],u_xpb_out[83][143],u_xpb_out[84][143],u_xpb_out[85][143],u_xpb_out[86][143],u_xpb_out[87][143],u_xpb_out[88][143],u_xpb_out[89][143],u_xpb_out[90][143],u_xpb_out[91][143],u_xpb_out[92][143],u_xpb_out[93][143],u_xpb_out[94][143],u_xpb_out[95][143],u_xpb_out[96][143],u_xpb_out[97][143],u_xpb_out[98][143],u_xpb_out[99][143],u_xpb_out[100][143],u_xpb_out[101][143],u_xpb_out[102][143],u_xpb_out[103][143],u_xpb_out[104][143],u_xpb_out[105][143]};

assign col_out_144 = {u_xpb_out[0][144],u_xpb_out[1][144],u_xpb_out[2][144],u_xpb_out[3][144],u_xpb_out[4][144],u_xpb_out[5][144],u_xpb_out[6][144],u_xpb_out[7][144],u_xpb_out[8][144],u_xpb_out[9][144],u_xpb_out[10][144],u_xpb_out[11][144],u_xpb_out[12][144],u_xpb_out[13][144],u_xpb_out[14][144],u_xpb_out[15][144],u_xpb_out[16][144],u_xpb_out[17][144],u_xpb_out[18][144],u_xpb_out[19][144],u_xpb_out[20][144],u_xpb_out[21][144],u_xpb_out[22][144],u_xpb_out[23][144],u_xpb_out[24][144],u_xpb_out[25][144],u_xpb_out[26][144],u_xpb_out[27][144],u_xpb_out[28][144],u_xpb_out[29][144],u_xpb_out[30][144],u_xpb_out[31][144],u_xpb_out[32][144],u_xpb_out[33][144],u_xpb_out[34][144],u_xpb_out[35][144],u_xpb_out[36][144],u_xpb_out[37][144],u_xpb_out[38][144],u_xpb_out[39][144],u_xpb_out[40][144],u_xpb_out[41][144],u_xpb_out[42][144],u_xpb_out[43][144],u_xpb_out[44][144],u_xpb_out[45][144],u_xpb_out[46][144],u_xpb_out[47][144],u_xpb_out[48][144],u_xpb_out[49][144],u_xpb_out[50][144],u_xpb_out[51][144],u_xpb_out[52][144],u_xpb_out[53][144],u_xpb_out[54][144],u_xpb_out[55][144],u_xpb_out[56][144],u_xpb_out[57][144],u_xpb_out[58][144],u_xpb_out[59][144],u_xpb_out[60][144],u_xpb_out[61][144],u_xpb_out[62][144],u_xpb_out[63][144],u_xpb_out[64][144],u_xpb_out[65][144],u_xpb_out[66][144],u_xpb_out[67][144],u_xpb_out[68][144],u_xpb_out[69][144],u_xpb_out[70][144],u_xpb_out[71][144],u_xpb_out[72][144],u_xpb_out[73][144],u_xpb_out[74][144],u_xpb_out[75][144],u_xpb_out[76][144],u_xpb_out[77][144],u_xpb_out[78][144],u_xpb_out[79][144],u_xpb_out[80][144],u_xpb_out[81][144],u_xpb_out[82][144],u_xpb_out[83][144],u_xpb_out[84][144],u_xpb_out[85][144],u_xpb_out[86][144],u_xpb_out[87][144],u_xpb_out[88][144],u_xpb_out[89][144],u_xpb_out[90][144],u_xpb_out[91][144],u_xpb_out[92][144],u_xpb_out[93][144],u_xpb_out[94][144],u_xpb_out[95][144],u_xpb_out[96][144],u_xpb_out[97][144],u_xpb_out[98][144],u_xpb_out[99][144],u_xpb_out[100][144],u_xpb_out[101][144],u_xpb_out[102][144],u_xpb_out[103][144],u_xpb_out[104][144],u_xpb_out[105][144]};

assign col_out_145 = {u_xpb_out[0][145],u_xpb_out[1][145],u_xpb_out[2][145],u_xpb_out[3][145],u_xpb_out[4][145],u_xpb_out[5][145],u_xpb_out[6][145],u_xpb_out[7][145],u_xpb_out[8][145],u_xpb_out[9][145],u_xpb_out[10][145],u_xpb_out[11][145],u_xpb_out[12][145],u_xpb_out[13][145],u_xpb_out[14][145],u_xpb_out[15][145],u_xpb_out[16][145],u_xpb_out[17][145],u_xpb_out[18][145],u_xpb_out[19][145],u_xpb_out[20][145],u_xpb_out[21][145],u_xpb_out[22][145],u_xpb_out[23][145],u_xpb_out[24][145],u_xpb_out[25][145],u_xpb_out[26][145],u_xpb_out[27][145],u_xpb_out[28][145],u_xpb_out[29][145],u_xpb_out[30][145],u_xpb_out[31][145],u_xpb_out[32][145],u_xpb_out[33][145],u_xpb_out[34][145],u_xpb_out[35][145],u_xpb_out[36][145],u_xpb_out[37][145],u_xpb_out[38][145],u_xpb_out[39][145],u_xpb_out[40][145],u_xpb_out[41][145],u_xpb_out[42][145],u_xpb_out[43][145],u_xpb_out[44][145],u_xpb_out[45][145],u_xpb_out[46][145],u_xpb_out[47][145],u_xpb_out[48][145],u_xpb_out[49][145],u_xpb_out[50][145],u_xpb_out[51][145],u_xpb_out[52][145],u_xpb_out[53][145],u_xpb_out[54][145],u_xpb_out[55][145],u_xpb_out[56][145],u_xpb_out[57][145],u_xpb_out[58][145],u_xpb_out[59][145],u_xpb_out[60][145],u_xpb_out[61][145],u_xpb_out[62][145],u_xpb_out[63][145],u_xpb_out[64][145],u_xpb_out[65][145],u_xpb_out[66][145],u_xpb_out[67][145],u_xpb_out[68][145],u_xpb_out[69][145],u_xpb_out[70][145],u_xpb_out[71][145],u_xpb_out[72][145],u_xpb_out[73][145],u_xpb_out[74][145],u_xpb_out[75][145],u_xpb_out[76][145],u_xpb_out[77][145],u_xpb_out[78][145],u_xpb_out[79][145],u_xpb_out[80][145],u_xpb_out[81][145],u_xpb_out[82][145],u_xpb_out[83][145],u_xpb_out[84][145],u_xpb_out[85][145],u_xpb_out[86][145],u_xpb_out[87][145],u_xpb_out[88][145],u_xpb_out[89][145],u_xpb_out[90][145],u_xpb_out[91][145],u_xpb_out[92][145],u_xpb_out[93][145],u_xpb_out[94][145],u_xpb_out[95][145],u_xpb_out[96][145],u_xpb_out[97][145],u_xpb_out[98][145],u_xpb_out[99][145],u_xpb_out[100][145],u_xpb_out[101][145],u_xpb_out[102][145],u_xpb_out[103][145],u_xpb_out[104][145],u_xpb_out[105][145]};

assign col_out_146 = {u_xpb_out[0][146],u_xpb_out[1][146],u_xpb_out[2][146],u_xpb_out[3][146],u_xpb_out[4][146],u_xpb_out[5][146],u_xpb_out[6][146],u_xpb_out[7][146],u_xpb_out[8][146],u_xpb_out[9][146],u_xpb_out[10][146],u_xpb_out[11][146],u_xpb_out[12][146],u_xpb_out[13][146],u_xpb_out[14][146],u_xpb_out[15][146],u_xpb_out[16][146],u_xpb_out[17][146],u_xpb_out[18][146],u_xpb_out[19][146],u_xpb_out[20][146],u_xpb_out[21][146],u_xpb_out[22][146],u_xpb_out[23][146],u_xpb_out[24][146],u_xpb_out[25][146],u_xpb_out[26][146],u_xpb_out[27][146],u_xpb_out[28][146],u_xpb_out[29][146],u_xpb_out[30][146],u_xpb_out[31][146],u_xpb_out[32][146],u_xpb_out[33][146],u_xpb_out[34][146],u_xpb_out[35][146],u_xpb_out[36][146],u_xpb_out[37][146],u_xpb_out[38][146],u_xpb_out[39][146],u_xpb_out[40][146],u_xpb_out[41][146],u_xpb_out[42][146],u_xpb_out[43][146],u_xpb_out[44][146],u_xpb_out[45][146],u_xpb_out[46][146],u_xpb_out[47][146],u_xpb_out[48][146],u_xpb_out[49][146],u_xpb_out[50][146],u_xpb_out[51][146],u_xpb_out[52][146],u_xpb_out[53][146],u_xpb_out[54][146],u_xpb_out[55][146],u_xpb_out[56][146],u_xpb_out[57][146],u_xpb_out[58][146],u_xpb_out[59][146],u_xpb_out[60][146],u_xpb_out[61][146],u_xpb_out[62][146],u_xpb_out[63][146],u_xpb_out[64][146],u_xpb_out[65][146],u_xpb_out[66][146],u_xpb_out[67][146],u_xpb_out[68][146],u_xpb_out[69][146],u_xpb_out[70][146],u_xpb_out[71][146],u_xpb_out[72][146],u_xpb_out[73][146],u_xpb_out[74][146],u_xpb_out[75][146],u_xpb_out[76][146],u_xpb_out[77][146],u_xpb_out[78][146],u_xpb_out[79][146],u_xpb_out[80][146],u_xpb_out[81][146],u_xpb_out[82][146],u_xpb_out[83][146],u_xpb_out[84][146],u_xpb_out[85][146],u_xpb_out[86][146],u_xpb_out[87][146],u_xpb_out[88][146],u_xpb_out[89][146],u_xpb_out[90][146],u_xpb_out[91][146],u_xpb_out[92][146],u_xpb_out[93][146],u_xpb_out[94][146],u_xpb_out[95][146],u_xpb_out[96][146],u_xpb_out[97][146],u_xpb_out[98][146],u_xpb_out[99][146],u_xpb_out[100][146],u_xpb_out[101][146],u_xpb_out[102][146],u_xpb_out[103][146],u_xpb_out[104][146],u_xpb_out[105][146]};

assign col_out_147 = {u_xpb_out[0][147],u_xpb_out[1][147],u_xpb_out[2][147],u_xpb_out[3][147],u_xpb_out[4][147],u_xpb_out[5][147],u_xpb_out[6][147],u_xpb_out[7][147],u_xpb_out[8][147],u_xpb_out[9][147],u_xpb_out[10][147],u_xpb_out[11][147],u_xpb_out[12][147],u_xpb_out[13][147],u_xpb_out[14][147],u_xpb_out[15][147],u_xpb_out[16][147],u_xpb_out[17][147],u_xpb_out[18][147],u_xpb_out[19][147],u_xpb_out[20][147],u_xpb_out[21][147],u_xpb_out[22][147],u_xpb_out[23][147],u_xpb_out[24][147],u_xpb_out[25][147],u_xpb_out[26][147],u_xpb_out[27][147],u_xpb_out[28][147],u_xpb_out[29][147],u_xpb_out[30][147],u_xpb_out[31][147],u_xpb_out[32][147],u_xpb_out[33][147],u_xpb_out[34][147],u_xpb_out[35][147],u_xpb_out[36][147],u_xpb_out[37][147],u_xpb_out[38][147],u_xpb_out[39][147],u_xpb_out[40][147],u_xpb_out[41][147],u_xpb_out[42][147],u_xpb_out[43][147],u_xpb_out[44][147],u_xpb_out[45][147],u_xpb_out[46][147],u_xpb_out[47][147],u_xpb_out[48][147],u_xpb_out[49][147],u_xpb_out[50][147],u_xpb_out[51][147],u_xpb_out[52][147],u_xpb_out[53][147],u_xpb_out[54][147],u_xpb_out[55][147],u_xpb_out[56][147],u_xpb_out[57][147],u_xpb_out[58][147],u_xpb_out[59][147],u_xpb_out[60][147],u_xpb_out[61][147],u_xpb_out[62][147],u_xpb_out[63][147],u_xpb_out[64][147],u_xpb_out[65][147],u_xpb_out[66][147],u_xpb_out[67][147],u_xpb_out[68][147],u_xpb_out[69][147],u_xpb_out[70][147],u_xpb_out[71][147],u_xpb_out[72][147],u_xpb_out[73][147],u_xpb_out[74][147],u_xpb_out[75][147],u_xpb_out[76][147],u_xpb_out[77][147],u_xpb_out[78][147],u_xpb_out[79][147],u_xpb_out[80][147],u_xpb_out[81][147],u_xpb_out[82][147],u_xpb_out[83][147],u_xpb_out[84][147],u_xpb_out[85][147],u_xpb_out[86][147],u_xpb_out[87][147],u_xpb_out[88][147],u_xpb_out[89][147],u_xpb_out[90][147],u_xpb_out[91][147],u_xpb_out[92][147],u_xpb_out[93][147],u_xpb_out[94][147],u_xpb_out[95][147],u_xpb_out[96][147],u_xpb_out[97][147],u_xpb_out[98][147],u_xpb_out[99][147],u_xpb_out[100][147],u_xpb_out[101][147],u_xpb_out[102][147],u_xpb_out[103][147],u_xpb_out[104][147],u_xpb_out[105][147]};

assign col_out_148 = {u_xpb_out[0][148],u_xpb_out[1][148],u_xpb_out[2][148],u_xpb_out[3][148],u_xpb_out[4][148],u_xpb_out[5][148],u_xpb_out[6][148],u_xpb_out[7][148],u_xpb_out[8][148],u_xpb_out[9][148],u_xpb_out[10][148],u_xpb_out[11][148],u_xpb_out[12][148],u_xpb_out[13][148],u_xpb_out[14][148],u_xpb_out[15][148],u_xpb_out[16][148],u_xpb_out[17][148],u_xpb_out[18][148],u_xpb_out[19][148],u_xpb_out[20][148],u_xpb_out[21][148],u_xpb_out[22][148],u_xpb_out[23][148],u_xpb_out[24][148],u_xpb_out[25][148],u_xpb_out[26][148],u_xpb_out[27][148],u_xpb_out[28][148],u_xpb_out[29][148],u_xpb_out[30][148],u_xpb_out[31][148],u_xpb_out[32][148],u_xpb_out[33][148],u_xpb_out[34][148],u_xpb_out[35][148],u_xpb_out[36][148],u_xpb_out[37][148],u_xpb_out[38][148],u_xpb_out[39][148],u_xpb_out[40][148],u_xpb_out[41][148],u_xpb_out[42][148],u_xpb_out[43][148],u_xpb_out[44][148],u_xpb_out[45][148],u_xpb_out[46][148],u_xpb_out[47][148],u_xpb_out[48][148],u_xpb_out[49][148],u_xpb_out[50][148],u_xpb_out[51][148],u_xpb_out[52][148],u_xpb_out[53][148],u_xpb_out[54][148],u_xpb_out[55][148],u_xpb_out[56][148],u_xpb_out[57][148],u_xpb_out[58][148],u_xpb_out[59][148],u_xpb_out[60][148],u_xpb_out[61][148],u_xpb_out[62][148],u_xpb_out[63][148],u_xpb_out[64][148],u_xpb_out[65][148],u_xpb_out[66][148],u_xpb_out[67][148],u_xpb_out[68][148],u_xpb_out[69][148],u_xpb_out[70][148],u_xpb_out[71][148],u_xpb_out[72][148],u_xpb_out[73][148],u_xpb_out[74][148],u_xpb_out[75][148],u_xpb_out[76][148],u_xpb_out[77][148],u_xpb_out[78][148],u_xpb_out[79][148],u_xpb_out[80][148],u_xpb_out[81][148],u_xpb_out[82][148],u_xpb_out[83][148],u_xpb_out[84][148],u_xpb_out[85][148],u_xpb_out[86][148],u_xpb_out[87][148],u_xpb_out[88][148],u_xpb_out[89][148],u_xpb_out[90][148],u_xpb_out[91][148],u_xpb_out[92][148],u_xpb_out[93][148],u_xpb_out[94][148],u_xpb_out[95][148],u_xpb_out[96][148],u_xpb_out[97][148],u_xpb_out[98][148],u_xpb_out[99][148],u_xpb_out[100][148],u_xpb_out[101][148],u_xpb_out[102][148],u_xpb_out[103][148],u_xpb_out[104][148],u_xpb_out[105][148]};

assign col_out_149 = {u_xpb_out[0][149],u_xpb_out[1][149],u_xpb_out[2][149],u_xpb_out[3][149],u_xpb_out[4][149],u_xpb_out[5][149],u_xpb_out[6][149],u_xpb_out[7][149],u_xpb_out[8][149],u_xpb_out[9][149],u_xpb_out[10][149],u_xpb_out[11][149],u_xpb_out[12][149],u_xpb_out[13][149],u_xpb_out[14][149],u_xpb_out[15][149],u_xpb_out[16][149],u_xpb_out[17][149],u_xpb_out[18][149],u_xpb_out[19][149],u_xpb_out[20][149],u_xpb_out[21][149],u_xpb_out[22][149],u_xpb_out[23][149],u_xpb_out[24][149],u_xpb_out[25][149],u_xpb_out[26][149],u_xpb_out[27][149],u_xpb_out[28][149],u_xpb_out[29][149],u_xpb_out[30][149],u_xpb_out[31][149],u_xpb_out[32][149],u_xpb_out[33][149],u_xpb_out[34][149],u_xpb_out[35][149],u_xpb_out[36][149],u_xpb_out[37][149],u_xpb_out[38][149],u_xpb_out[39][149],u_xpb_out[40][149],u_xpb_out[41][149],u_xpb_out[42][149],u_xpb_out[43][149],u_xpb_out[44][149],u_xpb_out[45][149],u_xpb_out[46][149],u_xpb_out[47][149],u_xpb_out[48][149],u_xpb_out[49][149],u_xpb_out[50][149],u_xpb_out[51][149],u_xpb_out[52][149],u_xpb_out[53][149],u_xpb_out[54][149],u_xpb_out[55][149],u_xpb_out[56][149],u_xpb_out[57][149],u_xpb_out[58][149],u_xpb_out[59][149],u_xpb_out[60][149],u_xpb_out[61][149],u_xpb_out[62][149],u_xpb_out[63][149],u_xpb_out[64][149],u_xpb_out[65][149],u_xpb_out[66][149],u_xpb_out[67][149],u_xpb_out[68][149],u_xpb_out[69][149],u_xpb_out[70][149],u_xpb_out[71][149],u_xpb_out[72][149],u_xpb_out[73][149],u_xpb_out[74][149],u_xpb_out[75][149],u_xpb_out[76][149],u_xpb_out[77][149],u_xpb_out[78][149],u_xpb_out[79][149],u_xpb_out[80][149],u_xpb_out[81][149],u_xpb_out[82][149],u_xpb_out[83][149],u_xpb_out[84][149],u_xpb_out[85][149],u_xpb_out[86][149],u_xpb_out[87][149],u_xpb_out[88][149],u_xpb_out[89][149],u_xpb_out[90][149],u_xpb_out[91][149],u_xpb_out[92][149],u_xpb_out[93][149],u_xpb_out[94][149],u_xpb_out[95][149],u_xpb_out[96][149],u_xpb_out[97][149],u_xpb_out[98][149],u_xpb_out[99][149],u_xpb_out[100][149],u_xpb_out[101][149],u_xpb_out[102][149],u_xpb_out[103][149],u_xpb_out[104][149],u_xpb_out[105][149]};

assign col_out_150 = {u_xpb_out[0][150],u_xpb_out[1][150],u_xpb_out[2][150],u_xpb_out[3][150],u_xpb_out[4][150],u_xpb_out[5][150],u_xpb_out[6][150],u_xpb_out[7][150],u_xpb_out[8][150],u_xpb_out[9][150],u_xpb_out[10][150],u_xpb_out[11][150],u_xpb_out[12][150],u_xpb_out[13][150],u_xpb_out[14][150],u_xpb_out[15][150],u_xpb_out[16][150],u_xpb_out[17][150],u_xpb_out[18][150],u_xpb_out[19][150],u_xpb_out[20][150],u_xpb_out[21][150],u_xpb_out[22][150],u_xpb_out[23][150],u_xpb_out[24][150],u_xpb_out[25][150],u_xpb_out[26][150],u_xpb_out[27][150],u_xpb_out[28][150],u_xpb_out[29][150],u_xpb_out[30][150],u_xpb_out[31][150],u_xpb_out[32][150],u_xpb_out[33][150],u_xpb_out[34][150],u_xpb_out[35][150],u_xpb_out[36][150],u_xpb_out[37][150],u_xpb_out[38][150],u_xpb_out[39][150],u_xpb_out[40][150],u_xpb_out[41][150],u_xpb_out[42][150],u_xpb_out[43][150],u_xpb_out[44][150],u_xpb_out[45][150],u_xpb_out[46][150],u_xpb_out[47][150],u_xpb_out[48][150],u_xpb_out[49][150],u_xpb_out[50][150],u_xpb_out[51][150],u_xpb_out[52][150],u_xpb_out[53][150],u_xpb_out[54][150],u_xpb_out[55][150],u_xpb_out[56][150],u_xpb_out[57][150],u_xpb_out[58][150],u_xpb_out[59][150],u_xpb_out[60][150],u_xpb_out[61][150],u_xpb_out[62][150],u_xpb_out[63][150],u_xpb_out[64][150],u_xpb_out[65][150],u_xpb_out[66][150],u_xpb_out[67][150],u_xpb_out[68][150],u_xpb_out[69][150],u_xpb_out[70][150],u_xpb_out[71][150],u_xpb_out[72][150],u_xpb_out[73][150],u_xpb_out[74][150],u_xpb_out[75][150],u_xpb_out[76][150],u_xpb_out[77][150],u_xpb_out[78][150],u_xpb_out[79][150],u_xpb_out[80][150],u_xpb_out[81][150],u_xpb_out[82][150],u_xpb_out[83][150],u_xpb_out[84][150],u_xpb_out[85][150],u_xpb_out[86][150],u_xpb_out[87][150],u_xpb_out[88][150],u_xpb_out[89][150],u_xpb_out[90][150],u_xpb_out[91][150],u_xpb_out[92][150],u_xpb_out[93][150],u_xpb_out[94][150],u_xpb_out[95][150],u_xpb_out[96][150],u_xpb_out[97][150],u_xpb_out[98][150],u_xpb_out[99][150],u_xpb_out[100][150],u_xpb_out[101][150],u_xpb_out[102][150],u_xpb_out[103][150],u_xpb_out[104][150],u_xpb_out[105][150]};

assign col_out_151 = {u_xpb_out[0][151],u_xpb_out[1][151],u_xpb_out[2][151],u_xpb_out[3][151],u_xpb_out[4][151],u_xpb_out[5][151],u_xpb_out[6][151],u_xpb_out[7][151],u_xpb_out[8][151],u_xpb_out[9][151],u_xpb_out[10][151],u_xpb_out[11][151],u_xpb_out[12][151],u_xpb_out[13][151],u_xpb_out[14][151],u_xpb_out[15][151],u_xpb_out[16][151],u_xpb_out[17][151],u_xpb_out[18][151],u_xpb_out[19][151],u_xpb_out[20][151],u_xpb_out[21][151],u_xpb_out[22][151],u_xpb_out[23][151],u_xpb_out[24][151],u_xpb_out[25][151],u_xpb_out[26][151],u_xpb_out[27][151],u_xpb_out[28][151],u_xpb_out[29][151],u_xpb_out[30][151],u_xpb_out[31][151],u_xpb_out[32][151],u_xpb_out[33][151],u_xpb_out[34][151],u_xpb_out[35][151],u_xpb_out[36][151],u_xpb_out[37][151],u_xpb_out[38][151],u_xpb_out[39][151],u_xpb_out[40][151],u_xpb_out[41][151],u_xpb_out[42][151],u_xpb_out[43][151],u_xpb_out[44][151],u_xpb_out[45][151],u_xpb_out[46][151],u_xpb_out[47][151],u_xpb_out[48][151],u_xpb_out[49][151],u_xpb_out[50][151],u_xpb_out[51][151],u_xpb_out[52][151],u_xpb_out[53][151],u_xpb_out[54][151],u_xpb_out[55][151],u_xpb_out[56][151],u_xpb_out[57][151],u_xpb_out[58][151],u_xpb_out[59][151],u_xpb_out[60][151],u_xpb_out[61][151],u_xpb_out[62][151],u_xpb_out[63][151],u_xpb_out[64][151],u_xpb_out[65][151],u_xpb_out[66][151],u_xpb_out[67][151],u_xpb_out[68][151],u_xpb_out[69][151],u_xpb_out[70][151],u_xpb_out[71][151],u_xpb_out[72][151],u_xpb_out[73][151],u_xpb_out[74][151],u_xpb_out[75][151],u_xpb_out[76][151],u_xpb_out[77][151],u_xpb_out[78][151],u_xpb_out[79][151],u_xpb_out[80][151],u_xpb_out[81][151],u_xpb_out[82][151],u_xpb_out[83][151],u_xpb_out[84][151],u_xpb_out[85][151],u_xpb_out[86][151],u_xpb_out[87][151],u_xpb_out[88][151],u_xpb_out[89][151],u_xpb_out[90][151],u_xpb_out[91][151],u_xpb_out[92][151],u_xpb_out[93][151],u_xpb_out[94][151],u_xpb_out[95][151],u_xpb_out[96][151],u_xpb_out[97][151],u_xpb_out[98][151],u_xpb_out[99][151],u_xpb_out[100][151],u_xpb_out[101][151],u_xpb_out[102][151],u_xpb_out[103][151],u_xpb_out[104][151],u_xpb_out[105][151]};

assign col_out_152 = {u_xpb_out[0][152],u_xpb_out[1][152],u_xpb_out[2][152],u_xpb_out[3][152],u_xpb_out[4][152],u_xpb_out[5][152],u_xpb_out[6][152],u_xpb_out[7][152],u_xpb_out[8][152],u_xpb_out[9][152],u_xpb_out[10][152],u_xpb_out[11][152],u_xpb_out[12][152],u_xpb_out[13][152],u_xpb_out[14][152],u_xpb_out[15][152],u_xpb_out[16][152],u_xpb_out[17][152],u_xpb_out[18][152],u_xpb_out[19][152],u_xpb_out[20][152],u_xpb_out[21][152],u_xpb_out[22][152],u_xpb_out[23][152],u_xpb_out[24][152],u_xpb_out[25][152],u_xpb_out[26][152],u_xpb_out[27][152],u_xpb_out[28][152],u_xpb_out[29][152],u_xpb_out[30][152],u_xpb_out[31][152],u_xpb_out[32][152],u_xpb_out[33][152],u_xpb_out[34][152],u_xpb_out[35][152],u_xpb_out[36][152],u_xpb_out[37][152],u_xpb_out[38][152],u_xpb_out[39][152],u_xpb_out[40][152],u_xpb_out[41][152],u_xpb_out[42][152],u_xpb_out[43][152],u_xpb_out[44][152],u_xpb_out[45][152],u_xpb_out[46][152],u_xpb_out[47][152],u_xpb_out[48][152],u_xpb_out[49][152],u_xpb_out[50][152],u_xpb_out[51][152],u_xpb_out[52][152],u_xpb_out[53][152],u_xpb_out[54][152],u_xpb_out[55][152],u_xpb_out[56][152],u_xpb_out[57][152],u_xpb_out[58][152],u_xpb_out[59][152],u_xpb_out[60][152],u_xpb_out[61][152],u_xpb_out[62][152],u_xpb_out[63][152],u_xpb_out[64][152],u_xpb_out[65][152],u_xpb_out[66][152],u_xpb_out[67][152],u_xpb_out[68][152],u_xpb_out[69][152],u_xpb_out[70][152],u_xpb_out[71][152],u_xpb_out[72][152],u_xpb_out[73][152],u_xpb_out[74][152],u_xpb_out[75][152],u_xpb_out[76][152],u_xpb_out[77][152],u_xpb_out[78][152],u_xpb_out[79][152],u_xpb_out[80][152],u_xpb_out[81][152],u_xpb_out[82][152],u_xpb_out[83][152],u_xpb_out[84][152],u_xpb_out[85][152],u_xpb_out[86][152],u_xpb_out[87][152],u_xpb_out[88][152],u_xpb_out[89][152],u_xpb_out[90][152],u_xpb_out[91][152],u_xpb_out[92][152],u_xpb_out[93][152],u_xpb_out[94][152],u_xpb_out[95][152],u_xpb_out[96][152],u_xpb_out[97][152],u_xpb_out[98][152],u_xpb_out[99][152],u_xpb_out[100][152],u_xpb_out[101][152],u_xpb_out[102][152],u_xpb_out[103][152],u_xpb_out[104][152],u_xpb_out[105][152]};

assign col_out_153 = {u_xpb_out[0][153],u_xpb_out[1][153],u_xpb_out[2][153],u_xpb_out[3][153],u_xpb_out[4][153],u_xpb_out[5][153],u_xpb_out[6][153],u_xpb_out[7][153],u_xpb_out[8][153],u_xpb_out[9][153],u_xpb_out[10][153],u_xpb_out[11][153],u_xpb_out[12][153],u_xpb_out[13][153],u_xpb_out[14][153],u_xpb_out[15][153],u_xpb_out[16][153],u_xpb_out[17][153],u_xpb_out[18][153],u_xpb_out[19][153],u_xpb_out[20][153],u_xpb_out[21][153],u_xpb_out[22][153],u_xpb_out[23][153],u_xpb_out[24][153],u_xpb_out[25][153],u_xpb_out[26][153],u_xpb_out[27][153],u_xpb_out[28][153],u_xpb_out[29][153],u_xpb_out[30][153],u_xpb_out[31][153],u_xpb_out[32][153],u_xpb_out[33][153],u_xpb_out[34][153],u_xpb_out[35][153],u_xpb_out[36][153],u_xpb_out[37][153],u_xpb_out[38][153],u_xpb_out[39][153],u_xpb_out[40][153],u_xpb_out[41][153],u_xpb_out[42][153],u_xpb_out[43][153],u_xpb_out[44][153],u_xpb_out[45][153],u_xpb_out[46][153],u_xpb_out[47][153],u_xpb_out[48][153],u_xpb_out[49][153],u_xpb_out[50][153],u_xpb_out[51][153],u_xpb_out[52][153],u_xpb_out[53][153],u_xpb_out[54][153],u_xpb_out[55][153],u_xpb_out[56][153],u_xpb_out[57][153],u_xpb_out[58][153],u_xpb_out[59][153],u_xpb_out[60][153],u_xpb_out[61][153],u_xpb_out[62][153],u_xpb_out[63][153],u_xpb_out[64][153],u_xpb_out[65][153],u_xpb_out[66][153],u_xpb_out[67][153],u_xpb_out[68][153],u_xpb_out[69][153],u_xpb_out[70][153],u_xpb_out[71][153],u_xpb_out[72][153],u_xpb_out[73][153],u_xpb_out[74][153],u_xpb_out[75][153],u_xpb_out[76][153],u_xpb_out[77][153],u_xpb_out[78][153],u_xpb_out[79][153],u_xpb_out[80][153],u_xpb_out[81][153],u_xpb_out[82][153],u_xpb_out[83][153],u_xpb_out[84][153],u_xpb_out[85][153],u_xpb_out[86][153],u_xpb_out[87][153],u_xpb_out[88][153],u_xpb_out[89][153],u_xpb_out[90][153],u_xpb_out[91][153],u_xpb_out[92][153],u_xpb_out[93][153],u_xpb_out[94][153],u_xpb_out[95][153],u_xpb_out[96][153],u_xpb_out[97][153],u_xpb_out[98][153],u_xpb_out[99][153],u_xpb_out[100][153],u_xpb_out[101][153],u_xpb_out[102][153],u_xpb_out[103][153],u_xpb_out[104][153],u_xpb_out[105][153]};

assign col_out_154 = {u_xpb_out[0][154],u_xpb_out[1][154],u_xpb_out[2][154],u_xpb_out[3][154],u_xpb_out[4][154],u_xpb_out[5][154],u_xpb_out[6][154],u_xpb_out[7][154],u_xpb_out[8][154],u_xpb_out[9][154],u_xpb_out[10][154],u_xpb_out[11][154],u_xpb_out[12][154],u_xpb_out[13][154],u_xpb_out[14][154],u_xpb_out[15][154],u_xpb_out[16][154],u_xpb_out[17][154],u_xpb_out[18][154],u_xpb_out[19][154],u_xpb_out[20][154],u_xpb_out[21][154],u_xpb_out[22][154],u_xpb_out[23][154],u_xpb_out[24][154],u_xpb_out[25][154],u_xpb_out[26][154],u_xpb_out[27][154],u_xpb_out[28][154],u_xpb_out[29][154],u_xpb_out[30][154],u_xpb_out[31][154],u_xpb_out[32][154],u_xpb_out[33][154],u_xpb_out[34][154],u_xpb_out[35][154],u_xpb_out[36][154],u_xpb_out[37][154],u_xpb_out[38][154],u_xpb_out[39][154],u_xpb_out[40][154],u_xpb_out[41][154],u_xpb_out[42][154],u_xpb_out[43][154],u_xpb_out[44][154],u_xpb_out[45][154],u_xpb_out[46][154],u_xpb_out[47][154],u_xpb_out[48][154],u_xpb_out[49][154],u_xpb_out[50][154],u_xpb_out[51][154],u_xpb_out[52][154],u_xpb_out[53][154],u_xpb_out[54][154],u_xpb_out[55][154],u_xpb_out[56][154],u_xpb_out[57][154],u_xpb_out[58][154],u_xpb_out[59][154],u_xpb_out[60][154],u_xpb_out[61][154],u_xpb_out[62][154],u_xpb_out[63][154],u_xpb_out[64][154],u_xpb_out[65][154],u_xpb_out[66][154],u_xpb_out[67][154],u_xpb_out[68][154],u_xpb_out[69][154],u_xpb_out[70][154],u_xpb_out[71][154],u_xpb_out[72][154],u_xpb_out[73][154],u_xpb_out[74][154],u_xpb_out[75][154],u_xpb_out[76][154],u_xpb_out[77][154],u_xpb_out[78][154],u_xpb_out[79][154],u_xpb_out[80][154],u_xpb_out[81][154],u_xpb_out[82][154],u_xpb_out[83][154],u_xpb_out[84][154],u_xpb_out[85][154],u_xpb_out[86][154],u_xpb_out[87][154],u_xpb_out[88][154],u_xpb_out[89][154],u_xpb_out[90][154],u_xpb_out[91][154],u_xpb_out[92][154],u_xpb_out[93][154],u_xpb_out[94][154],u_xpb_out[95][154],u_xpb_out[96][154],u_xpb_out[97][154],u_xpb_out[98][154],u_xpb_out[99][154],u_xpb_out[100][154],u_xpb_out[101][154],u_xpb_out[102][154],u_xpb_out[103][154],u_xpb_out[104][154],u_xpb_out[105][154]};

assign col_out_155 = {u_xpb_out[0][155],u_xpb_out[1][155],u_xpb_out[2][155],u_xpb_out[3][155],u_xpb_out[4][155],u_xpb_out[5][155],u_xpb_out[6][155],u_xpb_out[7][155],u_xpb_out[8][155],u_xpb_out[9][155],u_xpb_out[10][155],u_xpb_out[11][155],u_xpb_out[12][155],u_xpb_out[13][155],u_xpb_out[14][155],u_xpb_out[15][155],u_xpb_out[16][155],u_xpb_out[17][155],u_xpb_out[18][155],u_xpb_out[19][155],u_xpb_out[20][155],u_xpb_out[21][155],u_xpb_out[22][155],u_xpb_out[23][155],u_xpb_out[24][155],u_xpb_out[25][155],u_xpb_out[26][155],u_xpb_out[27][155],u_xpb_out[28][155],u_xpb_out[29][155],u_xpb_out[30][155],u_xpb_out[31][155],u_xpb_out[32][155],u_xpb_out[33][155],u_xpb_out[34][155],u_xpb_out[35][155],u_xpb_out[36][155],u_xpb_out[37][155],u_xpb_out[38][155],u_xpb_out[39][155],u_xpb_out[40][155],u_xpb_out[41][155],u_xpb_out[42][155],u_xpb_out[43][155],u_xpb_out[44][155],u_xpb_out[45][155],u_xpb_out[46][155],u_xpb_out[47][155],u_xpb_out[48][155],u_xpb_out[49][155],u_xpb_out[50][155],u_xpb_out[51][155],u_xpb_out[52][155],u_xpb_out[53][155],u_xpb_out[54][155],u_xpb_out[55][155],u_xpb_out[56][155],u_xpb_out[57][155],u_xpb_out[58][155],u_xpb_out[59][155],u_xpb_out[60][155],u_xpb_out[61][155],u_xpb_out[62][155],u_xpb_out[63][155],u_xpb_out[64][155],u_xpb_out[65][155],u_xpb_out[66][155],u_xpb_out[67][155],u_xpb_out[68][155],u_xpb_out[69][155],u_xpb_out[70][155],u_xpb_out[71][155],u_xpb_out[72][155],u_xpb_out[73][155],u_xpb_out[74][155],u_xpb_out[75][155],u_xpb_out[76][155],u_xpb_out[77][155],u_xpb_out[78][155],u_xpb_out[79][155],u_xpb_out[80][155],u_xpb_out[81][155],u_xpb_out[82][155],u_xpb_out[83][155],u_xpb_out[84][155],u_xpb_out[85][155],u_xpb_out[86][155],u_xpb_out[87][155],u_xpb_out[88][155],u_xpb_out[89][155],u_xpb_out[90][155],u_xpb_out[91][155],u_xpb_out[92][155],u_xpb_out[93][155],u_xpb_out[94][155],u_xpb_out[95][155],u_xpb_out[96][155],u_xpb_out[97][155],u_xpb_out[98][155],u_xpb_out[99][155],u_xpb_out[100][155],u_xpb_out[101][155],u_xpb_out[102][155],u_xpb_out[103][155],u_xpb_out[104][155],u_xpb_out[105][155]};

assign col_out_156 = {u_xpb_out[0][156],u_xpb_out[1][156],u_xpb_out[2][156],u_xpb_out[3][156],u_xpb_out[4][156],u_xpb_out[5][156],u_xpb_out[6][156],u_xpb_out[7][156],u_xpb_out[8][156],u_xpb_out[9][156],u_xpb_out[10][156],u_xpb_out[11][156],u_xpb_out[12][156],u_xpb_out[13][156],u_xpb_out[14][156],u_xpb_out[15][156],u_xpb_out[16][156],u_xpb_out[17][156],u_xpb_out[18][156],u_xpb_out[19][156],u_xpb_out[20][156],u_xpb_out[21][156],u_xpb_out[22][156],u_xpb_out[23][156],u_xpb_out[24][156],u_xpb_out[25][156],u_xpb_out[26][156],u_xpb_out[27][156],u_xpb_out[28][156],u_xpb_out[29][156],u_xpb_out[30][156],u_xpb_out[31][156],u_xpb_out[32][156],u_xpb_out[33][156],u_xpb_out[34][156],u_xpb_out[35][156],u_xpb_out[36][156],u_xpb_out[37][156],u_xpb_out[38][156],u_xpb_out[39][156],u_xpb_out[40][156],u_xpb_out[41][156],u_xpb_out[42][156],u_xpb_out[43][156],u_xpb_out[44][156],u_xpb_out[45][156],u_xpb_out[46][156],u_xpb_out[47][156],u_xpb_out[48][156],u_xpb_out[49][156],u_xpb_out[50][156],u_xpb_out[51][156],u_xpb_out[52][156],u_xpb_out[53][156],u_xpb_out[54][156],u_xpb_out[55][156],u_xpb_out[56][156],u_xpb_out[57][156],u_xpb_out[58][156],u_xpb_out[59][156],u_xpb_out[60][156],u_xpb_out[61][156],u_xpb_out[62][156],u_xpb_out[63][156],u_xpb_out[64][156],u_xpb_out[65][156],u_xpb_out[66][156],u_xpb_out[67][156],u_xpb_out[68][156],u_xpb_out[69][156],u_xpb_out[70][156],u_xpb_out[71][156],u_xpb_out[72][156],u_xpb_out[73][156],u_xpb_out[74][156],u_xpb_out[75][156],u_xpb_out[76][156],u_xpb_out[77][156],u_xpb_out[78][156],u_xpb_out[79][156],u_xpb_out[80][156],u_xpb_out[81][156],u_xpb_out[82][156],u_xpb_out[83][156],u_xpb_out[84][156],u_xpb_out[85][156],u_xpb_out[86][156],u_xpb_out[87][156],u_xpb_out[88][156],u_xpb_out[89][156],u_xpb_out[90][156],u_xpb_out[91][156],u_xpb_out[92][156],u_xpb_out[93][156],u_xpb_out[94][156],u_xpb_out[95][156],u_xpb_out[96][156],u_xpb_out[97][156],u_xpb_out[98][156],u_xpb_out[99][156],u_xpb_out[100][156],u_xpb_out[101][156],u_xpb_out[102][156],u_xpb_out[103][156],u_xpb_out[104][156],u_xpb_out[105][156]};

assign col_out_157 = {u_xpb_out[0][157],u_xpb_out[1][157],u_xpb_out[2][157],u_xpb_out[3][157],u_xpb_out[4][157],u_xpb_out[5][157],u_xpb_out[6][157],u_xpb_out[7][157],u_xpb_out[8][157],u_xpb_out[9][157],u_xpb_out[10][157],u_xpb_out[11][157],u_xpb_out[12][157],u_xpb_out[13][157],u_xpb_out[14][157],u_xpb_out[15][157],u_xpb_out[16][157],u_xpb_out[17][157],u_xpb_out[18][157],u_xpb_out[19][157],u_xpb_out[20][157],u_xpb_out[21][157],u_xpb_out[22][157],u_xpb_out[23][157],u_xpb_out[24][157],u_xpb_out[25][157],u_xpb_out[26][157],u_xpb_out[27][157],u_xpb_out[28][157],u_xpb_out[29][157],u_xpb_out[30][157],u_xpb_out[31][157],u_xpb_out[32][157],u_xpb_out[33][157],u_xpb_out[34][157],u_xpb_out[35][157],u_xpb_out[36][157],u_xpb_out[37][157],u_xpb_out[38][157],u_xpb_out[39][157],u_xpb_out[40][157],u_xpb_out[41][157],u_xpb_out[42][157],u_xpb_out[43][157],u_xpb_out[44][157],u_xpb_out[45][157],u_xpb_out[46][157],u_xpb_out[47][157],u_xpb_out[48][157],u_xpb_out[49][157],u_xpb_out[50][157],u_xpb_out[51][157],u_xpb_out[52][157],u_xpb_out[53][157],u_xpb_out[54][157],u_xpb_out[55][157],u_xpb_out[56][157],u_xpb_out[57][157],u_xpb_out[58][157],u_xpb_out[59][157],u_xpb_out[60][157],u_xpb_out[61][157],u_xpb_out[62][157],u_xpb_out[63][157],u_xpb_out[64][157],u_xpb_out[65][157],u_xpb_out[66][157],u_xpb_out[67][157],u_xpb_out[68][157],u_xpb_out[69][157],u_xpb_out[70][157],u_xpb_out[71][157],u_xpb_out[72][157],u_xpb_out[73][157],u_xpb_out[74][157],u_xpb_out[75][157],u_xpb_out[76][157],u_xpb_out[77][157],u_xpb_out[78][157],u_xpb_out[79][157],u_xpb_out[80][157],u_xpb_out[81][157],u_xpb_out[82][157],u_xpb_out[83][157],u_xpb_out[84][157],u_xpb_out[85][157],u_xpb_out[86][157],u_xpb_out[87][157],u_xpb_out[88][157],u_xpb_out[89][157],u_xpb_out[90][157],u_xpb_out[91][157],u_xpb_out[92][157],u_xpb_out[93][157],u_xpb_out[94][157],u_xpb_out[95][157],u_xpb_out[96][157],u_xpb_out[97][157],u_xpb_out[98][157],u_xpb_out[99][157],u_xpb_out[100][157],u_xpb_out[101][157],u_xpb_out[102][157],u_xpb_out[103][157],u_xpb_out[104][157],u_xpb_out[105][157]};

assign col_out_158 = {u_xpb_out[0][158],u_xpb_out[1][158],u_xpb_out[2][158],u_xpb_out[3][158],u_xpb_out[4][158],u_xpb_out[5][158],u_xpb_out[6][158],u_xpb_out[7][158],u_xpb_out[8][158],u_xpb_out[9][158],u_xpb_out[10][158],u_xpb_out[11][158],u_xpb_out[12][158],u_xpb_out[13][158],u_xpb_out[14][158],u_xpb_out[15][158],u_xpb_out[16][158],u_xpb_out[17][158],u_xpb_out[18][158],u_xpb_out[19][158],u_xpb_out[20][158],u_xpb_out[21][158],u_xpb_out[22][158],u_xpb_out[23][158],u_xpb_out[24][158],u_xpb_out[25][158],u_xpb_out[26][158],u_xpb_out[27][158],u_xpb_out[28][158],u_xpb_out[29][158],u_xpb_out[30][158],u_xpb_out[31][158],u_xpb_out[32][158],u_xpb_out[33][158],u_xpb_out[34][158],u_xpb_out[35][158],u_xpb_out[36][158],u_xpb_out[37][158],u_xpb_out[38][158],u_xpb_out[39][158],u_xpb_out[40][158],u_xpb_out[41][158],u_xpb_out[42][158],u_xpb_out[43][158],u_xpb_out[44][158],u_xpb_out[45][158],u_xpb_out[46][158],u_xpb_out[47][158],u_xpb_out[48][158],u_xpb_out[49][158],u_xpb_out[50][158],u_xpb_out[51][158],u_xpb_out[52][158],u_xpb_out[53][158],u_xpb_out[54][158],u_xpb_out[55][158],u_xpb_out[56][158],u_xpb_out[57][158],u_xpb_out[58][158],u_xpb_out[59][158],u_xpb_out[60][158],u_xpb_out[61][158],u_xpb_out[62][158],u_xpb_out[63][158],u_xpb_out[64][158],u_xpb_out[65][158],u_xpb_out[66][158],u_xpb_out[67][158],u_xpb_out[68][158],u_xpb_out[69][158],u_xpb_out[70][158],u_xpb_out[71][158],u_xpb_out[72][158],u_xpb_out[73][158],u_xpb_out[74][158],u_xpb_out[75][158],u_xpb_out[76][158],u_xpb_out[77][158],u_xpb_out[78][158],u_xpb_out[79][158],u_xpb_out[80][158],u_xpb_out[81][158],u_xpb_out[82][158],u_xpb_out[83][158],u_xpb_out[84][158],u_xpb_out[85][158],u_xpb_out[86][158],u_xpb_out[87][158],u_xpb_out[88][158],u_xpb_out[89][158],u_xpb_out[90][158],u_xpb_out[91][158],u_xpb_out[92][158],u_xpb_out[93][158],u_xpb_out[94][158],u_xpb_out[95][158],u_xpb_out[96][158],u_xpb_out[97][158],u_xpb_out[98][158],u_xpb_out[99][158],u_xpb_out[100][158],u_xpb_out[101][158],u_xpb_out[102][158],u_xpb_out[103][158],u_xpb_out[104][158],u_xpb_out[105][158]};

assign col_out_159 = {u_xpb_out[0][159],u_xpb_out[1][159],u_xpb_out[2][159],u_xpb_out[3][159],u_xpb_out[4][159],u_xpb_out[5][159],u_xpb_out[6][159],u_xpb_out[7][159],u_xpb_out[8][159],u_xpb_out[9][159],u_xpb_out[10][159],u_xpb_out[11][159],u_xpb_out[12][159],u_xpb_out[13][159],u_xpb_out[14][159],u_xpb_out[15][159],u_xpb_out[16][159],u_xpb_out[17][159],u_xpb_out[18][159],u_xpb_out[19][159],u_xpb_out[20][159],u_xpb_out[21][159],u_xpb_out[22][159],u_xpb_out[23][159],u_xpb_out[24][159],u_xpb_out[25][159],u_xpb_out[26][159],u_xpb_out[27][159],u_xpb_out[28][159],u_xpb_out[29][159],u_xpb_out[30][159],u_xpb_out[31][159],u_xpb_out[32][159],u_xpb_out[33][159],u_xpb_out[34][159],u_xpb_out[35][159],u_xpb_out[36][159],u_xpb_out[37][159],u_xpb_out[38][159],u_xpb_out[39][159],u_xpb_out[40][159],u_xpb_out[41][159],u_xpb_out[42][159],u_xpb_out[43][159],u_xpb_out[44][159],u_xpb_out[45][159],u_xpb_out[46][159],u_xpb_out[47][159],u_xpb_out[48][159],u_xpb_out[49][159],u_xpb_out[50][159],u_xpb_out[51][159],u_xpb_out[52][159],u_xpb_out[53][159],u_xpb_out[54][159],u_xpb_out[55][159],u_xpb_out[56][159],u_xpb_out[57][159],u_xpb_out[58][159],u_xpb_out[59][159],u_xpb_out[60][159],u_xpb_out[61][159],u_xpb_out[62][159],u_xpb_out[63][159],u_xpb_out[64][159],u_xpb_out[65][159],u_xpb_out[66][159],u_xpb_out[67][159],u_xpb_out[68][159],u_xpb_out[69][159],u_xpb_out[70][159],u_xpb_out[71][159],u_xpb_out[72][159],u_xpb_out[73][159],u_xpb_out[74][159],u_xpb_out[75][159],u_xpb_out[76][159],u_xpb_out[77][159],u_xpb_out[78][159],u_xpb_out[79][159],u_xpb_out[80][159],u_xpb_out[81][159],u_xpb_out[82][159],u_xpb_out[83][159],u_xpb_out[84][159],u_xpb_out[85][159],u_xpb_out[86][159],u_xpb_out[87][159],u_xpb_out[88][159],u_xpb_out[89][159],u_xpb_out[90][159],u_xpb_out[91][159],u_xpb_out[92][159],u_xpb_out[93][159],u_xpb_out[94][159],u_xpb_out[95][159],u_xpb_out[96][159],u_xpb_out[97][159],u_xpb_out[98][159],u_xpb_out[99][159],u_xpb_out[100][159],u_xpb_out[101][159],u_xpb_out[102][159],u_xpb_out[103][159],u_xpb_out[104][159],u_xpb_out[105][159]};

assign col_out_160 = {u_xpb_out[0][160],u_xpb_out[1][160],u_xpb_out[2][160],u_xpb_out[3][160],u_xpb_out[4][160],u_xpb_out[5][160],u_xpb_out[6][160],u_xpb_out[7][160],u_xpb_out[8][160],u_xpb_out[9][160],u_xpb_out[10][160],u_xpb_out[11][160],u_xpb_out[12][160],u_xpb_out[13][160],u_xpb_out[14][160],u_xpb_out[15][160],u_xpb_out[16][160],u_xpb_out[17][160],u_xpb_out[18][160],u_xpb_out[19][160],u_xpb_out[20][160],u_xpb_out[21][160],u_xpb_out[22][160],u_xpb_out[23][160],u_xpb_out[24][160],u_xpb_out[25][160],u_xpb_out[26][160],u_xpb_out[27][160],u_xpb_out[28][160],u_xpb_out[29][160],u_xpb_out[30][160],u_xpb_out[31][160],u_xpb_out[32][160],u_xpb_out[33][160],u_xpb_out[34][160],u_xpb_out[35][160],u_xpb_out[36][160],u_xpb_out[37][160],u_xpb_out[38][160],u_xpb_out[39][160],u_xpb_out[40][160],u_xpb_out[41][160],u_xpb_out[42][160],u_xpb_out[43][160],u_xpb_out[44][160],u_xpb_out[45][160],u_xpb_out[46][160],u_xpb_out[47][160],u_xpb_out[48][160],u_xpb_out[49][160],u_xpb_out[50][160],u_xpb_out[51][160],u_xpb_out[52][160],u_xpb_out[53][160],u_xpb_out[54][160],u_xpb_out[55][160],u_xpb_out[56][160],u_xpb_out[57][160],u_xpb_out[58][160],u_xpb_out[59][160],u_xpb_out[60][160],u_xpb_out[61][160],u_xpb_out[62][160],u_xpb_out[63][160],u_xpb_out[64][160],u_xpb_out[65][160],u_xpb_out[66][160],u_xpb_out[67][160],u_xpb_out[68][160],u_xpb_out[69][160],u_xpb_out[70][160],u_xpb_out[71][160],u_xpb_out[72][160],u_xpb_out[73][160],u_xpb_out[74][160],u_xpb_out[75][160],u_xpb_out[76][160],u_xpb_out[77][160],u_xpb_out[78][160],u_xpb_out[79][160],u_xpb_out[80][160],u_xpb_out[81][160],u_xpb_out[82][160],u_xpb_out[83][160],u_xpb_out[84][160],u_xpb_out[85][160],u_xpb_out[86][160],u_xpb_out[87][160],u_xpb_out[88][160],u_xpb_out[89][160],u_xpb_out[90][160],u_xpb_out[91][160],u_xpb_out[92][160],u_xpb_out[93][160],u_xpb_out[94][160],u_xpb_out[95][160],u_xpb_out[96][160],u_xpb_out[97][160],u_xpb_out[98][160],u_xpb_out[99][160],u_xpb_out[100][160],u_xpb_out[101][160],u_xpb_out[102][160],u_xpb_out[103][160],u_xpb_out[104][160],u_xpb_out[105][160]};

assign col_out_161 = {u_xpb_out[0][161],u_xpb_out[1][161],u_xpb_out[2][161],u_xpb_out[3][161],u_xpb_out[4][161],u_xpb_out[5][161],u_xpb_out[6][161],u_xpb_out[7][161],u_xpb_out[8][161],u_xpb_out[9][161],u_xpb_out[10][161],u_xpb_out[11][161],u_xpb_out[12][161],u_xpb_out[13][161],u_xpb_out[14][161],u_xpb_out[15][161],u_xpb_out[16][161],u_xpb_out[17][161],u_xpb_out[18][161],u_xpb_out[19][161],u_xpb_out[20][161],u_xpb_out[21][161],u_xpb_out[22][161],u_xpb_out[23][161],u_xpb_out[24][161],u_xpb_out[25][161],u_xpb_out[26][161],u_xpb_out[27][161],u_xpb_out[28][161],u_xpb_out[29][161],u_xpb_out[30][161],u_xpb_out[31][161],u_xpb_out[32][161],u_xpb_out[33][161],u_xpb_out[34][161],u_xpb_out[35][161],u_xpb_out[36][161],u_xpb_out[37][161],u_xpb_out[38][161],u_xpb_out[39][161],u_xpb_out[40][161],u_xpb_out[41][161],u_xpb_out[42][161],u_xpb_out[43][161],u_xpb_out[44][161],u_xpb_out[45][161],u_xpb_out[46][161],u_xpb_out[47][161],u_xpb_out[48][161],u_xpb_out[49][161],u_xpb_out[50][161],u_xpb_out[51][161],u_xpb_out[52][161],u_xpb_out[53][161],u_xpb_out[54][161],u_xpb_out[55][161],u_xpb_out[56][161],u_xpb_out[57][161],u_xpb_out[58][161],u_xpb_out[59][161],u_xpb_out[60][161],u_xpb_out[61][161],u_xpb_out[62][161],u_xpb_out[63][161],u_xpb_out[64][161],u_xpb_out[65][161],u_xpb_out[66][161],u_xpb_out[67][161],u_xpb_out[68][161],u_xpb_out[69][161],u_xpb_out[70][161],u_xpb_out[71][161],u_xpb_out[72][161],u_xpb_out[73][161],u_xpb_out[74][161],u_xpb_out[75][161],u_xpb_out[76][161],u_xpb_out[77][161],u_xpb_out[78][161],u_xpb_out[79][161],u_xpb_out[80][161],u_xpb_out[81][161],u_xpb_out[82][161],u_xpb_out[83][161],u_xpb_out[84][161],u_xpb_out[85][161],u_xpb_out[86][161],u_xpb_out[87][161],u_xpb_out[88][161],u_xpb_out[89][161],u_xpb_out[90][161],u_xpb_out[91][161],u_xpb_out[92][161],u_xpb_out[93][161],u_xpb_out[94][161],u_xpb_out[95][161],u_xpb_out[96][161],u_xpb_out[97][161],u_xpb_out[98][161],u_xpb_out[99][161],u_xpb_out[100][161],u_xpb_out[101][161],u_xpb_out[102][161],u_xpb_out[103][161],u_xpb_out[104][161],u_xpb_out[105][161]};

assign col_out_162 = {u_xpb_out[0][162],u_xpb_out[1][162],u_xpb_out[2][162],u_xpb_out[3][162],u_xpb_out[4][162],u_xpb_out[5][162],u_xpb_out[6][162],u_xpb_out[7][162],u_xpb_out[8][162],u_xpb_out[9][162],u_xpb_out[10][162],u_xpb_out[11][162],u_xpb_out[12][162],u_xpb_out[13][162],u_xpb_out[14][162],u_xpb_out[15][162],u_xpb_out[16][162],u_xpb_out[17][162],u_xpb_out[18][162],u_xpb_out[19][162],u_xpb_out[20][162],u_xpb_out[21][162],u_xpb_out[22][162],u_xpb_out[23][162],u_xpb_out[24][162],u_xpb_out[25][162],u_xpb_out[26][162],u_xpb_out[27][162],u_xpb_out[28][162],u_xpb_out[29][162],u_xpb_out[30][162],u_xpb_out[31][162],u_xpb_out[32][162],u_xpb_out[33][162],u_xpb_out[34][162],u_xpb_out[35][162],u_xpb_out[36][162],u_xpb_out[37][162],u_xpb_out[38][162],u_xpb_out[39][162],u_xpb_out[40][162],u_xpb_out[41][162],u_xpb_out[42][162],u_xpb_out[43][162],u_xpb_out[44][162],u_xpb_out[45][162],u_xpb_out[46][162],u_xpb_out[47][162],u_xpb_out[48][162],u_xpb_out[49][162],u_xpb_out[50][162],u_xpb_out[51][162],u_xpb_out[52][162],u_xpb_out[53][162],u_xpb_out[54][162],u_xpb_out[55][162],u_xpb_out[56][162],u_xpb_out[57][162],u_xpb_out[58][162],u_xpb_out[59][162],u_xpb_out[60][162],u_xpb_out[61][162],u_xpb_out[62][162],u_xpb_out[63][162],u_xpb_out[64][162],u_xpb_out[65][162],u_xpb_out[66][162],u_xpb_out[67][162],u_xpb_out[68][162],u_xpb_out[69][162],u_xpb_out[70][162],u_xpb_out[71][162],u_xpb_out[72][162],u_xpb_out[73][162],u_xpb_out[74][162],u_xpb_out[75][162],u_xpb_out[76][162],u_xpb_out[77][162],u_xpb_out[78][162],u_xpb_out[79][162],u_xpb_out[80][162],u_xpb_out[81][162],u_xpb_out[82][162],u_xpb_out[83][162],u_xpb_out[84][162],u_xpb_out[85][162],u_xpb_out[86][162],u_xpb_out[87][162],u_xpb_out[88][162],u_xpb_out[89][162],u_xpb_out[90][162],u_xpb_out[91][162],u_xpb_out[92][162],u_xpb_out[93][162],u_xpb_out[94][162],u_xpb_out[95][162],u_xpb_out[96][162],u_xpb_out[97][162],u_xpb_out[98][162],u_xpb_out[99][162],u_xpb_out[100][162],u_xpb_out[101][162],u_xpb_out[102][162],u_xpb_out[103][162],u_xpb_out[104][162],u_xpb_out[105][162]};

assign col_out_163 = {u_xpb_out[0][163],u_xpb_out[1][163],u_xpb_out[2][163],u_xpb_out[3][163],u_xpb_out[4][163],u_xpb_out[5][163],u_xpb_out[6][163],u_xpb_out[7][163],u_xpb_out[8][163],u_xpb_out[9][163],u_xpb_out[10][163],u_xpb_out[11][163],u_xpb_out[12][163],u_xpb_out[13][163],u_xpb_out[14][163],u_xpb_out[15][163],u_xpb_out[16][163],u_xpb_out[17][163],u_xpb_out[18][163],u_xpb_out[19][163],u_xpb_out[20][163],u_xpb_out[21][163],u_xpb_out[22][163],u_xpb_out[23][163],u_xpb_out[24][163],u_xpb_out[25][163],u_xpb_out[26][163],u_xpb_out[27][163],u_xpb_out[28][163],u_xpb_out[29][163],u_xpb_out[30][163],u_xpb_out[31][163],u_xpb_out[32][163],u_xpb_out[33][163],u_xpb_out[34][163],u_xpb_out[35][163],u_xpb_out[36][163],u_xpb_out[37][163],u_xpb_out[38][163],u_xpb_out[39][163],u_xpb_out[40][163],u_xpb_out[41][163],u_xpb_out[42][163],u_xpb_out[43][163],u_xpb_out[44][163],u_xpb_out[45][163],u_xpb_out[46][163],u_xpb_out[47][163],u_xpb_out[48][163],u_xpb_out[49][163],u_xpb_out[50][163],u_xpb_out[51][163],u_xpb_out[52][163],u_xpb_out[53][163],u_xpb_out[54][163],u_xpb_out[55][163],u_xpb_out[56][163],u_xpb_out[57][163],u_xpb_out[58][163],u_xpb_out[59][163],u_xpb_out[60][163],u_xpb_out[61][163],u_xpb_out[62][163],u_xpb_out[63][163],u_xpb_out[64][163],u_xpb_out[65][163],u_xpb_out[66][163],u_xpb_out[67][163],u_xpb_out[68][163],u_xpb_out[69][163],u_xpb_out[70][163],u_xpb_out[71][163],u_xpb_out[72][163],u_xpb_out[73][163],u_xpb_out[74][163],u_xpb_out[75][163],u_xpb_out[76][163],u_xpb_out[77][163],u_xpb_out[78][163],u_xpb_out[79][163],u_xpb_out[80][163],u_xpb_out[81][163],u_xpb_out[82][163],u_xpb_out[83][163],u_xpb_out[84][163],u_xpb_out[85][163],u_xpb_out[86][163],u_xpb_out[87][163],u_xpb_out[88][163],u_xpb_out[89][163],u_xpb_out[90][163],u_xpb_out[91][163],u_xpb_out[92][163],u_xpb_out[93][163],u_xpb_out[94][163],u_xpb_out[95][163],u_xpb_out[96][163],u_xpb_out[97][163],u_xpb_out[98][163],u_xpb_out[99][163],u_xpb_out[100][163],u_xpb_out[101][163],u_xpb_out[102][163],u_xpb_out[103][163],u_xpb_out[104][163],u_xpb_out[105][163]};

assign col_out_164 = {u_xpb_out[0][164],u_xpb_out[1][164],u_xpb_out[2][164],u_xpb_out[3][164],u_xpb_out[4][164],u_xpb_out[5][164],u_xpb_out[6][164],u_xpb_out[7][164],u_xpb_out[8][164],u_xpb_out[9][164],u_xpb_out[10][164],u_xpb_out[11][164],u_xpb_out[12][164],u_xpb_out[13][164],u_xpb_out[14][164],u_xpb_out[15][164],u_xpb_out[16][164],u_xpb_out[17][164],u_xpb_out[18][164],u_xpb_out[19][164],u_xpb_out[20][164],u_xpb_out[21][164],u_xpb_out[22][164],u_xpb_out[23][164],u_xpb_out[24][164],u_xpb_out[25][164],u_xpb_out[26][164],u_xpb_out[27][164],u_xpb_out[28][164],u_xpb_out[29][164],u_xpb_out[30][164],u_xpb_out[31][164],u_xpb_out[32][164],u_xpb_out[33][164],u_xpb_out[34][164],u_xpb_out[35][164],u_xpb_out[36][164],u_xpb_out[37][164],u_xpb_out[38][164],u_xpb_out[39][164],u_xpb_out[40][164],u_xpb_out[41][164],u_xpb_out[42][164],u_xpb_out[43][164],u_xpb_out[44][164],u_xpb_out[45][164],u_xpb_out[46][164],u_xpb_out[47][164],u_xpb_out[48][164],u_xpb_out[49][164],u_xpb_out[50][164],u_xpb_out[51][164],u_xpb_out[52][164],u_xpb_out[53][164],u_xpb_out[54][164],u_xpb_out[55][164],u_xpb_out[56][164],u_xpb_out[57][164],u_xpb_out[58][164],u_xpb_out[59][164],u_xpb_out[60][164],u_xpb_out[61][164],u_xpb_out[62][164],u_xpb_out[63][164],u_xpb_out[64][164],u_xpb_out[65][164],u_xpb_out[66][164],u_xpb_out[67][164],u_xpb_out[68][164],u_xpb_out[69][164],u_xpb_out[70][164],u_xpb_out[71][164],u_xpb_out[72][164],u_xpb_out[73][164],u_xpb_out[74][164],u_xpb_out[75][164],u_xpb_out[76][164],u_xpb_out[77][164],u_xpb_out[78][164],u_xpb_out[79][164],u_xpb_out[80][164],u_xpb_out[81][164],u_xpb_out[82][164],u_xpb_out[83][164],u_xpb_out[84][164],u_xpb_out[85][164],u_xpb_out[86][164],u_xpb_out[87][164],u_xpb_out[88][164],u_xpb_out[89][164],u_xpb_out[90][164],u_xpb_out[91][164],u_xpb_out[92][164],u_xpb_out[93][164],u_xpb_out[94][164],u_xpb_out[95][164],u_xpb_out[96][164],u_xpb_out[97][164],u_xpb_out[98][164],u_xpb_out[99][164],u_xpb_out[100][164],u_xpb_out[101][164],u_xpb_out[102][164],u_xpb_out[103][164],u_xpb_out[104][164],u_xpb_out[105][164]};

assign col_out_165 = {u_xpb_out[0][165],u_xpb_out[1][165],u_xpb_out[2][165],u_xpb_out[3][165],u_xpb_out[4][165],u_xpb_out[5][165],u_xpb_out[6][165],u_xpb_out[7][165],u_xpb_out[8][165],u_xpb_out[9][165],u_xpb_out[10][165],u_xpb_out[11][165],u_xpb_out[12][165],u_xpb_out[13][165],u_xpb_out[14][165],u_xpb_out[15][165],u_xpb_out[16][165],u_xpb_out[17][165],u_xpb_out[18][165],u_xpb_out[19][165],u_xpb_out[20][165],u_xpb_out[21][165],u_xpb_out[22][165],u_xpb_out[23][165],u_xpb_out[24][165],u_xpb_out[25][165],u_xpb_out[26][165],u_xpb_out[27][165],u_xpb_out[28][165],u_xpb_out[29][165],u_xpb_out[30][165],u_xpb_out[31][165],u_xpb_out[32][165],u_xpb_out[33][165],u_xpb_out[34][165],u_xpb_out[35][165],u_xpb_out[36][165],u_xpb_out[37][165],u_xpb_out[38][165],u_xpb_out[39][165],u_xpb_out[40][165],u_xpb_out[41][165],u_xpb_out[42][165],u_xpb_out[43][165],u_xpb_out[44][165],u_xpb_out[45][165],u_xpb_out[46][165],u_xpb_out[47][165],u_xpb_out[48][165],u_xpb_out[49][165],u_xpb_out[50][165],u_xpb_out[51][165],u_xpb_out[52][165],u_xpb_out[53][165],u_xpb_out[54][165],u_xpb_out[55][165],u_xpb_out[56][165],u_xpb_out[57][165],u_xpb_out[58][165],u_xpb_out[59][165],u_xpb_out[60][165],u_xpb_out[61][165],u_xpb_out[62][165],u_xpb_out[63][165],u_xpb_out[64][165],u_xpb_out[65][165],u_xpb_out[66][165],u_xpb_out[67][165],u_xpb_out[68][165],u_xpb_out[69][165],u_xpb_out[70][165],u_xpb_out[71][165],u_xpb_out[72][165],u_xpb_out[73][165],u_xpb_out[74][165],u_xpb_out[75][165],u_xpb_out[76][165],u_xpb_out[77][165],u_xpb_out[78][165],u_xpb_out[79][165],u_xpb_out[80][165],u_xpb_out[81][165],u_xpb_out[82][165],u_xpb_out[83][165],u_xpb_out[84][165],u_xpb_out[85][165],u_xpb_out[86][165],u_xpb_out[87][165],u_xpb_out[88][165],u_xpb_out[89][165],u_xpb_out[90][165],u_xpb_out[91][165],u_xpb_out[92][165],u_xpb_out[93][165],u_xpb_out[94][165],u_xpb_out[95][165],u_xpb_out[96][165],u_xpb_out[97][165],u_xpb_out[98][165],u_xpb_out[99][165],u_xpb_out[100][165],u_xpb_out[101][165],u_xpb_out[102][165],u_xpb_out[103][165],u_xpb_out[104][165],u_xpb_out[105][165]};

assign col_out_166 = {u_xpb_out[0][166],u_xpb_out[1][166],u_xpb_out[2][166],u_xpb_out[3][166],u_xpb_out[4][166],u_xpb_out[5][166],u_xpb_out[6][166],u_xpb_out[7][166],u_xpb_out[8][166],u_xpb_out[9][166],u_xpb_out[10][166],u_xpb_out[11][166],u_xpb_out[12][166],u_xpb_out[13][166],u_xpb_out[14][166],u_xpb_out[15][166],u_xpb_out[16][166],u_xpb_out[17][166],u_xpb_out[18][166],u_xpb_out[19][166],u_xpb_out[20][166],u_xpb_out[21][166],u_xpb_out[22][166],u_xpb_out[23][166],u_xpb_out[24][166],u_xpb_out[25][166],u_xpb_out[26][166],u_xpb_out[27][166],u_xpb_out[28][166],u_xpb_out[29][166],u_xpb_out[30][166],u_xpb_out[31][166],u_xpb_out[32][166],u_xpb_out[33][166],u_xpb_out[34][166],u_xpb_out[35][166],u_xpb_out[36][166],u_xpb_out[37][166],u_xpb_out[38][166],u_xpb_out[39][166],u_xpb_out[40][166],u_xpb_out[41][166],u_xpb_out[42][166],u_xpb_out[43][166],u_xpb_out[44][166],u_xpb_out[45][166],u_xpb_out[46][166],u_xpb_out[47][166],u_xpb_out[48][166],u_xpb_out[49][166],u_xpb_out[50][166],u_xpb_out[51][166],u_xpb_out[52][166],u_xpb_out[53][166],u_xpb_out[54][166],u_xpb_out[55][166],u_xpb_out[56][166],u_xpb_out[57][166],u_xpb_out[58][166],u_xpb_out[59][166],u_xpb_out[60][166],u_xpb_out[61][166],u_xpb_out[62][166],u_xpb_out[63][166],u_xpb_out[64][166],u_xpb_out[65][166],u_xpb_out[66][166],u_xpb_out[67][166],u_xpb_out[68][166],u_xpb_out[69][166],u_xpb_out[70][166],u_xpb_out[71][166],u_xpb_out[72][166],u_xpb_out[73][166],u_xpb_out[74][166],u_xpb_out[75][166],u_xpb_out[76][166],u_xpb_out[77][166],u_xpb_out[78][166],u_xpb_out[79][166],u_xpb_out[80][166],u_xpb_out[81][166],u_xpb_out[82][166],u_xpb_out[83][166],u_xpb_out[84][166],u_xpb_out[85][166],u_xpb_out[86][166],u_xpb_out[87][166],u_xpb_out[88][166],u_xpb_out[89][166],u_xpb_out[90][166],u_xpb_out[91][166],u_xpb_out[92][166],u_xpb_out[93][166],u_xpb_out[94][166],u_xpb_out[95][166],u_xpb_out[96][166],u_xpb_out[97][166],u_xpb_out[98][166],u_xpb_out[99][166],u_xpb_out[100][166],u_xpb_out[101][166],u_xpb_out[102][166],u_xpb_out[103][166],u_xpb_out[104][166],u_xpb_out[105][166]};

assign col_out_167 = {u_xpb_out[0][167],u_xpb_out[1][167],u_xpb_out[2][167],u_xpb_out[3][167],u_xpb_out[4][167],u_xpb_out[5][167],u_xpb_out[6][167],u_xpb_out[7][167],u_xpb_out[8][167],u_xpb_out[9][167],u_xpb_out[10][167],u_xpb_out[11][167],u_xpb_out[12][167],u_xpb_out[13][167],u_xpb_out[14][167],u_xpb_out[15][167],u_xpb_out[16][167],u_xpb_out[17][167],u_xpb_out[18][167],u_xpb_out[19][167],u_xpb_out[20][167],u_xpb_out[21][167],u_xpb_out[22][167],u_xpb_out[23][167],u_xpb_out[24][167],u_xpb_out[25][167],u_xpb_out[26][167],u_xpb_out[27][167],u_xpb_out[28][167],u_xpb_out[29][167],u_xpb_out[30][167],u_xpb_out[31][167],u_xpb_out[32][167],u_xpb_out[33][167],u_xpb_out[34][167],u_xpb_out[35][167],u_xpb_out[36][167],u_xpb_out[37][167],u_xpb_out[38][167],u_xpb_out[39][167],u_xpb_out[40][167],u_xpb_out[41][167],u_xpb_out[42][167],u_xpb_out[43][167],u_xpb_out[44][167],u_xpb_out[45][167],u_xpb_out[46][167],u_xpb_out[47][167],u_xpb_out[48][167],u_xpb_out[49][167],u_xpb_out[50][167],u_xpb_out[51][167],u_xpb_out[52][167],u_xpb_out[53][167],u_xpb_out[54][167],u_xpb_out[55][167],u_xpb_out[56][167],u_xpb_out[57][167],u_xpb_out[58][167],u_xpb_out[59][167],u_xpb_out[60][167],u_xpb_out[61][167],u_xpb_out[62][167],u_xpb_out[63][167],u_xpb_out[64][167],u_xpb_out[65][167],u_xpb_out[66][167],u_xpb_out[67][167],u_xpb_out[68][167],u_xpb_out[69][167],u_xpb_out[70][167],u_xpb_out[71][167],u_xpb_out[72][167],u_xpb_out[73][167],u_xpb_out[74][167],u_xpb_out[75][167],u_xpb_out[76][167],u_xpb_out[77][167],u_xpb_out[78][167],u_xpb_out[79][167],u_xpb_out[80][167],u_xpb_out[81][167],u_xpb_out[82][167],u_xpb_out[83][167],u_xpb_out[84][167],u_xpb_out[85][167],u_xpb_out[86][167],u_xpb_out[87][167],u_xpb_out[88][167],u_xpb_out[89][167],u_xpb_out[90][167],u_xpb_out[91][167],u_xpb_out[92][167],u_xpb_out[93][167],u_xpb_out[94][167],u_xpb_out[95][167],u_xpb_out[96][167],u_xpb_out[97][167],u_xpb_out[98][167],u_xpb_out[99][167],u_xpb_out[100][167],u_xpb_out[101][167],u_xpb_out[102][167],u_xpb_out[103][167],u_xpb_out[104][167],u_xpb_out[105][167]};

assign col_out_168 = {u_xpb_out[0][168],u_xpb_out[1][168],u_xpb_out[2][168],u_xpb_out[3][168],u_xpb_out[4][168],u_xpb_out[5][168],u_xpb_out[6][168],u_xpb_out[7][168],u_xpb_out[8][168],u_xpb_out[9][168],u_xpb_out[10][168],u_xpb_out[11][168],u_xpb_out[12][168],u_xpb_out[13][168],u_xpb_out[14][168],u_xpb_out[15][168],u_xpb_out[16][168],u_xpb_out[17][168],u_xpb_out[18][168],u_xpb_out[19][168],u_xpb_out[20][168],u_xpb_out[21][168],u_xpb_out[22][168],u_xpb_out[23][168],u_xpb_out[24][168],u_xpb_out[25][168],u_xpb_out[26][168],u_xpb_out[27][168],u_xpb_out[28][168],u_xpb_out[29][168],u_xpb_out[30][168],u_xpb_out[31][168],u_xpb_out[32][168],u_xpb_out[33][168],u_xpb_out[34][168],u_xpb_out[35][168],u_xpb_out[36][168],u_xpb_out[37][168],u_xpb_out[38][168],u_xpb_out[39][168],u_xpb_out[40][168],u_xpb_out[41][168],u_xpb_out[42][168],u_xpb_out[43][168],u_xpb_out[44][168],u_xpb_out[45][168],u_xpb_out[46][168],u_xpb_out[47][168],u_xpb_out[48][168],u_xpb_out[49][168],u_xpb_out[50][168],u_xpb_out[51][168],u_xpb_out[52][168],u_xpb_out[53][168],u_xpb_out[54][168],u_xpb_out[55][168],u_xpb_out[56][168],u_xpb_out[57][168],u_xpb_out[58][168],u_xpb_out[59][168],u_xpb_out[60][168],u_xpb_out[61][168],u_xpb_out[62][168],u_xpb_out[63][168],u_xpb_out[64][168],u_xpb_out[65][168],u_xpb_out[66][168],u_xpb_out[67][168],u_xpb_out[68][168],u_xpb_out[69][168],u_xpb_out[70][168],u_xpb_out[71][168],u_xpb_out[72][168],u_xpb_out[73][168],u_xpb_out[74][168],u_xpb_out[75][168],u_xpb_out[76][168],u_xpb_out[77][168],u_xpb_out[78][168],u_xpb_out[79][168],u_xpb_out[80][168],u_xpb_out[81][168],u_xpb_out[82][168],u_xpb_out[83][168],u_xpb_out[84][168],u_xpb_out[85][168],u_xpb_out[86][168],u_xpb_out[87][168],u_xpb_out[88][168],u_xpb_out[89][168],u_xpb_out[90][168],u_xpb_out[91][168],u_xpb_out[92][168],u_xpb_out[93][168],u_xpb_out[94][168],u_xpb_out[95][168],u_xpb_out[96][168],u_xpb_out[97][168],u_xpb_out[98][168],u_xpb_out[99][168],u_xpb_out[100][168],u_xpb_out[101][168],u_xpb_out[102][168],u_xpb_out[103][168],u_xpb_out[104][168],u_xpb_out[105][168]};

assign col_out_169 = {u_xpb_out[0][169],u_xpb_out[1][169],u_xpb_out[2][169],u_xpb_out[3][169],u_xpb_out[4][169],u_xpb_out[5][169],u_xpb_out[6][169],u_xpb_out[7][169],u_xpb_out[8][169],u_xpb_out[9][169],u_xpb_out[10][169],u_xpb_out[11][169],u_xpb_out[12][169],u_xpb_out[13][169],u_xpb_out[14][169],u_xpb_out[15][169],u_xpb_out[16][169],u_xpb_out[17][169],u_xpb_out[18][169],u_xpb_out[19][169],u_xpb_out[20][169],u_xpb_out[21][169],u_xpb_out[22][169],u_xpb_out[23][169],u_xpb_out[24][169],u_xpb_out[25][169],u_xpb_out[26][169],u_xpb_out[27][169],u_xpb_out[28][169],u_xpb_out[29][169],u_xpb_out[30][169],u_xpb_out[31][169],u_xpb_out[32][169],u_xpb_out[33][169],u_xpb_out[34][169],u_xpb_out[35][169],u_xpb_out[36][169],u_xpb_out[37][169],u_xpb_out[38][169],u_xpb_out[39][169],u_xpb_out[40][169],u_xpb_out[41][169],u_xpb_out[42][169],u_xpb_out[43][169],u_xpb_out[44][169],u_xpb_out[45][169],u_xpb_out[46][169],u_xpb_out[47][169],u_xpb_out[48][169],u_xpb_out[49][169],u_xpb_out[50][169],u_xpb_out[51][169],u_xpb_out[52][169],u_xpb_out[53][169],u_xpb_out[54][169],u_xpb_out[55][169],u_xpb_out[56][169],u_xpb_out[57][169],u_xpb_out[58][169],u_xpb_out[59][169],u_xpb_out[60][169],u_xpb_out[61][169],u_xpb_out[62][169],u_xpb_out[63][169],u_xpb_out[64][169],u_xpb_out[65][169],u_xpb_out[66][169],u_xpb_out[67][169],u_xpb_out[68][169],u_xpb_out[69][169],u_xpb_out[70][169],u_xpb_out[71][169],u_xpb_out[72][169],u_xpb_out[73][169],u_xpb_out[74][169],u_xpb_out[75][169],u_xpb_out[76][169],u_xpb_out[77][169],u_xpb_out[78][169],u_xpb_out[79][169],u_xpb_out[80][169],u_xpb_out[81][169],u_xpb_out[82][169],u_xpb_out[83][169],u_xpb_out[84][169],u_xpb_out[85][169],u_xpb_out[86][169],u_xpb_out[87][169],u_xpb_out[88][169],u_xpb_out[89][169],u_xpb_out[90][169],u_xpb_out[91][169],u_xpb_out[92][169],u_xpb_out[93][169],u_xpb_out[94][169],u_xpb_out[95][169],u_xpb_out[96][169],u_xpb_out[97][169],u_xpb_out[98][169],u_xpb_out[99][169],u_xpb_out[100][169],u_xpb_out[101][169],u_xpb_out[102][169],u_xpb_out[103][169],u_xpb_out[104][169],u_xpb_out[105][169]};

assign col_out_170 = {u_xpb_out[0][170],u_xpb_out[1][170],u_xpb_out[2][170],u_xpb_out[3][170],u_xpb_out[4][170],u_xpb_out[5][170],u_xpb_out[6][170],u_xpb_out[7][170],u_xpb_out[8][170],u_xpb_out[9][170],u_xpb_out[10][170],u_xpb_out[11][170],u_xpb_out[12][170],u_xpb_out[13][170],u_xpb_out[14][170],u_xpb_out[15][170],u_xpb_out[16][170],u_xpb_out[17][170],u_xpb_out[18][170],u_xpb_out[19][170],u_xpb_out[20][170],u_xpb_out[21][170],u_xpb_out[22][170],u_xpb_out[23][170],u_xpb_out[24][170],u_xpb_out[25][170],u_xpb_out[26][170],u_xpb_out[27][170],u_xpb_out[28][170],u_xpb_out[29][170],u_xpb_out[30][170],u_xpb_out[31][170],u_xpb_out[32][170],u_xpb_out[33][170],u_xpb_out[34][170],u_xpb_out[35][170],u_xpb_out[36][170],u_xpb_out[37][170],u_xpb_out[38][170],u_xpb_out[39][170],u_xpb_out[40][170],u_xpb_out[41][170],u_xpb_out[42][170],u_xpb_out[43][170],u_xpb_out[44][170],u_xpb_out[45][170],u_xpb_out[46][170],u_xpb_out[47][170],u_xpb_out[48][170],u_xpb_out[49][170],u_xpb_out[50][170],u_xpb_out[51][170],u_xpb_out[52][170],u_xpb_out[53][170],u_xpb_out[54][170],u_xpb_out[55][170],u_xpb_out[56][170],u_xpb_out[57][170],u_xpb_out[58][170],u_xpb_out[59][170],u_xpb_out[60][170],u_xpb_out[61][170],u_xpb_out[62][170],u_xpb_out[63][170],u_xpb_out[64][170],u_xpb_out[65][170],u_xpb_out[66][170],u_xpb_out[67][170],u_xpb_out[68][170],u_xpb_out[69][170],u_xpb_out[70][170],u_xpb_out[71][170],u_xpb_out[72][170],u_xpb_out[73][170],u_xpb_out[74][170],u_xpb_out[75][170],u_xpb_out[76][170],u_xpb_out[77][170],u_xpb_out[78][170],u_xpb_out[79][170],u_xpb_out[80][170],u_xpb_out[81][170],u_xpb_out[82][170],u_xpb_out[83][170],u_xpb_out[84][170],u_xpb_out[85][170],u_xpb_out[86][170],u_xpb_out[87][170],u_xpb_out[88][170],u_xpb_out[89][170],u_xpb_out[90][170],u_xpb_out[91][170],u_xpb_out[92][170],u_xpb_out[93][170],u_xpb_out[94][170],u_xpb_out[95][170],u_xpb_out[96][170],u_xpb_out[97][170],u_xpb_out[98][170],u_xpb_out[99][170],u_xpb_out[100][170],u_xpb_out[101][170],u_xpb_out[102][170],u_xpb_out[103][170],u_xpb_out[104][170],u_xpb_out[105][170]};

assign col_out_171 = {u_xpb_out[0][171],u_xpb_out[1][171],u_xpb_out[2][171],u_xpb_out[3][171],u_xpb_out[4][171],u_xpb_out[5][171],u_xpb_out[6][171],u_xpb_out[7][171],u_xpb_out[8][171],u_xpb_out[9][171],u_xpb_out[10][171],u_xpb_out[11][171],u_xpb_out[12][171],u_xpb_out[13][171],u_xpb_out[14][171],u_xpb_out[15][171],u_xpb_out[16][171],u_xpb_out[17][171],u_xpb_out[18][171],u_xpb_out[19][171],u_xpb_out[20][171],u_xpb_out[21][171],u_xpb_out[22][171],u_xpb_out[23][171],u_xpb_out[24][171],u_xpb_out[25][171],u_xpb_out[26][171],u_xpb_out[27][171],u_xpb_out[28][171],u_xpb_out[29][171],u_xpb_out[30][171],u_xpb_out[31][171],u_xpb_out[32][171],u_xpb_out[33][171],u_xpb_out[34][171],u_xpb_out[35][171],u_xpb_out[36][171],u_xpb_out[37][171],u_xpb_out[38][171],u_xpb_out[39][171],u_xpb_out[40][171],u_xpb_out[41][171],u_xpb_out[42][171],u_xpb_out[43][171],u_xpb_out[44][171],u_xpb_out[45][171],u_xpb_out[46][171],u_xpb_out[47][171],u_xpb_out[48][171],u_xpb_out[49][171],u_xpb_out[50][171],u_xpb_out[51][171],u_xpb_out[52][171],u_xpb_out[53][171],u_xpb_out[54][171],u_xpb_out[55][171],u_xpb_out[56][171],u_xpb_out[57][171],u_xpb_out[58][171],u_xpb_out[59][171],u_xpb_out[60][171],u_xpb_out[61][171],u_xpb_out[62][171],u_xpb_out[63][171],u_xpb_out[64][171],u_xpb_out[65][171],u_xpb_out[66][171],u_xpb_out[67][171],u_xpb_out[68][171],u_xpb_out[69][171],u_xpb_out[70][171],u_xpb_out[71][171],u_xpb_out[72][171],u_xpb_out[73][171],u_xpb_out[74][171],u_xpb_out[75][171],u_xpb_out[76][171],u_xpb_out[77][171],u_xpb_out[78][171],u_xpb_out[79][171],u_xpb_out[80][171],u_xpb_out[81][171],u_xpb_out[82][171],u_xpb_out[83][171],u_xpb_out[84][171],u_xpb_out[85][171],u_xpb_out[86][171],u_xpb_out[87][171],u_xpb_out[88][171],u_xpb_out[89][171],u_xpb_out[90][171],u_xpb_out[91][171],u_xpb_out[92][171],u_xpb_out[93][171],u_xpb_out[94][171],u_xpb_out[95][171],u_xpb_out[96][171],u_xpb_out[97][171],u_xpb_out[98][171],u_xpb_out[99][171],u_xpb_out[100][171],u_xpb_out[101][171],u_xpb_out[102][171],u_xpb_out[103][171],u_xpb_out[104][171],u_xpb_out[105][171]};

assign col_out_172 = {u_xpb_out[0][172],u_xpb_out[1][172],u_xpb_out[2][172],u_xpb_out[3][172],u_xpb_out[4][172],u_xpb_out[5][172],u_xpb_out[6][172],u_xpb_out[7][172],u_xpb_out[8][172],u_xpb_out[9][172],u_xpb_out[10][172],u_xpb_out[11][172],u_xpb_out[12][172],u_xpb_out[13][172],u_xpb_out[14][172],u_xpb_out[15][172],u_xpb_out[16][172],u_xpb_out[17][172],u_xpb_out[18][172],u_xpb_out[19][172],u_xpb_out[20][172],u_xpb_out[21][172],u_xpb_out[22][172],u_xpb_out[23][172],u_xpb_out[24][172],u_xpb_out[25][172],u_xpb_out[26][172],u_xpb_out[27][172],u_xpb_out[28][172],u_xpb_out[29][172],u_xpb_out[30][172],u_xpb_out[31][172],u_xpb_out[32][172],u_xpb_out[33][172],u_xpb_out[34][172],u_xpb_out[35][172],u_xpb_out[36][172],u_xpb_out[37][172],u_xpb_out[38][172],u_xpb_out[39][172],u_xpb_out[40][172],u_xpb_out[41][172],u_xpb_out[42][172],u_xpb_out[43][172],u_xpb_out[44][172],u_xpb_out[45][172],u_xpb_out[46][172],u_xpb_out[47][172],u_xpb_out[48][172],u_xpb_out[49][172],u_xpb_out[50][172],u_xpb_out[51][172],u_xpb_out[52][172],u_xpb_out[53][172],u_xpb_out[54][172],u_xpb_out[55][172],u_xpb_out[56][172],u_xpb_out[57][172],u_xpb_out[58][172],u_xpb_out[59][172],u_xpb_out[60][172],u_xpb_out[61][172],u_xpb_out[62][172],u_xpb_out[63][172],u_xpb_out[64][172],u_xpb_out[65][172],u_xpb_out[66][172],u_xpb_out[67][172],u_xpb_out[68][172],u_xpb_out[69][172],u_xpb_out[70][172],u_xpb_out[71][172],u_xpb_out[72][172],u_xpb_out[73][172],u_xpb_out[74][172],u_xpb_out[75][172],u_xpb_out[76][172],u_xpb_out[77][172],u_xpb_out[78][172],u_xpb_out[79][172],u_xpb_out[80][172],u_xpb_out[81][172],u_xpb_out[82][172],u_xpb_out[83][172],u_xpb_out[84][172],u_xpb_out[85][172],u_xpb_out[86][172],u_xpb_out[87][172],u_xpb_out[88][172],u_xpb_out[89][172],u_xpb_out[90][172],u_xpb_out[91][172],u_xpb_out[92][172],u_xpb_out[93][172],u_xpb_out[94][172],u_xpb_out[95][172],u_xpb_out[96][172],u_xpb_out[97][172],u_xpb_out[98][172],u_xpb_out[99][172],u_xpb_out[100][172],u_xpb_out[101][172],u_xpb_out[102][172],u_xpb_out[103][172],u_xpb_out[104][172],u_xpb_out[105][172]};

assign col_out_173 = {u_xpb_out[0][173],u_xpb_out[1][173],u_xpb_out[2][173],u_xpb_out[3][173],u_xpb_out[4][173],u_xpb_out[5][173],u_xpb_out[6][173],u_xpb_out[7][173],u_xpb_out[8][173],u_xpb_out[9][173],u_xpb_out[10][173],u_xpb_out[11][173],u_xpb_out[12][173],u_xpb_out[13][173],u_xpb_out[14][173],u_xpb_out[15][173],u_xpb_out[16][173],u_xpb_out[17][173],u_xpb_out[18][173],u_xpb_out[19][173],u_xpb_out[20][173],u_xpb_out[21][173],u_xpb_out[22][173],u_xpb_out[23][173],u_xpb_out[24][173],u_xpb_out[25][173],u_xpb_out[26][173],u_xpb_out[27][173],u_xpb_out[28][173],u_xpb_out[29][173],u_xpb_out[30][173],u_xpb_out[31][173],u_xpb_out[32][173],u_xpb_out[33][173],u_xpb_out[34][173],u_xpb_out[35][173],u_xpb_out[36][173],u_xpb_out[37][173],u_xpb_out[38][173],u_xpb_out[39][173],u_xpb_out[40][173],u_xpb_out[41][173],u_xpb_out[42][173],u_xpb_out[43][173],u_xpb_out[44][173],u_xpb_out[45][173],u_xpb_out[46][173],u_xpb_out[47][173],u_xpb_out[48][173],u_xpb_out[49][173],u_xpb_out[50][173],u_xpb_out[51][173],u_xpb_out[52][173],u_xpb_out[53][173],u_xpb_out[54][173],u_xpb_out[55][173],u_xpb_out[56][173],u_xpb_out[57][173],u_xpb_out[58][173],u_xpb_out[59][173],u_xpb_out[60][173],u_xpb_out[61][173],u_xpb_out[62][173],u_xpb_out[63][173],u_xpb_out[64][173],u_xpb_out[65][173],u_xpb_out[66][173],u_xpb_out[67][173],u_xpb_out[68][173],u_xpb_out[69][173],u_xpb_out[70][173],u_xpb_out[71][173],u_xpb_out[72][173],u_xpb_out[73][173],u_xpb_out[74][173],u_xpb_out[75][173],u_xpb_out[76][173],u_xpb_out[77][173],u_xpb_out[78][173],u_xpb_out[79][173],u_xpb_out[80][173],u_xpb_out[81][173],u_xpb_out[82][173],u_xpb_out[83][173],u_xpb_out[84][173],u_xpb_out[85][173],u_xpb_out[86][173],u_xpb_out[87][173],u_xpb_out[88][173],u_xpb_out[89][173],u_xpb_out[90][173],u_xpb_out[91][173],u_xpb_out[92][173],u_xpb_out[93][173],u_xpb_out[94][173],u_xpb_out[95][173],u_xpb_out[96][173],u_xpb_out[97][173],u_xpb_out[98][173],u_xpb_out[99][173],u_xpb_out[100][173],u_xpb_out[101][173],u_xpb_out[102][173],u_xpb_out[103][173],u_xpb_out[104][173],u_xpb_out[105][173]};

assign col_out_174 = {u_xpb_out[0][174],u_xpb_out[1][174],u_xpb_out[2][174],u_xpb_out[3][174],u_xpb_out[4][174],u_xpb_out[5][174],u_xpb_out[6][174],u_xpb_out[7][174],u_xpb_out[8][174],u_xpb_out[9][174],u_xpb_out[10][174],u_xpb_out[11][174],u_xpb_out[12][174],u_xpb_out[13][174],u_xpb_out[14][174],u_xpb_out[15][174],u_xpb_out[16][174],u_xpb_out[17][174],u_xpb_out[18][174],u_xpb_out[19][174],u_xpb_out[20][174],u_xpb_out[21][174],u_xpb_out[22][174],u_xpb_out[23][174],u_xpb_out[24][174],u_xpb_out[25][174],u_xpb_out[26][174],u_xpb_out[27][174],u_xpb_out[28][174],u_xpb_out[29][174],u_xpb_out[30][174],u_xpb_out[31][174],u_xpb_out[32][174],u_xpb_out[33][174],u_xpb_out[34][174],u_xpb_out[35][174],u_xpb_out[36][174],u_xpb_out[37][174],u_xpb_out[38][174],u_xpb_out[39][174],u_xpb_out[40][174],u_xpb_out[41][174],u_xpb_out[42][174],u_xpb_out[43][174],u_xpb_out[44][174],u_xpb_out[45][174],u_xpb_out[46][174],u_xpb_out[47][174],u_xpb_out[48][174],u_xpb_out[49][174],u_xpb_out[50][174],u_xpb_out[51][174],u_xpb_out[52][174],u_xpb_out[53][174],u_xpb_out[54][174],u_xpb_out[55][174],u_xpb_out[56][174],u_xpb_out[57][174],u_xpb_out[58][174],u_xpb_out[59][174],u_xpb_out[60][174],u_xpb_out[61][174],u_xpb_out[62][174],u_xpb_out[63][174],u_xpb_out[64][174],u_xpb_out[65][174],u_xpb_out[66][174],u_xpb_out[67][174],u_xpb_out[68][174],u_xpb_out[69][174],u_xpb_out[70][174],u_xpb_out[71][174],u_xpb_out[72][174],u_xpb_out[73][174],u_xpb_out[74][174],u_xpb_out[75][174],u_xpb_out[76][174],u_xpb_out[77][174],u_xpb_out[78][174],u_xpb_out[79][174],u_xpb_out[80][174],u_xpb_out[81][174],u_xpb_out[82][174],u_xpb_out[83][174],u_xpb_out[84][174],u_xpb_out[85][174],u_xpb_out[86][174],u_xpb_out[87][174],u_xpb_out[88][174],u_xpb_out[89][174],u_xpb_out[90][174],u_xpb_out[91][174],u_xpb_out[92][174],u_xpb_out[93][174],u_xpb_out[94][174],u_xpb_out[95][174],u_xpb_out[96][174],u_xpb_out[97][174],u_xpb_out[98][174],u_xpb_out[99][174],u_xpb_out[100][174],u_xpb_out[101][174],u_xpb_out[102][174],u_xpb_out[103][174],u_xpb_out[104][174],u_xpb_out[105][174]};

assign col_out_175 = {u_xpb_out[0][175],u_xpb_out[1][175],u_xpb_out[2][175],u_xpb_out[3][175],u_xpb_out[4][175],u_xpb_out[5][175],u_xpb_out[6][175],u_xpb_out[7][175],u_xpb_out[8][175],u_xpb_out[9][175],u_xpb_out[10][175],u_xpb_out[11][175],u_xpb_out[12][175],u_xpb_out[13][175],u_xpb_out[14][175],u_xpb_out[15][175],u_xpb_out[16][175],u_xpb_out[17][175],u_xpb_out[18][175],u_xpb_out[19][175],u_xpb_out[20][175],u_xpb_out[21][175],u_xpb_out[22][175],u_xpb_out[23][175],u_xpb_out[24][175],u_xpb_out[25][175],u_xpb_out[26][175],u_xpb_out[27][175],u_xpb_out[28][175],u_xpb_out[29][175],u_xpb_out[30][175],u_xpb_out[31][175],u_xpb_out[32][175],u_xpb_out[33][175],u_xpb_out[34][175],u_xpb_out[35][175],u_xpb_out[36][175],u_xpb_out[37][175],u_xpb_out[38][175],u_xpb_out[39][175],u_xpb_out[40][175],u_xpb_out[41][175],u_xpb_out[42][175],u_xpb_out[43][175],u_xpb_out[44][175],u_xpb_out[45][175],u_xpb_out[46][175],u_xpb_out[47][175],u_xpb_out[48][175],u_xpb_out[49][175],u_xpb_out[50][175],u_xpb_out[51][175],u_xpb_out[52][175],u_xpb_out[53][175],u_xpb_out[54][175],u_xpb_out[55][175],u_xpb_out[56][175],u_xpb_out[57][175],u_xpb_out[58][175],u_xpb_out[59][175],u_xpb_out[60][175],u_xpb_out[61][175],u_xpb_out[62][175],u_xpb_out[63][175],u_xpb_out[64][175],u_xpb_out[65][175],u_xpb_out[66][175],u_xpb_out[67][175],u_xpb_out[68][175],u_xpb_out[69][175],u_xpb_out[70][175],u_xpb_out[71][175],u_xpb_out[72][175],u_xpb_out[73][175],u_xpb_out[74][175],u_xpb_out[75][175],u_xpb_out[76][175],u_xpb_out[77][175],u_xpb_out[78][175],u_xpb_out[79][175],u_xpb_out[80][175],u_xpb_out[81][175],u_xpb_out[82][175],u_xpb_out[83][175],u_xpb_out[84][175],u_xpb_out[85][175],u_xpb_out[86][175],u_xpb_out[87][175],u_xpb_out[88][175],u_xpb_out[89][175],u_xpb_out[90][175],u_xpb_out[91][175],u_xpb_out[92][175],u_xpb_out[93][175],u_xpb_out[94][175],u_xpb_out[95][175],u_xpb_out[96][175],u_xpb_out[97][175],u_xpb_out[98][175],u_xpb_out[99][175],u_xpb_out[100][175],u_xpb_out[101][175],u_xpb_out[102][175],u_xpb_out[103][175],u_xpb_out[104][175],u_xpb_out[105][175]};

assign col_out_176 = {u_xpb_out[0][176],u_xpb_out[1][176],u_xpb_out[2][176],u_xpb_out[3][176],u_xpb_out[4][176],u_xpb_out[5][176],u_xpb_out[6][176],u_xpb_out[7][176],u_xpb_out[8][176],u_xpb_out[9][176],u_xpb_out[10][176],u_xpb_out[11][176],u_xpb_out[12][176],u_xpb_out[13][176],u_xpb_out[14][176],u_xpb_out[15][176],u_xpb_out[16][176],u_xpb_out[17][176],u_xpb_out[18][176],u_xpb_out[19][176],u_xpb_out[20][176],u_xpb_out[21][176],u_xpb_out[22][176],u_xpb_out[23][176],u_xpb_out[24][176],u_xpb_out[25][176],u_xpb_out[26][176],u_xpb_out[27][176],u_xpb_out[28][176],u_xpb_out[29][176],u_xpb_out[30][176],u_xpb_out[31][176],u_xpb_out[32][176],u_xpb_out[33][176],u_xpb_out[34][176],u_xpb_out[35][176],u_xpb_out[36][176],u_xpb_out[37][176],u_xpb_out[38][176],u_xpb_out[39][176],u_xpb_out[40][176],u_xpb_out[41][176],u_xpb_out[42][176],u_xpb_out[43][176],u_xpb_out[44][176],u_xpb_out[45][176],u_xpb_out[46][176],u_xpb_out[47][176],u_xpb_out[48][176],u_xpb_out[49][176],u_xpb_out[50][176],u_xpb_out[51][176],u_xpb_out[52][176],u_xpb_out[53][176],u_xpb_out[54][176],u_xpb_out[55][176],u_xpb_out[56][176],u_xpb_out[57][176],u_xpb_out[58][176],u_xpb_out[59][176],u_xpb_out[60][176],u_xpb_out[61][176],u_xpb_out[62][176],u_xpb_out[63][176],u_xpb_out[64][176],u_xpb_out[65][176],u_xpb_out[66][176],u_xpb_out[67][176],u_xpb_out[68][176],u_xpb_out[69][176],u_xpb_out[70][176],u_xpb_out[71][176],u_xpb_out[72][176],u_xpb_out[73][176],u_xpb_out[74][176],u_xpb_out[75][176],u_xpb_out[76][176],u_xpb_out[77][176],u_xpb_out[78][176],u_xpb_out[79][176],u_xpb_out[80][176],u_xpb_out[81][176],u_xpb_out[82][176],u_xpb_out[83][176],u_xpb_out[84][176],u_xpb_out[85][176],u_xpb_out[86][176],u_xpb_out[87][176],u_xpb_out[88][176],u_xpb_out[89][176],u_xpb_out[90][176],u_xpb_out[91][176],u_xpb_out[92][176],u_xpb_out[93][176],u_xpb_out[94][176],u_xpb_out[95][176],u_xpb_out[96][176],u_xpb_out[97][176],u_xpb_out[98][176],u_xpb_out[99][176],u_xpb_out[100][176],u_xpb_out[101][176],u_xpb_out[102][176],u_xpb_out[103][176],u_xpb_out[104][176],u_xpb_out[105][176]};

assign col_out_177 = {u_xpb_out[0][177],u_xpb_out[1][177],u_xpb_out[2][177],u_xpb_out[3][177],u_xpb_out[4][177],u_xpb_out[5][177],u_xpb_out[6][177],u_xpb_out[7][177],u_xpb_out[8][177],u_xpb_out[9][177],u_xpb_out[10][177],u_xpb_out[11][177],u_xpb_out[12][177],u_xpb_out[13][177],u_xpb_out[14][177],u_xpb_out[15][177],u_xpb_out[16][177],u_xpb_out[17][177],u_xpb_out[18][177],u_xpb_out[19][177],u_xpb_out[20][177],u_xpb_out[21][177],u_xpb_out[22][177],u_xpb_out[23][177],u_xpb_out[24][177],u_xpb_out[25][177],u_xpb_out[26][177],u_xpb_out[27][177],u_xpb_out[28][177],u_xpb_out[29][177],u_xpb_out[30][177],u_xpb_out[31][177],u_xpb_out[32][177],u_xpb_out[33][177],u_xpb_out[34][177],u_xpb_out[35][177],u_xpb_out[36][177],u_xpb_out[37][177],u_xpb_out[38][177],u_xpb_out[39][177],u_xpb_out[40][177],u_xpb_out[41][177],u_xpb_out[42][177],u_xpb_out[43][177],u_xpb_out[44][177],u_xpb_out[45][177],u_xpb_out[46][177],u_xpb_out[47][177],u_xpb_out[48][177],u_xpb_out[49][177],u_xpb_out[50][177],u_xpb_out[51][177],u_xpb_out[52][177],u_xpb_out[53][177],u_xpb_out[54][177],u_xpb_out[55][177],u_xpb_out[56][177],u_xpb_out[57][177],u_xpb_out[58][177],u_xpb_out[59][177],u_xpb_out[60][177],u_xpb_out[61][177],u_xpb_out[62][177],u_xpb_out[63][177],u_xpb_out[64][177],u_xpb_out[65][177],u_xpb_out[66][177],u_xpb_out[67][177],u_xpb_out[68][177],u_xpb_out[69][177],u_xpb_out[70][177],u_xpb_out[71][177],u_xpb_out[72][177],u_xpb_out[73][177],u_xpb_out[74][177],u_xpb_out[75][177],u_xpb_out[76][177],u_xpb_out[77][177],u_xpb_out[78][177],u_xpb_out[79][177],u_xpb_out[80][177],u_xpb_out[81][177],u_xpb_out[82][177],u_xpb_out[83][177],u_xpb_out[84][177],u_xpb_out[85][177],u_xpb_out[86][177],u_xpb_out[87][177],u_xpb_out[88][177],u_xpb_out[89][177],u_xpb_out[90][177],u_xpb_out[91][177],u_xpb_out[92][177],u_xpb_out[93][177],u_xpb_out[94][177],u_xpb_out[95][177],u_xpb_out[96][177],u_xpb_out[97][177],u_xpb_out[98][177],u_xpb_out[99][177],u_xpb_out[100][177],u_xpb_out[101][177],u_xpb_out[102][177],u_xpb_out[103][177],u_xpb_out[104][177],u_xpb_out[105][177]};

assign col_out_178 = {u_xpb_out[0][178],u_xpb_out[1][178],u_xpb_out[2][178],u_xpb_out[3][178],u_xpb_out[4][178],u_xpb_out[5][178],u_xpb_out[6][178],u_xpb_out[7][178],u_xpb_out[8][178],u_xpb_out[9][178],u_xpb_out[10][178],u_xpb_out[11][178],u_xpb_out[12][178],u_xpb_out[13][178],u_xpb_out[14][178],u_xpb_out[15][178],u_xpb_out[16][178],u_xpb_out[17][178],u_xpb_out[18][178],u_xpb_out[19][178],u_xpb_out[20][178],u_xpb_out[21][178],u_xpb_out[22][178],u_xpb_out[23][178],u_xpb_out[24][178],u_xpb_out[25][178],u_xpb_out[26][178],u_xpb_out[27][178],u_xpb_out[28][178],u_xpb_out[29][178],u_xpb_out[30][178],u_xpb_out[31][178],u_xpb_out[32][178],u_xpb_out[33][178],u_xpb_out[34][178],u_xpb_out[35][178],u_xpb_out[36][178],u_xpb_out[37][178],u_xpb_out[38][178],u_xpb_out[39][178],u_xpb_out[40][178],u_xpb_out[41][178],u_xpb_out[42][178],u_xpb_out[43][178],u_xpb_out[44][178],u_xpb_out[45][178],u_xpb_out[46][178],u_xpb_out[47][178],u_xpb_out[48][178],u_xpb_out[49][178],u_xpb_out[50][178],u_xpb_out[51][178],u_xpb_out[52][178],u_xpb_out[53][178],u_xpb_out[54][178],u_xpb_out[55][178],u_xpb_out[56][178],u_xpb_out[57][178],u_xpb_out[58][178],u_xpb_out[59][178],u_xpb_out[60][178],u_xpb_out[61][178],u_xpb_out[62][178],u_xpb_out[63][178],u_xpb_out[64][178],u_xpb_out[65][178],u_xpb_out[66][178],u_xpb_out[67][178],u_xpb_out[68][178],u_xpb_out[69][178],u_xpb_out[70][178],u_xpb_out[71][178],u_xpb_out[72][178],u_xpb_out[73][178],u_xpb_out[74][178],u_xpb_out[75][178],u_xpb_out[76][178],u_xpb_out[77][178],u_xpb_out[78][178],u_xpb_out[79][178],u_xpb_out[80][178],u_xpb_out[81][178],u_xpb_out[82][178],u_xpb_out[83][178],u_xpb_out[84][178],u_xpb_out[85][178],u_xpb_out[86][178],u_xpb_out[87][178],u_xpb_out[88][178],u_xpb_out[89][178],u_xpb_out[90][178],u_xpb_out[91][178],u_xpb_out[92][178],u_xpb_out[93][178],u_xpb_out[94][178],u_xpb_out[95][178],u_xpb_out[96][178],u_xpb_out[97][178],u_xpb_out[98][178],u_xpb_out[99][178],u_xpb_out[100][178],u_xpb_out[101][178],u_xpb_out[102][178],u_xpb_out[103][178],u_xpb_out[104][178],u_xpb_out[105][178]};

assign col_out_179 = {u_xpb_out[0][179],u_xpb_out[1][179],u_xpb_out[2][179],u_xpb_out[3][179],u_xpb_out[4][179],u_xpb_out[5][179],u_xpb_out[6][179],u_xpb_out[7][179],u_xpb_out[8][179],u_xpb_out[9][179],u_xpb_out[10][179],u_xpb_out[11][179],u_xpb_out[12][179],u_xpb_out[13][179],u_xpb_out[14][179],u_xpb_out[15][179],u_xpb_out[16][179],u_xpb_out[17][179],u_xpb_out[18][179],u_xpb_out[19][179],u_xpb_out[20][179],u_xpb_out[21][179],u_xpb_out[22][179],u_xpb_out[23][179],u_xpb_out[24][179],u_xpb_out[25][179],u_xpb_out[26][179],u_xpb_out[27][179],u_xpb_out[28][179],u_xpb_out[29][179],u_xpb_out[30][179],u_xpb_out[31][179],u_xpb_out[32][179],u_xpb_out[33][179],u_xpb_out[34][179],u_xpb_out[35][179],u_xpb_out[36][179],u_xpb_out[37][179],u_xpb_out[38][179],u_xpb_out[39][179],u_xpb_out[40][179],u_xpb_out[41][179],u_xpb_out[42][179],u_xpb_out[43][179],u_xpb_out[44][179],u_xpb_out[45][179],u_xpb_out[46][179],u_xpb_out[47][179],u_xpb_out[48][179],u_xpb_out[49][179],u_xpb_out[50][179],u_xpb_out[51][179],u_xpb_out[52][179],u_xpb_out[53][179],u_xpb_out[54][179],u_xpb_out[55][179],u_xpb_out[56][179],u_xpb_out[57][179],u_xpb_out[58][179],u_xpb_out[59][179],u_xpb_out[60][179],u_xpb_out[61][179],u_xpb_out[62][179],u_xpb_out[63][179],u_xpb_out[64][179],u_xpb_out[65][179],u_xpb_out[66][179],u_xpb_out[67][179],u_xpb_out[68][179],u_xpb_out[69][179],u_xpb_out[70][179],u_xpb_out[71][179],u_xpb_out[72][179],u_xpb_out[73][179],u_xpb_out[74][179],u_xpb_out[75][179],u_xpb_out[76][179],u_xpb_out[77][179],u_xpb_out[78][179],u_xpb_out[79][179],u_xpb_out[80][179],u_xpb_out[81][179],u_xpb_out[82][179],u_xpb_out[83][179],u_xpb_out[84][179],u_xpb_out[85][179],u_xpb_out[86][179],u_xpb_out[87][179],u_xpb_out[88][179],u_xpb_out[89][179],u_xpb_out[90][179],u_xpb_out[91][179],u_xpb_out[92][179],u_xpb_out[93][179],u_xpb_out[94][179],u_xpb_out[95][179],u_xpb_out[96][179],u_xpb_out[97][179],u_xpb_out[98][179],u_xpb_out[99][179],u_xpb_out[100][179],u_xpb_out[101][179],u_xpb_out[102][179],u_xpb_out[103][179],u_xpb_out[104][179],u_xpb_out[105][179]};

assign col_out_180 = {u_xpb_out[0][180],u_xpb_out[1][180],u_xpb_out[2][180],u_xpb_out[3][180],u_xpb_out[4][180],u_xpb_out[5][180],u_xpb_out[6][180],u_xpb_out[7][180],u_xpb_out[8][180],u_xpb_out[9][180],u_xpb_out[10][180],u_xpb_out[11][180],u_xpb_out[12][180],u_xpb_out[13][180],u_xpb_out[14][180],u_xpb_out[15][180],u_xpb_out[16][180],u_xpb_out[17][180],u_xpb_out[18][180],u_xpb_out[19][180],u_xpb_out[20][180],u_xpb_out[21][180],u_xpb_out[22][180],u_xpb_out[23][180],u_xpb_out[24][180],u_xpb_out[25][180],u_xpb_out[26][180],u_xpb_out[27][180],u_xpb_out[28][180],u_xpb_out[29][180],u_xpb_out[30][180],u_xpb_out[31][180],u_xpb_out[32][180],u_xpb_out[33][180],u_xpb_out[34][180],u_xpb_out[35][180],u_xpb_out[36][180],u_xpb_out[37][180],u_xpb_out[38][180],u_xpb_out[39][180],u_xpb_out[40][180],u_xpb_out[41][180],u_xpb_out[42][180],u_xpb_out[43][180],u_xpb_out[44][180],u_xpb_out[45][180],u_xpb_out[46][180],u_xpb_out[47][180],u_xpb_out[48][180],u_xpb_out[49][180],u_xpb_out[50][180],u_xpb_out[51][180],u_xpb_out[52][180],u_xpb_out[53][180],u_xpb_out[54][180],u_xpb_out[55][180],u_xpb_out[56][180],u_xpb_out[57][180],u_xpb_out[58][180],u_xpb_out[59][180],u_xpb_out[60][180],u_xpb_out[61][180],u_xpb_out[62][180],u_xpb_out[63][180],u_xpb_out[64][180],u_xpb_out[65][180],u_xpb_out[66][180],u_xpb_out[67][180],u_xpb_out[68][180],u_xpb_out[69][180],u_xpb_out[70][180],u_xpb_out[71][180],u_xpb_out[72][180],u_xpb_out[73][180],u_xpb_out[74][180],u_xpb_out[75][180],u_xpb_out[76][180],u_xpb_out[77][180],u_xpb_out[78][180],u_xpb_out[79][180],u_xpb_out[80][180],u_xpb_out[81][180],u_xpb_out[82][180],u_xpb_out[83][180],u_xpb_out[84][180],u_xpb_out[85][180],u_xpb_out[86][180],u_xpb_out[87][180],u_xpb_out[88][180],u_xpb_out[89][180],u_xpb_out[90][180],u_xpb_out[91][180],u_xpb_out[92][180],u_xpb_out[93][180],u_xpb_out[94][180],u_xpb_out[95][180],u_xpb_out[96][180],u_xpb_out[97][180],u_xpb_out[98][180],u_xpb_out[99][180],u_xpb_out[100][180],u_xpb_out[101][180],u_xpb_out[102][180],u_xpb_out[103][180],u_xpb_out[104][180],u_xpb_out[105][180]};

assign col_out_181 = {u_xpb_out[0][181],u_xpb_out[1][181],u_xpb_out[2][181],u_xpb_out[3][181],u_xpb_out[4][181],u_xpb_out[5][181],u_xpb_out[6][181],u_xpb_out[7][181],u_xpb_out[8][181],u_xpb_out[9][181],u_xpb_out[10][181],u_xpb_out[11][181],u_xpb_out[12][181],u_xpb_out[13][181],u_xpb_out[14][181],u_xpb_out[15][181],u_xpb_out[16][181],u_xpb_out[17][181],u_xpb_out[18][181],u_xpb_out[19][181],u_xpb_out[20][181],u_xpb_out[21][181],u_xpb_out[22][181],u_xpb_out[23][181],u_xpb_out[24][181],u_xpb_out[25][181],u_xpb_out[26][181],u_xpb_out[27][181],u_xpb_out[28][181],u_xpb_out[29][181],u_xpb_out[30][181],u_xpb_out[31][181],u_xpb_out[32][181],u_xpb_out[33][181],u_xpb_out[34][181],u_xpb_out[35][181],u_xpb_out[36][181],u_xpb_out[37][181],u_xpb_out[38][181],u_xpb_out[39][181],u_xpb_out[40][181],u_xpb_out[41][181],u_xpb_out[42][181],u_xpb_out[43][181],u_xpb_out[44][181],u_xpb_out[45][181],u_xpb_out[46][181],u_xpb_out[47][181],u_xpb_out[48][181],u_xpb_out[49][181],u_xpb_out[50][181],u_xpb_out[51][181],u_xpb_out[52][181],u_xpb_out[53][181],u_xpb_out[54][181],u_xpb_out[55][181],u_xpb_out[56][181],u_xpb_out[57][181],u_xpb_out[58][181],u_xpb_out[59][181],u_xpb_out[60][181],u_xpb_out[61][181],u_xpb_out[62][181],u_xpb_out[63][181],u_xpb_out[64][181],u_xpb_out[65][181],u_xpb_out[66][181],u_xpb_out[67][181],u_xpb_out[68][181],u_xpb_out[69][181],u_xpb_out[70][181],u_xpb_out[71][181],u_xpb_out[72][181],u_xpb_out[73][181],u_xpb_out[74][181],u_xpb_out[75][181],u_xpb_out[76][181],u_xpb_out[77][181],u_xpb_out[78][181],u_xpb_out[79][181],u_xpb_out[80][181],u_xpb_out[81][181],u_xpb_out[82][181],u_xpb_out[83][181],u_xpb_out[84][181],u_xpb_out[85][181],u_xpb_out[86][181],u_xpb_out[87][181],u_xpb_out[88][181],u_xpb_out[89][181],u_xpb_out[90][181],u_xpb_out[91][181],u_xpb_out[92][181],u_xpb_out[93][181],u_xpb_out[94][181],u_xpb_out[95][181],u_xpb_out[96][181],u_xpb_out[97][181],u_xpb_out[98][181],u_xpb_out[99][181],u_xpb_out[100][181],u_xpb_out[101][181],u_xpb_out[102][181],u_xpb_out[103][181],u_xpb_out[104][181],u_xpb_out[105][181]};

assign col_out_182 = {u_xpb_out[0][182],u_xpb_out[1][182],u_xpb_out[2][182],u_xpb_out[3][182],u_xpb_out[4][182],u_xpb_out[5][182],u_xpb_out[6][182],u_xpb_out[7][182],u_xpb_out[8][182],u_xpb_out[9][182],u_xpb_out[10][182],u_xpb_out[11][182],u_xpb_out[12][182],u_xpb_out[13][182],u_xpb_out[14][182],u_xpb_out[15][182],u_xpb_out[16][182],u_xpb_out[17][182],u_xpb_out[18][182],u_xpb_out[19][182],u_xpb_out[20][182],u_xpb_out[21][182],u_xpb_out[22][182],u_xpb_out[23][182],u_xpb_out[24][182],u_xpb_out[25][182],u_xpb_out[26][182],u_xpb_out[27][182],u_xpb_out[28][182],u_xpb_out[29][182],u_xpb_out[30][182],u_xpb_out[31][182],u_xpb_out[32][182],u_xpb_out[33][182],u_xpb_out[34][182],u_xpb_out[35][182],u_xpb_out[36][182],u_xpb_out[37][182],u_xpb_out[38][182],u_xpb_out[39][182],u_xpb_out[40][182],u_xpb_out[41][182],u_xpb_out[42][182],u_xpb_out[43][182],u_xpb_out[44][182],u_xpb_out[45][182],u_xpb_out[46][182],u_xpb_out[47][182],u_xpb_out[48][182],u_xpb_out[49][182],u_xpb_out[50][182],u_xpb_out[51][182],u_xpb_out[52][182],u_xpb_out[53][182],u_xpb_out[54][182],u_xpb_out[55][182],u_xpb_out[56][182],u_xpb_out[57][182],u_xpb_out[58][182],u_xpb_out[59][182],u_xpb_out[60][182],u_xpb_out[61][182],u_xpb_out[62][182],u_xpb_out[63][182],u_xpb_out[64][182],u_xpb_out[65][182],u_xpb_out[66][182],u_xpb_out[67][182],u_xpb_out[68][182],u_xpb_out[69][182],u_xpb_out[70][182],u_xpb_out[71][182],u_xpb_out[72][182],u_xpb_out[73][182],u_xpb_out[74][182],u_xpb_out[75][182],u_xpb_out[76][182],u_xpb_out[77][182],u_xpb_out[78][182],u_xpb_out[79][182],u_xpb_out[80][182],u_xpb_out[81][182],u_xpb_out[82][182],u_xpb_out[83][182],u_xpb_out[84][182],u_xpb_out[85][182],u_xpb_out[86][182],u_xpb_out[87][182],u_xpb_out[88][182],u_xpb_out[89][182],u_xpb_out[90][182],u_xpb_out[91][182],u_xpb_out[92][182],u_xpb_out[93][182],u_xpb_out[94][182],u_xpb_out[95][182],u_xpb_out[96][182],u_xpb_out[97][182],u_xpb_out[98][182],u_xpb_out[99][182],u_xpb_out[100][182],u_xpb_out[101][182],u_xpb_out[102][182],u_xpb_out[103][182],u_xpb_out[104][182],u_xpb_out[105][182]};

assign col_out_183 = {u_xpb_out[0][183],u_xpb_out[1][183],u_xpb_out[2][183],u_xpb_out[3][183],u_xpb_out[4][183],u_xpb_out[5][183],u_xpb_out[6][183],u_xpb_out[7][183],u_xpb_out[8][183],u_xpb_out[9][183],u_xpb_out[10][183],u_xpb_out[11][183],u_xpb_out[12][183],u_xpb_out[13][183],u_xpb_out[14][183],u_xpb_out[15][183],u_xpb_out[16][183],u_xpb_out[17][183],u_xpb_out[18][183],u_xpb_out[19][183],u_xpb_out[20][183],u_xpb_out[21][183],u_xpb_out[22][183],u_xpb_out[23][183],u_xpb_out[24][183],u_xpb_out[25][183],u_xpb_out[26][183],u_xpb_out[27][183],u_xpb_out[28][183],u_xpb_out[29][183],u_xpb_out[30][183],u_xpb_out[31][183],u_xpb_out[32][183],u_xpb_out[33][183],u_xpb_out[34][183],u_xpb_out[35][183],u_xpb_out[36][183],u_xpb_out[37][183],u_xpb_out[38][183],u_xpb_out[39][183],u_xpb_out[40][183],u_xpb_out[41][183],u_xpb_out[42][183],u_xpb_out[43][183],u_xpb_out[44][183],u_xpb_out[45][183],u_xpb_out[46][183],u_xpb_out[47][183],u_xpb_out[48][183],u_xpb_out[49][183],u_xpb_out[50][183],u_xpb_out[51][183],u_xpb_out[52][183],u_xpb_out[53][183],u_xpb_out[54][183],u_xpb_out[55][183],u_xpb_out[56][183],u_xpb_out[57][183],u_xpb_out[58][183],u_xpb_out[59][183],u_xpb_out[60][183],u_xpb_out[61][183],u_xpb_out[62][183],u_xpb_out[63][183],u_xpb_out[64][183],u_xpb_out[65][183],u_xpb_out[66][183],u_xpb_out[67][183],u_xpb_out[68][183],u_xpb_out[69][183],u_xpb_out[70][183],u_xpb_out[71][183],u_xpb_out[72][183],u_xpb_out[73][183],u_xpb_out[74][183],u_xpb_out[75][183],u_xpb_out[76][183],u_xpb_out[77][183],u_xpb_out[78][183],u_xpb_out[79][183],u_xpb_out[80][183],u_xpb_out[81][183],u_xpb_out[82][183],u_xpb_out[83][183],u_xpb_out[84][183],u_xpb_out[85][183],u_xpb_out[86][183],u_xpb_out[87][183],u_xpb_out[88][183],u_xpb_out[89][183],u_xpb_out[90][183],u_xpb_out[91][183],u_xpb_out[92][183],u_xpb_out[93][183],u_xpb_out[94][183],u_xpb_out[95][183],u_xpb_out[96][183],u_xpb_out[97][183],u_xpb_out[98][183],u_xpb_out[99][183],u_xpb_out[100][183],u_xpb_out[101][183],u_xpb_out[102][183],u_xpb_out[103][183],u_xpb_out[104][183],u_xpb_out[105][183]};

assign col_out_184 = {u_xpb_out[0][184],u_xpb_out[1][184],u_xpb_out[2][184],u_xpb_out[3][184],u_xpb_out[4][184],u_xpb_out[5][184],u_xpb_out[6][184],u_xpb_out[7][184],u_xpb_out[8][184],u_xpb_out[9][184],u_xpb_out[10][184],u_xpb_out[11][184],u_xpb_out[12][184],u_xpb_out[13][184],u_xpb_out[14][184],u_xpb_out[15][184],u_xpb_out[16][184],u_xpb_out[17][184],u_xpb_out[18][184],u_xpb_out[19][184],u_xpb_out[20][184],u_xpb_out[21][184],u_xpb_out[22][184],u_xpb_out[23][184],u_xpb_out[24][184],u_xpb_out[25][184],u_xpb_out[26][184],u_xpb_out[27][184],u_xpb_out[28][184],u_xpb_out[29][184],u_xpb_out[30][184],u_xpb_out[31][184],u_xpb_out[32][184],u_xpb_out[33][184],u_xpb_out[34][184],u_xpb_out[35][184],u_xpb_out[36][184],u_xpb_out[37][184],u_xpb_out[38][184],u_xpb_out[39][184],u_xpb_out[40][184],u_xpb_out[41][184],u_xpb_out[42][184],u_xpb_out[43][184],u_xpb_out[44][184],u_xpb_out[45][184],u_xpb_out[46][184],u_xpb_out[47][184],u_xpb_out[48][184],u_xpb_out[49][184],u_xpb_out[50][184],u_xpb_out[51][184],u_xpb_out[52][184],u_xpb_out[53][184],u_xpb_out[54][184],u_xpb_out[55][184],u_xpb_out[56][184],u_xpb_out[57][184],u_xpb_out[58][184],u_xpb_out[59][184],u_xpb_out[60][184],u_xpb_out[61][184],u_xpb_out[62][184],u_xpb_out[63][184],u_xpb_out[64][184],u_xpb_out[65][184],u_xpb_out[66][184],u_xpb_out[67][184],u_xpb_out[68][184],u_xpb_out[69][184],u_xpb_out[70][184],u_xpb_out[71][184],u_xpb_out[72][184],u_xpb_out[73][184],u_xpb_out[74][184],u_xpb_out[75][184],u_xpb_out[76][184],u_xpb_out[77][184],u_xpb_out[78][184],u_xpb_out[79][184],u_xpb_out[80][184],u_xpb_out[81][184],u_xpb_out[82][184],u_xpb_out[83][184],u_xpb_out[84][184],u_xpb_out[85][184],u_xpb_out[86][184],u_xpb_out[87][184],u_xpb_out[88][184],u_xpb_out[89][184],u_xpb_out[90][184],u_xpb_out[91][184],u_xpb_out[92][184],u_xpb_out[93][184],u_xpb_out[94][184],u_xpb_out[95][184],u_xpb_out[96][184],u_xpb_out[97][184],u_xpb_out[98][184],u_xpb_out[99][184],u_xpb_out[100][184],u_xpb_out[101][184],u_xpb_out[102][184],u_xpb_out[103][184],u_xpb_out[104][184],u_xpb_out[105][184]};

assign col_out_185 = {u_xpb_out[0][185],u_xpb_out[1][185],u_xpb_out[2][185],u_xpb_out[3][185],u_xpb_out[4][185],u_xpb_out[5][185],u_xpb_out[6][185],u_xpb_out[7][185],u_xpb_out[8][185],u_xpb_out[9][185],u_xpb_out[10][185],u_xpb_out[11][185],u_xpb_out[12][185],u_xpb_out[13][185],u_xpb_out[14][185],u_xpb_out[15][185],u_xpb_out[16][185],u_xpb_out[17][185],u_xpb_out[18][185],u_xpb_out[19][185],u_xpb_out[20][185],u_xpb_out[21][185],u_xpb_out[22][185],u_xpb_out[23][185],u_xpb_out[24][185],u_xpb_out[25][185],u_xpb_out[26][185],u_xpb_out[27][185],u_xpb_out[28][185],u_xpb_out[29][185],u_xpb_out[30][185],u_xpb_out[31][185],u_xpb_out[32][185],u_xpb_out[33][185],u_xpb_out[34][185],u_xpb_out[35][185],u_xpb_out[36][185],u_xpb_out[37][185],u_xpb_out[38][185],u_xpb_out[39][185],u_xpb_out[40][185],u_xpb_out[41][185],u_xpb_out[42][185],u_xpb_out[43][185],u_xpb_out[44][185],u_xpb_out[45][185],u_xpb_out[46][185],u_xpb_out[47][185],u_xpb_out[48][185],u_xpb_out[49][185],u_xpb_out[50][185],u_xpb_out[51][185],u_xpb_out[52][185],u_xpb_out[53][185],u_xpb_out[54][185],u_xpb_out[55][185],u_xpb_out[56][185],u_xpb_out[57][185],u_xpb_out[58][185],u_xpb_out[59][185],u_xpb_out[60][185],u_xpb_out[61][185],u_xpb_out[62][185],u_xpb_out[63][185],u_xpb_out[64][185],u_xpb_out[65][185],u_xpb_out[66][185],u_xpb_out[67][185],u_xpb_out[68][185],u_xpb_out[69][185],u_xpb_out[70][185],u_xpb_out[71][185],u_xpb_out[72][185],u_xpb_out[73][185],u_xpb_out[74][185],u_xpb_out[75][185],u_xpb_out[76][185],u_xpb_out[77][185],u_xpb_out[78][185],u_xpb_out[79][185],u_xpb_out[80][185],u_xpb_out[81][185],u_xpb_out[82][185],u_xpb_out[83][185],u_xpb_out[84][185],u_xpb_out[85][185],u_xpb_out[86][185],u_xpb_out[87][185],u_xpb_out[88][185],u_xpb_out[89][185],u_xpb_out[90][185],u_xpb_out[91][185],u_xpb_out[92][185],u_xpb_out[93][185],u_xpb_out[94][185],u_xpb_out[95][185],u_xpb_out[96][185],u_xpb_out[97][185],u_xpb_out[98][185],u_xpb_out[99][185],u_xpb_out[100][185],u_xpb_out[101][185],u_xpb_out[102][185],u_xpb_out[103][185],u_xpb_out[104][185],u_xpb_out[105][185]};

assign col_out_186 = {u_xpb_out[0][186],u_xpb_out[1][186],u_xpb_out[2][186],u_xpb_out[3][186],u_xpb_out[4][186],u_xpb_out[5][186],u_xpb_out[6][186],u_xpb_out[7][186],u_xpb_out[8][186],u_xpb_out[9][186],u_xpb_out[10][186],u_xpb_out[11][186],u_xpb_out[12][186],u_xpb_out[13][186],u_xpb_out[14][186],u_xpb_out[15][186],u_xpb_out[16][186],u_xpb_out[17][186],u_xpb_out[18][186],u_xpb_out[19][186],u_xpb_out[20][186],u_xpb_out[21][186],u_xpb_out[22][186],u_xpb_out[23][186],u_xpb_out[24][186],u_xpb_out[25][186],u_xpb_out[26][186],u_xpb_out[27][186],u_xpb_out[28][186],u_xpb_out[29][186],u_xpb_out[30][186],u_xpb_out[31][186],u_xpb_out[32][186],u_xpb_out[33][186],u_xpb_out[34][186],u_xpb_out[35][186],u_xpb_out[36][186],u_xpb_out[37][186],u_xpb_out[38][186],u_xpb_out[39][186],u_xpb_out[40][186],u_xpb_out[41][186],u_xpb_out[42][186],u_xpb_out[43][186],u_xpb_out[44][186],u_xpb_out[45][186],u_xpb_out[46][186],u_xpb_out[47][186],u_xpb_out[48][186],u_xpb_out[49][186],u_xpb_out[50][186],u_xpb_out[51][186],u_xpb_out[52][186],u_xpb_out[53][186],u_xpb_out[54][186],u_xpb_out[55][186],u_xpb_out[56][186],u_xpb_out[57][186],u_xpb_out[58][186],u_xpb_out[59][186],u_xpb_out[60][186],u_xpb_out[61][186],u_xpb_out[62][186],u_xpb_out[63][186],u_xpb_out[64][186],u_xpb_out[65][186],u_xpb_out[66][186],u_xpb_out[67][186],u_xpb_out[68][186],u_xpb_out[69][186],u_xpb_out[70][186],u_xpb_out[71][186],u_xpb_out[72][186],u_xpb_out[73][186],u_xpb_out[74][186],u_xpb_out[75][186],u_xpb_out[76][186],u_xpb_out[77][186],u_xpb_out[78][186],u_xpb_out[79][186],u_xpb_out[80][186],u_xpb_out[81][186],u_xpb_out[82][186],u_xpb_out[83][186],u_xpb_out[84][186],u_xpb_out[85][186],u_xpb_out[86][186],u_xpb_out[87][186],u_xpb_out[88][186],u_xpb_out[89][186],u_xpb_out[90][186],u_xpb_out[91][186],u_xpb_out[92][186],u_xpb_out[93][186],u_xpb_out[94][186],u_xpb_out[95][186],u_xpb_out[96][186],u_xpb_out[97][186],u_xpb_out[98][186],u_xpb_out[99][186],u_xpb_out[100][186],u_xpb_out[101][186],u_xpb_out[102][186],u_xpb_out[103][186],u_xpb_out[104][186],u_xpb_out[105][186]};

assign col_out_187 = {u_xpb_out[0][187],u_xpb_out[1][187],u_xpb_out[2][187],u_xpb_out[3][187],u_xpb_out[4][187],u_xpb_out[5][187],u_xpb_out[6][187],u_xpb_out[7][187],u_xpb_out[8][187],u_xpb_out[9][187],u_xpb_out[10][187],u_xpb_out[11][187],u_xpb_out[12][187],u_xpb_out[13][187],u_xpb_out[14][187],u_xpb_out[15][187],u_xpb_out[16][187],u_xpb_out[17][187],u_xpb_out[18][187],u_xpb_out[19][187],u_xpb_out[20][187],u_xpb_out[21][187],u_xpb_out[22][187],u_xpb_out[23][187],u_xpb_out[24][187],u_xpb_out[25][187],u_xpb_out[26][187],u_xpb_out[27][187],u_xpb_out[28][187],u_xpb_out[29][187],u_xpb_out[30][187],u_xpb_out[31][187],u_xpb_out[32][187],u_xpb_out[33][187],u_xpb_out[34][187],u_xpb_out[35][187],u_xpb_out[36][187],u_xpb_out[37][187],u_xpb_out[38][187],u_xpb_out[39][187],u_xpb_out[40][187],u_xpb_out[41][187],u_xpb_out[42][187],u_xpb_out[43][187],u_xpb_out[44][187],u_xpb_out[45][187],u_xpb_out[46][187],u_xpb_out[47][187],u_xpb_out[48][187],u_xpb_out[49][187],u_xpb_out[50][187],u_xpb_out[51][187],u_xpb_out[52][187],u_xpb_out[53][187],u_xpb_out[54][187],u_xpb_out[55][187],u_xpb_out[56][187],u_xpb_out[57][187],u_xpb_out[58][187],u_xpb_out[59][187],u_xpb_out[60][187],u_xpb_out[61][187],u_xpb_out[62][187],u_xpb_out[63][187],u_xpb_out[64][187],u_xpb_out[65][187],u_xpb_out[66][187],u_xpb_out[67][187],u_xpb_out[68][187],u_xpb_out[69][187],u_xpb_out[70][187],u_xpb_out[71][187],u_xpb_out[72][187],u_xpb_out[73][187],u_xpb_out[74][187],u_xpb_out[75][187],u_xpb_out[76][187],u_xpb_out[77][187],u_xpb_out[78][187],u_xpb_out[79][187],u_xpb_out[80][187],u_xpb_out[81][187],u_xpb_out[82][187],u_xpb_out[83][187],u_xpb_out[84][187],u_xpb_out[85][187],u_xpb_out[86][187],u_xpb_out[87][187],u_xpb_out[88][187],u_xpb_out[89][187],u_xpb_out[90][187],u_xpb_out[91][187],u_xpb_out[92][187],u_xpb_out[93][187],u_xpb_out[94][187],u_xpb_out[95][187],u_xpb_out[96][187],u_xpb_out[97][187],u_xpb_out[98][187],u_xpb_out[99][187],u_xpb_out[100][187],u_xpb_out[101][187],u_xpb_out[102][187],u_xpb_out[103][187],u_xpb_out[104][187],u_xpb_out[105][187]};

assign col_out_188 = {u_xpb_out[0][188],u_xpb_out[1][188],u_xpb_out[2][188],u_xpb_out[3][188],u_xpb_out[4][188],u_xpb_out[5][188],u_xpb_out[6][188],u_xpb_out[7][188],u_xpb_out[8][188],u_xpb_out[9][188],u_xpb_out[10][188],u_xpb_out[11][188],u_xpb_out[12][188],u_xpb_out[13][188],u_xpb_out[14][188],u_xpb_out[15][188],u_xpb_out[16][188],u_xpb_out[17][188],u_xpb_out[18][188],u_xpb_out[19][188],u_xpb_out[20][188],u_xpb_out[21][188],u_xpb_out[22][188],u_xpb_out[23][188],u_xpb_out[24][188],u_xpb_out[25][188],u_xpb_out[26][188],u_xpb_out[27][188],u_xpb_out[28][188],u_xpb_out[29][188],u_xpb_out[30][188],u_xpb_out[31][188],u_xpb_out[32][188],u_xpb_out[33][188],u_xpb_out[34][188],u_xpb_out[35][188],u_xpb_out[36][188],u_xpb_out[37][188],u_xpb_out[38][188],u_xpb_out[39][188],u_xpb_out[40][188],u_xpb_out[41][188],u_xpb_out[42][188],u_xpb_out[43][188],u_xpb_out[44][188],u_xpb_out[45][188],u_xpb_out[46][188],u_xpb_out[47][188],u_xpb_out[48][188],u_xpb_out[49][188],u_xpb_out[50][188],u_xpb_out[51][188],u_xpb_out[52][188],u_xpb_out[53][188],u_xpb_out[54][188],u_xpb_out[55][188],u_xpb_out[56][188],u_xpb_out[57][188],u_xpb_out[58][188],u_xpb_out[59][188],u_xpb_out[60][188],u_xpb_out[61][188],u_xpb_out[62][188],u_xpb_out[63][188],u_xpb_out[64][188],u_xpb_out[65][188],u_xpb_out[66][188],u_xpb_out[67][188],u_xpb_out[68][188],u_xpb_out[69][188],u_xpb_out[70][188],u_xpb_out[71][188],u_xpb_out[72][188],u_xpb_out[73][188],u_xpb_out[74][188],u_xpb_out[75][188],u_xpb_out[76][188],u_xpb_out[77][188],u_xpb_out[78][188],u_xpb_out[79][188],u_xpb_out[80][188],u_xpb_out[81][188],u_xpb_out[82][188],u_xpb_out[83][188],u_xpb_out[84][188],u_xpb_out[85][188],u_xpb_out[86][188],u_xpb_out[87][188],u_xpb_out[88][188],u_xpb_out[89][188],u_xpb_out[90][188],u_xpb_out[91][188],u_xpb_out[92][188],u_xpb_out[93][188],u_xpb_out[94][188],u_xpb_out[95][188],u_xpb_out[96][188],u_xpb_out[97][188],u_xpb_out[98][188],u_xpb_out[99][188],u_xpb_out[100][188],u_xpb_out[101][188],u_xpb_out[102][188],u_xpb_out[103][188],u_xpb_out[104][188],u_xpb_out[105][188]};

assign col_out_189 = {u_xpb_out[0][189],u_xpb_out[1][189],u_xpb_out[2][189],u_xpb_out[3][189],u_xpb_out[4][189],u_xpb_out[5][189],u_xpb_out[6][189],u_xpb_out[7][189],u_xpb_out[8][189],u_xpb_out[9][189],u_xpb_out[10][189],u_xpb_out[11][189],u_xpb_out[12][189],u_xpb_out[13][189],u_xpb_out[14][189],u_xpb_out[15][189],u_xpb_out[16][189],u_xpb_out[17][189],u_xpb_out[18][189],u_xpb_out[19][189],u_xpb_out[20][189],u_xpb_out[21][189],u_xpb_out[22][189],u_xpb_out[23][189],u_xpb_out[24][189],u_xpb_out[25][189],u_xpb_out[26][189],u_xpb_out[27][189],u_xpb_out[28][189],u_xpb_out[29][189],u_xpb_out[30][189],u_xpb_out[31][189],u_xpb_out[32][189],u_xpb_out[33][189],u_xpb_out[34][189],u_xpb_out[35][189],u_xpb_out[36][189],u_xpb_out[37][189],u_xpb_out[38][189],u_xpb_out[39][189],u_xpb_out[40][189],u_xpb_out[41][189],u_xpb_out[42][189],u_xpb_out[43][189],u_xpb_out[44][189],u_xpb_out[45][189],u_xpb_out[46][189],u_xpb_out[47][189],u_xpb_out[48][189],u_xpb_out[49][189],u_xpb_out[50][189],u_xpb_out[51][189],u_xpb_out[52][189],u_xpb_out[53][189],u_xpb_out[54][189],u_xpb_out[55][189],u_xpb_out[56][189],u_xpb_out[57][189],u_xpb_out[58][189],u_xpb_out[59][189],u_xpb_out[60][189],u_xpb_out[61][189],u_xpb_out[62][189],u_xpb_out[63][189],u_xpb_out[64][189],u_xpb_out[65][189],u_xpb_out[66][189],u_xpb_out[67][189],u_xpb_out[68][189],u_xpb_out[69][189],u_xpb_out[70][189],u_xpb_out[71][189],u_xpb_out[72][189],u_xpb_out[73][189],u_xpb_out[74][189],u_xpb_out[75][189],u_xpb_out[76][189],u_xpb_out[77][189],u_xpb_out[78][189],u_xpb_out[79][189],u_xpb_out[80][189],u_xpb_out[81][189],u_xpb_out[82][189],u_xpb_out[83][189],u_xpb_out[84][189],u_xpb_out[85][189],u_xpb_out[86][189],u_xpb_out[87][189],u_xpb_out[88][189],u_xpb_out[89][189],u_xpb_out[90][189],u_xpb_out[91][189],u_xpb_out[92][189],u_xpb_out[93][189],u_xpb_out[94][189],u_xpb_out[95][189],u_xpb_out[96][189],u_xpb_out[97][189],u_xpb_out[98][189],u_xpb_out[99][189],u_xpb_out[100][189],u_xpb_out[101][189],u_xpb_out[102][189],u_xpb_out[103][189],u_xpb_out[104][189],u_xpb_out[105][189]};

assign col_out_190 = {u_xpb_out[0][190],u_xpb_out[1][190],u_xpb_out[2][190],u_xpb_out[3][190],u_xpb_out[4][190],u_xpb_out[5][190],u_xpb_out[6][190],u_xpb_out[7][190],u_xpb_out[8][190],u_xpb_out[9][190],u_xpb_out[10][190],u_xpb_out[11][190],u_xpb_out[12][190],u_xpb_out[13][190],u_xpb_out[14][190],u_xpb_out[15][190],u_xpb_out[16][190],u_xpb_out[17][190],u_xpb_out[18][190],u_xpb_out[19][190],u_xpb_out[20][190],u_xpb_out[21][190],u_xpb_out[22][190],u_xpb_out[23][190],u_xpb_out[24][190],u_xpb_out[25][190],u_xpb_out[26][190],u_xpb_out[27][190],u_xpb_out[28][190],u_xpb_out[29][190],u_xpb_out[30][190],u_xpb_out[31][190],u_xpb_out[32][190],u_xpb_out[33][190],u_xpb_out[34][190],u_xpb_out[35][190],u_xpb_out[36][190],u_xpb_out[37][190],u_xpb_out[38][190],u_xpb_out[39][190],u_xpb_out[40][190],u_xpb_out[41][190],u_xpb_out[42][190],u_xpb_out[43][190],u_xpb_out[44][190],u_xpb_out[45][190],u_xpb_out[46][190],u_xpb_out[47][190],u_xpb_out[48][190],u_xpb_out[49][190],u_xpb_out[50][190],u_xpb_out[51][190],u_xpb_out[52][190],u_xpb_out[53][190],u_xpb_out[54][190],u_xpb_out[55][190],u_xpb_out[56][190],u_xpb_out[57][190],u_xpb_out[58][190],u_xpb_out[59][190],u_xpb_out[60][190],u_xpb_out[61][190],u_xpb_out[62][190],u_xpb_out[63][190],u_xpb_out[64][190],u_xpb_out[65][190],u_xpb_out[66][190],u_xpb_out[67][190],u_xpb_out[68][190],u_xpb_out[69][190],u_xpb_out[70][190],u_xpb_out[71][190],u_xpb_out[72][190],u_xpb_out[73][190],u_xpb_out[74][190],u_xpb_out[75][190],u_xpb_out[76][190],u_xpb_out[77][190],u_xpb_out[78][190],u_xpb_out[79][190],u_xpb_out[80][190],u_xpb_out[81][190],u_xpb_out[82][190],u_xpb_out[83][190],u_xpb_out[84][190],u_xpb_out[85][190],u_xpb_out[86][190],u_xpb_out[87][190],u_xpb_out[88][190],u_xpb_out[89][190],u_xpb_out[90][190],u_xpb_out[91][190],u_xpb_out[92][190],u_xpb_out[93][190],u_xpb_out[94][190],u_xpb_out[95][190],u_xpb_out[96][190],u_xpb_out[97][190],u_xpb_out[98][190],u_xpb_out[99][190],u_xpb_out[100][190],u_xpb_out[101][190],u_xpb_out[102][190],u_xpb_out[103][190],u_xpb_out[104][190],u_xpb_out[105][190]};

assign col_out_191 = {u_xpb_out[0][191],u_xpb_out[1][191],u_xpb_out[2][191],u_xpb_out[3][191],u_xpb_out[4][191],u_xpb_out[5][191],u_xpb_out[6][191],u_xpb_out[7][191],u_xpb_out[8][191],u_xpb_out[9][191],u_xpb_out[10][191],u_xpb_out[11][191],u_xpb_out[12][191],u_xpb_out[13][191],u_xpb_out[14][191],u_xpb_out[15][191],u_xpb_out[16][191],u_xpb_out[17][191],u_xpb_out[18][191],u_xpb_out[19][191],u_xpb_out[20][191],u_xpb_out[21][191],u_xpb_out[22][191],u_xpb_out[23][191],u_xpb_out[24][191],u_xpb_out[25][191],u_xpb_out[26][191],u_xpb_out[27][191],u_xpb_out[28][191],u_xpb_out[29][191],u_xpb_out[30][191],u_xpb_out[31][191],u_xpb_out[32][191],u_xpb_out[33][191],u_xpb_out[34][191],u_xpb_out[35][191],u_xpb_out[36][191],u_xpb_out[37][191],u_xpb_out[38][191],u_xpb_out[39][191],u_xpb_out[40][191],u_xpb_out[41][191],u_xpb_out[42][191],u_xpb_out[43][191],u_xpb_out[44][191],u_xpb_out[45][191],u_xpb_out[46][191],u_xpb_out[47][191],u_xpb_out[48][191],u_xpb_out[49][191],u_xpb_out[50][191],u_xpb_out[51][191],u_xpb_out[52][191],u_xpb_out[53][191],u_xpb_out[54][191],u_xpb_out[55][191],u_xpb_out[56][191],u_xpb_out[57][191],u_xpb_out[58][191],u_xpb_out[59][191],u_xpb_out[60][191],u_xpb_out[61][191],u_xpb_out[62][191],u_xpb_out[63][191],u_xpb_out[64][191],u_xpb_out[65][191],u_xpb_out[66][191],u_xpb_out[67][191],u_xpb_out[68][191],u_xpb_out[69][191],u_xpb_out[70][191],u_xpb_out[71][191],u_xpb_out[72][191],u_xpb_out[73][191],u_xpb_out[74][191],u_xpb_out[75][191],u_xpb_out[76][191],u_xpb_out[77][191],u_xpb_out[78][191],u_xpb_out[79][191],u_xpb_out[80][191],u_xpb_out[81][191],u_xpb_out[82][191],u_xpb_out[83][191],u_xpb_out[84][191],u_xpb_out[85][191],u_xpb_out[86][191],u_xpb_out[87][191],u_xpb_out[88][191],u_xpb_out[89][191],u_xpb_out[90][191],u_xpb_out[91][191],u_xpb_out[92][191],u_xpb_out[93][191],u_xpb_out[94][191],u_xpb_out[95][191],u_xpb_out[96][191],u_xpb_out[97][191],u_xpb_out[98][191],u_xpb_out[99][191],u_xpb_out[100][191],u_xpb_out[101][191],u_xpb_out[102][191],u_xpb_out[103][191],u_xpb_out[104][191],u_xpb_out[105][191]};

assign col_out_192 = {u_xpb_out[0][192],u_xpb_out[1][192],u_xpb_out[2][192],u_xpb_out[3][192],u_xpb_out[4][192],u_xpb_out[5][192],u_xpb_out[6][192],u_xpb_out[7][192],u_xpb_out[8][192],u_xpb_out[9][192],u_xpb_out[10][192],u_xpb_out[11][192],u_xpb_out[12][192],u_xpb_out[13][192],u_xpb_out[14][192],u_xpb_out[15][192],u_xpb_out[16][192],u_xpb_out[17][192],u_xpb_out[18][192],u_xpb_out[19][192],u_xpb_out[20][192],u_xpb_out[21][192],u_xpb_out[22][192],u_xpb_out[23][192],u_xpb_out[24][192],u_xpb_out[25][192],u_xpb_out[26][192],u_xpb_out[27][192],u_xpb_out[28][192],u_xpb_out[29][192],u_xpb_out[30][192],u_xpb_out[31][192],u_xpb_out[32][192],u_xpb_out[33][192],u_xpb_out[34][192],u_xpb_out[35][192],u_xpb_out[36][192],u_xpb_out[37][192],u_xpb_out[38][192],u_xpb_out[39][192],u_xpb_out[40][192],u_xpb_out[41][192],u_xpb_out[42][192],u_xpb_out[43][192],u_xpb_out[44][192],u_xpb_out[45][192],u_xpb_out[46][192],u_xpb_out[47][192],u_xpb_out[48][192],u_xpb_out[49][192],u_xpb_out[50][192],u_xpb_out[51][192],u_xpb_out[52][192],u_xpb_out[53][192],u_xpb_out[54][192],u_xpb_out[55][192],u_xpb_out[56][192],u_xpb_out[57][192],u_xpb_out[58][192],u_xpb_out[59][192],u_xpb_out[60][192],u_xpb_out[61][192],u_xpb_out[62][192],u_xpb_out[63][192],u_xpb_out[64][192],u_xpb_out[65][192],u_xpb_out[66][192],u_xpb_out[67][192],u_xpb_out[68][192],u_xpb_out[69][192],u_xpb_out[70][192],u_xpb_out[71][192],u_xpb_out[72][192],u_xpb_out[73][192],u_xpb_out[74][192],u_xpb_out[75][192],u_xpb_out[76][192],u_xpb_out[77][192],u_xpb_out[78][192],u_xpb_out[79][192],u_xpb_out[80][192],u_xpb_out[81][192],u_xpb_out[82][192],u_xpb_out[83][192],u_xpb_out[84][192],u_xpb_out[85][192],u_xpb_out[86][192],u_xpb_out[87][192],u_xpb_out[88][192],u_xpb_out[89][192],u_xpb_out[90][192],u_xpb_out[91][192],u_xpb_out[92][192],u_xpb_out[93][192],u_xpb_out[94][192],u_xpb_out[95][192],u_xpb_out[96][192],u_xpb_out[97][192],u_xpb_out[98][192],u_xpb_out[99][192],u_xpb_out[100][192],u_xpb_out[101][192],u_xpb_out[102][192],u_xpb_out[103][192],u_xpb_out[104][192],u_xpb_out[105][192]};

assign col_out_193 = {u_xpb_out[0][193],u_xpb_out[1][193],u_xpb_out[2][193],u_xpb_out[3][193],u_xpb_out[4][193],u_xpb_out[5][193],u_xpb_out[6][193],u_xpb_out[7][193],u_xpb_out[8][193],u_xpb_out[9][193],u_xpb_out[10][193],u_xpb_out[11][193],u_xpb_out[12][193],u_xpb_out[13][193],u_xpb_out[14][193],u_xpb_out[15][193],u_xpb_out[16][193],u_xpb_out[17][193],u_xpb_out[18][193],u_xpb_out[19][193],u_xpb_out[20][193],u_xpb_out[21][193],u_xpb_out[22][193],u_xpb_out[23][193],u_xpb_out[24][193],u_xpb_out[25][193],u_xpb_out[26][193],u_xpb_out[27][193],u_xpb_out[28][193],u_xpb_out[29][193],u_xpb_out[30][193],u_xpb_out[31][193],u_xpb_out[32][193],u_xpb_out[33][193],u_xpb_out[34][193],u_xpb_out[35][193],u_xpb_out[36][193],u_xpb_out[37][193],u_xpb_out[38][193],u_xpb_out[39][193],u_xpb_out[40][193],u_xpb_out[41][193],u_xpb_out[42][193],u_xpb_out[43][193],u_xpb_out[44][193],u_xpb_out[45][193],u_xpb_out[46][193],u_xpb_out[47][193],u_xpb_out[48][193],u_xpb_out[49][193],u_xpb_out[50][193],u_xpb_out[51][193],u_xpb_out[52][193],u_xpb_out[53][193],u_xpb_out[54][193],u_xpb_out[55][193],u_xpb_out[56][193],u_xpb_out[57][193],u_xpb_out[58][193],u_xpb_out[59][193],u_xpb_out[60][193],u_xpb_out[61][193],u_xpb_out[62][193],u_xpb_out[63][193],u_xpb_out[64][193],u_xpb_out[65][193],u_xpb_out[66][193],u_xpb_out[67][193],u_xpb_out[68][193],u_xpb_out[69][193],u_xpb_out[70][193],u_xpb_out[71][193],u_xpb_out[72][193],u_xpb_out[73][193],u_xpb_out[74][193],u_xpb_out[75][193],u_xpb_out[76][193],u_xpb_out[77][193],u_xpb_out[78][193],u_xpb_out[79][193],u_xpb_out[80][193],u_xpb_out[81][193],u_xpb_out[82][193],u_xpb_out[83][193],u_xpb_out[84][193],u_xpb_out[85][193],u_xpb_out[86][193],u_xpb_out[87][193],u_xpb_out[88][193],u_xpb_out[89][193],u_xpb_out[90][193],u_xpb_out[91][193],u_xpb_out[92][193],u_xpb_out[93][193],u_xpb_out[94][193],u_xpb_out[95][193],u_xpb_out[96][193],u_xpb_out[97][193],u_xpb_out[98][193],u_xpb_out[99][193],u_xpb_out[100][193],u_xpb_out[101][193],u_xpb_out[102][193],u_xpb_out[103][193],u_xpb_out[104][193],u_xpb_out[105][193]};

assign col_out_194 = {u_xpb_out[0][194],u_xpb_out[1][194],u_xpb_out[2][194],u_xpb_out[3][194],u_xpb_out[4][194],u_xpb_out[5][194],u_xpb_out[6][194],u_xpb_out[7][194],u_xpb_out[8][194],u_xpb_out[9][194],u_xpb_out[10][194],u_xpb_out[11][194],u_xpb_out[12][194],u_xpb_out[13][194],u_xpb_out[14][194],u_xpb_out[15][194],u_xpb_out[16][194],u_xpb_out[17][194],u_xpb_out[18][194],u_xpb_out[19][194],u_xpb_out[20][194],u_xpb_out[21][194],u_xpb_out[22][194],u_xpb_out[23][194],u_xpb_out[24][194],u_xpb_out[25][194],u_xpb_out[26][194],u_xpb_out[27][194],u_xpb_out[28][194],u_xpb_out[29][194],u_xpb_out[30][194],u_xpb_out[31][194],u_xpb_out[32][194],u_xpb_out[33][194],u_xpb_out[34][194],u_xpb_out[35][194],u_xpb_out[36][194],u_xpb_out[37][194],u_xpb_out[38][194],u_xpb_out[39][194],u_xpb_out[40][194],u_xpb_out[41][194],u_xpb_out[42][194],u_xpb_out[43][194],u_xpb_out[44][194],u_xpb_out[45][194],u_xpb_out[46][194],u_xpb_out[47][194],u_xpb_out[48][194],u_xpb_out[49][194],u_xpb_out[50][194],u_xpb_out[51][194],u_xpb_out[52][194],u_xpb_out[53][194],u_xpb_out[54][194],u_xpb_out[55][194],u_xpb_out[56][194],u_xpb_out[57][194],u_xpb_out[58][194],u_xpb_out[59][194],u_xpb_out[60][194],u_xpb_out[61][194],u_xpb_out[62][194],u_xpb_out[63][194],u_xpb_out[64][194],u_xpb_out[65][194],u_xpb_out[66][194],u_xpb_out[67][194],u_xpb_out[68][194],u_xpb_out[69][194],u_xpb_out[70][194],u_xpb_out[71][194],u_xpb_out[72][194],u_xpb_out[73][194],u_xpb_out[74][194],u_xpb_out[75][194],u_xpb_out[76][194],u_xpb_out[77][194],u_xpb_out[78][194],u_xpb_out[79][194],u_xpb_out[80][194],u_xpb_out[81][194],u_xpb_out[82][194],u_xpb_out[83][194],u_xpb_out[84][194],u_xpb_out[85][194],u_xpb_out[86][194],u_xpb_out[87][194],u_xpb_out[88][194],u_xpb_out[89][194],u_xpb_out[90][194],u_xpb_out[91][194],u_xpb_out[92][194],u_xpb_out[93][194],u_xpb_out[94][194],u_xpb_out[95][194],u_xpb_out[96][194],u_xpb_out[97][194],u_xpb_out[98][194],u_xpb_out[99][194],u_xpb_out[100][194],u_xpb_out[101][194],u_xpb_out[102][194],u_xpb_out[103][194],u_xpb_out[104][194],u_xpb_out[105][194]};

assign col_out_195 = {u_xpb_out[0][195],u_xpb_out[1][195],u_xpb_out[2][195],u_xpb_out[3][195],u_xpb_out[4][195],u_xpb_out[5][195],u_xpb_out[6][195],u_xpb_out[7][195],u_xpb_out[8][195],u_xpb_out[9][195],u_xpb_out[10][195],u_xpb_out[11][195],u_xpb_out[12][195],u_xpb_out[13][195],u_xpb_out[14][195],u_xpb_out[15][195],u_xpb_out[16][195],u_xpb_out[17][195],u_xpb_out[18][195],u_xpb_out[19][195],u_xpb_out[20][195],u_xpb_out[21][195],u_xpb_out[22][195],u_xpb_out[23][195],u_xpb_out[24][195],u_xpb_out[25][195],u_xpb_out[26][195],u_xpb_out[27][195],u_xpb_out[28][195],u_xpb_out[29][195],u_xpb_out[30][195],u_xpb_out[31][195],u_xpb_out[32][195],u_xpb_out[33][195],u_xpb_out[34][195],u_xpb_out[35][195],u_xpb_out[36][195],u_xpb_out[37][195],u_xpb_out[38][195],u_xpb_out[39][195],u_xpb_out[40][195],u_xpb_out[41][195],u_xpb_out[42][195],u_xpb_out[43][195],u_xpb_out[44][195],u_xpb_out[45][195],u_xpb_out[46][195],u_xpb_out[47][195],u_xpb_out[48][195],u_xpb_out[49][195],u_xpb_out[50][195],u_xpb_out[51][195],u_xpb_out[52][195],u_xpb_out[53][195],u_xpb_out[54][195],u_xpb_out[55][195],u_xpb_out[56][195],u_xpb_out[57][195],u_xpb_out[58][195],u_xpb_out[59][195],u_xpb_out[60][195],u_xpb_out[61][195],u_xpb_out[62][195],u_xpb_out[63][195],u_xpb_out[64][195],u_xpb_out[65][195],u_xpb_out[66][195],u_xpb_out[67][195],u_xpb_out[68][195],u_xpb_out[69][195],u_xpb_out[70][195],u_xpb_out[71][195],u_xpb_out[72][195],u_xpb_out[73][195],u_xpb_out[74][195],u_xpb_out[75][195],u_xpb_out[76][195],u_xpb_out[77][195],u_xpb_out[78][195],u_xpb_out[79][195],u_xpb_out[80][195],u_xpb_out[81][195],u_xpb_out[82][195],u_xpb_out[83][195],u_xpb_out[84][195],u_xpb_out[85][195],u_xpb_out[86][195],u_xpb_out[87][195],u_xpb_out[88][195],u_xpb_out[89][195],u_xpb_out[90][195],u_xpb_out[91][195],u_xpb_out[92][195],u_xpb_out[93][195],u_xpb_out[94][195],u_xpb_out[95][195],u_xpb_out[96][195],u_xpb_out[97][195],u_xpb_out[98][195],u_xpb_out[99][195],u_xpb_out[100][195],u_xpb_out[101][195],u_xpb_out[102][195],u_xpb_out[103][195],u_xpb_out[104][195],u_xpb_out[105][195]};

assign col_out_196 = {u_xpb_out[0][196],u_xpb_out[1][196],u_xpb_out[2][196],u_xpb_out[3][196],u_xpb_out[4][196],u_xpb_out[5][196],u_xpb_out[6][196],u_xpb_out[7][196],u_xpb_out[8][196],u_xpb_out[9][196],u_xpb_out[10][196],u_xpb_out[11][196],u_xpb_out[12][196],u_xpb_out[13][196],u_xpb_out[14][196],u_xpb_out[15][196],u_xpb_out[16][196],u_xpb_out[17][196],u_xpb_out[18][196],u_xpb_out[19][196],u_xpb_out[20][196],u_xpb_out[21][196],u_xpb_out[22][196],u_xpb_out[23][196],u_xpb_out[24][196],u_xpb_out[25][196],u_xpb_out[26][196],u_xpb_out[27][196],u_xpb_out[28][196],u_xpb_out[29][196],u_xpb_out[30][196],u_xpb_out[31][196],u_xpb_out[32][196],u_xpb_out[33][196],u_xpb_out[34][196],u_xpb_out[35][196],u_xpb_out[36][196],u_xpb_out[37][196],u_xpb_out[38][196],u_xpb_out[39][196],u_xpb_out[40][196],u_xpb_out[41][196],u_xpb_out[42][196],u_xpb_out[43][196],u_xpb_out[44][196],u_xpb_out[45][196],u_xpb_out[46][196],u_xpb_out[47][196],u_xpb_out[48][196],u_xpb_out[49][196],u_xpb_out[50][196],u_xpb_out[51][196],u_xpb_out[52][196],u_xpb_out[53][196],u_xpb_out[54][196],u_xpb_out[55][196],u_xpb_out[56][196],u_xpb_out[57][196],u_xpb_out[58][196],u_xpb_out[59][196],u_xpb_out[60][196],u_xpb_out[61][196],u_xpb_out[62][196],u_xpb_out[63][196],u_xpb_out[64][196],u_xpb_out[65][196],u_xpb_out[66][196],u_xpb_out[67][196],u_xpb_out[68][196],u_xpb_out[69][196],u_xpb_out[70][196],u_xpb_out[71][196],u_xpb_out[72][196],u_xpb_out[73][196],u_xpb_out[74][196],u_xpb_out[75][196],u_xpb_out[76][196],u_xpb_out[77][196],u_xpb_out[78][196],u_xpb_out[79][196],u_xpb_out[80][196],u_xpb_out[81][196],u_xpb_out[82][196],u_xpb_out[83][196],u_xpb_out[84][196],u_xpb_out[85][196],u_xpb_out[86][196],u_xpb_out[87][196],u_xpb_out[88][196],u_xpb_out[89][196],u_xpb_out[90][196],u_xpb_out[91][196],u_xpb_out[92][196],u_xpb_out[93][196],u_xpb_out[94][196],u_xpb_out[95][196],u_xpb_out[96][196],u_xpb_out[97][196],u_xpb_out[98][196],u_xpb_out[99][196],u_xpb_out[100][196],u_xpb_out[101][196],u_xpb_out[102][196],u_xpb_out[103][196],u_xpb_out[104][196],u_xpb_out[105][196]};

assign col_out_197 = {u_xpb_out[0][197],u_xpb_out[1][197],u_xpb_out[2][197],u_xpb_out[3][197],u_xpb_out[4][197],u_xpb_out[5][197],u_xpb_out[6][197],u_xpb_out[7][197],u_xpb_out[8][197],u_xpb_out[9][197],u_xpb_out[10][197],u_xpb_out[11][197],u_xpb_out[12][197],u_xpb_out[13][197],u_xpb_out[14][197],u_xpb_out[15][197],u_xpb_out[16][197],u_xpb_out[17][197],u_xpb_out[18][197],u_xpb_out[19][197],u_xpb_out[20][197],u_xpb_out[21][197],u_xpb_out[22][197],u_xpb_out[23][197],u_xpb_out[24][197],u_xpb_out[25][197],u_xpb_out[26][197],u_xpb_out[27][197],u_xpb_out[28][197],u_xpb_out[29][197],u_xpb_out[30][197],u_xpb_out[31][197],u_xpb_out[32][197],u_xpb_out[33][197],u_xpb_out[34][197],u_xpb_out[35][197],u_xpb_out[36][197],u_xpb_out[37][197],u_xpb_out[38][197],u_xpb_out[39][197],u_xpb_out[40][197],u_xpb_out[41][197],u_xpb_out[42][197],u_xpb_out[43][197],u_xpb_out[44][197],u_xpb_out[45][197],u_xpb_out[46][197],u_xpb_out[47][197],u_xpb_out[48][197],u_xpb_out[49][197],u_xpb_out[50][197],u_xpb_out[51][197],u_xpb_out[52][197],u_xpb_out[53][197],u_xpb_out[54][197],u_xpb_out[55][197],u_xpb_out[56][197],u_xpb_out[57][197],u_xpb_out[58][197],u_xpb_out[59][197],u_xpb_out[60][197],u_xpb_out[61][197],u_xpb_out[62][197],u_xpb_out[63][197],u_xpb_out[64][197],u_xpb_out[65][197],u_xpb_out[66][197],u_xpb_out[67][197],u_xpb_out[68][197],u_xpb_out[69][197],u_xpb_out[70][197],u_xpb_out[71][197],u_xpb_out[72][197],u_xpb_out[73][197],u_xpb_out[74][197],u_xpb_out[75][197],u_xpb_out[76][197],u_xpb_out[77][197],u_xpb_out[78][197],u_xpb_out[79][197],u_xpb_out[80][197],u_xpb_out[81][197],u_xpb_out[82][197],u_xpb_out[83][197],u_xpb_out[84][197],u_xpb_out[85][197],u_xpb_out[86][197],u_xpb_out[87][197],u_xpb_out[88][197],u_xpb_out[89][197],u_xpb_out[90][197],u_xpb_out[91][197],u_xpb_out[92][197],u_xpb_out[93][197],u_xpb_out[94][197],u_xpb_out[95][197],u_xpb_out[96][197],u_xpb_out[97][197],u_xpb_out[98][197],u_xpb_out[99][197],u_xpb_out[100][197],u_xpb_out[101][197],u_xpb_out[102][197],u_xpb_out[103][197],u_xpb_out[104][197],u_xpb_out[105][197]};

assign col_out_198 = {u_xpb_out[0][198],u_xpb_out[1][198],u_xpb_out[2][198],u_xpb_out[3][198],u_xpb_out[4][198],u_xpb_out[5][198],u_xpb_out[6][198],u_xpb_out[7][198],u_xpb_out[8][198],u_xpb_out[9][198],u_xpb_out[10][198],u_xpb_out[11][198],u_xpb_out[12][198],u_xpb_out[13][198],u_xpb_out[14][198],u_xpb_out[15][198],u_xpb_out[16][198],u_xpb_out[17][198],u_xpb_out[18][198],u_xpb_out[19][198],u_xpb_out[20][198],u_xpb_out[21][198],u_xpb_out[22][198],u_xpb_out[23][198],u_xpb_out[24][198],u_xpb_out[25][198],u_xpb_out[26][198],u_xpb_out[27][198],u_xpb_out[28][198],u_xpb_out[29][198],u_xpb_out[30][198],u_xpb_out[31][198],u_xpb_out[32][198],u_xpb_out[33][198],u_xpb_out[34][198],u_xpb_out[35][198],u_xpb_out[36][198],u_xpb_out[37][198],u_xpb_out[38][198],u_xpb_out[39][198],u_xpb_out[40][198],u_xpb_out[41][198],u_xpb_out[42][198],u_xpb_out[43][198],u_xpb_out[44][198],u_xpb_out[45][198],u_xpb_out[46][198],u_xpb_out[47][198],u_xpb_out[48][198],u_xpb_out[49][198],u_xpb_out[50][198],u_xpb_out[51][198],u_xpb_out[52][198],u_xpb_out[53][198],u_xpb_out[54][198],u_xpb_out[55][198],u_xpb_out[56][198],u_xpb_out[57][198],u_xpb_out[58][198],u_xpb_out[59][198],u_xpb_out[60][198],u_xpb_out[61][198],u_xpb_out[62][198],u_xpb_out[63][198],u_xpb_out[64][198],u_xpb_out[65][198],u_xpb_out[66][198],u_xpb_out[67][198],u_xpb_out[68][198],u_xpb_out[69][198],u_xpb_out[70][198],u_xpb_out[71][198],u_xpb_out[72][198],u_xpb_out[73][198],u_xpb_out[74][198],u_xpb_out[75][198],u_xpb_out[76][198],u_xpb_out[77][198],u_xpb_out[78][198],u_xpb_out[79][198],u_xpb_out[80][198],u_xpb_out[81][198],u_xpb_out[82][198],u_xpb_out[83][198],u_xpb_out[84][198],u_xpb_out[85][198],u_xpb_out[86][198],u_xpb_out[87][198],u_xpb_out[88][198],u_xpb_out[89][198],u_xpb_out[90][198],u_xpb_out[91][198],u_xpb_out[92][198],u_xpb_out[93][198],u_xpb_out[94][198],u_xpb_out[95][198],u_xpb_out[96][198],u_xpb_out[97][198],u_xpb_out[98][198],u_xpb_out[99][198],u_xpb_out[100][198],u_xpb_out[101][198],u_xpb_out[102][198],u_xpb_out[103][198],u_xpb_out[104][198],u_xpb_out[105][198]};

assign col_out_199 = {u_xpb_out[0][199],u_xpb_out[1][199],u_xpb_out[2][199],u_xpb_out[3][199],u_xpb_out[4][199],u_xpb_out[5][199],u_xpb_out[6][199],u_xpb_out[7][199],u_xpb_out[8][199],u_xpb_out[9][199],u_xpb_out[10][199],u_xpb_out[11][199],u_xpb_out[12][199],u_xpb_out[13][199],u_xpb_out[14][199],u_xpb_out[15][199],u_xpb_out[16][199],u_xpb_out[17][199],u_xpb_out[18][199],u_xpb_out[19][199],u_xpb_out[20][199],u_xpb_out[21][199],u_xpb_out[22][199],u_xpb_out[23][199],u_xpb_out[24][199],u_xpb_out[25][199],u_xpb_out[26][199],u_xpb_out[27][199],u_xpb_out[28][199],u_xpb_out[29][199],u_xpb_out[30][199],u_xpb_out[31][199],u_xpb_out[32][199],u_xpb_out[33][199],u_xpb_out[34][199],u_xpb_out[35][199],u_xpb_out[36][199],u_xpb_out[37][199],u_xpb_out[38][199],u_xpb_out[39][199],u_xpb_out[40][199],u_xpb_out[41][199],u_xpb_out[42][199],u_xpb_out[43][199],u_xpb_out[44][199],u_xpb_out[45][199],u_xpb_out[46][199],u_xpb_out[47][199],u_xpb_out[48][199],u_xpb_out[49][199],u_xpb_out[50][199],u_xpb_out[51][199],u_xpb_out[52][199],u_xpb_out[53][199],u_xpb_out[54][199],u_xpb_out[55][199],u_xpb_out[56][199],u_xpb_out[57][199],u_xpb_out[58][199],u_xpb_out[59][199],u_xpb_out[60][199],u_xpb_out[61][199],u_xpb_out[62][199],u_xpb_out[63][199],u_xpb_out[64][199],u_xpb_out[65][199],u_xpb_out[66][199],u_xpb_out[67][199],u_xpb_out[68][199],u_xpb_out[69][199],u_xpb_out[70][199],u_xpb_out[71][199],u_xpb_out[72][199],u_xpb_out[73][199],u_xpb_out[74][199],u_xpb_out[75][199],u_xpb_out[76][199],u_xpb_out[77][199],u_xpb_out[78][199],u_xpb_out[79][199],u_xpb_out[80][199],u_xpb_out[81][199],u_xpb_out[82][199],u_xpb_out[83][199],u_xpb_out[84][199],u_xpb_out[85][199],u_xpb_out[86][199],u_xpb_out[87][199],u_xpb_out[88][199],u_xpb_out[89][199],u_xpb_out[90][199],u_xpb_out[91][199],u_xpb_out[92][199],u_xpb_out[93][199],u_xpb_out[94][199],u_xpb_out[95][199],u_xpb_out[96][199],u_xpb_out[97][199],u_xpb_out[98][199],u_xpb_out[99][199],u_xpb_out[100][199],u_xpb_out[101][199],u_xpb_out[102][199],u_xpb_out[103][199],u_xpb_out[104][199],u_xpb_out[105][199]};

assign col_out_200 = {u_xpb_out[0][200],u_xpb_out[1][200],u_xpb_out[2][200],u_xpb_out[3][200],u_xpb_out[4][200],u_xpb_out[5][200],u_xpb_out[6][200],u_xpb_out[7][200],u_xpb_out[8][200],u_xpb_out[9][200],u_xpb_out[10][200],u_xpb_out[11][200],u_xpb_out[12][200],u_xpb_out[13][200],u_xpb_out[14][200],u_xpb_out[15][200],u_xpb_out[16][200],u_xpb_out[17][200],u_xpb_out[18][200],u_xpb_out[19][200],u_xpb_out[20][200],u_xpb_out[21][200],u_xpb_out[22][200],u_xpb_out[23][200],u_xpb_out[24][200],u_xpb_out[25][200],u_xpb_out[26][200],u_xpb_out[27][200],u_xpb_out[28][200],u_xpb_out[29][200],u_xpb_out[30][200],u_xpb_out[31][200],u_xpb_out[32][200],u_xpb_out[33][200],u_xpb_out[34][200],u_xpb_out[35][200],u_xpb_out[36][200],u_xpb_out[37][200],u_xpb_out[38][200],u_xpb_out[39][200],u_xpb_out[40][200],u_xpb_out[41][200],u_xpb_out[42][200],u_xpb_out[43][200],u_xpb_out[44][200],u_xpb_out[45][200],u_xpb_out[46][200],u_xpb_out[47][200],u_xpb_out[48][200],u_xpb_out[49][200],u_xpb_out[50][200],u_xpb_out[51][200],u_xpb_out[52][200],u_xpb_out[53][200],u_xpb_out[54][200],u_xpb_out[55][200],u_xpb_out[56][200],u_xpb_out[57][200],u_xpb_out[58][200],u_xpb_out[59][200],u_xpb_out[60][200],u_xpb_out[61][200],u_xpb_out[62][200],u_xpb_out[63][200],u_xpb_out[64][200],u_xpb_out[65][200],u_xpb_out[66][200],u_xpb_out[67][200],u_xpb_out[68][200],u_xpb_out[69][200],u_xpb_out[70][200],u_xpb_out[71][200],u_xpb_out[72][200],u_xpb_out[73][200],u_xpb_out[74][200],u_xpb_out[75][200],u_xpb_out[76][200],u_xpb_out[77][200],u_xpb_out[78][200],u_xpb_out[79][200],u_xpb_out[80][200],u_xpb_out[81][200],u_xpb_out[82][200],u_xpb_out[83][200],u_xpb_out[84][200],u_xpb_out[85][200],u_xpb_out[86][200],u_xpb_out[87][200],u_xpb_out[88][200],u_xpb_out[89][200],u_xpb_out[90][200],u_xpb_out[91][200],u_xpb_out[92][200],u_xpb_out[93][200],u_xpb_out[94][200],u_xpb_out[95][200],u_xpb_out[96][200],u_xpb_out[97][200],u_xpb_out[98][200],u_xpb_out[99][200],u_xpb_out[100][200],u_xpb_out[101][200],u_xpb_out[102][200],u_xpb_out[103][200],u_xpb_out[104][200],u_xpb_out[105][200]};

assign col_out_201 = {u_xpb_out[0][201],u_xpb_out[1][201],u_xpb_out[2][201],u_xpb_out[3][201],u_xpb_out[4][201],u_xpb_out[5][201],u_xpb_out[6][201],u_xpb_out[7][201],u_xpb_out[8][201],u_xpb_out[9][201],u_xpb_out[10][201],u_xpb_out[11][201],u_xpb_out[12][201],u_xpb_out[13][201],u_xpb_out[14][201],u_xpb_out[15][201],u_xpb_out[16][201],u_xpb_out[17][201],u_xpb_out[18][201],u_xpb_out[19][201],u_xpb_out[20][201],u_xpb_out[21][201],u_xpb_out[22][201],u_xpb_out[23][201],u_xpb_out[24][201],u_xpb_out[25][201],u_xpb_out[26][201],u_xpb_out[27][201],u_xpb_out[28][201],u_xpb_out[29][201],u_xpb_out[30][201],u_xpb_out[31][201],u_xpb_out[32][201],u_xpb_out[33][201],u_xpb_out[34][201],u_xpb_out[35][201],u_xpb_out[36][201],u_xpb_out[37][201],u_xpb_out[38][201],u_xpb_out[39][201],u_xpb_out[40][201],u_xpb_out[41][201],u_xpb_out[42][201],u_xpb_out[43][201],u_xpb_out[44][201],u_xpb_out[45][201],u_xpb_out[46][201],u_xpb_out[47][201],u_xpb_out[48][201],u_xpb_out[49][201],u_xpb_out[50][201],u_xpb_out[51][201],u_xpb_out[52][201],u_xpb_out[53][201],u_xpb_out[54][201],u_xpb_out[55][201],u_xpb_out[56][201],u_xpb_out[57][201],u_xpb_out[58][201],u_xpb_out[59][201],u_xpb_out[60][201],u_xpb_out[61][201],u_xpb_out[62][201],u_xpb_out[63][201],u_xpb_out[64][201],u_xpb_out[65][201],u_xpb_out[66][201],u_xpb_out[67][201],u_xpb_out[68][201],u_xpb_out[69][201],u_xpb_out[70][201],u_xpb_out[71][201],u_xpb_out[72][201],u_xpb_out[73][201],u_xpb_out[74][201],u_xpb_out[75][201],u_xpb_out[76][201],u_xpb_out[77][201],u_xpb_out[78][201],u_xpb_out[79][201],u_xpb_out[80][201],u_xpb_out[81][201],u_xpb_out[82][201],u_xpb_out[83][201],u_xpb_out[84][201],u_xpb_out[85][201],u_xpb_out[86][201],u_xpb_out[87][201],u_xpb_out[88][201],u_xpb_out[89][201],u_xpb_out[90][201],u_xpb_out[91][201],u_xpb_out[92][201],u_xpb_out[93][201],u_xpb_out[94][201],u_xpb_out[95][201],u_xpb_out[96][201],u_xpb_out[97][201],u_xpb_out[98][201],u_xpb_out[99][201],u_xpb_out[100][201],u_xpb_out[101][201],u_xpb_out[102][201],u_xpb_out[103][201],u_xpb_out[104][201],u_xpb_out[105][201]};

assign col_out_202 = {u_xpb_out[0][202],u_xpb_out[1][202],u_xpb_out[2][202],u_xpb_out[3][202],u_xpb_out[4][202],u_xpb_out[5][202],u_xpb_out[6][202],u_xpb_out[7][202],u_xpb_out[8][202],u_xpb_out[9][202],u_xpb_out[10][202],u_xpb_out[11][202],u_xpb_out[12][202],u_xpb_out[13][202],u_xpb_out[14][202],u_xpb_out[15][202],u_xpb_out[16][202],u_xpb_out[17][202],u_xpb_out[18][202],u_xpb_out[19][202],u_xpb_out[20][202],u_xpb_out[21][202],u_xpb_out[22][202],u_xpb_out[23][202],u_xpb_out[24][202],u_xpb_out[25][202],u_xpb_out[26][202],u_xpb_out[27][202],u_xpb_out[28][202],u_xpb_out[29][202],u_xpb_out[30][202],u_xpb_out[31][202],u_xpb_out[32][202],u_xpb_out[33][202],u_xpb_out[34][202],u_xpb_out[35][202],u_xpb_out[36][202],u_xpb_out[37][202],u_xpb_out[38][202],u_xpb_out[39][202],u_xpb_out[40][202],u_xpb_out[41][202],u_xpb_out[42][202],u_xpb_out[43][202],u_xpb_out[44][202],u_xpb_out[45][202],u_xpb_out[46][202],u_xpb_out[47][202],u_xpb_out[48][202],u_xpb_out[49][202],u_xpb_out[50][202],u_xpb_out[51][202],u_xpb_out[52][202],u_xpb_out[53][202],u_xpb_out[54][202],u_xpb_out[55][202],u_xpb_out[56][202],u_xpb_out[57][202],u_xpb_out[58][202],u_xpb_out[59][202],u_xpb_out[60][202],u_xpb_out[61][202],u_xpb_out[62][202],u_xpb_out[63][202],u_xpb_out[64][202],u_xpb_out[65][202],u_xpb_out[66][202],u_xpb_out[67][202],u_xpb_out[68][202],u_xpb_out[69][202],u_xpb_out[70][202],u_xpb_out[71][202],u_xpb_out[72][202],u_xpb_out[73][202],u_xpb_out[74][202],u_xpb_out[75][202],u_xpb_out[76][202],u_xpb_out[77][202],u_xpb_out[78][202],u_xpb_out[79][202],u_xpb_out[80][202],u_xpb_out[81][202],u_xpb_out[82][202],u_xpb_out[83][202],u_xpb_out[84][202],u_xpb_out[85][202],u_xpb_out[86][202],u_xpb_out[87][202],u_xpb_out[88][202],u_xpb_out[89][202],u_xpb_out[90][202],u_xpb_out[91][202],u_xpb_out[92][202],u_xpb_out[93][202],u_xpb_out[94][202],u_xpb_out[95][202],u_xpb_out[96][202],u_xpb_out[97][202],u_xpb_out[98][202],u_xpb_out[99][202],u_xpb_out[100][202],u_xpb_out[101][202],u_xpb_out[102][202],u_xpb_out[103][202],u_xpb_out[104][202],u_xpb_out[105][202]};

assign col_out_203 = {u_xpb_out[0][203],u_xpb_out[1][203],u_xpb_out[2][203],u_xpb_out[3][203],u_xpb_out[4][203],u_xpb_out[5][203],u_xpb_out[6][203],u_xpb_out[7][203],u_xpb_out[8][203],u_xpb_out[9][203],u_xpb_out[10][203],u_xpb_out[11][203],u_xpb_out[12][203],u_xpb_out[13][203],u_xpb_out[14][203],u_xpb_out[15][203],u_xpb_out[16][203],u_xpb_out[17][203],u_xpb_out[18][203],u_xpb_out[19][203],u_xpb_out[20][203],u_xpb_out[21][203],u_xpb_out[22][203],u_xpb_out[23][203],u_xpb_out[24][203],u_xpb_out[25][203],u_xpb_out[26][203],u_xpb_out[27][203],u_xpb_out[28][203],u_xpb_out[29][203],u_xpb_out[30][203],u_xpb_out[31][203],u_xpb_out[32][203],u_xpb_out[33][203],u_xpb_out[34][203],u_xpb_out[35][203],u_xpb_out[36][203],u_xpb_out[37][203],u_xpb_out[38][203],u_xpb_out[39][203],u_xpb_out[40][203],u_xpb_out[41][203],u_xpb_out[42][203],u_xpb_out[43][203],u_xpb_out[44][203],u_xpb_out[45][203],u_xpb_out[46][203],u_xpb_out[47][203],u_xpb_out[48][203],u_xpb_out[49][203],u_xpb_out[50][203],u_xpb_out[51][203],u_xpb_out[52][203],u_xpb_out[53][203],u_xpb_out[54][203],u_xpb_out[55][203],u_xpb_out[56][203],u_xpb_out[57][203],u_xpb_out[58][203],u_xpb_out[59][203],u_xpb_out[60][203],u_xpb_out[61][203],u_xpb_out[62][203],u_xpb_out[63][203],u_xpb_out[64][203],u_xpb_out[65][203],u_xpb_out[66][203],u_xpb_out[67][203],u_xpb_out[68][203],u_xpb_out[69][203],u_xpb_out[70][203],u_xpb_out[71][203],u_xpb_out[72][203],u_xpb_out[73][203],u_xpb_out[74][203],u_xpb_out[75][203],u_xpb_out[76][203],u_xpb_out[77][203],u_xpb_out[78][203],u_xpb_out[79][203],u_xpb_out[80][203],u_xpb_out[81][203],u_xpb_out[82][203],u_xpb_out[83][203],u_xpb_out[84][203],u_xpb_out[85][203],u_xpb_out[86][203],u_xpb_out[87][203],u_xpb_out[88][203],u_xpb_out[89][203],u_xpb_out[90][203],u_xpb_out[91][203],u_xpb_out[92][203],u_xpb_out[93][203],u_xpb_out[94][203],u_xpb_out[95][203],u_xpb_out[96][203],u_xpb_out[97][203],u_xpb_out[98][203],u_xpb_out[99][203],u_xpb_out[100][203],u_xpb_out[101][203],u_xpb_out[102][203],u_xpb_out[103][203],u_xpb_out[104][203],u_xpb_out[105][203]};

assign col_out_204 = {u_xpb_out[0][204],u_xpb_out[1][204],u_xpb_out[2][204],u_xpb_out[3][204],u_xpb_out[4][204],u_xpb_out[5][204],u_xpb_out[6][204],u_xpb_out[7][204],u_xpb_out[8][204],u_xpb_out[9][204],u_xpb_out[10][204],u_xpb_out[11][204],u_xpb_out[12][204],u_xpb_out[13][204],u_xpb_out[14][204],u_xpb_out[15][204],u_xpb_out[16][204],u_xpb_out[17][204],u_xpb_out[18][204],u_xpb_out[19][204],u_xpb_out[20][204],u_xpb_out[21][204],u_xpb_out[22][204],u_xpb_out[23][204],u_xpb_out[24][204],u_xpb_out[25][204],u_xpb_out[26][204],u_xpb_out[27][204],u_xpb_out[28][204],u_xpb_out[29][204],u_xpb_out[30][204],u_xpb_out[31][204],u_xpb_out[32][204],u_xpb_out[33][204],u_xpb_out[34][204],u_xpb_out[35][204],u_xpb_out[36][204],u_xpb_out[37][204],u_xpb_out[38][204],u_xpb_out[39][204],u_xpb_out[40][204],u_xpb_out[41][204],u_xpb_out[42][204],u_xpb_out[43][204],u_xpb_out[44][204],u_xpb_out[45][204],u_xpb_out[46][204],u_xpb_out[47][204],u_xpb_out[48][204],u_xpb_out[49][204],u_xpb_out[50][204],u_xpb_out[51][204],u_xpb_out[52][204],u_xpb_out[53][204],u_xpb_out[54][204],u_xpb_out[55][204],u_xpb_out[56][204],u_xpb_out[57][204],u_xpb_out[58][204],u_xpb_out[59][204],u_xpb_out[60][204],u_xpb_out[61][204],u_xpb_out[62][204],u_xpb_out[63][204],u_xpb_out[64][204],u_xpb_out[65][204],u_xpb_out[66][204],u_xpb_out[67][204],u_xpb_out[68][204],u_xpb_out[69][204],u_xpb_out[70][204],u_xpb_out[71][204],u_xpb_out[72][204],u_xpb_out[73][204],u_xpb_out[74][204],u_xpb_out[75][204],u_xpb_out[76][204],u_xpb_out[77][204],u_xpb_out[78][204],u_xpb_out[79][204],u_xpb_out[80][204],u_xpb_out[81][204],u_xpb_out[82][204],u_xpb_out[83][204],u_xpb_out[84][204],u_xpb_out[85][204],u_xpb_out[86][204],u_xpb_out[87][204],u_xpb_out[88][204],u_xpb_out[89][204],u_xpb_out[90][204],u_xpb_out[91][204],u_xpb_out[92][204],u_xpb_out[93][204],u_xpb_out[94][204],u_xpb_out[95][204],u_xpb_out[96][204],u_xpb_out[97][204],u_xpb_out[98][204],u_xpb_out[99][204],u_xpb_out[100][204],u_xpb_out[101][204],u_xpb_out[102][204],u_xpb_out[103][204],u_xpb_out[104][204],u_xpb_out[105][204]};

assign col_out_205 = {u_xpb_out[0][205],u_xpb_out[1][205],u_xpb_out[2][205],u_xpb_out[3][205],u_xpb_out[4][205],u_xpb_out[5][205],u_xpb_out[6][205],u_xpb_out[7][205],u_xpb_out[8][205],u_xpb_out[9][205],u_xpb_out[10][205],u_xpb_out[11][205],u_xpb_out[12][205],u_xpb_out[13][205],u_xpb_out[14][205],u_xpb_out[15][205],u_xpb_out[16][205],u_xpb_out[17][205],u_xpb_out[18][205],u_xpb_out[19][205],u_xpb_out[20][205],u_xpb_out[21][205],u_xpb_out[22][205],u_xpb_out[23][205],u_xpb_out[24][205],u_xpb_out[25][205],u_xpb_out[26][205],u_xpb_out[27][205],u_xpb_out[28][205],u_xpb_out[29][205],u_xpb_out[30][205],u_xpb_out[31][205],u_xpb_out[32][205],u_xpb_out[33][205],u_xpb_out[34][205],u_xpb_out[35][205],u_xpb_out[36][205],u_xpb_out[37][205],u_xpb_out[38][205],u_xpb_out[39][205],u_xpb_out[40][205],u_xpb_out[41][205],u_xpb_out[42][205],u_xpb_out[43][205],u_xpb_out[44][205],u_xpb_out[45][205],u_xpb_out[46][205],u_xpb_out[47][205],u_xpb_out[48][205],u_xpb_out[49][205],u_xpb_out[50][205],u_xpb_out[51][205],u_xpb_out[52][205],u_xpb_out[53][205],u_xpb_out[54][205],u_xpb_out[55][205],u_xpb_out[56][205],u_xpb_out[57][205],u_xpb_out[58][205],u_xpb_out[59][205],u_xpb_out[60][205],u_xpb_out[61][205],u_xpb_out[62][205],u_xpb_out[63][205],u_xpb_out[64][205],u_xpb_out[65][205],u_xpb_out[66][205],u_xpb_out[67][205],u_xpb_out[68][205],u_xpb_out[69][205],u_xpb_out[70][205],u_xpb_out[71][205],u_xpb_out[72][205],u_xpb_out[73][205],u_xpb_out[74][205],u_xpb_out[75][205],u_xpb_out[76][205],u_xpb_out[77][205],u_xpb_out[78][205],u_xpb_out[79][205],u_xpb_out[80][205],u_xpb_out[81][205],u_xpb_out[82][205],u_xpb_out[83][205],u_xpb_out[84][205],u_xpb_out[85][205],u_xpb_out[86][205],u_xpb_out[87][205],u_xpb_out[88][205],u_xpb_out[89][205],u_xpb_out[90][205],u_xpb_out[91][205],u_xpb_out[92][205],u_xpb_out[93][205],u_xpb_out[94][205],u_xpb_out[95][205],u_xpb_out[96][205],u_xpb_out[97][205],u_xpb_out[98][205],u_xpb_out[99][205],u_xpb_out[100][205],u_xpb_out[101][205],u_xpb_out[102][205],u_xpb_out[103][205],u_xpb_out[104][205],u_xpb_out[105][205]};

assign col_out_206 = {u_xpb_out[0][206],u_xpb_out[1][206],u_xpb_out[2][206],u_xpb_out[3][206],u_xpb_out[4][206],u_xpb_out[5][206],u_xpb_out[6][206],u_xpb_out[7][206],u_xpb_out[8][206],u_xpb_out[9][206],u_xpb_out[10][206],u_xpb_out[11][206],u_xpb_out[12][206],u_xpb_out[13][206],u_xpb_out[14][206],u_xpb_out[15][206],u_xpb_out[16][206],u_xpb_out[17][206],u_xpb_out[18][206],u_xpb_out[19][206],u_xpb_out[20][206],u_xpb_out[21][206],u_xpb_out[22][206],u_xpb_out[23][206],u_xpb_out[24][206],u_xpb_out[25][206],u_xpb_out[26][206],u_xpb_out[27][206],u_xpb_out[28][206],u_xpb_out[29][206],u_xpb_out[30][206],u_xpb_out[31][206],u_xpb_out[32][206],u_xpb_out[33][206],u_xpb_out[34][206],u_xpb_out[35][206],u_xpb_out[36][206],u_xpb_out[37][206],u_xpb_out[38][206],u_xpb_out[39][206],u_xpb_out[40][206],u_xpb_out[41][206],u_xpb_out[42][206],u_xpb_out[43][206],u_xpb_out[44][206],u_xpb_out[45][206],u_xpb_out[46][206],u_xpb_out[47][206],u_xpb_out[48][206],u_xpb_out[49][206],u_xpb_out[50][206],u_xpb_out[51][206],u_xpb_out[52][206],u_xpb_out[53][206],u_xpb_out[54][206],u_xpb_out[55][206],u_xpb_out[56][206],u_xpb_out[57][206],u_xpb_out[58][206],u_xpb_out[59][206],u_xpb_out[60][206],u_xpb_out[61][206],u_xpb_out[62][206],u_xpb_out[63][206],u_xpb_out[64][206],u_xpb_out[65][206],u_xpb_out[66][206],u_xpb_out[67][206],u_xpb_out[68][206],u_xpb_out[69][206],u_xpb_out[70][206],u_xpb_out[71][206],u_xpb_out[72][206],u_xpb_out[73][206],u_xpb_out[74][206],u_xpb_out[75][206],u_xpb_out[76][206],u_xpb_out[77][206],u_xpb_out[78][206],u_xpb_out[79][206],u_xpb_out[80][206],u_xpb_out[81][206],u_xpb_out[82][206],u_xpb_out[83][206],u_xpb_out[84][206],u_xpb_out[85][206],u_xpb_out[86][206],u_xpb_out[87][206],u_xpb_out[88][206],u_xpb_out[89][206],u_xpb_out[90][206],u_xpb_out[91][206],u_xpb_out[92][206],u_xpb_out[93][206],u_xpb_out[94][206],u_xpb_out[95][206],u_xpb_out[96][206],u_xpb_out[97][206],u_xpb_out[98][206],u_xpb_out[99][206],u_xpb_out[100][206],u_xpb_out[101][206],u_xpb_out[102][206],u_xpb_out[103][206],u_xpb_out[104][206],u_xpb_out[105][206]};

assign col_out_207 = {u_xpb_out[0][207],u_xpb_out[1][207],u_xpb_out[2][207],u_xpb_out[3][207],u_xpb_out[4][207],u_xpb_out[5][207],u_xpb_out[6][207],u_xpb_out[7][207],u_xpb_out[8][207],u_xpb_out[9][207],u_xpb_out[10][207],u_xpb_out[11][207],u_xpb_out[12][207],u_xpb_out[13][207],u_xpb_out[14][207],u_xpb_out[15][207],u_xpb_out[16][207],u_xpb_out[17][207],u_xpb_out[18][207],u_xpb_out[19][207],u_xpb_out[20][207],u_xpb_out[21][207],u_xpb_out[22][207],u_xpb_out[23][207],u_xpb_out[24][207],u_xpb_out[25][207],u_xpb_out[26][207],u_xpb_out[27][207],u_xpb_out[28][207],u_xpb_out[29][207],u_xpb_out[30][207],u_xpb_out[31][207],u_xpb_out[32][207],u_xpb_out[33][207],u_xpb_out[34][207],u_xpb_out[35][207],u_xpb_out[36][207],u_xpb_out[37][207],u_xpb_out[38][207],u_xpb_out[39][207],u_xpb_out[40][207],u_xpb_out[41][207],u_xpb_out[42][207],u_xpb_out[43][207],u_xpb_out[44][207],u_xpb_out[45][207],u_xpb_out[46][207],u_xpb_out[47][207],u_xpb_out[48][207],u_xpb_out[49][207],u_xpb_out[50][207],u_xpb_out[51][207],u_xpb_out[52][207],u_xpb_out[53][207],u_xpb_out[54][207],u_xpb_out[55][207],u_xpb_out[56][207],u_xpb_out[57][207],u_xpb_out[58][207],u_xpb_out[59][207],u_xpb_out[60][207],u_xpb_out[61][207],u_xpb_out[62][207],u_xpb_out[63][207],u_xpb_out[64][207],u_xpb_out[65][207],u_xpb_out[66][207],u_xpb_out[67][207],u_xpb_out[68][207],u_xpb_out[69][207],u_xpb_out[70][207],u_xpb_out[71][207],u_xpb_out[72][207],u_xpb_out[73][207],u_xpb_out[74][207],u_xpb_out[75][207],u_xpb_out[76][207],u_xpb_out[77][207],u_xpb_out[78][207],u_xpb_out[79][207],u_xpb_out[80][207],u_xpb_out[81][207],u_xpb_out[82][207],u_xpb_out[83][207],u_xpb_out[84][207],u_xpb_out[85][207],u_xpb_out[86][207],u_xpb_out[87][207],u_xpb_out[88][207],u_xpb_out[89][207],u_xpb_out[90][207],u_xpb_out[91][207],u_xpb_out[92][207],u_xpb_out[93][207],u_xpb_out[94][207],u_xpb_out[95][207],u_xpb_out[96][207],u_xpb_out[97][207],u_xpb_out[98][207],u_xpb_out[99][207],u_xpb_out[100][207],u_xpb_out[101][207],u_xpb_out[102][207],u_xpb_out[103][207],u_xpb_out[104][207],u_xpb_out[105][207]};

assign col_out_208 = {u_xpb_out[0][208],u_xpb_out[1][208],u_xpb_out[2][208],u_xpb_out[3][208],u_xpb_out[4][208],u_xpb_out[5][208],u_xpb_out[6][208],u_xpb_out[7][208],u_xpb_out[8][208],u_xpb_out[9][208],u_xpb_out[10][208],u_xpb_out[11][208],u_xpb_out[12][208],u_xpb_out[13][208],u_xpb_out[14][208],u_xpb_out[15][208],u_xpb_out[16][208],u_xpb_out[17][208],u_xpb_out[18][208],u_xpb_out[19][208],u_xpb_out[20][208],u_xpb_out[21][208],u_xpb_out[22][208],u_xpb_out[23][208],u_xpb_out[24][208],u_xpb_out[25][208],u_xpb_out[26][208],u_xpb_out[27][208],u_xpb_out[28][208],u_xpb_out[29][208],u_xpb_out[30][208],u_xpb_out[31][208],u_xpb_out[32][208],u_xpb_out[33][208],u_xpb_out[34][208],u_xpb_out[35][208],u_xpb_out[36][208],u_xpb_out[37][208],u_xpb_out[38][208],u_xpb_out[39][208],u_xpb_out[40][208],u_xpb_out[41][208],u_xpb_out[42][208],u_xpb_out[43][208],u_xpb_out[44][208],u_xpb_out[45][208],u_xpb_out[46][208],u_xpb_out[47][208],u_xpb_out[48][208],u_xpb_out[49][208],u_xpb_out[50][208],u_xpb_out[51][208],u_xpb_out[52][208],u_xpb_out[53][208],u_xpb_out[54][208],u_xpb_out[55][208],u_xpb_out[56][208],u_xpb_out[57][208],u_xpb_out[58][208],u_xpb_out[59][208],u_xpb_out[60][208],u_xpb_out[61][208],u_xpb_out[62][208],u_xpb_out[63][208],u_xpb_out[64][208],u_xpb_out[65][208],u_xpb_out[66][208],u_xpb_out[67][208],u_xpb_out[68][208],u_xpb_out[69][208],u_xpb_out[70][208],u_xpb_out[71][208],u_xpb_out[72][208],u_xpb_out[73][208],u_xpb_out[74][208],u_xpb_out[75][208],u_xpb_out[76][208],u_xpb_out[77][208],u_xpb_out[78][208],u_xpb_out[79][208],u_xpb_out[80][208],u_xpb_out[81][208],u_xpb_out[82][208],u_xpb_out[83][208],u_xpb_out[84][208],u_xpb_out[85][208],u_xpb_out[86][208],u_xpb_out[87][208],u_xpb_out[88][208],u_xpb_out[89][208],u_xpb_out[90][208],u_xpb_out[91][208],u_xpb_out[92][208],u_xpb_out[93][208],u_xpb_out[94][208],u_xpb_out[95][208],u_xpb_out[96][208],u_xpb_out[97][208],u_xpb_out[98][208],u_xpb_out[99][208],u_xpb_out[100][208],u_xpb_out[101][208],u_xpb_out[102][208],u_xpb_out[103][208],u_xpb_out[104][208],u_xpb_out[105][208]};

assign col_out_209 = {u_xpb_out[0][209],u_xpb_out[1][209],u_xpb_out[2][209],u_xpb_out[3][209],u_xpb_out[4][209],u_xpb_out[5][209],u_xpb_out[6][209],u_xpb_out[7][209],u_xpb_out[8][209],u_xpb_out[9][209],u_xpb_out[10][209],u_xpb_out[11][209],u_xpb_out[12][209],u_xpb_out[13][209],u_xpb_out[14][209],u_xpb_out[15][209],u_xpb_out[16][209],u_xpb_out[17][209],u_xpb_out[18][209],u_xpb_out[19][209],u_xpb_out[20][209],u_xpb_out[21][209],u_xpb_out[22][209],u_xpb_out[23][209],u_xpb_out[24][209],u_xpb_out[25][209],u_xpb_out[26][209],u_xpb_out[27][209],u_xpb_out[28][209],u_xpb_out[29][209],u_xpb_out[30][209],u_xpb_out[31][209],u_xpb_out[32][209],u_xpb_out[33][209],u_xpb_out[34][209],u_xpb_out[35][209],u_xpb_out[36][209],u_xpb_out[37][209],u_xpb_out[38][209],u_xpb_out[39][209],u_xpb_out[40][209],u_xpb_out[41][209],u_xpb_out[42][209],u_xpb_out[43][209],u_xpb_out[44][209],u_xpb_out[45][209],u_xpb_out[46][209],u_xpb_out[47][209],u_xpb_out[48][209],u_xpb_out[49][209],u_xpb_out[50][209],u_xpb_out[51][209],u_xpb_out[52][209],u_xpb_out[53][209],u_xpb_out[54][209],u_xpb_out[55][209],u_xpb_out[56][209],u_xpb_out[57][209],u_xpb_out[58][209],u_xpb_out[59][209],u_xpb_out[60][209],u_xpb_out[61][209],u_xpb_out[62][209],u_xpb_out[63][209],u_xpb_out[64][209],u_xpb_out[65][209],u_xpb_out[66][209],u_xpb_out[67][209],u_xpb_out[68][209],u_xpb_out[69][209],u_xpb_out[70][209],u_xpb_out[71][209],u_xpb_out[72][209],u_xpb_out[73][209],u_xpb_out[74][209],u_xpb_out[75][209],u_xpb_out[76][209],u_xpb_out[77][209],u_xpb_out[78][209],u_xpb_out[79][209],u_xpb_out[80][209],u_xpb_out[81][209],u_xpb_out[82][209],u_xpb_out[83][209],u_xpb_out[84][209],u_xpb_out[85][209],u_xpb_out[86][209],u_xpb_out[87][209],u_xpb_out[88][209],u_xpb_out[89][209],u_xpb_out[90][209],u_xpb_out[91][209],u_xpb_out[92][209],u_xpb_out[93][209],u_xpb_out[94][209],u_xpb_out[95][209],u_xpb_out[96][209],u_xpb_out[97][209],u_xpb_out[98][209],u_xpb_out[99][209],u_xpb_out[100][209],u_xpb_out[101][209],u_xpb_out[102][209],u_xpb_out[103][209],u_xpb_out[104][209],u_xpb_out[105][209]};

assign col_out_210 = {u_xpb_out[0][210],u_xpb_out[1][210],u_xpb_out[2][210],u_xpb_out[3][210],u_xpb_out[4][210],u_xpb_out[5][210],u_xpb_out[6][210],u_xpb_out[7][210],u_xpb_out[8][210],u_xpb_out[9][210],u_xpb_out[10][210],u_xpb_out[11][210],u_xpb_out[12][210],u_xpb_out[13][210],u_xpb_out[14][210],u_xpb_out[15][210],u_xpb_out[16][210],u_xpb_out[17][210],u_xpb_out[18][210],u_xpb_out[19][210],u_xpb_out[20][210],u_xpb_out[21][210],u_xpb_out[22][210],u_xpb_out[23][210],u_xpb_out[24][210],u_xpb_out[25][210],u_xpb_out[26][210],u_xpb_out[27][210],u_xpb_out[28][210],u_xpb_out[29][210],u_xpb_out[30][210],u_xpb_out[31][210],u_xpb_out[32][210],u_xpb_out[33][210],u_xpb_out[34][210],u_xpb_out[35][210],u_xpb_out[36][210],u_xpb_out[37][210],u_xpb_out[38][210],u_xpb_out[39][210],u_xpb_out[40][210],u_xpb_out[41][210],u_xpb_out[42][210],u_xpb_out[43][210],u_xpb_out[44][210],u_xpb_out[45][210],u_xpb_out[46][210],u_xpb_out[47][210],u_xpb_out[48][210],u_xpb_out[49][210],u_xpb_out[50][210],u_xpb_out[51][210],u_xpb_out[52][210],u_xpb_out[53][210],u_xpb_out[54][210],u_xpb_out[55][210],u_xpb_out[56][210],u_xpb_out[57][210],u_xpb_out[58][210],u_xpb_out[59][210],u_xpb_out[60][210],u_xpb_out[61][210],u_xpb_out[62][210],u_xpb_out[63][210],u_xpb_out[64][210],u_xpb_out[65][210],u_xpb_out[66][210],u_xpb_out[67][210],u_xpb_out[68][210],u_xpb_out[69][210],u_xpb_out[70][210],u_xpb_out[71][210],u_xpb_out[72][210],u_xpb_out[73][210],u_xpb_out[74][210],u_xpb_out[75][210],u_xpb_out[76][210],u_xpb_out[77][210],u_xpb_out[78][210],u_xpb_out[79][210],u_xpb_out[80][210],u_xpb_out[81][210],u_xpb_out[82][210],u_xpb_out[83][210],u_xpb_out[84][210],u_xpb_out[85][210],u_xpb_out[86][210],u_xpb_out[87][210],u_xpb_out[88][210],u_xpb_out[89][210],u_xpb_out[90][210],u_xpb_out[91][210],u_xpb_out[92][210],u_xpb_out[93][210],u_xpb_out[94][210],u_xpb_out[95][210],u_xpb_out[96][210],u_xpb_out[97][210],u_xpb_out[98][210],u_xpb_out[99][210],u_xpb_out[100][210],u_xpb_out[101][210],u_xpb_out[102][210],u_xpb_out[103][210],u_xpb_out[104][210],u_xpb_out[105][210]};

assign col_out_211 = {u_xpb_out[0][211],u_xpb_out[1][211],u_xpb_out[2][211],u_xpb_out[3][211],u_xpb_out[4][211],u_xpb_out[5][211],u_xpb_out[6][211],u_xpb_out[7][211],u_xpb_out[8][211],u_xpb_out[9][211],u_xpb_out[10][211],u_xpb_out[11][211],u_xpb_out[12][211],u_xpb_out[13][211],u_xpb_out[14][211],u_xpb_out[15][211],u_xpb_out[16][211],u_xpb_out[17][211],u_xpb_out[18][211],u_xpb_out[19][211],u_xpb_out[20][211],u_xpb_out[21][211],u_xpb_out[22][211],u_xpb_out[23][211],u_xpb_out[24][211],u_xpb_out[25][211],u_xpb_out[26][211],u_xpb_out[27][211],u_xpb_out[28][211],u_xpb_out[29][211],u_xpb_out[30][211],u_xpb_out[31][211],u_xpb_out[32][211],u_xpb_out[33][211],u_xpb_out[34][211],u_xpb_out[35][211],u_xpb_out[36][211],u_xpb_out[37][211],u_xpb_out[38][211],u_xpb_out[39][211],u_xpb_out[40][211],u_xpb_out[41][211],u_xpb_out[42][211],u_xpb_out[43][211],u_xpb_out[44][211],u_xpb_out[45][211],u_xpb_out[46][211],u_xpb_out[47][211],u_xpb_out[48][211],u_xpb_out[49][211],u_xpb_out[50][211],u_xpb_out[51][211],u_xpb_out[52][211],u_xpb_out[53][211],u_xpb_out[54][211],u_xpb_out[55][211],u_xpb_out[56][211],u_xpb_out[57][211],u_xpb_out[58][211],u_xpb_out[59][211],u_xpb_out[60][211],u_xpb_out[61][211],u_xpb_out[62][211],u_xpb_out[63][211],u_xpb_out[64][211],u_xpb_out[65][211],u_xpb_out[66][211],u_xpb_out[67][211],u_xpb_out[68][211],u_xpb_out[69][211],u_xpb_out[70][211],u_xpb_out[71][211],u_xpb_out[72][211],u_xpb_out[73][211],u_xpb_out[74][211],u_xpb_out[75][211],u_xpb_out[76][211],u_xpb_out[77][211],u_xpb_out[78][211],u_xpb_out[79][211],u_xpb_out[80][211],u_xpb_out[81][211],u_xpb_out[82][211],u_xpb_out[83][211],u_xpb_out[84][211],u_xpb_out[85][211],u_xpb_out[86][211],u_xpb_out[87][211],u_xpb_out[88][211],u_xpb_out[89][211],u_xpb_out[90][211],u_xpb_out[91][211],u_xpb_out[92][211],u_xpb_out[93][211],u_xpb_out[94][211],u_xpb_out[95][211],u_xpb_out[96][211],u_xpb_out[97][211],u_xpb_out[98][211],u_xpb_out[99][211],u_xpb_out[100][211],u_xpb_out[101][211],u_xpb_out[102][211],u_xpb_out[103][211],u_xpb_out[104][211],u_xpb_out[105][211]};

assign col_out_212 = {u_xpb_out[0][212],u_xpb_out[1][212],u_xpb_out[2][212],u_xpb_out[3][212],u_xpb_out[4][212],u_xpb_out[5][212],u_xpb_out[6][212],u_xpb_out[7][212],u_xpb_out[8][212],u_xpb_out[9][212],u_xpb_out[10][212],u_xpb_out[11][212],u_xpb_out[12][212],u_xpb_out[13][212],u_xpb_out[14][212],u_xpb_out[15][212],u_xpb_out[16][212],u_xpb_out[17][212],u_xpb_out[18][212],u_xpb_out[19][212],u_xpb_out[20][212],u_xpb_out[21][212],u_xpb_out[22][212],u_xpb_out[23][212],u_xpb_out[24][212],u_xpb_out[25][212],u_xpb_out[26][212],u_xpb_out[27][212],u_xpb_out[28][212],u_xpb_out[29][212],u_xpb_out[30][212],u_xpb_out[31][212],u_xpb_out[32][212],u_xpb_out[33][212],u_xpb_out[34][212],u_xpb_out[35][212],u_xpb_out[36][212],u_xpb_out[37][212],u_xpb_out[38][212],u_xpb_out[39][212],u_xpb_out[40][212],u_xpb_out[41][212],u_xpb_out[42][212],u_xpb_out[43][212],u_xpb_out[44][212],u_xpb_out[45][212],u_xpb_out[46][212],u_xpb_out[47][212],u_xpb_out[48][212],u_xpb_out[49][212],u_xpb_out[50][212],u_xpb_out[51][212],u_xpb_out[52][212],u_xpb_out[53][212],u_xpb_out[54][212],u_xpb_out[55][212],u_xpb_out[56][212],u_xpb_out[57][212],u_xpb_out[58][212],u_xpb_out[59][212],u_xpb_out[60][212],u_xpb_out[61][212],u_xpb_out[62][212],u_xpb_out[63][212],u_xpb_out[64][212],u_xpb_out[65][212],u_xpb_out[66][212],u_xpb_out[67][212],u_xpb_out[68][212],u_xpb_out[69][212],u_xpb_out[70][212],u_xpb_out[71][212],u_xpb_out[72][212],u_xpb_out[73][212],u_xpb_out[74][212],u_xpb_out[75][212],u_xpb_out[76][212],u_xpb_out[77][212],u_xpb_out[78][212],u_xpb_out[79][212],u_xpb_out[80][212],u_xpb_out[81][212],u_xpb_out[82][212],u_xpb_out[83][212],u_xpb_out[84][212],u_xpb_out[85][212],u_xpb_out[86][212],u_xpb_out[87][212],u_xpb_out[88][212],u_xpb_out[89][212],u_xpb_out[90][212],u_xpb_out[91][212],u_xpb_out[92][212],u_xpb_out[93][212],u_xpb_out[94][212],u_xpb_out[95][212],u_xpb_out[96][212],u_xpb_out[97][212],u_xpb_out[98][212],u_xpb_out[99][212],u_xpb_out[100][212],u_xpb_out[101][212],u_xpb_out[102][212],u_xpb_out[103][212],u_xpb_out[104][212],u_xpb_out[105][212]};

assign col_out_213 = {u_xpb_out[0][213],u_xpb_out[1][213],u_xpb_out[2][213],u_xpb_out[3][213],u_xpb_out[4][213],u_xpb_out[5][213],u_xpb_out[6][213],u_xpb_out[7][213],u_xpb_out[8][213],u_xpb_out[9][213],u_xpb_out[10][213],u_xpb_out[11][213],u_xpb_out[12][213],u_xpb_out[13][213],u_xpb_out[14][213],u_xpb_out[15][213],u_xpb_out[16][213],u_xpb_out[17][213],u_xpb_out[18][213],u_xpb_out[19][213],u_xpb_out[20][213],u_xpb_out[21][213],u_xpb_out[22][213],u_xpb_out[23][213],u_xpb_out[24][213],u_xpb_out[25][213],u_xpb_out[26][213],u_xpb_out[27][213],u_xpb_out[28][213],u_xpb_out[29][213],u_xpb_out[30][213],u_xpb_out[31][213],u_xpb_out[32][213],u_xpb_out[33][213],u_xpb_out[34][213],u_xpb_out[35][213],u_xpb_out[36][213],u_xpb_out[37][213],u_xpb_out[38][213],u_xpb_out[39][213],u_xpb_out[40][213],u_xpb_out[41][213],u_xpb_out[42][213],u_xpb_out[43][213],u_xpb_out[44][213],u_xpb_out[45][213],u_xpb_out[46][213],u_xpb_out[47][213],u_xpb_out[48][213],u_xpb_out[49][213],u_xpb_out[50][213],u_xpb_out[51][213],u_xpb_out[52][213],u_xpb_out[53][213],u_xpb_out[54][213],u_xpb_out[55][213],u_xpb_out[56][213],u_xpb_out[57][213],u_xpb_out[58][213],u_xpb_out[59][213],u_xpb_out[60][213],u_xpb_out[61][213],u_xpb_out[62][213],u_xpb_out[63][213],u_xpb_out[64][213],u_xpb_out[65][213],u_xpb_out[66][213],u_xpb_out[67][213],u_xpb_out[68][213],u_xpb_out[69][213],u_xpb_out[70][213],u_xpb_out[71][213],u_xpb_out[72][213],u_xpb_out[73][213],u_xpb_out[74][213],u_xpb_out[75][213],u_xpb_out[76][213],u_xpb_out[77][213],u_xpb_out[78][213],u_xpb_out[79][213],u_xpb_out[80][213],u_xpb_out[81][213],u_xpb_out[82][213],u_xpb_out[83][213],u_xpb_out[84][213],u_xpb_out[85][213],u_xpb_out[86][213],u_xpb_out[87][213],u_xpb_out[88][213],u_xpb_out[89][213],u_xpb_out[90][213],u_xpb_out[91][213],u_xpb_out[92][213],u_xpb_out[93][213],u_xpb_out[94][213],u_xpb_out[95][213],u_xpb_out[96][213],u_xpb_out[97][213],u_xpb_out[98][213],u_xpb_out[99][213],u_xpb_out[100][213],u_xpb_out[101][213],u_xpb_out[102][213],u_xpb_out[103][213],u_xpb_out[104][213],u_xpb_out[105][213]};

assign col_out_214 = {u_xpb_out[0][214],u_xpb_out[1][214],u_xpb_out[2][214],u_xpb_out[3][214],u_xpb_out[4][214],u_xpb_out[5][214],u_xpb_out[6][214],u_xpb_out[7][214],u_xpb_out[8][214],u_xpb_out[9][214],u_xpb_out[10][214],u_xpb_out[11][214],u_xpb_out[12][214],u_xpb_out[13][214],u_xpb_out[14][214],u_xpb_out[15][214],u_xpb_out[16][214],u_xpb_out[17][214],u_xpb_out[18][214],u_xpb_out[19][214],u_xpb_out[20][214],u_xpb_out[21][214],u_xpb_out[22][214],u_xpb_out[23][214],u_xpb_out[24][214],u_xpb_out[25][214],u_xpb_out[26][214],u_xpb_out[27][214],u_xpb_out[28][214],u_xpb_out[29][214],u_xpb_out[30][214],u_xpb_out[31][214],u_xpb_out[32][214],u_xpb_out[33][214],u_xpb_out[34][214],u_xpb_out[35][214],u_xpb_out[36][214],u_xpb_out[37][214],u_xpb_out[38][214],u_xpb_out[39][214],u_xpb_out[40][214],u_xpb_out[41][214],u_xpb_out[42][214],u_xpb_out[43][214],u_xpb_out[44][214],u_xpb_out[45][214],u_xpb_out[46][214],u_xpb_out[47][214],u_xpb_out[48][214],u_xpb_out[49][214],u_xpb_out[50][214],u_xpb_out[51][214],u_xpb_out[52][214],u_xpb_out[53][214],u_xpb_out[54][214],u_xpb_out[55][214],u_xpb_out[56][214],u_xpb_out[57][214],u_xpb_out[58][214],u_xpb_out[59][214],u_xpb_out[60][214],u_xpb_out[61][214],u_xpb_out[62][214],u_xpb_out[63][214],u_xpb_out[64][214],u_xpb_out[65][214],u_xpb_out[66][214],u_xpb_out[67][214],u_xpb_out[68][214],u_xpb_out[69][214],u_xpb_out[70][214],u_xpb_out[71][214],u_xpb_out[72][214],u_xpb_out[73][214],u_xpb_out[74][214],u_xpb_out[75][214],u_xpb_out[76][214],u_xpb_out[77][214],u_xpb_out[78][214],u_xpb_out[79][214],u_xpb_out[80][214],u_xpb_out[81][214],u_xpb_out[82][214],u_xpb_out[83][214],u_xpb_out[84][214],u_xpb_out[85][214],u_xpb_out[86][214],u_xpb_out[87][214],u_xpb_out[88][214],u_xpb_out[89][214],u_xpb_out[90][214],u_xpb_out[91][214],u_xpb_out[92][214],u_xpb_out[93][214],u_xpb_out[94][214],u_xpb_out[95][214],u_xpb_out[96][214],u_xpb_out[97][214],u_xpb_out[98][214],u_xpb_out[99][214],u_xpb_out[100][214],u_xpb_out[101][214],u_xpb_out[102][214],u_xpb_out[103][214],u_xpb_out[104][214],u_xpb_out[105][214]};

assign col_out_215 = {u_xpb_out[0][215],u_xpb_out[1][215],u_xpb_out[2][215],u_xpb_out[3][215],u_xpb_out[4][215],u_xpb_out[5][215],u_xpb_out[6][215],u_xpb_out[7][215],u_xpb_out[8][215],u_xpb_out[9][215],u_xpb_out[10][215],u_xpb_out[11][215],u_xpb_out[12][215],u_xpb_out[13][215],u_xpb_out[14][215],u_xpb_out[15][215],u_xpb_out[16][215],u_xpb_out[17][215],u_xpb_out[18][215],u_xpb_out[19][215],u_xpb_out[20][215],u_xpb_out[21][215],u_xpb_out[22][215],u_xpb_out[23][215],u_xpb_out[24][215],u_xpb_out[25][215],u_xpb_out[26][215],u_xpb_out[27][215],u_xpb_out[28][215],u_xpb_out[29][215],u_xpb_out[30][215],u_xpb_out[31][215],u_xpb_out[32][215],u_xpb_out[33][215],u_xpb_out[34][215],u_xpb_out[35][215],u_xpb_out[36][215],u_xpb_out[37][215],u_xpb_out[38][215],u_xpb_out[39][215],u_xpb_out[40][215],u_xpb_out[41][215],u_xpb_out[42][215],u_xpb_out[43][215],u_xpb_out[44][215],u_xpb_out[45][215],u_xpb_out[46][215],u_xpb_out[47][215],u_xpb_out[48][215],u_xpb_out[49][215],u_xpb_out[50][215],u_xpb_out[51][215],u_xpb_out[52][215],u_xpb_out[53][215],u_xpb_out[54][215],u_xpb_out[55][215],u_xpb_out[56][215],u_xpb_out[57][215],u_xpb_out[58][215],u_xpb_out[59][215],u_xpb_out[60][215],u_xpb_out[61][215],u_xpb_out[62][215],u_xpb_out[63][215],u_xpb_out[64][215],u_xpb_out[65][215],u_xpb_out[66][215],u_xpb_out[67][215],u_xpb_out[68][215],u_xpb_out[69][215],u_xpb_out[70][215],u_xpb_out[71][215],u_xpb_out[72][215],u_xpb_out[73][215],u_xpb_out[74][215],u_xpb_out[75][215],u_xpb_out[76][215],u_xpb_out[77][215],u_xpb_out[78][215],u_xpb_out[79][215],u_xpb_out[80][215],u_xpb_out[81][215],u_xpb_out[82][215],u_xpb_out[83][215],u_xpb_out[84][215],u_xpb_out[85][215],u_xpb_out[86][215],u_xpb_out[87][215],u_xpb_out[88][215],u_xpb_out[89][215],u_xpb_out[90][215],u_xpb_out[91][215],u_xpb_out[92][215],u_xpb_out[93][215],u_xpb_out[94][215],u_xpb_out[95][215],u_xpb_out[96][215],u_xpb_out[97][215],u_xpb_out[98][215],u_xpb_out[99][215],u_xpb_out[100][215],u_xpb_out[101][215],u_xpb_out[102][215],u_xpb_out[103][215],u_xpb_out[104][215],u_xpb_out[105][215]};

assign col_out_216 = {u_xpb_out[0][216],u_xpb_out[1][216],u_xpb_out[2][216],u_xpb_out[3][216],u_xpb_out[4][216],u_xpb_out[5][216],u_xpb_out[6][216],u_xpb_out[7][216],u_xpb_out[8][216],u_xpb_out[9][216],u_xpb_out[10][216],u_xpb_out[11][216],u_xpb_out[12][216],u_xpb_out[13][216],u_xpb_out[14][216],u_xpb_out[15][216],u_xpb_out[16][216],u_xpb_out[17][216],u_xpb_out[18][216],u_xpb_out[19][216],u_xpb_out[20][216],u_xpb_out[21][216],u_xpb_out[22][216],u_xpb_out[23][216],u_xpb_out[24][216],u_xpb_out[25][216],u_xpb_out[26][216],u_xpb_out[27][216],u_xpb_out[28][216],u_xpb_out[29][216],u_xpb_out[30][216],u_xpb_out[31][216],u_xpb_out[32][216],u_xpb_out[33][216],u_xpb_out[34][216],u_xpb_out[35][216],u_xpb_out[36][216],u_xpb_out[37][216],u_xpb_out[38][216],u_xpb_out[39][216],u_xpb_out[40][216],u_xpb_out[41][216],u_xpb_out[42][216],u_xpb_out[43][216],u_xpb_out[44][216],u_xpb_out[45][216],u_xpb_out[46][216],u_xpb_out[47][216],u_xpb_out[48][216],u_xpb_out[49][216],u_xpb_out[50][216],u_xpb_out[51][216],u_xpb_out[52][216],u_xpb_out[53][216],u_xpb_out[54][216],u_xpb_out[55][216],u_xpb_out[56][216],u_xpb_out[57][216],u_xpb_out[58][216],u_xpb_out[59][216],u_xpb_out[60][216],u_xpb_out[61][216],u_xpb_out[62][216],u_xpb_out[63][216],u_xpb_out[64][216],u_xpb_out[65][216],u_xpb_out[66][216],u_xpb_out[67][216],u_xpb_out[68][216],u_xpb_out[69][216],u_xpb_out[70][216],u_xpb_out[71][216],u_xpb_out[72][216],u_xpb_out[73][216],u_xpb_out[74][216],u_xpb_out[75][216],u_xpb_out[76][216],u_xpb_out[77][216],u_xpb_out[78][216],u_xpb_out[79][216],u_xpb_out[80][216],u_xpb_out[81][216],u_xpb_out[82][216],u_xpb_out[83][216],u_xpb_out[84][216],u_xpb_out[85][216],u_xpb_out[86][216],u_xpb_out[87][216],u_xpb_out[88][216],u_xpb_out[89][216],u_xpb_out[90][216],u_xpb_out[91][216],u_xpb_out[92][216],u_xpb_out[93][216],u_xpb_out[94][216],u_xpb_out[95][216],u_xpb_out[96][216],u_xpb_out[97][216],u_xpb_out[98][216],u_xpb_out[99][216],u_xpb_out[100][216],u_xpb_out[101][216],u_xpb_out[102][216],u_xpb_out[103][216],u_xpb_out[104][216],u_xpb_out[105][216]};

assign col_out_217 = {u_xpb_out[0][217],u_xpb_out[1][217],u_xpb_out[2][217],u_xpb_out[3][217],u_xpb_out[4][217],u_xpb_out[5][217],u_xpb_out[6][217],u_xpb_out[7][217],u_xpb_out[8][217],u_xpb_out[9][217],u_xpb_out[10][217],u_xpb_out[11][217],u_xpb_out[12][217],u_xpb_out[13][217],u_xpb_out[14][217],u_xpb_out[15][217],u_xpb_out[16][217],u_xpb_out[17][217],u_xpb_out[18][217],u_xpb_out[19][217],u_xpb_out[20][217],u_xpb_out[21][217],u_xpb_out[22][217],u_xpb_out[23][217],u_xpb_out[24][217],u_xpb_out[25][217],u_xpb_out[26][217],u_xpb_out[27][217],u_xpb_out[28][217],u_xpb_out[29][217],u_xpb_out[30][217],u_xpb_out[31][217],u_xpb_out[32][217],u_xpb_out[33][217],u_xpb_out[34][217],u_xpb_out[35][217],u_xpb_out[36][217],u_xpb_out[37][217],u_xpb_out[38][217],u_xpb_out[39][217],u_xpb_out[40][217],u_xpb_out[41][217],u_xpb_out[42][217],u_xpb_out[43][217],u_xpb_out[44][217],u_xpb_out[45][217],u_xpb_out[46][217],u_xpb_out[47][217],u_xpb_out[48][217],u_xpb_out[49][217],u_xpb_out[50][217],u_xpb_out[51][217],u_xpb_out[52][217],u_xpb_out[53][217],u_xpb_out[54][217],u_xpb_out[55][217],u_xpb_out[56][217],u_xpb_out[57][217],u_xpb_out[58][217],u_xpb_out[59][217],u_xpb_out[60][217],u_xpb_out[61][217],u_xpb_out[62][217],u_xpb_out[63][217],u_xpb_out[64][217],u_xpb_out[65][217],u_xpb_out[66][217],u_xpb_out[67][217],u_xpb_out[68][217],u_xpb_out[69][217],u_xpb_out[70][217],u_xpb_out[71][217],u_xpb_out[72][217],u_xpb_out[73][217],u_xpb_out[74][217],u_xpb_out[75][217],u_xpb_out[76][217],u_xpb_out[77][217],u_xpb_out[78][217],u_xpb_out[79][217],u_xpb_out[80][217],u_xpb_out[81][217],u_xpb_out[82][217],u_xpb_out[83][217],u_xpb_out[84][217],u_xpb_out[85][217],u_xpb_out[86][217],u_xpb_out[87][217],u_xpb_out[88][217],u_xpb_out[89][217],u_xpb_out[90][217],u_xpb_out[91][217],u_xpb_out[92][217],u_xpb_out[93][217],u_xpb_out[94][217],u_xpb_out[95][217],u_xpb_out[96][217],u_xpb_out[97][217],u_xpb_out[98][217],u_xpb_out[99][217],u_xpb_out[100][217],u_xpb_out[101][217],u_xpb_out[102][217],u_xpb_out[103][217],u_xpb_out[104][217],u_xpb_out[105][217]};

assign col_out_218 = {u_xpb_out[0][218],u_xpb_out[1][218],u_xpb_out[2][218],u_xpb_out[3][218],u_xpb_out[4][218],u_xpb_out[5][218],u_xpb_out[6][218],u_xpb_out[7][218],u_xpb_out[8][218],u_xpb_out[9][218],u_xpb_out[10][218],u_xpb_out[11][218],u_xpb_out[12][218],u_xpb_out[13][218],u_xpb_out[14][218],u_xpb_out[15][218],u_xpb_out[16][218],u_xpb_out[17][218],u_xpb_out[18][218],u_xpb_out[19][218],u_xpb_out[20][218],u_xpb_out[21][218],u_xpb_out[22][218],u_xpb_out[23][218],u_xpb_out[24][218],u_xpb_out[25][218],u_xpb_out[26][218],u_xpb_out[27][218],u_xpb_out[28][218],u_xpb_out[29][218],u_xpb_out[30][218],u_xpb_out[31][218],u_xpb_out[32][218],u_xpb_out[33][218],u_xpb_out[34][218],u_xpb_out[35][218],u_xpb_out[36][218],u_xpb_out[37][218],u_xpb_out[38][218],u_xpb_out[39][218],u_xpb_out[40][218],u_xpb_out[41][218],u_xpb_out[42][218],u_xpb_out[43][218],u_xpb_out[44][218],u_xpb_out[45][218],u_xpb_out[46][218],u_xpb_out[47][218],u_xpb_out[48][218],u_xpb_out[49][218],u_xpb_out[50][218],u_xpb_out[51][218],u_xpb_out[52][218],u_xpb_out[53][218],u_xpb_out[54][218],u_xpb_out[55][218],u_xpb_out[56][218],u_xpb_out[57][218],u_xpb_out[58][218],u_xpb_out[59][218],u_xpb_out[60][218],u_xpb_out[61][218],u_xpb_out[62][218],u_xpb_out[63][218],u_xpb_out[64][218],u_xpb_out[65][218],u_xpb_out[66][218],u_xpb_out[67][218],u_xpb_out[68][218],u_xpb_out[69][218],u_xpb_out[70][218],u_xpb_out[71][218],u_xpb_out[72][218],u_xpb_out[73][218],u_xpb_out[74][218],u_xpb_out[75][218],u_xpb_out[76][218],u_xpb_out[77][218],u_xpb_out[78][218],u_xpb_out[79][218],u_xpb_out[80][218],u_xpb_out[81][218],u_xpb_out[82][218],u_xpb_out[83][218],u_xpb_out[84][218],u_xpb_out[85][218],u_xpb_out[86][218],u_xpb_out[87][218],u_xpb_out[88][218],u_xpb_out[89][218],u_xpb_out[90][218],u_xpb_out[91][218],u_xpb_out[92][218],u_xpb_out[93][218],u_xpb_out[94][218],u_xpb_out[95][218],u_xpb_out[96][218],u_xpb_out[97][218],u_xpb_out[98][218],u_xpb_out[99][218],u_xpb_out[100][218],u_xpb_out[101][218],u_xpb_out[102][218],u_xpb_out[103][218],u_xpb_out[104][218],u_xpb_out[105][218]};

assign col_out_219 = {u_xpb_out[0][219],u_xpb_out[1][219],u_xpb_out[2][219],u_xpb_out[3][219],u_xpb_out[4][219],u_xpb_out[5][219],u_xpb_out[6][219],u_xpb_out[7][219],u_xpb_out[8][219],u_xpb_out[9][219],u_xpb_out[10][219],u_xpb_out[11][219],u_xpb_out[12][219],u_xpb_out[13][219],u_xpb_out[14][219],u_xpb_out[15][219],u_xpb_out[16][219],u_xpb_out[17][219],u_xpb_out[18][219],u_xpb_out[19][219],u_xpb_out[20][219],u_xpb_out[21][219],u_xpb_out[22][219],u_xpb_out[23][219],u_xpb_out[24][219],u_xpb_out[25][219],u_xpb_out[26][219],u_xpb_out[27][219],u_xpb_out[28][219],u_xpb_out[29][219],u_xpb_out[30][219],u_xpb_out[31][219],u_xpb_out[32][219],u_xpb_out[33][219],u_xpb_out[34][219],u_xpb_out[35][219],u_xpb_out[36][219],u_xpb_out[37][219],u_xpb_out[38][219],u_xpb_out[39][219],u_xpb_out[40][219],u_xpb_out[41][219],u_xpb_out[42][219],u_xpb_out[43][219],u_xpb_out[44][219],u_xpb_out[45][219],u_xpb_out[46][219],u_xpb_out[47][219],u_xpb_out[48][219],u_xpb_out[49][219],u_xpb_out[50][219],u_xpb_out[51][219],u_xpb_out[52][219],u_xpb_out[53][219],u_xpb_out[54][219],u_xpb_out[55][219],u_xpb_out[56][219],u_xpb_out[57][219],u_xpb_out[58][219],u_xpb_out[59][219],u_xpb_out[60][219],u_xpb_out[61][219],u_xpb_out[62][219],u_xpb_out[63][219],u_xpb_out[64][219],u_xpb_out[65][219],u_xpb_out[66][219],u_xpb_out[67][219],u_xpb_out[68][219],u_xpb_out[69][219],u_xpb_out[70][219],u_xpb_out[71][219],u_xpb_out[72][219],u_xpb_out[73][219],u_xpb_out[74][219],u_xpb_out[75][219],u_xpb_out[76][219],u_xpb_out[77][219],u_xpb_out[78][219],u_xpb_out[79][219],u_xpb_out[80][219],u_xpb_out[81][219],u_xpb_out[82][219],u_xpb_out[83][219],u_xpb_out[84][219],u_xpb_out[85][219],u_xpb_out[86][219],u_xpb_out[87][219],u_xpb_out[88][219],u_xpb_out[89][219],u_xpb_out[90][219],u_xpb_out[91][219],u_xpb_out[92][219],u_xpb_out[93][219],u_xpb_out[94][219],u_xpb_out[95][219],u_xpb_out[96][219],u_xpb_out[97][219],u_xpb_out[98][219],u_xpb_out[99][219],u_xpb_out[100][219],u_xpb_out[101][219],u_xpb_out[102][219],u_xpb_out[103][219],u_xpb_out[104][219],u_xpb_out[105][219]};

assign col_out_220 = {u_xpb_out[0][220],u_xpb_out[1][220],u_xpb_out[2][220],u_xpb_out[3][220],u_xpb_out[4][220],u_xpb_out[5][220],u_xpb_out[6][220],u_xpb_out[7][220],u_xpb_out[8][220],u_xpb_out[9][220],u_xpb_out[10][220],u_xpb_out[11][220],u_xpb_out[12][220],u_xpb_out[13][220],u_xpb_out[14][220],u_xpb_out[15][220],u_xpb_out[16][220],u_xpb_out[17][220],u_xpb_out[18][220],u_xpb_out[19][220],u_xpb_out[20][220],u_xpb_out[21][220],u_xpb_out[22][220],u_xpb_out[23][220],u_xpb_out[24][220],u_xpb_out[25][220],u_xpb_out[26][220],u_xpb_out[27][220],u_xpb_out[28][220],u_xpb_out[29][220],u_xpb_out[30][220],u_xpb_out[31][220],u_xpb_out[32][220],u_xpb_out[33][220],u_xpb_out[34][220],u_xpb_out[35][220],u_xpb_out[36][220],u_xpb_out[37][220],u_xpb_out[38][220],u_xpb_out[39][220],u_xpb_out[40][220],u_xpb_out[41][220],u_xpb_out[42][220],u_xpb_out[43][220],u_xpb_out[44][220],u_xpb_out[45][220],u_xpb_out[46][220],u_xpb_out[47][220],u_xpb_out[48][220],u_xpb_out[49][220],u_xpb_out[50][220],u_xpb_out[51][220],u_xpb_out[52][220],u_xpb_out[53][220],u_xpb_out[54][220],u_xpb_out[55][220],u_xpb_out[56][220],u_xpb_out[57][220],u_xpb_out[58][220],u_xpb_out[59][220],u_xpb_out[60][220],u_xpb_out[61][220],u_xpb_out[62][220],u_xpb_out[63][220],u_xpb_out[64][220],u_xpb_out[65][220],u_xpb_out[66][220],u_xpb_out[67][220],u_xpb_out[68][220],u_xpb_out[69][220],u_xpb_out[70][220],u_xpb_out[71][220],u_xpb_out[72][220],u_xpb_out[73][220],u_xpb_out[74][220],u_xpb_out[75][220],u_xpb_out[76][220],u_xpb_out[77][220],u_xpb_out[78][220],u_xpb_out[79][220],u_xpb_out[80][220],u_xpb_out[81][220],u_xpb_out[82][220],u_xpb_out[83][220],u_xpb_out[84][220],u_xpb_out[85][220],u_xpb_out[86][220],u_xpb_out[87][220],u_xpb_out[88][220],u_xpb_out[89][220],u_xpb_out[90][220],u_xpb_out[91][220],u_xpb_out[92][220],u_xpb_out[93][220],u_xpb_out[94][220],u_xpb_out[95][220],u_xpb_out[96][220],u_xpb_out[97][220],u_xpb_out[98][220],u_xpb_out[99][220],u_xpb_out[100][220],u_xpb_out[101][220],u_xpb_out[102][220],u_xpb_out[103][220],u_xpb_out[104][220],u_xpb_out[105][220]};

assign col_out_221 = {u_xpb_out[0][221],u_xpb_out[1][221],u_xpb_out[2][221],u_xpb_out[3][221],u_xpb_out[4][221],u_xpb_out[5][221],u_xpb_out[6][221],u_xpb_out[7][221],u_xpb_out[8][221],u_xpb_out[9][221],u_xpb_out[10][221],u_xpb_out[11][221],u_xpb_out[12][221],u_xpb_out[13][221],u_xpb_out[14][221],u_xpb_out[15][221],u_xpb_out[16][221],u_xpb_out[17][221],u_xpb_out[18][221],u_xpb_out[19][221],u_xpb_out[20][221],u_xpb_out[21][221],u_xpb_out[22][221],u_xpb_out[23][221],u_xpb_out[24][221],u_xpb_out[25][221],u_xpb_out[26][221],u_xpb_out[27][221],u_xpb_out[28][221],u_xpb_out[29][221],u_xpb_out[30][221],u_xpb_out[31][221],u_xpb_out[32][221],u_xpb_out[33][221],u_xpb_out[34][221],u_xpb_out[35][221],u_xpb_out[36][221],u_xpb_out[37][221],u_xpb_out[38][221],u_xpb_out[39][221],u_xpb_out[40][221],u_xpb_out[41][221],u_xpb_out[42][221],u_xpb_out[43][221],u_xpb_out[44][221],u_xpb_out[45][221],u_xpb_out[46][221],u_xpb_out[47][221],u_xpb_out[48][221],u_xpb_out[49][221],u_xpb_out[50][221],u_xpb_out[51][221],u_xpb_out[52][221],u_xpb_out[53][221],u_xpb_out[54][221],u_xpb_out[55][221],u_xpb_out[56][221],u_xpb_out[57][221],u_xpb_out[58][221],u_xpb_out[59][221],u_xpb_out[60][221],u_xpb_out[61][221],u_xpb_out[62][221],u_xpb_out[63][221],u_xpb_out[64][221],u_xpb_out[65][221],u_xpb_out[66][221],u_xpb_out[67][221],u_xpb_out[68][221],u_xpb_out[69][221],u_xpb_out[70][221],u_xpb_out[71][221],u_xpb_out[72][221],u_xpb_out[73][221],u_xpb_out[74][221],u_xpb_out[75][221],u_xpb_out[76][221],u_xpb_out[77][221],u_xpb_out[78][221],u_xpb_out[79][221],u_xpb_out[80][221],u_xpb_out[81][221],u_xpb_out[82][221],u_xpb_out[83][221],u_xpb_out[84][221],u_xpb_out[85][221],u_xpb_out[86][221],u_xpb_out[87][221],u_xpb_out[88][221],u_xpb_out[89][221],u_xpb_out[90][221],u_xpb_out[91][221],u_xpb_out[92][221],u_xpb_out[93][221],u_xpb_out[94][221],u_xpb_out[95][221],u_xpb_out[96][221],u_xpb_out[97][221],u_xpb_out[98][221],u_xpb_out[99][221],u_xpb_out[100][221],u_xpb_out[101][221],u_xpb_out[102][221],u_xpb_out[103][221],u_xpb_out[104][221],u_xpb_out[105][221]};

assign col_out_222 = {u_xpb_out[0][222],u_xpb_out[1][222],u_xpb_out[2][222],u_xpb_out[3][222],u_xpb_out[4][222],u_xpb_out[5][222],u_xpb_out[6][222],u_xpb_out[7][222],u_xpb_out[8][222],u_xpb_out[9][222],u_xpb_out[10][222],u_xpb_out[11][222],u_xpb_out[12][222],u_xpb_out[13][222],u_xpb_out[14][222],u_xpb_out[15][222],u_xpb_out[16][222],u_xpb_out[17][222],u_xpb_out[18][222],u_xpb_out[19][222],u_xpb_out[20][222],u_xpb_out[21][222],u_xpb_out[22][222],u_xpb_out[23][222],u_xpb_out[24][222],u_xpb_out[25][222],u_xpb_out[26][222],u_xpb_out[27][222],u_xpb_out[28][222],u_xpb_out[29][222],u_xpb_out[30][222],u_xpb_out[31][222],u_xpb_out[32][222],u_xpb_out[33][222],u_xpb_out[34][222],u_xpb_out[35][222],u_xpb_out[36][222],u_xpb_out[37][222],u_xpb_out[38][222],u_xpb_out[39][222],u_xpb_out[40][222],u_xpb_out[41][222],u_xpb_out[42][222],u_xpb_out[43][222],u_xpb_out[44][222],u_xpb_out[45][222],u_xpb_out[46][222],u_xpb_out[47][222],u_xpb_out[48][222],u_xpb_out[49][222],u_xpb_out[50][222],u_xpb_out[51][222],u_xpb_out[52][222],u_xpb_out[53][222],u_xpb_out[54][222],u_xpb_out[55][222],u_xpb_out[56][222],u_xpb_out[57][222],u_xpb_out[58][222],u_xpb_out[59][222],u_xpb_out[60][222],u_xpb_out[61][222],u_xpb_out[62][222],u_xpb_out[63][222],u_xpb_out[64][222],u_xpb_out[65][222],u_xpb_out[66][222],u_xpb_out[67][222],u_xpb_out[68][222],u_xpb_out[69][222],u_xpb_out[70][222],u_xpb_out[71][222],u_xpb_out[72][222],u_xpb_out[73][222],u_xpb_out[74][222],u_xpb_out[75][222],u_xpb_out[76][222],u_xpb_out[77][222],u_xpb_out[78][222],u_xpb_out[79][222],u_xpb_out[80][222],u_xpb_out[81][222],u_xpb_out[82][222],u_xpb_out[83][222],u_xpb_out[84][222],u_xpb_out[85][222],u_xpb_out[86][222],u_xpb_out[87][222],u_xpb_out[88][222],u_xpb_out[89][222],u_xpb_out[90][222],u_xpb_out[91][222],u_xpb_out[92][222],u_xpb_out[93][222],u_xpb_out[94][222],u_xpb_out[95][222],u_xpb_out[96][222],u_xpb_out[97][222],u_xpb_out[98][222],u_xpb_out[99][222],u_xpb_out[100][222],u_xpb_out[101][222],u_xpb_out[102][222],u_xpb_out[103][222],u_xpb_out[104][222],u_xpb_out[105][222]};

assign col_out_223 = {u_xpb_out[0][223],u_xpb_out[1][223],u_xpb_out[2][223],u_xpb_out[3][223],u_xpb_out[4][223],u_xpb_out[5][223],u_xpb_out[6][223],u_xpb_out[7][223],u_xpb_out[8][223],u_xpb_out[9][223],u_xpb_out[10][223],u_xpb_out[11][223],u_xpb_out[12][223],u_xpb_out[13][223],u_xpb_out[14][223],u_xpb_out[15][223],u_xpb_out[16][223],u_xpb_out[17][223],u_xpb_out[18][223],u_xpb_out[19][223],u_xpb_out[20][223],u_xpb_out[21][223],u_xpb_out[22][223],u_xpb_out[23][223],u_xpb_out[24][223],u_xpb_out[25][223],u_xpb_out[26][223],u_xpb_out[27][223],u_xpb_out[28][223],u_xpb_out[29][223],u_xpb_out[30][223],u_xpb_out[31][223],u_xpb_out[32][223],u_xpb_out[33][223],u_xpb_out[34][223],u_xpb_out[35][223],u_xpb_out[36][223],u_xpb_out[37][223],u_xpb_out[38][223],u_xpb_out[39][223],u_xpb_out[40][223],u_xpb_out[41][223],u_xpb_out[42][223],u_xpb_out[43][223],u_xpb_out[44][223],u_xpb_out[45][223],u_xpb_out[46][223],u_xpb_out[47][223],u_xpb_out[48][223],u_xpb_out[49][223],u_xpb_out[50][223],u_xpb_out[51][223],u_xpb_out[52][223],u_xpb_out[53][223],u_xpb_out[54][223],u_xpb_out[55][223],u_xpb_out[56][223],u_xpb_out[57][223],u_xpb_out[58][223],u_xpb_out[59][223],u_xpb_out[60][223],u_xpb_out[61][223],u_xpb_out[62][223],u_xpb_out[63][223],u_xpb_out[64][223],u_xpb_out[65][223],u_xpb_out[66][223],u_xpb_out[67][223],u_xpb_out[68][223],u_xpb_out[69][223],u_xpb_out[70][223],u_xpb_out[71][223],u_xpb_out[72][223],u_xpb_out[73][223],u_xpb_out[74][223],u_xpb_out[75][223],u_xpb_out[76][223],u_xpb_out[77][223],u_xpb_out[78][223],u_xpb_out[79][223],u_xpb_out[80][223],u_xpb_out[81][223],u_xpb_out[82][223],u_xpb_out[83][223],u_xpb_out[84][223],u_xpb_out[85][223],u_xpb_out[86][223],u_xpb_out[87][223],u_xpb_out[88][223],u_xpb_out[89][223],u_xpb_out[90][223],u_xpb_out[91][223],u_xpb_out[92][223],u_xpb_out[93][223],u_xpb_out[94][223],u_xpb_out[95][223],u_xpb_out[96][223],u_xpb_out[97][223],u_xpb_out[98][223],u_xpb_out[99][223],u_xpb_out[100][223],u_xpb_out[101][223],u_xpb_out[102][223],u_xpb_out[103][223],u_xpb_out[104][223],u_xpb_out[105][223]};

assign col_out_224 = {u_xpb_out[0][224],u_xpb_out[1][224],u_xpb_out[2][224],u_xpb_out[3][224],u_xpb_out[4][224],u_xpb_out[5][224],u_xpb_out[6][224],u_xpb_out[7][224],u_xpb_out[8][224],u_xpb_out[9][224],u_xpb_out[10][224],u_xpb_out[11][224],u_xpb_out[12][224],u_xpb_out[13][224],u_xpb_out[14][224],u_xpb_out[15][224],u_xpb_out[16][224],u_xpb_out[17][224],u_xpb_out[18][224],u_xpb_out[19][224],u_xpb_out[20][224],u_xpb_out[21][224],u_xpb_out[22][224],u_xpb_out[23][224],u_xpb_out[24][224],u_xpb_out[25][224],u_xpb_out[26][224],u_xpb_out[27][224],u_xpb_out[28][224],u_xpb_out[29][224],u_xpb_out[30][224],u_xpb_out[31][224],u_xpb_out[32][224],u_xpb_out[33][224],u_xpb_out[34][224],u_xpb_out[35][224],u_xpb_out[36][224],u_xpb_out[37][224],u_xpb_out[38][224],u_xpb_out[39][224],u_xpb_out[40][224],u_xpb_out[41][224],u_xpb_out[42][224],u_xpb_out[43][224],u_xpb_out[44][224],u_xpb_out[45][224],u_xpb_out[46][224],u_xpb_out[47][224],u_xpb_out[48][224],u_xpb_out[49][224],u_xpb_out[50][224],u_xpb_out[51][224],u_xpb_out[52][224],u_xpb_out[53][224],u_xpb_out[54][224],u_xpb_out[55][224],u_xpb_out[56][224],u_xpb_out[57][224],u_xpb_out[58][224],u_xpb_out[59][224],u_xpb_out[60][224],u_xpb_out[61][224],u_xpb_out[62][224],u_xpb_out[63][224],u_xpb_out[64][224],u_xpb_out[65][224],u_xpb_out[66][224],u_xpb_out[67][224],u_xpb_out[68][224],u_xpb_out[69][224],u_xpb_out[70][224],u_xpb_out[71][224],u_xpb_out[72][224],u_xpb_out[73][224],u_xpb_out[74][224],u_xpb_out[75][224],u_xpb_out[76][224],u_xpb_out[77][224],u_xpb_out[78][224],u_xpb_out[79][224],u_xpb_out[80][224],u_xpb_out[81][224],u_xpb_out[82][224],u_xpb_out[83][224],u_xpb_out[84][224],u_xpb_out[85][224],u_xpb_out[86][224],u_xpb_out[87][224],u_xpb_out[88][224],u_xpb_out[89][224],u_xpb_out[90][224],u_xpb_out[91][224],u_xpb_out[92][224],u_xpb_out[93][224],u_xpb_out[94][224],u_xpb_out[95][224],u_xpb_out[96][224],u_xpb_out[97][224],u_xpb_out[98][224],u_xpb_out[99][224],u_xpb_out[100][224],u_xpb_out[101][224],u_xpb_out[102][224],u_xpb_out[103][224],u_xpb_out[104][224],u_xpb_out[105][224]};

assign col_out_225 = {u_xpb_out[0][225],u_xpb_out[1][225],u_xpb_out[2][225],u_xpb_out[3][225],u_xpb_out[4][225],u_xpb_out[5][225],u_xpb_out[6][225],u_xpb_out[7][225],u_xpb_out[8][225],u_xpb_out[9][225],u_xpb_out[10][225],u_xpb_out[11][225],u_xpb_out[12][225],u_xpb_out[13][225],u_xpb_out[14][225],u_xpb_out[15][225],u_xpb_out[16][225],u_xpb_out[17][225],u_xpb_out[18][225],u_xpb_out[19][225],u_xpb_out[20][225],u_xpb_out[21][225],u_xpb_out[22][225],u_xpb_out[23][225],u_xpb_out[24][225],u_xpb_out[25][225],u_xpb_out[26][225],u_xpb_out[27][225],u_xpb_out[28][225],u_xpb_out[29][225],u_xpb_out[30][225],u_xpb_out[31][225],u_xpb_out[32][225],u_xpb_out[33][225],u_xpb_out[34][225],u_xpb_out[35][225],u_xpb_out[36][225],u_xpb_out[37][225],u_xpb_out[38][225],u_xpb_out[39][225],u_xpb_out[40][225],u_xpb_out[41][225],u_xpb_out[42][225],u_xpb_out[43][225],u_xpb_out[44][225],u_xpb_out[45][225],u_xpb_out[46][225],u_xpb_out[47][225],u_xpb_out[48][225],u_xpb_out[49][225],u_xpb_out[50][225],u_xpb_out[51][225],u_xpb_out[52][225],u_xpb_out[53][225],u_xpb_out[54][225],u_xpb_out[55][225],u_xpb_out[56][225],u_xpb_out[57][225],u_xpb_out[58][225],u_xpb_out[59][225],u_xpb_out[60][225],u_xpb_out[61][225],u_xpb_out[62][225],u_xpb_out[63][225],u_xpb_out[64][225],u_xpb_out[65][225],u_xpb_out[66][225],u_xpb_out[67][225],u_xpb_out[68][225],u_xpb_out[69][225],u_xpb_out[70][225],u_xpb_out[71][225],u_xpb_out[72][225],u_xpb_out[73][225],u_xpb_out[74][225],u_xpb_out[75][225],u_xpb_out[76][225],u_xpb_out[77][225],u_xpb_out[78][225],u_xpb_out[79][225],u_xpb_out[80][225],u_xpb_out[81][225],u_xpb_out[82][225],u_xpb_out[83][225],u_xpb_out[84][225],u_xpb_out[85][225],u_xpb_out[86][225],u_xpb_out[87][225],u_xpb_out[88][225],u_xpb_out[89][225],u_xpb_out[90][225],u_xpb_out[91][225],u_xpb_out[92][225],u_xpb_out[93][225],u_xpb_out[94][225],u_xpb_out[95][225],u_xpb_out[96][225],u_xpb_out[97][225],u_xpb_out[98][225],u_xpb_out[99][225],u_xpb_out[100][225],u_xpb_out[101][225],u_xpb_out[102][225],u_xpb_out[103][225],u_xpb_out[104][225],u_xpb_out[105][225]};

assign col_out_226 = {u_xpb_out[0][226],u_xpb_out[1][226],u_xpb_out[2][226],u_xpb_out[3][226],u_xpb_out[4][226],u_xpb_out[5][226],u_xpb_out[6][226],u_xpb_out[7][226],u_xpb_out[8][226],u_xpb_out[9][226],u_xpb_out[10][226],u_xpb_out[11][226],u_xpb_out[12][226],u_xpb_out[13][226],u_xpb_out[14][226],u_xpb_out[15][226],u_xpb_out[16][226],u_xpb_out[17][226],u_xpb_out[18][226],u_xpb_out[19][226],u_xpb_out[20][226],u_xpb_out[21][226],u_xpb_out[22][226],u_xpb_out[23][226],u_xpb_out[24][226],u_xpb_out[25][226],u_xpb_out[26][226],u_xpb_out[27][226],u_xpb_out[28][226],u_xpb_out[29][226],u_xpb_out[30][226],u_xpb_out[31][226],u_xpb_out[32][226],u_xpb_out[33][226],u_xpb_out[34][226],u_xpb_out[35][226],u_xpb_out[36][226],u_xpb_out[37][226],u_xpb_out[38][226],u_xpb_out[39][226],u_xpb_out[40][226],u_xpb_out[41][226],u_xpb_out[42][226],u_xpb_out[43][226],u_xpb_out[44][226],u_xpb_out[45][226],u_xpb_out[46][226],u_xpb_out[47][226],u_xpb_out[48][226],u_xpb_out[49][226],u_xpb_out[50][226],u_xpb_out[51][226],u_xpb_out[52][226],u_xpb_out[53][226],u_xpb_out[54][226],u_xpb_out[55][226],u_xpb_out[56][226],u_xpb_out[57][226],u_xpb_out[58][226],u_xpb_out[59][226],u_xpb_out[60][226],u_xpb_out[61][226],u_xpb_out[62][226],u_xpb_out[63][226],u_xpb_out[64][226],u_xpb_out[65][226],u_xpb_out[66][226],u_xpb_out[67][226],u_xpb_out[68][226],u_xpb_out[69][226],u_xpb_out[70][226],u_xpb_out[71][226],u_xpb_out[72][226],u_xpb_out[73][226],u_xpb_out[74][226],u_xpb_out[75][226],u_xpb_out[76][226],u_xpb_out[77][226],u_xpb_out[78][226],u_xpb_out[79][226],u_xpb_out[80][226],u_xpb_out[81][226],u_xpb_out[82][226],u_xpb_out[83][226],u_xpb_out[84][226],u_xpb_out[85][226],u_xpb_out[86][226],u_xpb_out[87][226],u_xpb_out[88][226],u_xpb_out[89][226],u_xpb_out[90][226],u_xpb_out[91][226],u_xpb_out[92][226],u_xpb_out[93][226],u_xpb_out[94][226],u_xpb_out[95][226],u_xpb_out[96][226],u_xpb_out[97][226],u_xpb_out[98][226],u_xpb_out[99][226],u_xpb_out[100][226],u_xpb_out[101][226],u_xpb_out[102][226],u_xpb_out[103][226],u_xpb_out[104][226],u_xpb_out[105][226]};

assign col_out_227 = {u_xpb_out[0][227],u_xpb_out[1][227],u_xpb_out[2][227],u_xpb_out[3][227],u_xpb_out[4][227],u_xpb_out[5][227],u_xpb_out[6][227],u_xpb_out[7][227],u_xpb_out[8][227],u_xpb_out[9][227],u_xpb_out[10][227],u_xpb_out[11][227],u_xpb_out[12][227],u_xpb_out[13][227],u_xpb_out[14][227],u_xpb_out[15][227],u_xpb_out[16][227],u_xpb_out[17][227],u_xpb_out[18][227],u_xpb_out[19][227],u_xpb_out[20][227],u_xpb_out[21][227],u_xpb_out[22][227],u_xpb_out[23][227],u_xpb_out[24][227],u_xpb_out[25][227],u_xpb_out[26][227],u_xpb_out[27][227],u_xpb_out[28][227],u_xpb_out[29][227],u_xpb_out[30][227],u_xpb_out[31][227],u_xpb_out[32][227],u_xpb_out[33][227],u_xpb_out[34][227],u_xpb_out[35][227],u_xpb_out[36][227],u_xpb_out[37][227],u_xpb_out[38][227],u_xpb_out[39][227],u_xpb_out[40][227],u_xpb_out[41][227],u_xpb_out[42][227],u_xpb_out[43][227],u_xpb_out[44][227],u_xpb_out[45][227],u_xpb_out[46][227],u_xpb_out[47][227],u_xpb_out[48][227],u_xpb_out[49][227],u_xpb_out[50][227],u_xpb_out[51][227],u_xpb_out[52][227],u_xpb_out[53][227],u_xpb_out[54][227],u_xpb_out[55][227],u_xpb_out[56][227],u_xpb_out[57][227],u_xpb_out[58][227],u_xpb_out[59][227],u_xpb_out[60][227],u_xpb_out[61][227],u_xpb_out[62][227],u_xpb_out[63][227],u_xpb_out[64][227],u_xpb_out[65][227],u_xpb_out[66][227],u_xpb_out[67][227],u_xpb_out[68][227],u_xpb_out[69][227],u_xpb_out[70][227],u_xpb_out[71][227],u_xpb_out[72][227],u_xpb_out[73][227],u_xpb_out[74][227],u_xpb_out[75][227],u_xpb_out[76][227],u_xpb_out[77][227],u_xpb_out[78][227],u_xpb_out[79][227],u_xpb_out[80][227],u_xpb_out[81][227],u_xpb_out[82][227],u_xpb_out[83][227],u_xpb_out[84][227],u_xpb_out[85][227],u_xpb_out[86][227],u_xpb_out[87][227],u_xpb_out[88][227],u_xpb_out[89][227],u_xpb_out[90][227],u_xpb_out[91][227],u_xpb_out[92][227],u_xpb_out[93][227],u_xpb_out[94][227],u_xpb_out[95][227],u_xpb_out[96][227],u_xpb_out[97][227],u_xpb_out[98][227],u_xpb_out[99][227],u_xpb_out[100][227],u_xpb_out[101][227],u_xpb_out[102][227],u_xpb_out[103][227],u_xpb_out[104][227],u_xpb_out[105][227]};

assign col_out_228 = {u_xpb_out[0][228],u_xpb_out[1][228],u_xpb_out[2][228],u_xpb_out[3][228],u_xpb_out[4][228],u_xpb_out[5][228],u_xpb_out[6][228],u_xpb_out[7][228],u_xpb_out[8][228],u_xpb_out[9][228],u_xpb_out[10][228],u_xpb_out[11][228],u_xpb_out[12][228],u_xpb_out[13][228],u_xpb_out[14][228],u_xpb_out[15][228],u_xpb_out[16][228],u_xpb_out[17][228],u_xpb_out[18][228],u_xpb_out[19][228],u_xpb_out[20][228],u_xpb_out[21][228],u_xpb_out[22][228],u_xpb_out[23][228],u_xpb_out[24][228],u_xpb_out[25][228],u_xpb_out[26][228],u_xpb_out[27][228],u_xpb_out[28][228],u_xpb_out[29][228],u_xpb_out[30][228],u_xpb_out[31][228],u_xpb_out[32][228],u_xpb_out[33][228],u_xpb_out[34][228],u_xpb_out[35][228],u_xpb_out[36][228],u_xpb_out[37][228],u_xpb_out[38][228],u_xpb_out[39][228],u_xpb_out[40][228],u_xpb_out[41][228],u_xpb_out[42][228],u_xpb_out[43][228],u_xpb_out[44][228],u_xpb_out[45][228],u_xpb_out[46][228],u_xpb_out[47][228],u_xpb_out[48][228],u_xpb_out[49][228],u_xpb_out[50][228],u_xpb_out[51][228],u_xpb_out[52][228],u_xpb_out[53][228],u_xpb_out[54][228],u_xpb_out[55][228],u_xpb_out[56][228],u_xpb_out[57][228],u_xpb_out[58][228],u_xpb_out[59][228],u_xpb_out[60][228],u_xpb_out[61][228],u_xpb_out[62][228],u_xpb_out[63][228],u_xpb_out[64][228],u_xpb_out[65][228],u_xpb_out[66][228],u_xpb_out[67][228],u_xpb_out[68][228],u_xpb_out[69][228],u_xpb_out[70][228],u_xpb_out[71][228],u_xpb_out[72][228],u_xpb_out[73][228],u_xpb_out[74][228],u_xpb_out[75][228],u_xpb_out[76][228],u_xpb_out[77][228],u_xpb_out[78][228],u_xpb_out[79][228],u_xpb_out[80][228],u_xpb_out[81][228],u_xpb_out[82][228],u_xpb_out[83][228],u_xpb_out[84][228],u_xpb_out[85][228],u_xpb_out[86][228],u_xpb_out[87][228],u_xpb_out[88][228],u_xpb_out[89][228],u_xpb_out[90][228],u_xpb_out[91][228],u_xpb_out[92][228],u_xpb_out[93][228],u_xpb_out[94][228],u_xpb_out[95][228],u_xpb_out[96][228],u_xpb_out[97][228],u_xpb_out[98][228],u_xpb_out[99][228],u_xpb_out[100][228],u_xpb_out[101][228],u_xpb_out[102][228],u_xpb_out[103][228],u_xpb_out[104][228],u_xpb_out[105][228]};

assign col_out_229 = {u_xpb_out[0][229],u_xpb_out[1][229],u_xpb_out[2][229],u_xpb_out[3][229],u_xpb_out[4][229],u_xpb_out[5][229],u_xpb_out[6][229],u_xpb_out[7][229],u_xpb_out[8][229],u_xpb_out[9][229],u_xpb_out[10][229],u_xpb_out[11][229],u_xpb_out[12][229],u_xpb_out[13][229],u_xpb_out[14][229],u_xpb_out[15][229],u_xpb_out[16][229],u_xpb_out[17][229],u_xpb_out[18][229],u_xpb_out[19][229],u_xpb_out[20][229],u_xpb_out[21][229],u_xpb_out[22][229],u_xpb_out[23][229],u_xpb_out[24][229],u_xpb_out[25][229],u_xpb_out[26][229],u_xpb_out[27][229],u_xpb_out[28][229],u_xpb_out[29][229],u_xpb_out[30][229],u_xpb_out[31][229],u_xpb_out[32][229],u_xpb_out[33][229],u_xpb_out[34][229],u_xpb_out[35][229],u_xpb_out[36][229],u_xpb_out[37][229],u_xpb_out[38][229],u_xpb_out[39][229],u_xpb_out[40][229],u_xpb_out[41][229],u_xpb_out[42][229],u_xpb_out[43][229],u_xpb_out[44][229],u_xpb_out[45][229],u_xpb_out[46][229],u_xpb_out[47][229],u_xpb_out[48][229],u_xpb_out[49][229],u_xpb_out[50][229],u_xpb_out[51][229],u_xpb_out[52][229],u_xpb_out[53][229],u_xpb_out[54][229],u_xpb_out[55][229],u_xpb_out[56][229],u_xpb_out[57][229],u_xpb_out[58][229],u_xpb_out[59][229],u_xpb_out[60][229],u_xpb_out[61][229],u_xpb_out[62][229],u_xpb_out[63][229],u_xpb_out[64][229],u_xpb_out[65][229],u_xpb_out[66][229],u_xpb_out[67][229],u_xpb_out[68][229],u_xpb_out[69][229],u_xpb_out[70][229],u_xpb_out[71][229],u_xpb_out[72][229],u_xpb_out[73][229],u_xpb_out[74][229],u_xpb_out[75][229],u_xpb_out[76][229],u_xpb_out[77][229],u_xpb_out[78][229],u_xpb_out[79][229],u_xpb_out[80][229],u_xpb_out[81][229],u_xpb_out[82][229],u_xpb_out[83][229],u_xpb_out[84][229],u_xpb_out[85][229],u_xpb_out[86][229],u_xpb_out[87][229],u_xpb_out[88][229],u_xpb_out[89][229],u_xpb_out[90][229],u_xpb_out[91][229],u_xpb_out[92][229],u_xpb_out[93][229],u_xpb_out[94][229],u_xpb_out[95][229],u_xpb_out[96][229],u_xpb_out[97][229],u_xpb_out[98][229],u_xpb_out[99][229],u_xpb_out[100][229],u_xpb_out[101][229],u_xpb_out[102][229],u_xpb_out[103][229],u_xpb_out[104][229],u_xpb_out[105][229]};

assign col_out_230 = {u_xpb_out[0][230],u_xpb_out[1][230],u_xpb_out[2][230],u_xpb_out[3][230],u_xpb_out[4][230],u_xpb_out[5][230],u_xpb_out[6][230],u_xpb_out[7][230],u_xpb_out[8][230],u_xpb_out[9][230],u_xpb_out[10][230],u_xpb_out[11][230],u_xpb_out[12][230],u_xpb_out[13][230],u_xpb_out[14][230],u_xpb_out[15][230],u_xpb_out[16][230],u_xpb_out[17][230],u_xpb_out[18][230],u_xpb_out[19][230],u_xpb_out[20][230],u_xpb_out[21][230],u_xpb_out[22][230],u_xpb_out[23][230],u_xpb_out[24][230],u_xpb_out[25][230],u_xpb_out[26][230],u_xpb_out[27][230],u_xpb_out[28][230],u_xpb_out[29][230],u_xpb_out[30][230],u_xpb_out[31][230],u_xpb_out[32][230],u_xpb_out[33][230],u_xpb_out[34][230],u_xpb_out[35][230],u_xpb_out[36][230],u_xpb_out[37][230],u_xpb_out[38][230],u_xpb_out[39][230],u_xpb_out[40][230],u_xpb_out[41][230],u_xpb_out[42][230],u_xpb_out[43][230],u_xpb_out[44][230],u_xpb_out[45][230],u_xpb_out[46][230],u_xpb_out[47][230],u_xpb_out[48][230],u_xpb_out[49][230],u_xpb_out[50][230],u_xpb_out[51][230],u_xpb_out[52][230],u_xpb_out[53][230],u_xpb_out[54][230],u_xpb_out[55][230],u_xpb_out[56][230],u_xpb_out[57][230],u_xpb_out[58][230],u_xpb_out[59][230],u_xpb_out[60][230],u_xpb_out[61][230],u_xpb_out[62][230],u_xpb_out[63][230],u_xpb_out[64][230],u_xpb_out[65][230],u_xpb_out[66][230],u_xpb_out[67][230],u_xpb_out[68][230],u_xpb_out[69][230],u_xpb_out[70][230],u_xpb_out[71][230],u_xpb_out[72][230],u_xpb_out[73][230],u_xpb_out[74][230],u_xpb_out[75][230],u_xpb_out[76][230],u_xpb_out[77][230],u_xpb_out[78][230],u_xpb_out[79][230],u_xpb_out[80][230],u_xpb_out[81][230],u_xpb_out[82][230],u_xpb_out[83][230],u_xpb_out[84][230],u_xpb_out[85][230],u_xpb_out[86][230],u_xpb_out[87][230],u_xpb_out[88][230],u_xpb_out[89][230],u_xpb_out[90][230],u_xpb_out[91][230],u_xpb_out[92][230],u_xpb_out[93][230],u_xpb_out[94][230],u_xpb_out[95][230],u_xpb_out[96][230],u_xpb_out[97][230],u_xpb_out[98][230],u_xpb_out[99][230],u_xpb_out[100][230],u_xpb_out[101][230],u_xpb_out[102][230],u_xpb_out[103][230],u_xpb_out[104][230],u_xpb_out[105][230]};

assign col_out_231 = {u_xpb_out[0][231],u_xpb_out[1][231],u_xpb_out[2][231],u_xpb_out[3][231],u_xpb_out[4][231],u_xpb_out[5][231],u_xpb_out[6][231],u_xpb_out[7][231],u_xpb_out[8][231],u_xpb_out[9][231],u_xpb_out[10][231],u_xpb_out[11][231],u_xpb_out[12][231],u_xpb_out[13][231],u_xpb_out[14][231],u_xpb_out[15][231],u_xpb_out[16][231],u_xpb_out[17][231],u_xpb_out[18][231],u_xpb_out[19][231],u_xpb_out[20][231],u_xpb_out[21][231],u_xpb_out[22][231],u_xpb_out[23][231],u_xpb_out[24][231],u_xpb_out[25][231],u_xpb_out[26][231],u_xpb_out[27][231],u_xpb_out[28][231],u_xpb_out[29][231],u_xpb_out[30][231],u_xpb_out[31][231],u_xpb_out[32][231],u_xpb_out[33][231],u_xpb_out[34][231],u_xpb_out[35][231],u_xpb_out[36][231],u_xpb_out[37][231],u_xpb_out[38][231],u_xpb_out[39][231],u_xpb_out[40][231],u_xpb_out[41][231],u_xpb_out[42][231],u_xpb_out[43][231],u_xpb_out[44][231],u_xpb_out[45][231],u_xpb_out[46][231],u_xpb_out[47][231],u_xpb_out[48][231],u_xpb_out[49][231],u_xpb_out[50][231],u_xpb_out[51][231],u_xpb_out[52][231],u_xpb_out[53][231],u_xpb_out[54][231],u_xpb_out[55][231],u_xpb_out[56][231],u_xpb_out[57][231],u_xpb_out[58][231],u_xpb_out[59][231],u_xpb_out[60][231],u_xpb_out[61][231],u_xpb_out[62][231],u_xpb_out[63][231],u_xpb_out[64][231],u_xpb_out[65][231],u_xpb_out[66][231],u_xpb_out[67][231],u_xpb_out[68][231],u_xpb_out[69][231],u_xpb_out[70][231],u_xpb_out[71][231],u_xpb_out[72][231],u_xpb_out[73][231],u_xpb_out[74][231],u_xpb_out[75][231],u_xpb_out[76][231],u_xpb_out[77][231],u_xpb_out[78][231],u_xpb_out[79][231],u_xpb_out[80][231],u_xpb_out[81][231],u_xpb_out[82][231],u_xpb_out[83][231],u_xpb_out[84][231],u_xpb_out[85][231],u_xpb_out[86][231],u_xpb_out[87][231],u_xpb_out[88][231],u_xpb_out[89][231],u_xpb_out[90][231],u_xpb_out[91][231],u_xpb_out[92][231],u_xpb_out[93][231],u_xpb_out[94][231],u_xpb_out[95][231],u_xpb_out[96][231],u_xpb_out[97][231],u_xpb_out[98][231],u_xpb_out[99][231],u_xpb_out[100][231],u_xpb_out[101][231],u_xpb_out[102][231],u_xpb_out[103][231],u_xpb_out[104][231],u_xpb_out[105][231]};

assign col_out_232 = {u_xpb_out[0][232],u_xpb_out[1][232],u_xpb_out[2][232],u_xpb_out[3][232],u_xpb_out[4][232],u_xpb_out[5][232],u_xpb_out[6][232],u_xpb_out[7][232],u_xpb_out[8][232],u_xpb_out[9][232],u_xpb_out[10][232],u_xpb_out[11][232],u_xpb_out[12][232],u_xpb_out[13][232],u_xpb_out[14][232],u_xpb_out[15][232],u_xpb_out[16][232],u_xpb_out[17][232],u_xpb_out[18][232],u_xpb_out[19][232],u_xpb_out[20][232],u_xpb_out[21][232],u_xpb_out[22][232],u_xpb_out[23][232],u_xpb_out[24][232],u_xpb_out[25][232],u_xpb_out[26][232],u_xpb_out[27][232],u_xpb_out[28][232],u_xpb_out[29][232],u_xpb_out[30][232],u_xpb_out[31][232],u_xpb_out[32][232],u_xpb_out[33][232],u_xpb_out[34][232],u_xpb_out[35][232],u_xpb_out[36][232],u_xpb_out[37][232],u_xpb_out[38][232],u_xpb_out[39][232],u_xpb_out[40][232],u_xpb_out[41][232],u_xpb_out[42][232],u_xpb_out[43][232],u_xpb_out[44][232],u_xpb_out[45][232],u_xpb_out[46][232],u_xpb_out[47][232],u_xpb_out[48][232],u_xpb_out[49][232],u_xpb_out[50][232],u_xpb_out[51][232],u_xpb_out[52][232],u_xpb_out[53][232],u_xpb_out[54][232],u_xpb_out[55][232],u_xpb_out[56][232],u_xpb_out[57][232],u_xpb_out[58][232],u_xpb_out[59][232],u_xpb_out[60][232],u_xpb_out[61][232],u_xpb_out[62][232],u_xpb_out[63][232],u_xpb_out[64][232],u_xpb_out[65][232],u_xpb_out[66][232],u_xpb_out[67][232],u_xpb_out[68][232],u_xpb_out[69][232],u_xpb_out[70][232],u_xpb_out[71][232],u_xpb_out[72][232],u_xpb_out[73][232],u_xpb_out[74][232],u_xpb_out[75][232],u_xpb_out[76][232],u_xpb_out[77][232],u_xpb_out[78][232],u_xpb_out[79][232],u_xpb_out[80][232],u_xpb_out[81][232],u_xpb_out[82][232],u_xpb_out[83][232],u_xpb_out[84][232],u_xpb_out[85][232],u_xpb_out[86][232],u_xpb_out[87][232],u_xpb_out[88][232],u_xpb_out[89][232],u_xpb_out[90][232],u_xpb_out[91][232],u_xpb_out[92][232],u_xpb_out[93][232],u_xpb_out[94][232],u_xpb_out[95][232],u_xpb_out[96][232],u_xpb_out[97][232],u_xpb_out[98][232],u_xpb_out[99][232],u_xpb_out[100][232],u_xpb_out[101][232],u_xpb_out[102][232],u_xpb_out[103][232],u_xpb_out[104][232],u_xpb_out[105][232]};

assign col_out_233 = {u_xpb_out[0][233],u_xpb_out[1][233],u_xpb_out[2][233],u_xpb_out[3][233],u_xpb_out[4][233],u_xpb_out[5][233],u_xpb_out[6][233],u_xpb_out[7][233],u_xpb_out[8][233],u_xpb_out[9][233],u_xpb_out[10][233],u_xpb_out[11][233],u_xpb_out[12][233],u_xpb_out[13][233],u_xpb_out[14][233],u_xpb_out[15][233],u_xpb_out[16][233],u_xpb_out[17][233],u_xpb_out[18][233],u_xpb_out[19][233],u_xpb_out[20][233],u_xpb_out[21][233],u_xpb_out[22][233],u_xpb_out[23][233],u_xpb_out[24][233],u_xpb_out[25][233],u_xpb_out[26][233],u_xpb_out[27][233],u_xpb_out[28][233],u_xpb_out[29][233],u_xpb_out[30][233],u_xpb_out[31][233],u_xpb_out[32][233],u_xpb_out[33][233],u_xpb_out[34][233],u_xpb_out[35][233],u_xpb_out[36][233],u_xpb_out[37][233],u_xpb_out[38][233],u_xpb_out[39][233],u_xpb_out[40][233],u_xpb_out[41][233],u_xpb_out[42][233],u_xpb_out[43][233],u_xpb_out[44][233],u_xpb_out[45][233],u_xpb_out[46][233],u_xpb_out[47][233],u_xpb_out[48][233],u_xpb_out[49][233],u_xpb_out[50][233],u_xpb_out[51][233],u_xpb_out[52][233],u_xpb_out[53][233],u_xpb_out[54][233],u_xpb_out[55][233],u_xpb_out[56][233],u_xpb_out[57][233],u_xpb_out[58][233],u_xpb_out[59][233],u_xpb_out[60][233],u_xpb_out[61][233],u_xpb_out[62][233],u_xpb_out[63][233],u_xpb_out[64][233],u_xpb_out[65][233],u_xpb_out[66][233],u_xpb_out[67][233],u_xpb_out[68][233],u_xpb_out[69][233],u_xpb_out[70][233],u_xpb_out[71][233],u_xpb_out[72][233],u_xpb_out[73][233],u_xpb_out[74][233],u_xpb_out[75][233],u_xpb_out[76][233],u_xpb_out[77][233],u_xpb_out[78][233],u_xpb_out[79][233],u_xpb_out[80][233],u_xpb_out[81][233],u_xpb_out[82][233],u_xpb_out[83][233],u_xpb_out[84][233],u_xpb_out[85][233],u_xpb_out[86][233],u_xpb_out[87][233],u_xpb_out[88][233],u_xpb_out[89][233],u_xpb_out[90][233],u_xpb_out[91][233],u_xpb_out[92][233],u_xpb_out[93][233],u_xpb_out[94][233],u_xpb_out[95][233],u_xpb_out[96][233],u_xpb_out[97][233],u_xpb_out[98][233],u_xpb_out[99][233],u_xpb_out[100][233],u_xpb_out[101][233],u_xpb_out[102][233],u_xpb_out[103][233],u_xpb_out[104][233],u_xpb_out[105][233]};

assign col_out_234 = {u_xpb_out[0][234],u_xpb_out[1][234],u_xpb_out[2][234],u_xpb_out[3][234],u_xpb_out[4][234],u_xpb_out[5][234],u_xpb_out[6][234],u_xpb_out[7][234],u_xpb_out[8][234],u_xpb_out[9][234],u_xpb_out[10][234],u_xpb_out[11][234],u_xpb_out[12][234],u_xpb_out[13][234],u_xpb_out[14][234],u_xpb_out[15][234],u_xpb_out[16][234],u_xpb_out[17][234],u_xpb_out[18][234],u_xpb_out[19][234],u_xpb_out[20][234],u_xpb_out[21][234],u_xpb_out[22][234],u_xpb_out[23][234],u_xpb_out[24][234],u_xpb_out[25][234],u_xpb_out[26][234],u_xpb_out[27][234],u_xpb_out[28][234],u_xpb_out[29][234],u_xpb_out[30][234],u_xpb_out[31][234],u_xpb_out[32][234],u_xpb_out[33][234],u_xpb_out[34][234],u_xpb_out[35][234],u_xpb_out[36][234],u_xpb_out[37][234],u_xpb_out[38][234],u_xpb_out[39][234],u_xpb_out[40][234],u_xpb_out[41][234],u_xpb_out[42][234],u_xpb_out[43][234],u_xpb_out[44][234],u_xpb_out[45][234],u_xpb_out[46][234],u_xpb_out[47][234],u_xpb_out[48][234],u_xpb_out[49][234],u_xpb_out[50][234],u_xpb_out[51][234],u_xpb_out[52][234],u_xpb_out[53][234],u_xpb_out[54][234],u_xpb_out[55][234],u_xpb_out[56][234],u_xpb_out[57][234],u_xpb_out[58][234],u_xpb_out[59][234],u_xpb_out[60][234],u_xpb_out[61][234],u_xpb_out[62][234],u_xpb_out[63][234],u_xpb_out[64][234],u_xpb_out[65][234],u_xpb_out[66][234],u_xpb_out[67][234],u_xpb_out[68][234],u_xpb_out[69][234],u_xpb_out[70][234],u_xpb_out[71][234],u_xpb_out[72][234],u_xpb_out[73][234],u_xpb_out[74][234],u_xpb_out[75][234],u_xpb_out[76][234],u_xpb_out[77][234],u_xpb_out[78][234],u_xpb_out[79][234],u_xpb_out[80][234],u_xpb_out[81][234],u_xpb_out[82][234],u_xpb_out[83][234],u_xpb_out[84][234],u_xpb_out[85][234],u_xpb_out[86][234],u_xpb_out[87][234],u_xpb_out[88][234],u_xpb_out[89][234],u_xpb_out[90][234],u_xpb_out[91][234],u_xpb_out[92][234],u_xpb_out[93][234],u_xpb_out[94][234],u_xpb_out[95][234],u_xpb_out[96][234],u_xpb_out[97][234],u_xpb_out[98][234],u_xpb_out[99][234],u_xpb_out[100][234],u_xpb_out[101][234],u_xpb_out[102][234],u_xpb_out[103][234],u_xpb_out[104][234],u_xpb_out[105][234]};

assign col_out_235 = {u_xpb_out[0][235],u_xpb_out[1][235],u_xpb_out[2][235],u_xpb_out[3][235],u_xpb_out[4][235],u_xpb_out[5][235],u_xpb_out[6][235],u_xpb_out[7][235],u_xpb_out[8][235],u_xpb_out[9][235],u_xpb_out[10][235],u_xpb_out[11][235],u_xpb_out[12][235],u_xpb_out[13][235],u_xpb_out[14][235],u_xpb_out[15][235],u_xpb_out[16][235],u_xpb_out[17][235],u_xpb_out[18][235],u_xpb_out[19][235],u_xpb_out[20][235],u_xpb_out[21][235],u_xpb_out[22][235],u_xpb_out[23][235],u_xpb_out[24][235],u_xpb_out[25][235],u_xpb_out[26][235],u_xpb_out[27][235],u_xpb_out[28][235],u_xpb_out[29][235],u_xpb_out[30][235],u_xpb_out[31][235],u_xpb_out[32][235],u_xpb_out[33][235],u_xpb_out[34][235],u_xpb_out[35][235],u_xpb_out[36][235],u_xpb_out[37][235],u_xpb_out[38][235],u_xpb_out[39][235],u_xpb_out[40][235],u_xpb_out[41][235],u_xpb_out[42][235],u_xpb_out[43][235],u_xpb_out[44][235],u_xpb_out[45][235],u_xpb_out[46][235],u_xpb_out[47][235],u_xpb_out[48][235],u_xpb_out[49][235],u_xpb_out[50][235],u_xpb_out[51][235],u_xpb_out[52][235],u_xpb_out[53][235],u_xpb_out[54][235],u_xpb_out[55][235],u_xpb_out[56][235],u_xpb_out[57][235],u_xpb_out[58][235],u_xpb_out[59][235],u_xpb_out[60][235],u_xpb_out[61][235],u_xpb_out[62][235],u_xpb_out[63][235],u_xpb_out[64][235],u_xpb_out[65][235],u_xpb_out[66][235],u_xpb_out[67][235],u_xpb_out[68][235],u_xpb_out[69][235],u_xpb_out[70][235],u_xpb_out[71][235],u_xpb_out[72][235],u_xpb_out[73][235],u_xpb_out[74][235],u_xpb_out[75][235],u_xpb_out[76][235],u_xpb_out[77][235],u_xpb_out[78][235],u_xpb_out[79][235],u_xpb_out[80][235],u_xpb_out[81][235],u_xpb_out[82][235],u_xpb_out[83][235],u_xpb_out[84][235],u_xpb_out[85][235],u_xpb_out[86][235],u_xpb_out[87][235],u_xpb_out[88][235],u_xpb_out[89][235],u_xpb_out[90][235],u_xpb_out[91][235],u_xpb_out[92][235],u_xpb_out[93][235],u_xpb_out[94][235],u_xpb_out[95][235],u_xpb_out[96][235],u_xpb_out[97][235],u_xpb_out[98][235],u_xpb_out[99][235],u_xpb_out[100][235],u_xpb_out[101][235],u_xpb_out[102][235],u_xpb_out[103][235],u_xpb_out[104][235],u_xpb_out[105][235]};

assign col_out_236 = {u_xpb_out[0][236],u_xpb_out[1][236],u_xpb_out[2][236],u_xpb_out[3][236],u_xpb_out[4][236],u_xpb_out[5][236],u_xpb_out[6][236],u_xpb_out[7][236],u_xpb_out[8][236],u_xpb_out[9][236],u_xpb_out[10][236],u_xpb_out[11][236],u_xpb_out[12][236],u_xpb_out[13][236],u_xpb_out[14][236],u_xpb_out[15][236],u_xpb_out[16][236],u_xpb_out[17][236],u_xpb_out[18][236],u_xpb_out[19][236],u_xpb_out[20][236],u_xpb_out[21][236],u_xpb_out[22][236],u_xpb_out[23][236],u_xpb_out[24][236],u_xpb_out[25][236],u_xpb_out[26][236],u_xpb_out[27][236],u_xpb_out[28][236],u_xpb_out[29][236],u_xpb_out[30][236],u_xpb_out[31][236],u_xpb_out[32][236],u_xpb_out[33][236],u_xpb_out[34][236],u_xpb_out[35][236],u_xpb_out[36][236],u_xpb_out[37][236],u_xpb_out[38][236],u_xpb_out[39][236],u_xpb_out[40][236],u_xpb_out[41][236],u_xpb_out[42][236],u_xpb_out[43][236],u_xpb_out[44][236],u_xpb_out[45][236],u_xpb_out[46][236],u_xpb_out[47][236],u_xpb_out[48][236],u_xpb_out[49][236],u_xpb_out[50][236],u_xpb_out[51][236],u_xpb_out[52][236],u_xpb_out[53][236],u_xpb_out[54][236],u_xpb_out[55][236],u_xpb_out[56][236],u_xpb_out[57][236],u_xpb_out[58][236],u_xpb_out[59][236],u_xpb_out[60][236],u_xpb_out[61][236],u_xpb_out[62][236],u_xpb_out[63][236],u_xpb_out[64][236],u_xpb_out[65][236],u_xpb_out[66][236],u_xpb_out[67][236],u_xpb_out[68][236],u_xpb_out[69][236],u_xpb_out[70][236],u_xpb_out[71][236],u_xpb_out[72][236],u_xpb_out[73][236],u_xpb_out[74][236],u_xpb_out[75][236],u_xpb_out[76][236],u_xpb_out[77][236],u_xpb_out[78][236],u_xpb_out[79][236],u_xpb_out[80][236],u_xpb_out[81][236],u_xpb_out[82][236],u_xpb_out[83][236],u_xpb_out[84][236],u_xpb_out[85][236],u_xpb_out[86][236],u_xpb_out[87][236],u_xpb_out[88][236],u_xpb_out[89][236],u_xpb_out[90][236],u_xpb_out[91][236],u_xpb_out[92][236],u_xpb_out[93][236],u_xpb_out[94][236],u_xpb_out[95][236],u_xpb_out[96][236],u_xpb_out[97][236],u_xpb_out[98][236],u_xpb_out[99][236],u_xpb_out[100][236],u_xpb_out[101][236],u_xpb_out[102][236],u_xpb_out[103][236],u_xpb_out[104][236],u_xpb_out[105][236]};

assign col_out_237 = {u_xpb_out[0][237],u_xpb_out[1][237],u_xpb_out[2][237],u_xpb_out[3][237],u_xpb_out[4][237],u_xpb_out[5][237],u_xpb_out[6][237],u_xpb_out[7][237],u_xpb_out[8][237],u_xpb_out[9][237],u_xpb_out[10][237],u_xpb_out[11][237],u_xpb_out[12][237],u_xpb_out[13][237],u_xpb_out[14][237],u_xpb_out[15][237],u_xpb_out[16][237],u_xpb_out[17][237],u_xpb_out[18][237],u_xpb_out[19][237],u_xpb_out[20][237],u_xpb_out[21][237],u_xpb_out[22][237],u_xpb_out[23][237],u_xpb_out[24][237],u_xpb_out[25][237],u_xpb_out[26][237],u_xpb_out[27][237],u_xpb_out[28][237],u_xpb_out[29][237],u_xpb_out[30][237],u_xpb_out[31][237],u_xpb_out[32][237],u_xpb_out[33][237],u_xpb_out[34][237],u_xpb_out[35][237],u_xpb_out[36][237],u_xpb_out[37][237],u_xpb_out[38][237],u_xpb_out[39][237],u_xpb_out[40][237],u_xpb_out[41][237],u_xpb_out[42][237],u_xpb_out[43][237],u_xpb_out[44][237],u_xpb_out[45][237],u_xpb_out[46][237],u_xpb_out[47][237],u_xpb_out[48][237],u_xpb_out[49][237],u_xpb_out[50][237],u_xpb_out[51][237],u_xpb_out[52][237],u_xpb_out[53][237],u_xpb_out[54][237],u_xpb_out[55][237],u_xpb_out[56][237],u_xpb_out[57][237],u_xpb_out[58][237],u_xpb_out[59][237],u_xpb_out[60][237],u_xpb_out[61][237],u_xpb_out[62][237],u_xpb_out[63][237],u_xpb_out[64][237],u_xpb_out[65][237],u_xpb_out[66][237],u_xpb_out[67][237],u_xpb_out[68][237],u_xpb_out[69][237],u_xpb_out[70][237],u_xpb_out[71][237],u_xpb_out[72][237],u_xpb_out[73][237],u_xpb_out[74][237],u_xpb_out[75][237],u_xpb_out[76][237],u_xpb_out[77][237],u_xpb_out[78][237],u_xpb_out[79][237],u_xpb_out[80][237],u_xpb_out[81][237],u_xpb_out[82][237],u_xpb_out[83][237],u_xpb_out[84][237],u_xpb_out[85][237],u_xpb_out[86][237],u_xpb_out[87][237],u_xpb_out[88][237],u_xpb_out[89][237],u_xpb_out[90][237],u_xpb_out[91][237],u_xpb_out[92][237],u_xpb_out[93][237],u_xpb_out[94][237],u_xpb_out[95][237],u_xpb_out[96][237],u_xpb_out[97][237],u_xpb_out[98][237],u_xpb_out[99][237],u_xpb_out[100][237],u_xpb_out[101][237],u_xpb_out[102][237],u_xpb_out[103][237],u_xpb_out[104][237],u_xpb_out[105][237]};

assign col_out_238 = {u_xpb_out[0][238],u_xpb_out[1][238],u_xpb_out[2][238],u_xpb_out[3][238],u_xpb_out[4][238],u_xpb_out[5][238],u_xpb_out[6][238],u_xpb_out[7][238],u_xpb_out[8][238],u_xpb_out[9][238],u_xpb_out[10][238],u_xpb_out[11][238],u_xpb_out[12][238],u_xpb_out[13][238],u_xpb_out[14][238],u_xpb_out[15][238],u_xpb_out[16][238],u_xpb_out[17][238],u_xpb_out[18][238],u_xpb_out[19][238],u_xpb_out[20][238],u_xpb_out[21][238],u_xpb_out[22][238],u_xpb_out[23][238],u_xpb_out[24][238],u_xpb_out[25][238],u_xpb_out[26][238],u_xpb_out[27][238],u_xpb_out[28][238],u_xpb_out[29][238],u_xpb_out[30][238],u_xpb_out[31][238],u_xpb_out[32][238],u_xpb_out[33][238],u_xpb_out[34][238],u_xpb_out[35][238],u_xpb_out[36][238],u_xpb_out[37][238],u_xpb_out[38][238],u_xpb_out[39][238],u_xpb_out[40][238],u_xpb_out[41][238],u_xpb_out[42][238],u_xpb_out[43][238],u_xpb_out[44][238],u_xpb_out[45][238],u_xpb_out[46][238],u_xpb_out[47][238],u_xpb_out[48][238],u_xpb_out[49][238],u_xpb_out[50][238],u_xpb_out[51][238],u_xpb_out[52][238],u_xpb_out[53][238],u_xpb_out[54][238],u_xpb_out[55][238],u_xpb_out[56][238],u_xpb_out[57][238],u_xpb_out[58][238],u_xpb_out[59][238],u_xpb_out[60][238],u_xpb_out[61][238],u_xpb_out[62][238],u_xpb_out[63][238],u_xpb_out[64][238],u_xpb_out[65][238],u_xpb_out[66][238],u_xpb_out[67][238],u_xpb_out[68][238],u_xpb_out[69][238],u_xpb_out[70][238],u_xpb_out[71][238],u_xpb_out[72][238],u_xpb_out[73][238],u_xpb_out[74][238],u_xpb_out[75][238],u_xpb_out[76][238],u_xpb_out[77][238],u_xpb_out[78][238],u_xpb_out[79][238],u_xpb_out[80][238],u_xpb_out[81][238],u_xpb_out[82][238],u_xpb_out[83][238],u_xpb_out[84][238],u_xpb_out[85][238],u_xpb_out[86][238],u_xpb_out[87][238],u_xpb_out[88][238],u_xpb_out[89][238],u_xpb_out[90][238],u_xpb_out[91][238],u_xpb_out[92][238],u_xpb_out[93][238],u_xpb_out[94][238],u_xpb_out[95][238],u_xpb_out[96][238],u_xpb_out[97][238],u_xpb_out[98][238],u_xpb_out[99][238],u_xpb_out[100][238],u_xpb_out[101][238],u_xpb_out[102][238],u_xpb_out[103][238],u_xpb_out[104][238],u_xpb_out[105][238]};

assign col_out_239 = {u_xpb_out[0][239],u_xpb_out[1][239],u_xpb_out[2][239],u_xpb_out[3][239],u_xpb_out[4][239],u_xpb_out[5][239],u_xpb_out[6][239],u_xpb_out[7][239],u_xpb_out[8][239],u_xpb_out[9][239],u_xpb_out[10][239],u_xpb_out[11][239],u_xpb_out[12][239],u_xpb_out[13][239],u_xpb_out[14][239],u_xpb_out[15][239],u_xpb_out[16][239],u_xpb_out[17][239],u_xpb_out[18][239],u_xpb_out[19][239],u_xpb_out[20][239],u_xpb_out[21][239],u_xpb_out[22][239],u_xpb_out[23][239],u_xpb_out[24][239],u_xpb_out[25][239],u_xpb_out[26][239],u_xpb_out[27][239],u_xpb_out[28][239],u_xpb_out[29][239],u_xpb_out[30][239],u_xpb_out[31][239],u_xpb_out[32][239],u_xpb_out[33][239],u_xpb_out[34][239],u_xpb_out[35][239],u_xpb_out[36][239],u_xpb_out[37][239],u_xpb_out[38][239],u_xpb_out[39][239],u_xpb_out[40][239],u_xpb_out[41][239],u_xpb_out[42][239],u_xpb_out[43][239],u_xpb_out[44][239],u_xpb_out[45][239],u_xpb_out[46][239],u_xpb_out[47][239],u_xpb_out[48][239],u_xpb_out[49][239],u_xpb_out[50][239],u_xpb_out[51][239],u_xpb_out[52][239],u_xpb_out[53][239],u_xpb_out[54][239],u_xpb_out[55][239],u_xpb_out[56][239],u_xpb_out[57][239],u_xpb_out[58][239],u_xpb_out[59][239],u_xpb_out[60][239],u_xpb_out[61][239],u_xpb_out[62][239],u_xpb_out[63][239],u_xpb_out[64][239],u_xpb_out[65][239],u_xpb_out[66][239],u_xpb_out[67][239],u_xpb_out[68][239],u_xpb_out[69][239],u_xpb_out[70][239],u_xpb_out[71][239],u_xpb_out[72][239],u_xpb_out[73][239],u_xpb_out[74][239],u_xpb_out[75][239],u_xpb_out[76][239],u_xpb_out[77][239],u_xpb_out[78][239],u_xpb_out[79][239],u_xpb_out[80][239],u_xpb_out[81][239],u_xpb_out[82][239],u_xpb_out[83][239],u_xpb_out[84][239],u_xpb_out[85][239],u_xpb_out[86][239],u_xpb_out[87][239],u_xpb_out[88][239],u_xpb_out[89][239],u_xpb_out[90][239],u_xpb_out[91][239],u_xpb_out[92][239],u_xpb_out[93][239],u_xpb_out[94][239],u_xpb_out[95][239],u_xpb_out[96][239],u_xpb_out[97][239],u_xpb_out[98][239],u_xpb_out[99][239],u_xpb_out[100][239],u_xpb_out[101][239],u_xpb_out[102][239],u_xpb_out[103][239],u_xpb_out[104][239],u_xpb_out[105][239]};

assign col_out_240 = {u_xpb_out[0][240],u_xpb_out[1][240],u_xpb_out[2][240],u_xpb_out[3][240],u_xpb_out[4][240],u_xpb_out[5][240],u_xpb_out[6][240],u_xpb_out[7][240],u_xpb_out[8][240],u_xpb_out[9][240],u_xpb_out[10][240],u_xpb_out[11][240],u_xpb_out[12][240],u_xpb_out[13][240],u_xpb_out[14][240],u_xpb_out[15][240],u_xpb_out[16][240],u_xpb_out[17][240],u_xpb_out[18][240],u_xpb_out[19][240],u_xpb_out[20][240],u_xpb_out[21][240],u_xpb_out[22][240],u_xpb_out[23][240],u_xpb_out[24][240],u_xpb_out[25][240],u_xpb_out[26][240],u_xpb_out[27][240],u_xpb_out[28][240],u_xpb_out[29][240],u_xpb_out[30][240],u_xpb_out[31][240],u_xpb_out[32][240],u_xpb_out[33][240],u_xpb_out[34][240],u_xpb_out[35][240],u_xpb_out[36][240],u_xpb_out[37][240],u_xpb_out[38][240],u_xpb_out[39][240],u_xpb_out[40][240],u_xpb_out[41][240],u_xpb_out[42][240],u_xpb_out[43][240],u_xpb_out[44][240],u_xpb_out[45][240],u_xpb_out[46][240],u_xpb_out[47][240],u_xpb_out[48][240],u_xpb_out[49][240],u_xpb_out[50][240],u_xpb_out[51][240],u_xpb_out[52][240],u_xpb_out[53][240],u_xpb_out[54][240],u_xpb_out[55][240],u_xpb_out[56][240],u_xpb_out[57][240],u_xpb_out[58][240],u_xpb_out[59][240],u_xpb_out[60][240],u_xpb_out[61][240],u_xpb_out[62][240],u_xpb_out[63][240],u_xpb_out[64][240],u_xpb_out[65][240],u_xpb_out[66][240],u_xpb_out[67][240],u_xpb_out[68][240],u_xpb_out[69][240],u_xpb_out[70][240],u_xpb_out[71][240],u_xpb_out[72][240],u_xpb_out[73][240],u_xpb_out[74][240],u_xpb_out[75][240],u_xpb_out[76][240],u_xpb_out[77][240],u_xpb_out[78][240],u_xpb_out[79][240],u_xpb_out[80][240],u_xpb_out[81][240],u_xpb_out[82][240],u_xpb_out[83][240],u_xpb_out[84][240],u_xpb_out[85][240],u_xpb_out[86][240],u_xpb_out[87][240],u_xpb_out[88][240],u_xpb_out[89][240],u_xpb_out[90][240],u_xpb_out[91][240],u_xpb_out[92][240],u_xpb_out[93][240],u_xpb_out[94][240],u_xpb_out[95][240],u_xpb_out[96][240],u_xpb_out[97][240],u_xpb_out[98][240],u_xpb_out[99][240],u_xpb_out[100][240],u_xpb_out[101][240],u_xpb_out[102][240],u_xpb_out[103][240],u_xpb_out[104][240],u_xpb_out[105][240]};

assign col_out_241 = {u_xpb_out[0][241],u_xpb_out[1][241],u_xpb_out[2][241],u_xpb_out[3][241],u_xpb_out[4][241],u_xpb_out[5][241],u_xpb_out[6][241],u_xpb_out[7][241],u_xpb_out[8][241],u_xpb_out[9][241],u_xpb_out[10][241],u_xpb_out[11][241],u_xpb_out[12][241],u_xpb_out[13][241],u_xpb_out[14][241],u_xpb_out[15][241],u_xpb_out[16][241],u_xpb_out[17][241],u_xpb_out[18][241],u_xpb_out[19][241],u_xpb_out[20][241],u_xpb_out[21][241],u_xpb_out[22][241],u_xpb_out[23][241],u_xpb_out[24][241],u_xpb_out[25][241],u_xpb_out[26][241],u_xpb_out[27][241],u_xpb_out[28][241],u_xpb_out[29][241],u_xpb_out[30][241],u_xpb_out[31][241],u_xpb_out[32][241],u_xpb_out[33][241],u_xpb_out[34][241],u_xpb_out[35][241],u_xpb_out[36][241],u_xpb_out[37][241],u_xpb_out[38][241],u_xpb_out[39][241],u_xpb_out[40][241],u_xpb_out[41][241],u_xpb_out[42][241],u_xpb_out[43][241],u_xpb_out[44][241],u_xpb_out[45][241],u_xpb_out[46][241],u_xpb_out[47][241],u_xpb_out[48][241],u_xpb_out[49][241],u_xpb_out[50][241],u_xpb_out[51][241],u_xpb_out[52][241],u_xpb_out[53][241],u_xpb_out[54][241],u_xpb_out[55][241],u_xpb_out[56][241],u_xpb_out[57][241],u_xpb_out[58][241],u_xpb_out[59][241],u_xpb_out[60][241],u_xpb_out[61][241],u_xpb_out[62][241],u_xpb_out[63][241],u_xpb_out[64][241],u_xpb_out[65][241],u_xpb_out[66][241],u_xpb_out[67][241],u_xpb_out[68][241],u_xpb_out[69][241],u_xpb_out[70][241],u_xpb_out[71][241],u_xpb_out[72][241],u_xpb_out[73][241],u_xpb_out[74][241],u_xpb_out[75][241],u_xpb_out[76][241],u_xpb_out[77][241],u_xpb_out[78][241],u_xpb_out[79][241],u_xpb_out[80][241],u_xpb_out[81][241],u_xpb_out[82][241],u_xpb_out[83][241],u_xpb_out[84][241],u_xpb_out[85][241],u_xpb_out[86][241],u_xpb_out[87][241],u_xpb_out[88][241],u_xpb_out[89][241],u_xpb_out[90][241],u_xpb_out[91][241],u_xpb_out[92][241],u_xpb_out[93][241],u_xpb_out[94][241],u_xpb_out[95][241],u_xpb_out[96][241],u_xpb_out[97][241],u_xpb_out[98][241],u_xpb_out[99][241],u_xpb_out[100][241],u_xpb_out[101][241],u_xpb_out[102][241],u_xpb_out[103][241],u_xpb_out[104][241],u_xpb_out[105][241]};

assign col_out_242 = {u_xpb_out[0][242],u_xpb_out[1][242],u_xpb_out[2][242],u_xpb_out[3][242],u_xpb_out[4][242],u_xpb_out[5][242],u_xpb_out[6][242],u_xpb_out[7][242],u_xpb_out[8][242],u_xpb_out[9][242],u_xpb_out[10][242],u_xpb_out[11][242],u_xpb_out[12][242],u_xpb_out[13][242],u_xpb_out[14][242],u_xpb_out[15][242],u_xpb_out[16][242],u_xpb_out[17][242],u_xpb_out[18][242],u_xpb_out[19][242],u_xpb_out[20][242],u_xpb_out[21][242],u_xpb_out[22][242],u_xpb_out[23][242],u_xpb_out[24][242],u_xpb_out[25][242],u_xpb_out[26][242],u_xpb_out[27][242],u_xpb_out[28][242],u_xpb_out[29][242],u_xpb_out[30][242],u_xpb_out[31][242],u_xpb_out[32][242],u_xpb_out[33][242],u_xpb_out[34][242],u_xpb_out[35][242],u_xpb_out[36][242],u_xpb_out[37][242],u_xpb_out[38][242],u_xpb_out[39][242],u_xpb_out[40][242],u_xpb_out[41][242],u_xpb_out[42][242],u_xpb_out[43][242],u_xpb_out[44][242],u_xpb_out[45][242],u_xpb_out[46][242],u_xpb_out[47][242],u_xpb_out[48][242],u_xpb_out[49][242],u_xpb_out[50][242],u_xpb_out[51][242],u_xpb_out[52][242],u_xpb_out[53][242],u_xpb_out[54][242],u_xpb_out[55][242],u_xpb_out[56][242],u_xpb_out[57][242],u_xpb_out[58][242],u_xpb_out[59][242],u_xpb_out[60][242],u_xpb_out[61][242],u_xpb_out[62][242],u_xpb_out[63][242],u_xpb_out[64][242],u_xpb_out[65][242],u_xpb_out[66][242],u_xpb_out[67][242],u_xpb_out[68][242],u_xpb_out[69][242],u_xpb_out[70][242],u_xpb_out[71][242],u_xpb_out[72][242],u_xpb_out[73][242],u_xpb_out[74][242],u_xpb_out[75][242],u_xpb_out[76][242],u_xpb_out[77][242],u_xpb_out[78][242],u_xpb_out[79][242],u_xpb_out[80][242],u_xpb_out[81][242],u_xpb_out[82][242],u_xpb_out[83][242],u_xpb_out[84][242],u_xpb_out[85][242],u_xpb_out[86][242],u_xpb_out[87][242],u_xpb_out[88][242],u_xpb_out[89][242],u_xpb_out[90][242],u_xpb_out[91][242],u_xpb_out[92][242],u_xpb_out[93][242],u_xpb_out[94][242],u_xpb_out[95][242],u_xpb_out[96][242],u_xpb_out[97][242],u_xpb_out[98][242],u_xpb_out[99][242],u_xpb_out[100][242],u_xpb_out[101][242],u_xpb_out[102][242],u_xpb_out[103][242],u_xpb_out[104][242],u_xpb_out[105][242]};

assign col_out_243 = {u_xpb_out[0][243],u_xpb_out[1][243],u_xpb_out[2][243],u_xpb_out[3][243],u_xpb_out[4][243],u_xpb_out[5][243],u_xpb_out[6][243],u_xpb_out[7][243],u_xpb_out[8][243],u_xpb_out[9][243],u_xpb_out[10][243],u_xpb_out[11][243],u_xpb_out[12][243],u_xpb_out[13][243],u_xpb_out[14][243],u_xpb_out[15][243],u_xpb_out[16][243],u_xpb_out[17][243],u_xpb_out[18][243],u_xpb_out[19][243],u_xpb_out[20][243],u_xpb_out[21][243],u_xpb_out[22][243],u_xpb_out[23][243],u_xpb_out[24][243],u_xpb_out[25][243],u_xpb_out[26][243],u_xpb_out[27][243],u_xpb_out[28][243],u_xpb_out[29][243],u_xpb_out[30][243],u_xpb_out[31][243],u_xpb_out[32][243],u_xpb_out[33][243],u_xpb_out[34][243],u_xpb_out[35][243],u_xpb_out[36][243],u_xpb_out[37][243],u_xpb_out[38][243],u_xpb_out[39][243],u_xpb_out[40][243],u_xpb_out[41][243],u_xpb_out[42][243],u_xpb_out[43][243],u_xpb_out[44][243],u_xpb_out[45][243],u_xpb_out[46][243],u_xpb_out[47][243],u_xpb_out[48][243],u_xpb_out[49][243],u_xpb_out[50][243],u_xpb_out[51][243],u_xpb_out[52][243],u_xpb_out[53][243],u_xpb_out[54][243],u_xpb_out[55][243],u_xpb_out[56][243],u_xpb_out[57][243],u_xpb_out[58][243],u_xpb_out[59][243],u_xpb_out[60][243],u_xpb_out[61][243],u_xpb_out[62][243],u_xpb_out[63][243],u_xpb_out[64][243],u_xpb_out[65][243],u_xpb_out[66][243],u_xpb_out[67][243],u_xpb_out[68][243],u_xpb_out[69][243],u_xpb_out[70][243],u_xpb_out[71][243],u_xpb_out[72][243],u_xpb_out[73][243],u_xpb_out[74][243],u_xpb_out[75][243],u_xpb_out[76][243],u_xpb_out[77][243],u_xpb_out[78][243],u_xpb_out[79][243],u_xpb_out[80][243],u_xpb_out[81][243],u_xpb_out[82][243],u_xpb_out[83][243],u_xpb_out[84][243],u_xpb_out[85][243],u_xpb_out[86][243],u_xpb_out[87][243],u_xpb_out[88][243],u_xpb_out[89][243],u_xpb_out[90][243],u_xpb_out[91][243],u_xpb_out[92][243],u_xpb_out[93][243],u_xpb_out[94][243],u_xpb_out[95][243],u_xpb_out[96][243],u_xpb_out[97][243],u_xpb_out[98][243],u_xpb_out[99][243],u_xpb_out[100][243],u_xpb_out[101][243],u_xpb_out[102][243],u_xpb_out[103][243],u_xpb_out[104][243],u_xpb_out[105][243]};

assign col_out_244 = {u_xpb_out[0][244],u_xpb_out[1][244],u_xpb_out[2][244],u_xpb_out[3][244],u_xpb_out[4][244],u_xpb_out[5][244],u_xpb_out[6][244],u_xpb_out[7][244],u_xpb_out[8][244],u_xpb_out[9][244],u_xpb_out[10][244],u_xpb_out[11][244],u_xpb_out[12][244],u_xpb_out[13][244],u_xpb_out[14][244],u_xpb_out[15][244],u_xpb_out[16][244],u_xpb_out[17][244],u_xpb_out[18][244],u_xpb_out[19][244],u_xpb_out[20][244],u_xpb_out[21][244],u_xpb_out[22][244],u_xpb_out[23][244],u_xpb_out[24][244],u_xpb_out[25][244],u_xpb_out[26][244],u_xpb_out[27][244],u_xpb_out[28][244],u_xpb_out[29][244],u_xpb_out[30][244],u_xpb_out[31][244],u_xpb_out[32][244],u_xpb_out[33][244],u_xpb_out[34][244],u_xpb_out[35][244],u_xpb_out[36][244],u_xpb_out[37][244],u_xpb_out[38][244],u_xpb_out[39][244],u_xpb_out[40][244],u_xpb_out[41][244],u_xpb_out[42][244],u_xpb_out[43][244],u_xpb_out[44][244],u_xpb_out[45][244],u_xpb_out[46][244],u_xpb_out[47][244],u_xpb_out[48][244],u_xpb_out[49][244],u_xpb_out[50][244],u_xpb_out[51][244],u_xpb_out[52][244],u_xpb_out[53][244],u_xpb_out[54][244],u_xpb_out[55][244],u_xpb_out[56][244],u_xpb_out[57][244],u_xpb_out[58][244],u_xpb_out[59][244],u_xpb_out[60][244],u_xpb_out[61][244],u_xpb_out[62][244],u_xpb_out[63][244],u_xpb_out[64][244],u_xpb_out[65][244],u_xpb_out[66][244],u_xpb_out[67][244],u_xpb_out[68][244],u_xpb_out[69][244],u_xpb_out[70][244],u_xpb_out[71][244],u_xpb_out[72][244],u_xpb_out[73][244],u_xpb_out[74][244],u_xpb_out[75][244],u_xpb_out[76][244],u_xpb_out[77][244],u_xpb_out[78][244],u_xpb_out[79][244],u_xpb_out[80][244],u_xpb_out[81][244],u_xpb_out[82][244],u_xpb_out[83][244],u_xpb_out[84][244],u_xpb_out[85][244],u_xpb_out[86][244],u_xpb_out[87][244],u_xpb_out[88][244],u_xpb_out[89][244],u_xpb_out[90][244],u_xpb_out[91][244],u_xpb_out[92][244],u_xpb_out[93][244],u_xpb_out[94][244],u_xpb_out[95][244],u_xpb_out[96][244],u_xpb_out[97][244],u_xpb_out[98][244],u_xpb_out[99][244],u_xpb_out[100][244],u_xpb_out[101][244],u_xpb_out[102][244],u_xpb_out[103][244],u_xpb_out[104][244],u_xpb_out[105][244]};

assign col_out_245 = {u_xpb_out[0][245],u_xpb_out[1][245],u_xpb_out[2][245],u_xpb_out[3][245],u_xpb_out[4][245],u_xpb_out[5][245],u_xpb_out[6][245],u_xpb_out[7][245],u_xpb_out[8][245],u_xpb_out[9][245],u_xpb_out[10][245],u_xpb_out[11][245],u_xpb_out[12][245],u_xpb_out[13][245],u_xpb_out[14][245],u_xpb_out[15][245],u_xpb_out[16][245],u_xpb_out[17][245],u_xpb_out[18][245],u_xpb_out[19][245],u_xpb_out[20][245],u_xpb_out[21][245],u_xpb_out[22][245],u_xpb_out[23][245],u_xpb_out[24][245],u_xpb_out[25][245],u_xpb_out[26][245],u_xpb_out[27][245],u_xpb_out[28][245],u_xpb_out[29][245],u_xpb_out[30][245],u_xpb_out[31][245],u_xpb_out[32][245],u_xpb_out[33][245],u_xpb_out[34][245],u_xpb_out[35][245],u_xpb_out[36][245],u_xpb_out[37][245],u_xpb_out[38][245],u_xpb_out[39][245],u_xpb_out[40][245],u_xpb_out[41][245],u_xpb_out[42][245],u_xpb_out[43][245],u_xpb_out[44][245],u_xpb_out[45][245],u_xpb_out[46][245],u_xpb_out[47][245],u_xpb_out[48][245],u_xpb_out[49][245],u_xpb_out[50][245],u_xpb_out[51][245],u_xpb_out[52][245],u_xpb_out[53][245],u_xpb_out[54][245],u_xpb_out[55][245],u_xpb_out[56][245],u_xpb_out[57][245],u_xpb_out[58][245],u_xpb_out[59][245],u_xpb_out[60][245],u_xpb_out[61][245],u_xpb_out[62][245],u_xpb_out[63][245],u_xpb_out[64][245],u_xpb_out[65][245],u_xpb_out[66][245],u_xpb_out[67][245],u_xpb_out[68][245],u_xpb_out[69][245],u_xpb_out[70][245],u_xpb_out[71][245],u_xpb_out[72][245],u_xpb_out[73][245],u_xpb_out[74][245],u_xpb_out[75][245],u_xpb_out[76][245],u_xpb_out[77][245],u_xpb_out[78][245],u_xpb_out[79][245],u_xpb_out[80][245],u_xpb_out[81][245],u_xpb_out[82][245],u_xpb_out[83][245],u_xpb_out[84][245],u_xpb_out[85][245],u_xpb_out[86][245],u_xpb_out[87][245],u_xpb_out[88][245],u_xpb_out[89][245],u_xpb_out[90][245],u_xpb_out[91][245],u_xpb_out[92][245],u_xpb_out[93][245],u_xpb_out[94][245],u_xpb_out[95][245],u_xpb_out[96][245],u_xpb_out[97][245],u_xpb_out[98][245],u_xpb_out[99][245],u_xpb_out[100][245],u_xpb_out[101][245],u_xpb_out[102][245],u_xpb_out[103][245],u_xpb_out[104][245],u_xpb_out[105][245]};

assign col_out_246 = {u_xpb_out[0][246],u_xpb_out[1][246],u_xpb_out[2][246],u_xpb_out[3][246],u_xpb_out[4][246],u_xpb_out[5][246],u_xpb_out[6][246],u_xpb_out[7][246],u_xpb_out[8][246],u_xpb_out[9][246],u_xpb_out[10][246],u_xpb_out[11][246],u_xpb_out[12][246],u_xpb_out[13][246],u_xpb_out[14][246],u_xpb_out[15][246],u_xpb_out[16][246],u_xpb_out[17][246],u_xpb_out[18][246],u_xpb_out[19][246],u_xpb_out[20][246],u_xpb_out[21][246],u_xpb_out[22][246],u_xpb_out[23][246],u_xpb_out[24][246],u_xpb_out[25][246],u_xpb_out[26][246],u_xpb_out[27][246],u_xpb_out[28][246],u_xpb_out[29][246],u_xpb_out[30][246],u_xpb_out[31][246],u_xpb_out[32][246],u_xpb_out[33][246],u_xpb_out[34][246],u_xpb_out[35][246],u_xpb_out[36][246],u_xpb_out[37][246],u_xpb_out[38][246],u_xpb_out[39][246],u_xpb_out[40][246],u_xpb_out[41][246],u_xpb_out[42][246],u_xpb_out[43][246],u_xpb_out[44][246],u_xpb_out[45][246],u_xpb_out[46][246],u_xpb_out[47][246],u_xpb_out[48][246],u_xpb_out[49][246],u_xpb_out[50][246],u_xpb_out[51][246],u_xpb_out[52][246],u_xpb_out[53][246],u_xpb_out[54][246],u_xpb_out[55][246],u_xpb_out[56][246],u_xpb_out[57][246],u_xpb_out[58][246],u_xpb_out[59][246],u_xpb_out[60][246],u_xpb_out[61][246],u_xpb_out[62][246],u_xpb_out[63][246],u_xpb_out[64][246],u_xpb_out[65][246],u_xpb_out[66][246],u_xpb_out[67][246],u_xpb_out[68][246],u_xpb_out[69][246],u_xpb_out[70][246],u_xpb_out[71][246],u_xpb_out[72][246],u_xpb_out[73][246],u_xpb_out[74][246],u_xpb_out[75][246],u_xpb_out[76][246],u_xpb_out[77][246],u_xpb_out[78][246],u_xpb_out[79][246],u_xpb_out[80][246],u_xpb_out[81][246],u_xpb_out[82][246],u_xpb_out[83][246],u_xpb_out[84][246],u_xpb_out[85][246],u_xpb_out[86][246],u_xpb_out[87][246],u_xpb_out[88][246],u_xpb_out[89][246],u_xpb_out[90][246],u_xpb_out[91][246],u_xpb_out[92][246],u_xpb_out[93][246],u_xpb_out[94][246],u_xpb_out[95][246],u_xpb_out[96][246],u_xpb_out[97][246],u_xpb_out[98][246],u_xpb_out[99][246],u_xpb_out[100][246],u_xpb_out[101][246],u_xpb_out[102][246],u_xpb_out[103][246],u_xpb_out[104][246],u_xpb_out[105][246]};

assign col_out_247 = {u_xpb_out[0][247],u_xpb_out[1][247],u_xpb_out[2][247],u_xpb_out[3][247],u_xpb_out[4][247],u_xpb_out[5][247],u_xpb_out[6][247],u_xpb_out[7][247],u_xpb_out[8][247],u_xpb_out[9][247],u_xpb_out[10][247],u_xpb_out[11][247],u_xpb_out[12][247],u_xpb_out[13][247],u_xpb_out[14][247],u_xpb_out[15][247],u_xpb_out[16][247],u_xpb_out[17][247],u_xpb_out[18][247],u_xpb_out[19][247],u_xpb_out[20][247],u_xpb_out[21][247],u_xpb_out[22][247],u_xpb_out[23][247],u_xpb_out[24][247],u_xpb_out[25][247],u_xpb_out[26][247],u_xpb_out[27][247],u_xpb_out[28][247],u_xpb_out[29][247],u_xpb_out[30][247],u_xpb_out[31][247],u_xpb_out[32][247],u_xpb_out[33][247],u_xpb_out[34][247],u_xpb_out[35][247],u_xpb_out[36][247],u_xpb_out[37][247],u_xpb_out[38][247],u_xpb_out[39][247],u_xpb_out[40][247],u_xpb_out[41][247],u_xpb_out[42][247],u_xpb_out[43][247],u_xpb_out[44][247],u_xpb_out[45][247],u_xpb_out[46][247],u_xpb_out[47][247],u_xpb_out[48][247],u_xpb_out[49][247],u_xpb_out[50][247],u_xpb_out[51][247],u_xpb_out[52][247],u_xpb_out[53][247],u_xpb_out[54][247],u_xpb_out[55][247],u_xpb_out[56][247],u_xpb_out[57][247],u_xpb_out[58][247],u_xpb_out[59][247],u_xpb_out[60][247],u_xpb_out[61][247],u_xpb_out[62][247],u_xpb_out[63][247],u_xpb_out[64][247],u_xpb_out[65][247],u_xpb_out[66][247],u_xpb_out[67][247],u_xpb_out[68][247],u_xpb_out[69][247],u_xpb_out[70][247],u_xpb_out[71][247],u_xpb_out[72][247],u_xpb_out[73][247],u_xpb_out[74][247],u_xpb_out[75][247],u_xpb_out[76][247],u_xpb_out[77][247],u_xpb_out[78][247],u_xpb_out[79][247],u_xpb_out[80][247],u_xpb_out[81][247],u_xpb_out[82][247],u_xpb_out[83][247],u_xpb_out[84][247],u_xpb_out[85][247],u_xpb_out[86][247],u_xpb_out[87][247],u_xpb_out[88][247],u_xpb_out[89][247],u_xpb_out[90][247],u_xpb_out[91][247],u_xpb_out[92][247],u_xpb_out[93][247],u_xpb_out[94][247],u_xpb_out[95][247],u_xpb_out[96][247],u_xpb_out[97][247],u_xpb_out[98][247],u_xpb_out[99][247],u_xpb_out[100][247],u_xpb_out[101][247],u_xpb_out[102][247],u_xpb_out[103][247],u_xpb_out[104][247],u_xpb_out[105][247]};

assign col_out_248 = {u_xpb_out[0][248],u_xpb_out[1][248],u_xpb_out[2][248],u_xpb_out[3][248],u_xpb_out[4][248],u_xpb_out[5][248],u_xpb_out[6][248],u_xpb_out[7][248],u_xpb_out[8][248],u_xpb_out[9][248],u_xpb_out[10][248],u_xpb_out[11][248],u_xpb_out[12][248],u_xpb_out[13][248],u_xpb_out[14][248],u_xpb_out[15][248],u_xpb_out[16][248],u_xpb_out[17][248],u_xpb_out[18][248],u_xpb_out[19][248],u_xpb_out[20][248],u_xpb_out[21][248],u_xpb_out[22][248],u_xpb_out[23][248],u_xpb_out[24][248],u_xpb_out[25][248],u_xpb_out[26][248],u_xpb_out[27][248],u_xpb_out[28][248],u_xpb_out[29][248],u_xpb_out[30][248],u_xpb_out[31][248],u_xpb_out[32][248],u_xpb_out[33][248],u_xpb_out[34][248],u_xpb_out[35][248],u_xpb_out[36][248],u_xpb_out[37][248],u_xpb_out[38][248],u_xpb_out[39][248],u_xpb_out[40][248],u_xpb_out[41][248],u_xpb_out[42][248],u_xpb_out[43][248],u_xpb_out[44][248],u_xpb_out[45][248],u_xpb_out[46][248],u_xpb_out[47][248],u_xpb_out[48][248],u_xpb_out[49][248],u_xpb_out[50][248],u_xpb_out[51][248],u_xpb_out[52][248],u_xpb_out[53][248],u_xpb_out[54][248],u_xpb_out[55][248],u_xpb_out[56][248],u_xpb_out[57][248],u_xpb_out[58][248],u_xpb_out[59][248],u_xpb_out[60][248],u_xpb_out[61][248],u_xpb_out[62][248],u_xpb_out[63][248],u_xpb_out[64][248],u_xpb_out[65][248],u_xpb_out[66][248],u_xpb_out[67][248],u_xpb_out[68][248],u_xpb_out[69][248],u_xpb_out[70][248],u_xpb_out[71][248],u_xpb_out[72][248],u_xpb_out[73][248],u_xpb_out[74][248],u_xpb_out[75][248],u_xpb_out[76][248],u_xpb_out[77][248],u_xpb_out[78][248],u_xpb_out[79][248],u_xpb_out[80][248],u_xpb_out[81][248],u_xpb_out[82][248],u_xpb_out[83][248],u_xpb_out[84][248],u_xpb_out[85][248],u_xpb_out[86][248],u_xpb_out[87][248],u_xpb_out[88][248],u_xpb_out[89][248],u_xpb_out[90][248],u_xpb_out[91][248],u_xpb_out[92][248],u_xpb_out[93][248],u_xpb_out[94][248],u_xpb_out[95][248],u_xpb_out[96][248],u_xpb_out[97][248],u_xpb_out[98][248],u_xpb_out[99][248],u_xpb_out[100][248],u_xpb_out[101][248],u_xpb_out[102][248],u_xpb_out[103][248],u_xpb_out[104][248],u_xpb_out[105][248]};

assign col_out_249 = {u_xpb_out[0][249],u_xpb_out[1][249],u_xpb_out[2][249],u_xpb_out[3][249],u_xpb_out[4][249],u_xpb_out[5][249],u_xpb_out[6][249],u_xpb_out[7][249],u_xpb_out[8][249],u_xpb_out[9][249],u_xpb_out[10][249],u_xpb_out[11][249],u_xpb_out[12][249],u_xpb_out[13][249],u_xpb_out[14][249],u_xpb_out[15][249],u_xpb_out[16][249],u_xpb_out[17][249],u_xpb_out[18][249],u_xpb_out[19][249],u_xpb_out[20][249],u_xpb_out[21][249],u_xpb_out[22][249],u_xpb_out[23][249],u_xpb_out[24][249],u_xpb_out[25][249],u_xpb_out[26][249],u_xpb_out[27][249],u_xpb_out[28][249],u_xpb_out[29][249],u_xpb_out[30][249],u_xpb_out[31][249],u_xpb_out[32][249],u_xpb_out[33][249],u_xpb_out[34][249],u_xpb_out[35][249],u_xpb_out[36][249],u_xpb_out[37][249],u_xpb_out[38][249],u_xpb_out[39][249],u_xpb_out[40][249],u_xpb_out[41][249],u_xpb_out[42][249],u_xpb_out[43][249],u_xpb_out[44][249],u_xpb_out[45][249],u_xpb_out[46][249],u_xpb_out[47][249],u_xpb_out[48][249],u_xpb_out[49][249],u_xpb_out[50][249],u_xpb_out[51][249],u_xpb_out[52][249],u_xpb_out[53][249],u_xpb_out[54][249],u_xpb_out[55][249],u_xpb_out[56][249],u_xpb_out[57][249],u_xpb_out[58][249],u_xpb_out[59][249],u_xpb_out[60][249],u_xpb_out[61][249],u_xpb_out[62][249],u_xpb_out[63][249],u_xpb_out[64][249],u_xpb_out[65][249],u_xpb_out[66][249],u_xpb_out[67][249],u_xpb_out[68][249],u_xpb_out[69][249],u_xpb_out[70][249],u_xpb_out[71][249],u_xpb_out[72][249],u_xpb_out[73][249],u_xpb_out[74][249],u_xpb_out[75][249],u_xpb_out[76][249],u_xpb_out[77][249],u_xpb_out[78][249],u_xpb_out[79][249],u_xpb_out[80][249],u_xpb_out[81][249],u_xpb_out[82][249],u_xpb_out[83][249],u_xpb_out[84][249],u_xpb_out[85][249],u_xpb_out[86][249],u_xpb_out[87][249],u_xpb_out[88][249],u_xpb_out[89][249],u_xpb_out[90][249],u_xpb_out[91][249],u_xpb_out[92][249],u_xpb_out[93][249],u_xpb_out[94][249],u_xpb_out[95][249],u_xpb_out[96][249],u_xpb_out[97][249],u_xpb_out[98][249],u_xpb_out[99][249],u_xpb_out[100][249],u_xpb_out[101][249],u_xpb_out[102][249],u_xpb_out[103][249],u_xpb_out[104][249],u_xpb_out[105][249]};

assign col_out_250 = {u_xpb_out[0][250],u_xpb_out[1][250],u_xpb_out[2][250],u_xpb_out[3][250],u_xpb_out[4][250],u_xpb_out[5][250],u_xpb_out[6][250],u_xpb_out[7][250],u_xpb_out[8][250],u_xpb_out[9][250],u_xpb_out[10][250],u_xpb_out[11][250],u_xpb_out[12][250],u_xpb_out[13][250],u_xpb_out[14][250],u_xpb_out[15][250],u_xpb_out[16][250],u_xpb_out[17][250],u_xpb_out[18][250],u_xpb_out[19][250],u_xpb_out[20][250],u_xpb_out[21][250],u_xpb_out[22][250],u_xpb_out[23][250],u_xpb_out[24][250],u_xpb_out[25][250],u_xpb_out[26][250],u_xpb_out[27][250],u_xpb_out[28][250],u_xpb_out[29][250],u_xpb_out[30][250],u_xpb_out[31][250],u_xpb_out[32][250],u_xpb_out[33][250],u_xpb_out[34][250],u_xpb_out[35][250],u_xpb_out[36][250],u_xpb_out[37][250],u_xpb_out[38][250],u_xpb_out[39][250],u_xpb_out[40][250],u_xpb_out[41][250],u_xpb_out[42][250],u_xpb_out[43][250],u_xpb_out[44][250],u_xpb_out[45][250],u_xpb_out[46][250],u_xpb_out[47][250],u_xpb_out[48][250],u_xpb_out[49][250],u_xpb_out[50][250],u_xpb_out[51][250],u_xpb_out[52][250],u_xpb_out[53][250],u_xpb_out[54][250],u_xpb_out[55][250],u_xpb_out[56][250],u_xpb_out[57][250],u_xpb_out[58][250],u_xpb_out[59][250],u_xpb_out[60][250],u_xpb_out[61][250],u_xpb_out[62][250],u_xpb_out[63][250],u_xpb_out[64][250],u_xpb_out[65][250],u_xpb_out[66][250],u_xpb_out[67][250],u_xpb_out[68][250],u_xpb_out[69][250],u_xpb_out[70][250],u_xpb_out[71][250],u_xpb_out[72][250],u_xpb_out[73][250],u_xpb_out[74][250],u_xpb_out[75][250],u_xpb_out[76][250],u_xpb_out[77][250],u_xpb_out[78][250],u_xpb_out[79][250],u_xpb_out[80][250],u_xpb_out[81][250],u_xpb_out[82][250],u_xpb_out[83][250],u_xpb_out[84][250],u_xpb_out[85][250],u_xpb_out[86][250],u_xpb_out[87][250],u_xpb_out[88][250],u_xpb_out[89][250],u_xpb_out[90][250],u_xpb_out[91][250],u_xpb_out[92][250],u_xpb_out[93][250],u_xpb_out[94][250],u_xpb_out[95][250],u_xpb_out[96][250],u_xpb_out[97][250],u_xpb_out[98][250],u_xpb_out[99][250],u_xpb_out[100][250],u_xpb_out[101][250],u_xpb_out[102][250],u_xpb_out[103][250],u_xpb_out[104][250],u_xpb_out[105][250]};

assign col_out_251 = {u_xpb_out[0][251],u_xpb_out[1][251],u_xpb_out[2][251],u_xpb_out[3][251],u_xpb_out[4][251],u_xpb_out[5][251],u_xpb_out[6][251],u_xpb_out[7][251],u_xpb_out[8][251],u_xpb_out[9][251],u_xpb_out[10][251],u_xpb_out[11][251],u_xpb_out[12][251],u_xpb_out[13][251],u_xpb_out[14][251],u_xpb_out[15][251],u_xpb_out[16][251],u_xpb_out[17][251],u_xpb_out[18][251],u_xpb_out[19][251],u_xpb_out[20][251],u_xpb_out[21][251],u_xpb_out[22][251],u_xpb_out[23][251],u_xpb_out[24][251],u_xpb_out[25][251],u_xpb_out[26][251],u_xpb_out[27][251],u_xpb_out[28][251],u_xpb_out[29][251],u_xpb_out[30][251],u_xpb_out[31][251],u_xpb_out[32][251],u_xpb_out[33][251],u_xpb_out[34][251],u_xpb_out[35][251],u_xpb_out[36][251],u_xpb_out[37][251],u_xpb_out[38][251],u_xpb_out[39][251],u_xpb_out[40][251],u_xpb_out[41][251],u_xpb_out[42][251],u_xpb_out[43][251],u_xpb_out[44][251],u_xpb_out[45][251],u_xpb_out[46][251],u_xpb_out[47][251],u_xpb_out[48][251],u_xpb_out[49][251],u_xpb_out[50][251],u_xpb_out[51][251],u_xpb_out[52][251],u_xpb_out[53][251],u_xpb_out[54][251],u_xpb_out[55][251],u_xpb_out[56][251],u_xpb_out[57][251],u_xpb_out[58][251],u_xpb_out[59][251],u_xpb_out[60][251],u_xpb_out[61][251],u_xpb_out[62][251],u_xpb_out[63][251],u_xpb_out[64][251],u_xpb_out[65][251],u_xpb_out[66][251],u_xpb_out[67][251],u_xpb_out[68][251],u_xpb_out[69][251],u_xpb_out[70][251],u_xpb_out[71][251],u_xpb_out[72][251],u_xpb_out[73][251],u_xpb_out[74][251],u_xpb_out[75][251],u_xpb_out[76][251],u_xpb_out[77][251],u_xpb_out[78][251],u_xpb_out[79][251],u_xpb_out[80][251],u_xpb_out[81][251],u_xpb_out[82][251],u_xpb_out[83][251],u_xpb_out[84][251],u_xpb_out[85][251],u_xpb_out[86][251],u_xpb_out[87][251],u_xpb_out[88][251],u_xpb_out[89][251],u_xpb_out[90][251],u_xpb_out[91][251],u_xpb_out[92][251],u_xpb_out[93][251],u_xpb_out[94][251],u_xpb_out[95][251],u_xpb_out[96][251],u_xpb_out[97][251],u_xpb_out[98][251],u_xpb_out[99][251],u_xpb_out[100][251],u_xpb_out[101][251],u_xpb_out[102][251],u_xpb_out[103][251],u_xpb_out[104][251],u_xpb_out[105][251]};

assign col_out_252 = {u_xpb_out[0][252],u_xpb_out[1][252],u_xpb_out[2][252],u_xpb_out[3][252],u_xpb_out[4][252],u_xpb_out[5][252],u_xpb_out[6][252],u_xpb_out[7][252],u_xpb_out[8][252],u_xpb_out[9][252],u_xpb_out[10][252],u_xpb_out[11][252],u_xpb_out[12][252],u_xpb_out[13][252],u_xpb_out[14][252],u_xpb_out[15][252],u_xpb_out[16][252],u_xpb_out[17][252],u_xpb_out[18][252],u_xpb_out[19][252],u_xpb_out[20][252],u_xpb_out[21][252],u_xpb_out[22][252],u_xpb_out[23][252],u_xpb_out[24][252],u_xpb_out[25][252],u_xpb_out[26][252],u_xpb_out[27][252],u_xpb_out[28][252],u_xpb_out[29][252],u_xpb_out[30][252],u_xpb_out[31][252],u_xpb_out[32][252],u_xpb_out[33][252],u_xpb_out[34][252],u_xpb_out[35][252],u_xpb_out[36][252],u_xpb_out[37][252],u_xpb_out[38][252],u_xpb_out[39][252],u_xpb_out[40][252],u_xpb_out[41][252],u_xpb_out[42][252],u_xpb_out[43][252],u_xpb_out[44][252],u_xpb_out[45][252],u_xpb_out[46][252],u_xpb_out[47][252],u_xpb_out[48][252],u_xpb_out[49][252],u_xpb_out[50][252],u_xpb_out[51][252],u_xpb_out[52][252],u_xpb_out[53][252],u_xpb_out[54][252],u_xpb_out[55][252],u_xpb_out[56][252],u_xpb_out[57][252],u_xpb_out[58][252],u_xpb_out[59][252],u_xpb_out[60][252],u_xpb_out[61][252],u_xpb_out[62][252],u_xpb_out[63][252],u_xpb_out[64][252],u_xpb_out[65][252],u_xpb_out[66][252],u_xpb_out[67][252],u_xpb_out[68][252],u_xpb_out[69][252],u_xpb_out[70][252],u_xpb_out[71][252],u_xpb_out[72][252],u_xpb_out[73][252],u_xpb_out[74][252],u_xpb_out[75][252],u_xpb_out[76][252],u_xpb_out[77][252],u_xpb_out[78][252],u_xpb_out[79][252],u_xpb_out[80][252],u_xpb_out[81][252],u_xpb_out[82][252],u_xpb_out[83][252],u_xpb_out[84][252],u_xpb_out[85][252],u_xpb_out[86][252],u_xpb_out[87][252],u_xpb_out[88][252],u_xpb_out[89][252],u_xpb_out[90][252],u_xpb_out[91][252],u_xpb_out[92][252],u_xpb_out[93][252],u_xpb_out[94][252],u_xpb_out[95][252],u_xpb_out[96][252],u_xpb_out[97][252],u_xpb_out[98][252],u_xpb_out[99][252],u_xpb_out[100][252],u_xpb_out[101][252],u_xpb_out[102][252],u_xpb_out[103][252],u_xpb_out[104][252],u_xpb_out[105][252]};

assign col_out_253 = {u_xpb_out[0][253],u_xpb_out[1][253],u_xpb_out[2][253],u_xpb_out[3][253],u_xpb_out[4][253],u_xpb_out[5][253],u_xpb_out[6][253],u_xpb_out[7][253],u_xpb_out[8][253],u_xpb_out[9][253],u_xpb_out[10][253],u_xpb_out[11][253],u_xpb_out[12][253],u_xpb_out[13][253],u_xpb_out[14][253],u_xpb_out[15][253],u_xpb_out[16][253],u_xpb_out[17][253],u_xpb_out[18][253],u_xpb_out[19][253],u_xpb_out[20][253],u_xpb_out[21][253],u_xpb_out[22][253],u_xpb_out[23][253],u_xpb_out[24][253],u_xpb_out[25][253],u_xpb_out[26][253],u_xpb_out[27][253],u_xpb_out[28][253],u_xpb_out[29][253],u_xpb_out[30][253],u_xpb_out[31][253],u_xpb_out[32][253],u_xpb_out[33][253],u_xpb_out[34][253],u_xpb_out[35][253],u_xpb_out[36][253],u_xpb_out[37][253],u_xpb_out[38][253],u_xpb_out[39][253],u_xpb_out[40][253],u_xpb_out[41][253],u_xpb_out[42][253],u_xpb_out[43][253],u_xpb_out[44][253],u_xpb_out[45][253],u_xpb_out[46][253],u_xpb_out[47][253],u_xpb_out[48][253],u_xpb_out[49][253],u_xpb_out[50][253],u_xpb_out[51][253],u_xpb_out[52][253],u_xpb_out[53][253],u_xpb_out[54][253],u_xpb_out[55][253],u_xpb_out[56][253],u_xpb_out[57][253],u_xpb_out[58][253],u_xpb_out[59][253],u_xpb_out[60][253],u_xpb_out[61][253],u_xpb_out[62][253],u_xpb_out[63][253],u_xpb_out[64][253],u_xpb_out[65][253],u_xpb_out[66][253],u_xpb_out[67][253],u_xpb_out[68][253],u_xpb_out[69][253],u_xpb_out[70][253],u_xpb_out[71][253],u_xpb_out[72][253],u_xpb_out[73][253],u_xpb_out[74][253],u_xpb_out[75][253],u_xpb_out[76][253],u_xpb_out[77][253],u_xpb_out[78][253],u_xpb_out[79][253],u_xpb_out[80][253],u_xpb_out[81][253],u_xpb_out[82][253],u_xpb_out[83][253],u_xpb_out[84][253],u_xpb_out[85][253],u_xpb_out[86][253],u_xpb_out[87][253],u_xpb_out[88][253],u_xpb_out[89][253],u_xpb_out[90][253],u_xpb_out[91][253],u_xpb_out[92][253],u_xpb_out[93][253],u_xpb_out[94][253],u_xpb_out[95][253],u_xpb_out[96][253],u_xpb_out[97][253],u_xpb_out[98][253],u_xpb_out[99][253],u_xpb_out[100][253],u_xpb_out[101][253],u_xpb_out[102][253],u_xpb_out[103][253],u_xpb_out[104][253],u_xpb_out[105][253]};

assign col_out_254 = {u_xpb_out[0][254],u_xpb_out[1][254],u_xpb_out[2][254],u_xpb_out[3][254],u_xpb_out[4][254],u_xpb_out[5][254],u_xpb_out[6][254],u_xpb_out[7][254],u_xpb_out[8][254],u_xpb_out[9][254],u_xpb_out[10][254],u_xpb_out[11][254],u_xpb_out[12][254],u_xpb_out[13][254],u_xpb_out[14][254],u_xpb_out[15][254],u_xpb_out[16][254],u_xpb_out[17][254],u_xpb_out[18][254],u_xpb_out[19][254],u_xpb_out[20][254],u_xpb_out[21][254],u_xpb_out[22][254],u_xpb_out[23][254],u_xpb_out[24][254],u_xpb_out[25][254],u_xpb_out[26][254],u_xpb_out[27][254],u_xpb_out[28][254],u_xpb_out[29][254],u_xpb_out[30][254],u_xpb_out[31][254],u_xpb_out[32][254],u_xpb_out[33][254],u_xpb_out[34][254],u_xpb_out[35][254],u_xpb_out[36][254],u_xpb_out[37][254],u_xpb_out[38][254],u_xpb_out[39][254],u_xpb_out[40][254],u_xpb_out[41][254],u_xpb_out[42][254],u_xpb_out[43][254],u_xpb_out[44][254],u_xpb_out[45][254],u_xpb_out[46][254],u_xpb_out[47][254],u_xpb_out[48][254],u_xpb_out[49][254],u_xpb_out[50][254],u_xpb_out[51][254],u_xpb_out[52][254],u_xpb_out[53][254],u_xpb_out[54][254],u_xpb_out[55][254],u_xpb_out[56][254],u_xpb_out[57][254],u_xpb_out[58][254],u_xpb_out[59][254],u_xpb_out[60][254],u_xpb_out[61][254],u_xpb_out[62][254],u_xpb_out[63][254],u_xpb_out[64][254],u_xpb_out[65][254],u_xpb_out[66][254],u_xpb_out[67][254],u_xpb_out[68][254],u_xpb_out[69][254],u_xpb_out[70][254],u_xpb_out[71][254],u_xpb_out[72][254],u_xpb_out[73][254],u_xpb_out[74][254],u_xpb_out[75][254],u_xpb_out[76][254],u_xpb_out[77][254],u_xpb_out[78][254],u_xpb_out[79][254],u_xpb_out[80][254],u_xpb_out[81][254],u_xpb_out[82][254],u_xpb_out[83][254],u_xpb_out[84][254],u_xpb_out[85][254],u_xpb_out[86][254],u_xpb_out[87][254],u_xpb_out[88][254],u_xpb_out[89][254],u_xpb_out[90][254],u_xpb_out[91][254],u_xpb_out[92][254],u_xpb_out[93][254],u_xpb_out[94][254],u_xpb_out[95][254],u_xpb_out[96][254],u_xpb_out[97][254],u_xpb_out[98][254],u_xpb_out[99][254],u_xpb_out[100][254],u_xpb_out[101][254],u_xpb_out[102][254],u_xpb_out[103][254],u_xpb_out[104][254],u_xpb_out[105][254]};

assign col_out_255 = {u_xpb_out[0][255],u_xpb_out[1][255],u_xpb_out[2][255],u_xpb_out[3][255],u_xpb_out[4][255],u_xpb_out[5][255],u_xpb_out[6][255],u_xpb_out[7][255],u_xpb_out[8][255],u_xpb_out[9][255],u_xpb_out[10][255],u_xpb_out[11][255],u_xpb_out[12][255],u_xpb_out[13][255],u_xpb_out[14][255],u_xpb_out[15][255],u_xpb_out[16][255],u_xpb_out[17][255],u_xpb_out[18][255],u_xpb_out[19][255],u_xpb_out[20][255],u_xpb_out[21][255],u_xpb_out[22][255],u_xpb_out[23][255],u_xpb_out[24][255],u_xpb_out[25][255],u_xpb_out[26][255],u_xpb_out[27][255],u_xpb_out[28][255],u_xpb_out[29][255],u_xpb_out[30][255],u_xpb_out[31][255],u_xpb_out[32][255],u_xpb_out[33][255],u_xpb_out[34][255],u_xpb_out[35][255],u_xpb_out[36][255],u_xpb_out[37][255],u_xpb_out[38][255],u_xpb_out[39][255],u_xpb_out[40][255],u_xpb_out[41][255],u_xpb_out[42][255],u_xpb_out[43][255],u_xpb_out[44][255],u_xpb_out[45][255],u_xpb_out[46][255],u_xpb_out[47][255],u_xpb_out[48][255],u_xpb_out[49][255],u_xpb_out[50][255],u_xpb_out[51][255],u_xpb_out[52][255],u_xpb_out[53][255],u_xpb_out[54][255],u_xpb_out[55][255],u_xpb_out[56][255],u_xpb_out[57][255],u_xpb_out[58][255],u_xpb_out[59][255],u_xpb_out[60][255],u_xpb_out[61][255],u_xpb_out[62][255],u_xpb_out[63][255],u_xpb_out[64][255],u_xpb_out[65][255],u_xpb_out[66][255],u_xpb_out[67][255],u_xpb_out[68][255],u_xpb_out[69][255],u_xpb_out[70][255],u_xpb_out[71][255],u_xpb_out[72][255],u_xpb_out[73][255],u_xpb_out[74][255],u_xpb_out[75][255],u_xpb_out[76][255],u_xpb_out[77][255],u_xpb_out[78][255],u_xpb_out[79][255],u_xpb_out[80][255],u_xpb_out[81][255],u_xpb_out[82][255],u_xpb_out[83][255],u_xpb_out[84][255],u_xpb_out[85][255],u_xpb_out[86][255],u_xpb_out[87][255],u_xpb_out[88][255],u_xpb_out[89][255],u_xpb_out[90][255],u_xpb_out[91][255],u_xpb_out[92][255],u_xpb_out[93][255],u_xpb_out[94][255],u_xpb_out[95][255],u_xpb_out[96][255],u_xpb_out[97][255],u_xpb_out[98][255],u_xpb_out[99][255],u_xpb_out[100][255],u_xpb_out[101][255],u_xpb_out[102][255],u_xpb_out[103][255],u_xpb_out[104][255],u_xpb_out[105][255]};

assign col_out_256 = {u_xpb_out[0][256],u_xpb_out[1][256],u_xpb_out[2][256],u_xpb_out[3][256],u_xpb_out[4][256],u_xpb_out[5][256],u_xpb_out[6][256],u_xpb_out[7][256],u_xpb_out[8][256],u_xpb_out[9][256],u_xpb_out[10][256],u_xpb_out[11][256],u_xpb_out[12][256],u_xpb_out[13][256],u_xpb_out[14][256],u_xpb_out[15][256],u_xpb_out[16][256],u_xpb_out[17][256],u_xpb_out[18][256],u_xpb_out[19][256],u_xpb_out[20][256],u_xpb_out[21][256],u_xpb_out[22][256],u_xpb_out[23][256],u_xpb_out[24][256],u_xpb_out[25][256],u_xpb_out[26][256],u_xpb_out[27][256],u_xpb_out[28][256],u_xpb_out[29][256],u_xpb_out[30][256],u_xpb_out[31][256],u_xpb_out[32][256],u_xpb_out[33][256],u_xpb_out[34][256],u_xpb_out[35][256],u_xpb_out[36][256],u_xpb_out[37][256],u_xpb_out[38][256],u_xpb_out[39][256],u_xpb_out[40][256],u_xpb_out[41][256],u_xpb_out[42][256],u_xpb_out[43][256],u_xpb_out[44][256],u_xpb_out[45][256],u_xpb_out[46][256],u_xpb_out[47][256],u_xpb_out[48][256],u_xpb_out[49][256],u_xpb_out[50][256],u_xpb_out[51][256],u_xpb_out[52][256],u_xpb_out[53][256],u_xpb_out[54][256],u_xpb_out[55][256],u_xpb_out[56][256],u_xpb_out[57][256],u_xpb_out[58][256],u_xpb_out[59][256],u_xpb_out[60][256],u_xpb_out[61][256],u_xpb_out[62][256],u_xpb_out[63][256],u_xpb_out[64][256],u_xpb_out[65][256],u_xpb_out[66][256],u_xpb_out[67][256],u_xpb_out[68][256],u_xpb_out[69][256],u_xpb_out[70][256],u_xpb_out[71][256],u_xpb_out[72][256],u_xpb_out[73][256],u_xpb_out[74][256],u_xpb_out[75][256],u_xpb_out[76][256],u_xpb_out[77][256],u_xpb_out[78][256],u_xpb_out[79][256],u_xpb_out[80][256],u_xpb_out[81][256],u_xpb_out[82][256],u_xpb_out[83][256],u_xpb_out[84][256],u_xpb_out[85][256],u_xpb_out[86][256],u_xpb_out[87][256],u_xpb_out[88][256],u_xpb_out[89][256],u_xpb_out[90][256],u_xpb_out[91][256],u_xpb_out[92][256],u_xpb_out[93][256],u_xpb_out[94][256],u_xpb_out[95][256],u_xpb_out[96][256],u_xpb_out[97][256],u_xpb_out[98][256],u_xpb_out[99][256],u_xpb_out[100][256],u_xpb_out[101][256],u_xpb_out[102][256],u_xpb_out[103][256],u_xpb_out[104][256],u_xpb_out[105][256]};

assign col_out_257 = {u_xpb_out[0][257],u_xpb_out[1][257],u_xpb_out[2][257],u_xpb_out[3][257],u_xpb_out[4][257],u_xpb_out[5][257],u_xpb_out[6][257],u_xpb_out[7][257],u_xpb_out[8][257],u_xpb_out[9][257],u_xpb_out[10][257],u_xpb_out[11][257],u_xpb_out[12][257],u_xpb_out[13][257],u_xpb_out[14][257],u_xpb_out[15][257],u_xpb_out[16][257],u_xpb_out[17][257],u_xpb_out[18][257],u_xpb_out[19][257],u_xpb_out[20][257],u_xpb_out[21][257],u_xpb_out[22][257],u_xpb_out[23][257],u_xpb_out[24][257],u_xpb_out[25][257],u_xpb_out[26][257],u_xpb_out[27][257],u_xpb_out[28][257],u_xpb_out[29][257],u_xpb_out[30][257],u_xpb_out[31][257],u_xpb_out[32][257],u_xpb_out[33][257],u_xpb_out[34][257],u_xpb_out[35][257],u_xpb_out[36][257],u_xpb_out[37][257],u_xpb_out[38][257],u_xpb_out[39][257],u_xpb_out[40][257],u_xpb_out[41][257],u_xpb_out[42][257],u_xpb_out[43][257],u_xpb_out[44][257],u_xpb_out[45][257],u_xpb_out[46][257],u_xpb_out[47][257],u_xpb_out[48][257],u_xpb_out[49][257],u_xpb_out[50][257],u_xpb_out[51][257],u_xpb_out[52][257],u_xpb_out[53][257],u_xpb_out[54][257],u_xpb_out[55][257],u_xpb_out[56][257],u_xpb_out[57][257],u_xpb_out[58][257],u_xpb_out[59][257],u_xpb_out[60][257],u_xpb_out[61][257],u_xpb_out[62][257],u_xpb_out[63][257],u_xpb_out[64][257],u_xpb_out[65][257],u_xpb_out[66][257],u_xpb_out[67][257],u_xpb_out[68][257],u_xpb_out[69][257],u_xpb_out[70][257],u_xpb_out[71][257],u_xpb_out[72][257],u_xpb_out[73][257],u_xpb_out[74][257],u_xpb_out[75][257],u_xpb_out[76][257],u_xpb_out[77][257],u_xpb_out[78][257],u_xpb_out[79][257],u_xpb_out[80][257],u_xpb_out[81][257],u_xpb_out[82][257],u_xpb_out[83][257],u_xpb_out[84][257],u_xpb_out[85][257],u_xpb_out[86][257],u_xpb_out[87][257],u_xpb_out[88][257],u_xpb_out[89][257],u_xpb_out[90][257],u_xpb_out[91][257],u_xpb_out[92][257],u_xpb_out[93][257],u_xpb_out[94][257],u_xpb_out[95][257],u_xpb_out[96][257],u_xpb_out[97][257],u_xpb_out[98][257],u_xpb_out[99][257],u_xpb_out[100][257],u_xpb_out[101][257],u_xpb_out[102][257],u_xpb_out[103][257],u_xpb_out[104][257],u_xpb_out[105][257]};

assign col_out_258 = {u_xpb_out[0][258],u_xpb_out[1][258],u_xpb_out[2][258],u_xpb_out[3][258],u_xpb_out[4][258],u_xpb_out[5][258],u_xpb_out[6][258],u_xpb_out[7][258],u_xpb_out[8][258],u_xpb_out[9][258],u_xpb_out[10][258],u_xpb_out[11][258],u_xpb_out[12][258],u_xpb_out[13][258],u_xpb_out[14][258],u_xpb_out[15][258],u_xpb_out[16][258],u_xpb_out[17][258],u_xpb_out[18][258],u_xpb_out[19][258],u_xpb_out[20][258],u_xpb_out[21][258],u_xpb_out[22][258],u_xpb_out[23][258],u_xpb_out[24][258],u_xpb_out[25][258],u_xpb_out[26][258],u_xpb_out[27][258],u_xpb_out[28][258],u_xpb_out[29][258],u_xpb_out[30][258],u_xpb_out[31][258],u_xpb_out[32][258],u_xpb_out[33][258],u_xpb_out[34][258],u_xpb_out[35][258],u_xpb_out[36][258],u_xpb_out[37][258],u_xpb_out[38][258],u_xpb_out[39][258],u_xpb_out[40][258],u_xpb_out[41][258],u_xpb_out[42][258],u_xpb_out[43][258],u_xpb_out[44][258],u_xpb_out[45][258],u_xpb_out[46][258],u_xpb_out[47][258],u_xpb_out[48][258],u_xpb_out[49][258],u_xpb_out[50][258],u_xpb_out[51][258],u_xpb_out[52][258],u_xpb_out[53][258],u_xpb_out[54][258],u_xpb_out[55][258],u_xpb_out[56][258],u_xpb_out[57][258],u_xpb_out[58][258],u_xpb_out[59][258],u_xpb_out[60][258],u_xpb_out[61][258],u_xpb_out[62][258],u_xpb_out[63][258],u_xpb_out[64][258],u_xpb_out[65][258],u_xpb_out[66][258],u_xpb_out[67][258],u_xpb_out[68][258],u_xpb_out[69][258],u_xpb_out[70][258],u_xpb_out[71][258],u_xpb_out[72][258],u_xpb_out[73][258],u_xpb_out[74][258],u_xpb_out[75][258],u_xpb_out[76][258],u_xpb_out[77][258],u_xpb_out[78][258],u_xpb_out[79][258],u_xpb_out[80][258],u_xpb_out[81][258],u_xpb_out[82][258],u_xpb_out[83][258],u_xpb_out[84][258],u_xpb_out[85][258],u_xpb_out[86][258],u_xpb_out[87][258],u_xpb_out[88][258],u_xpb_out[89][258],u_xpb_out[90][258],u_xpb_out[91][258],u_xpb_out[92][258],u_xpb_out[93][258],u_xpb_out[94][258],u_xpb_out[95][258],u_xpb_out[96][258],u_xpb_out[97][258],u_xpb_out[98][258],u_xpb_out[99][258],u_xpb_out[100][258],u_xpb_out[101][258],u_xpb_out[102][258],u_xpb_out[103][258],u_xpb_out[104][258],u_xpb_out[105][258]};

assign col_out_259 = {u_xpb_out[0][259],u_xpb_out[1][259],u_xpb_out[2][259],u_xpb_out[3][259],u_xpb_out[4][259],u_xpb_out[5][259],u_xpb_out[6][259],u_xpb_out[7][259],u_xpb_out[8][259],u_xpb_out[9][259],u_xpb_out[10][259],u_xpb_out[11][259],u_xpb_out[12][259],u_xpb_out[13][259],u_xpb_out[14][259],u_xpb_out[15][259],u_xpb_out[16][259],u_xpb_out[17][259],u_xpb_out[18][259],u_xpb_out[19][259],u_xpb_out[20][259],u_xpb_out[21][259],u_xpb_out[22][259],u_xpb_out[23][259],u_xpb_out[24][259],u_xpb_out[25][259],u_xpb_out[26][259],u_xpb_out[27][259],u_xpb_out[28][259],u_xpb_out[29][259],u_xpb_out[30][259],u_xpb_out[31][259],u_xpb_out[32][259],u_xpb_out[33][259],u_xpb_out[34][259],u_xpb_out[35][259],u_xpb_out[36][259],u_xpb_out[37][259],u_xpb_out[38][259],u_xpb_out[39][259],u_xpb_out[40][259],u_xpb_out[41][259],u_xpb_out[42][259],u_xpb_out[43][259],u_xpb_out[44][259],u_xpb_out[45][259],u_xpb_out[46][259],u_xpb_out[47][259],u_xpb_out[48][259],u_xpb_out[49][259],u_xpb_out[50][259],u_xpb_out[51][259],u_xpb_out[52][259],u_xpb_out[53][259],u_xpb_out[54][259],u_xpb_out[55][259],u_xpb_out[56][259],u_xpb_out[57][259],u_xpb_out[58][259],u_xpb_out[59][259],u_xpb_out[60][259],u_xpb_out[61][259],u_xpb_out[62][259],u_xpb_out[63][259],u_xpb_out[64][259],u_xpb_out[65][259],u_xpb_out[66][259],u_xpb_out[67][259],u_xpb_out[68][259],u_xpb_out[69][259],u_xpb_out[70][259],u_xpb_out[71][259],u_xpb_out[72][259],u_xpb_out[73][259],u_xpb_out[74][259],u_xpb_out[75][259],u_xpb_out[76][259],u_xpb_out[77][259],u_xpb_out[78][259],u_xpb_out[79][259],u_xpb_out[80][259],u_xpb_out[81][259],u_xpb_out[82][259],u_xpb_out[83][259],u_xpb_out[84][259],u_xpb_out[85][259],u_xpb_out[86][259],u_xpb_out[87][259],u_xpb_out[88][259],u_xpb_out[89][259],u_xpb_out[90][259],u_xpb_out[91][259],u_xpb_out[92][259],u_xpb_out[93][259],u_xpb_out[94][259],u_xpb_out[95][259],u_xpb_out[96][259],u_xpb_out[97][259],u_xpb_out[98][259],u_xpb_out[99][259],u_xpb_out[100][259],u_xpb_out[101][259],u_xpb_out[102][259],u_xpb_out[103][259],u_xpb_out[104][259],u_xpb_out[105][259]};

assign col_out_260 = {u_xpb_out[0][260],u_xpb_out[1][260],u_xpb_out[2][260],u_xpb_out[3][260],u_xpb_out[4][260],u_xpb_out[5][260],u_xpb_out[6][260],u_xpb_out[7][260],u_xpb_out[8][260],u_xpb_out[9][260],u_xpb_out[10][260],u_xpb_out[11][260],u_xpb_out[12][260],u_xpb_out[13][260],u_xpb_out[14][260],u_xpb_out[15][260],u_xpb_out[16][260],u_xpb_out[17][260],u_xpb_out[18][260],u_xpb_out[19][260],u_xpb_out[20][260],u_xpb_out[21][260],u_xpb_out[22][260],u_xpb_out[23][260],u_xpb_out[24][260],u_xpb_out[25][260],u_xpb_out[26][260],u_xpb_out[27][260],u_xpb_out[28][260],u_xpb_out[29][260],u_xpb_out[30][260],u_xpb_out[31][260],u_xpb_out[32][260],u_xpb_out[33][260],u_xpb_out[34][260],u_xpb_out[35][260],u_xpb_out[36][260],u_xpb_out[37][260],u_xpb_out[38][260],u_xpb_out[39][260],u_xpb_out[40][260],u_xpb_out[41][260],u_xpb_out[42][260],u_xpb_out[43][260],u_xpb_out[44][260],u_xpb_out[45][260],u_xpb_out[46][260],u_xpb_out[47][260],u_xpb_out[48][260],u_xpb_out[49][260],u_xpb_out[50][260],u_xpb_out[51][260],u_xpb_out[52][260],u_xpb_out[53][260],u_xpb_out[54][260],u_xpb_out[55][260],u_xpb_out[56][260],u_xpb_out[57][260],u_xpb_out[58][260],u_xpb_out[59][260],u_xpb_out[60][260],u_xpb_out[61][260],u_xpb_out[62][260],u_xpb_out[63][260],u_xpb_out[64][260],u_xpb_out[65][260],u_xpb_out[66][260],u_xpb_out[67][260],u_xpb_out[68][260],u_xpb_out[69][260],u_xpb_out[70][260],u_xpb_out[71][260],u_xpb_out[72][260],u_xpb_out[73][260],u_xpb_out[74][260],u_xpb_out[75][260],u_xpb_out[76][260],u_xpb_out[77][260],u_xpb_out[78][260],u_xpb_out[79][260],u_xpb_out[80][260],u_xpb_out[81][260],u_xpb_out[82][260],u_xpb_out[83][260],u_xpb_out[84][260],u_xpb_out[85][260],u_xpb_out[86][260],u_xpb_out[87][260],u_xpb_out[88][260],u_xpb_out[89][260],u_xpb_out[90][260],u_xpb_out[91][260],u_xpb_out[92][260],u_xpb_out[93][260],u_xpb_out[94][260],u_xpb_out[95][260],u_xpb_out[96][260],u_xpb_out[97][260],u_xpb_out[98][260],u_xpb_out[99][260],u_xpb_out[100][260],u_xpb_out[101][260],u_xpb_out[102][260],u_xpb_out[103][260],u_xpb_out[104][260],u_xpb_out[105][260]};

assign col_out_261 = {u_xpb_out[0][261],u_xpb_out[1][261],u_xpb_out[2][261],u_xpb_out[3][261],u_xpb_out[4][261],u_xpb_out[5][261],u_xpb_out[6][261],u_xpb_out[7][261],u_xpb_out[8][261],u_xpb_out[9][261],u_xpb_out[10][261],u_xpb_out[11][261],u_xpb_out[12][261],u_xpb_out[13][261],u_xpb_out[14][261],u_xpb_out[15][261],u_xpb_out[16][261],u_xpb_out[17][261],u_xpb_out[18][261],u_xpb_out[19][261],u_xpb_out[20][261],u_xpb_out[21][261],u_xpb_out[22][261],u_xpb_out[23][261],u_xpb_out[24][261],u_xpb_out[25][261],u_xpb_out[26][261],u_xpb_out[27][261],u_xpb_out[28][261],u_xpb_out[29][261],u_xpb_out[30][261],u_xpb_out[31][261],u_xpb_out[32][261],u_xpb_out[33][261],u_xpb_out[34][261],u_xpb_out[35][261],u_xpb_out[36][261],u_xpb_out[37][261],u_xpb_out[38][261],u_xpb_out[39][261],u_xpb_out[40][261],u_xpb_out[41][261],u_xpb_out[42][261],u_xpb_out[43][261],u_xpb_out[44][261],u_xpb_out[45][261],u_xpb_out[46][261],u_xpb_out[47][261],u_xpb_out[48][261],u_xpb_out[49][261],u_xpb_out[50][261],u_xpb_out[51][261],u_xpb_out[52][261],u_xpb_out[53][261],u_xpb_out[54][261],u_xpb_out[55][261],u_xpb_out[56][261],u_xpb_out[57][261],u_xpb_out[58][261],u_xpb_out[59][261],u_xpb_out[60][261],u_xpb_out[61][261],u_xpb_out[62][261],u_xpb_out[63][261],u_xpb_out[64][261],u_xpb_out[65][261],u_xpb_out[66][261],u_xpb_out[67][261],u_xpb_out[68][261],u_xpb_out[69][261],u_xpb_out[70][261],u_xpb_out[71][261],u_xpb_out[72][261],u_xpb_out[73][261],u_xpb_out[74][261],u_xpb_out[75][261],u_xpb_out[76][261],u_xpb_out[77][261],u_xpb_out[78][261],u_xpb_out[79][261],u_xpb_out[80][261],u_xpb_out[81][261],u_xpb_out[82][261],u_xpb_out[83][261],u_xpb_out[84][261],u_xpb_out[85][261],u_xpb_out[86][261],u_xpb_out[87][261],u_xpb_out[88][261],u_xpb_out[89][261],u_xpb_out[90][261],u_xpb_out[91][261],u_xpb_out[92][261],u_xpb_out[93][261],u_xpb_out[94][261],u_xpb_out[95][261],u_xpb_out[96][261],u_xpb_out[97][261],u_xpb_out[98][261],u_xpb_out[99][261],u_xpb_out[100][261],u_xpb_out[101][261],u_xpb_out[102][261],u_xpb_out[103][261],u_xpb_out[104][261],u_xpb_out[105][261]};

assign col_out_262 = {u_xpb_out[0][262],u_xpb_out[1][262],u_xpb_out[2][262],u_xpb_out[3][262],u_xpb_out[4][262],u_xpb_out[5][262],u_xpb_out[6][262],u_xpb_out[7][262],u_xpb_out[8][262],u_xpb_out[9][262],u_xpb_out[10][262],u_xpb_out[11][262],u_xpb_out[12][262],u_xpb_out[13][262],u_xpb_out[14][262],u_xpb_out[15][262],u_xpb_out[16][262],u_xpb_out[17][262],u_xpb_out[18][262],u_xpb_out[19][262],u_xpb_out[20][262],u_xpb_out[21][262],u_xpb_out[22][262],u_xpb_out[23][262],u_xpb_out[24][262],u_xpb_out[25][262],u_xpb_out[26][262],u_xpb_out[27][262],u_xpb_out[28][262],u_xpb_out[29][262],u_xpb_out[30][262],u_xpb_out[31][262],u_xpb_out[32][262],u_xpb_out[33][262],u_xpb_out[34][262],u_xpb_out[35][262],u_xpb_out[36][262],u_xpb_out[37][262],u_xpb_out[38][262],u_xpb_out[39][262],u_xpb_out[40][262],u_xpb_out[41][262],u_xpb_out[42][262],u_xpb_out[43][262],u_xpb_out[44][262],u_xpb_out[45][262],u_xpb_out[46][262],u_xpb_out[47][262],u_xpb_out[48][262],u_xpb_out[49][262],u_xpb_out[50][262],u_xpb_out[51][262],u_xpb_out[52][262],u_xpb_out[53][262],u_xpb_out[54][262],u_xpb_out[55][262],u_xpb_out[56][262],u_xpb_out[57][262],u_xpb_out[58][262],u_xpb_out[59][262],u_xpb_out[60][262],u_xpb_out[61][262],u_xpb_out[62][262],u_xpb_out[63][262],u_xpb_out[64][262],u_xpb_out[65][262],u_xpb_out[66][262],u_xpb_out[67][262],u_xpb_out[68][262],u_xpb_out[69][262],u_xpb_out[70][262],u_xpb_out[71][262],u_xpb_out[72][262],u_xpb_out[73][262],u_xpb_out[74][262],u_xpb_out[75][262],u_xpb_out[76][262],u_xpb_out[77][262],u_xpb_out[78][262],u_xpb_out[79][262],u_xpb_out[80][262],u_xpb_out[81][262],u_xpb_out[82][262],u_xpb_out[83][262],u_xpb_out[84][262],u_xpb_out[85][262],u_xpb_out[86][262],u_xpb_out[87][262],u_xpb_out[88][262],u_xpb_out[89][262],u_xpb_out[90][262],u_xpb_out[91][262],u_xpb_out[92][262],u_xpb_out[93][262],u_xpb_out[94][262],u_xpb_out[95][262],u_xpb_out[96][262],u_xpb_out[97][262],u_xpb_out[98][262],u_xpb_out[99][262],u_xpb_out[100][262],u_xpb_out[101][262],u_xpb_out[102][262],u_xpb_out[103][262],u_xpb_out[104][262],u_xpb_out[105][262]};

assign col_out_263 = {u_xpb_out[0][263],u_xpb_out[1][263],u_xpb_out[2][263],u_xpb_out[3][263],u_xpb_out[4][263],u_xpb_out[5][263],u_xpb_out[6][263],u_xpb_out[7][263],u_xpb_out[8][263],u_xpb_out[9][263],u_xpb_out[10][263],u_xpb_out[11][263],u_xpb_out[12][263],u_xpb_out[13][263],u_xpb_out[14][263],u_xpb_out[15][263],u_xpb_out[16][263],u_xpb_out[17][263],u_xpb_out[18][263],u_xpb_out[19][263],u_xpb_out[20][263],u_xpb_out[21][263],u_xpb_out[22][263],u_xpb_out[23][263],u_xpb_out[24][263],u_xpb_out[25][263],u_xpb_out[26][263],u_xpb_out[27][263],u_xpb_out[28][263],u_xpb_out[29][263],u_xpb_out[30][263],u_xpb_out[31][263],u_xpb_out[32][263],u_xpb_out[33][263],u_xpb_out[34][263],u_xpb_out[35][263],u_xpb_out[36][263],u_xpb_out[37][263],u_xpb_out[38][263],u_xpb_out[39][263],u_xpb_out[40][263],u_xpb_out[41][263],u_xpb_out[42][263],u_xpb_out[43][263],u_xpb_out[44][263],u_xpb_out[45][263],u_xpb_out[46][263],u_xpb_out[47][263],u_xpb_out[48][263],u_xpb_out[49][263],u_xpb_out[50][263],u_xpb_out[51][263],u_xpb_out[52][263],u_xpb_out[53][263],u_xpb_out[54][263],u_xpb_out[55][263],u_xpb_out[56][263],u_xpb_out[57][263],u_xpb_out[58][263],u_xpb_out[59][263],u_xpb_out[60][263],u_xpb_out[61][263],u_xpb_out[62][263],u_xpb_out[63][263],u_xpb_out[64][263],u_xpb_out[65][263],u_xpb_out[66][263],u_xpb_out[67][263],u_xpb_out[68][263],u_xpb_out[69][263],u_xpb_out[70][263],u_xpb_out[71][263],u_xpb_out[72][263],u_xpb_out[73][263],u_xpb_out[74][263],u_xpb_out[75][263],u_xpb_out[76][263],u_xpb_out[77][263],u_xpb_out[78][263],u_xpb_out[79][263],u_xpb_out[80][263],u_xpb_out[81][263],u_xpb_out[82][263],u_xpb_out[83][263],u_xpb_out[84][263],u_xpb_out[85][263],u_xpb_out[86][263],u_xpb_out[87][263],u_xpb_out[88][263],u_xpb_out[89][263],u_xpb_out[90][263],u_xpb_out[91][263],u_xpb_out[92][263],u_xpb_out[93][263],u_xpb_out[94][263],u_xpb_out[95][263],u_xpb_out[96][263],u_xpb_out[97][263],u_xpb_out[98][263],u_xpb_out[99][263],u_xpb_out[100][263],u_xpb_out[101][263],u_xpb_out[102][263],u_xpb_out[103][263],u_xpb_out[104][263],u_xpb_out[105][263]};

assign col_out_264 = {u_xpb_out[0][264],u_xpb_out[1][264],u_xpb_out[2][264],u_xpb_out[3][264],u_xpb_out[4][264],u_xpb_out[5][264],u_xpb_out[6][264],u_xpb_out[7][264],u_xpb_out[8][264],u_xpb_out[9][264],u_xpb_out[10][264],u_xpb_out[11][264],u_xpb_out[12][264],u_xpb_out[13][264],u_xpb_out[14][264],u_xpb_out[15][264],u_xpb_out[16][264],u_xpb_out[17][264],u_xpb_out[18][264],u_xpb_out[19][264],u_xpb_out[20][264],u_xpb_out[21][264],u_xpb_out[22][264],u_xpb_out[23][264],u_xpb_out[24][264],u_xpb_out[25][264],u_xpb_out[26][264],u_xpb_out[27][264],u_xpb_out[28][264],u_xpb_out[29][264],u_xpb_out[30][264],u_xpb_out[31][264],u_xpb_out[32][264],u_xpb_out[33][264],u_xpb_out[34][264],u_xpb_out[35][264],u_xpb_out[36][264],u_xpb_out[37][264],u_xpb_out[38][264],u_xpb_out[39][264],u_xpb_out[40][264],u_xpb_out[41][264],u_xpb_out[42][264],u_xpb_out[43][264],u_xpb_out[44][264],u_xpb_out[45][264],u_xpb_out[46][264],u_xpb_out[47][264],u_xpb_out[48][264],u_xpb_out[49][264],u_xpb_out[50][264],u_xpb_out[51][264],u_xpb_out[52][264],u_xpb_out[53][264],u_xpb_out[54][264],u_xpb_out[55][264],u_xpb_out[56][264],u_xpb_out[57][264],u_xpb_out[58][264],u_xpb_out[59][264],u_xpb_out[60][264],u_xpb_out[61][264],u_xpb_out[62][264],u_xpb_out[63][264],u_xpb_out[64][264],u_xpb_out[65][264],u_xpb_out[66][264],u_xpb_out[67][264],u_xpb_out[68][264],u_xpb_out[69][264],u_xpb_out[70][264],u_xpb_out[71][264],u_xpb_out[72][264],u_xpb_out[73][264],u_xpb_out[74][264],u_xpb_out[75][264],u_xpb_out[76][264],u_xpb_out[77][264],u_xpb_out[78][264],u_xpb_out[79][264],u_xpb_out[80][264],u_xpb_out[81][264],u_xpb_out[82][264],u_xpb_out[83][264],u_xpb_out[84][264],u_xpb_out[85][264],u_xpb_out[86][264],u_xpb_out[87][264],u_xpb_out[88][264],u_xpb_out[89][264],u_xpb_out[90][264],u_xpb_out[91][264],u_xpb_out[92][264],u_xpb_out[93][264],u_xpb_out[94][264],u_xpb_out[95][264],u_xpb_out[96][264],u_xpb_out[97][264],u_xpb_out[98][264],u_xpb_out[99][264],u_xpb_out[100][264],u_xpb_out[101][264],u_xpb_out[102][264],u_xpb_out[103][264],u_xpb_out[104][264],u_xpb_out[105][264]};

assign col_out_265 = {u_xpb_out[0][265],u_xpb_out[1][265],u_xpb_out[2][265],u_xpb_out[3][265],u_xpb_out[4][265],u_xpb_out[5][265],u_xpb_out[6][265],u_xpb_out[7][265],u_xpb_out[8][265],u_xpb_out[9][265],u_xpb_out[10][265],u_xpb_out[11][265],u_xpb_out[12][265],u_xpb_out[13][265],u_xpb_out[14][265],u_xpb_out[15][265],u_xpb_out[16][265],u_xpb_out[17][265],u_xpb_out[18][265],u_xpb_out[19][265],u_xpb_out[20][265],u_xpb_out[21][265],u_xpb_out[22][265],u_xpb_out[23][265],u_xpb_out[24][265],u_xpb_out[25][265],u_xpb_out[26][265],u_xpb_out[27][265],u_xpb_out[28][265],u_xpb_out[29][265],u_xpb_out[30][265],u_xpb_out[31][265],u_xpb_out[32][265],u_xpb_out[33][265],u_xpb_out[34][265],u_xpb_out[35][265],u_xpb_out[36][265],u_xpb_out[37][265],u_xpb_out[38][265],u_xpb_out[39][265],u_xpb_out[40][265],u_xpb_out[41][265],u_xpb_out[42][265],u_xpb_out[43][265],u_xpb_out[44][265],u_xpb_out[45][265],u_xpb_out[46][265],u_xpb_out[47][265],u_xpb_out[48][265],u_xpb_out[49][265],u_xpb_out[50][265],u_xpb_out[51][265],u_xpb_out[52][265],u_xpb_out[53][265],u_xpb_out[54][265],u_xpb_out[55][265],u_xpb_out[56][265],u_xpb_out[57][265],u_xpb_out[58][265],u_xpb_out[59][265],u_xpb_out[60][265],u_xpb_out[61][265],u_xpb_out[62][265],u_xpb_out[63][265],u_xpb_out[64][265],u_xpb_out[65][265],u_xpb_out[66][265],u_xpb_out[67][265],u_xpb_out[68][265],u_xpb_out[69][265],u_xpb_out[70][265],u_xpb_out[71][265],u_xpb_out[72][265],u_xpb_out[73][265],u_xpb_out[74][265],u_xpb_out[75][265],u_xpb_out[76][265],u_xpb_out[77][265],u_xpb_out[78][265],u_xpb_out[79][265],u_xpb_out[80][265],u_xpb_out[81][265],u_xpb_out[82][265],u_xpb_out[83][265],u_xpb_out[84][265],u_xpb_out[85][265],u_xpb_out[86][265],u_xpb_out[87][265],u_xpb_out[88][265],u_xpb_out[89][265],u_xpb_out[90][265],u_xpb_out[91][265],u_xpb_out[92][265],u_xpb_out[93][265],u_xpb_out[94][265],u_xpb_out[95][265],u_xpb_out[96][265],u_xpb_out[97][265],u_xpb_out[98][265],u_xpb_out[99][265],u_xpb_out[100][265],u_xpb_out[101][265],u_xpb_out[102][265],u_xpb_out[103][265],u_xpb_out[104][265],u_xpb_out[105][265]};

assign col_out_266 = {u_xpb_out[0][266],u_xpb_out[1][266],u_xpb_out[2][266],u_xpb_out[3][266],u_xpb_out[4][266],u_xpb_out[5][266],u_xpb_out[6][266],u_xpb_out[7][266],u_xpb_out[8][266],u_xpb_out[9][266],u_xpb_out[10][266],u_xpb_out[11][266],u_xpb_out[12][266],u_xpb_out[13][266],u_xpb_out[14][266],u_xpb_out[15][266],u_xpb_out[16][266],u_xpb_out[17][266],u_xpb_out[18][266],u_xpb_out[19][266],u_xpb_out[20][266],u_xpb_out[21][266],u_xpb_out[22][266],u_xpb_out[23][266],u_xpb_out[24][266],u_xpb_out[25][266],u_xpb_out[26][266],u_xpb_out[27][266],u_xpb_out[28][266],u_xpb_out[29][266],u_xpb_out[30][266],u_xpb_out[31][266],u_xpb_out[32][266],u_xpb_out[33][266],u_xpb_out[34][266],u_xpb_out[35][266],u_xpb_out[36][266],u_xpb_out[37][266],u_xpb_out[38][266],u_xpb_out[39][266],u_xpb_out[40][266],u_xpb_out[41][266],u_xpb_out[42][266],u_xpb_out[43][266],u_xpb_out[44][266],u_xpb_out[45][266],u_xpb_out[46][266],u_xpb_out[47][266],u_xpb_out[48][266],u_xpb_out[49][266],u_xpb_out[50][266],u_xpb_out[51][266],u_xpb_out[52][266],u_xpb_out[53][266],u_xpb_out[54][266],u_xpb_out[55][266],u_xpb_out[56][266],u_xpb_out[57][266],u_xpb_out[58][266],u_xpb_out[59][266],u_xpb_out[60][266],u_xpb_out[61][266],u_xpb_out[62][266],u_xpb_out[63][266],u_xpb_out[64][266],u_xpb_out[65][266],u_xpb_out[66][266],u_xpb_out[67][266],u_xpb_out[68][266],u_xpb_out[69][266],u_xpb_out[70][266],u_xpb_out[71][266],u_xpb_out[72][266],u_xpb_out[73][266],u_xpb_out[74][266],u_xpb_out[75][266],u_xpb_out[76][266],u_xpb_out[77][266],u_xpb_out[78][266],u_xpb_out[79][266],u_xpb_out[80][266],u_xpb_out[81][266],u_xpb_out[82][266],u_xpb_out[83][266],u_xpb_out[84][266],u_xpb_out[85][266],u_xpb_out[86][266],u_xpb_out[87][266],u_xpb_out[88][266],u_xpb_out[89][266],u_xpb_out[90][266],u_xpb_out[91][266],u_xpb_out[92][266],u_xpb_out[93][266],u_xpb_out[94][266],u_xpb_out[95][266],u_xpb_out[96][266],u_xpb_out[97][266],u_xpb_out[98][266],u_xpb_out[99][266],u_xpb_out[100][266],u_xpb_out[101][266],u_xpb_out[102][266],u_xpb_out[103][266],u_xpb_out[104][266],u_xpb_out[105][266]};

assign col_out_267 = {u_xpb_out[0][267],u_xpb_out[1][267],u_xpb_out[2][267],u_xpb_out[3][267],u_xpb_out[4][267],u_xpb_out[5][267],u_xpb_out[6][267],u_xpb_out[7][267],u_xpb_out[8][267],u_xpb_out[9][267],u_xpb_out[10][267],u_xpb_out[11][267],u_xpb_out[12][267],u_xpb_out[13][267],u_xpb_out[14][267],u_xpb_out[15][267],u_xpb_out[16][267],u_xpb_out[17][267],u_xpb_out[18][267],u_xpb_out[19][267],u_xpb_out[20][267],u_xpb_out[21][267],u_xpb_out[22][267],u_xpb_out[23][267],u_xpb_out[24][267],u_xpb_out[25][267],u_xpb_out[26][267],u_xpb_out[27][267],u_xpb_out[28][267],u_xpb_out[29][267],u_xpb_out[30][267],u_xpb_out[31][267],u_xpb_out[32][267],u_xpb_out[33][267],u_xpb_out[34][267],u_xpb_out[35][267],u_xpb_out[36][267],u_xpb_out[37][267],u_xpb_out[38][267],u_xpb_out[39][267],u_xpb_out[40][267],u_xpb_out[41][267],u_xpb_out[42][267],u_xpb_out[43][267],u_xpb_out[44][267],u_xpb_out[45][267],u_xpb_out[46][267],u_xpb_out[47][267],u_xpb_out[48][267],u_xpb_out[49][267],u_xpb_out[50][267],u_xpb_out[51][267],u_xpb_out[52][267],u_xpb_out[53][267],u_xpb_out[54][267],u_xpb_out[55][267],u_xpb_out[56][267],u_xpb_out[57][267],u_xpb_out[58][267],u_xpb_out[59][267],u_xpb_out[60][267],u_xpb_out[61][267],u_xpb_out[62][267],u_xpb_out[63][267],u_xpb_out[64][267],u_xpb_out[65][267],u_xpb_out[66][267],u_xpb_out[67][267],u_xpb_out[68][267],u_xpb_out[69][267],u_xpb_out[70][267],u_xpb_out[71][267],u_xpb_out[72][267],u_xpb_out[73][267],u_xpb_out[74][267],u_xpb_out[75][267],u_xpb_out[76][267],u_xpb_out[77][267],u_xpb_out[78][267],u_xpb_out[79][267],u_xpb_out[80][267],u_xpb_out[81][267],u_xpb_out[82][267],u_xpb_out[83][267],u_xpb_out[84][267],u_xpb_out[85][267],u_xpb_out[86][267],u_xpb_out[87][267],u_xpb_out[88][267],u_xpb_out[89][267],u_xpb_out[90][267],u_xpb_out[91][267],u_xpb_out[92][267],u_xpb_out[93][267],u_xpb_out[94][267],u_xpb_out[95][267],u_xpb_out[96][267],u_xpb_out[97][267],u_xpb_out[98][267],u_xpb_out[99][267],u_xpb_out[100][267],u_xpb_out[101][267],u_xpb_out[102][267],u_xpb_out[103][267],u_xpb_out[104][267],u_xpb_out[105][267]};

assign col_out_268 = {u_xpb_out[0][268],u_xpb_out[1][268],u_xpb_out[2][268],u_xpb_out[3][268],u_xpb_out[4][268],u_xpb_out[5][268],u_xpb_out[6][268],u_xpb_out[7][268],u_xpb_out[8][268],u_xpb_out[9][268],u_xpb_out[10][268],u_xpb_out[11][268],u_xpb_out[12][268],u_xpb_out[13][268],u_xpb_out[14][268],u_xpb_out[15][268],u_xpb_out[16][268],u_xpb_out[17][268],u_xpb_out[18][268],u_xpb_out[19][268],u_xpb_out[20][268],u_xpb_out[21][268],u_xpb_out[22][268],u_xpb_out[23][268],u_xpb_out[24][268],u_xpb_out[25][268],u_xpb_out[26][268],u_xpb_out[27][268],u_xpb_out[28][268],u_xpb_out[29][268],u_xpb_out[30][268],u_xpb_out[31][268],u_xpb_out[32][268],u_xpb_out[33][268],u_xpb_out[34][268],u_xpb_out[35][268],u_xpb_out[36][268],u_xpb_out[37][268],u_xpb_out[38][268],u_xpb_out[39][268],u_xpb_out[40][268],u_xpb_out[41][268],u_xpb_out[42][268],u_xpb_out[43][268],u_xpb_out[44][268],u_xpb_out[45][268],u_xpb_out[46][268],u_xpb_out[47][268],u_xpb_out[48][268],u_xpb_out[49][268],u_xpb_out[50][268],u_xpb_out[51][268],u_xpb_out[52][268],u_xpb_out[53][268],u_xpb_out[54][268],u_xpb_out[55][268],u_xpb_out[56][268],u_xpb_out[57][268],u_xpb_out[58][268],u_xpb_out[59][268],u_xpb_out[60][268],u_xpb_out[61][268],u_xpb_out[62][268],u_xpb_out[63][268],u_xpb_out[64][268],u_xpb_out[65][268],u_xpb_out[66][268],u_xpb_out[67][268],u_xpb_out[68][268],u_xpb_out[69][268],u_xpb_out[70][268],u_xpb_out[71][268],u_xpb_out[72][268],u_xpb_out[73][268],u_xpb_out[74][268],u_xpb_out[75][268],u_xpb_out[76][268],u_xpb_out[77][268],u_xpb_out[78][268],u_xpb_out[79][268],u_xpb_out[80][268],u_xpb_out[81][268],u_xpb_out[82][268],u_xpb_out[83][268],u_xpb_out[84][268],u_xpb_out[85][268],u_xpb_out[86][268],u_xpb_out[87][268],u_xpb_out[88][268],u_xpb_out[89][268],u_xpb_out[90][268],u_xpb_out[91][268],u_xpb_out[92][268],u_xpb_out[93][268],u_xpb_out[94][268],u_xpb_out[95][268],u_xpb_out[96][268],u_xpb_out[97][268],u_xpb_out[98][268],u_xpb_out[99][268],u_xpb_out[100][268],u_xpb_out[101][268],u_xpb_out[102][268],u_xpb_out[103][268],u_xpb_out[104][268],u_xpb_out[105][268]};

assign col_out_269 = {u_xpb_out[0][269],u_xpb_out[1][269],u_xpb_out[2][269],u_xpb_out[3][269],u_xpb_out[4][269],u_xpb_out[5][269],u_xpb_out[6][269],u_xpb_out[7][269],u_xpb_out[8][269],u_xpb_out[9][269],u_xpb_out[10][269],u_xpb_out[11][269],u_xpb_out[12][269],u_xpb_out[13][269],u_xpb_out[14][269],u_xpb_out[15][269],u_xpb_out[16][269],u_xpb_out[17][269],u_xpb_out[18][269],u_xpb_out[19][269],u_xpb_out[20][269],u_xpb_out[21][269],u_xpb_out[22][269],u_xpb_out[23][269],u_xpb_out[24][269],u_xpb_out[25][269],u_xpb_out[26][269],u_xpb_out[27][269],u_xpb_out[28][269],u_xpb_out[29][269],u_xpb_out[30][269],u_xpb_out[31][269],u_xpb_out[32][269],u_xpb_out[33][269],u_xpb_out[34][269],u_xpb_out[35][269],u_xpb_out[36][269],u_xpb_out[37][269],u_xpb_out[38][269],u_xpb_out[39][269],u_xpb_out[40][269],u_xpb_out[41][269],u_xpb_out[42][269],u_xpb_out[43][269],u_xpb_out[44][269],u_xpb_out[45][269],u_xpb_out[46][269],u_xpb_out[47][269],u_xpb_out[48][269],u_xpb_out[49][269],u_xpb_out[50][269],u_xpb_out[51][269],u_xpb_out[52][269],u_xpb_out[53][269],u_xpb_out[54][269],u_xpb_out[55][269],u_xpb_out[56][269],u_xpb_out[57][269],u_xpb_out[58][269],u_xpb_out[59][269],u_xpb_out[60][269],u_xpb_out[61][269],u_xpb_out[62][269],u_xpb_out[63][269],u_xpb_out[64][269],u_xpb_out[65][269],u_xpb_out[66][269],u_xpb_out[67][269],u_xpb_out[68][269],u_xpb_out[69][269],u_xpb_out[70][269],u_xpb_out[71][269],u_xpb_out[72][269],u_xpb_out[73][269],u_xpb_out[74][269],u_xpb_out[75][269],u_xpb_out[76][269],u_xpb_out[77][269],u_xpb_out[78][269],u_xpb_out[79][269],u_xpb_out[80][269],u_xpb_out[81][269],u_xpb_out[82][269],u_xpb_out[83][269],u_xpb_out[84][269],u_xpb_out[85][269],u_xpb_out[86][269],u_xpb_out[87][269],u_xpb_out[88][269],u_xpb_out[89][269],u_xpb_out[90][269],u_xpb_out[91][269],u_xpb_out[92][269],u_xpb_out[93][269],u_xpb_out[94][269],u_xpb_out[95][269],u_xpb_out[96][269],u_xpb_out[97][269],u_xpb_out[98][269],u_xpb_out[99][269],u_xpb_out[100][269],u_xpb_out[101][269],u_xpb_out[102][269],u_xpb_out[103][269],u_xpb_out[104][269],u_xpb_out[105][269]};

assign col_out_270 = {u_xpb_out[0][270],u_xpb_out[1][270],u_xpb_out[2][270],u_xpb_out[3][270],u_xpb_out[4][270],u_xpb_out[5][270],u_xpb_out[6][270],u_xpb_out[7][270],u_xpb_out[8][270],u_xpb_out[9][270],u_xpb_out[10][270],u_xpb_out[11][270],u_xpb_out[12][270],u_xpb_out[13][270],u_xpb_out[14][270],u_xpb_out[15][270],u_xpb_out[16][270],u_xpb_out[17][270],u_xpb_out[18][270],u_xpb_out[19][270],u_xpb_out[20][270],u_xpb_out[21][270],u_xpb_out[22][270],u_xpb_out[23][270],u_xpb_out[24][270],u_xpb_out[25][270],u_xpb_out[26][270],u_xpb_out[27][270],u_xpb_out[28][270],u_xpb_out[29][270],u_xpb_out[30][270],u_xpb_out[31][270],u_xpb_out[32][270],u_xpb_out[33][270],u_xpb_out[34][270],u_xpb_out[35][270],u_xpb_out[36][270],u_xpb_out[37][270],u_xpb_out[38][270],u_xpb_out[39][270],u_xpb_out[40][270],u_xpb_out[41][270],u_xpb_out[42][270],u_xpb_out[43][270],u_xpb_out[44][270],u_xpb_out[45][270],u_xpb_out[46][270],u_xpb_out[47][270],u_xpb_out[48][270],u_xpb_out[49][270],u_xpb_out[50][270],u_xpb_out[51][270],u_xpb_out[52][270],u_xpb_out[53][270],u_xpb_out[54][270],u_xpb_out[55][270],u_xpb_out[56][270],u_xpb_out[57][270],u_xpb_out[58][270],u_xpb_out[59][270],u_xpb_out[60][270],u_xpb_out[61][270],u_xpb_out[62][270],u_xpb_out[63][270],u_xpb_out[64][270],u_xpb_out[65][270],u_xpb_out[66][270],u_xpb_out[67][270],u_xpb_out[68][270],u_xpb_out[69][270],u_xpb_out[70][270],u_xpb_out[71][270],u_xpb_out[72][270],u_xpb_out[73][270],u_xpb_out[74][270],u_xpb_out[75][270],u_xpb_out[76][270],u_xpb_out[77][270],u_xpb_out[78][270],u_xpb_out[79][270],u_xpb_out[80][270],u_xpb_out[81][270],u_xpb_out[82][270],u_xpb_out[83][270],u_xpb_out[84][270],u_xpb_out[85][270],u_xpb_out[86][270],u_xpb_out[87][270],u_xpb_out[88][270],u_xpb_out[89][270],u_xpb_out[90][270],u_xpb_out[91][270],u_xpb_out[92][270],u_xpb_out[93][270],u_xpb_out[94][270],u_xpb_out[95][270],u_xpb_out[96][270],u_xpb_out[97][270],u_xpb_out[98][270],u_xpb_out[99][270],u_xpb_out[100][270],u_xpb_out[101][270],u_xpb_out[102][270],u_xpb_out[103][270],u_xpb_out[104][270],u_xpb_out[105][270]};

assign col_out_271 = {u_xpb_out[0][271],u_xpb_out[1][271],u_xpb_out[2][271],u_xpb_out[3][271],u_xpb_out[4][271],u_xpb_out[5][271],u_xpb_out[6][271],u_xpb_out[7][271],u_xpb_out[8][271],u_xpb_out[9][271],u_xpb_out[10][271],u_xpb_out[11][271],u_xpb_out[12][271],u_xpb_out[13][271],u_xpb_out[14][271],u_xpb_out[15][271],u_xpb_out[16][271],u_xpb_out[17][271],u_xpb_out[18][271],u_xpb_out[19][271],u_xpb_out[20][271],u_xpb_out[21][271],u_xpb_out[22][271],u_xpb_out[23][271],u_xpb_out[24][271],u_xpb_out[25][271],u_xpb_out[26][271],u_xpb_out[27][271],u_xpb_out[28][271],u_xpb_out[29][271],u_xpb_out[30][271],u_xpb_out[31][271],u_xpb_out[32][271],u_xpb_out[33][271],u_xpb_out[34][271],u_xpb_out[35][271],u_xpb_out[36][271],u_xpb_out[37][271],u_xpb_out[38][271],u_xpb_out[39][271],u_xpb_out[40][271],u_xpb_out[41][271],u_xpb_out[42][271],u_xpb_out[43][271],u_xpb_out[44][271],u_xpb_out[45][271],u_xpb_out[46][271],u_xpb_out[47][271],u_xpb_out[48][271],u_xpb_out[49][271],u_xpb_out[50][271],u_xpb_out[51][271],u_xpb_out[52][271],u_xpb_out[53][271],u_xpb_out[54][271],u_xpb_out[55][271],u_xpb_out[56][271],u_xpb_out[57][271],u_xpb_out[58][271],u_xpb_out[59][271],u_xpb_out[60][271],u_xpb_out[61][271],u_xpb_out[62][271],u_xpb_out[63][271],u_xpb_out[64][271],u_xpb_out[65][271],u_xpb_out[66][271],u_xpb_out[67][271],u_xpb_out[68][271],u_xpb_out[69][271],u_xpb_out[70][271],u_xpb_out[71][271],u_xpb_out[72][271],u_xpb_out[73][271],u_xpb_out[74][271],u_xpb_out[75][271],u_xpb_out[76][271],u_xpb_out[77][271],u_xpb_out[78][271],u_xpb_out[79][271],u_xpb_out[80][271],u_xpb_out[81][271],u_xpb_out[82][271],u_xpb_out[83][271],u_xpb_out[84][271],u_xpb_out[85][271],u_xpb_out[86][271],u_xpb_out[87][271],u_xpb_out[88][271],u_xpb_out[89][271],u_xpb_out[90][271],u_xpb_out[91][271],u_xpb_out[92][271],u_xpb_out[93][271],u_xpb_out[94][271],u_xpb_out[95][271],u_xpb_out[96][271],u_xpb_out[97][271],u_xpb_out[98][271],u_xpb_out[99][271],u_xpb_out[100][271],u_xpb_out[101][271],u_xpb_out[102][271],u_xpb_out[103][271],u_xpb_out[104][271],u_xpb_out[105][271]};

assign col_out_272 = {u_xpb_out[0][272],u_xpb_out[1][272],u_xpb_out[2][272],u_xpb_out[3][272],u_xpb_out[4][272],u_xpb_out[5][272],u_xpb_out[6][272],u_xpb_out[7][272],u_xpb_out[8][272],u_xpb_out[9][272],u_xpb_out[10][272],u_xpb_out[11][272],u_xpb_out[12][272],u_xpb_out[13][272],u_xpb_out[14][272],u_xpb_out[15][272],u_xpb_out[16][272],u_xpb_out[17][272],u_xpb_out[18][272],u_xpb_out[19][272],u_xpb_out[20][272],u_xpb_out[21][272],u_xpb_out[22][272],u_xpb_out[23][272],u_xpb_out[24][272],u_xpb_out[25][272],u_xpb_out[26][272],u_xpb_out[27][272],u_xpb_out[28][272],u_xpb_out[29][272],u_xpb_out[30][272],u_xpb_out[31][272],u_xpb_out[32][272],u_xpb_out[33][272],u_xpb_out[34][272],u_xpb_out[35][272],u_xpb_out[36][272],u_xpb_out[37][272],u_xpb_out[38][272],u_xpb_out[39][272],u_xpb_out[40][272],u_xpb_out[41][272],u_xpb_out[42][272],u_xpb_out[43][272],u_xpb_out[44][272],u_xpb_out[45][272],u_xpb_out[46][272],u_xpb_out[47][272],u_xpb_out[48][272],u_xpb_out[49][272],u_xpb_out[50][272],u_xpb_out[51][272],u_xpb_out[52][272],u_xpb_out[53][272],u_xpb_out[54][272],u_xpb_out[55][272],u_xpb_out[56][272],u_xpb_out[57][272],u_xpb_out[58][272],u_xpb_out[59][272],u_xpb_out[60][272],u_xpb_out[61][272],u_xpb_out[62][272],u_xpb_out[63][272],u_xpb_out[64][272],u_xpb_out[65][272],u_xpb_out[66][272],u_xpb_out[67][272],u_xpb_out[68][272],u_xpb_out[69][272],u_xpb_out[70][272],u_xpb_out[71][272],u_xpb_out[72][272],u_xpb_out[73][272],u_xpb_out[74][272],u_xpb_out[75][272],u_xpb_out[76][272],u_xpb_out[77][272],u_xpb_out[78][272],u_xpb_out[79][272],u_xpb_out[80][272],u_xpb_out[81][272],u_xpb_out[82][272],u_xpb_out[83][272],u_xpb_out[84][272],u_xpb_out[85][272],u_xpb_out[86][272],u_xpb_out[87][272],u_xpb_out[88][272],u_xpb_out[89][272],u_xpb_out[90][272],u_xpb_out[91][272],u_xpb_out[92][272],u_xpb_out[93][272],u_xpb_out[94][272],u_xpb_out[95][272],u_xpb_out[96][272],u_xpb_out[97][272],u_xpb_out[98][272],u_xpb_out[99][272],u_xpb_out[100][272],u_xpb_out[101][272],u_xpb_out[102][272],u_xpb_out[103][272],u_xpb_out[104][272],u_xpb_out[105][272]};

assign col_out_273 = {u_xpb_out[0][273],u_xpb_out[1][273],u_xpb_out[2][273],u_xpb_out[3][273],u_xpb_out[4][273],u_xpb_out[5][273],u_xpb_out[6][273],u_xpb_out[7][273],u_xpb_out[8][273],u_xpb_out[9][273],u_xpb_out[10][273],u_xpb_out[11][273],u_xpb_out[12][273],u_xpb_out[13][273],u_xpb_out[14][273],u_xpb_out[15][273],u_xpb_out[16][273],u_xpb_out[17][273],u_xpb_out[18][273],u_xpb_out[19][273],u_xpb_out[20][273],u_xpb_out[21][273],u_xpb_out[22][273],u_xpb_out[23][273],u_xpb_out[24][273],u_xpb_out[25][273],u_xpb_out[26][273],u_xpb_out[27][273],u_xpb_out[28][273],u_xpb_out[29][273],u_xpb_out[30][273],u_xpb_out[31][273],u_xpb_out[32][273],u_xpb_out[33][273],u_xpb_out[34][273],u_xpb_out[35][273],u_xpb_out[36][273],u_xpb_out[37][273],u_xpb_out[38][273],u_xpb_out[39][273],u_xpb_out[40][273],u_xpb_out[41][273],u_xpb_out[42][273],u_xpb_out[43][273],u_xpb_out[44][273],u_xpb_out[45][273],u_xpb_out[46][273],u_xpb_out[47][273],u_xpb_out[48][273],u_xpb_out[49][273],u_xpb_out[50][273],u_xpb_out[51][273],u_xpb_out[52][273],u_xpb_out[53][273],u_xpb_out[54][273],u_xpb_out[55][273],u_xpb_out[56][273],u_xpb_out[57][273],u_xpb_out[58][273],u_xpb_out[59][273],u_xpb_out[60][273],u_xpb_out[61][273],u_xpb_out[62][273],u_xpb_out[63][273],u_xpb_out[64][273],u_xpb_out[65][273],u_xpb_out[66][273],u_xpb_out[67][273],u_xpb_out[68][273],u_xpb_out[69][273],u_xpb_out[70][273],u_xpb_out[71][273],u_xpb_out[72][273],u_xpb_out[73][273],u_xpb_out[74][273],u_xpb_out[75][273],u_xpb_out[76][273],u_xpb_out[77][273],u_xpb_out[78][273],u_xpb_out[79][273],u_xpb_out[80][273],u_xpb_out[81][273],u_xpb_out[82][273],u_xpb_out[83][273],u_xpb_out[84][273],u_xpb_out[85][273],u_xpb_out[86][273],u_xpb_out[87][273],u_xpb_out[88][273],u_xpb_out[89][273],u_xpb_out[90][273],u_xpb_out[91][273],u_xpb_out[92][273],u_xpb_out[93][273],u_xpb_out[94][273],u_xpb_out[95][273],u_xpb_out[96][273],u_xpb_out[97][273],u_xpb_out[98][273],u_xpb_out[99][273],u_xpb_out[100][273],u_xpb_out[101][273],u_xpb_out[102][273],u_xpb_out[103][273],u_xpb_out[104][273],u_xpb_out[105][273]};

assign col_out_274 = {u_xpb_out[0][274],u_xpb_out[1][274],u_xpb_out[2][274],u_xpb_out[3][274],u_xpb_out[4][274],u_xpb_out[5][274],u_xpb_out[6][274],u_xpb_out[7][274],u_xpb_out[8][274],u_xpb_out[9][274],u_xpb_out[10][274],u_xpb_out[11][274],u_xpb_out[12][274],u_xpb_out[13][274],u_xpb_out[14][274],u_xpb_out[15][274],u_xpb_out[16][274],u_xpb_out[17][274],u_xpb_out[18][274],u_xpb_out[19][274],u_xpb_out[20][274],u_xpb_out[21][274],u_xpb_out[22][274],u_xpb_out[23][274],u_xpb_out[24][274],u_xpb_out[25][274],u_xpb_out[26][274],u_xpb_out[27][274],u_xpb_out[28][274],u_xpb_out[29][274],u_xpb_out[30][274],u_xpb_out[31][274],u_xpb_out[32][274],u_xpb_out[33][274],u_xpb_out[34][274],u_xpb_out[35][274],u_xpb_out[36][274],u_xpb_out[37][274],u_xpb_out[38][274],u_xpb_out[39][274],u_xpb_out[40][274],u_xpb_out[41][274],u_xpb_out[42][274],u_xpb_out[43][274],u_xpb_out[44][274],u_xpb_out[45][274],u_xpb_out[46][274],u_xpb_out[47][274],u_xpb_out[48][274],u_xpb_out[49][274],u_xpb_out[50][274],u_xpb_out[51][274],u_xpb_out[52][274],u_xpb_out[53][274],u_xpb_out[54][274],u_xpb_out[55][274],u_xpb_out[56][274],u_xpb_out[57][274],u_xpb_out[58][274],u_xpb_out[59][274],u_xpb_out[60][274],u_xpb_out[61][274],u_xpb_out[62][274],u_xpb_out[63][274],u_xpb_out[64][274],u_xpb_out[65][274],u_xpb_out[66][274],u_xpb_out[67][274],u_xpb_out[68][274],u_xpb_out[69][274],u_xpb_out[70][274],u_xpb_out[71][274],u_xpb_out[72][274],u_xpb_out[73][274],u_xpb_out[74][274],u_xpb_out[75][274],u_xpb_out[76][274],u_xpb_out[77][274],u_xpb_out[78][274],u_xpb_out[79][274],u_xpb_out[80][274],u_xpb_out[81][274],u_xpb_out[82][274],u_xpb_out[83][274],u_xpb_out[84][274],u_xpb_out[85][274],u_xpb_out[86][274],u_xpb_out[87][274],u_xpb_out[88][274],u_xpb_out[89][274],u_xpb_out[90][274],u_xpb_out[91][274],u_xpb_out[92][274],u_xpb_out[93][274],u_xpb_out[94][274],u_xpb_out[95][274],u_xpb_out[96][274],u_xpb_out[97][274],u_xpb_out[98][274],u_xpb_out[99][274],u_xpb_out[100][274],u_xpb_out[101][274],u_xpb_out[102][274],u_xpb_out[103][274],u_xpb_out[104][274],u_xpb_out[105][274]};

assign col_out_275 = {u_xpb_out[0][275],u_xpb_out[1][275],u_xpb_out[2][275],u_xpb_out[3][275],u_xpb_out[4][275],u_xpb_out[5][275],u_xpb_out[6][275],u_xpb_out[7][275],u_xpb_out[8][275],u_xpb_out[9][275],u_xpb_out[10][275],u_xpb_out[11][275],u_xpb_out[12][275],u_xpb_out[13][275],u_xpb_out[14][275],u_xpb_out[15][275],u_xpb_out[16][275],u_xpb_out[17][275],u_xpb_out[18][275],u_xpb_out[19][275],u_xpb_out[20][275],u_xpb_out[21][275],u_xpb_out[22][275],u_xpb_out[23][275],u_xpb_out[24][275],u_xpb_out[25][275],u_xpb_out[26][275],u_xpb_out[27][275],u_xpb_out[28][275],u_xpb_out[29][275],u_xpb_out[30][275],u_xpb_out[31][275],u_xpb_out[32][275],u_xpb_out[33][275],u_xpb_out[34][275],u_xpb_out[35][275],u_xpb_out[36][275],u_xpb_out[37][275],u_xpb_out[38][275],u_xpb_out[39][275],u_xpb_out[40][275],u_xpb_out[41][275],u_xpb_out[42][275],u_xpb_out[43][275],u_xpb_out[44][275],u_xpb_out[45][275],u_xpb_out[46][275],u_xpb_out[47][275],u_xpb_out[48][275],u_xpb_out[49][275],u_xpb_out[50][275],u_xpb_out[51][275],u_xpb_out[52][275],u_xpb_out[53][275],u_xpb_out[54][275],u_xpb_out[55][275],u_xpb_out[56][275],u_xpb_out[57][275],u_xpb_out[58][275],u_xpb_out[59][275],u_xpb_out[60][275],u_xpb_out[61][275],u_xpb_out[62][275],u_xpb_out[63][275],u_xpb_out[64][275],u_xpb_out[65][275],u_xpb_out[66][275],u_xpb_out[67][275],u_xpb_out[68][275],u_xpb_out[69][275],u_xpb_out[70][275],u_xpb_out[71][275],u_xpb_out[72][275],u_xpb_out[73][275],u_xpb_out[74][275],u_xpb_out[75][275],u_xpb_out[76][275],u_xpb_out[77][275],u_xpb_out[78][275],u_xpb_out[79][275],u_xpb_out[80][275],u_xpb_out[81][275],u_xpb_out[82][275],u_xpb_out[83][275],u_xpb_out[84][275],u_xpb_out[85][275],u_xpb_out[86][275],u_xpb_out[87][275],u_xpb_out[88][275],u_xpb_out[89][275],u_xpb_out[90][275],u_xpb_out[91][275],u_xpb_out[92][275],u_xpb_out[93][275],u_xpb_out[94][275],u_xpb_out[95][275],u_xpb_out[96][275],u_xpb_out[97][275],u_xpb_out[98][275],u_xpb_out[99][275],u_xpb_out[100][275],u_xpb_out[101][275],u_xpb_out[102][275],u_xpb_out[103][275],u_xpb_out[104][275],u_xpb_out[105][275]};

assign col_out_276 = {u_xpb_out[0][276],u_xpb_out[1][276],u_xpb_out[2][276],u_xpb_out[3][276],u_xpb_out[4][276],u_xpb_out[5][276],u_xpb_out[6][276],u_xpb_out[7][276],u_xpb_out[8][276],u_xpb_out[9][276],u_xpb_out[10][276],u_xpb_out[11][276],u_xpb_out[12][276],u_xpb_out[13][276],u_xpb_out[14][276],u_xpb_out[15][276],u_xpb_out[16][276],u_xpb_out[17][276],u_xpb_out[18][276],u_xpb_out[19][276],u_xpb_out[20][276],u_xpb_out[21][276],u_xpb_out[22][276],u_xpb_out[23][276],u_xpb_out[24][276],u_xpb_out[25][276],u_xpb_out[26][276],u_xpb_out[27][276],u_xpb_out[28][276],u_xpb_out[29][276],u_xpb_out[30][276],u_xpb_out[31][276],u_xpb_out[32][276],u_xpb_out[33][276],u_xpb_out[34][276],u_xpb_out[35][276],u_xpb_out[36][276],u_xpb_out[37][276],u_xpb_out[38][276],u_xpb_out[39][276],u_xpb_out[40][276],u_xpb_out[41][276],u_xpb_out[42][276],u_xpb_out[43][276],u_xpb_out[44][276],u_xpb_out[45][276],u_xpb_out[46][276],u_xpb_out[47][276],u_xpb_out[48][276],u_xpb_out[49][276],u_xpb_out[50][276],u_xpb_out[51][276],u_xpb_out[52][276],u_xpb_out[53][276],u_xpb_out[54][276],u_xpb_out[55][276],u_xpb_out[56][276],u_xpb_out[57][276],u_xpb_out[58][276],u_xpb_out[59][276],u_xpb_out[60][276],u_xpb_out[61][276],u_xpb_out[62][276],u_xpb_out[63][276],u_xpb_out[64][276],u_xpb_out[65][276],u_xpb_out[66][276],u_xpb_out[67][276],u_xpb_out[68][276],u_xpb_out[69][276],u_xpb_out[70][276],u_xpb_out[71][276],u_xpb_out[72][276],u_xpb_out[73][276],u_xpb_out[74][276],u_xpb_out[75][276],u_xpb_out[76][276],u_xpb_out[77][276],u_xpb_out[78][276],u_xpb_out[79][276],u_xpb_out[80][276],u_xpb_out[81][276],u_xpb_out[82][276],u_xpb_out[83][276],u_xpb_out[84][276],u_xpb_out[85][276],u_xpb_out[86][276],u_xpb_out[87][276],u_xpb_out[88][276],u_xpb_out[89][276],u_xpb_out[90][276],u_xpb_out[91][276],u_xpb_out[92][276],u_xpb_out[93][276],u_xpb_out[94][276],u_xpb_out[95][276],u_xpb_out[96][276],u_xpb_out[97][276],u_xpb_out[98][276],u_xpb_out[99][276],u_xpb_out[100][276],u_xpb_out[101][276],u_xpb_out[102][276],u_xpb_out[103][276],u_xpb_out[104][276],u_xpb_out[105][276]};

assign col_out_277 = {u_xpb_out[0][277],u_xpb_out[1][277],u_xpb_out[2][277],u_xpb_out[3][277],u_xpb_out[4][277],u_xpb_out[5][277],u_xpb_out[6][277],u_xpb_out[7][277],u_xpb_out[8][277],u_xpb_out[9][277],u_xpb_out[10][277],u_xpb_out[11][277],u_xpb_out[12][277],u_xpb_out[13][277],u_xpb_out[14][277],u_xpb_out[15][277],u_xpb_out[16][277],u_xpb_out[17][277],u_xpb_out[18][277],u_xpb_out[19][277],u_xpb_out[20][277],u_xpb_out[21][277],u_xpb_out[22][277],u_xpb_out[23][277],u_xpb_out[24][277],u_xpb_out[25][277],u_xpb_out[26][277],u_xpb_out[27][277],u_xpb_out[28][277],u_xpb_out[29][277],u_xpb_out[30][277],u_xpb_out[31][277],u_xpb_out[32][277],u_xpb_out[33][277],u_xpb_out[34][277],u_xpb_out[35][277],u_xpb_out[36][277],u_xpb_out[37][277],u_xpb_out[38][277],u_xpb_out[39][277],u_xpb_out[40][277],u_xpb_out[41][277],u_xpb_out[42][277],u_xpb_out[43][277],u_xpb_out[44][277],u_xpb_out[45][277],u_xpb_out[46][277],u_xpb_out[47][277],u_xpb_out[48][277],u_xpb_out[49][277],u_xpb_out[50][277],u_xpb_out[51][277],u_xpb_out[52][277],u_xpb_out[53][277],u_xpb_out[54][277],u_xpb_out[55][277],u_xpb_out[56][277],u_xpb_out[57][277],u_xpb_out[58][277],u_xpb_out[59][277],u_xpb_out[60][277],u_xpb_out[61][277],u_xpb_out[62][277],u_xpb_out[63][277],u_xpb_out[64][277],u_xpb_out[65][277],u_xpb_out[66][277],u_xpb_out[67][277],u_xpb_out[68][277],u_xpb_out[69][277],u_xpb_out[70][277],u_xpb_out[71][277],u_xpb_out[72][277],u_xpb_out[73][277],u_xpb_out[74][277],u_xpb_out[75][277],u_xpb_out[76][277],u_xpb_out[77][277],u_xpb_out[78][277],u_xpb_out[79][277],u_xpb_out[80][277],u_xpb_out[81][277],u_xpb_out[82][277],u_xpb_out[83][277],u_xpb_out[84][277],u_xpb_out[85][277],u_xpb_out[86][277],u_xpb_out[87][277],u_xpb_out[88][277],u_xpb_out[89][277],u_xpb_out[90][277],u_xpb_out[91][277],u_xpb_out[92][277],u_xpb_out[93][277],u_xpb_out[94][277],u_xpb_out[95][277],u_xpb_out[96][277],u_xpb_out[97][277],u_xpb_out[98][277],u_xpb_out[99][277],u_xpb_out[100][277],u_xpb_out[101][277],u_xpb_out[102][277],u_xpb_out[103][277],u_xpb_out[104][277],u_xpb_out[105][277]};

assign col_out_278 = {u_xpb_out[0][278],u_xpb_out[1][278],u_xpb_out[2][278],u_xpb_out[3][278],u_xpb_out[4][278],u_xpb_out[5][278],u_xpb_out[6][278],u_xpb_out[7][278],u_xpb_out[8][278],u_xpb_out[9][278],u_xpb_out[10][278],u_xpb_out[11][278],u_xpb_out[12][278],u_xpb_out[13][278],u_xpb_out[14][278],u_xpb_out[15][278],u_xpb_out[16][278],u_xpb_out[17][278],u_xpb_out[18][278],u_xpb_out[19][278],u_xpb_out[20][278],u_xpb_out[21][278],u_xpb_out[22][278],u_xpb_out[23][278],u_xpb_out[24][278],u_xpb_out[25][278],u_xpb_out[26][278],u_xpb_out[27][278],u_xpb_out[28][278],u_xpb_out[29][278],u_xpb_out[30][278],u_xpb_out[31][278],u_xpb_out[32][278],u_xpb_out[33][278],u_xpb_out[34][278],u_xpb_out[35][278],u_xpb_out[36][278],u_xpb_out[37][278],u_xpb_out[38][278],u_xpb_out[39][278],u_xpb_out[40][278],u_xpb_out[41][278],u_xpb_out[42][278],u_xpb_out[43][278],u_xpb_out[44][278],u_xpb_out[45][278],u_xpb_out[46][278],u_xpb_out[47][278],u_xpb_out[48][278],u_xpb_out[49][278],u_xpb_out[50][278],u_xpb_out[51][278],u_xpb_out[52][278],u_xpb_out[53][278],u_xpb_out[54][278],u_xpb_out[55][278],u_xpb_out[56][278],u_xpb_out[57][278],u_xpb_out[58][278],u_xpb_out[59][278],u_xpb_out[60][278],u_xpb_out[61][278],u_xpb_out[62][278],u_xpb_out[63][278],u_xpb_out[64][278],u_xpb_out[65][278],u_xpb_out[66][278],u_xpb_out[67][278],u_xpb_out[68][278],u_xpb_out[69][278],u_xpb_out[70][278],u_xpb_out[71][278],u_xpb_out[72][278],u_xpb_out[73][278],u_xpb_out[74][278],u_xpb_out[75][278],u_xpb_out[76][278],u_xpb_out[77][278],u_xpb_out[78][278],u_xpb_out[79][278],u_xpb_out[80][278],u_xpb_out[81][278],u_xpb_out[82][278],u_xpb_out[83][278],u_xpb_out[84][278],u_xpb_out[85][278],u_xpb_out[86][278],u_xpb_out[87][278],u_xpb_out[88][278],u_xpb_out[89][278],u_xpb_out[90][278],u_xpb_out[91][278],u_xpb_out[92][278],u_xpb_out[93][278],u_xpb_out[94][278],u_xpb_out[95][278],u_xpb_out[96][278],u_xpb_out[97][278],u_xpb_out[98][278],u_xpb_out[99][278],u_xpb_out[100][278],u_xpb_out[101][278],u_xpb_out[102][278],u_xpb_out[103][278],u_xpb_out[104][278],u_xpb_out[105][278]};

assign col_out_279 = {u_xpb_out[0][279],u_xpb_out[1][279],u_xpb_out[2][279],u_xpb_out[3][279],u_xpb_out[4][279],u_xpb_out[5][279],u_xpb_out[6][279],u_xpb_out[7][279],u_xpb_out[8][279],u_xpb_out[9][279],u_xpb_out[10][279],u_xpb_out[11][279],u_xpb_out[12][279],u_xpb_out[13][279],u_xpb_out[14][279],u_xpb_out[15][279],u_xpb_out[16][279],u_xpb_out[17][279],u_xpb_out[18][279],u_xpb_out[19][279],u_xpb_out[20][279],u_xpb_out[21][279],u_xpb_out[22][279],u_xpb_out[23][279],u_xpb_out[24][279],u_xpb_out[25][279],u_xpb_out[26][279],u_xpb_out[27][279],u_xpb_out[28][279],u_xpb_out[29][279],u_xpb_out[30][279],u_xpb_out[31][279],u_xpb_out[32][279],u_xpb_out[33][279],u_xpb_out[34][279],u_xpb_out[35][279],u_xpb_out[36][279],u_xpb_out[37][279],u_xpb_out[38][279],u_xpb_out[39][279],u_xpb_out[40][279],u_xpb_out[41][279],u_xpb_out[42][279],u_xpb_out[43][279],u_xpb_out[44][279],u_xpb_out[45][279],u_xpb_out[46][279],u_xpb_out[47][279],u_xpb_out[48][279],u_xpb_out[49][279],u_xpb_out[50][279],u_xpb_out[51][279],u_xpb_out[52][279],u_xpb_out[53][279],u_xpb_out[54][279],u_xpb_out[55][279],u_xpb_out[56][279],u_xpb_out[57][279],u_xpb_out[58][279],u_xpb_out[59][279],u_xpb_out[60][279],u_xpb_out[61][279],u_xpb_out[62][279],u_xpb_out[63][279],u_xpb_out[64][279],u_xpb_out[65][279],u_xpb_out[66][279],u_xpb_out[67][279],u_xpb_out[68][279],u_xpb_out[69][279],u_xpb_out[70][279],u_xpb_out[71][279],u_xpb_out[72][279],u_xpb_out[73][279],u_xpb_out[74][279],u_xpb_out[75][279],u_xpb_out[76][279],u_xpb_out[77][279],u_xpb_out[78][279],u_xpb_out[79][279],u_xpb_out[80][279],u_xpb_out[81][279],u_xpb_out[82][279],u_xpb_out[83][279],u_xpb_out[84][279],u_xpb_out[85][279],u_xpb_out[86][279],u_xpb_out[87][279],u_xpb_out[88][279],u_xpb_out[89][279],u_xpb_out[90][279],u_xpb_out[91][279],u_xpb_out[92][279],u_xpb_out[93][279],u_xpb_out[94][279],u_xpb_out[95][279],u_xpb_out[96][279],u_xpb_out[97][279],u_xpb_out[98][279],u_xpb_out[99][279],u_xpb_out[100][279],u_xpb_out[101][279],u_xpb_out[102][279],u_xpb_out[103][279],u_xpb_out[104][279],u_xpb_out[105][279]};

assign col_out_280 = {u_xpb_out[0][280],u_xpb_out[1][280],u_xpb_out[2][280],u_xpb_out[3][280],u_xpb_out[4][280],u_xpb_out[5][280],u_xpb_out[6][280],u_xpb_out[7][280],u_xpb_out[8][280],u_xpb_out[9][280],u_xpb_out[10][280],u_xpb_out[11][280],u_xpb_out[12][280],u_xpb_out[13][280],u_xpb_out[14][280],u_xpb_out[15][280],u_xpb_out[16][280],u_xpb_out[17][280],u_xpb_out[18][280],u_xpb_out[19][280],u_xpb_out[20][280],u_xpb_out[21][280],u_xpb_out[22][280],u_xpb_out[23][280],u_xpb_out[24][280],u_xpb_out[25][280],u_xpb_out[26][280],u_xpb_out[27][280],u_xpb_out[28][280],u_xpb_out[29][280],u_xpb_out[30][280],u_xpb_out[31][280],u_xpb_out[32][280],u_xpb_out[33][280],u_xpb_out[34][280],u_xpb_out[35][280],u_xpb_out[36][280],u_xpb_out[37][280],u_xpb_out[38][280],u_xpb_out[39][280],u_xpb_out[40][280],u_xpb_out[41][280],u_xpb_out[42][280],u_xpb_out[43][280],u_xpb_out[44][280],u_xpb_out[45][280],u_xpb_out[46][280],u_xpb_out[47][280],u_xpb_out[48][280],u_xpb_out[49][280],u_xpb_out[50][280],u_xpb_out[51][280],u_xpb_out[52][280],u_xpb_out[53][280],u_xpb_out[54][280],u_xpb_out[55][280],u_xpb_out[56][280],u_xpb_out[57][280],u_xpb_out[58][280],u_xpb_out[59][280],u_xpb_out[60][280],u_xpb_out[61][280],u_xpb_out[62][280],u_xpb_out[63][280],u_xpb_out[64][280],u_xpb_out[65][280],u_xpb_out[66][280],u_xpb_out[67][280],u_xpb_out[68][280],u_xpb_out[69][280],u_xpb_out[70][280],u_xpb_out[71][280],u_xpb_out[72][280],u_xpb_out[73][280],u_xpb_out[74][280],u_xpb_out[75][280],u_xpb_out[76][280],u_xpb_out[77][280],u_xpb_out[78][280],u_xpb_out[79][280],u_xpb_out[80][280],u_xpb_out[81][280],u_xpb_out[82][280],u_xpb_out[83][280],u_xpb_out[84][280],u_xpb_out[85][280],u_xpb_out[86][280],u_xpb_out[87][280],u_xpb_out[88][280],u_xpb_out[89][280],u_xpb_out[90][280],u_xpb_out[91][280],u_xpb_out[92][280],u_xpb_out[93][280],u_xpb_out[94][280],u_xpb_out[95][280],u_xpb_out[96][280],u_xpb_out[97][280],u_xpb_out[98][280],u_xpb_out[99][280],u_xpb_out[100][280],u_xpb_out[101][280],u_xpb_out[102][280],u_xpb_out[103][280],u_xpb_out[104][280],u_xpb_out[105][280]};

assign col_out_281 = {u_xpb_out[0][281],u_xpb_out[1][281],u_xpb_out[2][281],u_xpb_out[3][281],u_xpb_out[4][281],u_xpb_out[5][281],u_xpb_out[6][281],u_xpb_out[7][281],u_xpb_out[8][281],u_xpb_out[9][281],u_xpb_out[10][281],u_xpb_out[11][281],u_xpb_out[12][281],u_xpb_out[13][281],u_xpb_out[14][281],u_xpb_out[15][281],u_xpb_out[16][281],u_xpb_out[17][281],u_xpb_out[18][281],u_xpb_out[19][281],u_xpb_out[20][281],u_xpb_out[21][281],u_xpb_out[22][281],u_xpb_out[23][281],u_xpb_out[24][281],u_xpb_out[25][281],u_xpb_out[26][281],u_xpb_out[27][281],u_xpb_out[28][281],u_xpb_out[29][281],u_xpb_out[30][281],u_xpb_out[31][281],u_xpb_out[32][281],u_xpb_out[33][281],u_xpb_out[34][281],u_xpb_out[35][281],u_xpb_out[36][281],u_xpb_out[37][281],u_xpb_out[38][281],u_xpb_out[39][281],u_xpb_out[40][281],u_xpb_out[41][281],u_xpb_out[42][281],u_xpb_out[43][281],u_xpb_out[44][281],u_xpb_out[45][281],u_xpb_out[46][281],u_xpb_out[47][281],u_xpb_out[48][281],u_xpb_out[49][281],u_xpb_out[50][281],u_xpb_out[51][281],u_xpb_out[52][281],u_xpb_out[53][281],u_xpb_out[54][281],u_xpb_out[55][281],u_xpb_out[56][281],u_xpb_out[57][281],u_xpb_out[58][281],u_xpb_out[59][281],u_xpb_out[60][281],u_xpb_out[61][281],u_xpb_out[62][281],u_xpb_out[63][281],u_xpb_out[64][281],u_xpb_out[65][281],u_xpb_out[66][281],u_xpb_out[67][281],u_xpb_out[68][281],u_xpb_out[69][281],u_xpb_out[70][281],u_xpb_out[71][281],u_xpb_out[72][281],u_xpb_out[73][281],u_xpb_out[74][281],u_xpb_out[75][281],u_xpb_out[76][281],u_xpb_out[77][281],u_xpb_out[78][281],u_xpb_out[79][281],u_xpb_out[80][281],u_xpb_out[81][281],u_xpb_out[82][281],u_xpb_out[83][281],u_xpb_out[84][281],u_xpb_out[85][281],u_xpb_out[86][281],u_xpb_out[87][281],u_xpb_out[88][281],u_xpb_out[89][281],u_xpb_out[90][281],u_xpb_out[91][281],u_xpb_out[92][281],u_xpb_out[93][281],u_xpb_out[94][281],u_xpb_out[95][281],u_xpb_out[96][281],u_xpb_out[97][281],u_xpb_out[98][281],u_xpb_out[99][281],u_xpb_out[100][281],u_xpb_out[101][281],u_xpb_out[102][281],u_xpb_out[103][281],u_xpb_out[104][281],u_xpb_out[105][281]};

assign col_out_282 = {u_xpb_out[0][282],u_xpb_out[1][282],u_xpb_out[2][282],u_xpb_out[3][282],u_xpb_out[4][282],u_xpb_out[5][282],u_xpb_out[6][282],u_xpb_out[7][282],u_xpb_out[8][282],u_xpb_out[9][282],u_xpb_out[10][282],u_xpb_out[11][282],u_xpb_out[12][282],u_xpb_out[13][282],u_xpb_out[14][282],u_xpb_out[15][282],u_xpb_out[16][282],u_xpb_out[17][282],u_xpb_out[18][282],u_xpb_out[19][282],u_xpb_out[20][282],u_xpb_out[21][282],u_xpb_out[22][282],u_xpb_out[23][282],u_xpb_out[24][282],u_xpb_out[25][282],u_xpb_out[26][282],u_xpb_out[27][282],u_xpb_out[28][282],u_xpb_out[29][282],u_xpb_out[30][282],u_xpb_out[31][282],u_xpb_out[32][282],u_xpb_out[33][282],u_xpb_out[34][282],u_xpb_out[35][282],u_xpb_out[36][282],u_xpb_out[37][282],u_xpb_out[38][282],u_xpb_out[39][282],u_xpb_out[40][282],u_xpb_out[41][282],u_xpb_out[42][282],u_xpb_out[43][282],u_xpb_out[44][282],u_xpb_out[45][282],u_xpb_out[46][282],u_xpb_out[47][282],u_xpb_out[48][282],u_xpb_out[49][282],u_xpb_out[50][282],u_xpb_out[51][282],u_xpb_out[52][282],u_xpb_out[53][282],u_xpb_out[54][282],u_xpb_out[55][282],u_xpb_out[56][282],u_xpb_out[57][282],u_xpb_out[58][282],u_xpb_out[59][282],u_xpb_out[60][282],u_xpb_out[61][282],u_xpb_out[62][282],u_xpb_out[63][282],u_xpb_out[64][282],u_xpb_out[65][282],u_xpb_out[66][282],u_xpb_out[67][282],u_xpb_out[68][282],u_xpb_out[69][282],u_xpb_out[70][282],u_xpb_out[71][282],u_xpb_out[72][282],u_xpb_out[73][282],u_xpb_out[74][282],u_xpb_out[75][282],u_xpb_out[76][282],u_xpb_out[77][282],u_xpb_out[78][282],u_xpb_out[79][282],u_xpb_out[80][282],u_xpb_out[81][282],u_xpb_out[82][282],u_xpb_out[83][282],u_xpb_out[84][282],u_xpb_out[85][282],u_xpb_out[86][282],u_xpb_out[87][282],u_xpb_out[88][282],u_xpb_out[89][282],u_xpb_out[90][282],u_xpb_out[91][282],u_xpb_out[92][282],u_xpb_out[93][282],u_xpb_out[94][282],u_xpb_out[95][282],u_xpb_out[96][282],u_xpb_out[97][282],u_xpb_out[98][282],u_xpb_out[99][282],u_xpb_out[100][282],u_xpb_out[101][282],u_xpb_out[102][282],u_xpb_out[103][282],u_xpb_out[104][282],u_xpb_out[105][282]};

assign col_out_283 = {u_xpb_out[0][283],u_xpb_out[1][283],u_xpb_out[2][283],u_xpb_out[3][283],u_xpb_out[4][283],u_xpb_out[5][283],u_xpb_out[6][283],u_xpb_out[7][283],u_xpb_out[8][283],u_xpb_out[9][283],u_xpb_out[10][283],u_xpb_out[11][283],u_xpb_out[12][283],u_xpb_out[13][283],u_xpb_out[14][283],u_xpb_out[15][283],u_xpb_out[16][283],u_xpb_out[17][283],u_xpb_out[18][283],u_xpb_out[19][283],u_xpb_out[20][283],u_xpb_out[21][283],u_xpb_out[22][283],u_xpb_out[23][283],u_xpb_out[24][283],u_xpb_out[25][283],u_xpb_out[26][283],u_xpb_out[27][283],u_xpb_out[28][283],u_xpb_out[29][283],u_xpb_out[30][283],u_xpb_out[31][283],u_xpb_out[32][283],u_xpb_out[33][283],u_xpb_out[34][283],u_xpb_out[35][283],u_xpb_out[36][283],u_xpb_out[37][283],u_xpb_out[38][283],u_xpb_out[39][283],u_xpb_out[40][283],u_xpb_out[41][283],u_xpb_out[42][283],u_xpb_out[43][283],u_xpb_out[44][283],u_xpb_out[45][283],u_xpb_out[46][283],u_xpb_out[47][283],u_xpb_out[48][283],u_xpb_out[49][283],u_xpb_out[50][283],u_xpb_out[51][283],u_xpb_out[52][283],u_xpb_out[53][283],u_xpb_out[54][283],u_xpb_out[55][283],u_xpb_out[56][283],u_xpb_out[57][283],u_xpb_out[58][283],u_xpb_out[59][283],u_xpb_out[60][283],u_xpb_out[61][283],u_xpb_out[62][283],u_xpb_out[63][283],u_xpb_out[64][283],u_xpb_out[65][283],u_xpb_out[66][283],u_xpb_out[67][283],u_xpb_out[68][283],u_xpb_out[69][283],u_xpb_out[70][283],u_xpb_out[71][283],u_xpb_out[72][283],u_xpb_out[73][283],u_xpb_out[74][283],u_xpb_out[75][283],u_xpb_out[76][283],u_xpb_out[77][283],u_xpb_out[78][283],u_xpb_out[79][283],u_xpb_out[80][283],u_xpb_out[81][283],u_xpb_out[82][283],u_xpb_out[83][283],u_xpb_out[84][283],u_xpb_out[85][283],u_xpb_out[86][283],u_xpb_out[87][283],u_xpb_out[88][283],u_xpb_out[89][283],u_xpb_out[90][283],u_xpb_out[91][283],u_xpb_out[92][283],u_xpb_out[93][283],u_xpb_out[94][283],u_xpb_out[95][283],u_xpb_out[96][283],u_xpb_out[97][283],u_xpb_out[98][283],u_xpb_out[99][283],u_xpb_out[100][283],u_xpb_out[101][283],u_xpb_out[102][283],u_xpb_out[103][283],u_xpb_out[104][283],u_xpb_out[105][283]};

assign col_out_284 = {u_xpb_out[0][284],u_xpb_out[1][284],u_xpb_out[2][284],u_xpb_out[3][284],u_xpb_out[4][284],u_xpb_out[5][284],u_xpb_out[6][284],u_xpb_out[7][284],u_xpb_out[8][284],u_xpb_out[9][284],u_xpb_out[10][284],u_xpb_out[11][284],u_xpb_out[12][284],u_xpb_out[13][284],u_xpb_out[14][284],u_xpb_out[15][284],u_xpb_out[16][284],u_xpb_out[17][284],u_xpb_out[18][284],u_xpb_out[19][284],u_xpb_out[20][284],u_xpb_out[21][284],u_xpb_out[22][284],u_xpb_out[23][284],u_xpb_out[24][284],u_xpb_out[25][284],u_xpb_out[26][284],u_xpb_out[27][284],u_xpb_out[28][284],u_xpb_out[29][284],u_xpb_out[30][284],u_xpb_out[31][284],u_xpb_out[32][284],u_xpb_out[33][284],u_xpb_out[34][284],u_xpb_out[35][284],u_xpb_out[36][284],u_xpb_out[37][284],u_xpb_out[38][284],u_xpb_out[39][284],u_xpb_out[40][284],u_xpb_out[41][284],u_xpb_out[42][284],u_xpb_out[43][284],u_xpb_out[44][284],u_xpb_out[45][284],u_xpb_out[46][284],u_xpb_out[47][284],u_xpb_out[48][284],u_xpb_out[49][284],u_xpb_out[50][284],u_xpb_out[51][284],u_xpb_out[52][284],u_xpb_out[53][284],u_xpb_out[54][284],u_xpb_out[55][284],u_xpb_out[56][284],u_xpb_out[57][284],u_xpb_out[58][284],u_xpb_out[59][284],u_xpb_out[60][284],u_xpb_out[61][284],u_xpb_out[62][284],u_xpb_out[63][284],u_xpb_out[64][284],u_xpb_out[65][284],u_xpb_out[66][284],u_xpb_out[67][284],u_xpb_out[68][284],u_xpb_out[69][284],u_xpb_out[70][284],u_xpb_out[71][284],u_xpb_out[72][284],u_xpb_out[73][284],u_xpb_out[74][284],u_xpb_out[75][284],u_xpb_out[76][284],u_xpb_out[77][284],u_xpb_out[78][284],u_xpb_out[79][284],u_xpb_out[80][284],u_xpb_out[81][284],u_xpb_out[82][284],u_xpb_out[83][284],u_xpb_out[84][284],u_xpb_out[85][284],u_xpb_out[86][284],u_xpb_out[87][284],u_xpb_out[88][284],u_xpb_out[89][284],u_xpb_out[90][284],u_xpb_out[91][284],u_xpb_out[92][284],u_xpb_out[93][284],u_xpb_out[94][284],u_xpb_out[95][284],u_xpb_out[96][284],u_xpb_out[97][284],u_xpb_out[98][284],u_xpb_out[99][284],u_xpb_out[100][284],u_xpb_out[101][284],u_xpb_out[102][284],u_xpb_out[103][284],u_xpb_out[104][284],u_xpb_out[105][284]};

assign col_out_285 = {u_xpb_out[0][285],u_xpb_out[1][285],u_xpb_out[2][285],u_xpb_out[3][285],u_xpb_out[4][285],u_xpb_out[5][285],u_xpb_out[6][285],u_xpb_out[7][285],u_xpb_out[8][285],u_xpb_out[9][285],u_xpb_out[10][285],u_xpb_out[11][285],u_xpb_out[12][285],u_xpb_out[13][285],u_xpb_out[14][285],u_xpb_out[15][285],u_xpb_out[16][285],u_xpb_out[17][285],u_xpb_out[18][285],u_xpb_out[19][285],u_xpb_out[20][285],u_xpb_out[21][285],u_xpb_out[22][285],u_xpb_out[23][285],u_xpb_out[24][285],u_xpb_out[25][285],u_xpb_out[26][285],u_xpb_out[27][285],u_xpb_out[28][285],u_xpb_out[29][285],u_xpb_out[30][285],u_xpb_out[31][285],u_xpb_out[32][285],u_xpb_out[33][285],u_xpb_out[34][285],u_xpb_out[35][285],u_xpb_out[36][285],u_xpb_out[37][285],u_xpb_out[38][285],u_xpb_out[39][285],u_xpb_out[40][285],u_xpb_out[41][285],u_xpb_out[42][285],u_xpb_out[43][285],u_xpb_out[44][285],u_xpb_out[45][285],u_xpb_out[46][285],u_xpb_out[47][285],u_xpb_out[48][285],u_xpb_out[49][285],u_xpb_out[50][285],u_xpb_out[51][285],u_xpb_out[52][285],u_xpb_out[53][285],u_xpb_out[54][285],u_xpb_out[55][285],u_xpb_out[56][285],u_xpb_out[57][285],u_xpb_out[58][285],u_xpb_out[59][285],u_xpb_out[60][285],u_xpb_out[61][285],u_xpb_out[62][285],u_xpb_out[63][285],u_xpb_out[64][285],u_xpb_out[65][285],u_xpb_out[66][285],u_xpb_out[67][285],u_xpb_out[68][285],u_xpb_out[69][285],u_xpb_out[70][285],u_xpb_out[71][285],u_xpb_out[72][285],u_xpb_out[73][285],u_xpb_out[74][285],u_xpb_out[75][285],u_xpb_out[76][285],u_xpb_out[77][285],u_xpb_out[78][285],u_xpb_out[79][285],u_xpb_out[80][285],u_xpb_out[81][285],u_xpb_out[82][285],u_xpb_out[83][285],u_xpb_out[84][285],u_xpb_out[85][285],u_xpb_out[86][285],u_xpb_out[87][285],u_xpb_out[88][285],u_xpb_out[89][285],u_xpb_out[90][285],u_xpb_out[91][285],u_xpb_out[92][285],u_xpb_out[93][285],u_xpb_out[94][285],u_xpb_out[95][285],u_xpb_out[96][285],u_xpb_out[97][285],u_xpb_out[98][285],u_xpb_out[99][285],u_xpb_out[100][285],u_xpb_out[101][285],u_xpb_out[102][285],u_xpb_out[103][285],u_xpb_out[104][285],u_xpb_out[105][285]};

assign col_out_286 = {u_xpb_out[0][286],u_xpb_out[1][286],u_xpb_out[2][286],u_xpb_out[3][286],u_xpb_out[4][286],u_xpb_out[5][286],u_xpb_out[6][286],u_xpb_out[7][286],u_xpb_out[8][286],u_xpb_out[9][286],u_xpb_out[10][286],u_xpb_out[11][286],u_xpb_out[12][286],u_xpb_out[13][286],u_xpb_out[14][286],u_xpb_out[15][286],u_xpb_out[16][286],u_xpb_out[17][286],u_xpb_out[18][286],u_xpb_out[19][286],u_xpb_out[20][286],u_xpb_out[21][286],u_xpb_out[22][286],u_xpb_out[23][286],u_xpb_out[24][286],u_xpb_out[25][286],u_xpb_out[26][286],u_xpb_out[27][286],u_xpb_out[28][286],u_xpb_out[29][286],u_xpb_out[30][286],u_xpb_out[31][286],u_xpb_out[32][286],u_xpb_out[33][286],u_xpb_out[34][286],u_xpb_out[35][286],u_xpb_out[36][286],u_xpb_out[37][286],u_xpb_out[38][286],u_xpb_out[39][286],u_xpb_out[40][286],u_xpb_out[41][286],u_xpb_out[42][286],u_xpb_out[43][286],u_xpb_out[44][286],u_xpb_out[45][286],u_xpb_out[46][286],u_xpb_out[47][286],u_xpb_out[48][286],u_xpb_out[49][286],u_xpb_out[50][286],u_xpb_out[51][286],u_xpb_out[52][286],u_xpb_out[53][286],u_xpb_out[54][286],u_xpb_out[55][286],u_xpb_out[56][286],u_xpb_out[57][286],u_xpb_out[58][286],u_xpb_out[59][286],u_xpb_out[60][286],u_xpb_out[61][286],u_xpb_out[62][286],u_xpb_out[63][286],u_xpb_out[64][286],u_xpb_out[65][286],u_xpb_out[66][286],u_xpb_out[67][286],u_xpb_out[68][286],u_xpb_out[69][286],u_xpb_out[70][286],u_xpb_out[71][286],u_xpb_out[72][286],u_xpb_out[73][286],u_xpb_out[74][286],u_xpb_out[75][286],u_xpb_out[76][286],u_xpb_out[77][286],u_xpb_out[78][286],u_xpb_out[79][286],u_xpb_out[80][286],u_xpb_out[81][286],u_xpb_out[82][286],u_xpb_out[83][286],u_xpb_out[84][286],u_xpb_out[85][286],u_xpb_out[86][286],u_xpb_out[87][286],u_xpb_out[88][286],u_xpb_out[89][286],u_xpb_out[90][286],u_xpb_out[91][286],u_xpb_out[92][286],u_xpb_out[93][286],u_xpb_out[94][286],u_xpb_out[95][286],u_xpb_out[96][286],u_xpb_out[97][286],u_xpb_out[98][286],u_xpb_out[99][286],u_xpb_out[100][286],u_xpb_out[101][286],u_xpb_out[102][286],u_xpb_out[103][286],u_xpb_out[104][286],u_xpb_out[105][286]};

assign col_out_287 = {u_xpb_out[0][287],u_xpb_out[1][287],u_xpb_out[2][287],u_xpb_out[3][287],u_xpb_out[4][287],u_xpb_out[5][287],u_xpb_out[6][287],u_xpb_out[7][287],u_xpb_out[8][287],u_xpb_out[9][287],u_xpb_out[10][287],u_xpb_out[11][287],u_xpb_out[12][287],u_xpb_out[13][287],u_xpb_out[14][287],u_xpb_out[15][287],u_xpb_out[16][287],u_xpb_out[17][287],u_xpb_out[18][287],u_xpb_out[19][287],u_xpb_out[20][287],u_xpb_out[21][287],u_xpb_out[22][287],u_xpb_out[23][287],u_xpb_out[24][287],u_xpb_out[25][287],u_xpb_out[26][287],u_xpb_out[27][287],u_xpb_out[28][287],u_xpb_out[29][287],u_xpb_out[30][287],u_xpb_out[31][287],u_xpb_out[32][287],u_xpb_out[33][287],u_xpb_out[34][287],u_xpb_out[35][287],u_xpb_out[36][287],u_xpb_out[37][287],u_xpb_out[38][287],u_xpb_out[39][287],u_xpb_out[40][287],u_xpb_out[41][287],u_xpb_out[42][287],u_xpb_out[43][287],u_xpb_out[44][287],u_xpb_out[45][287],u_xpb_out[46][287],u_xpb_out[47][287],u_xpb_out[48][287],u_xpb_out[49][287],u_xpb_out[50][287],u_xpb_out[51][287],u_xpb_out[52][287],u_xpb_out[53][287],u_xpb_out[54][287],u_xpb_out[55][287],u_xpb_out[56][287],u_xpb_out[57][287],u_xpb_out[58][287],u_xpb_out[59][287],u_xpb_out[60][287],u_xpb_out[61][287],u_xpb_out[62][287],u_xpb_out[63][287],u_xpb_out[64][287],u_xpb_out[65][287],u_xpb_out[66][287],u_xpb_out[67][287],u_xpb_out[68][287],u_xpb_out[69][287],u_xpb_out[70][287],u_xpb_out[71][287],u_xpb_out[72][287],u_xpb_out[73][287],u_xpb_out[74][287],u_xpb_out[75][287],u_xpb_out[76][287],u_xpb_out[77][287],u_xpb_out[78][287],u_xpb_out[79][287],u_xpb_out[80][287],u_xpb_out[81][287],u_xpb_out[82][287],u_xpb_out[83][287],u_xpb_out[84][287],u_xpb_out[85][287],u_xpb_out[86][287],u_xpb_out[87][287],u_xpb_out[88][287],u_xpb_out[89][287],u_xpb_out[90][287],u_xpb_out[91][287],u_xpb_out[92][287],u_xpb_out[93][287],u_xpb_out[94][287],u_xpb_out[95][287],u_xpb_out[96][287],u_xpb_out[97][287],u_xpb_out[98][287],u_xpb_out[99][287],u_xpb_out[100][287],u_xpb_out[101][287],u_xpb_out[102][287],u_xpb_out[103][287],u_xpb_out[104][287],u_xpb_out[105][287]};

assign col_out_288 = {u_xpb_out[0][288],u_xpb_out[1][288],u_xpb_out[2][288],u_xpb_out[3][288],u_xpb_out[4][288],u_xpb_out[5][288],u_xpb_out[6][288],u_xpb_out[7][288],u_xpb_out[8][288],u_xpb_out[9][288],u_xpb_out[10][288],u_xpb_out[11][288],u_xpb_out[12][288],u_xpb_out[13][288],u_xpb_out[14][288],u_xpb_out[15][288],u_xpb_out[16][288],u_xpb_out[17][288],u_xpb_out[18][288],u_xpb_out[19][288],u_xpb_out[20][288],u_xpb_out[21][288],u_xpb_out[22][288],u_xpb_out[23][288],u_xpb_out[24][288],u_xpb_out[25][288],u_xpb_out[26][288],u_xpb_out[27][288],u_xpb_out[28][288],u_xpb_out[29][288],u_xpb_out[30][288],u_xpb_out[31][288],u_xpb_out[32][288],u_xpb_out[33][288],u_xpb_out[34][288],u_xpb_out[35][288],u_xpb_out[36][288],u_xpb_out[37][288],u_xpb_out[38][288],u_xpb_out[39][288],u_xpb_out[40][288],u_xpb_out[41][288],u_xpb_out[42][288],u_xpb_out[43][288],u_xpb_out[44][288],u_xpb_out[45][288],u_xpb_out[46][288],u_xpb_out[47][288],u_xpb_out[48][288],u_xpb_out[49][288],u_xpb_out[50][288],u_xpb_out[51][288],u_xpb_out[52][288],u_xpb_out[53][288],u_xpb_out[54][288],u_xpb_out[55][288],u_xpb_out[56][288],u_xpb_out[57][288],u_xpb_out[58][288],u_xpb_out[59][288],u_xpb_out[60][288],u_xpb_out[61][288],u_xpb_out[62][288],u_xpb_out[63][288],u_xpb_out[64][288],u_xpb_out[65][288],u_xpb_out[66][288],u_xpb_out[67][288],u_xpb_out[68][288],u_xpb_out[69][288],u_xpb_out[70][288],u_xpb_out[71][288],u_xpb_out[72][288],u_xpb_out[73][288],u_xpb_out[74][288],u_xpb_out[75][288],u_xpb_out[76][288],u_xpb_out[77][288],u_xpb_out[78][288],u_xpb_out[79][288],u_xpb_out[80][288],u_xpb_out[81][288],u_xpb_out[82][288],u_xpb_out[83][288],u_xpb_out[84][288],u_xpb_out[85][288],u_xpb_out[86][288],u_xpb_out[87][288],u_xpb_out[88][288],u_xpb_out[89][288],u_xpb_out[90][288],u_xpb_out[91][288],u_xpb_out[92][288],u_xpb_out[93][288],u_xpb_out[94][288],u_xpb_out[95][288],u_xpb_out[96][288],u_xpb_out[97][288],u_xpb_out[98][288],u_xpb_out[99][288],u_xpb_out[100][288],u_xpb_out[101][288],u_xpb_out[102][288],u_xpb_out[103][288],u_xpb_out[104][288],u_xpb_out[105][288]};

assign col_out_289 = {u_xpb_out[0][289],u_xpb_out[1][289],u_xpb_out[2][289],u_xpb_out[3][289],u_xpb_out[4][289],u_xpb_out[5][289],u_xpb_out[6][289],u_xpb_out[7][289],u_xpb_out[8][289],u_xpb_out[9][289],u_xpb_out[10][289],u_xpb_out[11][289],u_xpb_out[12][289],u_xpb_out[13][289],u_xpb_out[14][289],u_xpb_out[15][289],u_xpb_out[16][289],u_xpb_out[17][289],u_xpb_out[18][289],u_xpb_out[19][289],u_xpb_out[20][289],u_xpb_out[21][289],u_xpb_out[22][289],u_xpb_out[23][289],u_xpb_out[24][289],u_xpb_out[25][289],u_xpb_out[26][289],u_xpb_out[27][289],u_xpb_out[28][289],u_xpb_out[29][289],u_xpb_out[30][289],u_xpb_out[31][289],u_xpb_out[32][289],u_xpb_out[33][289],u_xpb_out[34][289],u_xpb_out[35][289],u_xpb_out[36][289],u_xpb_out[37][289],u_xpb_out[38][289],u_xpb_out[39][289],u_xpb_out[40][289],u_xpb_out[41][289],u_xpb_out[42][289],u_xpb_out[43][289],u_xpb_out[44][289],u_xpb_out[45][289],u_xpb_out[46][289],u_xpb_out[47][289],u_xpb_out[48][289],u_xpb_out[49][289],u_xpb_out[50][289],u_xpb_out[51][289],u_xpb_out[52][289],u_xpb_out[53][289],u_xpb_out[54][289],u_xpb_out[55][289],u_xpb_out[56][289],u_xpb_out[57][289],u_xpb_out[58][289],u_xpb_out[59][289],u_xpb_out[60][289],u_xpb_out[61][289],u_xpb_out[62][289],u_xpb_out[63][289],u_xpb_out[64][289],u_xpb_out[65][289],u_xpb_out[66][289],u_xpb_out[67][289],u_xpb_out[68][289],u_xpb_out[69][289],u_xpb_out[70][289],u_xpb_out[71][289],u_xpb_out[72][289],u_xpb_out[73][289],u_xpb_out[74][289],u_xpb_out[75][289],u_xpb_out[76][289],u_xpb_out[77][289],u_xpb_out[78][289],u_xpb_out[79][289],u_xpb_out[80][289],u_xpb_out[81][289],u_xpb_out[82][289],u_xpb_out[83][289],u_xpb_out[84][289],u_xpb_out[85][289],u_xpb_out[86][289],u_xpb_out[87][289],u_xpb_out[88][289],u_xpb_out[89][289],u_xpb_out[90][289],u_xpb_out[91][289],u_xpb_out[92][289],u_xpb_out[93][289],u_xpb_out[94][289],u_xpb_out[95][289],u_xpb_out[96][289],u_xpb_out[97][289],u_xpb_out[98][289],u_xpb_out[99][289],u_xpb_out[100][289],u_xpb_out[101][289],u_xpb_out[102][289],u_xpb_out[103][289],u_xpb_out[104][289],u_xpb_out[105][289]};

assign col_out_290 = {u_xpb_out[0][290],u_xpb_out[1][290],u_xpb_out[2][290],u_xpb_out[3][290],u_xpb_out[4][290],u_xpb_out[5][290],u_xpb_out[6][290],u_xpb_out[7][290],u_xpb_out[8][290],u_xpb_out[9][290],u_xpb_out[10][290],u_xpb_out[11][290],u_xpb_out[12][290],u_xpb_out[13][290],u_xpb_out[14][290],u_xpb_out[15][290],u_xpb_out[16][290],u_xpb_out[17][290],u_xpb_out[18][290],u_xpb_out[19][290],u_xpb_out[20][290],u_xpb_out[21][290],u_xpb_out[22][290],u_xpb_out[23][290],u_xpb_out[24][290],u_xpb_out[25][290],u_xpb_out[26][290],u_xpb_out[27][290],u_xpb_out[28][290],u_xpb_out[29][290],u_xpb_out[30][290],u_xpb_out[31][290],u_xpb_out[32][290],u_xpb_out[33][290],u_xpb_out[34][290],u_xpb_out[35][290],u_xpb_out[36][290],u_xpb_out[37][290],u_xpb_out[38][290],u_xpb_out[39][290],u_xpb_out[40][290],u_xpb_out[41][290],u_xpb_out[42][290],u_xpb_out[43][290],u_xpb_out[44][290],u_xpb_out[45][290],u_xpb_out[46][290],u_xpb_out[47][290],u_xpb_out[48][290],u_xpb_out[49][290],u_xpb_out[50][290],u_xpb_out[51][290],u_xpb_out[52][290],u_xpb_out[53][290],u_xpb_out[54][290],u_xpb_out[55][290],u_xpb_out[56][290],u_xpb_out[57][290],u_xpb_out[58][290],u_xpb_out[59][290],u_xpb_out[60][290],u_xpb_out[61][290],u_xpb_out[62][290],u_xpb_out[63][290],u_xpb_out[64][290],u_xpb_out[65][290],u_xpb_out[66][290],u_xpb_out[67][290],u_xpb_out[68][290],u_xpb_out[69][290],u_xpb_out[70][290],u_xpb_out[71][290],u_xpb_out[72][290],u_xpb_out[73][290],u_xpb_out[74][290],u_xpb_out[75][290],u_xpb_out[76][290],u_xpb_out[77][290],u_xpb_out[78][290],u_xpb_out[79][290],u_xpb_out[80][290],u_xpb_out[81][290],u_xpb_out[82][290],u_xpb_out[83][290],u_xpb_out[84][290],u_xpb_out[85][290],u_xpb_out[86][290],u_xpb_out[87][290],u_xpb_out[88][290],u_xpb_out[89][290],u_xpb_out[90][290],u_xpb_out[91][290],u_xpb_out[92][290],u_xpb_out[93][290],u_xpb_out[94][290],u_xpb_out[95][290],u_xpb_out[96][290],u_xpb_out[97][290],u_xpb_out[98][290],u_xpb_out[99][290],u_xpb_out[100][290],u_xpb_out[101][290],u_xpb_out[102][290],u_xpb_out[103][290],u_xpb_out[104][290],u_xpb_out[105][290]};

assign col_out_291 = {u_xpb_out[0][291],u_xpb_out[1][291],u_xpb_out[2][291],u_xpb_out[3][291],u_xpb_out[4][291],u_xpb_out[5][291],u_xpb_out[6][291],u_xpb_out[7][291],u_xpb_out[8][291],u_xpb_out[9][291],u_xpb_out[10][291],u_xpb_out[11][291],u_xpb_out[12][291],u_xpb_out[13][291],u_xpb_out[14][291],u_xpb_out[15][291],u_xpb_out[16][291],u_xpb_out[17][291],u_xpb_out[18][291],u_xpb_out[19][291],u_xpb_out[20][291],u_xpb_out[21][291],u_xpb_out[22][291],u_xpb_out[23][291],u_xpb_out[24][291],u_xpb_out[25][291],u_xpb_out[26][291],u_xpb_out[27][291],u_xpb_out[28][291],u_xpb_out[29][291],u_xpb_out[30][291],u_xpb_out[31][291],u_xpb_out[32][291],u_xpb_out[33][291],u_xpb_out[34][291],u_xpb_out[35][291],u_xpb_out[36][291],u_xpb_out[37][291],u_xpb_out[38][291],u_xpb_out[39][291],u_xpb_out[40][291],u_xpb_out[41][291],u_xpb_out[42][291],u_xpb_out[43][291],u_xpb_out[44][291],u_xpb_out[45][291],u_xpb_out[46][291],u_xpb_out[47][291],u_xpb_out[48][291],u_xpb_out[49][291],u_xpb_out[50][291],u_xpb_out[51][291],u_xpb_out[52][291],u_xpb_out[53][291],u_xpb_out[54][291],u_xpb_out[55][291],u_xpb_out[56][291],u_xpb_out[57][291],u_xpb_out[58][291],u_xpb_out[59][291],u_xpb_out[60][291],u_xpb_out[61][291],u_xpb_out[62][291],u_xpb_out[63][291],u_xpb_out[64][291],u_xpb_out[65][291],u_xpb_out[66][291],u_xpb_out[67][291],u_xpb_out[68][291],u_xpb_out[69][291],u_xpb_out[70][291],u_xpb_out[71][291],u_xpb_out[72][291],u_xpb_out[73][291],u_xpb_out[74][291],u_xpb_out[75][291],u_xpb_out[76][291],u_xpb_out[77][291],u_xpb_out[78][291],u_xpb_out[79][291],u_xpb_out[80][291],u_xpb_out[81][291],u_xpb_out[82][291],u_xpb_out[83][291],u_xpb_out[84][291],u_xpb_out[85][291],u_xpb_out[86][291],u_xpb_out[87][291],u_xpb_out[88][291],u_xpb_out[89][291],u_xpb_out[90][291],u_xpb_out[91][291],u_xpb_out[92][291],u_xpb_out[93][291],u_xpb_out[94][291],u_xpb_out[95][291],u_xpb_out[96][291],u_xpb_out[97][291],u_xpb_out[98][291],u_xpb_out[99][291],u_xpb_out[100][291],u_xpb_out[101][291],u_xpb_out[102][291],u_xpb_out[103][291],u_xpb_out[104][291],u_xpb_out[105][291]};

assign col_out_292 = {u_xpb_out[0][292],u_xpb_out[1][292],u_xpb_out[2][292],u_xpb_out[3][292],u_xpb_out[4][292],u_xpb_out[5][292],u_xpb_out[6][292],u_xpb_out[7][292],u_xpb_out[8][292],u_xpb_out[9][292],u_xpb_out[10][292],u_xpb_out[11][292],u_xpb_out[12][292],u_xpb_out[13][292],u_xpb_out[14][292],u_xpb_out[15][292],u_xpb_out[16][292],u_xpb_out[17][292],u_xpb_out[18][292],u_xpb_out[19][292],u_xpb_out[20][292],u_xpb_out[21][292],u_xpb_out[22][292],u_xpb_out[23][292],u_xpb_out[24][292],u_xpb_out[25][292],u_xpb_out[26][292],u_xpb_out[27][292],u_xpb_out[28][292],u_xpb_out[29][292],u_xpb_out[30][292],u_xpb_out[31][292],u_xpb_out[32][292],u_xpb_out[33][292],u_xpb_out[34][292],u_xpb_out[35][292],u_xpb_out[36][292],u_xpb_out[37][292],u_xpb_out[38][292],u_xpb_out[39][292],u_xpb_out[40][292],u_xpb_out[41][292],u_xpb_out[42][292],u_xpb_out[43][292],u_xpb_out[44][292],u_xpb_out[45][292],u_xpb_out[46][292],u_xpb_out[47][292],u_xpb_out[48][292],u_xpb_out[49][292],u_xpb_out[50][292],u_xpb_out[51][292],u_xpb_out[52][292],u_xpb_out[53][292],u_xpb_out[54][292],u_xpb_out[55][292],u_xpb_out[56][292],u_xpb_out[57][292],u_xpb_out[58][292],u_xpb_out[59][292],u_xpb_out[60][292],u_xpb_out[61][292],u_xpb_out[62][292],u_xpb_out[63][292],u_xpb_out[64][292],u_xpb_out[65][292],u_xpb_out[66][292],u_xpb_out[67][292],u_xpb_out[68][292],u_xpb_out[69][292],u_xpb_out[70][292],u_xpb_out[71][292],u_xpb_out[72][292],u_xpb_out[73][292],u_xpb_out[74][292],u_xpb_out[75][292],u_xpb_out[76][292],u_xpb_out[77][292],u_xpb_out[78][292],u_xpb_out[79][292],u_xpb_out[80][292],u_xpb_out[81][292],u_xpb_out[82][292],u_xpb_out[83][292],u_xpb_out[84][292],u_xpb_out[85][292],u_xpb_out[86][292],u_xpb_out[87][292],u_xpb_out[88][292],u_xpb_out[89][292],u_xpb_out[90][292],u_xpb_out[91][292],u_xpb_out[92][292],u_xpb_out[93][292],u_xpb_out[94][292],u_xpb_out[95][292],u_xpb_out[96][292],u_xpb_out[97][292],u_xpb_out[98][292],u_xpb_out[99][292],u_xpb_out[100][292],u_xpb_out[101][292],u_xpb_out[102][292],u_xpb_out[103][292],u_xpb_out[104][292],u_xpb_out[105][292]};

assign col_out_293 = {u_xpb_out[0][293],u_xpb_out[1][293],u_xpb_out[2][293],u_xpb_out[3][293],u_xpb_out[4][293],u_xpb_out[5][293],u_xpb_out[6][293],u_xpb_out[7][293],u_xpb_out[8][293],u_xpb_out[9][293],u_xpb_out[10][293],u_xpb_out[11][293],u_xpb_out[12][293],u_xpb_out[13][293],u_xpb_out[14][293],u_xpb_out[15][293],u_xpb_out[16][293],u_xpb_out[17][293],u_xpb_out[18][293],u_xpb_out[19][293],u_xpb_out[20][293],u_xpb_out[21][293],u_xpb_out[22][293],u_xpb_out[23][293],u_xpb_out[24][293],u_xpb_out[25][293],u_xpb_out[26][293],u_xpb_out[27][293],u_xpb_out[28][293],u_xpb_out[29][293],u_xpb_out[30][293],u_xpb_out[31][293],u_xpb_out[32][293],u_xpb_out[33][293],u_xpb_out[34][293],u_xpb_out[35][293],u_xpb_out[36][293],u_xpb_out[37][293],u_xpb_out[38][293],u_xpb_out[39][293],u_xpb_out[40][293],u_xpb_out[41][293],u_xpb_out[42][293],u_xpb_out[43][293],u_xpb_out[44][293],u_xpb_out[45][293],u_xpb_out[46][293],u_xpb_out[47][293],u_xpb_out[48][293],u_xpb_out[49][293],u_xpb_out[50][293],u_xpb_out[51][293],u_xpb_out[52][293],u_xpb_out[53][293],u_xpb_out[54][293],u_xpb_out[55][293],u_xpb_out[56][293],u_xpb_out[57][293],u_xpb_out[58][293],u_xpb_out[59][293],u_xpb_out[60][293],u_xpb_out[61][293],u_xpb_out[62][293],u_xpb_out[63][293],u_xpb_out[64][293],u_xpb_out[65][293],u_xpb_out[66][293],u_xpb_out[67][293],u_xpb_out[68][293],u_xpb_out[69][293],u_xpb_out[70][293],u_xpb_out[71][293],u_xpb_out[72][293],u_xpb_out[73][293],u_xpb_out[74][293],u_xpb_out[75][293],u_xpb_out[76][293],u_xpb_out[77][293],u_xpb_out[78][293],u_xpb_out[79][293],u_xpb_out[80][293],u_xpb_out[81][293],u_xpb_out[82][293],u_xpb_out[83][293],u_xpb_out[84][293],u_xpb_out[85][293],u_xpb_out[86][293],u_xpb_out[87][293],u_xpb_out[88][293],u_xpb_out[89][293],u_xpb_out[90][293],u_xpb_out[91][293],u_xpb_out[92][293],u_xpb_out[93][293],u_xpb_out[94][293],u_xpb_out[95][293],u_xpb_out[96][293],u_xpb_out[97][293],u_xpb_out[98][293],u_xpb_out[99][293],u_xpb_out[100][293],u_xpb_out[101][293],u_xpb_out[102][293],u_xpb_out[103][293],u_xpb_out[104][293],u_xpb_out[105][293]};

assign col_out_294 = {u_xpb_out[0][294],u_xpb_out[1][294],u_xpb_out[2][294],u_xpb_out[3][294],u_xpb_out[4][294],u_xpb_out[5][294],u_xpb_out[6][294],u_xpb_out[7][294],u_xpb_out[8][294],u_xpb_out[9][294],u_xpb_out[10][294],u_xpb_out[11][294],u_xpb_out[12][294],u_xpb_out[13][294],u_xpb_out[14][294],u_xpb_out[15][294],u_xpb_out[16][294],u_xpb_out[17][294],u_xpb_out[18][294],u_xpb_out[19][294],u_xpb_out[20][294],u_xpb_out[21][294],u_xpb_out[22][294],u_xpb_out[23][294],u_xpb_out[24][294],u_xpb_out[25][294],u_xpb_out[26][294],u_xpb_out[27][294],u_xpb_out[28][294],u_xpb_out[29][294],u_xpb_out[30][294],u_xpb_out[31][294],u_xpb_out[32][294],u_xpb_out[33][294],u_xpb_out[34][294],u_xpb_out[35][294],u_xpb_out[36][294],u_xpb_out[37][294],u_xpb_out[38][294],u_xpb_out[39][294],u_xpb_out[40][294],u_xpb_out[41][294],u_xpb_out[42][294],u_xpb_out[43][294],u_xpb_out[44][294],u_xpb_out[45][294],u_xpb_out[46][294],u_xpb_out[47][294],u_xpb_out[48][294],u_xpb_out[49][294],u_xpb_out[50][294],u_xpb_out[51][294],u_xpb_out[52][294],u_xpb_out[53][294],u_xpb_out[54][294],u_xpb_out[55][294],u_xpb_out[56][294],u_xpb_out[57][294],u_xpb_out[58][294],u_xpb_out[59][294],u_xpb_out[60][294],u_xpb_out[61][294],u_xpb_out[62][294],u_xpb_out[63][294],u_xpb_out[64][294],u_xpb_out[65][294],u_xpb_out[66][294],u_xpb_out[67][294],u_xpb_out[68][294],u_xpb_out[69][294],u_xpb_out[70][294],u_xpb_out[71][294],u_xpb_out[72][294],u_xpb_out[73][294],u_xpb_out[74][294],u_xpb_out[75][294],u_xpb_out[76][294],u_xpb_out[77][294],u_xpb_out[78][294],u_xpb_out[79][294],u_xpb_out[80][294],u_xpb_out[81][294],u_xpb_out[82][294],u_xpb_out[83][294],u_xpb_out[84][294],u_xpb_out[85][294],u_xpb_out[86][294],u_xpb_out[87][294],u_xpb_out[88][294],u_xpb_out[89][294],u_xpb_out[90][294],u_xpb_out[91][294],u_xpb_out[92][294],u_xpb_out[93][294],u_xpb_out[94][294],u_xpb_out[95][294],u_xpb_out[96][294],u_xpb_out[97][294],u_xpb_out[98][294],u_xpb_out[99][294],u_xpb_out[100][294],u_xpb_out[101][294],u_xpb_out[102][294],u_xpb_out[103][294],u_xpb_out[104][294],u_xpb_out[105][294]};

assign col_out_295 = {u_xpb_out[0][295],u_xpb_out[1][295],u_xpb_out[2][295],u_xpb_out[3][295],u_xpb_out[4][295],u_xpb_out[5][295],u_xpb_out[6][295],u_xpb_out[7][295],u_xpb_out[8][295],u_xpb_out[9][295],u_xpb_out[10][295],u_xpb_out[11][295],u_xpb_out[12][295],u_xpb_out[13][295],u_xpb_out[14][295],u_xpb_out[15][295],u_xpb_out[16][295],u_xpb_out[17][295],u_xpb_out[18][295],u_xpb_out[19][295],u_xpb_out[20][295],u_xpb_out[21][295],u_xpb_out[22][295],u_xpb_out[23][295],u_xpb_out[24][295],u_xpb_out[25][295],u_xpb_out[26][295],u_xpb_out[27][295],u_xpb_out[28][295],u_xpb_out[29][295],u_xpb_out[30][295],u_xpb_out[31][295],u_xpb_out[32][295],u_xpb_out[33][295],u_xpb_out[34][295],u_xpb_out[35][295],u_xpb_out[36][295],u_xpb_out[37][295],u_xpb_out[38][295],u_xpb_out[39][295],u_xpb_out[40][295],u_xpb_out[41][295],u_xpb_out[42][295],u_xpb_out[43][295],u_xpb_out[44][295],u_xpb_out[45][295],u_xpb_out[46][295],u_xpb_out[47][295],u_xpb_out[48][295],u_xpb_out[49][295],u_xpb_out[50][295],u_xpb_out[51][295],u_xpb_out[52][295],u_xpb_out[53][295],u_xpb_out[54][295],u_xpb_out[55][295],u_xpb_out[56][295],u_xpb_out[57][295],u_xpb_out[58][295],u_xpb_out[59][295],u_xpb_out[60][295],u_xpb_out[61][295],u_xpb_out[62][295],u_xpb_out[63][295],u_xpb_out[64][295],u_xpb_out[65][295],u_xpb_out[66][295],u_xpb_out[67][295],u_xpb_out[68][295],u_xpb_out[69][295],u_xpb_out[70][295],u_xpb_out[71][295],u_xpb_out[72][295],u_xpb_out[73][295],u_xpb_out[74][295],u_xpb_out[75][295],u_xpb_out[76][295],u_xpb_out[77][295],u_xpb_out[78][295],u_xpb_out[79][295],u_xpb_out[80][295],u_xpb_out[81][295],u_xpb_out[82][295],u_xpb_out[83][295],u_xpb_out[84][295],u_xpb_out[85][295],u_xpb_out[86][295],u_xpb_out[87][295],u_xpb_out[88][295],u_xpb_out[89][295],u_xpb_out[90][295],u_xpb_out[91][295],u_xpb_out[92][295],u_xpb_out[93][295],u_xpb_out[94][295],u_xpb_out[95][295],u_xpb_out[96][295],u_xpb_out[97][295],u_xpb_out[98][295],u_xpb_out[99][295],u_xpb_out[100][295],u_xpb_out[101][295],u_xpb_out[102][295],u_xpb_out[103][295],u_xpb_out[104][295],u_xpb_out[105][295]};

assign col_out_296 = {u_xpb_out[0][296],u_xpb_out[1][296],u_xpb_out[2][296],u_xpb_out[3][296],u_xpb_out[4][296],u_xpb_out[5][296],u_xpb_out[6][296],u_xpb_out[7][296],u_xpb_out[8][296],u_xpb_out[9][296],u_xpb_out[10][296],u_xpb_out[11][296],u_xpb_out[12][296],u_xpb_out[13][296],u_xpb_out[14][296],u_xpb_out[15][296],u_xpb_out[16][296],u_xpb_out[17][296],u_xpb_out[18][296],u_xpb_out[19][296],u_xpb_out[20][296],u_xpb_out[21][296],u_xpb_out[22][296],u_xpb_out[23][296],u_xpb_out[24][296],u_xpb_out[25][296],u_xpb_out[26][296],u_xpb_out[27][296],u_xpb_out[28][296],u_xpb_out[29][296],u_xpb_out[30][296],u_xpb_out[31][296],u_xpb_out[32][296],u_xpb_out[33][296],u_xpb_out[34][296],u_xpb_out[35][296],u_xpb_out[36][296],u_xpb_out[37][296],u_xpb_out[38][296],u_xpb_out[39][296],u_xpb_out[40][296],u_xpb_out[41][296],u_xpb_out[42][296],u_xpb_out[43][296],u_xpb_out[44][296],u_xpb_out[45][296],u_xpb_out[46][296],u_xpb_out[47][296],u_xpb_out[48][296],u_xpb_out[49][296],u_xpb_out[50][296],u_xpb_out[51][296],u_xpb_out[52][296],u_xpb_out[53][296],u_xpb_out[54][296],u_xpb_out[55][296],u_xpb_out[56][296],u_xpb_out[57][296],u_xpb_out[58][296],u_xpb_out[59][296],u_xpb_out[60][296],u_xpb_out[61][296],u_xpb_out[62][296],u_xpb_out[63][296],u_xpb_out[64][296],u_xpb_out[65][296],u_xpb_out[66][296],u_xpb_out[67][296],u_xpb_out[68][296],u_xpb_out[69][296],u_xpb_out[70][296],u_xpb_out[71][296],u_xpb_out[72][296],u_xpb_out[73][296],u_xpb_out[74][296],u_xpb_out[75][296],u_xpb_out[76][296],u_xpb_out[77][296],u_xpb_out[78][296],u_xpb_out[79][296],u_xpb_out[80][296],u_xpb_out[81][296],u_xpb_out[82][296],u_xpb_out[83][296],u_xpb_out[84][296],u_xpb_out[85][296],u_xpb_out[86][296],u_xpb_out[87][296],u_xpb_out[88][296],u_xpb_out[89][296],u_xpb_out[90][296],u_xpb_out[91][296],u_xpb_out[92][296],u_xpb_out[93][296],u_xpb_out[94][296],u_xpb_out[95][296],u_xpb_out[96][296],u_xpb_out[97][296],u_xpb_out[98][296],u_xpb_out[99][296],u_xpb_out[100][296],u_xpb_out[101][296],u_xpb_out[102][296],u_xpb_out[103][296],u_xpb_out[104][296],u_xpb_out[105][296]};

assign col_out_297 = {u_xpb_out[0][297],u_xpb_out[1][297],u_xpb_out[2][297],u_xpb_out[3][297],u_xpb_out[4][297],u_xpb_out[5][297],u_xpb_out[6][297],u_xpb_out[7][297],u_xpb_out[8][297],u_xpb_out[9][297],u_xpb_out[10][297],u_xpb_out[11][297],u_xpb_out[12][297],u_xpb_out[13][297],u_xpb_out[14][297],u_xpb_out[15][297],u_xpb_out[16][297],u_xpb_out[17][297],u_xpb_out[18][297],u_xpb_out[19][297],u_xpb_out[20][297],u_xpb_out[21][297],u_xpb_out[22][297],u_xpb_out[23][297],u_xpb_out[24][297],u_xpb_out[25][297],u_xpb_out[26][297],u_xpb_out[27][297],u_xpb_out[28][297],u_xpb_out[29][297],u_xpb_out[30][297],u_xpb_out[31][297],u_xpb_out[32][297],u_xpb_out[33][297],u_xpb_out[34][297],u_xpb_out[35][297],u_xpb_out[36][297],u_xpb_out[37][297],u_xpb_out[38][297],u_xpb_out[39][297],u_xpb_out[40][297],u_xpb_out[41][297],u_xpb_out[42][297],u_xpb_out[43][297],u_xpb_out[44][297],u_xpb_out[45][297],u_xpb_out[46][297],u_xpb_out[47][297],u_xpb_out[48][297],u_xpb_out[49][297],u_xpb_out[50][297],u_xpb_out[51][297],u_xpb_out[52][297],u_xpb_out[53][297],u_xpb_out[54][297],u_xpb_out[55][297],u_xpb_out[56][297],u_xpb_out[57][297],u_xpb_out[58][297],u_xpb_out[59][297],u_xpb_out[60][297],u_xpb_out[61][297],u_xpb_out[62][297],u_xpb_out[63][297],u_xpb_out[64][297],u_xpb_out[65][297],u_xpb_out[66][297],u_xpb_out[67][297],u_xpb_out[68][297],u_xpb_out[69][297],u_xpb_out[70][297],u_xpb_out[71][297],u_xpb_out[72][297],u_xpb_out[73][297],u_xpb_out[74][297],u_xpb_out[75][297],u_xpb_out[76][297],u_xpb_out[77][297],u_xpb_out[78][297],u_xpb_out[79][297],u_xpb_out[80][297],u_xpb_out[81][297],u_xpb_out[82][297],u_xpb_out[83][297],u_xpb_out[84][297],u_xpb_out[85][297],u_xpb_out[86][297],u_xpb_out[87][297],u_xpb_out[88][297],u_xpb_out[89][297],u_xpb_out[90][297],u_xpb_out[91][297],u_xpb_out[92][297],u_xpb_out[93][297],u_xpb_out[94][297],u_xpb_out[95][297],u_xpb_out[96][297],u_xpb_out[97][297],u_xpb_out[98][297],u_xpb_out[99][297],u_xpb_out[100][297],u_xpb_out[101][297],u_xpb_out[102][297],u_xpb_out[103][297],u_xpb_out[104][297],u_xpb_out[105][297]};

assign col_out_298 = {u_xpb_out[0][298],u_xpb_out[1][298],u_xpb_out[2][298],u_xpb_out[3][298],u_xpb_out[4][298],u_xpb_out[5][298],u_xpb_out[6][298],u_xpb_out[7][298],u_xpb_out[8][298],u_xpb_out[9][298],u_xpb_out[10][298],u_xpb_out[11][298],u_xpb_out[12][298],u_xpb_out[13][298],u_xpb_out[14][298],u_xpb_out[15][298],u_xpb_out[16][298],u_xpb_out[17][298],u_xpb_out[18][298],u_xpb_out[19][298],u_xpb_out[20][298],u_xpb_out[21][298],u_xpb_out[22][298],u_xpb_out[23][298],u_xpb_out[24][298],u_xpb_out[25][298],u_xpb_out[26][298],u_xpb_out[27][298],u_xpb_out[28][298],u_xpb_out[29][298],u_xpb_out[30][298],u_xpb_out[31][298],u_xpb_out[32][298],u_xpb_out[33][298],u_xpb_out[34][298],u_xpb_out[35][298],u_xpb_out[36][298],u_xpb_out[37][298],u_xpb_out[38][298],u_xpb_out[39][298],u_xpb_out[40][298],u_xpb_out[41][298],u_xpb_out[42][298],u_xpb_out[43][298],u_xpb_out[44][298],u_xpb_out[45][298],u_xpb_out[46][298],u_xpb_out[47][298],u_xpb_out[48][298],u_xpb_out[49][298],u_xpb_out[50][298],u_xpb_out[51][298],u_xpb_out[52][298],u_xpb_out[53][298],u_xpb_out[54][298],u_xpb_out[55][298],u_xpb_out[56][298],u_xpb_out[57][298],u_xpb_out[58][298],u_xpb_out[59][298],u_xpb_out[60][298],u_xpb_out[61][298],u_xpb_out[62][298],u_xpb_out[63][298],u_xpb_out[64][298],u_xpb_out[65][298],u_xpb_out[66][298],u_xpb_out[67][298],u_xpb_out[68][298],u_xpb_out[69][298],u_xpb_out[70][298],u_xpb_out[71][298],u_xpb_out[72][298],u_xpb_out[73][298],u_xpb_out[74][298],u_xpb_out[75][298],u_xpb_out[76][298],u_xpb_out[77][298],u_xpb_out[78][298],u_xpb_out[79][298],u_xpb_out[80][298],u_xpb_out[81][298],u_xpb_out[82][298],u_xpb_out[83][298],u_xpb_out[84][298],u_xpb_out[85][298],u_xpb_out[86][298],u_xpb_out[87][298],u_xpb_out[88][298],u_xpb_out[89][298],u_xpb_out[90][298],u_xpb_out[91][298],u_xpb_out[92][298],u_xpb_out[93][298],u_xpb_out[94][298],u_xpb_out[95][298],u_xpb_out[96][298],u_xpb_out[97][298],u_xpb_out[98][298],u_xpb_out[99][298],u_xpb_out[100][298],u_xpb_out[101][298],u_xpb_out[102][298],u_xpb_out[103][298],u_xpb_out[104][298],u_xpb_out[105][298]};

assign col_out_299 = {u_xpb_out[0][299],u_xpb_out[1][299],u_xpb_out[2][299],u_xpb_out[3][299],u_xpb_out[4][299],u_xpb_out[5][299],u_xpb_out[6][299],u_xpb_out[7][299],u_xpb_out[8][299],u_xpb_out[9][299],u_xpb_out[10][299],u_xpb_out[11][299],u_xpb_out[12][299],u_xpb_out[13][299],u_xpb_out[14][299],u_xpb_out[15][299],u_xpb_out[16][299],u_xpb_out[17][299],u_xpb_out[18][299],u_xpb_out[19][299],u_xpb_out[20][299],u_xpb_out[21][299],u_xpb_out[22][299],u_xpb_out[23][299],u_xpb_out[24][299],u_xpb_out[25][299],u_xpb_out[26][299],u_xpb_out[27][299],u_xpb_out[28][299],u_xpb_out[29][299],u_xpb_out[30][299],u_xpb_out[31][299],u_xpb_out[32][299],u_xpb_out[33][299],u_xpb_out[34][299],u_xpb_out[35][299],u_xpb_out[36][299],u_xpb_out[37][299],u_xpb_out[38][299],u_xpb_out[39][299],u_xpb_out[40][299],u_xpb_out[41][299],u_xpb_out[42][299],u_xpb_out[43][299],u_xpb_out[44][299],u_xpb_out[45][299],u_xpb_out[46][299],u_xpb_out[47][299],u_xpb_out[48][299],u_xpb_out[49][299],u_xpb_out[50][299],u_xpb_out[51][299],u_xpb_out[52][299],u_xpb_out[53][299],u_xpb_out[54][299],u_xpb_out[55][299],u_xpb_out[56][299],u_xpb_out[57][299],u_xpb_out[58][299],u_xpb_out[59][299],u_xpb_out[60][299],u_xpb_out[61][299],u_xpb_out[62][299],u_xpb_out[63][299],u_xpb_out[64][299],u_xpb_out[65][299],u_xpb_out[66][299],u_xpb_out[67][299],u_xpb_out[68][299],u_xpb_out[69][299],u_xpb_out[70][299],u_xpb_out[71][299],u_xpb_out[72][299],u_xpb_out[73][299],u_xpb_out[74][299],u_xpb_out[75][299],u_xpb_out[76][299],u_xpb_out[77][299],u_xpb_out[78][299],u_xpb_out[79][299],u_xpb_out[80][299],u_xpb_out[81][299],u_xpb_out[82][299],u_xpb_out[83][299],u_xpb_out[84][299],u_xpb_out[85][299],u_xpb_out[86][299],u_xpb_out[87][299],u_xpb_out[88][299],u_xpb_out[89][299],u_xpb_out[90][299],u_xpb_out[91][299],u_xpb_out[92][299],u_xpb_out[93][299],u_xpb_out[94][299],u_xpb_out[95][299],u_xpb_out[96][299],u_xpb_out[97][299],u_xpb_out[98][299],u_xpb_out[99][299],u_xpb_out[100][299],u_xpb_out[101][299],u_xpb_out[102][299],u_xpb_out[103][299],u_xpb_out[104][299],u_xpb_out[105][299]};

assign col_out_300 = {u_xpb_out[0][300],u_xpb_out[1][300],u_xpb_out[2][300],u_xpb_out[3][300],u_xpb_out[4][300],u_xpb_out[5][300],u_xpb_out[6][300],u_xpb_out[7][300],u_xpb_out[8][300],u_xpb_out[9][300],u_xpb_out[10][300],u_xpb_out[11][300],u_xpb_out[12][300],u_xpb_out[13][300],u_xpb_out[14][300],u_xpb_out[15][300],u_xpb_out[16][300],u_xpb_out[17][300],u_xpb_out[18][300],u_xpb_out[19][300],u_xpb_out[20][300],u_xpb_out[21][300],u_xpb_out[22][300],u_xpb_out[23][300],u_xpb_out[24][300],u_xpb_out[25][300],u_xpb_out[26][300],u_xpb_out[27][300],u_xpb_out[28][300],u_xpb_out[29][300],u_xpb_out[30][300],u_xpb_out[31][300],u_xpb_out[32][300],u_xpb_out[33][300],u_xpb_out[34][300],u_xpb_out[35][300],u_xpb_out[36][300],u_xpb_out[37][300],u_xpb_out[38][300],u_xpb_out[39][300],u_xpb_out[40][300],u_xpb_out[41][300],u_xpb_out[42][300],u_xpb_out[43][300],u_xpb_out[44][300],u_xpb_out[45][300],u_xpb_out[46][300],u_xpb_out[47][300],u_xpb_out[48][300],u_xpb_out[49][300],u_xpb_out[50][300],u_xpb_out[51][300],u_xpb_out[52][300],u_xpb_out[53][300],u_xpb_out[54][300],u_xpb_out[55][300],u_xpb_out[56][300],u_xpb_out[57][300],u_xpb_out[58][300],u_xpb_out[59][300],u_xpb_out[60][300],u_xpb_out[61][300],u_xpb_out[62][300],u_xpb_out[63][300],u_xpb_out[64][300],u_xpb_out[65][300],u_xpb_out[66][300],u_xpb_out[67][300],u_xpb_out[68][300],u_xpb_out[69][300],u_xpb_out[70][300],u_xpb_out[71][300],u_xpb_out[72][300],u_xpb_out[73][300],u_xpb_out[74][300],u_xpb_out[75][300],u_xpb_out[76][300],u_xpb_out[77][300],u_xpb_out[78][300],u_xpb_out[79][300],u_xpb_out[80][300],u_xpb_out[81][300],u_xpb_out[82][300],u_xpb_out[83][300],u_xpb_out[84][300],u_xpb_out[85][300],u_xpb_out[86][300],u_xpb_out[87][300],u_xpb_out[88][300],u_xpb_out[89][300],u_xpb_out[90][300],u_xpb_out[91][300],u_xpb_out[92][300],u_xpb_out[93][300],u_xpb_out[94][300],u_xpb_out[95][300],u_xpb_out[96][300],u_xpb_out[97][300],u_xpb_out[98][300],u_xpb_out[99][300],u_xpb_out[100][300],u_xpb_out[101][300],u_xpb_out[102][300],u_xpb_out[103][300],u_xpb_out[104][300],u_xpb_out[105][300]};

assign col_out_301 = {u_xpb_out[0][301],u_xpb_out[1][301],u_xpb_out[2][301],u_xpb_out[3][301],u_xpb_out[4][301],u_xpb_out[5][301],u_xpb_out[6][301],u_xpb_out[7][301],u_xpb_out[8][301],u_xpb_out[9][301],u_xpb_out[10][301],u_xpb_out[11][301],u_xpb_out[12][301],u_xpb_out[13][301],u_xpb_out[14][301],u_xpb_out[15][301],u_xpb_out[16][301],u_xpb_out[17][301],u_xpb_out[18][301],u_xpb_out[19][301],u_xpb_out[20][301],u_xpb_out[21][301],u_xpb_out[22][301],u_xpb_out[23][301],u_xpb_out[24][301],u_xpb_out[25][301],u_xpb_out[26][301],u_xpb_out[27][301],u_xpb_out[28][301],u_xpb_out[29][301],u_xpb_out[30][301],u_xpb_out[31][301],u_xpb_out[32][301],u_xpb_out[33][301],u_xpb_out[34][301],u_xpb_out[35][301],u_xpb_out[36][301],u_xpb_out[37][301],u_xpb_out[38][301],u_xpb_out[39][301],u_xpb_out[40][301],u_xpb_out[41][301],u_xpb_out[42][301],u_xpb_out[43][301],u_xpb_out[44][301],u_xpb_out[45][301],u_xpb_out[46][301],u_xpb_out[47][301],u_xpb_out[48][301],u_xpb_out[49][301],u_xpb_out[50][301],u_xpb_out[51][301],u_xpb_out[52][301],u_xpb_out[53][301],u_xpb_out[54][301],u_xpb_out[55][301],u_xpb_out[56][301],u_xpb_out[57][301],u_xpb_out[58][301],u_xpb_out[59][301],u_xpb_out[60][301],u_xpb_out[61][301],u_xpb_out[62][301],u_xpb_out[63][301],u_xpb_out[64][301],u_xpb_out[65][301],u_xpb_out[66][301],u_xpb_out[67][301],u_xpb_out[68][301],u_xpb_out[69][301],u_xpb_out[70][301],u_xpb_out[71][301],u_xpb_out[72][301],u_xpb_out[73][301],u_xpb_out[74][301],u_xpb_out[75][301],u_xpb_out[76][301],u_xpb_out[77][301],u_xpb_out[78][301],u_xpb_out[79][301],u_xpb_out[80][301],u_xpb_out[81][301],u_xpb_out[82][301],u_xpb_out[83][301],u_xpb_out[84][301],u_xpb_out[85][301],u_xpb_out[86][301],u_xpb_out[87][301],u_xpb_out[88][301],u_xpb_out[89][301],u_xpb_out[90][301],u_xpb_out[91][301],u_xpb_out[92][301],u_xpb_out[93][301],u_xpb_out[94][301],u_xpb_out[95][301],u_xpb_out[96][301],u_xpb_out[97][301],u_xpb_out[98][301],u_xpb_out[99][301],u_xpb_out[100][301],u_xpb_out[101][301],u_xpb_out[102][301],u_xpb_out[103][301],u_xpb_out[104][301],u_xpb_out[105][301]};

assign col_out_302 = {u_xpb_out[0][302],u_xpb_out[1][302],u_xpb_out[2][302],u_xpb_out[3][302],u_xpb_out[4][302],u_xpb_out[5][302],u_xpb_out[6][302],u_xpb_out[7][302],u_xpb_out[8][302],u_xpb_out[9][302],u_xpb_out[10][302],u_xpb_out[11][302],u_xpb_out[12][302],u_xpb_out[13][302],u_xpb_out[14][302],u_xpb_out[15][302],u_xpb_out[16][302],u_xpb_out[17][302],u_xpb_out[18][302],u_xpb_out[19][302],u_xpb_out[20][302],u_xpb_out[21][302],u_xpb_out[22][302],u_xpb_out[23][302],u_xpb_out[24][302],u_xpb_out[25][302],u_xpb_out[26][302],u_xpb_out[27][302],u_xpb_out[28][302],u_xpb_out[29][302],u_xpb_out[30][302],u_xpb_out[31][302],u_xpb_out[32][302],u_xpb_out[33][302],u_xpb_out[34][302],u_xpb_out[35][302],u_xpb_out[36][302],u_xpb_out[37][302],u_xpb_out[38][302],u_xpb_out[39][302],u_xpb_out[40][302],u_xpb_out[41][302],u_xpb_out[42][302],u_xpb_out[43][302],u_xpb_out[44][302],u_xpb_out[45][302],u_xpb_out[46][302],u_xpb_out[47][302],u_xpb_out[48][302],u_xpb_out[49][302],u_xpb_out[50][302],u_xpb_out[51][302],u_xpb_out[52][302],u_xpb_out[53][302],u_xpb_out[54][302],u_xpb_out[55][302],u_xpb_out[56][302],u_xpb_out[57][302],u_xpb_out[58][302],u_xpb_out[59][302],u_xpb_out[60][302],u_xpb_out[61][302],u_xpb_out[62][302],u_xpb_out[63][302],u_xpb_out[64][302],u_xpb_out[65][302],u_xpb_out[66][302],u_xpb_out[67][302],u_xpb_out[68][302],u_xpb_out[69][302],u_xpb_out[70][302],u_xpb_out[71][302],u_xpb_out[72][302],u_xpb_out[73][302],u_xpb_out[74][302],u_xpb_out[75][302],u_xpb_out[76][302],u_xpb_out[77][302],u_xpb_out[78][302],u_xpb_out[79][302],u_xpb_out[80][302],u_xpb_out[81][302],u_xpb_out[82][302],u_xpb_out[83][302],u_xpb_out[84][302],u_xpb_out[85][302],u_xpb_out[86][302],u_xpb_out[87][302],u_xpb_out[88][302],u_xpb_out[89][302],u_xpb_out[90][302],u_xpb_out[91][302],u_xpb_out[92][302],u_xpb_out[93][302],u_xpb_out[94][302],u_xpb_out[95][302],u_xpb_out[96][302],u_xpb_out[97][302],u_xpb_out[98][302],u_xpb_out[99][302],u_xpb_out[100][302],u_xpb_out[101][302],u_xpb_out[102][302],u_xpb_out[103][302],u_xpb_out[104][302],u_xpb_out[105][302]};

assign col_out_303 = {u_xpb_out[0][303],u_xpb_out[1][303],u_xpb_out[2][303],u_xpb_out[3][303],u_xpb_out[4][303],u_xpb_out[5][303],u_xpb_out[6][303],u_xpb_out[7][303],u_xpb_out[8][303],u_xpb_out[9][303],u_xpb_out[10][303],u_xpb_out[11][303],u_xpb_out[12][303],u_xpb_out[13][303],u_xpb_out[14][303],u_xpb_out[15][303],u_xpb_out[16][303],u_xpb_out[17][303],u_xpb_out[18][303],u_xpb_out[19][303],u_xpb_out[20][303],u_xpb_out[21][303],u_xpb_out[22][303],u_xpb_out[23][303],u_xpb_out[24][303],u_xpb_out[25][303],u_xpb_out[26][303],u_xpb_out[27][303],u_xpb_out[28][303],u_xpb_out[29][303],u_xpb_out[30][303],u_xpb_out[31][303],u_xpb_out[32][303],u_xpb_out[33][303],u_xpb_out[34][303],u_xpb_out[35][303],u_xpb_out[36][303],u_xpb_out[37][303],u_xpb_out[38][303],u_xpb_out[39][303],u_xpb_out[40][303],u_xpb_out[41][303],u_xpb_out[42][303],u_xpb_out[43][303],u_xpb_out[44][303],u_xpb_out[45][303],u_xpb_out[46][303],u_xpb_out[47][303],u_xpb_out[48][303],u_xpb_out[49][303],u_xpb_out[50][303],u_xpb_out[51][303],u_xpb_out[52][303],u_xpb_out[53][303],u_xpb_out[54][303],u_xpb_out[55][303],u_xpb_out[56][303],u_xpb_out[57][303],u_xpb_out[58][303],u_xpb_out[59][303],u_xpb_out[60][303],u_xpb_out[61][303],u_xpb_out[62][303],u_xpb_out[63][303],u_xpb_out[64][303],u_xpb_out[65][303],u_xpb_out[66][303],u_xpb_out[67][303],u_xpb_out[68][303],u_xpb_out[69][303],u_xpb_out[70][303],u_xpb_out[71][303],u_xpb_out[72][303],u_xpb_out[73][303],u_xpb_out[74][303],u_xpb_out[75][303],u_xpb_out[76][303],u_xpb_out[77][303],u_xpb_out[78][303],u_xpb_out[79][303],u_xpb_out[80][303],u_xpb_out[81][303],u_xpb_out[82][303],u_xpb_out[83][303],u_xpb_out[84][303],u_xpb_out[85][303],u_xpb_out[86][303],u_xpb_out[87][303],u_xpb_out[88][303],u_xpb_out[89][303],u_xpb_out[90][303],u_xpb_out[91][303],u_xpb_out[92][303],u_xpb_out[93][303],u_xpb_out[94][303],u_xpb_out[95][303],u_xpb_out[96][303],u_xpb_out[97][303],u_xpb_out[98][303],u_xpb_out[99][303],u_xpb_out[100][303],u_xpb_out[101][303],u_xpb_out[102][303],u_xpb_out[103][303],u_xpb_out[104][303],u_xpb_out[105][303]};

assign col_out_304 = {u_xpb_out[0][304],u_xpb_out[1][304],u_xpb_out[2][304],u_xpb_out[3][304],u_xpb_out[4][304],u_xpb_out[5][304],u_xpb_out[6][304],u_xpb_out[7][304],u_xpb_out[8][304],u_xpb_out[9][304],u_xpb_out[10][304],u_xpb_out[11][304],u_xpb_out[12][304],u_xpb_out[13][304],u_xpb_out[14][304],u_xpb_out[15][304],u_xpb_out[16][304],u_xpb_out[17][304],u_xpb_out[18][304],u_xpb_out[19][304],u_xpb_out[20][304],u_xpb_out[21][304],u_xpb_out[22][304],u_xpb_out[23][304],u_xpb_out[24][304],u_xpb_out[25][304],u_xpb_out[26][304],u_xpb_out[27][304],u_xpb_out[28][304],u_xpb_out[29][304],u_xpb_out[30][304],u_xpb_out[31][304],u_xpb_out[32][304],u_xpb_out[33][304],u_xpb_out[34][304],u_xpb_out[35][304],u_xpb_out[36][304],u_xpb_out[37][304],u_xpb_out[38][304],u_xpb_out[39][304],u_xpb_out[40][304],u_xpb_out[41][304],u_xpb_out[42][304],u_xpb_out[43][304],u_xpb_out[44][304],u_xpb_out[45][304],u_xpb_out[46][304],u_xpb_out[47][304],u_xpb_out[48][304],u_xpb_out[49][304],u_xpb_out[50][304],u_xpb_out[51][304],u_xpb_out[52][304],u_xpb_out[53][304],u_xpb_out[54][304],u_xpb_out[55][304],u_xpb_out[56][304],u_xpb_out[57][304],u_xpb_out[58][304],u_xpb_out[59][304],u_xpb_out[60][304],u_xpb_out[61][304],u_xpb_out[62][304],u_xpb_out[63][304],u_xpb_out[64][304],u_xpb_out[65][304],u_xpb_out[66][304],u_xpb_out[67][304],u_xpb_out[68][304],u_xpb_out[69][304],u_xpb_out[70][304],u_xpb_out[71][304],u_xpb_out[72][304],u_xpb_out[73][304],u_xpb_out[74][304],u_xpb_out[75][304],u_xpb_out[76][304],u_xpb_out[77][304],u_xpb_out[78][304],u_xpb_out[79][304],u_xpb_out[80][304],u_xpb_out[81][304],u_xpb_out[82][304],u_xpb_out[83][304],u_xpb_out[84][304],u_xpb_out[85][304],u_xpb_out[86][304],u_xpb_out[87][304],u_xpb_out[88][304],u_xpb_out[89][304],u_xpb_out[90][304],u_xpb_out[91][304],u_xpb_out[92][304],u_xpb_out[93][304],u_xpb_out[94][304],u_xpb_out[95][304],u_xpb_out[96][304],u_xpb_out[97][304],u_xpb_out[98][304],u_xpb_out[99][304],u_xpb_out[100][304],u_xpb_out[101][304],u_xpb_out[102][304],u_xpb_out[103][304],u_xpb_out[104][304],u_xpb_out[105][304]};

assign col_out_305 = {u_xpb_out[0][305],u_xpb_out[1][305],u_xpb_out[2][305],u_xpb_out[3][305],u_xpb_out[4][305],u_xpb_out[5][305],u_xpb_out[6][305],u_xpb_out[7][305],u_xpb_out[8][305],u_xpb_out[9][305],u_xpb_out[10][305],u_xpb_out[11][305],u_xpb_out[12][305],u_xpb_out[13][305],u_xpb_out[14][305],u_xpb_out[15][305],u_xpb_out[16][305],u_xpb_out[17][305],u_xpb_out[18][305],u_xpb_out[19][305],u_xpb_out[20][305],u_xpb_out[21][305],u_xpb_out[22][305],u_xpb_out[23][305],u_xpb_out[24][305],u_xpb_out[25][305],u_xpb_out[26][305],u_xpb_out[27][305],u_xpb_out[28][305],u_xpb_out[29][305],u_xpb_out[30][305],u_xpb_out[31][305],u_xpb_out[32][305],u_xpb_out[33][305],u_xpb_out[34][305],u_xpb_out[35][305],u_xpb_out[36][305],u_xpb_out[37][305],u_xpb_out[38][305],u_xpb_out[39][305],u_xpb_out[40][305],u_xpb_out[41][305],u_xpb_out[42][305],u_xpb_out[43][305],u_xpb_out[44][305],u_xpb_out[45][305],u_xpb_out[46][305],u_xpb_out[47][305],u_xpb_out[48][305],u_xpb_out[49][305],u_xpb_out[50][305],u_xpb_out[51][305],u_xpb_out[52][305],u_xpb_out[53][305],u_xpb_out[54][305],u_xpb_out[55][305],u_xpb_out[56][305],u_xpb_out[57][305],u_xpb_out[58][305],u_xpb_out[59][305],u_xpb_out[60][305],u_xpb_out[61][305],u_xpb_out[62][305],u_xpb_out[63][305],u_xpb_out[64][305],u_xpb_out[65][305],u_xpb_out[66][305],u_xpb_out[67][305],u_xpb_out[68][305],u_xpb_out[69][305],u_xpb_out[70][305],u_xpb_out[71][305],u_xpb_out[72][305],u_xpb_out[73][305],u_xpb_out[74][305],u_xpb_out[75][305],u_xpb_out[76][305],u_xpb_out[77][305],u_xpb_out[78][305],u_xpb_out[79][305],u_xpb_out[80][305],u_xpb_out[81][305],u_xpb_out[82][305],u_xpb_out[83][305],u_xpb_out[84][305],u_xpb_out[85][305],u_xpb_out[86][305],u_xpb_out[87][305],u_xpb_out[88][305],u_xpb_out[89][305],u_xpb_out[90][305],u_xpb_out[91][305],u_xpb_out[92][305],u_xpb_out[93][305],u_xpb_out[94][305],u_xpb_out[95][305],u_xpb_out[96][305],u_xpb_out[97][305],u_xpb_out[98][305],u_xpb_out[99][305],u_xpb_out[100][305],u_xpb_out[101][305],u_xpb_out[102][305],u_xpb_out[103][305],u_xpb_out[104][305],u_xpb_out[105][305]};

assign col_out_306 = {u_xpb_out[0][306],u_xpb_out[1][306],u_xpb_out[2][306],u_xpb_out[3][306],u_xpb_out[4][306],u_xpb_out[5][306],u_xpb_out[6][306],u_xpb_out[7][306],u_xpb_out[8][306],u_xpb_out[9][306],u_xpb_out[10][306],u_xpb_out[11][306],u_xpb_out[12][306],u_xpb_out[13][306],u_xpb_out[14][306],u_xpb_out[15][306],u_xpb_out[16][306],u_xpb_out[17][306],u_xpb_out[18][306],u_xpb_out[19][306],u_xpb_out[20][306],u_xpb_out[21][306],u_xpb_out[22][306],u_xpb_out[23][306],u_xpb_out[24][306],u_xpb_out[25][306],u_xpb_out[26][306],u_xpb_out[27][306],u_xpb_out[28][306],u_xpb_out[29][306],u_xpb_out[30][306],u_xpb_out[31][306],u_xpb_out[32][306],u_xpb_out[33][306],u_xpb_out[34][306],u_xpb_out[35][306],u_xpb_out[36][306],u_xpb_out[37][306],u_xpb_out[38][306],u_xpb_out[39][306],u_xpb_out[40][306],u_xpb_out[41][306],u_xpb_out[42][306],u_xpb_out[43][306],u_xpb_out[44][306],u_xpb_out[45][306],u_xpb_out[46][306],u_xpb_out[47][306],u_xpb_out[48][306],u_xpb_out[49][306],u_xpb_out[50][306],u_xpb_out[51][306],u_xpb_out[52][306],u_xpb_out[53][306],u_xpb_out[54][306],u_xpb_out[55][306],u_xpb_out[56][306],u_xpb_out[57][306],u_xpb_out[58][306],u_xpb_out[59][306],u_xpb_out[60][306],u_xpb_out[61][306],u_xpb_out[62][306],u_xpb_out[63][306],u_xpb_out[64][306],u_xpb_out[65][306],u_xpb_out[66][306],u_xpb_out[67][306],u_xpb_out[68][306],u_xpb_out[69][306],u_xpb_out[70][306],u_xpb_out[71][306],u_xpb_out[72][306],u_xpb_out[73][306],u_xpb_out[74][306],u_xpb_out[75][306],u_xpb_out[76][306],u_xpb_out[77][306],u_xpb_out[78][306],u_xpb_out[79][306],u_xpb_out[80][306],u_xpb_out[81][306],u_xpb_out[82][306],u_xpb_out[83][306],u_xpb_out[84][306],u_xpb_out[85][306],u_xpb_out[86][306],u_xpb_out[87][306],u_xpb_out[88][306],u_xpb_out[89][306],u_xpb_out[90][306],u_xpb_out[91][306],u_xpb_out[92][306],u_xpb_out[93][306],u_xpb_out[94][306],u_xpb_out[95][306],u_xpb_out[96][306],u_xpb_out[97][306],u_xpb_out[98][306],u_xpb_out[99][306],u_xpb_out[100][306],u_xpb_out[101][306],u_xpb_out[102][306],u_xpb_out[103][306],u_xpb_out[104][306],u_xpb_out[105][306]};

assign col_out_307 = {u_xpb_out[0][307],u_xpb_out[1][307],u_xpb_out[2][307],u_xpb_out[3][307],u_xpb_out[4][307],u_xpb_out[5][307],u_xpb_out[6][307],u_xpb_out[7][307],u_xpb_out[8][307],u_xpb_out[9][307],u_xpb_out[10][307],u_xpb_out[11][307],u_xpb_out[12][307],u_xpb_out[13][307],u_xpb_out[14][307],u_xpb_out[15][307],u_xpb_out[16][307],u_xpb_out[17][307],u_xpb_out[18][307],u_xpb_out[19][307],u_xpb_out[20][307],u_xpb_out[21][307],u_xpb_out[22][307],u_xpb_out[23][307],u_xpb_out[24][307],u_xpb_out[25][307],u_xpb_out[26][307],u_xpb_out[27][307],u_xpb_out[28][307],u_xpb_out[29][307],u_xpb_out[30][307],u_xpb_out[31][307],u_xpb_out[32][307],u_xpb_out[33][307],u_xpb_out[34][307],u_xpb_out[35][307],u_xpb_out[36][307],u_xpb_out[37][307],u_xpb_out[38][307],u_xpb_out[39][307],u_xpb_out[40][307],u_xpb_out[41][307],u_xpb_out[42][307],u_xpb_out[43][307],u_xpb_out[44][307],u_xpb_out[45][307],u_xpb_out[46][307],u_xpb_out[47][307],u_xpb_out[48][307],u_xpb_out[49][307],u_xpb_out[50][307],u_xpb_out[51][307],u_xpb_out[52][307],u_xpb_out[53][307],u_xpb_out[54][307],u_xpb_out[55][307],u_xpb_out[56][307],u_xpb_out[57][307],u_xpb_out[58][307],u_xpb_out[59][307],u_xpb_out[60][307],u_xpb_out[61][307],u_xpb_out[62][307],u_xpb_out[63][307],u_xpb_out[64][307],u_xpb_out[65][307],u_xpb_out[66][307],u_xpb_out[67][307],u_xpb_out[68][307],u_xpb_out[69][307],u_xpb_out[70][307],u_xpb_out[71][307],u_xpb_out[72][307],u_xpb_out[73][307],u_xpb_out[74][307],u_xpb_out[75][307],u_xpb_out[76][307],u_xpb_out[77][307],u_xpb_out[78][307],u_xpb_out[79][307],u_xpb_out[80][307],u_xpb_out[81][307],u_xpb_out[82][307],u_xpb_out[83][307],u_xpb_out[84][307],u_xpb_out[85][307],u_xpb_out[86][307],u_xpb_out[87][307],u_xpb_out[88][307],u_xpb_out[89][307],u_xpb_out[90][307],u_xpb_out[91][307],u_xpb_out[92][307],u_xpb_out[93][307],u_xpb_out[94][307],u_xpb_out[95][307],u_xpb_out[96][307],u_xpb_out[97][307],u_xpb_out[98][307],u_xpb_out[99][307],u_xpb_out[100][307],u_xpb_out[101][307],u_xpb_out[102][307],u_xpb_out[103][307],u_xpb_out[104][307],u_xpb_out[105][307]};

assign col_out_308 = {u_xpb_out[0][308],u_xpb_out[1][308],u_xpb_out[2][308],u_xpb_out[3][308],u_xpb_out[4][308],u_xpb_out[5][308],u_xpb_out[6][308],u_xpb_out[7][308],u_xpb_out[8][308],u_xpb_out[9][308],u_xpb_out[10][308],u_xpb_out[11][308],u_xpb_out[12][308],u_xpb_out[13][308],u_xpb_out[14][308],u_xpb_out[15][308],u_xpb_out[16][308],u_xpb_out[17][308],u_xpb_out[18][308],u_xpb_out[19][308],u_xpb_out[20][308],u_xpb_out[21][308],u_xpb_out[22][308],u_xpb_out[23][308],u_xpb_out[24][308],u_xpb_out[25][308],u_xpb_out[26][308],u_xpb_out[27][308],u_xpb_out[28][308],u_xpb_out[29][308],u_xpb_out[30][308],u_xpb_out[31][308],u_xpb_out[32][308],u_xpb_out[33][308],u_xpb_out[34][308],u_xpb_out[35][308],u_xpb_out[36][308],u_xpb_out[37][308],u_xpb_out[38][308],u_xpb_out[39][308],u_xpb_out[40][308],u_xpb_out[41][308],u_xpb_out[42][308],u_xpb_out[43][308],u_xpb_out[44][308],u_xpb_out[45][308],u_xpb_out[46][308],u_xpb_out[47][308],u_xpb_out[48][308],u_xpb_out[49][308],u_xpb_out[50][308],u_xpb_out[51][308],u_xpb_out[52][308],u_xpb_out[53][308],u_xpb_out[54][308],u_xpb_out[55][308],u_xpb_out[56][308],u_xpb_out[57][308],u_xpb_out[58][308],u_xpb_out[59][308],u_xpb_out[60][308],u_xpb_out[61][308],u_xpb_out[62][308],u_xpb_out[63][308],u_xpb_out[64][308],u_xpb_out[65][308],u_xpb_out[66][308],u_xpb_out[67][308],u_xpb_out[68][308],u_xpb_out[69][308],u_xpb_out[70][308],u_xpb_out[71][308],u_xpb_out[72][308],u_xpb_out[73][308],u_xpb_out[74][308],u_xpb_out[75][308],u_xpb_out[76][308],u_xpb_out[77][308],u_xpb_out[78][308],u_xpb_out[79][308],u_xpb_out[80][308],u_xpb_out[81][308],u_xpb_out[82][308],u_xpb_out[83][308],u_xpb_out[84][308],u_xpb_out[85][308],u_xpb_out[86][308],u_xpb_out[87][308],u_xpb_out[88][308],u_xpb_out[89][308],u_xpb_out[90][308],u_xpb_out[91][308],u_xpb_out[92][308],u_xpb_out[93][308],u_xpb_out[94][308],u_xpb_out[95][308],u_xpb_out[96][308],u_xpb_out[97][308],u_xpb_out[98][308],u_xpb_out[99][308],u_xpb_out[100][308],u_xpb_out[101][308],u_xpb_out[102][308],u_xpb_out[103][308],u_xpb_out[104][308],u_xpb_out[105][308]};

assign col_out_309 = {u_xpb_out[0][309],u_xpb_out[1][309],u_xpb_out[2][309],u_xpb_out[3][309],u_xpb_out[4][309],u_xpb_out[5][309],u_xpb_out[6][309],u_xpb_out[7][309],u_xpb_out[8][309],u_xpb_out[9][309],u_xpb_out[10][309],u_xpb_out[11][309],u_xpb_out[12][309],u_xpb_out[13][309],u_xpb_out[14][309],u_xpb_out[15][309],u_xpb_out[16][309],u_xpb_out[17][309],u_xpb_out[18][309],u_xpb_out[19][309],u_xpb_out[20][309],u_xpb_out[21][309],u_xpb_out[22][309],u_xpb_out[23][309],u_xpb_out[24][309],u_xpb_out[25][309],u_xpb_out[26][309],u_xpb_out[27][309],u_xpb_out[28][309],u_xpb_out[29][309],u_xpb_out[30][309],u_xpb_out[31][309],u_xpb_out[32][309],u_xpb_out[33][309],u_xpb_out[34][309],u_xpb_out[35][309],u_xpb_out[36][309],u_xpb_out[37][309],u_xpb_out[38][309],u_xpb_out[39][309],u_xpb_out[40][309],u_xpb_out[41][309],u_xpb_out[42][309],u_xpb_out[43][309],u_xpb_out[44][309],u_xpb_out[45][309],u_xpb_out[46][309],u_xpb_out[47][309],u_xpb_out[48][309],u_xpb_out[49][309],u_xpb_out[50][309],u_xpb_out[51][309],u_xpb_out[52][309],u_xpb_out[53][309],u_xpb_out[54][309],u_xpb_out[55][309],u_xpb_out[56][309],u_xpb_out[57][309],u_xpb_out[58][309],u_xpb_out[59][309],u_xpb_out[60][309],u_xpb_out[61][309],u_xpb_out[62][309],u_xpb_out[63][309],u_xpb_out[64][309],u_xpb_out[65][309],u_xpb_out[66][309],u_xpb_out[67][309],u_xpb_out[68][309],u_xpb_out[69][309],u_xpb_out[70][309],u_xpb_out[71][309],u_xpb_out[72][309],u_xpb_out[73][309],u_xpb_out[74][309],u_xpb_out[75][309],u_xpb_out[76][309],u_xpb_out[77][309],u_xpb_out[78][309],u_xpb_out[79][309],u_xpb_out[80][309],u_xpb_out[81][309],u_xpb_out[82][309],u_xpb_out[83][309],u_xpb_out[84][309],u_xpb_out[85][309],u_xpb_out[86][309],u_xpb_out[87][309],u_xpb_out[88][309],u_xpb_out[89][309],u_xpb_out[90][309],u_xpb_out[91][309],u_xpb_out[92][309],u_xpb_out[93][309],u_xpb_out[94][309],u_xpb_out[95][309],u_xpb_out[96][309],u_xpb_out[97][309],u_xpb_out[98][309],u_xpb_out[99][309],u_xpb_out[100][309],u_xpb_out[101][309],u_xpb_out[102][309],u_xpb_out[103][309],u_xpb_out[104][309],u_xpb_out[105][309]};

assign col_out_310 = {u_xpb_out[0][310],u_xpb_out[1][310],u_xpb_out[2][310],u_xpb_out[3][310],u_xpb_out[4][310],u_xpb_out[5][310],u_xpb_out[6][310],u_xpb_out[7][310],u_xpb_out[8][310],u_xpb_out[9][310],u_xpb_out[10][310],u_xpb_out[11][310],u_xpb_out[12][310],u_xpb_out[13][310],u_xpb_out[14][310],u_xpb_out[15][310],u_xpb_out[16][310],u_xpb_out[17][310],u_xpb_out[18][310],u_xpb_out[19][310],u_xpb_out[20][310],u_xpb_out[21][310],u_xpb_out[22][310],u_xpb_out[23][310],u_xpb_out[24][310],u_xpb_out[25][310],u_xpb_out[26][310],u_xpb_out[27][310],u_xpb_out[28][310],u_xpb_out[29][310],u_xpb_out[30][310],u_xpb_out[31][310],u_xpb_out[32][310],u_xpb_out[33][310],u_xpb_out[34][310],u_xpb_out[35][310],u_xpb_out[36][310],u_xpb_out[37][310],u_xpb_out[38][310],u_xpb_out[39][310],u_xpb_out[40][310],u_xpb_out[41][310],u_xpb_out[42][310],u_xpb_out[43][310],u_xpb_out[44][310],u_xpb_out[45][310],u_xpb_out[46][310],u_xpb_out[47][310],u_xpb_out[48][310],u_xpb_out[49][310],u_xpb_out[50][310],u_xpb_out[51][310],u_xpb_out[52][310],u_xpb_out[53][310],u_xpb_out[54][310],u_xpb_out[55][310],u_xpb_out[56][310],u_xpb_out[57][310],u_xpb_out[58][310],u_xpb_out[59][310],u_xpb_out[60][310],u_xpb_out[61][310],u_xpb_out[62][310],u_xpb_out[63][310],u_xpb_out[64][310],u_xpb_out[65][310],u_xpb_out[66][310],u_xpb_out[67][310],u_xpb_out[68][310],u_xpb_out[69][310],u_xpb_out[70][310],u_xpb_out[71][310],u_xpb_out[72][310],u_xpb_out[73][310],u_xpb_out[74][310],u_xpb_out[75][310],u_xpb_out[76][310],u_xpb_out[77][310],u_xpb_out[78][310],u_xpb_out[79][310],u_xpb_out[80][310],u_xpb_out[81][310],u_xpb_out[82][310],u_xpb_out[83][310],u_xpb_out[84][310],u_xpb_out[85][310],u_xpb_out[86][310],u_xpb_out[87][310],u_xpb_out[88][310],u_xpb_out[89][310],u_xpb_out[90][310],u_xpb_out[91][310],u_xpb_out[92][310],u_xpb_out[93][310],u_xpb_out[94][310],u_xpb_out[95][310],u_xpb_out[96][310],u_xpb_out[97][310],u_xpb_out[98][310],u_xpb_out[99][310],u_xpb_out[100][310],u_xpb_out[101][310],u_xpb_out[102][310],u_xpb_out[103][310],u_xpb_out[104][310],u_xpb_out[105][310]};

assign col_out_311 = {u_xpb_out[0][311],u_xpb_out[1][311],u_xpb_out[2][311],u_xpb_out[3][311],u_xpb_out[4][311],u_xpb_out[5][311],u_xpb_out[6][311],u_xpb_out[7][311],u_xpb_out[8][311],u_xpb_out[9][311],u_xpb_out[10][311],u_xpb_out[11][311],u_xpb_out[12][311],u_xpb_out[13][311],u_xpb_out[14][311],u_xpb_out[15][311],u_xpb_out[16][311],u_xpb_out[17][311],u_xpb_out[18][311],u_xpb_out[19][311],u_xpb_out[20][311],u_xpb_out[21][311],u_xpb_out[22][311],u_xpb_out[23][311],u_xpb_out[24][311],u_xpb_out[25][311],u_xpb_out[26][311],u_xpb_out[27][311],u_xpb_out[28][311],u_xpb_out[29][311],u_xpb_out[30][311],u_xpb_out[31][311],u_xpb_out[32][311],u_xpb_out[33][311],u_xpb_out[34][311],u_xpb_out[35][311],u_xpb_out[36][311],u_xpb_out[37][311],u_xpb_out[38][311],u_xpb_out[39][311],u_xpb_out[40][311],u_xpb_out[41][311],u_xpb_out[42][311],u_xpb_out[43][311],u_xpb_out[44][311],u_xpb_out[45][311],u_xpb_out[46][311],u_xpb_out[47][311],u_xpb_out[48][311],u_xpb_out[49][311],u_xpb_out[50][311],u_xpb_out[51][311],u_xpb_out[52][311],u_xpb_out[53][311],u_xpb_out[54][311],u_xpb_out[55][311],u_xpb_out[56][311],u_xpb_out[57][311],u_xpb_out[58][311],u_xpb_out[59][311],u_xpb_out[60][311],u_xpb_out[61][311],u_xpb_out[62][311],u_xpb_out[63][311],u_xpb_out[64][311],u_xpb_out[65][311],u_xpb_out[66][311],u_xpb_out[67][311],u_xpb_out[68][311],u_xpb_out[69][311],u_xpb_out[70][311],u_xpb_out[71][311],u_xpb_out[72][311],u_xpb_out[73][311],u_xpb_out[74][311],u_xpb_out[75][311],u_xpb_out[76][311],u_xpb_out[77][311],u_xpb_out[78][311],u_xpb_out[79][311],u_xpb_out[80][311],u_xpb_out[81][311],u_xpb_out[82][311],u_xpb_out[83][311],u_xpb_out[84][311],u_xpb_out[85][311],u_xpb_out[86][311],u_xpb_out[87][311],u_xpb_out[88][311],u_xpb_out[89][311],u_xpb_out[90][311],u_xpb_out[91][311],u_xpb_out[92][311],u_xpb_out[93][311],u_xpb_out[94][311],u_xpb_out[95][311],u_xpb_out[96][311],u_xpb_out[97][311],u_xpb_out[98][311],u_xpb_out[99][311],u_xpb_out[100][311],u_xpb_out[101][311],u_xpb_out[102][311],u_xpb_out[103][311],u_xpb_out[104][311],u_xpb_out[105][311]};

assign col_out_312 = {u_xpb_out[0][312],u_xpb_out[1][312],u_xpb_out[2][312],u_xpb_out[3][312],u_xpb_out[4][312],u_xpb_out[5][312],u_xpb_out[6][312],u_xpb_out[7][312],u_xpb_out[8][312],u_xpb_out[9][312],u_xpb_out[10][312],u_xpb_out[11][312],u_xpb_out[12][312],u_xpb_out[13][312],u_xpb_out[14][312],u_xpb_out[15][312],u_xpb_out[16][312],u_xpb_out[17][312],u_xpb_out[18][312],u_xpb_out[19][312],u_xpb_out[20][312],u_xpb_out[21][312],u_xpb_out[22][312],u_xpb_out[23][312],u_xpb_out[24][312],u_xpb_out[25][312],u_xpb_out[26][312],u_xpb_out[27][312],u_xpb_out[28][312],u_xpb_out[29][312],u_xpb_out[30][312],u_xpb_out[31][312],u_xpb_out[32][312],u_xpb_out[33][312],u_xpb_out[34][312],u_xpb_out[35][312],u_xpb_out[36][312],u_xpb_out[37][312],u_xpb_out[38][312],u_xpb_out[39][312],u_xpb_out[40][312],u_xpb_out[41][312],u_xpb_out[42][312],u_xpb_out[43][312],u_xpb_out[44][312],u_xpb_out[45][312],u_xpb_out[46][312],u_xpb_out[47][312],u_xpb_out[48][312],u_xpb_out[49][312],u_xpb_out[50][312],u_xpb_out[51][312],u_xpb_out[52][312],u_xpb_out[53][312],u_xpb_out[54][312],u_xpb_out[55][312],u_xpb_out[56][312],u_xpb_out[57][312],u_xpb_out[58][312],u_xpb_out[59][312],u_xpb_out[60][312],u_xpb_out[61][312],u_xpb_out[62][312],u_xpb_out[63][312],u_xpb_out[64][312],u_xpb_out[65][312],u_xpb_out[66][312],u_xpb_out[67][312],u_xpb_out[68][312],u_xpb_out[69][312],u_xpb_out[70][312],u_xpb_out[71][312],u_xpb_out[72][312],u_xpb_out[73][312],u_xpb_out[74][312],u_xpb_out[75][312],u_xpb_out[76][312],u_xpb_out[77][312],u_xpb_out[78][312],u_xpb_out[79][312],u_xpb_out[80][312],u_xpb_out[81][312],u_xpb_out[82][312],u_xpb_out[83][312],u_xpb_out[84][312],u_xpb_out[85][312],u_xpb_out[86][312],u_xpb_out[87][312],u_xpb_out[88][312],u_xpb_out[89][312],u_xpb_out[90][312],u_xpb_out[91][312],u_xpb_out[92][312],u_xpb_out[93][312],u_xpb_out[94][312],u_xpb_out[95][312],u_xpb_out[96][312],u_xpb_out[97][312],u_xpb_out[98][312],u_xpb_out[99][312],u_xpb_out[100][312],u_xpb_out[101][312],u_xpb_out[102][312],u_xpb_out[103][312],u_xpb_out[104][312],u_xpb_out[105][312]};

assign col_out_313 = {u_xpb_out[0][313],u_xpb_out[1][313],u_xpb_out[2][313],u_xpb_out[3][313],u_xpb_out[4][313],u_xpb_out[5][313],u_xpb_out[6][313],u_xpb_out[7][313],u_xpb_out[8][313],u_xpb_out[9][313],u_xpb_out[10][313],u_xpb_out[11][313],u_xpb_out[12][313],u_xpb_out[13][313],u_xpb_out[14][313],u_xpb_out[15][313],u_xpb_out[16][313],u_xpb_out[17][313],u_xpb_out[18][313],u_xpb_out[19][313],u_xpb_out[20][313],u_xpb_out[21][313],u_xpb_out[22][313],u_xpb_out[23][313],u_xpb_out[24][313],u_xpb_out[25][313],u_xpb_out[26][313],u_xpb_out[27][313],u_xpb_out[28][313],u_xpb_out[29][313],u_xpb_out[30][313],u_xpb_out[31][313],u_xpb_out[32][313],u_xpb_out[33][313],u_xpb_out[34][313],u_xpb_out[35][313],u_xpb_out[36][313],u_xpb_out[37][313],u_xpb_out[38][313],u_xpb_out[39][313],u_xpb_out[40][313],u_xpb_out[41][313],u_xpb_out[42][313],u_xpb_out[43][313],u_xpb_out[44][313],u_xpb_out[45][313],u_xpb_out[46][313],u_xpb_out[47][313],u_xpb_out[48][313],u_xpb_out[49][313],u_xpb_out[50][313],u_xpb_out[51][313],u_xpb_out[52][313],u_xpb_out[53][313],u_xpb_out[54][313],u_xpb_out[55][313],u_xpb_out[56][313],u_xpb_out[57][313],u_xpb_out[58][313],u_xpb_out[59][313],u_xpb_out[60][313],u_xpb_out[61][313],u_xpb_out[62][313],u_xpb_out[63][313],u_xpb_out[64][313],u_xpb_out[65][313],u_xpb_out[66][313],u_xpb_out[67][313],u_xpb_out[68][313],u_xpb_out[69][313],u_xpb_out[70][313],u_xpb_out[71][313],u_xpb_out[72][313],u_xpb_out[73][313],u_xpb_out[74][313],u_xpb_out[75][313],u_xpb_out[76][313],u_xpb_out[77][313],u_xpb_out[78][313],u_xpb_out[79][313],u_xpb_out[80][313],u_xpb_out[81][313],u_xpb_out[82][313],u_xpb_out[83][313],u_xpb_out[84][313],u_xpb_out[85][313],u_xpb_out[86][313],u_xpb_out[87][313],u_xpb_out[88][313],u_xpb_out[89][313],u_xpb_out[90][313],u_xpb_out[91][313],u_xpb_out[92][313],u_xpb_out[93][313],u_xpb_out[94][313],u_xpb_out[95][313],u_xpb_out[96][313],u_xpb_out[97][313],u_xpb_out[98][313],u_xpb_out[99][313],u_xpb_out[100][313],u_xpb_out[101][313],u_xpb_out[102][313],u_xpb_out[103][313],u_xpb_out[104][313],u_xpb_out[105][313]};

assign col_out_314 = {u_xpb_out[0][314],u_xpb_out[1][314],u_xpb_out[2][314],u_xpb_out[3][314],u_xpb_out[4][314],u_xpb_out[5][314],u_xpb_out[6][314],u_xpb_out[7][314],u_xpb_out[8][314],u_xpb_out[9][314],u_xpb_out[10][314],u_xpb_out[11][314],u_xpb_out[12][314],u_xpb_out[13][314],u_xpb_out[14][314],u_xpb_out[15][314],u_xpb_out[16][314],u_xpb_out[17][314],u_xpb_out[18][314],u_xpb_out[19][314],u_xpb_out[20][314],u_xpb_out[21][314],u_xpb_out[22][314],u_xpb_out[23][314],u_xpb_out[24][314],u_xpb_out[25][314],u_xpb_out[26][314],u_xpb_out[27][314],u_xpb_out[28][314],u_xpb_out[29][314],u_xpb_out[30][314],u_xpb_out[31][314],u_xpb_out[32][314],u_xpb_out[33][314],u_xpb_out[34][314],u_xpb_out[35][314],u_xpb_out[36][314],u_xpb_out[37][314],u_xpb_out[38][314],u_xpb_out[39][314],u_xpb_out[40][314],u_xpb_out[41][314],u_xpb_out[42][314],u_xpb_out[43][314],u_xpb_out[44][314],u_xpb_out[45][314],u_xpb_out[46][314],u_xpb_out[47][314],u_xpb_out[48][314],u_xpb_out[49][314],u_xpb_out[50][314],u_xpb_out[51][314],u_xpb_out[52][314],u_xpb_out[53][314],u_xpb_out[54][314],u_xpb_out[55][314],u_xpb_out[56][314],u_xpb_out[57][314],u_xpb_out[58][314],u_xpb_out[59][314],u_xpb_out[60][314],u_xpb_out[61][314],u_xpb_out[62][314],u_xpb_out[63][314],u_xpb_out[64][314],u_xpb_out[65][314],u_xpb_out[66][314],u_xpb_out[67][314],u_xpb_out[68][314],u_xpb_out[69][314],u_xpb_out[70][314],u_xpb_out[71][314],u_xpb_out[72][314],u_xpb_out[73][314],u_xpb_out[74][314],u_xpb_out[75][314],u_xpb_out[76][314],u_xpb_out[77][314],u_xpb_out[78][314],u_xpb_out[79][314],u_xpb_out[80][314],u_xpb_out[81][314],u_xpb_out[82][314],u_xpb_out[83][314],u_xpb_out[84][314],u_xpb_out[85][314],u_xpb_out[86][314],u_xpb_out[87][314],u_xpb_out[88][314],u_xpb_out[89][314],u_xpb_out[90][314],u_xpb_out[91][314],u_xpb_out[92][314],u_xpb_out[93][314],u_xpb_out[94][314],u_xpb_out[95][314],u_xpb_out[96][314],u_xpb_out[97][314],u_xpb_out[98][314],u_xpb_out[99][314],u_xpb_out[100][314],u_xpb_out[101][314],u_xpb_out[102][314],u_xpb_out[103][314],u_xpb_out[104][314],u_xpb_out[105][314]};

assign col_out_315 = {u_xpb_out[0][315],u_xpb_out[1][315],u_xpb_out[2][315],u_xpb_out[3][315],u_xpb_out[4][315],u_xpb_out[5][315],u_xpb_out[6][315],u_xpb_out[7][315],u_xpb_out[8][315],u_xpb_out[9][315],u_xpb_out[10][315],u_xpb_out[11][315],u_xpb_out[12][315],u_xpb_out[13][315],u_xpb_out[14][315],u_xpb_out[15][315],u_xpb_out[16][315],u_xpb_out[17][315],u_xpb_out[18][315],u_xpb_out[19][315],u_xpb_out[20][315],u_xpb_out[21][315],u_xpb_out[22][315],u_xpb_out[23][315],u_xpb_out[24][315],u_xpb_out[25][315],u_xpb_out[26][315],u_xpb_out[27][315],u_xpb_out[28][315],u_xpb_out[29][315],u_xpb_out[30][315],u_xpb_out[31][315],u_xpb_out[32][315],u_xpb_out[33][315],u_xpb_out[34][315],u_xpb_out[35][315],u_xpb_out[36][315],u_xpb_out[37][315],u_xpb_out[38][315],u_xpb_out[39][315],u_xpb_out[40][315],u_xpb_out[41][315],u_xpb_out[42][315],u_xpb_out[43][315],u_xpb_out[44][315],u_xpb_out[45][315],u_xpb_out[46][315],u_xpb_out[47][315],u_xpb_out[48][315],u_xpb_out[49][315],u_xpb_out[50][315],u_xpb_out[51][315],u_xpb_out[52][315],u_xpb_out[53][315],u_xpb_out[54][315],u_xpb_out[55][315],u_xpb_out[56][315],u_xpb_out[57][315],u_xpb_out[58][315],u_xpb_out[59][315],u_xpb_out[60][315],u_xpb_out[61][315],u_xpb_out[62][315],u_xpb_out[63][315],u_xpb_out[64][315],u_xpb_out[65][315],u_xpb_out[66][315],u_xpb_out[67][315],u_xpb_out[68][315],u_xpb_out[69][315],u_xpb_out[70][315],u_xpb_out[71][315],u_xpb_out[72][315],u_xpb_out[73][315],u_xpb_out[74][315],u_xpb_out[75][315],u_xpb_out[76][315],u_xpb_out[77][315],u_xpb_out[78][315],u_xpb_out[79][315],u_xpb_out[80][315],u_xpb_out[81][315],u_xpb_out[82][315],u_xpb_out[83][315],u_xpb_out[84][315],u_xpb_out[85][315],u_xpb_out[86][315],u_xpb_out[87][315],u_xpb_out[88][315],u_xpb_out[89][315],u_xpb_out[90][315],u_xpb_out[91][315],u_xpb_out[92][315],u_xpb_out[93][315],u_xpb_out[94][315],u_xpb_out[95][315],u_xpb_out[96][315],u_xpb_out[97][315],u_xpb_out[98][315],u_xpb_out[99][315],u_xpb_out[100][315],u_xpb_out[101][315],u_xpb_out[102][315],u_xpb_out[103][315],u_xpb_out[104][315],u_xpb_out[105][315]};

assign col_out_316 = {u_xpb_out[0][316],u_xpb_out[1][316],u_xpb_out[2][316],u_xpb_out[3][316],u_xpb_out[4][316],u_xpb_out[5][316],u_xpb_out[6][316],u_xpb_out[7][316],u_xpb_out[8][316],u_xpb_out[9][316],u_xpb_out[10][316],u_xpb_out[11][316],u_xpb_out[12][316],u_xpb_out[13][316],u_xpb_out[14][316],u_xpb_out[15][316],u_xpb_out[16][316],u_xpb_out[17][316],u_xpb_out[18][316],u_xpb_out[19][316],u_xpb_out[20][316],u_xpb_out[21][316],u_xpb_out[22][316],u_xpb_out[23][316],u_xpb_out[24][316],u_xpb_out[25][316],u_xpb_out[26][316],u_xpb_out[27][316],u_xpb_out[28][316],u_xpb_out[29][316],u_xpb_out[30][316],u_xpb_out[31][316],u_xpb_out[32][316],u_xpb_out[33][316],u_xpb_out[34][316],u_xpb_out[35][316],u_xpb_out[36][316],u_xpb_out[37][316],u_xpb_out[38][316],u_xpb_out[39][316],u_xpb_out[40][316],u_xpb_out[41][316],u_xpb_out[42][316],u_xpb_out[43][316],u_xpb_out[44][316],u_xpb_out[45][316],u_xpb_out[46][316],u_xpb_out[47][316],u_xpb_out[48][316],u_xpb_out[49][316],u_xpb_out[50][316],u_xpb_out[51][316],u_xpb_out[52][316],u_xpb_out[53][316],u_xpb_out[54][316],u_xpb_out[55][316],u_xpb_out[56][316],u_xpb_out[57][316],u_xpb_out[58][316],u_xpb_out[59][316],u_xpb_out[60][316],u_xpb_out[61][316],u_xpb_out[62][316],u_xpb_out[63][316],u_xpb_out[64][316],u_xpb_out[65][316],u_xpb_out[66][316],u_xpb_out[67][316],u_xpb_out[68][316],u_xpb_out[69][316],u_xpb_out[70][316],u_xpb_out[71][316],u_xpb_out[72][316],u_xpb_out[73][316],u_xpb_out[74][316],u_xpb_out[75][316],u_xpb_out[76][316],u_xpb_out[77][316],u_xpb_out[78][316],u_xpb_out[79][316],u_xpb_out[80][316],u_xpb_out[81][316],u_xpb_out[82][316],u_xpb_out[83][316],u_xpb_out[84][316],u_xpb_out[85][316],u_xpb_out[86][316],u_xpb_out[87][316],u_xpb_out[88][316],u_xpb_out[89][316],u_xpb_out[90][316],u_xpb_out[91][316],u_xpb_out[92][316],u_xpb_out[93][316],u_xpb_out[94][316],u_xpb_out[95][316],u_xpb_out[96][316],u_xpb_out[97][316],u_xpb_out[98][316],u_xpb_out[99][316],u_xpb_out[100][316],u_xpb_out[101][316],u_xpb_out[102][316],u_xpb_out[103][316],u_xpb_out[104][316],u_xpb_out[105][316]};

assign col_out_317 = {u_xpb_out[0][317],u_xpb_out[1][317],u_xpb_out[2][317],u_xpb_out[3][317],u_xpb_out[4][317],u_xpb_out[5][317],u_xpb_out[6][317],u_xpb_out[7][317],u_xpb_out[8][317],u_xpb_out[9][317],u_xpb_out[10][317],u_xpb_out[11][317],u_xpb_out[12][317],u_xpb_out[13][317],u_xpb_out[14][317],u_xpb_out[15][317],u_xpb_out[16][317],u_xpb_out[17][317],u_xpb_out[18][317],u_xpb_out[19][317],u_xpb_out[20][317],u_xpb_out[21][317],u_xpb_out[22][317],u_xpb_out[23][317],u_xpb_out[24][317],u_xpb_out[25][317],u_xpb_out[26][317],u_xpb_out[27][317],u_xpb_out[28][317],u_xpb_out[29][317],u_xpb_out[30][317],u_xpb_out[31][317],u_xpb_out[32][317],u_xpb_out[33][317],u_xpb_out[34][317],u_xpb_out[35][317],u_xpb_out[36][317],u_xpb_out[37][317],u_xpb_out[38][317],u_xpb_out[39][317],u_xpb_out[40][317],u_xpb_out[41][317],u_xpb_out[42][317],u_xpb_out[43][317],u_xpb_out[44][317],u_xpb_out[45][317],u_xpb_out[46][317],u_xpb_out[47][317],u_xpb_out[48][317],u_xpb_out[49][317],u_xpb_out[50][317],u_xpb_out[51][317],u_xpb_out[52][317],u_xpb_out[53][317],u_xpb_out[54][317],u_xpb_out[55][317],u_xpb_out[56][317],u_xpb_out[57][317],u_xpb_out[58][317],u_xpb_out[59][317],u_xpb_out[60][317],u_xpb_out[61][317],u_xpb_out[62][317],u_xpb_out[63][317],u_xpb_out[64][317],u_xpb_out[65][317],u_xpb_out[66][317],u_xpb_out[67][317],u_xpb_out[68][317],u_xpb_out[69][317],u_xpb_out[70][317],u_xpb_out[71][317],u_xpb_out[72][317],u_xpb_out[73][317],u_xpb_out[74][317],u_xpb_out[75][317],u_xpb_out[76][317],u_xpb_out[77][317],u_xpb_out[78][317],u_xpb_out[79][317],u_xpb_out[80][317],u_xpb_out[81][317],u_xpb_out[82][317],u_xpb_out[83][317],u_xpb_out[84][317],u_xpb_out[85][317],u_xpb_out[86][317],u_xpb_out[87][317],u_xpb_out[88][317],u_xpb_out[89][317],u_xpb_out[90][317],u_xpb_out[91][317],u_xpb_out[92][317],u_xpb_out[93][317],u_xpb_out[94][317],u_xpb_out[95][317],u_xpb_out[96][317],u_xpb_out[97][317],u_xpb_out[98][317],u_xpb_out[99][317],u_xpb_out[100][317],u_xpb_out[101][317],u_xpb_out[102][317],u_xpb_out[103][317],u_xpb_out[104][317],u_xpb_out[105][317]};

assign col_out_318 = {u_xpb_out[0][318],u_xpb_out[1][318],u_xpb_out[2][318],u_xpb_out[3][318],u_xpb_out[4][318],u_xpb_out[5][318],u_xpb_out[6][318],u_xpb_out[7][318],u_xpb_out[8][318],u_xpb_out[9][318],u_xpb_out[10][318],u_xpb_out[11][318],u_xpb_out[12][318],u_xpb_out[13][318],u_xpb_out[14][318],u_xpb_out[15][318],u_xpb_out[16][318],u_xpb_out[17][318],u_xpb_out[18][318],u_xpb_out[19][318],u_xpb_out[20][318],u_xpb_out[21][318],u_xpb_out[22][318],u_xpb_out[23][318],u_xpb_out[24][318],u_xpb_out[25][318],u_xpb_out[26][318],u_xpb_out[27][318],u_xpb_out[28][318],u_xpb_out[29][318],u_xpb_out[30][318],u_xpb_out[31][318],u_xpb_out[32][318],u_xpb_out[33][318],u_xpb_out[34][318],u_xpb_out[35][318],u_xpb_out[36][318],u_xpb_out[37][318],u_xpb_out[38][318],u_xpb_out[39][318],u_xpb_out[40][318],u_xpb_out[41][318],u_xpb_out[42][318],u_xpb_out[43][318],u_xpb_out[44][318],u_xpb_out[45][318],u_xpb_out[46][318],u_xpb_out[47][318],u_xpb_out[48][318],u_xpb_out[49][318],u_xpb_out[50][318],u_xpb_out[51][318],u_xpb_out[52][318],u_xpb_out[53][318],u_xpb_out[54][318],u_xpb_out[55][318],u_xpb_out[56][318],u_xpb_out[57][318],u_xpb_out[58][318],u_xpb_out[59][318],u_xpb_out[60][318],u_xpb_out[61][318],u_xpb_out[62][318],u_xpb_out[63][318],u_xpb_out[64][318],u_xpb_out[65][318],u_xpb_out[66][318],u_xpb_out[67][318],u_xpb_out[68][318],u_xpb_out[69][318],u_xpb_out[70][318],u_xpb_out[71][318],u_xpb_out[72][318],u_xpb_out[73][318],u_xpb_out[74][318],u_xpb_out[75][318],u_xpb_out[76][318],u_xpb_out[77][318],u_xpb_out[78][318],u_xpb_out[79][318],u_xpb_out[80][318],u_xpb_out[81][318],u_xpb_out[82][318],u_xpb_out[83][318],u_xpb_out[84][318],u_xpb_out[85][318],u_xpb_out[86][318],u_xpb_out[87][318],u_xpb_out[88][318],u_xpb_out[89][318],u_xpb_out[90][318],u_xpb_out[91][318],u_xpb_out[92][318],u_xpb_out[93][318],u_xpb_out[94][318],u_xpb_out[95][318],u_xpb_out[96][318],u_xpb_out[97][318],u_xpb_out[98][318],u_xpb_out[99][318],u_xpb_out[100][318],u_xpb_out[101][318],u_xpb_out[102][318],u_xpb_out[103][318],u_xpb_out[104][318],u_xpb_out[105][318]};

assign col_out_319 = {u_xpb_out[0][319],u_xpb_out[1][319],u_xpb_out[2][319],u_xpb_out[3][319],u_xpb_out[4][319],u_xpb_out[5][319],u_xpb_out[6][319],u_xpb_out[7][319],u_xpb_out[8][319],u_xpb_out[9][319],u_xpb_out[10][319],u_xpb_out[11][319],u_xpb_out[12][319],u_xpb_out[13][319],u_xpb_out[14][319],u_xpb_out[15][319],u_xpb_out[16][319],u_xpb_out[17][319],u_xpb_out[18][319],u_xpb_out[19][319],u_xpb_out[20][319],u_xpb_out[21][319],u_xpb_out[22][319],u_xpb_out[23][319],u_xpb_out[24][319],u_xpb_out[25][319],u_xpb_out[26][319],u_xpb_out[27][319],u_xpb_out[28][319],u_xpb_out[29][319],u_xpb_out[30][319],u_xpb_out[31][319],u_xpb_out[32][319],u_xpb_out[33][319],u_xpb_out[34][319],u_xpb_out[35][319],u_xpb_out[36][319],u_xpb_out[37][319],u_xpb_out[38][319],u_xpb_out[39][319],u_xpb_out[40][319],u_xpb_out[41][319],u_xpb_out[42][319],u_xpb_out[43][319],u_xpb_out[44][319],u_xpb_out[45][319],u_xpb_out[46][319],u_xpb_out[47][319],u_xpb_out[48][319],u_xpb_out[49][319],u_xpb_out[50][319],u_xpb_out[51][319],u_xpb_out[52][319],u_xpb_out[53][319],u_xpb_out[54][319],u_xpb_out[55][319],u_xpb_out[56][319],u_xpb_out[57][319],u_xpb_out[58][319],u_xpb_out[59][319],u_xpb_out[60][319],u_xpb_out[61][319],u_xpb_out[62][319],u_xpb_out[63][319],u_xpb_out[64][319],u_xpb_out[65][319],u_xpb_out[66][319],u_xpb_out[67][319],u_xpb_out[68][319],u_xpb_out[69][319],u_xpb_out[70][319],u_xpb_out[71][319],u_xpb_out[72][319],u_xpb_out[73][319],u_xpb_out[74][319],u_xpb_out[75][319],u_xpb_out[76][319],u_xpb_out[77][319],u_xpb_out[78][319],u_xpb_out[79][319],u_xpb_out[80][319],u_xpb_out[81][319],u_xpb_out[82][319],u_xpb_out[83][319],u_xpb_out[84][319],u_xpb_out[85][319],u_xpb_out[86][319],u_xpb_out[87][319],u_xpb_out[88][319],u_xpb_out[89][319],u_xpb_out[90][319],u_xpb_out[91][319],u_xpb_out[92][319],u_xpb_out[93][319],u_xpb_out[94][319],u_xpb_out[95][319],u_xpb_out[96][319],u_xpb_out[97][319],u_xpb_out[98][319],u_xpb_out[99][319],u_xpb_out[100][319],u_xpb_out[101][319],u_xpb_out[102][319],u_xpb_out[103][319],u_xpb_out[104][319],u_xpb_out[105][319]};

assign col_out_320 = {u_xpb_out[0][320],u_xpb_out[1][320],u_xpb_out[2][320],u_xpb_out[3][320],u_xpb_out[4][320],u_xpb_out[5][320],u_xpb_out[6][320],u_xpb_out[7][320],u_xpb_out[8][320],u_xpb_out[9][320],u_xpb_out[10][320],u_xpb_out[11][320],u_xpb_out[12][320],u_xpb_out[13][320],u_xpb_out[14][320],u_xpb_out[15][320],u_xpb_out[16][320],u_xpb_out[17][320],u_xpb_out[18][320],u_xpb_out[19][320],u_xpb_out[20][320],u_xpb_out[21][320],u_xpb_out[22][320],u_xpb_out[23][320],u_xpb_out[24][320],u_xpb_out[25][320],u_xpb_out[26][320],u_xpb_out[27][320],u_xpb_out[28][320],u_xpb_out[29][320],u_xpb_out[30][320],u_xpb_out[31][320],u_xpb_out[32][320],u_xpb_out[33][320],u_xpb_out[34][320],u_xpb_out[35][320],u_xpb_out[36][320],u_xpb_out[37][320],u_xpb_out[38][320],u_xpb_out[39][320],u_xpb_out[40][320],u_xpb_out[41][320],u_xpb_out[42][320],u_xpb_out[43][320],u_xpb_out[44][320],u_xpb_out[45][320],u_xpb_out[46][320],u_xpb_out[47][320],u_xpb_out[48][320],u_xpb_out[49][320],u_xpb_out[50][320],u_xpb_out[51][320],u_xpb_out[52][320],u_xpb_out[53][320],u_xpb_out[54][320],u_xpb_out[55][320],u_xpb_out[56][320],u_xpb_out[57][320],u_xpb_out[58][320],u_xpb_out[59][320],u_xpb_out[60][320],u_xpb_out[61][320],u_xpb_out[62][320],u_xpb_out[63][320],u_xpb_out[64][320],u_xpb_out[65][320],u_xpb_out[66][320],u_xpb_out[67][320],u_xpb_out[68][320],u_xpb_out[69][320],u_xpb_out[70][320],u_xpb_out[71][320],u_xpb_out[72][320],u_xpb_out[73][320],u_xpb_out[74][320],u_xpb_out[75][320],u_xpb_out[76][320],u_xpb_out[77][320],u_xpb_out[78][320],u_xpb_out[79][320],u_xpb_out[80][320],u_xpb_out[81][320],u_xpb_out[82][320],u_xpb_out[83][320],u_xpb_out[84][320],u_xpb_out[85][320],u_xpb_out[86][320],u_xpb_out[87][320],u_xpb_out[88][320],u_xpb_out[89][320],u_xpb_out[90][320],u_xpb_out[91][320],u_xpb_out[92][320],u_xpb_out[93][320],u_xpb_out[94][320],u_xpb_out[95][320],u_xpb_out[96][320],u_xpb_out[97][320],u_xpb_out[98][320],u_xpb_out[99][320],u_xpb_out[100][320],u_xpb_out[101][320],u_xpb_out[102][320],u_xpb_out[103][320],u_xpb_out[104][320],u_xpb_out[105][320]};

assign col_out_321 = {u_xpb_out[0][321],u_xpb_out[1][321],u_xpb_out[2][321],u_xpb_out[3][321],u_xpb_out[4][321],u_xpb_out[5][321],u_xpb_out[6][321],u_xpb_out[7][321],u_xpb_out[8][321],u_xpb_out[9][321],u_xpb_out[10][321],u_xpb_out[11][321],u_xpb_out[12][321],u_xpb_out[13][321],u_xpb_out[14][321],u_xpb_out[15][321],u_xpb_out[16][321],u_xpb_out[17][321],u_xpb_out[18][321],u_xpb_out[19][321],u_xpb_out[20][321],u_xpb_out[21][321],u_xpb_out[22][321],u_xpb_out[23][321],u_xpb_out[24][321],u_xpb_out[25][321],u_xpb_out[26][321],u_xpb_out[27][321],u_xpb_out[28][321],u_xpb_out[29][321],u_xpb_out[30][321],u_xpb_out[31][321],u_xpb_out[32][321],u_xpb_out[33][321],u_xpb_out[34][321],u_xpb_out[35][321],u_xpb_out[36][321],u_xpb_out[37][321],u_xpb_out[38][321],u_xpb_out[39][321],u_xpb_out[40][321],u_xpb_out[41][321],u_xpb_out[42][321],u_xpb_out[43][321],u_xpb_out[44][321],u_xpb_out[45][321],u_xpb_out[46][321],u_xpb_out[47][321],u_xpb_out[48][321],u_xpb_out[49][321],u_xpb_out[50][321],u_xpb_out[51][321],u_xpb_out[52][321],u_xpb_out[53][321],u_xpb_out[54][321],u_xpb_out[55][321],u_xpb_out[56][321],u_xpb_out[57][321],u_xpb_out[58][321],u_xpb_out[59][321],u_xpb_out[60][321],u_xpb_out[61][321],u_xpb_out[62][321],u_xpb_out[63][321],u_xpb_out[64][321],u_xpb_out[65][321],u_xpb_out[66][321],u_xpb_out[67][321],u_xpb_out[68][321],u_xpb_out[69][321],u_xpb_out[70][321],u_xpb_out[71][321],u_xpb_out[72][321],u_xpb_out[73][321],u_xpb_out[74][321],u_xpb_out[75][321],u_xpb_out[76][321],u_xpb_out[77][321],u_xpb_out[78][321],u_xpb_out[79][321],u_xpb_out[80][321],u_xpb_out[81][321],u_xpb_out[82][321],u_xpb_out[83][321],u_xpb_out[84][321],u_xpb_out[85][321],u_xpb_out[86][321],u_xpb_out[87][321],u_xpb_out[88][321],u_xpb_out[89][321],u_xpb_out[90][321],u_xpb_out[91][321],u_xpb_out[92][321],u_xpb_out[93][321],u_xpb_out[94][321],u_xpb_out[95][321],u_xpb_out[96][321],u_xpb_out[97][321],u_xpb_out[98][321],u_xpb_out[99][321],u_xpb_out[100][321],u_xpb_out[101][321],u_xpb_out[102][321],u_xpb_out[103][321],u_xpb_out[104][321],u_xpb_out[105][321]};

assign col_out_322 = {u_xpb_out[0][322],u_xpb_out[1][322],u_xpb_out[2][322],u_xpb_out[3][322],u_xpb_out[4][322],u_xpb_out[5][322],u_xpb_out[6][322],u_xpb_out[7][322],u_xpb_out[8][322],u_xpb_out[9][322],u_xpb_out[10][322],u_xpb_out[11][322],u_xpb_out[12][322],u_xpb_out[13][322],u_xpb_out[14][322],u_xpb_out[15][322],u_xpb_out[16][322],u_xpb_out[17][322],u_xpb_out[18][322],u_xpb_out[19][322],u_xpb_out[20][322],u_xpb_out[21][322],u_xpb_out[22][322],u_xpb_out[23][322],u_xpb_out[24][322],u_xpb_out[25][322],u_xpb_out[26][322],u_xpb_out[27][322],u_xpb_out[28][322],u_xpb_out[29][322],u_xpb_out[30][322],u_xpb_out[31][322],u_xpb_out[32][322],u_xpb_out[33][322],u_xpb_out[34][322],u_xpb_out[35][322],u_xpb_out[36][322],u_xpb_out[37][322],u_xpb_out[38][322],u_xpb_out[39][322],u_xpb_out[40][322],u_xpb_out[41][322],u_xpb_out[42][322],u_xpb_out[43][322],u_xpb_out[44][322],u_xpb_out[45][322],u_xpb_out[46][322],u_xpb_out[47][322],u_xpb_out[48][322],u_xpb_out[49][322],u_xpb_out[50][322],u_xpb_out[51][322],u_xpb_out[52][322],u_xpb_out[53][322],u_xpb_out[54][322],u_xpb_out[55][322],u_xpb_out[56][322],u_xpb_out[57][322],u_xpb_out[58][322],u_xpb_out[59][322],u_xpb_out[60][322],u_xpb_out[61][322],u_xpb_out[62][322],u_xpb_out[63][322],u_xpb_out[64][322],u_xpb_out[65][322],u_xpb_out[66][322],u_xpb_out[67][322],u_xpb_out[68][322],u_xpb_out[69][322],u_xpb_out[70][322],u_xpb_out[71][322],u_xpb_out[72][322],u_xpb_out[73][322],u_xpb_out[74][322],u_xpb_out[75][322],u_xpb_out[76][322],u_xpb_out[77][322],u_xpb_out[78][322],u_xpb_out[79][322],u_xpb_out[80][322],u_xpb_out[81][322],u_xpb_out[82][322],u_xpb_out[83][322],u_xpb_out[84][322],u_xpb_out[85][322],u_xpb_out[86][322],u_xpb_out[87][322],u_xpb_out[88][322],u_xpb_out[89][322],u_xpb_out[90][322],u_xpb_out[91][322],u_xpb_out[92][322],u_xpb_out[93][322],u_xpb_out[94][322],u_xpb_out[95][322],u_xpb_out[96][322],u_xpb_out[97][322],u_xpb_out[98][322],u_xpb_out[99][322],u_xpb_out[100][322],u_xpb_out[101][322],u_xpb_out[102][322],u_xpb_out[103][322],u_xpb_out[104][322],u_xpb_out[105][322]};

assign col_out_323 = {u_xpb_out[0][323],u_xpb_out[1][323],u_xpb_out[2][323],u_xpb_out[3][323],u_xpb_out[4][323],u_xpb_out[5][323],u_xpb_out[6][323],u_xpb_out[7][323],u_xpb_out[8][323],u_xpb_out[9][323],u_xpb_out[10][323],u_xpb_out[11][323],u_xpb_out[12][323],u_xpb_out[13][323],u_xpb_out[14][323],u_xpb_out[15][323],u_xpb_out[16][323],u_xpb_out[17][323],u_xpb_out[18][323],u_xpb_out[19][323],u_xpb_out[20][323],u_xpb_out[21][323],u_xpb_out[22][323],u_xpb_out[23][323],u_xpb_out[24][323],u_xpb_out[25][323],u_xpb_out[26][323],u_xpb_out[27][323],u_xpb_out[28][323],u_xpb_out[29][323],u_xpb_out[30][323],u_xpb_out[31][323],u_xpb_out[32][323],u_xpb_out[33][323],u_xpb_out[34][323],u_xpb_out[35][323],u_xpb_out[36][323],u_xpb_out[37][323],u_xpb_out[38][323],u_xpb_out[39][323],u_xpb_out[40][323],u_xpb_out[41][323],u_xpb_out[42][323],u_xpb_out[43][323],u_xpb_out[44][323],u_xpb_out[45][323],u_xpb_out[46][323],u_xpb_out[47][323],u_xpb_out[48][323],u_xpb_out[49][323],u_xpb_out[50][323],u_xpb_out[51][323],u_xpb_out[52][323],u_xpb_out[53][323],u_xpb_out[54][323],u_xpb_out[55][323],u_xpb_out[56][323],u_xpb_out[57][323],u_xpb_out[58][323],u_xpb_out[59][323],u_xpb_out[60][323],u_xpb_out[61][323],u_xpb_out[62][323],u_xpb_out[63][323],u_xpb_out[64][323],u_xpb_out[65][323],u_xpb_out[66][323],u_xpb_out[67][323],u_xpb_out[68][323],u_xpb_out[69][323],u_xpb_out[70][323],u_xpb_out[71][323],u_xpb_out[72][323],u_xpb_out[73][323],u_xpb_out[74][323],u_xpb_out[75][323],u_xpb_out[76][323],u_xpb_out[77][323],u_xpb_out[78][323],u_xpb_out[79][323],u_xpb_out[80][323],u_xpb_out[81][323],u_xpb_out[82][323],u_xpb_out[83][323],u_xpb_out[84][323],u_xpb_out[85][323],u_xpb_out[86][323],u_xpb_out[87][323],u_xpb_out[88][323],u_xpb_out[89][323],u_xpb_out[90][323],u_xpb_out[91][323],u_xpb_out[92][323],u_xpb_out[93][323],u_xpb_out[94][323],u_xpb_out[95][323],u_xpb_out[96][323],u_xpb_out[97][323],u_xpb_out[98][323],u_xpb_out[99][323],u_xpb_out[100][323],u_xpb_out[101][323],u_xpb_out[102][323],u_xpb_out[103][323],u_xpb_out[104][323],u_xpb_out[105][323]};

assign col_out_324 = {u_xpb_out[0][324],u_xpb_out[1][324],u_xpb_out[2][324],u_xpb_out[3][324],u_xpb_out[4][324],u_xpb_out[5][324],u_xpb_out[6][324],u_xpb_out[7][324],u_xpb_out[8][324],u_xpb_out[9][324],u_xpb_out[10][324],u_xpb_out[11][324],u_xpb_out[12][324],u_xpb_out[13][324],u_xpb_out[14][324],u_xpb_out[15][324],u_xpb_out[16][324],u_xpb_out[17][324],u_xpb_out[18][324],u_xpb_out[19][324],u_xpb_out[20][324],u_xpb_out[21][324],u_xpb_out[22][324],u_xpb_out[23][324],u_xpb_out[24][324],u_xpb_out[25][324],u_xpb_out[26][324],u_xpb_out[27][324],u_xpb_out[28][324],u_xpb_out[29][324],u_xpb_out[30][324],u_xpb_out[31][324],u_xpb_out[32][324],u_xpb_out[33][324],u_xpb_out[34][324],u_xpb_out[35][324],u_xpb_out[36][324],u_xpb_out[37][324],u_xpb_out[38][324],u_xpb_out[39][324],u_xpb_out[40][324],u_xpb_out[41][324],u_xpb_out[42][324],u_xpb_out[43][324],u_xpb_out[44][324],u_xpb_out[45][324],u_xpb_out[46][324],u_xpb_out[47][324],u_xpb_out[48][324],u_xpb_out[49][324],u_xpb_out[50][324],u_xpb_out[51][324],u_xpb_out[52][324],u_xpb_out[53][324],u_xpb_out[54][324],u_xpb_out[55][324],u_xpb_out[56][324],u_xpb_out[57][324],u_xpb_out[58][324],u_xpb_out[59][324],u_xpb_out[60][324],u_xpb_out[61][324],u_xpb_out[62][324],u_xpb_out[63][324],u_xpb_out[64][324],u_xpb_out[65][324],u_xpb_out[66][324],u_xpb_out[67][324],u_xpb_out[68][324],u_xpb_out[69][324],u_xpb_out[70][324],u_xpb_out[71][324],u_xpb_out[72][324],u_xpb_out[73][324],u_xpb_out[74][324],u_xpb_out[75][324],u_xpb_out[76][324],u_xpb_out[77][324],u_xpb_out[78][324],u_xpb_out[79][324],u_xpb_out[80][324],u_xpb_out[81][324],u_xpb_out[82][324],u_xpb_out[83][324],u_xpb_out[84][324],u_xpb_out[85][324],u_xpb_out[86][324],u_xpb_out[87][324],u_xpb_out[88][324],u_xpb_out[89][324],u_xpb_out[90][324],u_xpb_out[91][324],u_xpb_out[92][324],u_xpb_out[93][324],u_xpb_out[94][324],u_xpb_out[95][324],u_xpb_out[96][324],u_xpb_out[97][324],u_xpb_out[98][324],u_xpb_out[99][324],u_xpb_out[100][324],u_xpb_out[101][324],u_xpb_out[102][324],u_xpb_out[103][324],u_xpb_out[104][324],u_xpb_out[105][324]};

assign col_out_325 = {u_xpb_out[0][325],u_xpb_out[1][325],u_xpb_out[2][325],u_xpb_out[3][325],u_xpb_out[4][325],u_xpb_out[5][325],u_xpb_out[6][325],u_xpb_out[7][325],u_xpb_out[8][325],u_xpb_out[9][325],u_xpb_out[10][325],u_xpb_out[11][325],u_xpb_out[12][325],u_xpb_out[13][325],u_xpb_out[14][325],u_xpb_out[15][325],u_xpb_out[16][325],u_xpb_out[17][325],u_xpb_out[18][325],u_xpb_out[19][325],u_xpb_out[20][325],u_xpb_out[21][325],u_xpb_out[22][325],u_xpb_out[23][325],u_xpb_out[24][325],u_xpb_out[25][325],u_xpb_out[26][325],u_xpb_out[27][325],u_xpb_out[28][325],u_xpb_out[29][325],u_xpb_out[30][325],u_xpb_out[31][325],u_xpb_out[32][325],u_xpb_out[33][325],u_xpb_out[34][325],u_xpb_out[35][325],u_xpb_out[36][325],u_xpb_out[37][325],u_xpb_out[38][325],u_xpb_out[39][325],u_xpb_out[40][325],u_xpb_out[41][325],u_xpb_out[42][325],u_xpb_out[43][325],u_xpb_out[44][325],u_xpb_out[45][325],u_xpb_out[46][325],u_xpb_out[47][325],u_xpb_out[48][325],u_xpb_out[49][325],u_xpb_out[50][325],u_xpb_out[51][325],u_xpb_out[52][325],u_xpb_out[53][325],u_xpb_out[54][325],u_xpb_out[55][325],u_xpb_out[56][325],u_xpb_out[57][325],u_xpb_out[58][325],u_xpb_out[59][325],u_xpb_out[60][325],u_xpb_out[61][325],u_xpb_out[62][325],u_xpb_out[63][325],u_xpb_out[64][325],u_xpb_out[65][325],u_xpb_out[66][325],u_xpb_out[67][325],u_xpb_out[68][325],u_xpb_out[69][325],u_xpb_out[70][325],u_xpb_out[71][325],u_xpb_out[72][325],u_xpb_out[73][325],u_xpb_out[74][325],u_xpb_out[75][325],u_xpb_out[76][325],u_xpb_out[77][325],u_xpb_out[78][325],u_xpb_out[79][325],u_xpb_out[80][325],u_xpb_out[81][325],u_xpb_out[82][325],u_xpb_out[83][325],u_xpb_out[84][325],u_xpb_out[85][325],u_xpb_out[86][325],u_xpb_out[87][325],u_xpb_out[88][325],u_xpb_out[89][325],u_xpb_out[90][325],u_xpb_out[91][325],u_xpb_out[92][325],u_xpb_out[93][325],u_xpb_out[94][325],u_xpb_out[95][325],u_xpb_out[96][325],u_xpb_out[97][325],u_xpb_out[98][325],u_xpb_out[99][325],u_xpb_out[100][325],u_xpb_out[101][325],u_xpb_out[102][325],u_xpb_out[103][325],u_xpb_out[104][325],u_xpb_out[105][325]};

assign col_out_326 = {u_xpb_out[0][326],u_xpb_out[1][326],u_xpb_out[2][326],u_xpb_out[3][326],u_xpb_out[4][326],u_xpb_out[5][326],u_xpb_out[6][326],u_xpb_out[7][326],u_xpb_out[8][326],u_xpb_out[9][326],u_xpb_out[10][326],u_xpb_out[11][326],u_xpb_out[12][326],u_xpb_out[13][326],u_xpb_out[14][326],u_xpb_out[15][326],u_xpb_out[16][326],u_xpb_out[17][326],u_xpb_out[18][326],u_xpb_out[19][326],u_xpb_out[20][326],u_xpb_out[21][326],u_xpb_out[22][326],u_xpb_out[23][326],u_xpb_out[24][326],u_xpb_out[25][326],u_xpb_out[26][326],u_xpb_out[27][326],u_xpb_out[28][326],u_xpb_out[29][326],u_xpb_out[30][326],u_xpb_out[31][326],u_xpb_out[32][326],u_xpb_out[33][326],u_xpb_out[34][326],u_xpb_out[35][326],u_xpb_out[36][326],u_xpb_out[37][326],u_xpb_out[38][326],u_xpb_out[39][326],u_xpb_out[40][326],u_xpb_out[41][326],u_xpb_out[42][326],u_xpb_out[43][326],u_xpb_out[44][326],u_xpb_out[45][326],u_xpb_out[46][326],u_xpb_out[47][326],u_xpb_out[48][326],u_xpb_out[49][326],u_xpb_out[50][326],u_xpb_out[51][326],u_xpb_out[52][326],u_xpb_out[53][326],u_xpb_out[54][326],u_xpb_out[55][326],u_xpb_out[56][326],u_xpb_out[57][326],u_xpb_out[58][326],u_xpb_out[59][326],u_xpb_out[60][326],u_xpb_out[61][326],u_xpb_out[62][326],u_xpb_out[63][326],u_xpb_out[64][326],u_xpb_out[65][326],u_xpb_out[66][326],u_xpb_out[67][326],u_xpb_out[68][326],u_xpb_out[69][326],u_xpb_out[70][326],u_xpb_out[71][326],u_xpb_out[72][326],u_xpb_out[73][326],u_xpb_out[74][326],u_xpb_out[75][326],u_xpb_out[76][326],u_xpb_out[77][326],u_xpb_out[78][326],u_xpb_out[79][326],u_xpb_out[80][326],u_xpb_out[81][326],u_xpb_out[82][326],u_xpb_out[83][326],u_xpb_out[84][326],u_xpb_out[85][326],u_xpb_out[86][326],u_xpb_out[87][326],u_xpb_out[88][326],u_xpb_out[89][326],u_xpb_out[90][326],u_xpb_out[91][326],u_xpb_out[92][326],u_xpb_out[93][326],u_xpb_out[94][326],u_xpb_out[95][326],u_xpb_out[96][326],u_xpb_out[97][326],u_xpb_out[98][326],u_xpb_out[99][326],u_xpb_out[100][326],u_xpb_out[101][326],u_xpb_out[102][326],u_xpb_out[103][326],u_xpb_out[104][326],u_xpb_out[105][326]};

assign col_out_327 = {u_xpb_out[0][327],u_xpb_out[1][327],u_xpb_out[2][327],u_xpb_out[3][327],u_xpb_out[4][327],u_xpb_out[5][327],u_xpb_out[6][327],u_xpb_out[7][327],u_xpb_out[8][327],u_xpb_out[9][327],u_xpb_out[10][327],u_xpb_out[11][327],u_xpb_out[12][327],u_xpb_out[13][327],u_xpb_out[14][327],u_xpb_out[15][327],u_xpb_out[16][327],u_xpb_out[17][327],u_xpb_out[18][327],u_xpb_out[19][327],u_xpb_out[20][327],u_xpb_out[21][327],u_xpb_out[22][327],u_xpb_out[23][327],u_xpb_out[24][327],u_xpb_out[25][327],u_xpb_out[26][327],u_xpb_out[27][327],u_xpb_out[28][327],u_xpb_out[29][327],u_xpb_out[30][327],u_xpb_out[31][327],u_xpb_out[32][327],u_xpb_out[33][327],u_xpb_out[34][327],u_xpb_out[35][327],u_xpb_out[36][327],u_xpb_out[37][327],u_xpb_out[38][327],u_xpb_out[39][327],u_xpb_out[40][327],u_xpb_out[41][327],u_xpb_out[42][327],u_xpb_out[43][327],u_xpb_out[44][327],u_xpb_out[45][327],u_xpb_out[46][327],u_xpb_out[47][327],u_xpb_out[48][327],u_xpb_out[49][327],u_xpb_out[50][327],u_xpb_out[51][327],u_xpb_out[52][327],u_xpb_out[53][327],u_xpb_out[54][327],u_xpb_out[55][327],u_xpb_out[56][327],u_xpb_out[57][327],u_xpb_out[58][327],u_xpb_out[59][327],u_xpb_out[60][327],u_xpb_out[61][327],u_xpb_out[62][327],u_xpb_out[63][327],u_xpb_out[64][327],u_xpb_out[65][327],u_xpb_out[66][327],u_xpb_out[67][327],u_xpb_out[68][327],u_xpb_out[69][327],u_xpb_out[70][327],u_xpb_out[71][327],u_xpb_out[72][327],u_xpb_out[73][327],u_xpb_out[74][327],u_xpb_out[75][327],u_xpb_out[76][327],u_xpb_out[77][327],u_xpb_out[78][327],u_xpb_out[79][327],u_xpb_out[80][327],u_xpb_out[81][327],u_xpb_out[82][327],u_xpb_out[83][327],u_xpb_out[84][327],u_xpb_out[85][327],u_xpb_out[86][327],u_xpb_out[87][327],u_xpb_out[88][327],u_xpb_out[89][327],u_xpb_out[90][327],u_xpb_out[91][327],u_xpb_out[92][327],u_xpb_out[93][327],u_xpb_out[94][327],u_xpb_out[95][327],u_xpb_out[96][327],u_xpb_out[97][327],u_xpb_out[98][327],u_xpb_out[99][327],u_xpb_out[100][327],u_xpb_out[101][327],u_xpb_out[102][327],u_xpb_out[103][327],u_xpb_out[104][327],u_xpb_out[105][327]};

assign col_out_328 = {u_xpb_out[0][328],u_xpb_out[1][328],u_xpb_out[2][328],u_xpb_out[3][328],u_xpb_out[4][328],u_xpb_out[5][328],u_xpb_out[6][328],u_xpb_out[7][328],u_xpb_out[8][328],u_xpb_out[9][328],u_xpb_out[10][328],u_xpb_out[11][328],u_xpb_out[12][328],u_xpb_out[13][328],u_xpb_out[14][328],u_xpb_out[15][328],u_xpb_out[16][328],u_xpb_out[17][328],u_xpb_out[18][328],u_xpb_out[19][328],u_xpb_out[20][328],u_xpb_out[21][328],u_xpb_out[22][328],u_xpb_out[23][328],u_xpb_out[24][328],u_xpb_out[25][328],u_xpb_out[26][328],u_xpb_out[27][328],u_xpb_out[28][328],u_xpb_out[29][328],u_xpb_out[30][328],u_xpb_out[31][328],u_xpb_out[32][328],u_xpb_out[33][328],u_xpb_out[34][328],u_xpb_out[35][328],u_xpb_out[36][328],u_xpb_out[37][328],u_xpb_out[38][328],u_xpb_out[39][328],u_xpb_out[40][328],u_xpb_out[41][328],u_xpb_out[42][328],u_xpb_out[43][328],u_xpb_out[44][328],u_xpb_out[45][328],u_xpb_out[46][328],u_xpb_out[47][328],u_xpb_out[48][328],u_xpb_out[49][328],u_xpb_out[50][328],u_xpb_out[51][328],u_xpb_out[52][328],u_xpb_out[53][328],u_xpb_out[54][328],u_xpb_out[55][328],u_xpb_out[56][328],u_xpb_out[57][328],u_xpb_out[58][328],u_xpb_out[59][328],u_xpb_out[60][328],u_xpb_out[61][328],u_xpb_out[62][328],u_xpb_out[63][328],u_xpb_out[64][328],u_xpb_out[65][328],u_xpb_out[66][328],u_xpb_out[67][328],u_xpb_out[68][328],u_xpb_out[69][328],u_xpb_out[70][328],u_xpb_out[71][328],u_xpb_out[72][328],u_xpb_out[73][328],u_xpb_out[74][328],u_xpb_out[75][328],u_xpb_out[76][328],u_xpb_out[77][328],u_xpb_out[78][328],u_xpb_out[79][328],u_xpb_out[80][328],u_xpb_out[81][328],u_xpb_out[82][328],u_xpb_out[83][328],u_xpb_out[84][328],u_xpb_out[85][328],u_xpb_out[86][328],u_xpb_out[87][328],u_xpb_out[88][328],u_xpb_out[89][328],u_xpb_out[90][328],u_xpb_out[91][328],u_xpb_out[92][328],u_xpb_out[93][328],u_xpb_out[94][328],u_xpb_out[95][328],u_xpb_out[96][328],u_xpb_out[97][328],u_xpb_out[98][328],u_xpb_out[99][328],u_xpb_out[100][328],u_xpb_out[101][328],u_xpb_out[102][328],u_xpb_out[103][328],u_xpb_out[104][328],u_xpb_out[105][328]};

assign col_out_329 = {u_xpb_out[0][329],u_xpb_out[1][329],u_xpb_out[2][329],u_xpb_out[3][329],u_xpb_out[4][329],u_xpb_out[5][329],u_xpb_out[6][329],u_xpb_out[7][329],u_xpb_out[8][329],u_xpb_out[9][329],u_xpb_out[10][329],u_xpb_out[11][329],u_xpb_out[12][329],u_xpb_out[13][329],u_xpb_out[14][329],u_xpb_out[15][329],u_xpb_out[16][329],u_xpb_out[17][329],u_xpb_out[18][329],u_xpb_out[19][329],u_xpb_out[20][329],u_xpb_out[21][329],u_xpb_out[22][329],u_xpb_out[23][329],u_xpb_out[24][329],u_xpb_out[25][329],u_xpb_out[26][329],u_xpb_out[27][329],u_xpb_out[28][329],u_xpb_out[29][329],u_xpb_out[30][329],u_xpb_out[31][329],u_xpb_out[32][329],u_xpb_out[33][329],u_xpb_out[34][329],u_xpb_out[35][329],u_xpb_out[36][329],u_xpb_out[37][329],u_xpb_out[38][329],u_xpb_out[39][329],u_xpb_out[40][329],u_xpb_out[41][329],u_xpb_out[42][329],u_xpb_out[43][329],u_xpb_out[44][329],u_xpb_out[45][329],u_xpb_out[46][329],u_xpb_out[47][329],u_xpb_out[48][329],u_xpb_out[49][329],u_xpb_out[50][329],u_xpb_out[51][329],u_xpb_out[52][329],u_xpb_out[53][329],u_xpb_out[54][329],u_xpb_out[55][329],u_xpb_out[56][329],u_xpb_out[57][329],u_xpb_out[58][329],u_xpb_out[59][329],u_xpb_out[60][329],u_xpb_out[61][329],u_xpb_out[62][329],u_xpb_out[63][329],u_xpb_out[64][329],u_xpb_out[65][329],u_xpb_out[66][329],u_xpb_out[67][329],u_xpb_out[68][329],u_xpb_out[69][329],u_xpb_out[70][329],u_xpb_out[71][329],u_xpb_out[72][329],u_xpb_out[73][329],u_xpb_out[74][329],u_xpb_out[75][329],u_xpb_out[76][329],u_xpb_out[77][329],u_xpb_out[78][329],u_xpb_out[79][329],u_xpb_out[80][329],u_xpb_out[81][329],u_xpb_out[82][329],u_xpb_out[83][329],u_xpb_out[84][329],u_xpb_out[85][329],u_xpb_out[86][329],u_xpb_out[87][329],u_xpb_out[88][329],u_xpb_out[89][329],u_xpb_out[90][329],u_xpb_out[91][329],u_xpb_out[92][329],u_xpb_out[93][329],u_xpb_out[94][329],u_xpb_out[95][329],u_xpb_out[96][329],u_xpb_out[97][329],u_xpb_out[98][329],u_xpb_out[99][329],u_xpb_out[100][329],u_xpb_out[101][329],u_xpb_out[102][329],u_xpb_out[103][329],u_xpb_out[104][329],u_xpb_out[105][329]};

assign col_out_330 = {u_xpb_out[0][330],u_xpb_out[1][330],u_xpb_out[2][330],u_xpb_out[3][330],u_xpb_out[4][330],u_xpb_out[5][330],u_xpb_out[6][330],u_xpb_out[7][330],u_xpb_out[8][330],u_xpb_out[9][330],u_xpb_out[10][330],u_xpb_out[11][330],u_xpb_out[12][330],u_xpb_out[13][330],u_xpb_out[14][330],u_xpb_out[15][330],u_xpb_out[16][330],u_xpb_out[17][330],u_xpb_out[18][330],u_xpb_out[19][330],u_xpb_out[20][330],u_xpb_out[21][330],u_xpb_out[22][330],u_xpb_out[23][330],u_xpb_out[24][330],u_xpb_out[25][330],u_xpb_out[26][330],u_xpb_out[27][330],u_xpb_out[28][330],u_xpb_out[29][330],u_xpb_out[30][330],u_xpb_out[31][330],u_xpb_out[32][330],u_xpb_out[33][330],u_xpb_out[34][330],u_xpb_out[35][330],u_xpb_out[36][330],u_xpb_out[37][330],u_xpb_out[38][330],u_xpb_out[39][330],u_xpb_out[40][330],u_xpb_out[41][330],u_xpb_out[42][330],u_xpb_out[43][330],u_xpb_out[44][330],u_xpb_out[45][330],u_xpb_out[46][330],u_xpb_out[47][330],u_xpb_out[48][330],u_xpb_out[49][330],u_xpb_out[50][330],u_xpb_out[51][330],u_xpb_out[52][330],u_xpb_out[53][330],u_xpb_out[54][330],u_xpb_out[55][330],u_xpb_out[56][330],u_xpb_out[57][330],u_xpb_out[58][330],u_xpb_out[59][330],u_xpb_out[60][330],u_xpb_out[61][330],u_xpb_out[62][330],u_xpb_out[63][330],u_xpb_out[64][330],u_xpb_out[65][330],u_xpb_out[66][330],u_xpb_out[67][330],u_xpb_out[68][330],u_xpb_out[69][330],u_xpb_out[70][330],u_xpb_out[71][330],u_xpb_out[72][330],u_xpb_out[73][330],u_xpb_out[74][330],u_xpb_out[75][330],u_xpb_out[76][330],u_xpb_out[77][330],u_xpb_out[78][330],u_xpb_out[79][330],u_xpb_out[80][330],u_xpb_out[81][330],u_xpb_out[82][330],u_xpb_out[83][330],u_xpb_out[84][330],u_xpb_out[85][330],u_xpb_out[86][330],u_xpb_out[87][330],u_xpb_out[88][330],u_xpb_out[89][330],u_xpb_out[90][330],u_xpb_out[91][330],u_xpb_out[92][330],u_xpb_out[93][330],u_xpb_out[94][330],u_xpb_out[95][330],u_xpb_out[96][330],u_xpb_out[97][330],u_xpb_out[98][330],u_xpb_out[99][330],u_xpb_out[100][330],u_xpb_out[101][330],u_xpb_out[102][330],u_xpb_out[103][330],u_xpb_out[104][330],u_xpb_out[105][330]};

assign col_out_331 = {u_xpb_out[0][331],u_xpb_out[1][331],u_xpb_out[2][331],u_xpb_out[3][331],u_xpb_out[4][331],u_xpb_out[5][331],u_xpb_out[6][331],u_xpb_out[7][331],u_xpb_out[8][331],u_xpb_out[9][331],u_xpb_out[10][331],u_xpb_out[11][331],u_xpb_out[12][331],u_xpb_out[13][331],u_xpb_out[14][331],u_xpb_out[15][331],u_xpb_out[16][331],u_xpb_out[17][331],u_xpb_out[18][331],u_xpb_out[19][331],u_xpb_out[20][331],u_xpb_out[21][331],u_xpb_out[22][331],u_xpb_out[23][331],u_xpb_out[24][331],u_xpb_out[25][331],u_xpb_out[26][331],u_xpb_out[27][331],u_xpb_out[28][331],u_xpb_out[29][331],u_xpb_out[30][331],u_xpb_out[31][331],u_xpb_out[32][331],u_xpb_out[33][331],u_xpb_out[34][331],u_xpb_out[35][331],u_xpb_out[36][331],u_xpb_out[37][331],u_xpb_out[38][331],u_xpb_out[39][331],u_xpb_out[40][331],u_xpb_out[41][331],u_xpb_out[42][331],u_xpb_out[43][331],u_xpb_out[44][331],u_xpb_out[45][331],u_xpb_out[46][331],u_xpb_out[47][331],u_xpb_out[48][331],u_xpb_out[49][331],u_xpb_out[50][331],u_xpb_out[51][331],u_xpb_out[52][331],u_xpb_out[53][331],u_xpb_out[54][331],u_xpb_out[55][331],u_xpb_out[56][331],u_xpb_out[57][331],u_xpb_out[58][331],u_xpb_out[59][331],u_xpb_out[60][331],u_xpb_out[61][331],u_xpb_out[62][331],u_xpb_out[63][331],u_xpb_out[64][331],u_xpb_out[65][331],u_xpb_out[66][331],u_xpb_out[67][331],u_xpb_out[68][331],u_xpb_out[69][331],u_xpb_out[70][331],u_xpb_out[71][331],u_xpb_out[72][331],u_xpb_out[73][331],u_xpb_out[74][331],u_xpb_out[75][331],u_xpb_out[76][331],u_xpb_out[77][331],u_xpb_out[78][331],u_xpb_out[79][331],u_xpb_out[80][331],u_xpb_out[81][331],u_xpb_out[82][331],u_xpb_out[83][331],u_xpb_out[84][331],u_xpb_out[85][331],u_xpb_out[86][331],u_xpb_out[87][331],u_xpb_out[88][331],u_xpb_out[89][331],u_xpb_out[90][331],u_xpb_out[91][331],u_xpb_out[92][331],u_xpb_out[93][331],u_xpb_out[94][331],u_xpb_out[95][331],u_xpb_out[96][331],u_xpb_out[97][331],u_xpb_out[98][331],u_xpb_out[99][331],u_xpb_out[100][331],u_xpb_out[101][331],u_xpb_out[102][331],u_xpb_out[103][331],u_xpb_out[104][331],u_xpb_out[105][331]};

assign col_out_332 = {u_xpb_out[0][332],u_xpb_out[1][332],u_xpb_out[2][332],u_xpb_out[3][332],u_xpb_out[4][332],u_xpb_out[5][332],u_xpb_out[6][332],u_xpb_out[7][332],u_xpb_out[8][332],u_xpb_out[9][332],u_xpb_out[10][332],u_xpb_out[11][332],u_xpb_out[12][332],u_xpb_out[13][332],u_xpb_out[14][332],u_xpb_out[15][332],u_xpb_out[16][332],u_xpb_out[17][332],u_xpb_out[18][332],u_xpb_out[19][332],u_xpb_out[20][332],u_xpb_out[21][332],u_xpb_out[22][332],u_xpb_out[23][332],u_xpb_out[24][332],u_xpb_out[25][332],u_xpb_out[26][332],u_xpb_out[27][332],u_xpb_out[28][332],u_xpb_out[29][332],u_xpb_out[30][332],u_xpb_out[31][332],u_xpb_out[32][332],u_xpb_out[33][332],u_xpb_out[34][332],u_xpb_out[35][332],u_xpb_out[36][332],u_xpb_out[37][332],u_xpb_out[38][332],u_xpb_out[39][332],u_xpb_out[40][332],u_xpb_out[41][332],u_xpb_out[42][332],u_xpb_out[43][332],u_xpb_out[44][332],u_xpb_out[45][332],u_xpb_out[46][332],u_xpb_out[47][332],u_xpb_out[48][332],u_xpb_out[49][332],u_xpb_out[50][332],u_xpb_out[51][332],u_xpb_out[52][332],u_xpb_out[53][332],u_xpb_out[54][332],u_xpb_out[55][332],u_xpb_out[56][332],u_xpb_out[57][332],u_xpb_out[58][332],u_xpb_out[59][332],u_xpb_out[60][332],u_xpb_out[61][332],u_xpb_out[62][332],u_xpb_out[63][332],u_xpb_out[64][332],u_xpb_out[65][332],u_xpb_out[66][332],u_xpb_out[67][332],u_xpb_out[68][332],u_xpb_out[69][332],u_xpb_out[70][332],u_xpb_out[71][332],u_xpb_out[72][332],u_xpb_out[73][332],u_xpb_out[74][332],u_xpb_out[75][332],u_xpb_out[76][332],u_xpb_out[77][332],u_xpb_out[78][332],u_xpb_out[79][332],u_xpb_out[80][332],u_xpb_out[81][332],u_xpb_out[82][332],u_xpb_out[83][332],u_xpb_out[84][332],u_xpb_out[85][332],u_xpb_out[86][332],u_xpb_out[87][332],u_xpb_out[88][332],u_xpb_out[89][332],u_xpb_out[90][332],u_xpb_out[91][332],u_xpb_out[92][332],u_xpb_out[93][332],u_xpb_out[94][332],u_xpb_out[95][332],u_xpb_out[96][332],u_xpb_out[97][332],u_xpb_out[98][332],u_xpb_out[99][332],u_xpb_out[100][332],u_xpb_out[101][332],u_xpb_out[102][332],u_xpb_out[103][332],u_xpb_out[104][332],u_xpb_out[105][332]};

assign col_out_333 = {u_xpb_out[0][333],u_xpb_out[1][333],u_xpb_out[2][333],u_xpb_out[3][333],u_xpb_out[4][333],u_xpb_out[5][333],u_xpb_out[6][333],u_xpb_out[7][333],u_xpb_out[8][333],u_xpb_out[9][333],u_xpb_out[10][333],u_xpb_out[11][333],u_xpb_out[12][333],u_xpb_out[13][333],u_xpb_out[14][333],u_xpb_out[15][333],u_xpb_out[16][333],u_xpb_out[17][333],u_xpb_out[18][333],u_xpb_out[19][333],u_xpb_out[20][333],u_xpb_out[21][333],u_xpb_out[22][333],u_xpb_out[23][333],u_xpb_out[24][333],u_xpb_out[25][333],u_xpb_out[26][333],u_xpb_out[27][333],u_xpb_out[28][333],u_xpb_out[29][333],u_xpb_out[30][333],u_xpb_out[31][333],u_xpb_out[32][333],u_xpb_out[33][333],u_xpb_out[34][333],u_xpb_out[35][333],u_xpb_out[36][333],u_xpb_out[37][333],u_xpb_out[38][333],u_xpb_out[39][333],u_xpb_out[40][333],u_xpb_out[41][333],u_xpb_out[42][333],u_xpb_out[43][333],u_xpb_out[44][333],u_xpb_out[45][333],u_xpb_out[46][333],u_xpb_out[47][333],u_xpb_out[48][333],u_xpb_out[49][333],u_xpb_out[50][333],u_xpb_out[51][333],u_xpb_out[52][333],u_xpb_out[53][333],u_xpb_out[54][333],u_xpb_out[55][333],u_xpb_out[56][333],u_xpb_out[57][333],u_xpb_out[58][333],u_xpb_out[59][333],u_xpb_out[60][333],u_xpb_out[61][333],u_xpb_out[62][333],u_xpb_out[63][333],u_xpb_out[64][333],u_xpb_out[65][333],u_xpb_out[66][333],u_xpb_out[67][333],u_xpb_out[68][333],u_xpb_out[69][333],u_xpb_out[70][333],u_xpb_out[71][333],u_xpb_out[72][333],u_xpb_out[73][333],u_xpb_out[74][333],u_xpb_out[75][333],u_xpb_out[76][333],u_xpb_out[77][333],u_xpb_out[78][333],u_xpb_out[79][333],u_xpb_out[80][333],u_xpb_out[81][333],u_xpb_out[82][333],u_xpb_out[83][333],u_xpb_out[84][333],u_xpb_out[85][333],u_xpb_out[86][333],u_xpb_out[87][333],u_xpb_out[88][333],u_xpb_out[89][333],u_xpb_out[90][333],u_xpb_out[91][333],u_xpb_out[92][333],u_xpb_out[93][333],u_xpb_out[94][333],u_xpb_out[95][333],u_xpb_out[96][333],u_xpb_out[97][333],u_xpb_out[98][333],u_xpb_out[99][333],u_xpb_out[100][333],u_xpb_out[101][333],u_xpb_out[102][333],u_xpb_out[103][333],u_xpb_out[104][333],u_xpb_out[105][333]};

assign col_out_334 = {u_xpb_out[0][334],u_xpb_out[1][334],u_xpb_out[2][334],u_xpb_out[3][334],u_xpb_out[4][334],u_xpb_out[5][334],u_xpb_out[6][334],u_xpb_out[7][334],u_xpb_out[8][334],u_xpb_out[9][334],u_xpb_out[10][334],u_xpb_out[11][334],u_xpb_out[12][334],u_xpb_out[13][334],u_xpb_out[14][334],u_xpb_out[15][334],u_xpb_out[16][334],u_xpb_out[17][334],u_xpb_out[18][334],u_xpb_out[19][334],u_xpb_out[20][334],u_xpb_out[21][334],u_xpb_out[22][334],u_xpb_out[23][334],u_xpb_out[24][334],u_xpb_out[25][334],u_xpb_out[26][334],u_xpb_out[27][334],u_xpb_out[28][334],u_xpb_out[29][334],u_xpb_out[30][334],u_xpb_out[31][334],u_xpb_out[32][334],u_xpb_out[33][334],u_xpb_out[34][334],u_xpb_out[35][334],u_xpb_out[36][334],u_xpb_out[37][334],u_xpb_out[38][334],u_xpb_out[39][334],u_xpb_out[40][334],u_xpb_out[41][334],u_xpb_out[42][334],u_xpb_out[43][334],u_xpb_out[44][334],u_xpb_out[45][334],u_xpb_out[46][334],u_xpb_out[47][334],u_xpb_out[48][334],u_xpb_out[49][334],u_xpb_out[50][334],u_xpb_out[51][334],u_xpb_out[52][334],u_xpb_out[53][334],u_xpb_out[54][334],u_xpb_out[55][334],u_xpb_out[56][334],u_xpb_out[57][334],u_xpb_out[58][334],u_xpb_out[59][334],u_xpb_out[60][334],u_xpb_out[61][334],u_xpb_out[62][334],u_xpb_out[63][334],u_xpb_out[64][334],u_xpb_out[65][334],u_xpb_out[66][334],u_xpb_out[67][334],u_xpb_out[68][334],u_xpb_out[69][334],u_xpb_out[70][334],u_xpb_out[71][334],u_xpb_out[72][334],u_xpb_out[73][334],u_xpb_out[74][334],u_xpb_out[75][334],u_xpb_out[76][334],u_xpb_out[77][334],u_xpb_out[78][334],u_xpb_out[79][334],u_xpb_out[80][334],u_xpb_out[81][334],u_xpb_out[82][334],u_xpb_out[83][334],u_xpb_out[84][334],u_xpb_out[85][334],u_xpb_out[86][334],u_xpb_out[87][334],u_xpb_out[88][334],u_xpb_out[89][334],u_xpb_out[90][334],u_xpb_out[91][334],u_xpb_out[92][334],u_xpb_out[93][334],u_xpb_out[94][334],u_xpb_out[95][334],u_xpb_out[96][334],u_xpb_out[97][334],u_xpb_out[98][334],u_xpb_out[99][334],u_xpb_out[100][334],u_xpb_out[101][334],u_xpb_out[102][334],u_xpb_out[103][334],u_xpb_out[104][334],u_xpb_out[105][334]};

assign col_out_335 = {u_xpb_out[0][335],u_xpb_out[1][335],u_xpb_out[2][335],u_xpb_out[3][335],u_xpb_out[4][335],u_xpb_out[5][335],u_xpb_out[6][335],u_xpb_out[7][335],u_xpb_out[8][335],u_xpb_out[9][335],u_xpb_out[10][335],u_xpb_out[11][335],u_xpb_out[12][335],u_xpb_out[13][335],u_xpb_out[14][335],u_xpb_out[15][335],u_xpb_out[16][335],u_xpb_out[17][335],u_xpb_out[18][335],u_xpb_out[19][335],u_xpb_out[20][335],u_xpb_out[21][335],u_xpb_out[22][335],u_xpb_out[23][335],u_xpb_out[24][335],u_xpb_out[25][335],u_xpb_out[26][335],u_xpb_out[27][335],u_xpb_out[28][335],u_xpb_out[29][335],u_xpb_out[30][335],u_xpb_out[31][335],u_xpb_out[32][335],u_xpb_out[33][335],u_xpb_out[34][335],u_xpb_out[35][335],u_xpb_out[36][335],u_xpb_out[37][335],u_xpb_out[38][335],u_xpb_out[39][335],u_xpb_out[40][335],u_xpb_out[41][335],u_xpb_out[42][335],u_xpb_out[43][335],u_xpb_out[44][335],u_xpb_out[45][335],u_xpb_out[46][335],u_xpb_out[47][335],u_xpb_out[48][335],u_xpb_out[49][335],u_xpb_out[50][335],u_xpb_out[51][335],u_xpb_out[52][335],u_xpb_out[53][335],u_xpb_out[54][335],u_xpb_out[55][335],u_xpb_out[56][335],u_xpb_out[57][335],u_xpb_out[58][335],u_xpb_out[59][335],u_xpb_out[60][335],u_xpb_out[61][335],u_xpb_out[62][335],u_xpb_out[63][335],u_xpb_out[64][335],u_xpb_out[65][335],u_xpb_out[66][335],u_xpb_out[67][335],u_xpb_out[68][335],u_xpb_out[69][335],u_xpb_out[70][335],u_xpb_out[71][335],u_xpb_out[72][335],u_xpb_out[73][335],u_xpb_out[74][335],u_xpb_out[75][335],u_xpb_out[76][335],u_xpb_out[77][335],u_xpb_out[78][335],u_xpb_out[79][335],u_xpb_out[80][335],u_xpb_out[81][335],u_xpb_out[82][335],u_xpb_out[83][335],u_xpb_out[84][335],u_xpb_out[85][335],u_xpb_out[86][335],u_xpb_out[87][335],u_xpb_out[88][335],u_xpb_out[89][335],u_xpb_out[90][335],u_xpb_out[91][335],u_xpb_out[92][335],u_xpb_out[93][335],u_xpb_out[94][335],u_xpb_out[95][335],u_xpb_out[96][335],u_xpb_out[97][335],u_xpb_out[98][335],u_xpb_out[99][335],u_xpb_out[100][335],u_xpb_out[101][335],u_xpb_out[102][335],u_xpb_out[103][335],u_xpb_out[104][335],u_xpb_out[105][335]};

assign col_out_336 = {u_xpb_out[0][336],u_xpb_out[1][336],u_xpb_out[2][336],u_xpb_out[3][336],u_xpb_out[4][336],u_xpb_out[5][336],u_xpb_out[6][336],u_xpb_out[7][336],u_xpb_out[8][336],u_xpb_out[9][336],u_xpb_out[10][336],u_xpb_out[11][336],u_xpb_out[12][336],u_xpb_out[13][336],u_xpb_out[14][336],u_xpb_out[15][336],u_xpb_out[16][336],u_xpb_out[17][336],u_xpb_out[18][336],u_xpb_out[19][336],u_xpb_out[20][336],u_xpb_out[21][336],u_xpb_out[22][336],u_xpb_out[23][336],u_xpb_out[24][336],u_xpb_out[25][336],u_xpb_out[26][336],u_xpb_out[27][336],u_xpb_out[28][336],u_xpb_out[29][336],u_xpb_out[30][336],u_xpb_out[31][336],u_xpb_out[32][336],u_xpb_out[33][336],u_xpb_out[34][336],u_xpb_out[35][336],u_xpb_out[36][336],u_xpb_out[37][336],u_xpb_out[38][336],u_xpb_out[39][336],u_xpb_out[40][336],u_xpb_out[41][336],u_xpb_out[42][336],u_xpb_out[43][336],u_xpb_out[44][336],u_xpb_out[45][336],u_xpb_out[46][336],u_xpb_out[47][336],u_xpb_out[48][336],u_xpb_out[49][336],u_xpb_out[50][336],u_xpb_out[51][336],u_xpb_out[52][336],u_xpb_out[53][336],u_xpb_out[54][336],u_xpb_out[55][336],u_xpb_out[56][336],u_xpb_out[57][336],u_xpb_out[58][336],u_xpb_out[59][336],u_xpb_out[60][336],u_xpb_out[61][336],u_xpb_out[62][336],u_xpb_out[63][336],u_xpb_out[64][336],u_xpb_out[65][336],u_xpb_out[66][336],u_xpb_out[67][336],u_xpb_out[68][336],u_xpb_out[69][336],u_xpb_out[70][336],u_xpb_out[71][336],u_xpb_out[72][336],u_xpb_out[73][336],u_xpb_out[74][336],u_xpb_out[75][336],u_xpb_out[76][336],u_xpb_out[77][336],u_xpb_out[78][336],u_xpb_out[79][336],u_xpb_out[80][336],u_xpb_out[81][336],u_xpb_out[82][336],u_xpb_out[83][336],u_xpb_out[84][336],u_xpb_out[85][336],u_xpb_out[86][336],u_xpb_out[87][336],u_xpb_out[88][336],u_xpb_out[89][336],u_xpb_out[90][336],u_xpb_out[91][336],u_xpb_out[92][336],u_xpb_out[93][336],u_xpb_out[94][336],u_xpb_out[95][336],u_xpb_out[96][336],u_xpb_out[97][336],u_xpb_out[98][336],u_xpb_out[99][336],u_xpb_out[100][336],u_xpb_out[101][336],u_xpb_out[102][336],u_xpb_out[103][336],u_xpb_out[104][336],u_xpb_out[105][336]};

assign col_out_337 = {u_xpb_out[0][337],u_xpb_out[1][337],u_xpb_out[2][337],u_xpb_out[3][337],u_xpb_out[4][337],u_xpb_out[5][337],u_xpb_out[6][337],u_xpb_out[7][337],u_xpb_out[8][337],u_xpb_out[9][337],u_xpb_out[10][337],u_xpb_out[11][337],u_xpb_out[12][337],u_xpb_out[13][337],u_xpb_out[14][337],u_xpb_out[15][337],u_xpb_out[16][337],u_xpb_out[17][337],u_xpb_out[18][337],u_xpb_out[19][337],u_xpb_out[20][337],u_xpb_out[21][337],u_xpb_out[22][337],u_xpb_out[23][337],u_xpb_out[24][337],u_xpb_out[25][337],u_xpb_out[26][337],u_xpb_out[27][337],u_xpb_out[28][337],u_xpb_out[29][337],u_xpb_out[30][337],u_xpb_out[31][337],u_xpb_out[32][337],u_xpb_out[33][337],u_xpb_out[34][337],u_xpb_out[35][337],u_xpb_out[36][337],u_xpb_out[37][337],u_xpb_out[38][337],u_xpb_out[39][337],u_xpb_out[40][337],u_xpb_out[41][337],u_xpb_out[42][337],u_xpb_out[43][337],u_xpb_out[44][337],u_xpb_out[45][337],u_xpb_out[46][337],u_xpb_out[47][337],u_xpb_out[48][337],u_xpb_out[49][337],u_xpb_out[50][337],u_xpb_out[51][337],u_xpb_out[52][337],u_xpb_out[53][337],u_xpb_out[54][337],u_xpb_out[55][337],u_xpb_out[56][337],u_xpb_out[57][337],u_xpb_out[58][337],u_xpb_out[59][337],u_xpb_out[60][337],u_xpb_out[61][337],u_xpb_out[62][337],u_xpb_out[63][337],u_xpb_out[64][337],u_xpb_out[65][337],u_xpb_out[66][337],u_xpb_out[67][337],u_xpb_out[68][337],u_xpb_out[69][337],u_xpb_out[70][337],u_xpb_out[71][337],u_xpb_out[72][337],u_xpb_out[73][337],u_xpb_out[74][337],u_xpb_out[75][337],u_xpb_out[76][337],u_xpb_out[77][337],u_xpb_out[78][337],u_xpb_out[79][337],u_xpb_out[80][337],u_xpb_out[81][337],u_xpb_out[82][337],u_xpb_out[83][337],u_xpb_out[84][337],u_xpb_out[85][337],u_xpb_out[86][337],u_xpb_out[87][337],u_xpb_out[88][337],u_xpb_out[89][337],u_xpb_out[90][337],u_xpb_out[91][337],u_xpb_out[92][337],u_xpb_out[93][337],u_xpb_out[94][337],u_xpb_out[95][337],u_xpb_out[96][337],u_xpb_out[97][337],u_xpb_out[98][337],u_xpb_out[99][337],u_xpb_out[100][337],u_xpb_out[101][337],u_xpb_out[102][337],u_xpb_out[103][337],u_xpb_out[104][337],u_xpb_out[105][337]};

assign col_out_338 = {u_xpb_out[0][338],u_xpb_out[1][338],u_xpb_out[2][338],u_xpb_out[3][338],u_xpb_out[4][338],u_xpb_out[5][338],u_xpb_out[6][338],u_xpb_out[7][338],u_xpb_out[8][338],u_xpb_out[9][338],u_xpb_out[10][338],u_xpb_out[11][338],u_xpb_out[12][338],u_xpb_out[13][338],u_xpb_out[14][338],u_xpb_out[15][338],u_xpb_out[16][338],u_xpb_out[17][338],u_xpb_out[18][338],u_xpb_out[19][338],u_xpb_out[20][338],u_xpb_out[21][338],u_xpb_out[22][338],u_xpb_out[23][338],u_xpb_out[24][338],u_xpb_out[25][338],u_xpb_out[26][338],u_xpb_out[27][338],u_xpb_out[28][338],u_xpb_out[29][338],u_xpb_out[30][338],u_xpb_out[31][338],u_xpb_out[32][338],u_xpb_out[33][338],u_xpb_out[34][338],u_xpb_out[35][338],u_xpb_out[36][338],u_xpb_out[37][338],u_xpb_out[38][338],u_xpb_out[39][338],u_xpb_out[40][338],u_xpb_out[41][338],u_xpb_out[42][338],u_xpb_out[43][338],u_xpb_out[44][338],u_xpb_out[45][338],u_xpb_out[46][338],u_xpb_out[47][338],u_xpb_out[48][338],u_xpb_out[49][338],u_xpb_out[50][338],u_xpb_out[51][338],u_xpb_out[52][338],u_xpb_out[53][338],u_xpb_out[54][338],u_xpb_out[55][338],u_xpb_out[56][338],u_xpb_out[57][338],u_xpb_out[58][338],u_xpb_out[59][338],u_xpb_out[60][338],u_xpb_out[61][338],u_xpb_out[62][338],u_xpb_out[63][338],u_xpb_out[64][338],u_xpb_out[65][338],u_xpb_out[66][338],u_xpb_out[67][338],u_xpb_out[68][338],u_xpb_out[69][338],u_xpb_out[70][338],u_xpb_out[71][338],u_xpb_out[72][338],u_xpb_out[73][338],u_xpb_out[74][338],u_xpb_out[75][338],u_xpb_out[76][338],u_xpb_out[77][338],u_xpb_out[78][338],u_xpb_out[79][338],u_xpb_out[80][338],u_xpb_out[81][338],u_xpb_out[82][338],u_xpb_out[83][338],u_xpb_out[84][338],u_xpb_out[85][338],u_xpb_out[86][338],u_xpb_out[87][338],u_xpb_out[88][338],u_xpb_out[89][338],u_xpb_out[90][338],u_xpb_out[91][338],u_xpb_out[92][338],u_xpb_out[93][338],u_xpb_out[94][338],u_xpb_out[95][338],u_xpb_out[96][338],u_xpb_out[97][338],u_xpb_out[98][338],u_xpb_out[99][338],u_xpb_out[100][338],u_xpb_out[101][338],u_xpb_out[102][338],u_xpb_out[103][338],u_xpb_out[104][338],u_xpb_out[105][338]};

assign col_out_339 = {u_xpb_out[0][339],u_xpb_out[1][339],u_xpb_out[2][339],u_xpb_out[3][339],u_xpb_out[4][339],u_xpb_out[5][339],u_xpb_out[6][339],u_xpb_out[7][339],u_xpb_out[8][339],u_xpb_out[9][339],u_xpb_out[10][339],u_xpb_out[11][339],u_xpb_out[12][339],u_xpb_out[13][339],u_xpb_out[14][339],u_xpb_out[15][339],u_xpb_out[16][339],u_xpb_out[17][339],u_xpb_out[18][339],u_xpb_out[19][339],u_xpb_out[20][339],u_xpb_out[21][339],u_xpb_out[22][339],u_xpb_out[23][339],u_xpb_out[24][339],u_xpb_out[25][339],u_xpb_out[26][339],u_xpb_out[27][339],u_xpb_out[28][339],u_xpb_out[29][339],u_xpb_out[30][339],u_xpb_out[31][339],u_xpb_out[32][339],u_xpb_out[33][339],u_xpb_out[34][339],u_xpb_out[35][339],u_xpb_out[36][339],u_xpb_out[37][339],u_xpb_out[38][339],u_xpb_out[39][339],u_xpb_out[40][339],u_xpb_out[41][339],u_xpb_out[42][339],u_xpb_out[43][339],u_xpb_out[44][339],u_xpb_out[45][339],u_xpb_out[46][339],u_xpb_out[47][339],u_xpb_out[48][339],u_xpb_out[49][339],u_xpb_out[50][339],u_xpb_out[51][339],u_xpb_out[52][339],u_xpb_out[53][339],u_xpb_out[54][339],u_xpb_out[55][339],u_xpb_out[56][339],u_xpb_out[57][339],u_xpb_out[58][339],u_xpb_out[59][339],u_xpb_out[60][339],u_xpb_out[61][339],u_xpb_out[62][339],u_xpb_out[63][339],u_xpb_out[64][339],u_xpb_out[65][339],u_xpb_out[66][339],u_xpb_out[67][339],u_xpb_out[68][339],u_xpb_out[69][339],u_xpb_out[70][339],u_xpb_out[71][339],u_xpb_out[72][339],u_xpb_out[73][339],u_xpb_out[74][339],u_xpb_out[75][339],u_xpb_out[76][339],u_xpb_out[77][339],u_xpb_out[78][339],u_xpb_out[79][339],u_xpb_out[80][339],u_xpb_out[81][339],u_xpb_out[82][339],u_xpb_out[83][339],u_xpb_out[84][339],u_xpb_out[85][339],u_xpb_out[86][339],u_xpb_out[87][339],u_xpb_out[88][339],u_xpb_out[89][339],u_xpb_out[90][339],u_xpb_out[91][339],u_xpb_out[92][339],u_xpb_out[93][339],u_xpb_out[94][339],u_xpb_out[95][339],u_xpb_out[96][339],u_xpb_out[97][339],u_xpb_out[98][339],u_xpb_out[99][339],u_xpb_out[100][339],u_xpb_out[101][339],u_xpb_out[102][339],u_xpb_out[103][339],u_xpb_out[104][339],u_xpb_out[105][339]};

assign col_out_340 = {u_xpb_out[0][340],u_xpb_out[1][340],u_xpb_out[2][340],u_xpb_out[3][340],u_xpb_out[4][340],u_xpb_out[5][340],u_xpb_out[6][340],u_xpb_out[7][340],u_xpb_out[8][340],u_xpb_out[9][340],u_xpb_out[10][340],u_xpb_out[11][340],u_xpb_out[12][340],u_xpb_out[13][340],u_xpb_out[14][340],u_xpb_out[15][340],u_xpb_out[16][340],u_xpb_out[17][340],u_xpb_out[18][340],u_xpb_out[19][340],u_xpb_out[20][340],u_xpb_out[21][340],u_xpb_out[22][340],u_xpb_out[23][340],u_xpb_out[24][340],u_xpb_out[25][340],u_xpb_out[26][340],u_xpb_out[27][340],u_xpb_out[28][340],u_xpb_out[29][340],u_xpb_out[30][340],u_xpb_out[31][340],u_xpb_out[32][340],u_xpb_out[33][340],u_xpb_out[34][340],u_xpb_out[35][340],u_xpb_out[36][340],u_xpb_out[37][340],u_xpb_out[38][340],u_xpb_out[39][340],u_xpb_out[40][340],u_xpb_out[41][340],u_xpb_out[42][340],u_xpb_out[43][340],u_xpb_out[44][340],u_xpb_out[45][340],u_xpb_out[46][340],u_xpb_out[47][340],u_xpb_out[48][340],u_xpb_out[49][340],u_xpb_out[50][340],u_xpb_out[51][340],u_xpb_out[52][340],u_xpb_out[53][340],u_xpb_out[54][340],u_xpb_out[55][340],u_xpb_out[56][340],u_xpb_out[57][340],u_xpb_out[58][340],u_xpb_out[59][340],u_xpb_out[60][340],u_xpb_out[61][340],u_xpb_out[62][340],u_xpb_out[63][340],u_xpb_out[64][340],u_xpb_out[65][340],u_xpb_out[66][340],u_xpb_out[67][340],u_xpb_out[68][340],u_xpb_out[69][340],u_xpb_out[70][340],u_xpb_out[71][340],u_xpb_out[72][340],u_xpb_out[73][340],u_xpb_out[74][340],u_xpb_out[75][340],u_xpb_out[76][340],u_xpb_out[77][340],u_xpb_out[78][340],u_xpb_out[79][340],u_xpb_out[80][340],u_xpb_out[81][340],u_xpb_out[82][340],u_xpb_out[83][340],u_xpb_out[84][340],u_xpb_out[85][340],u_xpb_out[86][340],u_xpb_out[87][340],u_xpb_out[88][340],u_xpb_out[89][340],u_xpb_out[90][340],u_xpb_out[91][340],u_xpb_out[92][340],u_xpb_out[93][340],u_xpb_out[94][340],u_xpb_out[95][340],u_xpb_out[96][340],u_xpb_out[97][340],u_xpb_out[98][340],u_xpb_out[99][340],u_xpb_out[100][340],u_xpb_out[101][340],u_xpb_out[102][340],u_xpb_out[103][340],u_xpb_out[104][340],u_xpb_out[105][340]};

assign col_out_341 = {u_xpb_out[0][341],u_xpb_out[1][341],u_xpb_out[2][341],u_xpb_out[3][341],u_xpb_out[4][341],u_xpb_out[5][341],u_xpb_out[6][341],u_xpb_out[7][341],u_xpb_out[8][341],u_xpb_out[9][341],u_xpb_out[10][341],u_xpb_out[11][341],u_xpb_out[12][341],u_xpb_out[13][341],u_xpb_out[14][341],u_xpb_out[15][341],u_xpb_out[16][341],u_xpb_out[17][341],u_xpb_out[18][341],u_xpb_out[19][341],u_xpb_out[20][341],u_xpb_out[21][341],u_xpb_out[22][341],u_xpb_out[23][341],u_xpb_out[24][341],u_xpb_out[25][341],u_xpb_out[26][341],u_xpb_out[27][341],u_xpb_out[28][341],u_xpb_out[29][341],u_xpb_out[30][341],u_xpb_out[31][341],u_xpb_out[32][341],u_xpb_out[33][341],u_xpb_out[34][341],u_xpb_out[35][341],u_xpb_out[36][341],u_xpb_out[37][341],u_xpb_out[38][341],u_xpb_out[39][341],u_xpb_out[40][341],u_xpb_out[41][341],u_xpb_out[42][341],u_xpb_out[43][341],u_xpb_out[44][341],u_xpb_out[45][341],u_xpb_out[46][341],u_xpb_out[47][341],u_xpb_out[48][341],u_xpb_out[49][341],u_xpb_out[50][341],u_xpb_out[51][341],u_xpb_out[52][341],u_xpb_out[53][341],u_xpb_out[54][341],u_xpb_out[55][341],u_xpb_out[56][341],u_xpb_out[57][341],u_xpb_out[58][341],u_xpb_out[59][341],u_xpb_out[60][341],u_xpb_out[61][341],u_xpb_out[62][341],u_xpb_out[63][341],u_xpb_out[64][341],u_xpb_out[65][341],u_xpb_out[66][341],u_xpb_out[67][341],u_xpb_out[68][341],u_xpb_out[69][341],u_xpb_out[70][341],u_xpb_out[71][341],u_xpb_out[72][341],u_xpb_out[73][341],u_xpb_out[74][341],u_xpb_out[75][341],u_xpb_out[76][341],u_xpb_out[77][341],u_xpb_out[78][341],u_xpb_out[79][341],u_xpb_out[80][341],u_xpb_out[81][341],u_xpb_out[82][341],u_xpb_out[83][341],u_xpb_out[84][341],u_xpb_out[85][341],u_xpb_out[86][341],u_xpb_out[87][341],u_xpb_out[88][341],u_xpb_out[89][341],u_xpb_out[90][341],u_xpb_out[91][341],u_xpb_out[92][341],u_xpb_out[93][341],u_xpb_out[94][341],u_xpb_out[95][341],u_xpb_out[96][341],u_xpb_out[97][341],u_xpb_out[98][341],u_xpb_out[99][341],u_xpb_out[100][341],u_xpb_out[101][341],u_xpb_out[102][341],u_xpb_out[103][341],u_xpb_out[104][341],u_xpb_out[105][341]};

assign col_out_342 = {u_xpb_out[0][342],u_xpb_out[1][342],u_xpb_out[2][342],u_xpb_out[3][342],u_xpb_out[4][342],u_xpb_out[5][342],u_xpb_out[6][342],u_xpb_out[7][342],u_xpb_out[8][342],u_xpb_out[9][342],u_xpb_out[10][342],u_xpb_out[11][342],u_xpb_out[12][342],u_xpb_out[13][342],u_xpb_out[14][342],u_xpb_out[15][342],u_xpb_out[16][342],u_xpb_out[17][342],u_xpb_out[18][342],u_xpb_out[19][342],u_xpb_out[20][342],u_xpb_out[21][342],u_xpb_out[22][342],u_xpb_out[23][342],u_xpb_out[24][342],u_xpb_out[25][342],u_xpb_out[26][342],u_xpb_out[27][342],u_xpb_out[28][342],u_xpb_out[29][342],u_xpb_out[30][342],u_xpb_out[31][342],u_xpb_out[32][342],u_xpb_out[33][342],u_xpb_out[34][342],u_xpb_out[35][342],u_xpb_out[36][342],u_xpb_out[37][342],u_xpb_out[38][342],u_xpb_out[39][342],u_xpb_out[40][342],u_xpb_out[41][342],u_xpb_out[42][342],u_xpb_out[43][342],u_xpb_out[44][342],u_xpb_out[45][342],u_xpb_out[46][342],u_xpb_out[47][342],u_xpb_out[48][342],u_xpb_out[49][342],u_xpb_out[50][342],u_xpb_out[51][342],u_xpb_out[52][342],u_xpb_out[53][342],u_xpb_out[54][342],u_xpb_out[55][342],u_xpb_out[56][342],u_xpb_out[57][342],u_xpb_out[58][342],u_xpb_out[59][342],u_xpb_out[60][342],u_xpb_out[61][342],u_xpb_out[62][342],u_xpb_out[63][342],u_xpb_out[64][342],u_xpb_out[65][342],u_xpb_out[66][342],u_xpb_out[67][342],u_xpb_out[68][342],u_xpb_out[69][342],u_xpb_out[70][342],u_xpb_out[71][342],u_xpb_out[72][342],u_xpb_out[73][342],u_xpb_out[74][342],u_xpb_out[75][342],u_xpb_out[76][342],u_xpb_out[77][342],u_xpb_out[78][342],u_xpb_out[79][342],u_xpb_out[80][342],u_xpb_out[81][342],u_xpb_out[82][342],u_xpb_out[83][342],u_xpb_out[84][342],u_xpb_out[85][342],u_xpb_out[86][342],u_xpb_out[87][342],u_xpb_out[88][342],u_xpb_out[89][342],u_xpb_out[90][342],u_xpb_out[91][342],u_xpb_out[92][342],u_xpb_out[93][342],u_xpb_out[94][342],u_xpb_out[95][342],u_xpb_out[96][342],u_xpb_out[97][342],u_xpb_out[98][342],u_xpb_out[99][342],u_xpb_out[100][342],u_xpb_out[101][342],u_xpb_out[102][342],u_xpb_out[103][342],u_xpb_out[104][342],u_xpb_out[105][342]};

assign col_out_343 = {u_xpb_out[0][343],u_xpb_out[1][343],u_xpb_out[2][343],u_xpb_out[3][343],u_xpb_out[4][343],u_xpb_out[5][343],u_xpb_out[6][343],u_xpb_out[7][343],u_xpb_out[8][343],u_xpb_out[9][343],u_xpb_out[10][343],u_xpb_out[11][343],u_xpb_out[12][343],u_xpb_out[13][343],u_xpb_out[14][343],u_xpb_out[15][343],u_xpb_out[16][343],u_xpb_out[17][343],u_xpb_out[18][343],u_xpb_out[19][343],u_xpb_out[20][343],u_xpb_out[21][343],u_xpb_out[22][343],u_xpb_out[23][343],u_xpb_out[24][343],u_xpb_out[25][343],u_xpb_out[26][343],u_xpb_out[27][343],u_xpb_out[28][343],u_xpb_out[29][343],u_xpb_out[30][343],u_xpb_out[31][343],u_xpb_out[32][343],u_xpb_out[33][343],u_xpb_out[34][343],u_xpb_out[35][343],u_xpb_out[36][343],u_xpb_out[37][343],u_xpb_out[38][343],u_xpb_out[39][343],u_xpb_out[40][343],u_xpb_out[41][343],u_xpb_out[42][343],u_xpb_out[43][343],u_xpb_out[44][343],u_xpb_out[45][343],u_xpb_out[46][343],u_xpb_out[47][343],u_xpb_out[48][343],u_xpb_out[49][343],u_xpb_out[50][343],u_xpb_out[51][343],u_xpb_out[52][343],u_xpb_out[53][343],u_xpb_out[54][343],u_xpb_out[55][343],u_xpb_out[56][343],u_xpb_out[57][343],u_xpb_out[58][343],u_xpb_out[59][343],u_xpb_out[60][343],u_xpb_out[61][343],u_xpb_out[62][343],u_xpb_out[63][343],u_xpb_out[64][343],u_xpb_out[65][343],u_xpb_out[66][343],u_xpb_out[67][343],u_xpb_out[68][343],u_xpb_out[69][343],u_xpb_out[70][343],u_xpb_out[71][343],u_xpb_out[72][343],u_xpb_out[73][343],u_xpb_out[74][343],u_xpb_out[75][343],u_xpb_out[76][343],u_xpb_out[77][343],u_xpb_out[78][343],u_xpb_out[79][343],u_xpb_out[80][343],u_xpb_out[81][343],u_xpb_out[82][343],u_xpb_out[83][343],u_xpb_out[84][343],u_xpb_out[85][343],u_xpb_out[86][343],u_xpb_out[87][343],u_xpb_out[88][343],u_xpb_out[89][343],u_xpb_out[90][343],u_xpb_out[91][343],u_xpb_out[92][343],u_xpb_out[93][343],u_xpb_out[94][343],u_xpb_out[95][343],u_xpb_out[96][343],u_xpb_out[97][343],u_xpb_out[98][343],u_xpb_out[99][343],u_xpb_out[100][343],u_xpb_out[101][343],u_xpb_out[102][343],u_xpb_out[103][343],u_xpb_out[104][343],u_xpb_out[105][343]};

assign col_out_344 = {u_xpb_out[0][344],u_xpb_out[1][344],u_xpb_out[2][344],u_xpb_out[3][344],u_xpb_out[4][344],u_xpb_out[5][344],u_xpb_out[6][344],u_xpb_out[7][344],u_xpb_out[8][344],u_xpb_out[9][344],u_xpb_out[10][344],u_xpb_out[11][344],u_xpb_out[12][344],u_xpb_out[13][344],u_xpb_out[14][344],u_xpb_out[15][344],u_xpb_out[16][344],u_xpb_out[17][344],u_xpb_out[18][344],u_xpb_out[19][344],u_xpb_out[20][344],u_xpb_out[21][344],u_xpb_out[22][344],u_xpb_out[23][344],u_xpb_out[24][344],u_xpb_out[25][344],u_xpb_out[26][344],u_xpb_out[27][344],u_xpb_out[28][344],u_xpb_out[29][344],u_xpb_out[30][344],u_xpb_out[31][344],u_xpb_out[32][344],u_xpb_out[33][344],u_xpb_out[34][344],u_xpb_out[35][344],u_xpb_out[36][344],u_xpb_out[37][344],u_xpb_out[38][344],u_xpb_out[39][344],u_xpb_out[40][344],u_xpb_out[41][344],u_xpb_out[42][344],u_xpb_out[43][344],u_xpb_out[44][344],u_xpb_out[45][344],u_xpb_out[46][344],u_xpb_out[47][344],u_xpb_out[48][344],u_xpb_out[49][344],u_xpb_out[50][344],u_xpb_out[51][344],u_xpb_out[52][344],u_xpb_out[53][344],u_xpb_out[54][344],u_xpb_out[55][344],u_xpb_out[56][344],u_xpb_out[57][344],u_xpb_out[58][344],u_xpb_out[59][344],u_xpb_out[60][344],u_xpb_out[61][344],u_xpb_out[62][344],u_xpb_out[63][344],u_xpb_out[64][344],u_xpb_out[65][344],u_xpb_out[66][344],u_xpb_out[67][344],u_xpb_out[68][344],u_xpb_out[69][344],u_xpb_out[70][344],u_xpb_out[71][344],u_xpb_out[72][344],u_xpb_out[73][344],u_xpb_out[74][344],u_xpb_out[75][344],u_xpb_out[76][344],u_xpb_out[77][344],u_xpb_out[78][344],u_xpb_out[79][344],u_xpb_out[80][344],u_xpb_out[81][344],u_xpb_out[82][344],u_xpb_out[83][344],u_xpb_out[84][344],u_xpb_out[85][344],u_xpb_out[86][344],u_xpb_out[87][344],u_xpb_out[88][344],u_xpb_out[89][344],u_xpb_out[90][344],u_xpb_out[91][344],u_xpb_out[92][344],u_xpb_out[93][344],u_xpb_out[94][344],u_xpb_out[95][344],u_xpb_out[96][344],u_xpb_out[97][344],u_xpb_out[98][344],u_xpb_out[99][344],u_xpb_out[100][344],u_xpb_out[101][344],u_xpb_out[102][344],u_xpb_out[103][344],u_xpb_out[104][344],u_xpb_out[105][344]};

assign col_out_345 = {u_xpb_out[0][345],u_xpb_out[1][345],u_xpb_out[2][345],u_xpb_out[3][345],u_xpb_out[4][345],u_xpb_out[5][345],u_xpb_out[6][345],u_xpb_out[7][345],u_xpb_out[8][345],u_xpb_out[9][345],u_xpb_out[10][345],u_xpb_out[11][345],u_xpb_out[12][345],u_xpb_out[13][345],u_xpb_out[14][345],u_xpb_out[15][345],u_xpb_out[16][345],u_xpb_out[17][345],u_xpb_out[18][345],u_xpb_out[19][345],u_xpb_out[20][345],u_xpb_out[21][345],u_xpb_out[22][345],u_xpb_out[23][345],u_xpb_out[24][345],u_xpb_out[25][345],u_xpb_out[26][345],u_xpb_out[27][345],u_xpb_out[28][345],u_xpb_out[29][345],u_xpb_out[30][345],u_xpb_out[31][345],u_xpb_out[32][345],u_xpb_out[33][345],u_xpb_out[34][345],u_xpb_out[35][345],u_xpb_out[36][345],u_xpb_out[37][345],u_xpb_out[38][345],u_xpb_out[39][345],u_xpb_out[40][345],u_xpb_out[41][345],u_xpb_out[42][345],u_xpb_out[43][345],u_xpb_out[44][345],u_xpb_out[45][345],u_xpb_out[46][345],u_xpb_out[47][345],u_xpb_out[48][345],u_xpb_out[49][345],u_xpb_out[50][345],u_xpb_out[51][345],u_xpb_out[52][345],u_xpb_out[53][345],u_xpb_out[54][345],u_xpb_out[55][345],u_xpb_out[56][345],u_xpb_out[57][345],u_xpb_out[58][345],u_xpb_out[59][345],u_xpb_out[60][345],u_xpb_out[61][345],u_xpb_out[62][345],u_xpb_out[63][345],u_xpb_out[64][345],u_xpb_out[65][345],u_xpb_out[66][345],u_xpb_out[67][345],u_xpb_out[68][345],u_xpb_out[69][345],u_xpb_out[70][345],u_xpb_out[71][345],u_xpb_out[72][345],u_xpb_out[73][345],u_xpb_out[74][345],u_xpb_out[75][345],u_xpb_out[76][345],u_xpb_out[77][345],u_xpb_out[78][345],u_xpb_out[79][345],u_xpb_out[80][345],u_xpb_out[81][345],u_xpb_out[82][345],u_xpb_out[83][345],u_xpb_out[84][345],u_xpb_out[85][345],u_xpb_out[86][345],u_xpb_out[87][345],u_xpb_out[88][345],u_xpb_out[89][345],u_xpb_out[90][345],u_xpb_out[91][345],u_xpb_out[92][345],u_xpb_out[93][345],u_xpb_out[94][345],u_xpb_out[95][345],u_xpb_out[96][345],u_xpb_out[97][345],u_xpb_out[98][345],u_xpb_out[99][345],u_xpb_out[100][345],u_xpb_out[101][345],u_xpb_out[102][345],u_xpb_out[103][345],u_xpb_out[104][345],u_xpb_out[105][345]};

assign col_out_346 = {u_xpb_out[0][346],u_xpb_out[1][346],u_xpb_out[2][346],u_xpb_out[3][346],u_xpb_out[4][346],u_xpb_out[5][346],u_xpb_out[6][346],u_xpb_out[7][346],u_xpb_out[8][346],u_xpb_out[9][346],u_xpb_out[10][346],u_xpb_out[11][346],u_xpb_out[12][346],u_xpb_out[13][346],u_xpb_out[14][346],u_xpb_out[15][346],u_xpb_out[16][346],u_xpb_out[17][346],u_xpb_out[18][346],u_xpb_out[19][346],u_xpb_out[20][346],u_xpb_out[21][346],u_xpb_out[22][346],u_xpb_out[23][346],u_xpb_out[24][346],u_xpb_out[25][346],u_xpb_out[26][346],u_xpb_out[27][346],u_xpb_out[28][346],u_xpb_out[29][346],u_xpb_out[30][346],u_xpb_out[31][346],u_xpb_out[32][346],u_xpb_out[33][346],u_xpb_out[34][346],u_xpb_out[35][346],u_xpb_out[36][346],u_xpb_out[37][346],u_xpb_out[38][346],u_xpb_out[39][346],u_xpb_out[40][346],u_xpb_out[41][346],u_xpb_out[42][346],u_xpb_out[43][346],u_xpb_out[44][346],u_xpb_out[45][346],u_xpb_out[46][346],u_xpb_out[47][346],u_xpb_out[48][346],u_xpb_out[49][346],u_xpb_out[50][346],u_xpb_out[51][346],u_xpb_out[52][346],u_xpb_out[53][346],u_xpb_out[54][346],u_xpb_out[55][346],u_xpb_out[56][346],u_xpb_out[57][346],u_xpb_out[58][346],u_xpb_out[59][346],u_xpb_out[60][346],u_xpb_out[61][346],u_xpb_out[62][346],u_xpb_out[63][346],u_xpb_out[64][346],u_xpb_out[65][346],u_xpb_out[66][346],u_xpb_out[67][346],u_xpb_out[68][346],u_xpb_out[69][346],u_xpb_out[70][346],u_xpb_out[71][346],u_xpb_out[72][346],u_xpb_out[73][346],u_xpb_out[74][346],u_xpb_out[75][346],u_xpb_out[76][346],u_xpb_out[77][346],u_xpb_out[78][346],u_xpb_out[79][346],u_xpb_out[80][346],u_xpb_out[81][346],u_xpb_out[82][346],u_xpb_out[83][346],u_xpb_out[84][346],u_xpb_out[85][346],u_xpb_out[86][346],u_xpb_out[87][346],u_xpb_out[88][346],u_xpb_out[89][346],u_xpb_out[90][346],u_xpb_out[91][346],u_xpb_out[92][346],u_xpb_out[93][346],u_xpb_out[94][346],u_xpb_out[95][346],u_xpb_out[96][346],u_xpb_out[97][346],u_xpb_out[98][346],u_xpb_out[99][346],u_xpb_out[100][346],u_xpb_out[101][346],u_xpb_out[102][346],u_xpb_out[103][346],u_xpb_out[104][346],u_xpb_out[105][346]};

assign col_out_347 = {u_xpb_out[0][347],u_xpb_out[1][347],u_xpb_out[2][347],u_xpb_out[3][347],u_xpb_out[4][347],u_xpb_out[5][347],u_xpb_out[6][347],u_xpb_out[7][347],u_xpb_out[8][347],u_xpb_out[9][347],u_xpb_out[10][347],u_xpb_out[11][347],u_xpb_out[12][347],u_xpb_out[13][347],u_xpb_out[14][347],u_xpb_out[15][347],u_xpb_out[16][347],u_xpb_out[17][347],u_xpb_out[18][347],u_xpb_out[19][347],u_xpb_out[20][347],u_xpb_out[21][347],u_xpb_out[22][347],u_xpb_out[23][347],u_xpb_out[24][347],u_xpb_out[25][347],u_xpb_out[26][347],u_xpb_out[27][347],u_xpb_out[28][347],u_xpb_out[29][347],u_xpb_out[30][347],u_xpb_out[31][347],u_xpb_out[32][347],u_xpb_out[33][347],u_xpb_out[34][347],u_xpb_out[35][347],u_xpb_out[36][347],u_xpb_out[37][347],u_xpb_out[38][347],u_xpb_out[39][347],u_xpb_out[40][347],u_xpb_out[41][347],u_xpb_out[42][347],u_xpb_out[43][347],u_xpb_out[44][347],u_xpb_out[45][347],u_xpb_out[46][347],u_xpb_out[47][347],u_xpb_out[48][347],u_xpb_out[49][347],u_xpb_out[50][347],u_xpb_out[51][347],u_xpb_out[52][347],u_xpb_out[53][347],u_xpb_out[54][347],u_xpb_out[55][347],u_xpb_out[56][347],u_xpb_out[57][347],u_xpb_out[58][347],u_xpb_out[59][347],u_xpb_out[60][347],u_xpb_out[61][347],u_xpb_out[62][347],u_xpb_out[63][347],u_xpb_out[64][347],u_xpb_out[65][347],u_xpb_out[66][347],u_xpb_out[67][347],u_xpb_out[68][347],u_xpb_out[69][347],u_xpb_out[70][347],u_xpb_out[71][347],u_xpb_out[72][347],u_xpb_out[73][347],u_xpb_out[74][347],u_xpb_out[75][347],u_xpb_out[76][347],u_xpb_out[77][347],u_xpb_out[78][347],u_xpb_out[79][347],u_xpb_out[80][347],u_xpb_out[81][347],u_xpb_out[82][347],u_xpb_out[83][347],u_xpb_out[84][347],u_xpb_out[85][347],u_xpb_out[86][347],u_xpb_out[87][347],u_xpb_out[88][347],u_xpb_out[89][347],u_xpb_out[90][347],u_xpb_out[91][347],u_xpb_out[92][347],u_xpb_out[93][347],u_xpb_out[94][347],u_xpb_out[95][347],u_xpb_out[96][347],u_xpb_out[97][347],u_xpb_out[98][347],u_xpb_out[99][347],u_xpb_out[100][347],u_xpb_out[101][347],u_xpb_out[102][347],u_xpb_out[103][347],u_xpb_out[104][347],u_xpb_out[105][347]};

assign col_out_348 = {u_xpb_out[0][348],u_xpb_out[1][348],u_xpb_out[2][348],u_xpb_out[3][348],u_xpb_out[4][348],u_xpb_out[5][348],u_xpb_out[6][348],u_xpb_out[7][348],u_xpb_out[8][348],u_xpb_out[9][348],u_xpb_out[10][348],u_xpb_out[11][348],u_xpb_out[12][348],u_xpb_out[13][348],u_xpb_out[14][348],u_xpb_out[15][348],u_xpb_out[16][348],u_xpb_out[17][348],u_xpb_out[18][348],u_xpb_out[19][348],u_xpb_out[20][348],u_xpb_out[21][348],u_xpb_out[22][348],u_xpb_out[23][348],u_xpb_out[24][348],u_xpb_out[25][348],u_xpb_out[26][348],u_xpb_out[27][348],u_xpb_out[28][348],u_xpb_out[29][348],u_xpb_out[30][348],u_xpb_out[31][348],u_xpb_out[32][348],u_xpb_out[33][348],u_xpb_out[34][348],u_xpb_out[35][348],u_xpb_out[36][348],u_xpb_out[37][348],u_xpb_out[38][348],u_xpb_out[39][348],u_xpb_out[40][348],u_xpb_out[41][348],u_xpb_out[42][348],u_xpb_out[43][348],u_xpb_out[44][348],u_xpb_out[45][348],u_xpb_out[46][348],u_xpb_out[47][348],u_xpb_out[48][348],u_xpb_out[49][348],u_xpb_out[50][348],u_xpb_out[51][348],u_xpb_out[52][348],u_xpb_out[53][348],u_xpb_out[54][348],u_xpb_out[55][348],u_xpb_out[56][348],u_xpb_out[57][348],u_xpb_out[58][348],u_xpb_out[59][348],u_xpb_out[60][348],u_xpb_out[61][348],u_xpb_out[62][348],u_xpb_out[63][348],u_xpb_out[64][348],u_xpb_out[65][348],u_xpb_out[66][348],u_xpb_out[67][348],u_xpb_out[68][348],u_xpb_out[69][348],u_xpb_out[70][348],u_xpb_out[71][348],u_xpb_out[72][348],u_xpb_out[73][348],u_xpb_out[74][348],u_xpb_out[75][348],u_xpb_out[76][348],u_xpb_out[77][348],u_xpb_out[78][348],u_xpb_out[79][348],u_xpb_out[80][348],u_xpb_out[81][348],u_xpb_out[82][348],u_xpb_out[83][348],u_xpb_out[84][348],u_xpb_out[85][348],u_xpb_out[86][348],u_xpb_out[87][348],u_xpb_out[88][348],u_xpb_out[89][348],u_xpb_out[90][348],u_xpb_out[91][348],u_xpb_out[92][348],u_xpb_out[93][348],u_xpb_out[94][348],u_xpb_out[95][348],u_xpb_out[96][348],u_xpb_out[97][348],u_xpb_out[98][348],u_xpb_out[99][348],u_xpb_out[100][348],u_xpb_out[101][348],u_xpb_out[102][348],u_xpb_out[103][348],u_xpb_out[104][348],u_xpb_out[105][348]};

assign col_out_349 = {u_xpb_out[0][349],u_xpb_out[1][349],u_xpb_out[2][349],u_xpb_out[3][349],u_xpb_out[4][349],u_xpb_out[5][349],u_xpb_out[6][349],u_xpb_out[7][349],u_xpb_out[8][349],u_xpb_out[9][349],u_xpb_out[10][349],u_xpb_out[11][349],u_xpb_out[12][349],u_xpb_out[13][349],u_xpb_out[14][349],u_xpb_out[15][349],u_xpb_out[16][349],u_xpb_out[17][349],u_xpb_out[18][349],u_xpb_out[19][349],u_xpb_out[20][349],u_xpb_out[21][349],u_xpb_out[22][349],u_xpb_out[23][349],u_xpb_out[24][349],u_xpb_out[25][349],u_xpb_out[26][349],u_xpb_out[27][349],u_xpb_out[28][349],u_xpb_out[29][349],u_xpb_out[30][349],u_xpb_out[31][349],u_xpb_out[32][349],u_xpb_out[33][349],u_xpb_out[34][349],u_xpb_out[35][349],u_xpb_out[36][349],u_xpb_out[37][349],u_xpb_out[38][349],u_xpb_out[39][349],u_xpb_out[40][349],u_xpb_out[41][349],u_xpb_out[42][349],u_xpb_out[43][349],u_xpb_out[44][349],u_xpb_out[45][349],u_xpb_out[46][349],u_xpb_out[47][349],u_xpb_out[48][349],u_xpb_out[49][349],u_xpb_out[50][349],u_xpb_out[51][349],u_xpb_out[52][349],u_xpb_out[53][349],u_xpb_out[54][349],u_xpb_out[55][349],u_xpb_out[56][349],u_xpb_out[57][349],u_xpb_out[58][349],u_xpb_out[59][349],u_xpb_out[60][349],u_xpb_out[61][349],u_xpb_out[62][349],u_xpb_out[63][349],u_xpb_out[64][349],u_xpb_out[65][349],u_xpb_out[66][349],u_xpb_out[67][349],u_xpb_out[68][349],u_xpb_out[69][349],u_xpb_out[70][349],u_xpb_out[71][349],u_xpb_out[72][349],u_xpb_out[73][349],u_xpb_out[74][349],u_xpb_out[75][349],u_xpb_out[76][349],u_xpb_out[77][349],u_xpb_out[78][349],u_xpb_out[79][349],u_xpb_out[80][349],u_xpb_out[81][349],u_xpb_out[82][349],u_xpb_out[83][349],u_xpb_out[84][349],u_xpb_out[85][349],u_xpb_out[86][349],u_xpb_out[87][349],u_xpb_out[88][349],u_xpb_out[89][349],u_xpb_out[90][349],u_xpb_out[91][349],u_xpb_out[92][349],u_xpb_out[93][349],u_xpb_out[94][349],u_xpb_out[95][349],u_xpb_out[96][349],u_xpb_out[97][349],u_xpb_out[98][349],u_xpb_out[99][349],u_xpb_out[100][349],u_xpb_out[101][349],u_xpb_out[102][349],u_xpb_out[103][349],u_xpb_out[104][349],u_xpb_out[105][349]};

assign col_out_350 = {u_xpb_out[0][350],u_xpb_out[1][350],u_xpb_out[2][350],u_xpb_out[3][350],u_xpb_out[4][350],u_xpb_out[5][350],u_xpb_out[6][350],u_xpb_out[7][350],u_xpb_out[8][350],u_xpb_out[9][350],u_xpb_out[10][350],u_xpb_out[11][350],u_xpb_out[12][350],u_xpb_out[13][350],u_xpb_out[14][350],u_xpb_out[15][350],u_xpb_out[16][350],u_xpb_out[17][350],u_xpb_out[18][350],u_xpb_out[19][350],u_xpb_out[20][350],u_xpb_out[21][350],u_xpb_out[22][350],u_xpb_out[23][350],u_xpb_out[24][350],u_xpb_out[25][350],u_xpb_out[26][350],u_xpb_out[27][350],u_xpb_out[28][350],u_xpb_out[29][350],u_xpb_out[30][350],u_xpb_out[31][350],u_xpb_out[32][350],u_xpb_out[33][350],u_xpb_out[34][350],u_xpb_out[35][350],u_xpb_out[36][350],u_xpb_out[37][350],u_xpb_out[38][350],u_xpb_out[39][350],u_xpb_out[40][350],u_xpb_out[41][350],u_xpb_out[42][350],u_xpb_out[43][350],u_xpb_out[44][350],u_xpb_out[45][350],u_xpb_out[46][350],u_xpb_out[47][350],u_xpb_out[48][350],u_xpb_out[49][350],u_xpb_out[50][350],u_xpb_out[51][350],u_xpb_out[52][350],u_xpb_out[53][350],u_xpb_out[54][350],u_xpb_out[55][350],u_xpb_out[56][350],u_xpb_out[57][350],u_xpb_out[58][350],u_xpb_out[59][350],u_xpb_out[60][350],u_xpb_out[61][350],u_xpb_out[62][350],u_xpb_out[63][350],u_xpb_out[64][350],u_xpb_out[65][350],u_xpb_out[66][350],u_xpb_out[67][350],u_xpb_out[68][350],u_xpb_out[69][350],u_xpb_out[70][350],u_xpb_out[71][350],u_xpb_out[72][350],u_xpb_out[73][350],u_xpb_out[74][350],u_xpb_out[75][350],u_xpb_out[76][350],u_xpb_out[77][350],u_xpb_out[78][350],u_xpb_out[79][350],u_xpb_out[80][350],u_xpb_out[81][350],u_xpb_out[82][350],u_xpb_out[83][350],u_xpb_out[84][350],u_xpb_out[85][350],u_xpb_out[86][350],u_xpb_out[87][350],u_xpb_out[88][350],u_xpb_out[89][350],u_xpb_out[90][350],u_xpb_out[91][350],u_xpb_out[92][350],u_xpb_out[93][350],u_xpb_out[94][350],u_xpb_out[95][350],u_xpb_out[96][350],u_xpb_out[97][350],u_xpb_out[98][350],u_xpb_out[99][350],u_xpb_out[100][350],u_xpb_out[101][350],u_xpb_out[102][350],u_xpb_out[103][350],u_xpb_out[104][350],u_xpb_out[105][350]};

assign col_out_351 = {u_xpb_out[0][351],u_xpb_out[1][351],u_xpb_out[2][351],u_xpb_out[3][351],u_xpb_out[4][351],u_xpb_out[5][351],u_xpb_out[6][351],u_xpb_out[7][351],u_xpb_out[8][351],u_xpb_out[9][351],u_xpb_out[10][351],u_xpb_out[11][351],u_xpb_out[12][351],u_xpb_out[13][351],u_xpb_out[14][351],u_xpb_out[15][351],u_xpb_out[16][351],u_xpb_out[17][351],u_xpb_out[18][351],u_xpb_out[19][351],u_xpb_out[20][351],u_xpb_out[21][351],u_xpb_out[22][351],u_xpb_out[23][351],u_xpb_out[24][351],u_xpb_out[25][351],u_xpb_out[26][351],u_xpb_out[27][351],u_xpb_out[28][351],u_xpb_out[29][351],u_xpb_out[30][351],u_xpb_out[31][351],u_xpb_out[32][351],u_xpb_out[33][351],u_xpb_out[34][351],u_xpb_out[35][351],u_xpb_out[36][351],u_xpb_out[37][351],u_xpb_out[38][351],u_xpb_out[39][351],u_xpb_out[40][351],u_xpb_out[41][351],u_xpb_out[42][351],u_xpb_out[43][351],u_xpb_out[44][351],u_xpb_out[45][351],u_xpb_out[46][351],u_xpb_out[47][351],u_xpb_out[48][351],u_xpb_out[49][351],u_xpb_out[50][351],u_xpb_out[51][351],u_xpb_out[52][351],u_xpb_out[53][351],u_xpb_out[54][351],u_xpb_out[55][351],u_xpb_out[56][351],u_xpb_out[57][351],u_xpb_out[58][351],u_xpb_out[59][351],u_xpb_out[60][351],u_xpb_out[61][351],u_xpb_out[62][351],u_xpb_out[63][351],u_xpb_out[64][351],u_xpb_out[65][351],u_xpb_out[66][351],u_xpb_out[67][351],u_xpb_out[68][351],u_xpb_out[69][351],u_xpb_out[70][351],u_xpb_out[71][351],u_xpb_out[72][351],u_xpb_out[73][351],u_xpb_out[74][351],u_xpb_out[75][351],u_xpb_out[76][351],u_xpb_out[77][351],u_xpb_out[78][351],u_xpb_out[79][351],u_xpb_out[80][351],u_xpb_out[81][351],u_xpb_out[82][351],u_xpb_out[83][351],u_xpb_out[84][351],u_xpb_out[85][351],u_xpb_out[86][351],u_xpb_out[87][351],u_xpb_out[88][351],u_xpb_out[89][351],u_xpb_out[90][351],u_xpb_out[91][351],u_xpb_out[92][351],u_xpb_out[93][351],u_xpb_out[94][351],u_xpb_out[95][351],u_xpb_out[96][351],u_xpb_out[97][351],u_xpb_out[98][351],u_xpb_out[99][351],u_xpb_out[100][351],u_xpb_out[101][351],u_xpb_out[102][351],u_xpb_out[103][351],u_xpb_out[104][351],u_xpb_out[105][351]};

assign col_out_352 = {u_xpb_out[0][352],u_xpb_out[1][352],u_xpb_out[2][352],u_xpb_out[3][352],u_xpb_out[4][352],u_xpb_out[5][352],u_xpb_out[6][352],u_xpb_out[7][352],u_xpb_out[8][352],u_xpb_out[9][352],u_xpb_out[10][352],u_xpb_out[11][352],u_xpb_out[12][352],u_xpb_out[13][352],u_xpb_out[14][352],u_xpb_out[15][352],u_xpb_out[16][352],u_xpb_out[17][352],u_xpb_out[18][352],u_xpb_out[19][352],u_xpb_out[20][352],u_xpb_out[21][352],u_xpb_out[22][352],u_xpb_out[23][352],u_xpb_out[24][352],u_xpb_out[25][352],u_xpb_out[26][352],u_xpb_out[27][352],u_xpb_out[28][352],u_xpb_out[29][352],u_xpb_out[30][352],u_xpb_out[31][352],u_xpb_out[32][352],u_xpb_out[33][352],u_xpb_out[34][352],u_xpb_out[35][352],u_xpb_out[36][352],u_xpb_out[37][352],u_xpb_out[38][352],u_xpb_out[39][352],u_xpb_out[40][352],u_xpb_out[41][352],u_xpb_out[42][352],u_xpb_out[43][352],u_xpb_out[44][352],u_xpb_out[45][352],u_xpb_out[46][352],u_xpb_out[47][352],u_xpb_out[48][352],u_xpb_out[49][352],u_xpb_out[50][352],u_xpb_out[51][352],u_xpb_out[52][352],u_xpb_out[53][352],u_xpb_out[54][352],u_xpb_out[55][352],u_xpb_out[56][352],u_xpb_out[57][352],u_xpb_out[58][352],u_xpb_out[59][352],u_xpb_out[60][352],u_xpb_out[61][352],u_xpb_out[62][352],u_xpb_out[63][352],u_xpb_out[64][352],u_xpb_out[65][352],u_xpb_out[66][352],u_xpb_out[67][352],u_xpb_out[68][352],u_xpb_out[69][352],u_xpb_out[70][352],u_xpb_out[71][352],u_xpb_out[72][352],u_xpb_out[73][352],u_xpb_out[74][352],u_xpb_out[75][352],u_xpb_out[76][352],u_xpb_out[77][352],u_xpb_out[78][352],u_xpb_out[79][352],u_xpb_out[80][352],u_xpb_out[81][352],u_xpb_out[82][352],u_xpb_out[83][352],u_xpb_out[84][352],u_xpb_out[85][352],u_xpb_out[86][352],u_xpb_out[87][352],u_xpb_out[88][352],u_xpb_out[89][352],u_xpb_out[90][352],u_xpb_out[91][352],u_xpb_out[92][352],u_xpb_out[93][352],u_xpb_out[94][352],u_xpb_out[95][352],u_xpb_out[96][352],u_xpb_out[97][352],u_xpb_out[98][352],u_xpb_out[99][352],u_xpb_out[100][352],u_xpb_out[101][352],u_xpb_out[102][352],u_xpb_out[103][352],u_xpb_out[104][352],u_xpb_out[105][352]};

assign col_out_353 = {u_xpb_out[0][353],u_xpb_out[1][353],u_xpb_out[2][353],u_xpb_out[3][353],u_xpb_out[4][353],u_xpb_out[5][353],u_xpb_out[6][353],u_xpb_out[7][353],u_xpb_out[8][353],u_xpb_out[9][353],u_xpb_out[10][353],u_xpb_out[11][353],u_xpb_out[12][353],u_xpb_out[13][353],u_xpb_out[14][353],u_xpb_out[15][353],u_xpb_out[16][353],u_xpb_out[17][353],u_xpb_out[18][353],u_xpb_out[19][353],u_xpb_out[20][353],u_xpb_out[21][353],u_xpb_out[22][353],u_xpb_out[23][353],u_xpb_out[24][353],u_xpb_out[25][353],u_xpb_out[26][353],u_xpb_out[27][353],u_xpb_out[28][353],u_xpb_out[29][353],u_xpb_out[30][353],u_xpb_out[31][353],u_xpb_out[32][353],u_xpb_out[33][353],u_xpb_out[34][353],u_xpb_out[35][353],u_xpb_out[36][353],u_xpb_out[37][353],u_xpb_out[38][353],u_xpb_out[39][353],u_xpb_out[40][353],u_xpb_out[41][353],u_xpb_out[42][353],u_xpb_out[43][353],u_xpb_out[44][353],u_xpb_out[45][353],u_xpb_out[46][353],u_xpb_out[47][353],u_xpb_out[48][353],u_xpb_out[49][353],u_xpb_out[50][353],u_xpb_out[51][353],u_xpb_out[52][353],u_xpb_out[53][353],u_xpb_out[54][353],u_xpb_out[55][353],u_xpb_out[56][353],u_xpb_out[57][353],u_xpb_out[58][353],u_xpb_out[59][353],u_xpb_out[60][353],u_xpb_out[61][353],u_xpb_out[62][353],u_xpb_out[63][353],u_xpb_out[64][353],u_xpb_out[65][353],u_xpb_out[66][353],u_xpb_out[67][353],u_xpb_out[68][353],u_xpb_out[69][353],u_xpb_out[70][353],u_xpb_out[71][353],u_xpb_out[72][353],u_xpb_out[73][353],u_xpb_out[74][353],u_xpb_out[75][353],u_xpb_out[76][353],u_xpb_out[77][353],u_xpb_out[78][353],u_xpb_out[79][353],u_xpb_out[80][353],u_xpb_out[81][353],u_xpb_out[82][353],u_xpb_out[83][353],u_xpb_out[84][353],u_xpb_out[85][353],u_xpb_out[86][353],u_xpb_out[87][353],u_xpb_out[88][353],u_xpb_out[89][353],u_xpb_out[90][353],u_xpb_out[91][353],u_xpb_out[92][353],u_xpb_out[93][353],u_xpb_out[94][353],u_xpb_out[95][353],u_xpb_out[96][353],u_xpb_out[97][353],u_xpb_out[98][353],u_xpb_out[99][353],u_xpb_out[100][353],u_xpb_out[101][353],u_xpb_out[102][353],u_xpb_out[103][353],u_xpb_out[104][353],u_xpb_out[105][353]};

assign col_out_354 = {u_xpb_out[0][354],u_xpb_out[1][354],u_xpb_out[2][354],u_xpb_out[3][354],u_xpb_out[4][354],u_xpb_out[5][354],u_xpb_out[6][354],u_xpb_out[7][354],u_xpb_out[8][354],u_xpb_out[9][354],u_xpb_out[10][354],u_xpb_out[11][354],u_xpb_out[12][354],u_xpb_out[13][354],u_xpb_out[14][354],u_xpb_out[15][354],u_xpb_out[16][354],u_xpb_out[17][354],u_xpb_out[18][354],u_xpb_out[19][354],u_xpb_out[20][354],u_xpb_out[21][354],u_xpb_out[22][354],u_xpb_out[23][354],u_xpb_out[24][354],u_xpb_out[25][354],u_xpb_out[26][354],u_xpb_out[27][354],u_xpb_out[28][354],u_xpb_out[29][354],u_xpb_out[30][354],u_xpb_out[31][354],u_xpb_out[32][354],u_xpb_out[33][354],u_xpb_out[34][354],u_xpb_out[35][354],u_xpb_out[36][354],u_xpb_out[37][354],u_xpb_out[38][354],u_xpb_out[39][354],u_xpb_out[40][354],u_xpb_out[41][354],u_xpb_out[42][354],u_xpb_out[43][354],u_xpb_out[44][354],u_xpb_out[45][354],u_xpb_out[46][354],u_xpb_out[47][354],u_xpb_out[48][354],u_xpb_out[49][354],u_xpb_out[50][354],u_xpb_out[51][354],u_xpb_out[52][354],u_xpb_out[53][354],u_xpb_out[54][354],u_xpb_out[55][354],u_xpb_out[56][354],u_xpb_out[57][354],u_xpb_out[58][354],u_xpb_out[59][354],u_xpb_out[60][354],u_xpb_out[61][354],u_xpb_out[62][354],u_xpb_out[63][354],u_xpb_out[64][354],u_xpb_out[65][354],u_xpb_out[66][354],u_xpb_out[67][354],u_xpb_out[68][354],u_xpb_out[69][354],u_xpb_out[70][354],u_xpb_out[71][354],u_xpb_out[72][354],u_xpb_out[73][354],u_xpb_out[74][354],u_xpb_out[75][354],u_xpb_out[76][354],u_xpb_out[77][354],u_xpb_out[78][354],u_xpb_out[79][354],u_xpb_out[80][354],u_xpb_out[81][354],u_xpb_out[82][354],u_xpb_out[83][354],u_xpb_out[84][354],u_xpb_out[85][354],u_xpb_out[86][354],u_xpb_out[87][354],u_xpb_out[88][354],u_xpb_out[89][354],u_xpb_out[90][354],u_xpb_out[91][354],u_xpb_out[92][354],u_xpb_out[93][354],u_xpb_out[94][354],u_xpb_out[95][354],u_xpb_out[96][354],u_xpb_out[97][354],u_xpb_out[98][354],u_xpb_out[99][354],u_xpb_out[100][354],u_xpb_out[101][354],u_xpb_out[102][354],u_xpb_out[103][354],u_xpb_out[104][354],u_xpb_out[105][354]};

assign col_out_355 = {u_xpb_out[0][355],u_xpb_out[1][355],u_xpb_out[2][355],u_xpb_out[3][355],u_xpb_out[4][355],u_xpb_out[5][355],u_xpb_out[6][355],u_xpb_out[7][355],u_xpb_out[8][355],u_xpb_out[9][355],u_xpb_out[10][355],u_xpb_out[11][355],u_xpb_out[12][355],u_xpb_out[13][355],u_xpb_out[14][355],u_xpb_out[15][355],u_xpb_out[16][355],u_xpb_out[17][355],u_xpb_out[18][355],u_xpb_out[19][355],u_xpb_out[20][355],u_xpb_out[21][355],u_xpb_out[22][355],u_xpb_out[23][355],u_xpb_out[24][355],u_xpb_out[25][355],u_xpb_out[26][355],u_xpb_out[27][355],u_xpb_out[28][355],u_xpb_out[29][355],u_xpb_out[30][355],u_xpb_out[31][355],u_xpb_out[32][355],u_xpb_out[33][355],u_xpb_out[34][355],u_xpb_out[35][355],u_xpb_out[36][355],u_xpb_out[37][355],u_xpb_out[38][355],u_xpb_out[39][355],u_xpb_out[40][355],u_xpb_out[41][355],u_xpb_out[42][355],u_xpb_out[43][355],u_xpb_out[44][355],u_xpb_out[45][355],u_xpb_out[46][355],u_xpb_out[47][355],u_xpb_out[48][355],u_xpb_out[49][355],u_xpb_out[50][355],u_xpb_out[51][355],u_xpb_out[52][355],u_xpb_out[53][355],u_xpb_out[54][355],u_xpb_out[55][355],u_xpb_out[56][355],u_xpb_out[57][355],u_xpb_out[58][355],u_xpb_out[59][355],u_xpb_out[60][355],u_xpb_out[61][355],u_xpb_out[62][355],u_xpb_out[63][355],u_xpb_out[64][355],u_xpb_out[65][355],u_xpb_out[66][355],u_xpb_out[67][355],u_xpb_out[68][355],u_xpb_out[69][355],u_xpb_out[70][355],u_xpb_out[71][355],u_xpb_out[72][355],u_xpb_out[73][355],u_xpb_out[74][355],u_xpb_out[75][355],u_xpb_out[76][355],u_xpb_out[77][355],u_xpb_out[78][355],u_xpb_out[79][355],u_xpb_out[80][355],u_xpb_out[81][355],u_xpb_out[82][355],u_xpb_out[83][355],u_xpb_out[84][355],u_xpb_out[85][355],u_xpb_out[86][355],u_xpb_out[87][355],u_xpb_out[88][355],u_xpb_out[89][355],u_xpb_out[90][355],u_xpb_out[91][355],u_xpb_out[92][355],u_xpb_out[93][355],u_xpb_out[94][355],u_xpb_out[95][355],u_xpb_out[96][355],u_xpb_out[97][355],u_xpb_out[98][355],u_xpb_out[99][355],u_xpb_out[100][355],u_xpb_out[101][355],u_xpb_out[102][355],u_xpb_out[103][355],u_xpb_out[104][355],u_xpb_out[105][355]};

assign col_out_356 = {u_xpb_out[0][356],u_xpb_out[1][356],u_xpb_out[2][356],u_xpb_out[3][356],u_xpb_out[4][356],u_xpb_out[5][356],u_xpb_out[6][356],u_xpb_out[7][356],u_xpb_out[8][356],u_xpb_out[9][356],u_xpb_out[10][356],u_xpb_out[11][356],u_xpb_out[12][356],u_xpb_out[13][356],u_xpb_out[14][356],u_xpb_out[15][356],u_xpb_out[16][356],u_xpb_out[17][356],u_xpb_out[18][356],u_xpb_out[19][356],u_xpb_out[20][356],u_xpb_out[21][356],u_xpb_out[22][356],u_xpb_out[23][356],u_xpb_out[24][356],u_xpb_out[25][356],u_xpb_out[26][356],u_xpb_out[27][356],u_xpb_out[28][356],u_xpb_out[29][356],u_xpb_out[30][356],u_xpb_out[31][356],u_xpb_out[32][356],u_xpb_out[33][356],u_xpb_out[34][356],u_xpb_out[35][356],u_xpb_out[36][356],u_xpb_out[37][356],u_xpb_out[38][356],u_xpb_out[39][356],u_xpb_out[40][356],u_xpb_out[41][356],u_xpb_out[42][356],u_xpb_out[43][356],u_xpb_out[44][356],u_xpb_out[45][356],u_xpb_out[46][356],u_xpb_out[47][356],u_xpb_out[48][356],u_xpb_out[49][356],u_xpb_out[50][356],u_xpb_out[51][356],u_xpb_out[52][356],u_xpb_out[53][356],u_xpb_out[54][356],u_xpb_out[55][356],u_xpb_out[56][356],u_xpb_out[57][356],u_xpb_out[58][356],u_xpb_out[59][356],u_xpb_out[60][356],u_xpb_out[61][356],u_xpb_out[62][356],u_xpb_out[63][356],u_xpb_out[64][356],u_xpb_out[65][356],u_xpb_out[66][356],u_xpb_out[67][356],u_xpb_out[68][356],u_xpb_out[69][356],u_xpb_out[70][356],u_xpb_out[71][356],u_xpb_out[72][356],u_xpb_out[73][356],u_xpb_out[74][356],u_xpb_out[75][356],u_xpb_out[76][356],u_xpb_out[77][356],u_xpb_out[78][356],u_xpb_out[79][356],u_xpb_out[80][356],u_xpb_out[81][356],u_xpb_out[82][356],u_xpb_out[83][356],u_xpb_out[84][356],u_xpb_out[85][356],u_xpb_out[86][356],u_xpb_out[87][356],u_xpb_out[88][356],u_xpb_out[89][356],u_xpb_out[90][356],u_xpb_out[91][356],u_xpb_out[92][356],u_xpb_out[93][356],u_xpb_out[94][356],u_xpb_out[95][356],u_xpb_out[96][356],u_xpb_out[97][356],u_xpb_out[98][356],u_xpb_out[99][356],u_xpb_out[100][356],u_xpb_out[101][356],u_xpb_out[102][356],u_xpb_out[103][356],u_xpb_out[104][356],u_xpb_out[105][356]};

assign col_out_357 = {u_xpb_out[0][357],u_xpb_out[1][357],u_xpb_out[2][357],u_xpb_out[3][357],u_xpb_out[4][357],u_xpb_out[5][357],u_xpb_out[6][357],u_xpb_out[7][357],u_xpb_out[8][357],u_xpb_out[9][357],u_xpb_out[10][357],u_xpb_out[11][357],u_xpb_out[12][357],u_xpb_out[13][357],u_xpb_out[14][357],u_xpb_out[15][357],u_xpb_out[16][357],u_xpb_out[17][357],u_xpb_out[18][357],u_xpb_out[19][357],u_xpb_out[20][357],u_xpb_out[21][357],u_xpb_out[22][357],u_xpb_out[23][357],u_xpb_out[24][357],u_xpb_out[25][357],u_xpb_out[26][357],u_xpb_out[27][357],u_xpb_out[28][357],u_xpb_out[29][357],u_xpb_out[30][357],u_xpb_out[31][357],u_xpb_out[32][357],u_xpb_out[33][357],u_xpb_out[34][357],u_xpb_out[35][357],u_xpb_out[36][357],u_xpb_out[37][357],u_xpb_out[38][357],u_xpb_out[39][357],u_xpb_out[40][357],u_xpb_out[41][357],u_xpb_out[42][357],u_xpb_out[43][357],u_xpb_out[44][357],u_xpb_out[45][357],u_xpb_out[46][357],u_xpb_out[47][357],u_xpb_out[48][357],u_xpb_out[49][357],u_xpb_out[50][357],u_xpb_out[51][357],u_xpb_out[52][357],u_xpb_out[53][357],u_xpb_out[54][357],u_xpb_out[55][357],u_xpb_out[56][357],u_xpb_out[57][357],u_xpb_out[58][357],u_xpb_out[59][357],u_xpb_out[60][357],u_xpb_out[61][357],u_xpb_out[62][357],u_xpb_out[63][357],u_xpb_out[64][357],u_xpb_out[65][357],u_xpb_out[66][357],u_xpb_out[67][357],u_xpb_out[68][357],u_xpb_out[69][357],u_xpb_out[70][357],u_xpb_out[71][357],u_xpb_out[72][357],u_xpb_out[73][357],u_xpb_out[74][357],u_xpb_out[75][357],u_xpb_out[76][357],u_xpb_out[77][357],u_xpb_out[78][357],u_xpb_out[79][357],u_xpb_out[80][357],u_xpb_out[81][357],u_xpb_out[82][357],u_xpb_out[83][357],u_xpb_out[84][357],u_xpb_out[85][357],u_xpb_out[86][357],u_xpb_out[87][357],u_xpb_out[88][357],u_xpb_out[89][357],u_xpb_out[90][357],u_xpb_out[91][357],u_xpb_out[92][357],u_xpb_out[93][357],u_xpb_out[94][357],u_xpb_out[95][357],u_xpb_out[96][357],u_xpb_out[97][357],u_xpb_out[98][357],u_xpb_out[99][357],u_xpb_out[100][357],u_xpb_out[101][357],u_xpb_out[102][357],u_xpb_out[103][357],u_xpb_out[104][357],u_xpb_out[105][357]};

assign col_out_358 = {u_xpb_out[0][358],u_xpb_out[1][358],u_xpb_out[2][358],u_xpb_out[3][358],u_xpb_out[4][358],u_xpb_out[5][358],u_xpb_out[6][358],u_xpb_out[7][358],u_xpb_out[8][358],u_xpb_out[9][358],u_xpb_out[10][358],u_xpb_out[11][358],u_xpb_out[12][358],u_xpb_out[13][358],u_xpb_out[14][358],u_xpb_out[15][358],u_xpb_out[16][358],u_xpb_out[17][358],u_xpb_out[18][358],u_xpb_out[19][358],u_xpb_out[20][358],u_xpb_out[21][358],u_xpb_out[22][358],u_xpb_out[23][358],u_xpb_out[24][358],u_xpb_out[25][358],u_xpb_out[26][358],u_xpb_out[27][358],u_xpb_out[28][358],u_xpb_out[29][358],u_xpb_out[30][358],u_xpb_out[31][358],u_xpb_out[32][358],u_xpb_out[33][358],u_xpb_out[34][358],u_xpb_out[35][358],u_xpb_out[36][358],u_xpb_out[37][358],u_xpb_out[38][358],u_xpb_out[39][358],u_xpb_out[40][358],u_xpb_out[41][358],u_xpb_out[42][358],u_xpb_out[43][358],u_xpb_out[44][358],u_xpb_out[45][358],u_xpb_out[46][358],u_xpb_out[47][358],u_xpb_out[48][358],u_xpb_out[49][358],u_xpb_out[50][358],u_xpb_out[51][358],u_xpb_out[52][358],u_xpb_out[53][358],u_xpb_out[54][358],u_xpb_out[55][358],u_xpb_out[56][358],u_xpb_out[57][358],u_xpb_out[58][358],u_xpb_out[59][358],u_xpb_out[60][358],u_xpb_out[61][358],u_xpb_out[62][358],u_xpb_out[63][358],u_xpb_out[64][358],u_xpb_out[65][358],u_xpb_out[66][358],u_xpb_out[67][358],u_xpb_out[68][358],u_xpb_out[69][358],u_xpb_out[70][358],u_xpb_out[71][358],u_xpb_out[72][358],u_xpb_out[73][358],u_xpb_out[74][358],u_xpb_out[75][358],u_xpb_out[76][358],u_xpb_out[77][358],u_xpb_out[78][358],u_xpb_out[79][358],u_xpb_out[80][358],u_xpb_out[81][358],u_xpb_out[82][358],u_xpb_out[83][358],u_xpb_out[84][358],u_xpb_out[85][358],u_xpb_out[86][358],u_xpb_out[87][358],u_xpb_out[88][358],u_xpb_out[89][358],u_xpb_out[90][358],u_xpb_out[91][358],u_xpb_out[92][358],u_xpb_out[93][358],u_xpb_out[94][358],u_xpb_out[95][358],u_xpb_out[96][358],u_xpb_out[97][358],u_xpb_out[98][358],u_xpb_out[99][358],u_xpb_out[100][358],u_xpb_out[101][358],u_xpb_out[102][358],u_xpb_out[103][358],u_xpb_out[104][358],u_xpb_out[105][358]};

assign col_out_359 = {u_xpb_out[0][359],u_xpb_out[1][359],u_xpb_out[2][359],u_xpb_out[3][359],u_xpb_out[4][359],u_xpb_out[5][359],u_xpb_out[6][359],u_xpb_out[7][359],u_xpb_out[8][359],u_xpb_out[9][359],u_xpb_out[10][359],u_xpb_out[11][359],u_xpb_out[12][359],u_xpb_out[13][359],u_xpb_out[14][359],u_xpb_out[15][359],u_xpb_out[16][359],u_xpb_out[17][359],u_xpb_out[18][359],u_xpb_out[19][359],u_xpb_out[20][359],u_xpb_out[21][359],u_xpb_out[22][359],u_xpb_out[23][359],u_xpb_out[24][359],u_xpb_out[25][359],u_xpb_out[26][359],u_xpb_out[27][359],u_xpb_out[28][359],u_xpb_out[29][359],u_xpb_out[30][359],u_xpb_out[31][359],u_xpb_out[32][359],u_xpb_out[33][359],u_xpb_out[34][359],u_xpb_out[35][359],u_xpb_out[36][359],u_xpb_out[37][359],u_xpb_out[38][359],u_xpb_out[39][359],u_xpb_out[40][359],u_xpb_out[41][359],u_xpb_out[42][359],u_xpb_out[43][359],u_xpb_out[44][359],u_xpb_out[45][359],u_xpb_out[46][359],u_xpb_out[47][359],u_xpb_out[48][359],u_xpb_out[49][359],u_xpb_out[50][359],u_xpb_out[51][359],u_xpb_out[52][359],u_xpb_out[53][359],u_xpb_out[54][359],u_xpb_out[55][359],u_xpb_out[56][359],u_xpb_out[57][359],u_xpb_out[58][359],u_xpb_out[59][359],u_xpb_out[60][359],u_xpb_out[61][359],u_xpb_out[62][359],u_xpb_out[63][359],u_xpb_out[64][359],u_xpb_out[65][359],u_xpb_out[66][359],u_xpb_out[67][359],u_xpb_out[68][359],u_xpb_out[69][359],u_xpb_out[70][359],u_xpb_out[71][359],u_xpb_out[72][359],u_xpb_out[73][359],u_xpb_out[74][359],u_xpb_out[75][359],u_xpb_out[76][359],u_xpb_out[77][359],u_xpb_out[78][359],u_xpb_out[79][359],u_xpb_out[80][359],u_xpb_out[81][359],u_xpb_out[82][359],u_xpb_out[83][359],u_xpb_out[84][359],u_xpb_out[85][359],u_xpb_out[86][359],u_xpb_out[87][359],u_xpb_out[88][359],u_xpb_out[89][359],u_xpb_out[90][359],u_xpb_out[91][359],u_xpb_out[92][359],u_xpb_out[93][359],u_xpb_out[94][359],u_xpb_out[95][359],u_xpb_out[96][359],u_xpb_out[97][359],u_xpb_out[98][359],u_xpb_out[99][359],u_xpb_out[100][359],u_xpb_out[101][359],u_xpb_out[102][359],u_xpb_out[103][359],u_xpb_out[104][359],u_xpb_out[105][359]};

assign col_out_360 = {u_xpb_out[0][360],u_xpb_out[1][360],u_xpb_out[2][360],u_xpb_out[3][360],u_xpb_out[4][360],u_xpb_out[5][360],u_xpb_out[6][360],u_xpb_out[7][360],u_xpb_out[8][360],u_xpb_out[9][360],u_xpb_out[10][360],u_xpb_out[11][360],u_xpb_out[12][360],u_xpb_out[13][360],u_xpb_out[14][360],u_xpb_out[15][360],u_xpb_out[16][360],u_xpb_out[17][360],u_xpb_out[18][360],u_xpb_out[19][360],u_xpb_out[20][360],u_xpb_out[21][360],u_xpb_out[22][360],u_xpb_out[23][360],u_xpb_out[24][360],u_xpb_out[25][360],u_xpb_out[26][360],u_xpb_out[27][360],u_xpb_out[28][360],u_xpb_out[29][360],u_xpb_out[30][360],u_xpb_out[31][360],u_xpb_out[32][360],u_xpb_out[33][360],u_xpb_out[34][360],u_xpb_out[35][360],u_xpb_out[36][360],u_xpb_out[37][360],u_xpb_out[38][360],u_xpb_out[39][360],u_xpb_out[40][360],u_xpb_out[41][360],u_xpb_out[42][360],u_xpb_out[43][360],u_xpb_out[44][360],u_xpb_out[45][360],u_xpb_out[46][360],u_xpb_out[47][360],u_xpb_out[48][360],u_xpb_out[49][360],u_xpb_out[50][360],u_xpb_out[51][360],u_xpb_out[52][360],u_xpb_out[53][360],u_xpb_out[54][360],u_xpb_out[55][360],u_xpb_out[56][360],u_xpb_out[57][360],u_xpb_out[58][360],u_xpb_out[59][360],u_xpb_out[60][360],u_xpb_out[61][360],u_xpb_out[62][360],u_xpb_out[63][360],u_xpb_out[64][360],u_xpb_out[65][360],u_xpb_out[66][360],u_xpb_out[67][360],u_xpb_out[68][360],u_xpb_out[69][360],u_xpb_out[70][360],u_xpb_out[71][360],u_xpb_out[72][360],u_xpb_out[73][360],u_xpb_out[74][360],u_xpb_out[75][360],u_xpb_out[76][360],u_xpb_out[77][360],u_xpb_out[78][360],u_xpb_out[79][360],u_xpb_out[80][360],u_xpb_out[81][360],u_xpb_out[82][360],u_xpb_out[83][360],u_xpb_out[84][360],u_xpb_out[85][360],u_xpb_out[86][360],u_xpb_out[87][360],u_xpb_out[88][360],u_xpb_out[89][360],u_xpb_out[90][360],u_xpb_out[91][360],u_xpb_out[92][360],u_xpb_out[93][360],u_xpb_out[94][360],u_xpb_out[95][360],u_xpb_out[96][360],u_xpb_out[97][360],u_xpb_out[98][360],u_xpb_out[99][360],u_xpb_out[100][360],u_xpb_out[101][360],u_xpb_out[102][360],u_xpb_out[103][360],u_xpb_out[104][360],u_xpb_out[105][360]};

assign col_out_361 = {u_xpb_out[0][361],u_xpb_out[1][361],u_xpb_out[2][361],u_xpb_out[3][361],u_xpb_out[4][361],u_xpb_out[5][361],u_xpb_out[6][361],u_xpb_out[7][361],u_xpb_out[8][361],u_xpb_out[9][361],u_xpb_out[10][361],u_xpb_out[11][361],u_xpb_out[12][361],u_xpb_out[13][361],u_xpb_out[14][361],u_xpb_out[15][361],u_xpb_out[16][361],u_xpb_out[17][361],u_xpb_out[18][361],u_xpb_out[19][361],u_xpb_out[20][361],u_xpb_out[21][361],u_xpb_out[22][361],u_xpb_out[23][361],u_xpb_out[24][361],u_xpb_out[25][361],u_xpb_out[26][361],u_xpb_out[27][361],u_xpb_out[28][361],u_xpb_out[29][361],u_xpb_out[30][361],u_xpb_out[31][361],u_xpb_out[32][361],u_xpb_out[33][361],u_xpb_out[34][361],u_xpb_out[35][361],u_xpb_out[36][361],u_xpb_out[37][361],u_xpb_out[38][361],u_xpb_out[39][361],u_xpb_out[40][361],u_xpb_out[41][361],u_xpb_out[42][361],u_xpb_out[43][361],u_xpb_out[44][361],u_xpb_out[45][361],u_xpb_out[46][361],u_xpb_out[47][361],u_xpb_out[48][361],u_xpb_out[49][361],u_xpb_out[50][361],u_xpb_out[51][361],u_xpb_out[52][361],u_xpb_out[53][361],u_xpb_out[54][361],u_xpb_out[55][361],u_xpb_out[56][361],u_xpb_out[57][361],u_xpb_out[58][361],u_xpb_out[59][361],u_xpb_out[60][361],u_xpb_out[61][361],u_xpb_out[62][361],u_xpb_out[63][361],u_xpb_out[64][361],u_xpb_out[65][361],u_xpb_out[66][361],u_xpb_out[67][361],u_xpb_out[68][361],u_xpb_out[69][361],u_xpb_out[70][361],u_xpb_out[71][361],u_xpb_out[72][361],u_xpb_out[73][361],u_xpb_out[74][361],u_xpb_out[75][361],u_xpb_out[76][361],u_xpb_out[77][361],u_xpb_out[78][361],u_xpb_out[79][361],u_xpb_out[80][361],u_xpb_out[81][361],u_xpb_out[82][361],u_xpb_out[83][361],u_xpb_out[84][361],u_xpb_out[85][361],u_xpb_out[86][361],u_xpb_out[87][361],u_xpb_out[88][361],u_xpb_out[89][361],u_xpb_out[90][361],u_xpb_out[91][361],u_xpb_out[92][361],u_xpb_out[93][361],u_xpb_out[94][361],u_xpb_out[95][361],u_xpb_out[96][361],u_xpb_out[97][361],u_xpb_out[98][361],u_xpb_out[99][361],u_xpb_out[100][361],u_xpb_out[101][361],u_xpb_out[102][361],u_xpb_out[103][361],u_xpb_out[104][361],u_xpb_out[105][361]};

assign col_out_362 = {u_xpb_out[0][362],u_xpb_out[1][362],u_xpb_out[2][362],u_xpb_out[3][362],u_xpb_out[4][362],u_xpb_out[5][362],u_xpb_out[6][362],u_xpb_out[7][362],u_xpb_out[8][362],u_xpb_out[9][362],u_xpb_out[10][362],u_xpb_out[11][362],u_xpb_out[12][362],u_xpb_out[13][362],u_xpb_out[14][362],u_xpb_out[15][362],u_xpb_out[16][362],u_xpb_out[17][362],u_xpb_out[18][362],u_xpb_out[19][362],u_xpb_out[20][362],u_xpb_out[21][362],u_xpb_out[22][362],u_xpb_out[23][362],u_xpb_out[24][362],u_xpb_out[25][362],u_xpb_out[26][362],u_xpb_out[27][362],u_xpb_out[28][362],u_xpb_out[29][362],u_xpb_out[30][362],u_xpb_out[31][362],u_xpb_out[32][362],u_xpb_out[33][362],u_xpb_out[34][362],u_xpb_out[35][362],u_xpb_out[36][362],u_xpb_out[37][362],u_xpb_out[38][362],u_xpb_out[39][362],u_xpb_out[40][362],u_xpb_out[41][362],u_xpb_out[42][362],u_xpb_out[43][362],u_xpb_out[44][362],u_xpb_out[45][362],u_xpb_out[46][362],u_xpb_out[47][362],u_xpb_out[48][362],u_xpb_out[49][362],u_xpb_out[50][362],u_xpb_out[51][362],u_xpb_out[52][362],u_xpb_out[53][362],u_xpb_out[54][362],u_xpb_out[55][362],u_xpb_out[56][362],u_xpb_out[57][362],u_xpb_out[58][362],u_xpb_out[59][362],u_xpb_out[60][362],u_xpb_out[61][362],u_xpb_out[62][362],u_xpb_out[63][362],u_xpb_out[64][362],u_xpb_out[65][362],u_xpb_out[66][362],u_xpb_out[67][362],u_xpb_out[68][362],u_xpb_out[69][362],u_xpb_out[70][362],u_xpb_out[71][362],u_xpb_out[72][362],u_xpb_out[73][362],u_xpb_out[74][362],u_xpb_out[75][362],u_xpb_out[76][362],u_xpb_out[77][362],u_xpb_out[78][362],u_xpb_out[79][362],u_xpb_out[80][362],u_xpb_out[81][362],u_xpb_out[82][362],u_xpb_out[83][362],u_xpb_out[84][362],u_xpb_out[85][362],u_xpb_out[86][362],u_xpb_out[87][362],u_xpb_out[88][362],u_xpb_out[89][362],u_xpb_out[90][362],u_xpb_out[91][362],u_xpb_out[92][362],u_xpb_out[93][362],u_xpb_out[94][362],u_xpb_out[95][362],u_xpb_out[96][362],u_xpb_out[97][362],u_xpb_out[98][362],u_xpb_out[99][362],u_xpb_out[100][362],u_xpb_out[101][362],u_xpb_out[102][362],u_xpb_out[103][362],u_xpb_out[104][362],u_xpb_out[105][362]};

assign col_out_363 = {u_xpb_out[0][363],u_xpb_out[1][363],u_xpb_out[2][363],u_xpb_out[3][363],u_xpb_out[4][363],u_xpb_out[5][363],u_xpb_out[6][363],u_xpb_out[7][363],u_xpb_out[8][363],u_xpb_out[9][363],u_xpb_out[10][363],u_xpb_out[11][363],u_xpb_out[12][363],u_xpb_out[13][363],u_xpb_out[14][363],u_xpb_out[15][363],u_xpb_out[16][363],u_xpb_out[17][363],u_xpb_out[18][363],u_xpb_out[19][363],u_xpb_out[20][363],u_xpb_out[21][363],u_xpb_out[22][363],u_xpb_out[23][363],u_xpb_out[24][363],u_xpb_out[25][363],u_xpb_out[26][363],u_xpb_out[27][363],u_xpb_out[28][363],u_xpb_out[29][363],u_xpb_out[30][363],u_xpb_out[31][363],u_xpb_out[32][363],u_xpb_out[33][363],u_xpb_out[34][363],u_xpb_out[35][363],u_xpb_out[36][363],u_xpb_out[37][363],u_xpb_out[38][363],u_xpb_out[39][363],u_xpb_out[40][363],u_xpb_out[41][363],u_xpb_out[42][363],u_xpb_out[43][363],u_xpb_out[44][363],u_xpb_out[45][363],u_xpb_out[46][363],u_xpb_out[47][363],u_xpb_out[48][363],u_xpb_out[49][363],u_xpb_out[50][363],u_xpb_out[51][363],u_xpb_out[52][363],u_xpb_out[53][363],u_xpb_out[54][363],u_xpb_out[55][363],u_xpb_out[56][363],u_xpb_out[57][363],u_xpb_out[58][363],u_xpb_out[59][363],u_xpb_out[60][363],u_xpb_out[61][363],u_xpb_out[62][363],u_xpb_out[63][363],u_xpb_out[64][363],u_xpb_out[65][363],u_xpb_out[66][363],u_xpb_out[67][363],u_xpb_out[68][363],u_xpb_out[69][363],u_xpb_out[70][363],u_xpb_out[71][363],u_xpb_out[72][363],u_xpb_out[73][363],u_xpb_out[74][363],u_xpb_out[75][363],u_xpb_out[76][363],u_xpb_out[77][363],u_xpb_out[78][363],u_xpb_out[79][363],u_xpb_out[80][363],u_xpb_out[81][363],u_xpb_out[82][363],u_xpb_out[83][363],u_xpb_out[84][363],u_xpb_out[85][363],u_xpb_out[86][363],u_xpb_out[87][363],u_xpb_out[88][363],u_xpb_out[89][363],u_xpb_out[90][363],u_xpb_out[91][363],u_xpb_out[92][363],u_xpb_out[93][363],u_xpb_out[94][363],u_xpb_out[95][363],u_xpb_out[96][363],u_xpb_out[97][363],u_xpb_out[98][363],u_xpb_out[99][363],u_xpb_out[100][363],u_xpb_out[101][363],u_xpb_out[102][363],u_xpb_out[103][363],u_xpb_out[104][363],u_xpb_out[105][363]};

assign col_out_364 = {u_xpb_out[0][364],u_xpb_out[1][364],u_xpb_out[2][364],u_xpb_out[3][364],u_xpb_out[4][364],u_xpb_out[5][364],u_xpb_out[6][364],u_xpb_out[7][364],u_xpb_out[8][364],u_xpb_out[9][364],u_xpb_out[10][364],u_xpb_out[11][364],u_xpb_out[12][364],u_xpb_out[13][364],u_xpb_out[14][364],u_xpb_out[15][364],u_xpb_out[16][364],u_xpb_out[17][364],u_xpb_out[18][364],u_xpb_out[19][364],u_xpb_out[20][364],u_xpb_out[21][364],u_xpb_out[22][364],u_xpb_out[23][364],u_xpb_out[24][364],u_xpb_out[25][364],u_xpb_out[26][364],u_xpb_out[27][364],u_xpb_out[28][364],u_xpb_out[29][364],u_xpb_out[30][364],u_xpb_out[31][364],u_xpb_out[32][364],u_xpb_out[33][364],u_xpb_out[34][364],u_xpb_out[35][364],u_xpb_out[36][364],u_xpb_out[37][364],u_xpb_out[38][364],u_xpb_out[39][364],u_xpb_out[40][364],u_xpb_out[41][364],u_xpb_out[42][364],u_xpb_out[43][364],u_xpb_out[44][364],u_xpb_out[45][364],u_xpb_out[46][364],u_xpb_out[47][364],u_xpb_out[48][364],u_xpb_out[49][364],u_xpb_out[50][364],u_xpb_out[51][364],u_xpb_out[52][364],u_xpb_out[53][364],u_xpb_out[54][364],u_xpb_out[55][364],u_xpb_out[56][364],u_xpb_out[57][364],u_xpb_out[58][364],u_xpb_out[59][364],u_xpb_out[60][364],u_xpb_out[61][364],u_xpb_out[62][364],u_xpb_out[63][364],u_xpb_out[64][364],u_xpb_out[65][364],u_xpb_out[66][364],u_xpb_out[67][364],u_xpb_out[68][364],u_xpb_out[69][364],u_xpb_out[70][364],u_xpb_out[71][364],u_xpb_out[72][364],u_xpb_out[73][364],u_xpb_out[74][364],u_xpb_out[75][364],u_xpb_out[76][364],u_xpb_out[77][364],u_xpb_out[78][364],u_xpb_out[79][364],u_xpb_out[80][364],u_xpb_out[81][364],u_xpb_out[82][364],u_xpb_out[83][364],u_xpb_out[84][364],u_xpb_out[85][364],u_xpb_out[86][364],u_xpb_out[87][364],u_xpb_out[88][364],u_xpb_out[89][364],u_xpb_out[90][364],u_xpb_out[91][364],u_xpb_out[92][364],u_xpb_out[93][364],u_xpb_out[94][364],u_xpb_out[95][364],u_xpb_out[96][364],u_xpb_out[97][364],u_xpb_out[98][364],u_xpb_out[99][364],u_xpb_out[100][364],u_xpb_out[101][364],u_xpb_out[102][364],u_xpb_out[103][364],u_xpb_out[104][364],u_xpb_out[105][364]};

assign col_out_365 = {u_xpb_out[0][365],u_xpb_out[1][365],u_xpb_out[2][365],u_xpb_out[3][365],u_xpb_out[4][365],u_xpb_out[5][365],u_xpb_out[6][365],u_xpb_out[7][365],u_xpb_out[8][365],u_xpb_out[9][365],u_xpb_out[10][365],u_xpb_out[11][365],u_xpb_out[12][365],u_xpb_out[13][365],u_xpb_out[14][365],u_xpb_out[15][365],u_xpb_out[16][365],u_xpb_out[17][365],u_xpb_out[18][365],u_xpb_out[19][365],u_xpb_out[20][365],u_xpb_out[21][365],u_xpb_out[22][365],u_xpb_out[23][365],u_xpb_out[24][365],u_xpb_out[25][365],u_xpb_out[26][365],u_xpb_out[27][365],u_xpb_out[28][365],u_xpb_out[29][365],u_xpb_out[30][365],u_xpb_out[31][365],u_xpb_out[32][365],u_xpb_out[33][365],u_xpb_out[34][365],u_xpb_out[35][365],u_xpb_out[36][365],u_xpb_out[37][365],u_xpb_out[38][365],u_xpb_out[39][365],u_xpb_out[40][365],u_xpb_out[41][365],u_xpb_out[42][365],u_xpb_out[43][365],u_xpb_out[44][365],u_xpb_out[45][365],u_xpb_out[46][365],u_xpb_out[47][365],u_xpb_out[48][365],u_xpb_out[49][365],u_xpb_out[50][365],u_xpb_out[51][365],u_xpb_out[52][365],u_xpb_out[53][365],u_xpb_out[54][365],u_xpb_out[55][365],u_xpb_out[56][365],u_xpb_out[57][365],u_xpb_out[58][365],u_xpb_out[59][365],u_xpb_out[60][365],u_xpb_out[61][365],u_xpb_out[62][365],u_xpb_out[63][365],u_xpb_out[64][365],u_xpb_out[65][365],u_xpb_out[66][365],u_xpb_out[67][365],u_xpb_out[68][365],u_xpb_out[69][365],u_xpb_out[70][365],u_xpb_out[71][365],u_xpb_out[72][365],u_xpb_out[73][365],u_xpb_out[74][365],u_xpb_out[75][365],u_xpb_out[76][365],u_xpb_out[77][365],u_xpb_out[78][365],u_xpb_out[79][365],u_xpb_out[80][365],u_xpb_out[81][365],u_xpb_out[82][365],u_xpb_out[83][365],u_xpb_out[84][365],u_xpb_out[85][365],u_xpb_out[86][365],u_xpb_out[87][365],u_xpb_out[88][365],u_xpb_out[89][365],u_xpb_out[90][365],u_xpb_out[91][365],u_xpb_out[92][365],u_xpb_out[93][365],u_xpb_out[94][365],u_xpb_out[95][365],u_xpb_out[96][365],u_xpb_out[97][365],u_xpb_out[98][365],u_xpb_out[99][365],u_xpb_out[100][365],u_xpb_out[101][365],u_xpb_out[102][365],u_xpb_out[103][365],u_xpb_out[104][365],u_xpb_out[105][365]};

assign col_out_366 = {u_xpb_out[0][366],u_xpb_out[1][366],u_xpb_out[2][366],u_xpb_out[3][366],u_xpb_out[4][366],u_xpb_out[5][366],u_xpb_out[6][366],u_xpb_out[7][366],u_xpb_out[8][366],u_xpb_out[9][366],u_xpb_out[10][366],u_xpb_out[11][366],u_xpb_out[12][366],u_xpb_out[13][366],u_xpb_out[14][366],u_xpb_out[15][366],u_xpb_out[16][366],u_xpb_out[17][366],u_xpb_out[18][366],u_xpb_out[19][366],u_xpb_out[20][366],u_xpb_out[21][366],u_xpb_out[22][366],u_xpb_out[23][366],u_xpb_out[24][366],u_xpb_out[25][366],u_xpb_out[26][366],u_xpb_out[27][366],u_xpb_out[28][366],u_xpb_out[29][366],u_xpb_out[30][366],u_xpb_out[31][366],u_xpb_out[32][366],u_xpb_out[33][366],u_xpb_out[34][366],u_xpb_out[35][366],u_xpb_out[36][366],u_xpb_out[37][366],u_xpb_out[38][366],u_xpb_out[39][366],u_xpb_out[40][366],u_xpb_out[41][366],u_xpb_out[42][366],u_xpb_out[43][366],u_xpb_out[44][366],u_xpb_out[45][366],u_xpb_out[46][366],u_xpb_out[47][366],u_xpb_out[48][366],u_xpb_out[49][366],u_xpb_out[50][366],u_xpb_out[51][366],u_xpb_out[52][366],u_xpb_out[53][366],u_xpb_out[54][366],u_xpb_out[55][366],u_xpb_out[56][366],u_xpb_out[57][366],u_xpb_out[58][366],u_xpb_out[59][366],u_xpb_out[60][366],u_xpb_out[61][366],u_xpb_out[62][366],u_xpb_out[63][366],u_xpb_out[64][366],u_xpb_out[65][366],u_xpb_out[66][366],u_xpb_out[67][366],u_xpb_out[68][366],u_xpb_out[69][366],u_xpb_out[70][366],u_xpb_out[71][366],u_xpb_out[72][366],u_xpb_out[73][366],u_xpb_out[74][366],u_xpb_out[75][366],u_xpb_out[76][366],u_xpb_out[77][366],u_xpb_out[78][366],u_xpb_out[79][366],u_xpb_out[80][366],u_xpb_out[81][366],u_xpb_out[82][366],u_xpb_out[83][366],u_xpb_out[84][366],u_xpb_out[85][366],u_xpb_out[86][366],u_xpb_out[87][366],u_xpb_out[88][366],u_xpb_out[89][366],u_xpb_out[90][366],u_xpb_out[91][366],u_xpb_out[92][366],u_xpb_out[93][366],u_xpb_out[94][366],u_xpb_out[95][366],u_xpb_out[96][366],u_xpb_out[97][366],u_xpb_out[98][366],u_xpb_out[99][366],u_xpb_out[100][366],u_xpb_out[101][366],u_xpb_out[102][366],u_xpb_out[103][366],u_xpb_out[104][366],u_xpb_out[105][366]};

assign col_out_367 = {u_xpb_out[0][367],u_xpb_out[1][367],u_xpb_out[2][367],u_xpb_out[3][367],u_xpb_out[4][367],u_xpb_out[5][367],u_xpb_out[6][367],u_xpb_out[7][367],u_xpb_out[8][367],u_xpb_out[9][367],u_xpb_out[10][367],u_xpb_out[11][367],u_xpb_out[12][367],u_xpb_out[13][367],u_xpb_out[14][367],u_xpb_out[15][367],u_xpb_out[16][367],u_xpb_out[17][367],u_xpb_out[18][367],u_xpb_out[19][367],u_xpb_out[20][367],u_xpb_out[21][367],u_xpb_out[22][367],u_xpb_out[23][367],u_xpb_out[24][367],u_xpb_out[25][367],u_xpb_out[26][367],u_xpb_out[27][367],u_xpb_out[28][367],u_xpb_out[29][367],u_xpb_out[30][367],u_xpb_out[31][367],u_xpb_out[32][367],u_xpb_out[33][367],u_xpb_out[34][367],u_xpb_out[35][367],u_xpb_out[36][367],u_xpb_out[37][367],u_xpb_out[38][367],u_xpb_out[39][367],u_xpb_out[40][367],u_xpb_out[41][367],u_xpb_out[42][367],u_xpb_out[43][367],u_xpb_out[44][367],u_xpb_out[45][367],u_xpb_out[46][367],u_xpb_out[47][367],u_xpb_out[48][367],u_xpb_out[49][367],u_xpb_out[50][367],u_xpb_out[51][367],u_xpb_out[52][367],u_xpb_out[53][367],u_xpb_out[54][367],u_xpb_out[55][367],u_xpb_out[56][367],u_xpb_out[57][367],u_xpb_out[58][367],u_xpb_out[59][367],u_xpb_out[60][367],u_xpb_out[61][367],u_xpb_out[62][367],u_xpb_out[63][367],u_xpb_out[64][367],u_xpb_out[65][367],u_xpb_out[66][367],u_xpb_out[67][367],u_xpb_out[68][367],u_xpb_out[69][367],u_xpb_out[70][367],u_xpb_out[71][367],u_xpb_out[72][367],u_xpb_out[73][367],u_xpb_out[74][367],u_xpb_out[75][367],u_xpb_out[76][367],u_xpb_out[77][367],u_xpb_out[78][367],u_xpb_out[79][367],u_xpb_out[80][367],u_xpb_out[81][367],u_xpb_out[82][367],u_xpb_out[83][367],u_xpb_out[84][367],u_xpb_out[85][367],u_xpb_out[86][367],u_xpb_out[87][367],u_xpb_out[88][367],u_xpb_out[89][367],u_xpb_out[90][367],u_xpb_out[91][367],u_xpb_out[92][367],u_xpb_out[93][367],u_xpb_out[94][367],u_xpb_out[95][367],u_xpb_out[96][367],u_xpb_out[97][367],u_xpb_out[98][367],u_xpb_out[99][367],u_xpb_out[100][367],u_xpb_out[101][367],u_xpb_out[102][367],u_xpb_out[103][367],u_xpb_out[104][367],u_xpb_out[105][367]};

assign col_out_368 = {u_xpb_out[0][368],u_xpb_out[1][368],u_xpb_out[2][368],u_xpb_out[3][368],u_xpb_out[4][368],u_xpb_out[5][368],u_xpb_out[6][368],u_xpb_out[7][368],u_xpb_out[8][368],u_xpb_out[9][368],u_xpb_out[10][368],u_xpb_out[11][368],u_xpb_out[12][368],u_xpb_out[13][368],u_xpb_out[14][368],u_xpb_out[15][368],u_xpb_out[16][368],u_xpb_out[17][368],u_xpb_out[18][368],u_xpb_out[19][368],u_xpb_out[20][368],u_xpb_out[21][368],u_xpb_out[22][368],u_xpb_out[23][368],u_xpb_out[24][368],u_xpb_out[25][368],u_xpb_out[26][368],u_xpb_out[27][368],u_xpb_out[28][368],u_xpb_out[29][368],u_xpb_out[30][368],u_xpb_out[31][368],u_xpb_out[32][368],u_xpb_out[33][368],u_xpb_out[34][368],u_xpb_out[35][368],u_xpb_out[36][368],u_xpb_out[37][368],u_xpb_out[38][368],u_xpb_out[39][368],u_xpb_out[40][368],u_xpb_out[41][368],u_xpb_out[42][368],u_xpb_out[43][368],u_xpb_out[44][368],u_xpb_out[45][368],u_xpb_out[46][368],u_xpb_out[47][368],u_xpb_out[48][368],u_xpb_out[49][368],u_xpb_out[50][368],u_xpb_out[51][368],u_xpb_out[52][368],u_xpb_out[53][368],u_xpb_out[54][368],u_xpb_out[55][368],u_xpb_out[56][368],u_xpb_out[57][368],u_xpb_out[58][368],u_xpb_out[59][368],u_xpb_out[60][368],u_xpb_out[61][368],u_xpb_out[62][368],u_xpb_out[63][368],u_xpb_out[64][368],u_xpb_out[65][368],u_xpb_out[66][368],u_xpb_out[67][368],u_xpb_out[68][368],u_xpb_out[69][368],u_xpb_out[70][368],u_xpb_out[71][368],u_xpb_out[72][368],u_xpb_out[73][368],u_xpb_out[74][368],u_xpb_out[75][368],u_xpb_out[76][368],u_xpb_out[77][368],u_xpb_out[78][368],u_xpb_out[79][368],u_xpb_out[80][368],u_xpb_out[81][368],u_xpb_out[82][368],u_xpb_out[83][368],u_xpb_out[84][368],u_xpb_out[85][368],u_xpb_out[86][368],u_xpb_out[87][368],u_xpb_out[88][368],u_xpb_out[89][368],u_xpb_out[90][368],u_xpb_out[91][368],u_xpb_out[92][368],u_xpb_out[93][368],u_xpb_out[94][368],u_xpb_out[95][368],u_xpb_out[96][368],u_xpb_out[97][368],u_xpb_out[98][368],u_xpb_out[99][368],u_xpb_out[100][368],u_xpb_out[101][368],u_xpb_out[102][368],u_xpb_out[103][368],u_xpb_out[104][368],u_xpb_out[105][368]};

assign col_out_369 = {u_xpb_out[0][369],u_xpb_out[1][369],u_xpb_out[2][369],u_xpb_out[3][369],u_xpb_out[4][369],u_xpb_out[5][369],u_xpb_out[6][369],u_xpb_out[7][369],u_xpb_out[8][369],u_xpb_out[9][369],u_xpb_out[10][369],u_xpb_out[11][369],u_xpb_out[12][369],u_xpb_out[13][369],u_xpb_out[14][369],u_xpb_out[15][369],u_xpb_out[16][369],u_xpb_out[17][369],u_xpb_out[18][369],u_xpb_out[19][369],u_xpb_out[20][369],u_xpb_out[21][369],u_xpb_out[22][369],u_xpb_out[23][369],u_xpb_out[24][369],u_xpb_out[25][369],u_xpb_out[26][369],u_xpb_out[27][369],u_xpb_out[28][369],u_xpb_out[29][369],u_xpb_out[30][369],u_xpb_out[31][369],u_xpb_out[32][369],u_xpb_out[33][369],u_xpb_out[34][369],u_xpb_out[35][369],u_xpb_out[36][369],u_xpb_out[37][369],u_xpb_out[38][369],u_xpb_out[39][369],u_xpb_out[40][369],u_xpb_out[41][369],u_xpb_out[42][369],u_xpb_out[43][369],u_xpb_out[44][369],u_xpb_out[45][369],u_xpb_out[46][369],u_xpb_out[47][369],u_xpb_out[48][369],u_xpb_out[49][369],u_xpb_out[50][369],u_xpb_out[51][369],u_xpb_out[52][369],u_xpb_out[53][369],u_xpb_out[54][369],u_xpb_out[55][369],u_xpb_out[56][369],u_xpb_out[57][369],u_xpb_out[58][369],u_xpb_out[59][369],u_xpb_out[60][369],u_xpb_out[61][369],u_xpb_out[62][369],u_xpb_out[63][369],u_xpb_out[64][369],u_xpb_out[65][369],u_xpb_out[66][369],u_xpb_out[67][369],u_xpb_out[68][369],u_xpb_out[69][369],u_xpb_out[70][369],u_xpb_out[71][369],u_xpb_out[72][369],u_xpb_out[73][369],u_xpb_out[74][369],u_xpb_out[75][369],u_xpb_out[76][369],u_xpb_out[77][369],u_xpb_out[78][369],u_xpb_out[79][369],u_xpb_out[80][369],u_xpb_out[81][369],u_xpb_out[82][369],u_xpb_out[83][369],u_xpb_out[84][369],u_xpb_out[85][369],u_xpb_out[86][369],u_xpb_out[87][369],u_xpb_out[88][369],u_xpb_out[89][369],u_xpb_out[90][369],u_xpb_out[91][369],u_xpb_out[92][369],u_xpb_out[93][369],u_xpb_out[94][369],u_xpb_out[95][369],u_xpb_out[96][369],u_xpb_out[97][369],u_xpb_out[98][369],u_xpb_out[99][369],u_xpb_out[100][369],u_xpb_out[101][369],u_xpb_out[102][369],u_xpb_out[103][369],u_xpb_out[104][369],u_xpb_out[105][369]};

assign col_out_370 = {u_xpb_out[0][370],u_xpb_out[1][370],u_xpb_out[2][370],u_xpb_out[3][370],u_xpb_out[4][370],u_xpb_out[5][370],u_xpb_out[6][370],u_xpb_out[7][370],u_xpb_out[8][370],u_xpb_out[9][370],u_xpb_out[10][370],u_xpb_out[11][370],u_xpb_out[12][370],u_xpb_out[13][370],u_xpb_out[14][370],u_xpb_out[15][370],u_xpb_out[16][370],u_xpb_out[17][370],u_xpb_out[18][370],u_xpb_out[19][370],u_xpb_out[20][370],u_xpb_out[21][370],u_xpb_out[22][370],u_xpb_out[23][370],u_xpb_out[24][370],u_xpb_out[25][370],u_xpb_out[26][370],u_xpb_out[27][370],u_xpb_out[28][370],u_xpb_out[29][370],u_xpb_out[30][370],u_xpb_out[31][370],u_xpb_out[32][370],u_xpb_out[33][370],u_xpb_out[34][370],u_xpb_out[35][370],u_xpb_out[36][370],u_xpb_out[37][370],u_xpb_out[38][370],u_xpb_out[39][370],u_xpb_out[40][370],u_xpb_out[41][370],u_xpb_out[42][370],u_xpb_out[43][370],u_xpb_out[44][370],u_xpb_out[45][370],u_xpb_out[46][370],u_xpb_out[47][370],u_xpb_out[48][370],u_xpb_out[49][370],u_xpb_out[50][370],u_xpb_out[51][370],u_xpb_out[52][370],u_xpb_out[53][370],u_xpb_out[54][370],u_xpb_out[55][370],u_xpb_out[56][370],u_xpb_out[57][370],u_xpb_out[58][370],u_xpb_out[59][370],u_xpb_out[60][370],u_xpb_out[61][370],u_xpb_out[62][370],u_xpb_out[63][370],u_xpb_out[64][370],u_xpb_out[65][370],u_xpb_out[66][370],u_xpb_out[67][370],u_xpb_out[68][370],u_xpb_out[69][370],u_xpb_out[70][370],u_xpb_out[71][370],u_xpb_out[72][370],u_xpb_out[73][370],u_xpb_out[74][370],u_xpb_out[75][370],u_xpb_out[76][370],u_xpb_out[77][370],u_xpb_out[78][370],u_xpb_out[79][370],u_xpb_out[80][370],u_xpb_out[81][370],u_xpb_out[82][370],u_xpb_out[83][370],u_xpb_out[84][370],u_xpb_out[85][370],u_xpb_out[86][370],u_xpb_out[87][370],u_xpb_out[88][370],u_xpb_out[89][370],u_xpb_out[90][370],u_xpb_out[91][370],u_xpb_out[92][370],u_xpb_out[93][370],u_xpb_out[94][370],u_xpb_out[95][370],u_xpb_out[96][370],u_xpb_out[97][370],u_xpb_out[98][370],u_xpb_out[99][370],u_xpb_out[100][370],u_xpb_out[101][370],u_xpb_out[102][370],u_xpb_out[103][370],u_xpb_out[104][370],u_xpb_out[105][370]};

assign col_out_371 = {u_xpb_out[0][371],u_xpb_out[1][371],u_xpb_out[2][371],u_xpb_out[3][371],u_xpb_out[4][371],u_xpb_out[5][371],u_xpb_out[6][371],u_xpb_out[7][371],u_xpb_out[8][371],u_xpb_out[9][371],u_xpb_out[10][371],u_xpb_out[11][371],u_xpb_out[12][371],u_xpb_out[13][371],u_xpb_out[14][371],u_xpb_out[15][371],u_xpb_out[16][371],u_xpb_out[17][371],u_xpb_out[18][371],u_xpb_out[19][371],u_xpb_out[20][371],u_xpb_out[21][371],u_xpb_out[22][371],u_xpb_out[23][371],u_xpb_out[24][371],u_xpb_out[25][371],u_xpb_out[26][371],u_xpb_out[27][371],u_xpb_out[28][371],u_xpb_out[29][371],u_xpb_out[30][371],u_xpb_out[31][371],u_xpb_out[32][371],u_xpb_out[33][371],u_xpb_out[34][371],u_xpb_out[35][371],u_xpb_out[36][371],u_xpb_out[37][371],u_xpb_out[38][371],u_xpb_out[39][371],u_xpb_out[40][371],u_xpb_out[41][371],u_xpb_out[42][371],u_xpb_out[43][371],u_xpb_out[44][371],u_xpb_out[45][371],u_xpb_out[46][371],u_xpb_out[47][371],u_xpb_out[48][371],u_xpb_out[49][371],u_xpb_out[50][371],u_xpb_out[51][371],u_xpb_out[52][371],u_xpb_out[53][371],u_xpb_out[54][371],u_xpb_out[55][371],u_xpb_out[56][371],u_xpb_out[57][371],u_xpb_out[58][371],u_xpb_out[59][371],u_xpb_out[60][371],u_xpb_out[61][371],u_xpb_out[62][371],u_xpb_out[63][371],u_xpb_out[64][371],u_xpb_out[65][371],u_xpb_out[66][371],u_xpb_out[67][371],u_xpb_out[68][371],u_xpb_out[69][371],u_xpb_out[70][371],u_xpb_out[71][371],u_xpb_out[72][371],u_xpb_out[73][371],u_xpb_out[74][371],u_xpb_out[75][371],u_xpb_out[76][371],u_xpb_out[77][371],u_xpb_out[78][371],u_xpb_out[79][371],u_xpb_out[80][371],u_xpb_out[81][371],u_xpb_out[82][371],u_xpb_out[83][371],u_xpb_out[84][371],u_xpb_out[85][371],u_xpb_out[86][371],u_xpb_out[87][371],u_xpb_out[88][371],u_xpb_out[89][371],u_xpb_out[90][371],u_xpb_out[91][371],u_xpb_out[92][371],u_xpb_out[93][371],u_xpb_out[94][371],u_xpb_out[95][371],u_xpb_out[96][371],u_xpb_out[97][371],u_xpb_out[98][371],u_xpb_out[99][371],u_xpb_out[100][371],u_xpb_out[101][371],u_xpb_out[102][371],u_xpb_out[103][371],u_xpb_out[104][371],u_xpb_out[105][371]};

assign col_out_372 = {u_xpb_out[0][372],u_xpb_out[1][372],u_xpb_out[2][372],u_xpb_out[3][372],u_xpb_out[4][372],u_xpb_out[5][372],u_xpb_out[6][372],u_xpb_out[7][372],u_xpb_out[8][372],u_xpb_out[9][372],u_xpb_out[10][372],u_xpb_out[11][372],u_xpb_out[12][372],u_xpb_out[13][372],u_xpb_out[14][372],u_xpb_out[15][372],u_xpb_out[16][372],u_xpb_out[17][372],u_xpb_out[18][372],u_xpb_out[19][372],u_xpb_out[20][372],u_xpb_out[21][372],u_xpb_out[22][372],u_xpb_out[23][372],u_xpb_out[24][372],u_xpb_out[25][372],u_xpb_out[26][372],u_xpb_out[27][372],u_xpb_out[28][372],u_xpb_out[29][372],u_xpb_out[30][372],u_xpb_out[31][372],u_xpb_out[32][372],u_xpb_out[33][372],u_xpb_out[34][372],u_xpb_out[35][372],u_xpb_out[36][372],u_xpb_out[37][372],u_xpb_out[38][372],u_xpb_out[39][372],u_xpb_out[40][372],u_xpb_out[41][372],u_xpb_out[42][372],u_xpb_out[43][372],u_xpb_out[44][372],u_xpb_out[45][372],u_xpb_out[46][372],u_xpb_out[47][372],u_xpb_out[48][372],u_xpb_out[49][372],u_xpb_out[50][372],u_xpb_out[51][372],u_xpb_out[52][372],u_xpb_out[53][372],u_xpb_out[54][372],u_xpb_out[55][372],u_xpb_out[56][372],u_xpb_out[57][372],u_xpb_out[58][372],u_xpb_out[59][372],u_xpb_out[60][372],u_xpb_out[61][372],u_xpb_out[62][372],u_xpb_out[63][372],u_xpb_out[64][372],u_xpb_out[65][372],u_xpb_out[66][372],u_xpb_out[67][372],u_xpb_out[68][372],u_xpb_out[69][372],u_xpb_out[70][372],u_xpb_out[71][372],u_xpb_out[72][372],u_xpb_out[73][372],u_xpb_out[74][372],u_xpb_out[75][372],u_xpb_out[76][372],u_xpb_out[77][372],u_xpb_out[78][372],u_xpb_out[79][372],u_xpb_out[80][372],u_xpb_out[81][372],u_xpb_out[82][372],u_xpb_out[83][372],u_xpb_out[84][372],u_xpb_out[85][372],u_xpb_out[86][372],u_xpb_out[87][372],u_xpb_out[88][372],u_xpb_out[89][372],u_xpb_out[90][372],u_xpb_out[91][372],u_xpb_out[92][372],u_xpb_out[93][372],u_xpb_out[94][372],u_xpb_out[95][372],u_xpb_out[96][372],u_xpb_out[97][372],u_xpb_out[98][372],u_xpb_out[99][372],u_xpb_out[100][372],u_xpb_out[101][372],u_xpb_out[102][372],u_xpb_out[103][372],u_xpb_out[104][372],u_xpb_out[105][372]};

assign col_out_373 = {u_xpb_out[0][373],u_xpb_out[1][373],u_xpb_out[2][373],u_xpb_out[3][373],u_xpb_out[4][373],u_xpb_out[5][373],u_xpb_out[6][373],u_xpb_out[7][373],u_xpb_out[8][373],u_xpb_out[9][373],u_xpb_out[10][373],u_xpb_out[11][373],u_xpb_out[12][373],u_xpb_out[13][373],u_xpb_out[14][373],u_xpb_out[15][373],u_xpb_out[16][373],u_xpb_out[17][373],u_xpb_out[18][373],u_xpb_out[19][373],u_xpb_out[20][373],u_xpb_out[21][373],u_xpb_out[22][373],u_xpb_out[23][373],u_xpb_out[24][373],u_xpb_out[25][373],u_xpb_out[26][373],u_xpb_out[27][373],u_xpb_out[28][373],u_xpb_out[29][373],u_xpb_out[30][373],u_xpb_out[31][373],u_xpb_out[32][373],u_xpb_out[33][373],u_xpb_out[34][373],u_xpb_out[35][373],u_xpb_out[36][373],u_xpb_out[37][373],u_xpb_out[38][373],u_xpb_out[39][373],u_xpb_out[40][373],u_xpb_out[41][373],u_xpb_out[42][373],u_xpb_out[43][373],u_xpb_out[44][373],u_xpb_out[45][373],u_xpb_out[46][373],u_xpb_out[47][373],u_xpb_out[48][373],u_xpb_out[49][373],u_xpb_out[50][373],u_xpb_out[51][373],u_xpb_out[52][373],u_xpb_out[53][373],u_xpb_out[54][373],u_xpb_out[55][373],u_xpb_out[56][373],u_xpb_out[57][373],u_xpb_out[58][373],u_xpb_out[59][373],u_xpb_out[60][373],u_xpb_out[61][373],u_xpb_out[62][373],u_xpb_out[63][373],u_xpb_out[64][373],u_xpb_out[65][373],u_xpb_out[66][373],u_xpb_out[67][373],u_xpb_out[68][373],u_xpb_out[69][373],u_xpb_out[70][373],u_xpb_out[71][373],u_xpb_out[72][373],u_xpb_out[73][373],u_xpb_out[74][373],u_xpb_out[75][373],u_xpb_out[76][373],u_xpb_out[77][373],u_xpb_out[78][373],u_xpb_out[79][373],u_xpb_out[80][373],u_xpb_out[81][373],u_xpb_out[82][373],u_xpb_out[83][373],u_xpb_out[84][373],u_xpb_out[85][373],u_xpb_out[86][373],u_xpb_out[87][373],u_xpb_out[88][373],u_xpb_out[89][373],u_xpb_out[90][373],u_xpb_out[91][373],u_xpb_out[92][373],u_xpb_out[93][373],u_xpb_out[94][373],u_xpb_out[95][373],u_xpb_out[96][373],u_xpb_out[97][373],u_xpb_out[98][373],u_xpb_out[99][373],u_xpb_out[100][373],u_xpb_out[101][373],u_xpb_out[102][373],u_xpb_out[103][373],u_xpb_out[104][373],u_xpb_out[105][373]};

assign col_out_374 = {u_xpb_out[0][374],u_xpb_out[1][374],u_xpb_out[2][374],u_xpb_out[3][374],u_xpb_out[4][374],u_xpb_out[5][374],u_xpb_out[6][374],u_xpb_out[7][374],u_xpb_out[8][374],u_xpb_out[9][374],u_xpb_out[10][374],u_xpb_out[11][374],u_xpb_out[12][374],u_xpb_out[13][374],u_xpb_out[14][374],u_xpb_out[15][374],u_xpb_out[16][374],u_xpb_out[17][374],u_xpb_out[18][374],u_xpb_out[19][374],u_xpb_out[20][374],u_xpb_out[21][374],u_xpb_out[22][374],u_xpb_out[23][374],u_xpb_out[24][374],u_xpb_out[25][374],u_xpb_out[26][374],u_xpb_out[27][374],u_xpb_out[28][374],u_xpb_out[29][374],u_xpb_out[30][374],u_xpb_out[31][374],u_xpb_out[32][374],u_xpb_out[33][374],u_xpb_out[34][374],u_xpb_out[35][374],u_xpb_out[36][374],u_xpb_out[37][374],u_xpb_out[38][374],u_xpb_out[39][374],u_xpb_out[40][374],u_xpb_out[41][374],u_xpb_out[42][374],u_xpb_out[43][374],u_xpb_out[44][374],u_xpb_out[45][374],u_xpb_out[46][374],u_xpb_out[47][374],u_xpb_out[48][374],u_xpb_out[49][374],u_xpb_out[50][374],u_xpb_out[51][374],u_xpb_out[52][374],u_xpb_out[53][374],u_xpb_out[54][374],u_xpb_out[55][374],u_xpb_out[56][374],u_xpb_out[57][374],u_xpb_out[58][374],u_xpb_out[59][374],u_xpb_out[60][374],u_xpb_out[61][374],u_xpb_out[62][374],u_xpb_out[63][374],u_xpb_out[64][374],u_xpb_out[65][374],u_xpb_out[66][374],u_xpb_out[67][374],u_xpb_out[68][374],u_xpb_out[69][374],u_xpb_out[70][374],u_xpb_out[71][374],u_xpb_out[72][374],u_xpb_out[73][374],u_xpb_out[74][374],u_xpb_out[75][374],u_xpb_out[76][374],u_xpb_out[77][374],u_xpb_out[78][374],u_xpb_out[79][374],u_xpb_out[80][374],u_xpb_out[81][374],u_xpb_out[82][374],u_xpb_out[83][374],u_xpb_out[84][374],u_xpb_out[85][374],u_xpb_out[86][374],u_xpb_out[87][374],u_xpb_out[88][374],u_xpb_out[89][374],u_xpb_out[90][374],u_xpb_out[91][374],u_xpb_out[92][374],u_xpb_out[93][374],u_xpb_out[94][374],u_xpb_out[95][374],u_xpb_out[96][374],u_xpb_out[97][374],u_xpb_out[98][374],u_xpb_out[99][374],u_xpb_out[100][374],u_xpb_out[101][374],u_xpb_out[102][374],u_xpb_out[103][374],u_xpb_out[104][374],u_xpb_out[105][374]};

assign col_out_375 = {u_xpb_out[0][375],u_xpb_out[1][375],u_xpb_out[2][375],u_xpb_out[3][375],u_xpb_out[4][375],u_xpb_out[5][375],u_xpb_out[6][375],u_xpb_out[7][375],u_xpb_out[8][375],u_xpb_out[9][375],u_xpb_out[10][375],u_xpb_out[11][375],u_xpb_out[12][375],u_xpb_out[13][375],u_xpb_out[14][375],u_xpb_out[15][375],u_xpb_out[16][375],u_xpb_out[17][375],u_xpb_out[18][375],u_xpb_out[19][375],u_xpb_out[20][375],u_xpb_out[21][375],u_xpb_out[22][375],u_xpb_out[23][375],u_xpb_out[24][375],u_xpb_out[25][375],u_xpb_out[26][375],u_xpb_out[27][375],u_xpb_out[28][375],u_xpb_out[29][375],u_xpb_out[30][375],u_xpb_out[31][375],u_xpb_out[32][375],u_xpb_out[33][375],u_xpb_out[34][375],u_xpb_out[35][375],u_xpb_out[36][375],u_xpb_out[37][375],u_xpb_out[38][375],u_xpb_out[39][375],u_xpb_out[40][375],u_xpb_out[41][375],u_xpb_out[42][375],u_xpb_out[43][375],u_xpb_out[44][375],u_xpb_out[45][375],u_xpb_out[46][375],u_xpb_out[47][375],u_xpb_out[48][375],u_xpb_out[49][375],u_xpb_out[50][375],u_xpb_out[51][375],u_xpb_out[52][375],u_xpb_out[53][375],u_xpb_out[54][375],u_xpb_out[55][375],u_xpb_out[56][375],u_xpb_out[57][375],u_xpb_out[58][375],u_xpb_out[59][375],u_xpb_out[60][375],u_xpb_out[61][375],u_xpb_out[62][375],u_xpb_out[63][375],u_xpb_out[64][375],u_xpb_out[65][375],u_xpb_out[66][375],u_xpb_out[67][375],u_xpb_out[68][375],u_xpb_out[69][375],u_xpb_out[70][375],u_xpb_out[71][375],u_xpb_out[72][375],u_xpb_out[73][375],u_xpb_out[74][375],u_xpb_out[75][375],u_xpb_out[76][375],u_xpb_out[77][375],u_xpb_out[78][375],u_xpb_out[79][375],u_xpb_out[80][375],u_xpb_out[81][375],u_xpb_out[82][375],u_xpb_out[83][375],u_xpb_out[84][375],u_xpb_out[85][375],u_xpb_out[86][375],u_xpb_out[87][375],u_xpb_out[88][375],u_xpb_out[89][375],u_xpb_out[90][375],u_xpb_out[91][375],u_xpb_out[92][375],u_xpb_out[93][375],u_xpb_out[94][375],u_xpb_out[95][375],u_xpb_out[96][375],u_xpb_out[97][375],u_xpb_out[98][375],u_xpb_out[99][375],u_xpb_out[100][375],u_xpb_out[101][375],u_xpb_out[102][375],u_xpb_out[103][375],u_xpb_out[104][375],u_xpb_out[105][375]};

assign col_out_376 = {u_xpb_out[0][376],u_xpb_out[1][376],u_xpb_out[2][376],u_xpb_out[3][376],u_xpb_out[4][376],u_xpb_out[5][376],u_xpb_out[6][376],u_xpb_out[7][376],u_xpb_out[8][376],u_xpb_out[9][376],u_xpb_out[10][376],u_xpb_out[11][376],u_xpb_out[12][376],u_xpb_out[13][376],u_xpb_out[14][376],u_xpb_out[15][376],u_xpb_out[16][376],u_xpb_out[17][376],u_xpb_out[18][376],u_xpb_out[19][376],u_xpb_out[20][376],u_xpb_out[21][376],u_xpb_out[22][376],u_xpb_out[23][376],u_xpb_out[24][376],u_xpb_out[25][376],u_xpb_out[26][376],u_xpb_out[27][376],u_xpb_out[28][376],u_xpb_out[29][376],u_xpb_out[30][376],u_xpb_out[31][376],u_xpb_out[32][376],u_xpb_out[33][376],u_xpb_out[34][376],u_xpb_out[35][376],u_xpb_out[36][376],u_xpb_out[37][376],u_xpb_out[38][376],u_xpb_out[39][376],u_xpb_out[40][376],u_xpb_out[41][376],u_xpb_out[42][376],u_xpb_out[43][376],u_xpb_out[44][376],u_xpb_out[45][376],u_xpb_out[46][376],u_xpb_out[47][376],u_xpb_out[48][376],u_xpb_out[49][376],u_xpb_out[50][376],u_xpb_out[51][376],u_xpb_out[52][376],u_xpb_out[53][376],u_xpb_out[54][376],u_xpb_out[55][376],u_xpb_out[56][376],u_xpb_out[57][376],u_xpb_out[58][376],u_xpb_out[59][376],u_xpb_out[60][376],u_xpb_out[61][376],u_xpb_out[62][376],u_xpb_out[63][376],u_xpb_out[64][376],u_xpb_out[65][376],u_xpb_out[66][376],u_xpb_out[67][376],u_xpb_out[68][376],u_xpb_out[69][376],u_xpb_out[70][376],u_xpb_out[71][376],u_xpb_out[72][376],u_xpb_out[73][376],u_xpb_out[74][376],u_xpb_out[75][376],u_xpb_out[76][376],u_xpb_out[77][376],u_xpb_out[78][376],u_xpb_out[79][376],u_xpb_out[80][376],u_xpb_out[81][376],u_xpb_out[82][376],u_xpb_out[83][376],u_xpb_out[84][376],u_xpb_out[85][376],u_xpb_out[86][376],u_xpb_out[87][376],u_xpb_out[88][376],u_xpb_out[89][376],u_xpb_out[90][376],u_xpb_out[91][376],u_xpb_out[92][376],u_xpb_out[93][376],u_xpb_out[94][376],u_xpb_out[95][376],u_xpb_out[96][376],u_xpb_out[97][376],u_xpb_out[98][376],u_xpb_out[99][376],u_xpb_out[100][376],u_xpb_out[101][376],u_xpb_out[102][376],u_xpb_out[103][376],u_xpb_out[104][376],u_xpb_out[105][376]};

assign col_out_377 = {u_xpb_out[0][377],u_xpb_out[1][377],u_xpb_out[2][377],u_xpb_out[3][377],u_xpb_out[4][377],u_xpb_out[5][377],u_xpb_out[6][377],u_xpb_out[7][377],u_xpb_out[8][377],u_xpb_out[9][377],u_xpb_out[10][377],u_xpb_out[11][377],u_xpb_out[12][377],u_xpb_out[13][377],u_xpb_out[14][377],u_xpb_out[15][377],u_xpb_out[16][377],u_xpb_out[17][377],u_xpb_out[18][377],u_xpb_out[19][377],u_xpb_out[20][377],u_xpb_out[21][377],u_xpb_out[22][377],u_xpb_out[23][377],u_xpb_out[24][377],u_xpb_out[25][377],u_xpb_out[26][377],u_xpb_out[27][377],u_xpb_out[28][377],u_xpb_out[29][377],u_xpb_out[30][377],u_xpb_out[31][377],u_xpb_out[32][377],u_xpb_out[33][377],u_xpb_out[34][377],u_xpb_out[35][377],u_xpb_out[36][377],u_xpb_out[37][377],u_xpb_out[38][377],u_xpb_out[39][377],u_xpb_out[40][377],u_xpb_out[41][377],u_xpb_out[42][377],u_xpb_out[43][377],u_xpb_out[44][377],u_xpb_out[45][377],u_xpb_out[46][377],u_xpb_out[47][377],u_xpb_out[48][377],u_xpb_out[49][377],u_xpb_out[50][377],u_xpb_out[51][377],u_xpb_out[52][377],u_xpb_out[53][377],u_xpb_out[54][377],u_xpb_out[55][377],u_xpb_out[56][377],u_xpb_out[57][377],u_xpb_out[58][377],u_xpb_out[59][377],u_xpb_out[60][377],u_xpb_out[61][377],u_xpb_out[62][377],u_xpb_out[63][377],u_xpb_out[64][377],u_xpb_out[65][377],u_xpb_out[66][377],u_xpb_out[67][377],u_xpb_out[68][377],u_xpb_out[69][377],u_xpb_out[70][377],u_xpb_out[71][377],u_xpb_out[72][377],u_xpb_out[73][377],u_xpb_out[74][377],u_xpb_out[75][377],u_xpb_out[76][377],u_xpb_out[77][377],u_xpb_out[78][377],u_xpb_out[79][377],u_xpb_out[80][377],u_xpb_out[81][377],u_xpb_out[82][377],u_xpb_out[83][377],u_xpb_out[84][377],u_xpb_out[85][377],u_xpb_out[86][377],u_xpb_out[87][377],u_xpb_out[88][377],u_xpb_out[89][377],u_xpb_out[90][377],u_xpb_out[91][377],u_xpb_out[92][377],u_xpb_out[93][377],u_xpb_out[94][377],u_xpb_out[95][377],u_xpb_out[96][377],u_xpb_out[97][377],u_xpb_out[98][377],u_xpb_out[99][377],u_xpb_out[100][377],u_xpb_out[101][377],u_xpb_out[102][377],u_xpb_out[103][377],u_xpb_out[104][377],u_xpb_out[105][377]};

assign col_out_378 = {u_xpb_out[0][378],u_xpb_out[1][378],u_xpb_out[2][378],u_xpb_out[3][378],u_xpb_out[4][378],u_xpb_out[5][378],u_xpb_out[6][378],u_xpb_out[7][378],u_xpb_out[8][378],u_xpb_out[9][378],u_xpb_out[10][378],u_xpb_out[11][378],u_xpb_out[12][378],u_xpb_out[13][378],u_xpb_out[14][378],u_xpb_out[15][378],u_xpb_out[16][378],u_xpb_out[17][378],u_xpb_out[18][378],u_xpb_out[19][378],u_xpb_out[20][378],u_xpb_out[21][378],u_xpb_out[22][378],u_xpb_out[23][378],u_xpb_out[24][378],u_xpb_out[25][378],u_xpb_out[26][378],u_xpb_out[27][378],u_xpb_out[28][378],u_xpb_out[29][378],u_xpb_out[30][378],u_xpb_out[31][378],u_xpb_out[32][378],u_xpb_out[33][378],u_xpb_out[34][378],u_xpb_out[35][378],u_xpb_out[36][378],u_xpb_out[37][378],u_xpb_out[38][378],u_xpb_out[39][378],u_xpb_out[40][378],u_xpb_out[41][378],u_xpb_out[42][378],u_xpb_out[43][378],u_xpb_out[44][378],u_xpb_out[45][378],u_xpb_out[46][378],u_xpb_out[47][378],u_xpb_out[48][378],u_xpb_out[49][378],u_xpb_out[50][378],u_xpb_out[51][378],u_xpb_out[52][378],u_xpb_out[53][378],u_xpb_out[54][378],u_xpb_out[55][378],u_xpb_out[56][378],u_xpb_out[57][378],u_xpb_out[58][378],u_xpb_out[59][378],u_xpb_out[60][378],u_xpb_out[61][378],u_xpb_out[62][378],u_xpb_out[63][378],u_xpb_out[64][378],u_xpb_out[65][378],u_xpb_out[66][378],u_xpb_out[67][378],u_xpb_out[68][378],u_xpb_out[69][378],u_xpb_out[70][378],u_xpb_out[71][378],u_xpb_out[72][378],u_xpb_out[73][378],u_xpb_out[74][378],u_xpb_out[75][378],u_xpb_out[76][378],u_xpb_out[77][378],u_xpb_out[78][378],u_xpb_out[79][378],u_xpb_out[80][378],u_xpb_out[81][378],u_xpb_out[82][378],u_xpb_out[83][378],u_xpb_out[84][378],u_xpb_out[85][378],u_xpb_out[86][378],u_xpb_out[87][378],u_xpb_out[88][378],u_xpb_out[89][378],u_xpb_out[90][378],u_xpb_out[91][378],u_xpb_out[92][378],u_xpb_out[93][378],u_xpb_out[94][378],u_xpb_out[95][378],u_xpb_out[96][378],u_xpb_out[97][378],u_xpb_out[98][378],u_xpb_out[99][378],u_xpb_out[100][378],u_xpb_out[101][378],u_xpb_out[102][378],u_xpb_out[103][378],u_xpb_out[104][378],u_xpb_out[105][378]};

assign col_out_379 = {u_xpb_out[0][379],u_xpb_out[1][379],u_xpb_out[2][379],u_xpb_out[3][379],u_xpb_out[4][379],u_xpb_out[5][379],u_xpb_out[6][379],u_xpb_out[7][379],u_xpb_out[8][379],u_xpb_out[9][379],u_xpb_out[10][379],u_xpb_out[11][379],u_xpb_out[12][379],u_xpb_out[13][379],u_xpb_out[14][379],u_xpb_out[15][379],u_xpb_out[16][379],u_xpb_out[17][379],u_xpb_out[18][379],u_xpb_out[19][379],u_xpb_out[20][379],u_xpb_out[21][379],u_xpb_out[22][379],u_xpb_out[23][379],u_xpb_out[24][379],u_xpb_out[25][379],u_xpb_out[26][379],u_xpb_out[27][379],u_xpb_out[28][379],u_xpb_out[29][379],u_xpb_out[30][379],u_xpb_out[31][379],u_xpb_out[32][379],u_xpb_out[33][379],u_xpb_out[34][379],u_xpb_out[35][379],u_xpb_out[36][379],u_xpb_out[37][379],u_xpb_out[38][379],u_xpb_out[39][379],u_xpb_out[40][379],u_xpb_out[41][379],u_xpb_out[42][379],u_xpb_out[43][379],u_xpb_out[44][379],u_xpb_out[45][379],u_xpb_out[46][379],u_xpb_out[47][379],u_xpb_out[48][379],u_xpb_out[49][379],u_xpb_out[50][379],u_xpb_out[51][379],u_xpb_out[52][379],u_xpb_out[53][379],u_xpb_out[54][379],u_xpb_out[55][379],u_xpb_out[56][379],u_xpb_out[57][379],u_xpb_out[58][379],u_xpb_out[59][379],u_xpb_out[60][379],u_xpb_out[61][379],u_xpb_out[62][379],u_xpb_out[63][379],u_xpb_out[64][379],u_xpb_out[65][379],u_xpb_out[66][379],u_xpb_out[67][379],u_xpb_out[68][379],u_xpb_out[69][379],u_xpb_out[70][379],u_xpb_out[71][379],u_xpb_out[72][379],u_xpb_out[73][379],u_xpb_out[74][379],u_xpb_out[75][379],u_xpb_out[76][379],u_xpb_out[77][379],u_xpb_out[78][379],u_xpb_out[79][379],u_xpb_out[80][379],u_xpb_out[81][379],u_xpb_out[82][379],u_xpb_out[83][379],u_xpb_out[84][379],u_xpb_out[85][379],u_xpb_out[86][379],u_xpb_out[87][379],u_xpb_out[88][379],u_xpb_out[89][379],u_xpb_out[90][379],u_xpb_out[91][379],u_xpb_out[92][379],u_xpb_out[93][379],u_xpb_out[94][379],u_xpb_out[95][379],u_xpb_out[96][379],u_xpb_out[97][379],u_xpb_out[98][379],u_xpb_out[99][379],u_xpb_out[100][379],u_xpb_out[101][379],u_xpb_out[102][379],u_xpb_out[103][379],u_xpb_out[104][379],u_xpb_out[105][379]};

assign col_out_380 = {u_xpb_out[0][380],u_xpb_out[1][380],u_xpb_out[2][380],u_xpb_out[3][380],u_xpb_out[4][380],u_xpb_out[5][380],u_xpb_out[6][380],u_xpb_out[7][380],u_xpb_out[8][380],u_xpb_out[9][380],u_xpb_out[10][380],u_xpb_out[11][380],u_xpb_out[12][380],u_xpb_out[13][380],u_xpb_out[14][380],u_xpb_out[15][380],u_xpb_out[16][380],u_xpb_out[17][380],u_xpb_out[18][380],u_xpb_out[19][380],u_xpb_out[20][380],u_xpb_out[21][380],u_xpb_out[22][380],u_xpb_out[23][380],u_xpb_out[24][380],u_xpb_out[25][380],u_xpb_out[26][380],u_xpb_out[27][380],u_xpb_out[28][380],u_xpb_out[29][380],u_xpb_out[30][380],u_xpb_out[31][380],u_xpb_out[32][380],u_xpb_out[33][380],u_xpb_out[34][380],u_xpb_out[35][380],u_xpb_out[36][380],u_xpb_out[37][380],u_xpb_out[38][380],u_xpb_out[39][380],u_xpb_out[40][380],u_xpb_out[41][380],u_xpb_out[42][380],u_xpb_out[43][380],u_xpb_out[44][380],u_xpb_out[45][380],u_xpb_out[46][380],u_xpb_out[47][380],u_xpb_out[48][380],u_xpb_out[49][380],u_xpb_out[50][380],u_xpb_out[51][380],u_xpb_out[52][380],u_xpb_out[53][380],u_xpb_out[54][380],u_xpb_out[55][380],u_xpb_out[56][380],u_xpb_out[57][380],u_xpb_out[58][380],u_xpb_out[59][380],u_xpb_out[60][380],u_xpb_out[61][380],u_xpb_out[62][380],u_xpb_out[63][380],u_xpb_out[64][380],u_xpb_out[65][380],u_xpb_out[66][380],u_xpb_out[67][380],u_xpb_out[68][380],u_xpb_out[69][380],u_xpb_out[70][380],u_xpb_out[71][380],u_xpb_out[72][380],u_xpb_out[73][380],u_xpb_out[74][380],u_xpb_out[75][380],u_xpb_out[76][380],u_xpb_out[77][380],u_xpb_out[78][380],u_xpb_out[79][380],u_xpb_out[80][380],u_xpb_out[81][380],u_xpb_out[82][380],u_xpb_out[83][380],u_xpb_out[84][380],u_xpb_out[85][380],u_xpb_out[86][380],u_xpb_out[87][380],u_xpb_out[88][380],u_xpb_out[89][380],u_xpb_out[90][380],u_xpb_out[91][380],u_xpb_out[92][380],u_xpb_out[93][380],u_xpb_out[94][380],u_xpb_out[95][380],u_xpb_out[96][380],u_xpb_out[97][380],u_xpb_out[98][380],u_xpb_out[99][380],u_xpb_out[100][380],u_xpb_out[101][380],u_xpb_out[102][380],u_xpb_out[103][380],u_xpb_out[104][380],u_xpb_out[105][380]};

assign col_out_381 = {u_xpb_out[0][381],u_xpb_out[1][381],u_xpb_out[2][381],u_xpb_out[3][381],u_xpb_out[4][381],u_xpb_out[5][381],u_xpb_out[6][381],u_xpb_out[7][381],u_xpb_out[8][381],u_xpb_out[9][381],u_xpb_out[10][381],u_xpb_out[11][381],u_xpb_out[12][381],u_xpb_out[13][381],u_xpb_out[14][381],u_xpb_out[15][381],u_xpb_out[16][381],u_xpb_out[17][381],u_xpb_out[18][381],u_xpb_out[19][381],u_xpb_out[20][381],u_xpb_out[21][381],u_xpb_out[22][381],u_xpb_out[23][381],u_xpb_out[24][381],u_xpb_out[25][381],u_xpb_out[26][381],u_xpb_out[27][381],u_xpb_out[28][381],u_xpb_out[29][381],u_xpb_out[30][381],u_xpb_out[31][381],u_xpb_out[32][381],u_xpb_out[33][381],u_xpb_out[34][381],u_xpb_out[35][381],u_xpb_out[36][381],u_xpb_out[37][381],u_xpb_out[38][381],u_xpb_out[39][381],u_xpb_out[40][381],u_xpb_out[41][381],u_xpb_out[42][381],u_xpb_out[43][381],u_xpb_out[44][381],u_xpb_out[45][381],u_xpb_out[46][381],u_xpb_out[47][381],u_xpb_out[48][381],u_xpb_out[49][381],u_xpb_out[50][381],u_xpb_out[51][381],u_xpb_out[52][381],u_xpb_out[53][381],u_xpb_out[54][381],u_xpb_out[55][381],u_xpb_out[56][381],u_xpb_out[57][381],u_xpb_out[58][381],u_xpb_out[59][381],u_xpb_out[60][381],u_xpb_out[61][381],u_xpb_out[62][381],u_xpb_out[63][381],u_xpb_out[64][381],u_xpb_out[65][381],u_xpb_out[66][381],u_xpb_out[67][381],u_xpb_out[68][381],u_xpb_out[69][381],u_xpb_out[70][381],u_xpb_out[71][381],u_xpb_out[72][381],u_xpb_out[73][381],u_xpb_out[74][381],u_xpb_out[75][381],u_xpb_out[76][381],u_xpb_out[77][381],u_xpb_out[78][381],u_xpb_out[79][381],u_xpb_out[80][381],u_xpb_out[81][381],u_xpb_out[82][381],u_xpb_out[83][381],u_xpb_out[84][381],u_xpb_out[85][381],u_xpb_out[86][381],u_xpb_out[87][381],u_xpb_out[88][381],u_xpb_out[89][381],u_xpb_out[90][381],u_xpb_out[91][381],u_xpb_out[92][381],u_xpb_out[93][381],u_xpb_out[94][381],u_xpb_out[95][381],u_xpb_out[96][381],u_xpb_out[97][381],u_xpb_out[98][381],u_xpb_out[99][381],u_xpb_out[100][381],u_xpb_out[101][381],u_xpb_out[102][381],u_xpb_out[103][381],u_xpb_out[104][381],u_xpb_out[105][381]};

assign col_out_382 = {u_xpb_out[0][382],u_xpb_out[1][382],u_xpb_out[2][382],u_xpb_out[3][382],u_xpb_out[4][382],u_xpb_out[5][382],u_xpb_out[6][382],u_xpb_out[7][382],u_xpb_out[8][382],u_xpb_out[9][382],u_xpb_out[10][382],u_xpb_out[11][382],u_xpb_out[12][382],u_xpb_out[13][382],u_xpb_out[14][382],u_xpb_out[15][382],u_xpb_out[16][382],u_xpb_out[17][382],u_xpb_out[18][382],u_xpb_out[19][382],u_xpb_out[20][382],u_xpb_out[21][382],u_xpb_out[22][382],u_xpb_out[23][382],u_xpb_out[24][382],u_xpb_out[25][382],u_xpb_out[26][382],u_xpb_out[27][382],u_xpb_out[28][382],u_xpb_out[29][382],u_xpb_out[30][382],u_xpb_out[31][382],u_xpb_out[32][382],u_xpb_out[33][382],u_xpb_out[34][382],u_xpb_out[35][382],u_xpb_out[36][382],u_xpb_out[37][382],u_xpb_out[38][382],u_xpb_out[39][382],u_xpb_out[40][382],u_xpb_out[41][382],u_xpb_out[42][382],u_xpb_out[43][382],u_xpb_out[44][382],u_xpb_out[45][382],u_xpb_out[46][382],u_xpb_out[47][382],u_xpb_out[48][382],u_xpb_out[49][382],u_xpb_out[50][382],u_xpb_out[51][382],u_xpb_out[52][382],u_xpb_out[53][382],u_xpb_out[54][382],u_xpb_out[55][382],u_xpb_out[56][382],u_xpb_out[57][382],u_xpb_out[58][382],u_xpb_out[59][382],u_xpb_out[60][382],u_xpb_out[61][382],u_xpb_out[62][382],u_xpb_out[63][382],u_xpb_out[64][382],u_xpb_out[65][382],u_xpb_out[66][382],u_xpb_out[67][382],u_xpb_out[68][382],u_xpb_out[69][382],u_xpb_out[70][382],u_xpb_out[71][382],u_xpb_out[72][382],u_xpb_out[73][382],u_xpb_out[74][382],u_xpb_out[75][382],u_xpb_out[76][382],u_xpb_out[77][382],u_xpb_out[78][382],u_xpb_out[79][382],u_xpb_out[80][382],u_xpb_out[81][382],u_xpb_out[82][382],u_xpb_out[83][382],u_xpb_out[84][382],u_xpb_out[85][382],u_xpb_out[86][382],u_xpb_out[87][382],u_xpb_out[88][382],u_xpb_out[89][382],u_xpb_out[90][382],u_xpb_out[91][382],u_xpb_out[92][382],u_xpb_out[93][382],u_xpb_out[94][382],u_xpb_out[95][382],u_xpb_out[96][382],u_xpb_out[97][382],u_xpb_out[98][382],u_xpb_out[99][382],u_xpb_out[100][382],u_xpb_out[101][382],u_xpb_out[102][382],u_xpb_out[103][382],u_xpb_out[104][382],u_xpb_out[105][382]};

assign col_out_383 = {u_xpb_out[0][383],u_xpb_out[1][383],u_xpb_out[2][383],u_xpb_out[3][383],u_xpb_out[4][383],u_xpb_out[5][383],u_xpb_out[6][383],u_xpb_out[7][383],u_xpb_out[8][383],u_xpb_out[9][383],u_xpb_out[10][383],u_xpb_out[11][383],u_xpb_out[12][383],u_xpb_out[13][383],u_xpb_out[14][383],u_xpb_out[15][383],u_xpb_out[16][383],u_xpb_out[17][383],u_xpb_out[18][383],u_xpb_out[19][383],u_xpb_out[20][383],u_xpb_out[21][383],u_xpb_out[22][383],u_xpb_out[23][383],u_xpb_out[24][383],u_xpb_out[25][383],u_xpb_out[26][383],u_xpb_out[27][383],u_xpb_out[28][383],u_xpb_out[29][383],u_xpb_out[30][383],u_xpb_out[31][383],u_xpb_out[32][383],u_xpb_out[33][383],u_xpb_out[34][383],u_xpb_out[35][383],u_xpb_out[36][383],u_xpb_out[37][383],u_xpb_out[38][383],u_xpb_out[39][383],u_xpb_out[40][383],u_xpb_out[41][383],u_xpb_out[42][383],u_xpb_out[43][383],u_xpb_out[44][383],u_xpb_out[45][383],u_xpb_out[46][383],u_xpb_out[47][383],u_xpb_out[48][383],u_xpb_out[49][383],u_xpb_out[50][383],u_xpb_out[51][383],u_xpb_out[52][383],u_xpb_out[53][383],u_xpb_out[54][383],u_xpb_out[55][383],u_xpb_out[56][383],u_xpb_out[57][383],u_xpb_out[58][383],u_xpb_out[59][383],u_xpb_out[60][383],u_xpb_out[61][383],u_xpb_out[62][383],u_xpb_out[63][383],u_xpb_out[64][383],u_xpb_out[65][383],u_xpb_out[66][383],u_xpb_out[67][383],u_xpb_out[68][383],u_xpb_out[69][383],u_xpb_out[70][383],u_xpb_out[71][383],u_xpb_out[72][383],u_xpb_out[73][383],u_xpb_out[74][383],u_xpb_out[75][383],u_xpb_out[76][383],u_xpb_out[77][383],u_xpb_out[78][383],u_xpb_out[79][383],u_xpb_out[80][383],u_xpb_out[81][383],u_xpb_out[82][383],u_xpb_out[83][383],u_xpb_out[84][383],u_xpb_out[85][383],u_xpb_out[86][383],u_xpb_out[87][383],u_xpb_out[88][383],u_xpb_out[89][383],u_xpb_out[90][383],u_xpb_out[91][383],u_xpb_out[92][383],u_xpb_out[93][383],u_xpb_out[94][383],u_xpb_out[95][383],u_xpb_out[96][383],u_xpb_out[97][383],u_xpb_out[98][383],u_xpb_out[99][383],u_xpb_out[100][383],u_xpb_out[101][383],u_xpb_out[102][383],u_xpb_out[103][383],u_xpb_out[104][383],u_xpb_out[105][383]};

assign col_out_384 = {u_xpb_out[0][384],u_xpb_out[1][384],u_xpb_out[2][384],u_xpb_out[3][384],u_xpb_out[4][384],u_xpb_out[5][384],u_xpb_out[6][384],u_xpb_out[7][384],u_xpb_out[8][384],u_xpb_out[9][384],u_xpb_out[10][384],u_xpb_out[11][384],u_xpb_out[12][384],u_xpb_out[13][384],u_xpb_out[14][384],u_xpb_out[15][384],u_xpb_out[16][384],u_xpb_out[17][384],u_xpb_out[18][384],u_xpb_out[19][384],u_xpb_out[20][384],u_xpb_out[21][384],u_xpb_out[22][384],u_xpb_out[23][384],u_xpb_out[24][384],u_xpb_out[25][384],u_xpb_out[26][384],u_xpb_out[27][384],u_xpb_out[28][384],u_xpb_out[29][384],u_xpb_out[30][384],u_xpb_out[31][384],u_xpb_out[32][384],u_xpb_out[33][384],u_xpb_out[34][384],u_xpb_out[35][384],u_xpb_out[36][384],u_xpb_out[37][384],u_xpb_out[38][384],u_xpb_out[39][384],u_xpb_out[40][384],u_xpb_out[41][384],u_xpb_out[42][384],u_xpb_out[43][384],u_xpb_out[44][384],u_xpb_out[45][384],u_xpb_out[46][384],u_xpb_out[47][384],u_xpb_out[48][384],u_xpb_out[49][384],u_xpb_out[50][384],u_xpb_out[51][384],u_xpb_out[52][384],u_xpb_out[53][384],u_xpb_out[54][384],u_xpb_out[55][384],u_xpb_out[56][384],u_xpb_out[57][384],u_xpb_out[58][384],u_xpb_out[59][384],u_xpb_out[60][384],u_xpb_out[61][384],u_xpb_out[62][384],u_xpb_out[63][384],u_xpb_out[64][384],u_xpb_out[65][384],u_xpb_out[66][384],u_xpb_out[67][384],u_xpb_out[68][384],u_xpb_out[69][384],u_xpb_out[70][384],u_xpb_out[71][384],u_xpb_out[72][384],u_xpb_out[73][384],u_xpb_out[74][384],u_xpb_out[75][384],u_xpb_out[76][384],u_xpb_out[77][384],u_xpb_out[78][384],u_xpb_out[79][384],u_xpb_out[80][384],u_xpb_out[81][384],u_xpb_out[82][384],u_xpb_out[83][384],u_xpb_out[84][384],u_xpb_out[85][384],u_xpb_out[86][384],u_xpb_out[87][384],u_xpb_out[88][384],u_xpb_out[89][384],u_xpb_out[90][384],u_xpb_out[91][384],u_xpb_out[92][384],u_xpb_out[93][384],u_xpb_out[94][384],u_xpb_out[95][384],u_xpb_out[96][384],u_xpb_out[97][384],u_xpb_out[98][384],u_xpb_out[99][384],u_xpb_out[100][384],u_xpb_out[101][384],u_xpb_out[102][384],u_xpb_out[103][384],u_xpb_out[104][384],u_xpb_out[105][384]};

assign col_out_385 = {u_xpb_out[0][385],u_xpb_out[1][385],u_xpb_out[2][385],u_xpb_out[3][385],u_xpb_out[4][385],u_xpb_out[5][385],u_xpb_out[6][385],u_xpb_out[7][385],u_xpb_out[8][385],u_xpb_out[9][385],u_xpb_out[10][385],u_xpb_out[11][385],u_xpb_out[12][385],u_xpb_out[13][385],u_xpb_out[14][385],u_xpb_out[15][385],u_xpb_out[16][385],u_xpb_out[17][385],u_xpb_out[18][385],u_xpb_out[19][385],u_xpb_out[20][385],u_xpb_out[21][385],u_xpb_out[22][385],u_xpb_out[23][385],u_xpb_out[24][385],u_xpb_out[25][385],u_xpb_out[26][385],u_xpb_out[27][385],u_xpb_out[28][385],u_xpb_out[29][385],u_xpb_out[30][385],u_xpb_out[31][385],u_xpb_out[32][385],u_xpb_out[33][385],u_xpb_out[34][385],u_xpb_out[35][385],u_xpb_out[36][385],u_xpb_out[37][385],u_xpb_out[38][385],u_xpb_out[39][385],u_xpb_out[40][385],u_xpb_out[41][385],u_xpb_out[42][385],u_xpb_out[43][385],u_xpb_out[44][385],u_xpb_out[45][385],u_xpb_out[46][385],u_xpb_out[47][385],u_xpb_out[48][385],u_xpb_out[49][385],u_xpb_out[50][385],u_xpb_out[51][385],u_xpb_out[52][385],u_xpb_out[53][385],u_xpb_out[54][385],u_xpb_out[55][385],u_xpb_out[56][385],u_xpb_out[57][385],u_xpb_out[58][385],u_xpb_out[59][385],u_xpb_out[60][385],u_xpb_out[61][385],u_xpb_out[62][385],u_xpb_out[63][385],u_xpb_out[64][385],u_xpb_out[65][385],u_xpb_out[66][385],u_xpb_out[67][385],u_xpb_out[68][385],u_xpb_out[69][385],u_xpb_out[70][385],u_xpb_out[71][385],u_xpb_out[72][385],u_xpb_out[73][385],u_xpb_out[74][385],u_xpb_out[75][385],u_xpb_out[76][385],u_xpb_out[77][385],u_xpb_out[78][385],u_xpb_out[79][385],u_xpb_out[80][385],u_xpb_out[81][385],u_xpb_out[82][385],u_xpb_out[83][385],u_xpb_out[84][385],u_xpb_out[85][385],u_xpb_out[86][385],u_xpb_out[87][385],u_xpb_out[88][385],u_xpb_out[89][385],u_xpb_out[90][385],u_xpb_out[91][385],u_xpb_out[92][385],u_xpb_out[93][385],u_xpb_out[94][385],u_xpb_out[95][385],u_xpb_out[96][385],u_xpb_out[97][385],u_xpb_out[98][385],u_xpb_out[99][385],u_xpb_out[100][385],u_xpb_out[101][385],u_xpb_out[102][385],u_xpb_out[103][385],u_xpb_out[104][385],u_xpb_out[105][385]};

assign col_out_386 = {u_xpb_out[0][386],u_xpb_out[1][386],u_xpb_out[2][386],u_xpb_out[3][386],u_xpb_out[4][386],u_xpb_out[5][386],u_xpb_out[6][386],u_xpb_out[7][386],u_xpb_out[8][386],u_xpb_out[9][386],u_xpb_out[10][386],u_xpb_out[11][386],u_xpb_out[12][386],u_xpb_out[13][386],u_xpb_out[14][386],u_xpb_out[15][386],u_xpb_out[16][386],u_xpb_out[17][386],u_xpb_out[18][386],u_xpb_out[19][386],u_xpb_out[20][386],u_xpb_out[21][386],u_xpb_out[22][386],u_xpb_out[23][386],u_xpb_out[24][386],u_xpb_out[25][386],u_xpb_out[26][386],u_xpb_out[27][386],u_xpb_out[28][386],u_xpb_out[29][386],u_xpb_out[30][386],u_xpb_out[31][386],u_xpb_out[32][386],u_xpb_out[33][386],u_xpb_out[34][386],u_xpb_out[35][386],u_xpb_out[36][386],u_xpb_out[37][386],u_xpb_out[38][386],u_xpb_out[39][386],u_xpb_out[40][386],u_xpb_out[41][386],u_xpb_out[42][386],u_xpb_out[43][386],u_xpb_out[44][386],u_xpb_out[45][386],u_xpb_out[46][386],u_xpb_out[47][386],u_xpb_out[48][386],u_xpb_out[49][386],u_xpb_out[50][386],u_xpb_out[51][386],u_xpb_out[52][386],u_xpb_out[53][386],u_xpb_out[54][386],u_xpb_out[55][386],u_xpb_out[56][386],u_xpb_out[57][386],u_xpb_out[58][386],u_xpb_out[59][386],u_xpb_out[60][386],u_xpb_out[61][386],u_xpb_out[62][386],u_xpb_out[63][386],u_xpb_out[64][386],u_xpb_out[65][386],u_xpb_out[66][386],u_xpb_out[67][386],u_xpb_out[68][386],u_xpb_out[69][386],u_xpb_out[70][386],u_xpb_out[71][386],u_xpb_out[72][386],u_xpb_out[73][386],u_xpb_out[74][386],u_xpb_out[75][386],u_xpb_out[76][386],u_xpb_out[77][386],u_xpb_out[78][386],u_xpb_out[79][386],u_xpb_out[80][386],u_xpb_out[81][386],u_xpb_out[82][386],u_xpb_out[83][386],u_xpb_out[84][386],u_xpb_out[85][386],u_xpb_out[86][386],u_xpb_out[87][386],u_xpb_out[88][386],u_xpb_out[89][386],u_xpb_out[90][386],u_xpb_out[91][386],u_xpb_out[92][386],u_xpb_out[93][386],u_xpb_out[94][386],u_xpb_out[95][386],u_xpb_out[96][386],u_xpb_out[97][386],u_xpb_out[98][386],u_xpb_out[99][386],u_xpb_out[100][386],u_xpb_out[101][386],u_xpb_out[102][386],u_xpb_out[103][386],u_xpb_out[104][386],u_xpb_out[105][386]};

assign col_out_387 = {u_xpb_out[0][387],u_xpb_out[1][387],u_xpb_out[2][387],u_xpb_out[3][387],u_xpb_out[4][387],u_xpb_out[5][387],u_xpb_out[6][387],u_xpb_out[7][387],u_xpb_out[8][387],u_xpb_out[9][387],u_xpb_out[10][387],u_xpb_out[11][387],u_xpb_out[12][387],u_xpb_out[13][387],u_xpb_out[14][387],u_xpb_out[15][387],u_xpb_out[16][387],u_xpb_out[17][387],u_xpb_out[18][387],u_xpb_out[19][387],u_xpb_out[20][387],u_xpb_out[21][387],u_xpb_out[22][387],u_xpb_out[23][387],u_xpb_out[24][387],u_xpb_out[25][387],u_xpb_out[26][387],u_xpb_out[27][387],u_xpb_out[28][387],u_xpb_out[29][387],u_xpb_out[30][387],u_xpb_out[31][387],u_xpb_out[32][387],u_xpb_out[33][387],u_xpb_out[34][387],u_xpb_out[35][387],u_xpb_out[36][387],u_xpb_out[37][387],u_xpb_out[38][387],u_xpb_out[39][387],u_xpb_out[40][387],u_xpb_out[41][387],u_xpb_out[42][387],u_xpb_out[43][387],u_xpb_out[44][387],u_xpb_out[45][387],u_xpb_out[46][387],u_xpb_out[47][387],u_xpb_out[48][387],u_xpb_out[49][387],u_xpb_out[50][387],u_xpb_out[51][387],u_xpb_out[52][387],u_xpb_out[53][387],u_xpb_out[54][387],u_xpb_out[55][387],u_xpb_out[56][387],u_xpb_out[57][387],u_xpb_out[58][387],u_xpb_out[59][387],u_xpb_out[60][387],u_xpb_out[61][387],u_xpb_out[62][387],u_xpb_out[63][387],u_xpb_out[64][387],u_xpb_out[65][387],u_xpb_out[66][387],u_xpb_out[67][387],u_xpb_out[68][387],u_xpb_out[69][387],u_xpb_out[70][387],u_xpb_out[71][387],u_xpb_out[72][387],u_xpb_out[73][387],u_xpb_out[74][387],u_xpb_out[75][387],u_xpb_out[76][387],u_xpb_out[77][387],u_xpb_out[78][387],u_xpb_out[79][387],u_xpb_out[80][387],u_xpb_out[81][387],u_xpb_out[82][387],u_xpb_out[83][387],u_xpb_out[84][387],u_xpb_out[85][387],u_xpb_out[86][387],u_xpb_out[87][387],u_xpb_out[88][387],u_xpb_out[89][387],u_xpb_out[90][387],u_xpb_out[91][387],u_xpb_out[92][387],u_xpb_out[93][387],u_xpb_out[94][387],u_xpb_out[95][387],u_xpb_out[96][387],u_xpb_out[97][387],u_xpb_out[98][387],u_xpb_out[99][387],u_xpb_out[100][387],u_xpb_out[101][387],u_xpb_out[102][387],u_xpb_out[103][387],u_xpb_out[104][387],u_xpb_out[105][387]};

assign col_out_388 = {u_xpb_out[0][388],u_xpb_out[1][388],u_xpb_out[2][388],u_xpb_out[3][388],u_xpb_out[4][388],u_xpb_out[5][388],u_xpb_out[6][388],u_xpb_out[7][388],u_xpb_out[8][388],u_xpb_out[9][388],u_xpb_out[10][388],u_xpb_out[11][388],u_xpb_out[12][388],u_xpb_out[13][388],u_xpb_out[14][388],u_xpb_out[15][388],u_xpb_out[16][388],u_xpb_out[17][388],u_xpb_out[18][388],u_xpb_out[19][388],u_xpb_out[20][388],u_xpb_out[21][388],u_xpb_out[22][388],u_xpb_out[23][388],u_xpb_out[24][388],u_xpb_out[25][388],u_xpb_out[26][388],u_xpb_out[27][388],u_xpb_out[28][388],u_xpb_out[29][388],u_xpb_out[30][388],u_xpb_out[31][388],u_xpb_out[32][388],u_xpb_out[33][388],u_xpb_out[34][388],u_xpb_out[35][388],u_xpb_out[36][388],u_xpb_out[37][388],u_xpb_out[38][388],u_xpb_out[39][388],u_xpb_out[40][388],u_xpb_out[41][388],u_xpb_out[42][388],u_xpb_out[43][388],u_xpb_out[44][388],u_xpb_out[45][388],u_xpb_out[46][388],u_xpb_out[47][388],u_xpb_out[48][388],u_xpb_out[49][388],u_xpb_out[50][388],u_xpb_out[51][388],u_xpb_out[52][388],u_xpb_out[53][388],u_xpb_out[54][388],u_xpb_out[55][388],u_xpb_out[56][388],u_xpb_out[57][388],u_xpb_out[58][388],u_xpb_out[59][388],u_xpb_out[60][388],u_xpb_out[61][388],u_xpb_out[62][388],u_xpb_out[63][388],u_xpb_out[64][388],u_xpb_out[65][388],u_xpb_out[66][388],u_xpb_out[67][388],u_xpb_out[68][388],u_xpb_out[69][388],u_xpb_out[70][388],u_xpb_out[71][388],u_xpb_out[72][388],u_xpb_out[73][388],u_xpb_out[74][388],u_xpb_out[75][388],u_xpb_out[76][388],u_xpb_out[77][388],u_xpb_out[78][388],u_xpb_out[79][388],u_xpb_out[80][388],u_xpb_out[81][388],u_xpb_out[82][388],u_xpb_out[83][388],u_xpb_out[84][388],u_xpb_out[85][388],u_xpb_out[86][388],u_xpb_out[87][388],u_xpb_out[88][388],u_xpb_out[89][388],u_xpb_out[90][388],u_xpb_out[91][388],u_xpb_out[92][388],u_xpb_out[93][388],u_xpb_out[94][388],u_xpb_out[95][388],u_xpb_out[96][388],u_xpb_out[97][388],u_xpb_out[98][388],u_xpb_out[99][388],u_xpb_out[100][388],u_xpb_out[101][388],u_xpb_out[102][388],u_xpb_out[103][388],u_xpb_out[104][388],u_xpb_out[105][388]};

assign col_out_389 = {u_xpb_out[0][389],u_xpb_out[1][389],u_xpb_out[2][389],u_xpb_out[3][389],u_xpb_out[4][389],u_xpb_out[5][389],u_xpb_out[6][389],u_xpb_out[7][389],u_xpb_out[8][389],u_xpb_out[9][389],u_xpb_out[10][389],u_xpb_out[11][389],u_xpb_out[12][389],u_xpb_out[13][389],u_xpb_out[14][389],u_xpb_out[15][389],u_xpb_out[16][389],u_xpb_out[17][389],u_xpb_out[18][389],u_xpb_out[19][389],u_xpb_out[20][389],u_xpb_out[21][389],u_xpb_out[22][389],u_xpb_out[23][389],u_xpb_out[24][389],u_xpb_out[25][389],u_xpb_out[26][389],u_xpb_out[27][389],u_xpb_out[28][389],u_xpb_out[29][389],u_xpb_out[30][389],u_xpb_out[31][389],u_xpb_out[32][389],u_xpb_out[33][389],u_xpb_out[34][389],u_xpb_out[35][389],u_xpb_out[36][389],u_xpb_out[37][389],u_xpb_out[38][389],u_xpb_out[39][389],u_xpb_out[40][389],u_xpb_out[41][389],u_xpb_out[42][389],u_xpb_out[43][389],u_xpb_out[44][389],u_xpb_out[45][389],u_xpb_out[46][389],u_xpb_out[47][389],u_xpb_out[48][389],u_xpb_out[49][389],u_xpb_out[50][389],u_xpb_out[51][389],u_xpb_out[52][389],u_xpb_out[53][389],u_xpb_out[54][389],u_xpb_out[55][389],u_xpb_out[56][389],u_xpb_out[57][389],u_xpb_out[58][389],u_xpb_out[59][389],u_xpb_out[60][389],u_xpb_out[61][389],u_xpb_out[62][389],u_xpb_out[63][389],u_xpb_out[64][389],u_xpb_out[65][389],u_xpb_out[66][389],u_xpb_out[67][389],u_xpb_out[68][389],u_xpb_out[69][389],u_xpb_out[70][389],u_xpb_out[71][389],u_xpb_out[72][389],u_xpb_out[73][389],u_xpb_out[74][389],u_xpb_out[75][389],u_xpb_out[76][389],u_xpb_out[77][389],u_xpb_out[78][389],u_xpb_out[79][389],u_xpb_out[80][389],u_xpb_out[81][389],u_xpb_out[82][389],u_xpb_out[83][389],u_xpb_out[84][389],u_xpb_out[85][389],u_xpb_out[86][389],u_xpb_out[87][389],u_xpb_out[88][389],u_xpb_out[89][389],u_xpb_out[90][389],u_xpb_out[91][389],u_xpb_out[92][389],u_xpb_out[93][389],u_xpb_out[94][389],u_xpb_out[95][389],u_xpb_out[96][389],u_xpb_out[97][389],u_xpb_out[98][389],u_xpb_out[99][389],u_xpb_out[100][389],u_xpb_out[101][389],u_xpb_out[102][389],u_xpb_out[103][389],u_xpb_out[104][389],u_xpb_out[105][389]};

assign col_out_390 = {u_xpb_out[0][390],u_xpb_out[1][390],u_xpb_out[2][390],u_xpb_out[3][390],u_xpb_out[4][390],u_xpb_out[5][390],u_xpb_out[6][390],u_xpb_out[7][390],u_xpb_out[8][390],u_xpb_out[9][390],u_xpb_out[10][390],u_xpb_out[11][390],u_xpb_out[12][390],u_xpb_out[13][390],u_xpb_out[14][390],u_xpb_out[15][390],u_xpb_out[16][390],u_xpb_out[17][390],u_xpb_out[18][390],u_xpb_out[19][390],u_xpb_out[20][390],u_xpb_out[21][390],u_xpb_out[22][390],u_xpb_out[23][390],u_xpb_out[24][390],u_xpb_out[25][390],u_xpb_out[26][390],u_xpb_out[27][390],u_xpb_out[28][390],u_xpb_out[29][390],u_xpb_out[30][390],u_xpb_out[31][390],u_xpb_out[32][390],u_xpb_out[33][390],u_xpb_out[34][390],u_xpb_out[35][390],u_xpb_out[36][390],u_xpb_out[37][390],u_xpb_out[38][390],u_xpb_out[39][390],u_xpb_out[40][390],u_xpb_out[41][390],u_xpb_out[42][390],u_xpb_out[43][390],u_xpb_out[44][390],u_xpb_out[45][390],u_xpb_out[46][390],u_xpb_out[47][390],u_xpb_out[48][390],u_xpb_out[49][390],u_xpb_out[50][390],u_xpb_out[51][390],u_xpb_out[52][390],u_xpb_out[53][390],u_xpb_out[54][390],u_xpb_out[55][390],u_xpb_out[56][390],u_xpb_out[57][390],u_xpb_out[58][390],u_xpb_out[59][390],u_xpb_out[60][390],u_xpb_out[61][390],u_xpb_out[62][390],u_xpb_out[63][390],u_xpb_out[64][390],u_xpb_out[65][390],u_xpb_out[66][390],u_xpb_out[67][390],u_xpb_out[68][390],u_xpb_out[69][390],u_xpb_out[70][390],u_xpb_out[71][390],u_xpb_out[72][390],u_xpb_out[73][390],u_xpb_out[74][390],u_xpb_out[75][390],u_xpb_out[76][390],u_xpb_out[77][390],u_xpb_out[78][390],u_xpb_out[79][390],u_xpb_out[80][390],u_xpb_out[81][390],u_xpb_out[82][390],u_xpb_out[83][390],u_xpb_out[84][390],u_xpb_out[85][390],u_xpb_out[86][390],u_xpb_out[87][390],u_xpb_out[88][390],u_xpb_out[89][390],u_xpb_out[90][390],u_xpb_out[91][390],u_xpb_out[92][390],u_xpb_out[93][390],u_xpb_out[94][390],u_xpb_out[95][390],u_xpb_out[96][390],u_xpb_out[97][390],u_xpb_out[98][390],u_xpb_out[99][390],u_xpb_out[100][390],u_xpb_out[101][390],u_xpb_out[102][390],u_xpb_out[103][390],u_xpb_out[104][390],u_xpb_out[105][390]};

assign col_out_391 = {u_xpb_out[0][391],u_xpb_out[1][391],u_xpb_out[2][391],u_xpb_out[3][391],u_xpb_out[4][391],u_xpb_out[5][391],u_xpb_out[6][391],u_xpb_out[7][391],u_xpb_out[8][391],u_xpb_out[9][391],u_xpb_out[10][391],u_xpb_out[11][391],u_xpb_out[12][391],u_xpb_out[13][391],u_xpb_out[14][391],u_xpb_out[15][391],u_xpb_out[16][391],u_xpb_out[17][391],u_xpb_out[18][391],u_xpb_out[19][391],u_xpb_out[20][391],u_xpb_out[21][391],u_xpb_out[22][391],u_xpb_out[23][391],u_xpb_out[24][391],u_xpb_out[25][391],u_xpb_out[26][391],u_xpb_out[27][391],u_xpb_out[28][391],u_xpb_out[29][391],u_xpb_out[30][391],u_xpb_out[31][391],u_xpb_out[32][391],u_xpb_out[33][391],u_xpb_out[34][391],u_xpb_out[35][391],u_xpb_out[36][391],u_xpb_out[37][391],u_xpb_out[38][391],u_xpb_out[39][391],u_xpb_out[40][391],u_xpb_out[41][391],u_xpb_out[42][391],u_xpb_out[43][391],u_xpb_out[44][391],u_xpb_out[45][391],u_xpb_out[46][391],u_xpb_out[47][391],u_xpb_out[48][391],u_xpb_out[49][391],u_xpb_out[50][391],u_xpb_out[51][391],u_xpb_out[52][391],u_xpb_out[53][391],u_xpb_out[54][391],u_xpb_out[55][391],u_xpb_out[56][391],u_xpb_out[57][391],u_xpb_out[58][391],u_xpb_out[59][391],u_xpb_out[60][391],u_xpb_out[61][391],u_xpb_out[62][391],u_xpb_out[63][391],u_xpb_out[64][391],u_xpb_out[65][391],u_xpb_out[66][391],u_xpb_out[67][391],u_xpb_out[68][391],u_xpb_out[69][391],u_xpb_out[70][391],u_xpb_out[71][391],u_xpb_out[72][391],u_xpb_out[73][391],u_xpb_out[74][391],u_xpb_out[75][391],u_xpb_out[76][391],u_xpb_out[77][391],u_xpb_out[78][391],u_xpb_out[79][391],u_xpb_out[80][391],u_xpb_out[81][391],u_xpb_out[82][391],u_xpb_out[83][391],u_xpb_out[84][391],u_xpb_out[85][391],u_xpb_out[86][391],u_xpb_out[87][391],u_xpb_out[88][391],u_xpb_out[89][391],u_xpb_out[90][391],u_xpb_out[91][391],u_xpb_out[92][391],u_xpb_out[93][391],u_xpb_out[94][391],u_xpb_out[95][391],u_xpb_out[96][391],u_xpb_out[97][391],u_xpb_out[98][391],u_xpb_out[99][391],u_xpb_out[100][391],u_xpb_out[101][391],u_xpb_out[102][391],u_xpb_out[103][391],u_xpb_out[104][391],u_xpb_out[105][391]};

assign col_out_392 = {u_xpb_out[0][392],u_xpb_out[1][392],u_xpb_out[2][392],u_xpb_out[3][392],u_xpb_out[4][392],u_xpb_out[5][392],u_xpb_out[6][392],u_xpb_out[7][392],u_xpb_out[8][392],u_xpb_out[9][392],u_xpb_out[10][392],u_xpb_out[11][392],u_xpb_out[12][392],u_xpb_out[13][392],u_xpb_out[14][392],u_xpb_out[15][392],u_xpb_out[16][392],u_xpb_out[17][392],u_xpb_out[18][392],u_xpb_out[19][392],u_xpb_out[20][392],u_xpb_out[21][392],u_xpb_out[22][392],u_xpb_out[23][392],u_xpb_out[24][392],u_xpb_out[25][392],u_xpb_out[26][392],u_xpb_out[27][392],u_xpb_out[28][392],u_xpb_out[29][392],u_xpb_out[30][392],u_xpb_out[31][392],u_xpb_out[32][392],u_xpb_out[33][392],u_xpb_out[34][392],u_xpb_out[35][392],u_xpb_out[36][392],u_xpb_out[37][392],u_xpb_out[38][392],u_xpb_out[39][392],u_xpb_out[40][392],u_xpb_out[41][392],u_xpb_out[42][392],u_xpb_out[43][392],u_xpb_out[44][392],u_xpb_out[45][392],u_xpb_out[46][392],u_xpb_out[47][392],u_xpb_out[48][392],u_xpb_out[49][392],u_xpb_out[50][392],u_xpb_out[51][392],u_xpb_out[52][392],u_xpb_out[53][392],u_xpb_out[54][392],u_xpb_out[55][392],u_xpb_out[56][392],u_xpb_out[57][392],u_xpb_out[58][392],u_xpb_out[59][392],u_xpb_out[60][392],u_xpb_out[61][392],u_xpb_out[62][392],u_xpb_out[63][392],u_xpb_out[64][392],u_xpb_out[65][392],u_xpb_out[66][392],u_xpb_out[67][392],u_xpb_out[68][392],u_xpb_out[69][392],u_xpb_out[70][392],u_xpb_out[71][392],u_xpb_out[72][392],u_xpb_out[73][392],u_xpb_out[74][392],u_xpb_out[75][392],u_xpb_out[76][392],u_xpb_out[77][392],u_xpb_out[78][392],u_xpb_out[79][392],u_xpb_out[80][392],u_xpb_out[81][392],u_xpb_out[82][392],u_xpb_out[83][392],u_xpb_out[84][392],u_xpb_out[85][392],u_xpb_out[86][392],u_xpb_out[87][392],u_xpb_out[88][392],u_xpb_out[89][392],u_xpb_out[90][392],u_xpb_out[91][392],u_xpb_out[92][392],u_xpb_out[93][392],u_xpb_out[94][392],u_xpb_out[95][392],u_xpb_out[96][392],u_xpb_out[97][392],u_xpb_out[98][392],u_xpb_out[99][392],u_xpb_out[100][392],u_xpb_out[101][392],u_xpb_out[102][392],u_xpb_out[103][392],u_xpb_out[104][392],u_xpb_out[105][392]};

assign col_out_393 = {u_xpb_out[0][393],u_xpb_out[1][393],u_xpb_out[2][393],u_xpb_out[3][393],u_xpb_out[4][393],u_xpb_out[5][393],u_xpb_out[6][393],u_xpb_out[7][393],u_xpb_out[8][393],u_xpb_out[9][393],u_xpb_out[10][393],u_xpb_out[11][393],u_xpb_out[12][393],u_xpb_out[13][393],u_xpb_out[14][393],u_xpb_out[15][393],u_xpb_out[16][393],u_xpb_out[17][393],u_xpb_out[18][393],u_xpb_out[19][393],u_xpb_out[20][393],u_xpb_out[21][393],u_xpb_out[22][393],u_xpb_out[23][393],u_xpb_out[24][393],u_xpb_out[25][393],u_xpb_out[26][393],u_xpb_out[27][393],u_xpb_out[28][393],u_xpb_out[29][393],u_xpb_out[30][393],u_xpb_out[31][393],u_xpb_out[32][393],u_xpb_out[33][393],u_xpb_out[34][393],u_xpb_out[35][393],u_xpb_out[36][393],u_xpb_out[37][393],u_xpb_out[38][393],u_xpb_out[39][393],u_xpb_out[40][393],u_xpb_out[41][393],u_xpb_out[42][393],u_xpb_out[43][393],u_xpb_out[44][393],u_xpb_out[45][393],u_xpb_out[46][393],u_xpb_out[47][393],u_xpb_out[48][393],u_xpb_out[49][393],u_xpb_out[50][393],u_xpb_out[51][393],u_xpb_out[52][393],u_xpb_out[53][393],u_xpb_out[54][393],u_xpb_out[55][393],u_xpb_out[56][393],u_xpb_out[57][393],u_xpb_out[58][393],u_xpb_out[59][393],u_xpb_out[60][393],u_xpb_out[61][393],u_xpb_out[62][393],u_xpb_out[63][393],u_xpb_out[64][393],u_xpb_out[65][393],u_xpb_out[66][393],u_xpb_out[67][393],u_xpb_out[68][393],u_xpb_out[69][393],u_xpb_out[70][393],u_xpb_out[71][393],u_xpb_out[72][393],u_xpb_out[73][393],u_xpb_out[74][393],u_xpb_out[75][393],u_xpb_out[76][393],u_xpb_out[77][393],u_xpb_out[78][393],u_xpb_out[79][393],u_xpb_out[80][393],u_xpb_out[81][393],u_xpb_out[82][393],u_xpb_out[83][393],u_xpb_out[84][393],u_xpb_out[85][393],u_xpb_out[86][393],u_xpb_out[87][393],u_xpb_out[88][393],u_xpb_out[89][393],u_xpb_out[90][393],u_xpb_out[91][393],u_xpb_out[92][393],u_xpb_out[93][393],u_xpb_out[94][393],u_xpb_out[95][393],u_xpb_out[96][393],u_xpb_out[97][393],u_xpb_out[98][393],u_xpb_out[99][393],u_xpb_out[100][393],u_xpb_out[101][393],u_xpb_out[102][393],u_xpb_out[103][393],u_xpb_out[104][393],u_xpb_out[105][393]};

assign col_out_394 = {u_xpb_out[0][394],u_xpb_out[1][394],u_xpb_out[2][394],u_xpb_out[3][394],u_xpb_out[4][394],u_xpb_out[5][394],u_xpb_out[6][394],u_xpb_out[7][394],u_xpb_out[8][394],u_xpb_out[9][394],u_xpb_out[10][394],u_xpb_out[11][394],u_xpb_out[12][394],u_xpb_out[13][394],u_xpb_out[14][394],u_xpb_out[15][394],u_xpb_out[16][394],u_xpb_out[17][394],u_xpb_out[18][394],u_xpb_out[19][394],u_xpb_out[20][394],u_xpb_out[21][394],u_xpb_out[22][394],u_xpb_out[23][394],u_xpb_out[24][394],u_xpb_out[25][394],u_xpb_out[26][394],u_xpb_out[27][394],u_xpb_out[28][394],u_xpb_out[29][394],u_xpb_out[30][394],u_xpb_out[31][394],u_xpb_out[32][394],u_xpb_out[33][394],u_xpb_out[34][394],u_xpb_out[35][394],u_xpb_out[36][394],u_xpb_out[37][394],u_xpb_out[38][394],u_xpb_out[39][394],u_xpb_out[40][394],u_xpb_out[41][394],u_xpb_out[42][394],u_xpb_out[43][394],u_xpb_out[44][394],u_xpb_out[45][394],u_xpb_out[46][394],u_xpb_out[47][394],u_xpb_out[48][394],u_xpb_out[49][394],u_xpb_out[50][394],u_xpb_out[51][394],u_xpb_out[52][394],u_xpb_out[53][394],u_xpb_out[54][394],u_xpb_out[55][394],u_xpb_out[56][394],u_xpb_out[57][394],u_xpb_out[58][394],u_xpb_out[59][394],u_xpb_out[60][394],u_xpb_out[61][394],u_xpb_out[62][394],u_xpb_out[63][394],u_xpb_out[64][394],u_xpb_out[65][394],u_xpb_out[66][394],u_xpb_out[67][394],u_xpb_out[68][394],u_xpb_out[69][394],u_xpb_out[70][394],u_xpb_out[71][394],u_xpb_out[72][394],u_xpb_out[73][394],u_xpb_out[74][394],u_xpb_out[75][394],u_xpb_out[76][394],u_xpb_out[77][394],u_xpb_out[78][394],u_xpb_out[79][394],u_xpb_out[80][394],u_xpb_out[81][394],u_xpb_out[82][394],u_xpb_out[83][394],u_xpb_out[84][394],u_xpb_out[85][394],u_xpb_out[86][394],u_xpb_out[87][394],u_xpb_out[88][394],u_xpb_out[89][394],u_xpb_out[90][394],u_xpb_out[91][394],u_xpb_out[92][394],u_xpb_out[93][394],u_xpb_out[94][394],u_xpb_out[95][394],u_xpb_out[96][394],u_xpb_out[97][394],u_xpb_out[98][394],u_xpb_out[99][394],u_xpb_out[100][394],u_xpb_out[101][394],u_xpb_out[102][394],u_xpb_out[103][394],u_xpb_out[104][394],u_xpb_out[105][394]};

assign col_out_395 = {u_xpb_out[0][395],u_xpb_out[1][395],u_xpb_out[2][395],u_xpb_out[3][395],u_xpb_out[4][395],u_xpb_out[5][395],u_xpb_out[6][395],u_xpb_out[7][395],u_xpb_out[8][395],u_xpb_out[9][395],u_xpb_out[10][395],u_xpb_out[11][395],u_xpb_out[12][395],u_xpb_out[13][395],u_xpb_out[14][395],u_xpb_out[15][395],u_xpb_out[16][395],u_xpb_out[17][395],u_xpb_out[18][395],u_xpb_out[19][395],u_xpb_out[20][395],u_xpb_out[21][395],u_xpb_out[22][395],u_xpb_out[23][395],u_xpb_out[24][395],u_xpb_out[25][395],u_xpb_out[26][395],u_xpb_out[27][395],u_xpb_out[28][395],u_xpb_out[29][395],u_xpb_out[30][395],u_xpb_out[31][395],u_xpb_out[32][395],u_xpb_out[33][395],u_xpb_out[34][395],u_xpb_out[35][395],u_xpb_out[36][395],u_xpb_out[37][395],u_xpb_out[38][395],u_xpb_out[39][395],u_xpb_out[40][395],u_xpb_out[41][395],u_xpb_out[42][395],u_xpb_out[43][395],u_xpb_out[44][395],u_xpb_out[45][395],u_xpb_out[46][395],u_xpb_out[47][395],u_xpb_out[48][395],u_xpb_out[49][395],u_xpb_out[50][395],u_xpb_out[51][395],u_xpb_out[52][395],u_xpb_out[53][395],u_xpb_out[54][395],u_xpb_out[55][395],u_xpb_out[56][395],u_xpb_out[57][395],u_xpb_out[58][395],u_xpb_out[59][395],u_xpb_out[60][395],u_xpb_out[61][395],u_xpb_out[62][395],u_xpb_out[63][395],u_xpb_out[64][395],u_xpb_out[65][395],u_xpb_out[66][395],u_xpb_out[67][395],u_xpb_out[68][395],u_xpb_out[69][395],u_xpb_out[70][395],u_xpb_out[71][395],u_xpb_out[72][395],u_xpb_out[73][395],u_xpb_out[74][395],u_xpb_out[75][395],u_xpb_out[76][395],u_xpb_out[77][395],u_xpb_out[78][395],u_xpb_out[79][395],u_xpb_out[80][395],u_xpb_out[81][395],u_xpb_out[82][395],u_xpb_out[83][395],u_xpb_out[84][395],u_xpb_out[85][395],u_xpb_out[86][395],u_xpb_out[87][395],u_xpb_out[88][395],u_xpb_out[89][395],u_xpb_out[90][395],u_xpb_out[91][395],u_xpb_out[92][395],u_xpb_out[93][395],u_xpb_out[94][395],u_xpb_out[95][395],u_xpb_out[96][395],u_xpb_out[97][395],u_xpb_out[98][395],u_xpb_out[99][395],u_xpb_out[100][395],u_xpb_out[101][395],u_xpb_out[102][395],u_xpb_out[103][395],u_xpb_out[104][395],u_xpb_out[105][395]};

assign col_out_396 = {u_xpb_out[0][396],u_xpb_out[1][396],u_xpb_out[2][396],u_xpb_out[3][396],u_xpb_out[4][396],u_xpb_out[5][396],u_xpb_out[6][396],u_xpb_out[7][396],u_xpb_out[8][396],u_xpb_out[9][396],u_xpb_out[10][396],u_xpb_out[11][396],u_xpb_out[12][396],u_xpb_out[13][396],u_xpb_out[14][396],u_xpb_out[15][396],u_xpb_out[16][396],u_xpb_out[17][396],u_xpb_out[18][396],u_xpb_out[19][396],u_xpb_out[20][396],u_xpb_out[21][396],u_xpb_out[22][396],u_xpb_out[23][396],u_xpb_out[24][396],u_xpb_out[25][396],u_xpb_out[26][396],u_xpb_out[27][396],u_xpb_out[28][396],u_xpb_out[29][396],u_xpb_out[30][396],u_xpb_out[31][396],u_xpb_out[32][396],u_xpb_out[33][396],u_xpb_out[34][396],u_xpb_out[35][396],u_xpb_out[36][396],u_xpb_out[37][396],u_xpb_out[38][396],u_xpb_out[39][396],u_xpb_out[40][396],u_xpb_out[41][396],u_xpb_out[42][396],u_xpb_out[43][396],u_xpb_out[44][396],u_xpb_out[45][396],u_xpb_out[46][396],u_xpb_out[47][396],u_xpb_out[48][396],u_xpb_out[49][396],u_xpb_out[50][396],u_xpb_out[51][396],u_xpb_out[52][396],u_xpb_out[53][396],u_xpb_out[54][396],u_xpb_out[55][396],u_xpb_out[56][396],u_xpb_out[57][396],u_xpb_out[58][396],u_xpb_out[59][396],u_xpb_out[60][396],u_xpb_out[61][396],u_xpb_out[62][396],u_xpb_out[63][396],u_xpb_out[64][396],u_xpb_out[65][396],u_xpb_out[66][396],u_xpb_out[67][396],u_xpb_out[68][396],u_xpb_out[69][396],u_xpb_out[70][396],u_xpb_out[71][396],u_xpb_out[72][396],u_xpb_out[73][396],u_xpb_out[74][396],u_xpb_out[75][396],u_xpb_out[76][396],u_xpb_out[77][396],u_xpb_out[78][396],u_xpb_out[79][396],u_xpb_out[80][396],u_xpb_out[81][396],u_xpb_out[82][396],u_xpb_out[83][396],u_xpb_out[84][396],u_xpb_out[85][396],u_xpb_out[86][396],u_xpb_out[87][396],u_xpb_out[88][396],u_xpb_out[89][396],u_xpb_out[90][396],u_xpb_out[91][396],u_xpb_out[92][396],u_xpb_out[93][396],u_xpb_out[94][396],u_xpb_out[95][396],u_xpb_out[96][396],u_xpb_out[97][396],u_xpb_out[98][396],u_xpb_out[99][396],u_xpb_out[100][396],u_xpb_out[101][396],u_xpb_out[102][396],u_xpb_out[103][396],u_xpb_out[104][396],u_xpb_out[105][396]};

assign col_out_397 = {u_xpb_out[0][397],u_xpb_out[1][397],u_xpb_out[2][397],u_xpb_out[3][397],u_xpb_out[4][397],u_xpb_out[5][397],u_xpb_out[6][397],u_xpb_out[7][397],u_xpb_out[8][397],u_xpb_out[9][397],u_xpb_out[10][397],u_xpb_out[11][397],u_xpb_out[12][397],u_xpb_out[13][397],u_xpb_out[14][397],u_xpb_out[15][397],u_xpb_out[16][397],u_xpb_out[17][397],u_xpb_out[18][397],u_xpb_out[19][397],u_xpb_out[20][397],u_xpb_out[21][397],u_xpb_out[22][397],u_xpb_out[23][397],u_xpb_out[24][397],u_xpb_out[25][397],u_xpb_out[26][397],u_xpb_out[27][397],u_xpb_out[28][397],u_xpb_out[29][397],u_xpb_out[30][397],u_xpb_out[31][397],u_xpb_out[32][397],u_xpb_out[33][397],u_xpb_out[34][397],u_xpb_out[35][397],u_xpb_out[36][397],u_xpb_out[37][397],u_xpb_out[38][397],u_xpb_out[39][397],u_xpb_out[40][397],u_xpb_out[41][397],u_xpb_out[42][397],u_xpb_out[43][397],u_xpb_out[44][397],u_xpb_out[45][397],u_xpb_out[46][397],u_xpb_out[47][397],u_xpb_out[48][397],u_xpb_out[49][397],u_xpb_out[50][397],u_xpb_out[51][397],u_xpb_out[52][397],u_xpb_out[53][397],u_xpb_out[54][397],u_xpb_out[55][397],u_xpb_out[56][397],u_xpb_out[57][397],u_xpb_out[58][397],u_xpb_out[59][397],u_xpb_out[60][397],u_xpb_out[61][397],u_xpb_out[62][397],u_xpb_out[63][397],u_xpb_out[64][397],u_xpb_out[65][397],u_xpb_out[66][397],u_xpb_out[67][397],u_xpb_out[68][397],u_xpb_out[69][397],u_xpb_out[70][397],u_xpb_out[71][397],u_xpb_out[72][397],u_xpb_out[73][397],u_xpb_out[74][397],u_xpb_out[75][397],u_xpb_out[76][397],u_xpb_out[77][397],u_xpb_out[78][397],u_xpb_out[79][397],u_xpb_out[80][397],u_xpb_out[81][397],u_xpb_out[82][397],u_xpb_out[83][397],u_xpb_out[84][397],u_xpb_out[85][397],u_xpb_out[86][397],u_xpb_out[87][397],u_xpb_out[88][397],u_xpb_out[89][397],u_xpb_out[90][397],u_xpb_out[91][397],u_xpb_out[92][397],u_xpb_out[93][397],u_xpb_out[94][397],u_xpb_out[95][397],u_xpb_out[96][397],u_xpb_out[97][397],u_xpb_out[98][397],u_xpb_out[99][397],u_xpb_out[100][397],u_xpb_out[101][397],u_xpb_out[102][397],u_xpb_out[103][397],u_xpb_out[104][397],u_xpb_out[105][397]};

assign col_out_398 = {u_xpb_out[0][398],u_xpb_out[1][398],u_xpb_out[2][398],u_xpb_out[3][398],u_xpb_out[4][398],u_xpb_out[5][398],u_xpb_out[6][398],u_xpb_out[7][398],u_xpb_out[8][398],u_xpb_out[9][398],u_xpb_out[10][398],u_xpb_out[11][398],u_xpb_out[12][398],u_xpb_out[13][398],u_xpb_out[14][398],u_xpb_out[15][398],u_xpb_out[16][398],u_xpb_out[17][398],u_xpb_out[18][398],u_xpb_out[19][398],u_xpb_out[20][398],u_xpb_out[21][398],u_xpb_out[22][398],u_xpb_out[23][398],u_xpb_out[24][398],u_xpb_out[25][398],u_xpb_out[26][398],u_xpb_out[27][398],u_xpb_out[28][398],u_xpb_out[29][398],u_xpb_out[30][398],u_xpb_out[31][398],u_xpb_out[32][398],u_xpb_out[33][398],u_xpb_out[34][398],u_xpb_out[35][398],u_xpb_out[36][398],u_xpb_out[37][398],u_xpb_out[38][398],u_xpb_out[39][398],u_xpb_out[40][398],u_xpb_out[41][398],u_xpb_out[42][398],u_xpb_out[43][398],u_xpb_out[44][398],u_xpb_out[45][398],u_xpb_out[46][398],u_xpb_out[47][398],u_xpb_out[48][398],u_xpb_out[49][398],u_xpb_out[50][398],u_xpb_out[51][398],u_xpb_out[52][398],u_xpb_out[53][398],u_xpb_out[54][398],u_xpb_out[55][398],u_xpb_out[56][398],u_xpb_out[57][398],u_xpb_out[58][398],u_xpb_out[59][398],u_xpb_out[60][398],u_xpb_out[61][398],u_xpb_out[62][398],u_xpb_out[63][398],u_xpb_out[64][398],u_xpb_out[65][398],u_xpb_out[66][398],u_xpb_out[67][398],u_xpb_out[68][398],u_xpb_out[69][398],u_xpb_out[70][398],u_xpb_out[71][398],u_xpb_out[72][398],u_xpb_out[73][398],u_xpb_out[74][398],u_xpb_out[75][398],u_xpb_out[76][398],u_xpb_out[77][398],u_xpb_out[78][398],u_xpb_out[79][398],u_xpb_out[80][398],u_xpb_out[81][398],u_xpb_out[82][398],u_xpb_out[83][398],u_xpb_out[84][398],u_xpb_out[85][398],u_xpb_out[86][398],u_xpb_out[87][398],u_xpb_out[88][398],u_xpb_out[89][398],u_xpb_out[90][398],u_xpb_out[91][398],u_xpb_out[92][398],u_xpb_out[93][398],u_xpb_out[94][398],u_xpb_out[95][398],u_xpb_out[96][398],u_xpb_out[97][398],u_xpb_out[98][398],u_xpb_out[99][398],u_xpb_out[100][398],u_xpb_out[101][398],u_xpb_out[102][398],u_xpb_out[103][398],u_xpb_out[104][398],u_xpb_out[105][398]};

assign col_out_399 = {u_xpb_out[0][399],u_xpb_out[1][399],u_xpb_out[2][399],u_xpb_out[3][399],u_xpb_out[4][399],u_xpb_out[5][399],u_xpb_out[6][399],u_xpb_out[7][399],u_xpb_out[8][399],u_xpb_out[9][399],u_xpb_out[10][399],u_xpb_out[11][399],u_xpb_out[12][399],u_xpb_out[13][399],u_xpb_out[14][399],u_xpb_out[15][399],u_xpb_out[16][399],u_xpb_out[17][399],u_xpb_out[18][399],u_xpb_out[19][399],u_xpb_out[20][399],u_xpb_out[21][399],u_xpb_out[22][399],u_xpb_out[23][399],u_xpb_out[24][399],u_xpb_out[25][399],u_xpb_out[26][399],u_xpb_out[27][399],u_xpb_out[28][399],u_xpb_out[29][399],u_xpb_out[30][399],u_xpb_out[31][399],u_xpb_out[32][399],u_xpb_out[33][399],u_xpb_out[34][399],u_xpb_out[35][399],u_xpb_out[36][399],u_xpb_out[37][399],u_xpb_out[38][399],u_xpb_out[39][399],u_xpb_out[40][399],u_xpb_out[41][399],u_xpb_out[42][399],u_xpb_out[43][399],u_xpb_out[44][399],u_xpb_out[45][399],u_xpb_out[46][399],u_xpb_out[47][399],u_xpb_out[48][399],u_xpb_out[49][399],u_xpb_out[50][399],u_xpb_out[51][399],u_xpb_out[52][399],u_xpb_out[53][399],u_xpb_out[54][399],u_xpb_out[55][399],u_xpb_out[56][399],u_xpb_out[57][399],u_xpb_out[58][399],u_xpb_out[59][399],u_xpb_out[60][399],u_xpb_out[61][399],u_xpb_out[62][399],u_xpb_out[63][399],u_xpb_out[64][399],u_xpb_out[65][399],u_xpb_out[66][399],u_xpb_out[67][399],u_xpb_out[68][399],u_xpb_out[69][399],u_xpb_out[70][399],u_xpb_out[71][399],u_xpb_out[72][399],u_xpb_out[73][399],u_xpb_out[74][399],u_xpb_out[75][399],u_xpb_out[76][399],u_xpb_out[77][399],u_xpb_out[78][399],u_xpb_out[79][399],u_xpb_out[80][399],u_xpb_out[81][399],u_xpb_out[82][399],u_xpb_out[83][399],u_xpb_out[84][399],u_xpb_out[85][399],u_xpb_out[86][399],u_xpb_out[87][399],u_xpb_out[88][399],u_xpb_out[89][399],u_xpb_out[90][399],u_xpb_out[91][399],u_xpb_out[92][399],u_xpb_out[93][399],u_xpb_out[94][399],u_xpb_out[95][399],u_xpb_out[96][399],u_xpb_out[97][399],u_xpb_out[98][399],u_xpb_out[99][399],u_xpb_out[100][399],u_xpb_out[101][399],u_xpb_out[102][399],u_xpb_out[103][399],u_xpb_out[104][399],u_xpb_out[105][399]};

assign col_out_400 = {u_xpb_out[0][400],u_xpb_out[1][400],u_xpb_out[2][400],u_xpb_out[3][400],u_xpb_out[4][400],u_xpb_out[5][400],u_xpb_out[6][400],u_xpb_out[7][400],u_xpb_out[8][400],u_xpb_out[9][400],u_xpb_out[10][400],u_xpb_out[11][400],u_xpb_out[12][400],u_xpb_out[13][400],u_xpb_out[14][400],u_xpb_out[15][400],u_xpb_out[16][400],u_xpb_out[17][400],u_xpb_out[18][400],u_xpb_out[19][400],u_xpb_out[20][400],u_xpb_out[21][400],u_xpb_out[22][400],u_xpb_out[23][400],u_xpb_out[24][400],u_xpb_out[25][400],u_xpb_out[26][400],u_xpb_out[27][400],u_xpb_out[28][400],u_xpb_out[29][400],u_xpb_out[30][400],u_xpb_out[31][400],u_xpb_out[32][400],u_xpb_out[33][400],u_xpb_out[34][400],u_xpb_out[35][400],u_xpb_out[36][400],u_xpb_out[37][400],u_xpb_out[38][400],u_xpb_out[39][400],u_xpb_out[40][400],u_xpb_out[41][400],u_xpb_out[42][400],u_xpb_out[43][400],u_xpb_out[44][400],u_xpb_out[45][400],u_xpb_out[46][400],u_xpb_out[47][400],u_xpb_out[48][400],u_xpb_out[49][400],u_xpb_out[50][400],u_xpb_out[51][400],u_xpb_out[52][400],u_xpb_out[53][400],u_xpb_out[54][400],u_xpb_out[55][400],u_xpb_out[56][400],u_xpb_out[57][400],u_xpb_out[58][400],u_xpb_out[59][400],u_xpb_out[60][400],u_xpb_out[61][400],u_xpb_out[62][400],u_xpb_out[63][400],u_xpb_out[64][400],u_xpb_out[65][400],u_xpb_out[66][400],u_xpb_out[67][400],u_xpb_out[68][400],u_xpb_out[69][400],u_xpb_out[70][400],u_xpb_out[71][400],u_xpb_out[72][400],u_xpb_out[73][400],u_xpb_out[74][400],u_xpb_out[75][400],u_xpb_out[76][400],u_xpb_out[77][400],u_xpb_out[78][400],u_xpb_out[79][400],u_xpb_out[80][400],u_xpb_out[81][400],u_xpb_out[82][400],u_xpb_out[83][400],u_xpb_out[84][400],u_xpb_out[85][400],u_xpb_out[86][400],u_xpb_out[87][400],u_xpb_out[88][400],u_xpb_out[89][400],u_xpb_out[90][400],u_xpb_out[91][400],u_xpb_out[92][400],u_xpb_out[93][400],u_xpb_out[94][400],u_xpb_out[95][400],u_xpb_out[96][400],u_xpb_out[97][400],u_xpb_out[98][400],u_xpb_out[99][400],u_xpb_out[100][400],u_xpb_out[101][400],u_xpb_out[102][400],u_xpb_out[103][400],u_xpb_out[104][400],u_xpb_out[105][400]};

assign col_out_401 = {u_xpb_out[0][401],u_xpb_out[1][401],u_xpb_out[2][401],u_xpb_out[3][401],u_xpb_out[4][401],u_xpb_out[5][401],u_xpb_out[6][401],u_xpb_out[7][401],u_xpb_out[8][401],u_xpb_out[9][401],u_xpb_out[10][401],u_xpb_out[11][401],u_xpb_out[12][401],u_xpb_out[13][401],u_xpb_out[14][401],u_xpb_out[15][401],u_xpb_out[16][401],u_xpb_out[17][401],u_xpb_out[18][401],u_xpb_out[19][401],u_xpb_out[20][401],u_xpb_out[21][401],u_xpb_out[22][401],u_xpb_out[23][401],u_xpb_out[24][401],u_xpb_out[25][401],u_xpb_out[26][401],u_xpb_out[27][401],u_xpb_out[28][401],u_xpb_out[29][401],u_xpb_out[30][401],u_xpb_out[31][401],u_xpb_out[32][401],u_xpb_out[33][401],u_xpb_out[34][401],u_xpb_out[35][401],u_xpb_out[36][401],u_xpb_out[37][401],u_xpb_out[38][401],u_xpb_out[39][401],u_xpb_out[40][401],u_xpb_out[41][401],u_xpb_out[42][401],u_xpb_out[43][401],u_xpb_out[44][401],u_xpb_out[45][401],u_xpb_out[46][401],u_xpb_out[47][401],u_xpb_out[48][401],u_xpb_out[49][401],u_xpb_out[50][401],u_xpb_out[51][401],u_xpb_out[52][401],u_xpb_out[53][401],u_xpb_out[54][401],u_xpb_out[55][401],u_xpb_out[56][401],u_xpb_out[57][401],u_xpb_out[58][401],u_xpb_out[59][401],u_xpb_out[60][401],u_xpb_out[61][401],u_xpb_out[62][401],u_xpb_out[63][401],u_xpb_out[64][401],u_xpb_out[65][401],u_xpb_out[66][401],u_xpb_out[67][401],u_xpb_out[68][401],u_xpb_out[69][401],u_xpb_out[70][401],u_xpb_out[71][401],u_xpb_out[72][401],u_xpb_out[73][401],u_xpb_out[74][401],u_xpb_out[75][401],u_xpb_out[76][401],u_xpb_out[77][401],u_xpb_out[78][401],u_xpb_out[79][401],u_xpb_out[80][401],u_xpb_out[81][401],u_xpb_out[82][401],u_xpb_out[83][401],u_xpb_out[84][401],u_xpb_out[85][401],u_xpb_out[86][401],u_xpb_out[87][401],u_xpb_out[88][401],u_xpb_out[89][401],u_xpb_out[90][401],u_xpb_out[91][401],u_xpb_out[92][401],u_xpb_out[93][401],u_xpb_out[94][401],u_xpb_out[95][401],u_xpb_out[96][401],u_xpb_out[97][401],u_xpb_out[98][401],u_xpb_out[99][401],u_xpb_out[100][401],u_xpb_out[101][401],u_xpb_out[102][401],u_xpb_out[103][401],u_xpb_out[104][401],u_xpb_out[105][401]};

assign col_out_402 = {u_xpb_out[0][402],u_xpb_out[1][402],u_xpb_out[2][402],u_xpb_out[3][402],u_xpb_out[4][402],u_xpb_out[5][402],u_xpb_out[6][402],u_xpb_out[7][402],u_xpb_out[8][402],u_xpb_out[9][402],u_xpb_out[10][402],u_xpb_out[11][402],u_xpb_out[12][402],u_xpb_out[13][402],u_xpb_out[14][402],u_xpb_out[15][402],u_xpb_out[16][402],u_xpb_out[17][402],u_xpb_out[18][402],u_xpb_out[19][402],u_xpb_out[20][402],u_xpb_out[21][402],u_xpb_out[22][402],u_xpb_out[23][402],u_xpb_out[24][402],u_xpb_out[25][402],u_xpb_out[26][402],u_xpb_out[27][402],u_xpb_out[28][402],u_xpb_out[29][402],u_xpb_out[30][402],u_xpb_out[31][402],u_xpb_out[32][402],u_xpb_out[33][402],u_xpb_out[34][402],u_xpb_out[35][402],u_xpb_out[36][402],u_xpb_out[37][402],u_xpb_out[38][402],u_xpb_out[39][402],u_xpb_out[40][402],u_xpb_out[41][402],u_xpb_out[42][402],u_xpb_out[43][402],u_xpb_out[44][402],u_xpb_out[45][402],u_xpb_out[46][402],u_xpb_out[47][402],u_xpb_out[48][402],u_xpb_out[49][402],u_xpb_out[50][402],u_xpb_out[51][402],u_xpb_out[52][402],u_xpb_out[53][402],u_xpb_out[54][402],u_xpb_out[55][402],u_xpb_out[56][402],u_xpb_out[57][402],u_xpb_out[58][402],u_xpb_out[59][402],u_xpb_out[60][402],u_xpb_out[61][402],u_xpb_out[62][402],u_xpb_out[63][402],u_xpb_out[64][402],u_xpb_out[65][402],u_xpb_out[66][402],u_xpb_out[67][402],u_xpb_out[68][402],u_xpb_out[69][402],u_xpb_out[70][402],u_xpb_out[71][402],u_xpb_out[72][402],u_xpb_out[73][402],u_xpb_out[74][402],u_xpb_out[75][402],u_xpb_out[76][402],u_xpb_out[77][402],u_xpb_out[78][402],u_xpb_out[79][402],u_xpb_out[80][402],u_xpb_out[81][402],u_xpb_out[82][402],u_xpb_out[83][402],u_xpb_out[84][402],u_xpb_out[85][402],u_xpb_out[86][402],u_xpb_out[87][402],u_xpb_out[88][402],u_xpb_out[89][402],u_xpb_out[90][402],u_xpb_out[91][402],u_xpb_out[92][402],u_xpb_out[93][402],u_xpb_out[94][402],u_xpb_out[95][402],u_xpb_out[96][402],u_xpb_out[97][402],u_xpb_out[98][402],u_xpb_out[99][402],u_xpb_out[100][402],u_xpb_out[101][402],u_xpb_out[102][402],u_xpb_out[103][402],u_xpb_out[104][402],u_xpb_out[105][402]};

assign col_out_403 = {u_xpb_out[0][403],u_xpb_out[1][403],u_xpb_out[2][403],u_xpb_out[3][403],u_xpb_out[4][403],u_xpb_out[5][403],u_xpb_out[6][403],u_xpb_out[7][403],u_xpb_out[8][403],u_xpb_out[9][403],u_xpb_out[10][403],u_xpb_out[11][403],u_xpb_out[12][403],u_xpb_out[13][403],u_xpb_out[14][403],u_xpb_out[15][403],u_xpb_out[16][403],u_xpb_out[17][403],u_xpb_out[18][403],u_xpb_out[19][403],u_xpb_out[20][403],u_xpb_out[21][403],u_xpb_out[22][403],u_xpb_out[23][403],u_xpb_out[24][403],u_xpb_out[25][403],u_xpb_out[26][403],u_xpb_out[27][403],u_xpb_out[28][403],u_xpb_out[29][403],u_xpb_out[30][403],u_xpb_out[31][403],u_xpb_out[32][403],u_xpb_out[33][403],u_xpb_out[34][403],u_xpb_out[35][403],u_xpb_out[36][403],u_xpb_out[37][403],u_xpb_out[38][403],u_xpb_out[39][403],u_xpb_out[40][403],u_xpb_out[41][403],u_xpb_out[42][403],u_xpb_out[43][403],u_xpb_out[44][403],u_xpb_out[45][403],u_xpb_out[46][403],u_xpb_out[47][403],u_xpb_out[48][403],u_xpb_out[49][403],u_xpb_out[50][403],u_xpb_out[51][403],u_xpb_out[52][403],u_xpb_out[53][403],u_xpb_out[54][403],u_xpb_out[55][403],u_xpb_out[56][403],u_xpb_out[57][403],u_xpb_out[58][403],u_xpb_out[59][403],u_xpb_out[60][403],u_xpb_out[61][403],u_xpb_out[62][403],u_xpb_out[63][403],u_xpb_out[64][403],u_xpb_out[65][403],u_xpb_out[66][403],u_xpb_out[67][403],u_xpb_out[68][403],u_xpb_out[69][403],u_xpb_out[70][403],u_xpb_out[71][403],u_xpb_out[72][403],u_xpb_out[73][403],u_xpb_out[74][403],u_xpb_out[75][403],u_xpb_out[76][403],u_xpb_out[77][403],u_xpb_out[78][403],u_xpb_out[79][403],u_xpb_out[80][403],u_xpb_out[81][403],u_xpb_out[82][403],u_xpb_out[83][403],u_xpb_out[84][403],u_xpb_out[85][403],u_xpb_out[86][403],u_xpb_out[87][403],u_xpb_out[88][403],u_xpb_out[89][403],u_xpb_out[90][403],u_xpb_out[91][403],u_xpb_out[92][403],u_xpb_out[93][403],u_xpb_out[94][403],u_xpb_out[95][403],u_xpb_out[96][403],u_xpb_out[97][403],u_xpb_out[98][403],u_xpb_out[99][403],u_xpb_out[100][403],u_xpb_out[101][403],u_xpb_out[102][403],u_xpb_out[103][403],u_xpb_out[104][403],u_xpb_out[105][403]};

assign col_out_404 = {u_xpb_out[0][404],u_xpb_out[1][404],u_xpb_out[2][404],u_xpb_out[3][404],u_xpb_out[4][404],u_xpb_out[5][404],u_xpb_out[6][404],u_xpb_out[7][404],u_xpb_out[8][404],u_xpb_out[9][404],u_xpb_out[10][404],u_xpb_out[11][404],u_xpb_out[12][404],u_xpb_out[13][404],u_xpb_out[14][404],u_xpb_out[15][404],u_xpb_out[16][404],u_xpb_out[17][404],u_xpb_out[18][404],u_xpb_out[19][404],u_xpb_out[20][404],u_xpb_out[21][404],u_xpb_out[22][404],u_xpb_out[23][404],u_xpb_out[24][404],u_xpb_out[25][404],u_xpb_out[26][404],u_xpb_out[27][404],u_xpb_out[28][404],u_xpb_out[29][404],u_xpb_out[30][404],u_xpb_out[31][404],u_xpb_out[32][404],u_xpb_out[33][404],u_xpb_out[34][404],u_xpb_out[35][404],u_xpb_out[36][404],u_xpb_out[37][404],u_xpb_out[38][404],u_xpb_out[39][404],u_xpb_out[40][404],u_xpb_out[41][404],u_xpb_out[42][404],u_xpb_out[43][404],u_xpb_out[44][404],u_xpb_out[45][404],u_xpb_out[46][404],u_xpb_out[47][404],u_xpb_out[48][404],u_xpb_out[49][404],u_xpb_out[50][404],u_xpb_out[51][404],u_xpb_out[52][404],u_xpb_out[53][404],u_xpb_out[54][404],u_xpb_out[55][404],u_xpb_out[56][404],u_xpb_out[57][404],u_xpb_out[58][404],u_xpb_out[59][404],u_xpb_out[60][404],u_xpb_out[61][404],u_xpb_out[62][404],u_xpb_out[63][404],u_xpb_out[64][404],u_xpb_out[65][404],u_xpb_out[66][404],u_xpb_out[67][404],u_xpb_out[68][404],u_xpb_out[69][404],u_xpb_out[70][404],u_xpb_out[71][404],u_xpb_out[72][404],u_xpb_out[73][404],u_xpb_out[74][404],u_xpb_out[75][404],u_xpb_out[76][404],u_xpb_out[77][404],u_xpb_out[78][404],u_xpb_out[79][404],u_xpb_out[80][404],u_xpb_out[81][404],u_xpb_out[82][404],u_xpb_out[83][404],u_xpb_out[84][404],u_xpb_out[85][404],u_xpb_out[86][404],u_xpb_out[87][404],u_xpb_out[88][404],u_xpb_out[89][404],u_xpb_out[90][404],u_xpb_out[91][404],u_xpb_out[92][404],u_xpb_out[93][404],u_xpb_out[94][404],u_xpb_out[95][404],u_xpb_out[96][404],u_xpb_out[97][404],u_xpb_out[98][404],u_xpb_out[99][404],u_xpb_out[100][404],u_xpb_out[101][404],u_xpb_out[102][404],u_xpb_out[103][404],u_xpb_out[104][404],u_xpb_out[105][404]};

assign col_out_405 = {u_xpb_out[0][405],u_xpb_out[1][405],u_xpb_out[2][405],u_xpb_out[3][405],u_xpb_out[4][405],u_xpb_out[5][405],u_xpb_out[6][405],u_xpb_out[7][405],u_xpb_out[8][405],u_xpb_out[9][405],u_xpb_out[10][405],u_xpb_out[11][405],u_xpb_out[12][405],u_xpb_out[13][405],u_xpb_out[14][405],u_xpb_out[15][405],u_xpb_out[16][405],u_xpb_out[17][405],u_xpb_out[18][405],u_xpb_out[19][405],u_xpb_out[20][405],u_xpb_out[21][405],u_xpb_out[22][405],u_xpb_out[23][405],u_xpb_out[24][405],u_xpb_out[25][405],u_xpb_out[26][405],u_xpb_out[27][405],u_xpb_out[28][405],u_xpb_out[29][405],u_xpb_out[30][405],u_xpb_out[31][405],u_xpb_out[32][405],u_xpb_out[33][405],u_xpb_out[34][405],u_xpb_out[35][405],u_xpb_out[36][405],u_xpb_out[37][405],u_xpb_out[38][405],u_xpb_out[39][405],u_xpb_out[40][405],u_xpb_out[41][405],u_xpb_out[42][405],u_xpb_out[43][405],u_xpb_out[44][405],u_xpb_out[45][405],u_xpb_out[46][405],u_xpb_out[47][405],u_xpb_out[48][405],u_xpb_out[49][405],u_xpb_out[50][405],u_xpb_out[51][405],u_xpb_out[52][405],u_xpb_out[53][405],u_xpb_out[54][405],u_xpb_out[55][405],u_xpb_out[56][405],u_xpb_out[57][405],u_xpb_out[58][405],u_xpb_out[59][405],u_xpb_out[60][405],u_xpb_out[61][405],u_xpb_out[62][405],u_xpb_out[63][405],u_xpb_out[64][405],u_xpb_out[65][405],u_xpb_out[66][405],u_xpb_out[67][405],u_xpb_out[68][405],u_xpb_out[69][405],u_xpb_out[70][405],u_xpb_out[71][405],u_xpb_out[72][405],u_xpb_out[73][405],u_xpb_out[74][405],u_xpb_out[75][405],u_xpb_out[76][405],u_xpb_out[77][405],u_xpb_out[78][405],u_xpb_out[79][405],u_xpb_out[80][405],u_xpb_out[81][405],u_xpb_out[82][405],u_xpb_out[83][405],u_xpb_out[84][405],u_xpb_out[85][405],u_xpb_out[86][405],u_xpb_out[87][405],u_xpb_out[88][405],u_xpb_out[89][405],u_xpb_out[90][405],u_xpb_out[91][405],u_xpb_out[92][405],u_xpb_out[93][405],u_xpb_out[94][405],u_xpb_out[95][405],u_xpb_out[96][405],u_xpb_out[97][405],u_xpb_out[98][405],u_xpb_out[99][405],u_xpb_out[100][405],u_xpb_out[101][405],u_xpb_out[102][405],u_xpb_out[103][405],u_xpb_out[104][405],u_xpb_out[105][405]};

assign col_out_406 = {u_xpb_out[0][406],u_xpb_out[1][406],u_xpb_out[2][406],u_xpb_out[3][406],u_xpb_out[4][406],u_xpb_out[5][406],u_xpb_out[6][406],u_xpb_out[7][406],u_xpb_out[8][406],u_xpb_out[9][406],u_xpb_out[10][406],u_xpb_out[11][406],u_xpb_out[12][406],u_xpb_out[13][406],u_xpb_out[14][406],u_xpb_out[15][406],u_xpb_out[16][406],u_xpb_out[17][406],u_xpb_out[18][406],u_xpb_out[19][406],u_xpb_out[20][406],u_xpb_out[21][406],u_xpb_out[22][406],u_xpb_out[23][406],u_xpb_out[24][406],u_xpb_out[25][406],u_xpb_out[26][406],u_xpb_out[27][406],u_xpb_out[28][406],u_xpb_out[29][406],u_xpb_out[30][406],u_xpb_out[31][406],u_xpb_out[32][406],u_xpb_out[33][406],u_xpb_out[34][406],u_xpb_out[35][406],u_xpb_out[36][406],u_xpb_out[37][406],u_xpb_out[38][406],u_xpb_out[39][406],u_xpb_out[40][406],u_xpb_out[41][406],u_xpb_out[42][406],u_xpb_out[43][406],u_xpb_out[44][406],u_xpb_out[45][406],u_xpb_out[46][406],u_xpb_out[47][406],u_xpb_out[48][406],u_xpb_out[49][406],u_xpb_out[50][406],u_xpb_out[51][406],u_xpb_out[52][406],u_xpb_out[53][406],u_xpb_out[54][406],u_xpb_out[55][406],u_xpb_out[56][406],u_xpb_out[57][406],u_xpb_out[58][406],u_xpb_out[59][406],u_xpb_out[60][406],u_xpb_out[61][406],u_xpb_out[62][406],u_xpb_out[63][406],u_xpb_out[64][406],u_xpb_out[65][406],u_xpb_out[66][406],u_xpb_out[67][406],u_xpb_out[68][406],u_xpb_out[69][406],u_xpb_out[70][406],u_xpb_out[71][406],u_xpb_out[72][406],u_xpb_out[73][406],u_xpb_out[74][406],u_xpb_out[75][406],u_xpb_out[76][406],u_xpb_out[77][406],u_xpb_out[78][406],u_xpb_out[79][406],u_xpb_out[80][406],u_xpb_out[81][406],u_xpb_out[82][406],u_xpb_out[83][406],u_xpb_out[84][406],u_xpb_out[85][406],u_xpb_out[86][406],u_xpb_out[87][406],u_xpb_out[88][406],u_xpb_out[89][406],u_xpb_out[90][406],u_xpb_out[91][406],u_xpb_out[92][406],u_xpb_out[93][406],u_xpb_out[94][406],u_xpb_out[95][406],u_xpb_out[96][406],u_xpb_out[97][406],u_xpb_out[98][406],u_xpb_out[99][406],u_xpb_out[100][406],u_xpb_out[101][406],u_xpb_out[102][406],u_xpb_out[103][406],u_xpb_out[104][406],u_xpb_out[105][406]};

assign col_out_407 = {u_xpb_out[0][407],u_xpb_out[1][407],u_xpb_out[2][407],u_xpb_out[3][407],u_xpb_out[4][407],u_xpb_out[5][407],u_xpb_out[6][407],u_xpb_out[7][407],u_xpb_out[8][407],u_xpb_out[9][407],u_xpb_out[10][407],u_xpb_out[11][407],u_xpb_out[12][407],u_xpb_out[13][407],u_xpb_out[14][407],u_xpb_out[15][407],u_xpb_out[16][407],u_xpb_out[17][407],u_xpb_out[18][407],u_xpb_out[19][407],u_xpb_out[20][407],u_xpb_out[21][407],u_xpb_out[22][407],u_xpb_out[23][407],u_xpb_out[24][407],u_xpb_out[25][407],u_xpb_out[26][407],u_xpb_out[27][407],u_xpb_out[28][407],u_xpb_out[29][407],u_xpb_out[30][407],u_xpb_out[31][407],u_xpb_out[32][407],u_xpb_out[33][407],u_xpb_out[34][407],u_xpb_out[35][407],u_xpb_out[36][407],u_xpb_out[37][407],u_xpb_out[38][407],u_xpb_out[39][407],u_xpb_out[40][407],u_xpb_out[41][407],u_xpb_out[42][407],u_xpb_out[43][407],u_xpb_out[44][407],u_xpb_out[45][407],u_xpb_out[46][407],u_xpb_out[47][407],u_xpb_out[48][407],u_xpb_out[49][407],u_xpb_out[50][407],u_xpb_out[51][407],u_xpb_out[52][407],u_xpb_out[53][407],u_xpb_out[54][407],u_xpb_out[55][407],u_xpb_out[56][407],u_xpb_out[57][407],u_xpb_out[58][407],u_xpb_out[59][407],u_xpb_out[60][407],u_xpb_out[61][407],u_xpb_out[62][407],u_xpb_out[63][407],u_xpb_out[64][407],u_xpb_out[65][407],u_xpb_out[66][407],u_xpb_out[67][407],u_xpb_out[68][407],u_xpb_out[69][407],u_xpb_out[70][407],u_xpb_out[71][407],u_xpb_out[72][407],u_xpb_out[73][407],u_xpb_out[74][407],u_xpb_out[75][407],u_xpb_out[76][407],u_xpb_out[77][407],u_xpb_out[78][407],u_xpb_out[79][407],u_xpb_out[80][407],u_xpb_out[81][407],u_xpb_out[82][407],u_xpb_out[83][407],u_xpb_out[84][407],u_xpb_out[85][407],u_xpb_out[86][407],u_xpb_out[87][407],u_xpb_out[88][407],u_xpb_out[89][407],u_xpb_out[90][407],u_xpb_out[91][407],u_xpb_out[92][407],u_xpb_out[93][407],u_xpb_out[94][407],u_xpb_out[95][407],u_xpb_out[96][407],u_xpb_out[97][407],u_xpb_out[98][407],u_xpb_out[99][407],u_xpb_out[100][407],u_xpb_out[101][407],u_xpb_out[102][407],u_xpb_out[103][407],u_xpb_out[104][407],u_xpb_out[105][407]};

assign col_out_408 = {u_xpb_out[0][408],u_xpb_out[1][408],u_xpb_out[2][408],u_xpb_out[3][408],u_xpb_out[4][408],u_xpb_out[5][408],u_xpb_out[6][408],u_xpb_out[7][408],u_xpb_out[8][408],u_xpb_out[9][408],u_xpb_out[10][408],u_xpb_out[11][408],u_xpb_out[12][408],u_xpb_out[13][408],u_xpb_out[14][408],u_xpb_out[15][408],u_xpb_out[16][408],u_xpb_out[17][408],u_xpb_out[18][408],u_xpb_out[19][408],u_xpb_out[20][408],u_xpb_out[21][408],u_xpb_out[22][408],u_xpb_out[23][408],u_xpb_out[24][408],u_xpb_out[25][408],u_xpb_out[26][408],u_xpb_out[27][408],u_xpb_out[28][408],u_xpb_out[29][408],u_xpb_out[30][408],u_xpb_out[31][408],u_xpb_out[32][408],u_xpb_out[33][408],u_xpb_out[34][408],u_xpb_out[35][408],u_xpb_out[36][408],u_xpb_out[37][408],u_xpb_out[38][408],u_xpb_out[39][408],u_xpb_out[40][408],u_xpb_out[41][408],u_xpb_out[42][408],u_xpb_out[43][408],u_xpb_out[44][408],u_xpb_out[45][408],u_xpb_out[46][408],u_xpb_out[47][408],u_xpb_out[48][408],u_xpb_out[49][408],u_xpb_out[50][408],u_xpb_out[51][408],u_xpb_out[52][408],u_xpb_out[53][408],u_xpb_out[54][408],u_xpb_out[55][408],u_xpb_out[56][408],u_xpb_out[57][408],u_xpb_out[58][408],u_xpb_out[59][408],u_xpb_out[60][408],u_xpb_out[61][408],u_xpb_out[62][408],u_xpb_out[63][408],u_xpb_out[64][408],u_xpb_out[65][408],u_xpb_out[66][408],u_xpb_out[67][408],u_xpb_out[68][408],u_xpb_out[69][408],u_xpb_out[70][408],u_xpb_out[71][408],u_xpb_out[72][408],u_xpb_out[73][408],u_xpb_out[74][408],u_xpb_out[75][408],u_xpb_out[76][408],u_xpb_out[77][408],u_xpb_out[78][408],u_xpb_out[79][408],u_xpb_out[80][408],u_xpb_out[81][408],u_xpb_out[82][408],u_xpb_out[83][408],u_xpb_out[84][408],u_xpb_out[85][408],u_xpb_out[86][408],u_xpb_out[87][408],u_xpb_out[88][408],u_xpb_out[89][408],u_xpb_out[90][408],u_xpb_out[91][408],u_xpb_out[92][408],u_xpb_out[93][408],u_xpb_out[94][408],u_xpb_out[95][408],u_xpb_out[96][408],u_xpb_out[97][408],u_xpb_out[98][408],u_xpb_out[99][408],u_xpb_out[100][408],u_xpb_out[101][408],u_xpb_out[102][408],u_xpb_out[103][408],u_xpb_out[104][408],u_xpb_out[105][408]};

assign col_out_409 = {u_xpb_out[0][409],u_xpb_out[1][409],u_xpb_out[2][409],u_xpb_out[3][409],u_xpb_out[4][409],u_xpb_out[5][409],u_xpb_out[6][409],u_xpb_out[7][409],u_xpb_out[8][409],u_xpb_out[9][409],u_xpb_out[10][409],u_xpb_out[11][409],u_xpb_out[12][409],u_xpb_out[13][409],u_xpb_out[14][409],u_xpb_out[15][409],u_xpb_out[16][409],u_xpb_out[17][409],u_xpb_out[18][409],u_xpb_out[19][409],u_xpb_out[20][409],u_xpb_out[21][409],u_xpb_out[22][409],u_xpb_out[23][409],u_xpb_out[24][409],u_xpb_out[25][409],u_xpb_out[26][409],u_xpb_out[27][409],u_xpb_out[28][409],u_xpb_out[29][409],u_xpb_out[30][409],u_xpb_out[31][409],u_xpb_out[32][409],u_xpb_out[33][409],u_xpb_out[34][409],u_xpb_out[35][409],u_xpb_out[36][409],u_xpb_out[37][409],u_xpb_out[38][409],u_xpb_out[39][409],u_xpb_out[40][409],u_xpb_out[41][409],u_xpb_out[42][409],u_xpb_out[43][409],u_xpb_out[44][409],u_xpb_out[45][409],u_xpb_out[46][409],u_xpb_out[47][409],u_xpb_out[48][409],u_xpb_out[49][409],u_xpb_out[50][409],u_xpb_out[51][409],u_xpb_out[52][409],u_xpb_out[53][409],u_xpb_out[54][409],u_xpb_out[55][409],u_xpb_out[56][409],u_xpb_out[57][409],u_xpb_out[58][409],u_xpb_out[59][409],u_xpb_out[60][409],u_xpb_out[61][409],u_xpb_out[62][409],u_xpb_out[63][409],u_xpb_out[64][409],u_xpb_out[65][409],u_xpb_out[66][409],u_xpb_out[67][409],u_xpb_out[68][409],u_xpb_out[69][409],u_xpb_out[70][409],u_xpb_out[71][409],u_xpb_out[72][409],u_xpb_out[73][409],u_xpb_out[74][409],u_xpb_out[75][409],u_xpb_out[76][409],u_xpb_out[77][409],u_xpb_out[78][409],u_xpb_out[79][409],u_xpb_out[80][409],u_xpb_out[81][409],u_xpb_out[82][409],u_xpb_out[83][409],u_xpb_out[84][409],u_xpb_out[85][409],u_xpb_out[86][409],u_xpb_out[87][409],u_xpb_out[88][409],u_xpb_out[89][409],u_xpb_out[90][409],u_xpb_out[91][409],u_xpb_out[92][409],u_xpb_out[93][409],u_xpb_out[94][409],u_xpb_out[95][409],u_xpb_out[96][409],u_xpb_out[97][409],u_xpb_out[98][409],u_xpb_out[99][409],u_xpb_out[100][409],u_xpb_out[101][409],u_xpb_out[102][409],u_xpb_out[103][409],u_xpb_out[104][409],u_xpb_out[105][409]};

assign col_out_410 = {u_xpb_out[0][410],u_xpb_out[1][410],u_xpb_out[2][410],u_xpb_out[3][410],u_xpb_out[4][410],u_xpb_out[5][410],u_xpb_out[6][410],u_xpb_out[7][410],u_xpb_out[8][410],u_xpb_out[9][410],u_xpb_out[10][410],u_xpb_out[11][410],u_xpb_out[12][410],u_xpb_out[13][410],u_xpb_out[14][410],u_xpb_out[15][410],u_xpb_out[16][410],u_xpb_out[17][410],u_xpb_out[18][410],u_xpb_out[19][410],u_xpb_out[20][410],u_xpb_out[21][410],u_xpb_out[22][410],u_xpb_out[23][410],u_xpb_out[24][410],u_xpb_out[25][410],u_xpb_out[26][410],u_xpb_out[27][410],u_xpb_out[28][410],u_xpb_out[29][410],u_xpb_out[30][410],u_xpb_out[31][410],u_xpb_out[32][410],u_xpb_out[33][410],u_xpb_out[34][410],u_xpb_out[35][410],u_xpb_out[36][410],u_xpb_out[37][410],u_xpb_out[38][410],u_xpb_out[39][410],u_xpb_out[40][410],u_xpb_out[41][410],u_xpb_out[42][410],u_xpb_out[43][410],u_xpb_out[44][410],u_xpb_out[45][410],u_xpb_out[46][410],u_xpb_out[47][410],u_xpb_out[48][410],u_xpb_out[49][410],u_xpb_out[50][410],u_xpb_out[51][410],u_xpb_out[52][410],u_xpb_out[53][410],u_xpb_out[54][410],u_xpb_out[55][410],u_xpb_out[56][410],u_xpb_out[57][410],u_xpb_out[58][410],u_xpb_out[59][410],u_xpb_out[60][410],u_xpb_out[61][410],u_xpb_out[62][410],u_xpb_out[63][410],u_xpb_out[64][410],u_xpb_out[65][410],u_xpb_out[66][410],u_xpb_out[67][410],u_xpb_out[68][410],u_xpb_out[69][410],u_xpb_out[70][410],u_xpb_out[71][410],u_xpb_out[72][410],u_xpb_out[73][410],u_xpb_out[74][410],u_xpb_out[75][410],u_xpb_out[76][410],u_xpb_out[77][410],u_xpb_out[78][410],u_xpb_out[79][410],u_xpb_out[80][410],u_xpb_out[81][410],u_xpb_out[82][410],u_xpb_out[83][410],u_xpb_out[84][410],u_xpb_out[85][410],u_xpb_out[86][410],u_xpb_out[87][410],u_xpb_out[88][410],u_xpb_out[89][410],u_xpb_out[90][410],u_xpb_out[91][410],u_xpb_out[92][410],u_xpb_out[93][410],u_xpb_out[94][410],u_xpb_out[95][410],u_xpb_out[96][410],u_xpb_out[97][410],u_xpb_out[98][410],u_xpb_out[99][410],u_xpb_out[100][410],u_xpb_out[101][410],u_xpb_out[102][410],u_xpb_out[103][410],u_xpb_out[104][410],u_xpb_out[105][410]};

assign col_out_411 = {u_xpb_out[0][411],u_xpb_out[1][411],u_xpb_out[2][411],u_xpb_out[3][411],u_xpb_out[4][411],u_xpb_out[5][411],u_xpb_out[6][411],u_xpb_out[7][411],u_xpb_out[8][411],u_xpb_out[9][411],u_xpb_out[10][411],u_xpb_out[11][411],u_xpb_out[12][411],u_xpb_out[13][411],u_xpb_out[14][411],u_xpb_out[15][411],u_xpb_out[16][411],u_xpb_out[17][411],u_xpb_out[18][411],u_xpb_out[19][411],u_xpb_out[20][411],u_xpb_out[21][411],u_xpb_out[22][411],u_xpb_out[23][411],u_xpb_out[24][411],u_xpb_out[25][411],u_xpb_out[26][411],u_xpb_out[27][411],u_xpb_out[28][411],u_xpb_out[29][411],u_xpb_out[30][411],u_xpb_out[31][411],u_xpb_out[32][411],u_xpb_out[33][411],u_xpb_out[34][411],u_xpb_out[35][411],u_xpb_out[36][411],u_xpb_out[37][411],u_xpb_out[38][411],u_xpb_out[39][411],u_xpb_out[40][411],u_xpb_out[41][411],u_xpb_out[42][411],u_xpb_out[43][411],u_xpb_out[44][411],u_xpb_out[45][411],u_xpb_out[46][411],u_xpb_out[47][411],u_xpb_out[48][411],u_xpb_out[49][411],u_xpb_out[50][411],u_xpb_out[51][411],u_xpb_out[52][411],u_xpb_out[53][411],u_xpb_out[54][411],u_xpb_out[55][411],u_xpb_out[56][411],u_xpb_out[57][411],u_xpb_out[58][411],u_xpb_out[59][411],u_xpb_out[60][411],u_xpb_out[61][411],u_xpb_out[62][411],u_xpb_out[63][411],u_xpb_out[64][411],u_xpb_out[65][411],u_xpb_out[66][411],u_xpb_out[67][411],u_xpb_out[68][411],u_xpb_out[69][411],u_xpb_out[70][411],u_xpb_out[71][411],u_xpb_out[72][411],u_xpb_out[73][411],u_xpb_out[74][411],u_xpb_out[75][411],u_xpb_out[76][411],u_xpb_out[77][411],u_xpb_out[78][411],u_xpb_out[79][411],u_xpb_out[80][411],u_xpb_out[81][411],u_xpb_out[82][411],u_xpb_out[83][411],u_xpb_out[84][411],u_xpb_out[85][411],u_xpb_out[86][411],u_xpb_out[87][411],u_xpb_out[88][411],u_xpb_out[89][411],u_xpb_out[90][411],u_xpb_out[91][411],u_xpb_out[92][411],u_xpb_out[93][411],u_xpb_out[94][411],u_xpb_out[95][411],u_xpb_out[96][411],u_xpb_out[97][411],u_xpb_out[98][411],u_xpb_out[99][411],u_xpb_out[100][411],u_xpb_out[101][411],u_xpb_out[102][411],u_xpb_out[103][411],u_xpb_out[104][411],u_xpb_out[105][411]};

assign col_out_412 = {u_xpb_out[0][412],u_xpb_out[1][412],u_xpb_out[2][412],u_xpb_out[3][412],u_xpb_out[4][412],u_xpb_out[5][412],u_xpb_out[6][412],u_xpb_out[7][412],u_xpb_out[8][412],u_xpb_out[9][412],u_xpb_out[10][412],u_xpb_out[11][412],u_xpb_out[12][412],u_xpb_out[13][412],u_xpb_out[14][412],u_xpb_out[15][412],u_xpb_out[16][412],u_xpb_out[17][412],u_xpb_out[18][412],u_xpb_out[19][412],u_xpb_out[20][412],u_xpb_out[21][412],u_xpb_out[22][412],u_xpb_out[23][412],u_xpb_out[24][412],u_xpb_out[25][412],u_xpb_out[26][412],u_xpb_out[27][412],u_xpb_out[28][412],u_xpb_out[29][412],u_xpb_out[30][412],u_xpb_out[31][412],u_xpb_out[32][412],u_xpb_out[33][412],u_xpb_out[34][412],u_xpb_out[35][412],u_xpb_out[36][412],u_xpb_out[37][412],u_xpb_out[38][412],u_xpb_out[39][412],u_xpb_out[40][412],u_xpb_out[41][412],u_xpb_out[42][412],u_xpb_out[43][412],u_xpb_out[44][412],u_xpb_out[45][412],u_xpb_out[46][412],u_xpb_out[47][412],u_xpb_out[48][412],u_xpb_out[49][412],u_xpb_out[50][412],u_xpb_out[51][412],u_xpb_out[52][412],u_xpb_out[53][412],u_xpb_out[54][412],u_xpb_out[55][412],u_xpb_out[56][412],u_xpb_out[57][412],u_xpb_out[58][412],u_xpb_out[59][412],u_xpb_out[60][412],u_xpb_out[61][412],u_xpb_out[62][412],u_xpb_out[63][412],u_xpb_out[64][412],u_xpb_out[65][412],u_xpb_out[66][412],u_xpb_out[67][412],u_xpb_out[68][412],u_xpb_out[69][412],u_xpb_out[70][412],u_xpb_out[71][412],u_xpb_out[72][412],u_xpb_out[73][412],u_xpb_out[74][412],u_xpb_out[75][412],u_xpb_out[76][412],u_xpb_out[77][412],u_xpb_out[78][412],u_xpb_out[79][412],u_xpb_out[80][412],u_xpb_out[81][412],u_xpb_out[82][412],u_xpb_out[83][412],u_xpb_out[84][412],u_xpb_out[85][412],u_xpb_out[86][412],u_xpb_out[87][412],u_xpb_out[88][412],u_xpb_out[89][412],u_xpb_out[90][412],u_xpb_out[91][412],u_xpb_out[92][412],u_xpb_out[93][412],u_xpb_out[94][412],u_xpb_out[95][412],u_xpb_out[96][412],u_xpb_out[97][412],u_xpb_out[98][412],u_xpb_out[99][412],u_xpb_out[100][412],u_xpb_out[101][412],u_xpb_out[102][412],u_xpb_out[103][412],u_xpb_out[104][412],u_xpb_out[105][412]};

assign col_out_413 = {u_xpb_out[0][413],u_xpb_out[1][413],u_xpb_out[2][413],u_xpb_out[3][413],u_xpb_out[4][413],u_xpb_out[5][413],u_xpb_out[6][413],u_xpb_out[7][413],u_xpb_out[8][413],u_xpb_out[9][413],u_xpb_out[10][413],u_xpb_out[11][413],u_xpb_out[12][413],u_xpb_out[13][413],u_xpb_out[14][413],u_xpb_out[15][413],u_xpb_out[16][413],u_xpb_out[17][413],u_xpb_out[18][413],u_xpb_out[19][413],u_xpb_out[20][413],u_xpb_out[21][413],u_xpb_out[22][413],u_xpb_out[23][413],u_xpb_out[24][413],u_xpb_out[25][413],u_xpb_out[26][413],u_xpb_out[27][413],u_xpb_out[28][413],u_xpb_out[29][413],u_xpb_out[30][413],u_xpb_out[31][413],u_xpb_out[32][413],u_xpb_out[33][413],u_xpb_out[34][413],u_xpb_out[35][413],u_xpb_out[36][413],u_xpb_out[37][413],u_xpb_out[38][413],u_xpb_out[39][413],u_xpb_out[40][413],u_xpb_out[41][413],u_xpb_out[42][413],u_xpb_out[43][413],u_xpb_out[44][413],u_xpb_out[45][413],u_xpb_out[46][413],u_xpb_out[47][413],u_xpb_out[48][413],u_xpb_out[49][413],u_xpb_out[50][413],u_xpb_out[51][413],u_xpb_out[52][413],u_xpb_out[53][413],u_xpb_out[54][413],u_xpb_out[55][413],u_xpb_out[56][413],u_xpb_out[57][413],u_xpb_out[58][413],u_xpb_out[59][413],u_xpb_out[60][413],u_xpb_out[61][413],u_xpb_out[62][413],u_xpb_out[63][413],u_xpb_out[64][413],u_xpb_out[65][413],u_xpb_out[66][413],u_xpb_out[67][413],u_xpb_out[68][413],u_xpb_out[69][413],u_xpb_out[70][413],u_xpb_out[71][413],u_xpb_out[72][413],u_xpb_out[73][413],u_xpb_out[74][413],u_xpb_out[75][413],u_xpb_out[76][413],u_xpb_out[77][413],u_xpb_out[78][413],u_xpb_out[79][413],u_xpb_out[80][413],u_xpb_out[81][413],u_xpb_out[82][413],u_xpb_out[83][413],u_xpb_out[84][413],u_xpb_out[85][413],u_xpb_out[86][413],u_xpb_out[87][413],u_xpb_out[88][413],u_xpb_out[89][413],u_xpb_out[90][413],u_xpb_out[91][413],u_xpb_out[92][413],u_xpb_out[93][413],u_xpb_out[94][413],u_xpb_out[95][413],u_xpb_out[96][413],u_xpb_out[97][413],u_xpb_out[98][413],u_xpb_out[99][413],u_xpb_out[100][413],u_xpb_out[101][413],u_xpb_out[102][413],u_xpb_out[103][413],u_xpb_out[104][413],u_xpb_out[105][413]};

assign col_out_414 = {u_xpb_out[0][414],u_xpb_out[1][414],u_xpb_out[2][414],u_xpb_out[3][414],u_xpb_out[4][414],u_xpb_out[5][414],u_xpb_out[6][414],u_xpb_out[7][414],u_xpb_out[8][414],u_xpb_out[9][414],u_xpb_out[10][414],u_xpb_out[11][414],u_xpb_out[12][414],u_xpb_out[13][414],u_xpb_out[14][414],u_xpb_out[15][414],u_xpb_out[16][414],u_xpb_out[17][414],u_xpb_out[18][414],u_xpb_out[19][414],u_xpb_out[20][414],u_xpb_out[21][414],u_xpb_out[22][414],u_xpb_out[23][414],u_xpb_out[24][414],u_xpb_out[25][414],u_xpb_out[26][414],u_xpb_out[27][414],u_xpb_out[28][414],u_xpb_out[29][414],u_xpb_out[30][414],u_xpb_out[31][414],u_xpb_out[32][414],u_xpb_out[33][414],u_xpb_out[34][414],u_xpb_out[35][414],u_xpb_out[36][414],u_xpb_out[37][414],u_xpb_out[38][414],u_xpb_out[39][414],u_xpb_out[40][414],u_xpb_out[41][414],u_xpb_out[42][414],u_xpb_out[43][414],u_xpb_out[44][414],u_xpb_out[45][414],u_xpb_out[46][414],u_xpb_out[47][414],u_xpb_out[48][414],u_xpb_out[49][414],u_xpb_out[50][414],u_xpb_out[51][414],u_xpb_out[52][414],u_xpb_out[53][414],u_xpb_out[54][414],u_xpb_out[55][414],u_xpb_out[56][414],u_xpb_out[57][414],u_xpb_out[58][414],u_xpb_out[59][414],u_xpb_out[60][414],u_xpb_out[61][414],u_xpb_out[62][414],u_xpb_out[63][414],u_xpb_out[64][414],u_xpb_out[65][414],u_xpb_out[66][414],u_xpb_out[67][414],u_xpb_out[68][414],u_xpb_out[69][414],u_xpb_out[70][414],u_xpb_out[71][414],u_xpb_out[72][414],u_xpb_out[73][414],u_xpb_out[74][414],u_xpb_out[75][414],u_xpb_out[76][414],u_xpb_out[77][414],u_xpb_out[78][414],u_xpb_out[79][414],u_xpb_out[80][414],u_xpb_out[81][414],u_xpb_out[82][414],u_xpb_out[83][414],u_xpb_out[84][414],u_xpb_out[85][414],u_xpb_out[86][414],u_xpb_out[87][414],u_xpb_out[88][414],u_xpb_out[89][414],u_xpb_out[90][414],u_xpb_out[91][414],u_xpb_out[92][414],u_xpb_out[93][414],u_xpb_out[94][414],u_xpb_out[95][414],u_xpb_out[96][414],u_xpb_out[97][414],u_xpb_out[98][414],u_xpb_out[99][414],u_xpb_out[100][414],u_xpb_out[101][414],u_xpb_out[102][414],u_xpb_out[103][414],u_xpb_out[104][414],u_xpb_out[105][414]};

assign col_out_415 = {u_xpb_out[0][415],u_xpb_out[1][415],u_xpb_out[2][415],u_xpb_out[3][415],u_xpb_out[4][415],u_xpb_out[5][415],u_xpb_out[6][415],u_xpb_out[7][415],u_xpb_out[8][415],u_xpb_out[9][415],u_xpb_out[10][415],u_xpb_out[11][415],u_xpb_out[12][415],u_xpb_out[13][415],u_xpb_out[14][415],u_xpb_out[15][415],u_xpb_out[16][415],u_xpb_out[17][415],u_xpb_out[18][415],u_xpb_out[19][415],u_xpb_out[20][415],u_xpb_out[21][415],u_xpb_out[22][415],u_xpb_out[23][415],u_xpb_out[24][415],u_xpb_out[25][415],u_xpb_out[26][415],u_xpb_out[27][415],u_xpb_out[28][415],u_xpb_out[29][415],u_xpb_out[30][415],u_xpb_out[31][415],u_xpb_out[32][415],u_xpb_out[33][415],u_xpb_out[34][415],u_xpb_out[35][415],u_xpb_out[36][415],u_xpb_out[37][415],u_xpb_out[38][415],u_xpb_out[39][415],u_xpb_out[40][415],u_xpb_out[41][415],u_xpb_out[42][415],u_xpb_out[43][415],u_xpb_out[44][415],u_xpb_out[45][415],u_xpb_out[46][415],u_xpb_out[47][415],u_xpb_out[48][415],u_xpb_out[49][415],u_xpb_out[50][415],u_xpb_out[51][415],u_xpb_out[52][415],u_xpb_out[53][415],u_xpb_out[54][415],u_xpb_out[55][415],u_xpb_out[56][415],u_xpb_out[57][415],u_xpb_out[58][415],u_xpb_out[59][415],u_xpb_out[60][415],u_xpb_out[61][415],u_xpb_out[62][415],u_xpb_out[63][415],u_xpb_out[64][415],u_xpb_out[65][415],u_xpb_out[66][415],u_xpb_out[67][415],u_xpb_out[68][415],u_xpb_out[69][415],u_xpb_out[70][415],u_xpb_out[71][415],u_xpb_out[72][415],u_xpb_out[73][415],u_xpb_out[74][415],u_xpb_out[75][415],u_xpb_out[76][415],u_xpb_out[77][415],u_xpb_out[78][415],u_xpb_out[79][415],u_xpb_out[80][415],u_xpb_out[81][415],u_xpb_out[82][415],u_xpb_out[83][415],u_xpb_out[84][415],u_xpb_out[85][415],u_xpb_out[86][415],u_xpb_out[87][415],u_xpb_out[88][415],u_xpb_out[89][415],u_xpb_out[90][415],u_xpb_out[91][415],u_xpb_out[92][415],u_xpb_out[93][415],u_xpb_out[94][415],u_xpb_out[95][415],u_xpb_out[96][415],u_xpb_out[97][415],u_xpb_out[98][415],u_xpb_out[99][415],u_xpb_out[100][415],u_xpb_out[101][415],u_xpb_out[102][415],u_xpb_out[103][415],u_xpb_out[104][415],u_xpb_out[105][415]};

assign col_out_416 = {u_xpb_out[0][416],u_xpb_out[1][416],u_xpb_out[2][416],u_xpb_out[3][416],u_xpb_out[4][416],u_xpb_out[5][416],u_xpb_out[6][416],u_xpb_out[7][416],u_xpb_out[8][416],u_xpb_out[9][416],u_xpb_out[10][416],u_xpb_out[11][416],u_xpb_out[12][416],u_xpb_out[13][416],u_xpb_out[14][416],u_xpb_out[15][416],u_xpb_out[16][416],u_xpb_out[17][416],u_xpb_out[18][416],u_xpb_out[19][416],u_xpb_out[20][416],u_xpb_out[21][416],u_xpb_out[22][416],u_xpb_out[23][416],u_xpb_out[24][416],u_xpb_out[25][416],u_xpb_out[26][416],u_xpb_out[27][416],u_xpb_out[28][416],u_xpb_out[29][416],u_xpb_out[30][416],u_xpb_out[31][416],u_xpb_out[32][416],u_xpb_out[33][416],u_xpb_out[34][416],u_xpb_out[35][416],u_xpb_out[36][416],u_xpb_out[37][416],u_xpb_out[38][416],u_xpb_out[39][416],u_xpb_out[40][416],u_xpb_out[41][416],u_xpb_out[42][416],u_xpb_out[43][416],u_xpb_out[44][416],u_xpb_out[45][416],u_xpb_out[46][416],u_xpb_out[47][416],u_xpb_out[48][416],u_xpb_out[49][416],u_xpb_out[50][416],u_xpb_out[51][416],u_xpb_out[52][416],u_xpb_out[53][416],u_xpb_out[54][416],u_xpb_out[55][416],u_xpb_out[56][416],u_xpb_out[57][416],u_xpb_out[58][416],u_xpb_out[59][416],u_xpb_out[60][416],u_xpb_out[61][416],u_xpb_out[62][416],u_xpb_out[63][416],u_xpb_out[64][416],u_xpb_out[65][416],u_xpb_out[66][416],u_xpb_out[67][416],u_xpb_out[68][416],u_xpb_out[69][416],u_xpb_out[70][416],u_xpb_out[71][416],u_xpb_out[72][416],u_xpb_out[73][416],u_xpb_out[74][416],u_xpb_out[75][416],u_xpb_out[76][416],u_xpb_out[77][416],u_xpb_out[78][416],u_xpb_out[79][416],u_xpb_out[80][416],u_xpb_out[81][416],u_xpb_out[82][416],u_xpb_out[83][416],u_xpb_out[84][416],u_xpb_out[85][416],u_xpb_out[86][416],u_xpb_out[87][416],u_xpb_out[88][416],u_xpb_out[89][416],u_xpb_out[90][416],u_xpb_out[91][416],u_xpb_out[92][416],u_xpb_out[93][416],u_xpb_out[94][416],u_xpb_out[95][416],u_xpb_out[96][416],u_xpb_out[97][416],u_xpb_out[98][416],u_xpb_out[99][416],u_xpb_out[100][416],u_xpb_out[101][416],u_xpb_out[102][416],u_xpb_out[103][416],u_xpb_out[104][416],u_xpb_out[105][416]};

assign col_out_417 = {u_xpb_out[0][417],u_xpb_out[1][417],u_xpb_out[2][417],u_xpb_out[3][417],u_xpb_out[4][417],u_xpb_out[5][417],u_xpb_out[6][417],u_xpb_out[7][417],u_xpb_out[8][417],u_xpb_out[9][417],u_xpb_out[10][417],u_xpb_out[11][417],u_xpb_out[12][417],u_xpb_out[13][417],u_xpb_out[14][417],u_xpb_out[15][417],u_xpb_out[16][417],u_xpb_out[17][417],u_xpb_out[18][417],u_xpb_out[19][417],u_xpb_out[20][417],u_xpb_out[21][417],u_xpb_out[22][417],u_xpb_out[23][417],u_xpb_out[24][417],u_xpb_out[25][417],u_xpb_out[26][417],u_xpb_out[27][417],u_xpb_out[28][417],u_xpb_out[29][417],u_xpb_out[30][417],u_xpb_out[31][417],u_xpb_out[32][417],u_xpb_out[33][417],u_xpb_out[34][417],u_xpb_out[35][417],u_xpb_out[36][417],u_xpb_out[37][417],u_xpb_out[38][417],u_xpb_out[39][417],u_xpb_out[40][417],u_xpb_out[41][417],u_xpb_out[42][417],u_xpb_out[43][417],u_xpb_out[44][417],u_xpb_out[45][417],u_xpb_out[46][417],u_xpb_out[47][417],u_xpb_out[48][417],u_xpb_out[49][417],u_xpb_out[50][417],u_xpb_out[51][417],u_xpb_out[52][417],u_xpb_out[53][417],u_xpb_out[54][417],u_xpb_out[55][417],u_xpb_out[56][417],u_xpb_out[57][417],u_xpb_out[58][417],u_xpb_out[59][417],u_xpb_out[60][417],u_xpb_out[61][417],u_xpb_out[62][417],u_xpb_out[63][417],u_xpb_out[64][417],u_xpb_out[65][417],u_xpb_out[66][417],u_xpb_out[67][417],u_xpb_out[68][417],u_xpb_out[69][417],u_xpb_out[70][417],u_xpb_out[71][417],u_xpb_out[72][417],u_xpb_out[73][417],u_xpb_out[74][417],u_xpb_out[75][417],u_xpb_out[76][417],u_xpb_out[77][417],u_xpb_out[78][417],u_xpb_out[79][417],u_xpb_out[80][417],u_xpb_out[81][417],u_xpb_out[82][417],u_xpb_out[83][417],u_xpb_out[84][417],u_xpb_out[85][417],u_xpb_out[86][417],u_xpb_out[87][417],u_xpb_out[88][417],u_xpb_out[89][417],u_xpb_out[90][417],u_xpb_out[91][417],u_xpb_out[92][417],u_xpb_out[93][417],u_xpb_out[94][417],u_xpb_out[95][417],u_xpb_out[96][417],u_xpb_out[97][417],u_xpb_out[98][417],u_xpb_out[99][417],u_xpb_out[100][417],u_xpb_out[101][417],u_xpb_out[102][417],u_xpb_out[103][417],u_xpb_out[104][417],u_xpb_out[105][417]};

assign col_out_418 = {u_xpb_out[0][418],u_xpb_out[1][418],u_xpb_out[2][418],u_xpb_out[3][418],u_xpb_out[4][418],u_xpb_out[5][418],u_xpb_out[6][418],u_xpb_out[7][418],u_xpb_out[8][418],u_xpb_out[9][418],u_xpb_out[10][418],u_xpb_out[11][418],u_xpb_out[12][418],u_xpb_out[13][418],u_xpb_out[14][418],u_xpb_out[15][418],u_xpb_out[16][418],u_xpb_out[17][418],u_xpb_out[18][418],u_xpb_out[19][418],u_xpb_out[20][418],u_xpb_out[21][418],u_xpb_out[22][418],u_xpb_out[23][418],u_xpb_out[24][418],u_xpb_out[25][418],u_xpb_out[26][418],u_xpb_out[27][418],u_xpb_out[28][418],u_xpb_out[29][418],u_xpb_out[30][418],u_xpb_out[31][418],u_xpb_out[32][418],u_xpb_out[33][418],u_xpb_out[34][418],u_xpb_out[35][418],u_xpb_out[36][418],u_xpb_out[37][418],u_xpb_out[38][418],u_xpb_out[39][418],u_xpb_out[40][418],u_xpb_out[41][418],u_xpb_out[42][418],u_xpb_out[43][418],u_xpb_out[44][418],u_xpb_out[45][418],u_xpb_out[46][418],u_xpb_out[47][418],u_xpb_out[48][418],u_xpb_out[49][418],u_xpb_out[50][418],u_xpb_out[51][418],u_xpb_out[52][418],u_xpb_out[53][418],u_xpb_out[54][418],u_xpb_out[55][418],u_xpb_out[56][418],u_xpb_out[57][418],u_xpb_out[58][418],u_xpb_out[59][418],u_xpb_out[60][418],u_xpb_out[61][418],u_xpb_out[62][418],u_xpb_out[63][418],u_xpb_out[64][418],u_xpb_out[65][418],u_xpb_out[66][418],u_xpb_out[67][418],u_xpb_out[68][418],u_xpb_out[69][418],u_xpb_out[70][418],u_xpb_out[71][418],u_xpb_out[72][418],u_xpb_out[73][418],u_xpb_out[74][418],u_xpb_out[75][418],u_xpb_out[76][418],u_xpb_out[77][418],u_xpb_out[78][418],u_xpb_out[79][418],u_xpb_out[80][418],u_xpb_out[81][418],u_xpb_out[82][418],u_xpb_out[83][418],u_xpb_out[84][418],u_xpb_out[85][418],u_xpb_out[86][418],u_xpb_out[87][418],u_xpb_out[88][418],u_xpb_out[89][418],u_xpb_out[90][418],u_xpb_out[91][418],u_xpb_out[92][418],u_xpb_out[93][418],u_xpb_out[94][418],u_xpb_out[95][418],u_xpb_out[96][418],u_xpb_out[97][418],u_xpb_out[98][418],u_xpb_out[99][418],u_xpb_out[100][418],u_xpb_out[101][418],u_xpb_out[102][418],u_xpb_out[103][418],u_xpb_out[104][418],u_xpb_out[105][418]};

assign col_out_419 = {u_xpb_out[0][419],u_xpb_out[1][419],u_xpb_out[2][419],u_xpb_out[3][419],u_xpb_out[4][419],u_xpb_out[5][419],u_xpb_out[6][419],u_xpb_out[7][419],u_xpb_out[8][419],u_xpb_out[9][419],u_xpb_out[10][419],u_xpb_out[11][419],u_xpb_out[12][419],u_xpb_out[13][419],u_xpb_out[14][419],u_xpb_out[15][419],u_xpb_out[16][419],u_xpb_out[17][419],u_xpb_out[18][419],u_xpb_out[19][419],u_xpb_out[20][419],u_xpb_out[21][419],u_xpb_out[22][419],u_xpb_out[23][419],u_xpb_out[24][419],u_xpb_out[25][419],u_xpb_out[26][419],u_xpb_out[27][419],u_xpb_out[28][419],u_xpb_out[29][419],u_xpb_out[30][419],u_xpb_out[31][419],u_xpb_out[32][419],u_xpb_out[33][419],u_xpb_out[34][419],u_xpb_out[35][419],u_xpb_out[36][419],u_xpb_out[37][419],u_xpb_out[38][419],u_xpb_out[39][419],u_xpb_out[40][419],u_xpb_out[41][419],u_xpb_out[42][419],u_xpb_out[43][419],u_xpb_out[44][419],u_xpb_out[45][419],u_xpb_out[46][419],u_xpb_out[47][419],u_xpb_out[48][419],u_xpb_out[49][419],u_xpb_out[50][419],u_xpb_out[51][419],u_xpb_out[52][419],u_xpb_out[53][419],u_xpb_out[54][419],u_xpb_out[55][419],u_xpb_out[56][419],u_xpb_out[57][419],u_xpb_out[58][419],u_xpb_out[59][419],u_xpb_out[60][419],u_xpb_out[61][419],u_xpb_out[62][419],u_xpb_out[63][419],u_xpb_out[64][419],u_xpb_out[65][419],u_xpb_out[66][419],u_xpb_out[67][419],u_xpb_out[68][419],u_xpb_out[69][419],u_xpb_out[70][419],u_xpb_out[71][419],u_xpb_out[72][419],u_xpb_out[73][419],u_xpb_out[74][419],u_xpb_out[75][419],u_xpb_out[76][419],u_xpb_out[77][419],u_xpb_out[78][419],u_xpb_out[79][419],u_xpb_out[80][419],u_xpb_out[81][419],u_xpb_out[82][419],u_xpb_out[83][419],u_xpb_out[84][419],u_xpb_out[85][419],u_xpb_out[86][419],u_xpb_out[87][419],u_xpb_out[88][419],u_xpb_out[89][419],u_xpb_out[90][419],u_xpb_out[91][419],u_xpb_out[92][419],u_xpb_out[93][419],u_xpb_out[94][419],u_xpb_out[95][419],u_xpb_out[96][419],u_xpb_out[97][419],u_xpb_out[98][419],u_xpb_out[99][419],u_xpb_out[100][419],u_xpb_out[101][419],u_xpb_out[102][419],u_xpb_out[103][419],u_xpb_out[104][419],u_xpb_out[105][419]};

assign col_out_420 = {u_xpb_out[0][420],u_xpb_out[1][420],u_xpb_out[2][420],u_xpb_out[3][420],u_xpb_out[4][420],u_xpb_out[5][420],u_xpb_out[6][420],u_xpb_out[7][420],u_xpb_out[8][420],u_xpb_out[9][420],u_xpb_out[10][420],u_xpb_out[11][420],u_xpb_out[12][420],u_xpb_out[13][420],u_xpb_out[14][420],u_xpb_out[15][420],u_xpb_out[16][420],u_xpb_out[17][420],u_xpb_out[18][420],u_xpb_out[19][420],u_xpb_out[20][420],u_xpb_out[21][420],u_xpb_out[22][420],u_xpb_out[23][420],u_xpb_out[24][420],u_xpb_out[25][420],u_xpb_out[26][420],u_xpb_out[27][420],u_xpb_out[28][420],u_xpb_out[29][420],u_xpb_out[30][420],u_xpb_out[31][420],u_xpb_out[32][420],u_xpb_out[33][420],u_xpb_out[34][420],u_xpb_out[35][420],u_xpb_out[36][420],u_xpb_out[37][420],u_xpb_out[38][420],u_xpb_out[39][420],u_xpb_out[40][420],u_xpb_out[41][420],u_xpb_out[42][420],u_xpb_out[43][420],u_xpb_out[44][420],u_xpb_out[45][420],u_xpb_out[46][420],u_xpb_out[47][420],u_xpb_out[48][420],u_xpb_out[49][420],u_xpb_out[50][420],u_xpb_out[51][420],u_xpb_out[52][420],u_xpb_out[53][420],u_xpb_out[54][420],u_xpb_out[55][420],u_xpb_out[56][420],u_xpb_out[57][420],u_xpb_out[58][420],u_xpb_out[59][420],u_xpb_out[60][420],u_xpb_out[61][420],u_xpb_out[62][420],u_xpb_out[63][420],u_xpb_out[64][420],u_xpb_out[65][420],u_xpb_out[66][420],u_xpb_out[67][420],u_xpb_out[68][420],u_xpb_out[69][420],u_xpb_out[70][420],u_xpb_out[71][420],u_xpb_out[72][420],u_xpb_out[73][420],u_xpb_out[74][420],u_xpb_out[75][420],u_xpb_out[76][420],u_xpb_out[77][420],u_xpb_out[78][420],u_xpb_out[79][420],u_xpb_out[80][420],u_xpb_out[81][420],u_xpb_out[82][420],u_xpb_out[83][420],u_xpb_out[84][420],u_xpb_out[85][420],u_xpb_out[86][420],u_xpb_out[87][420],u_xpb_out[88][420],u_xpb_out[89][420],u_xpb_out[90][420],u_xpb_out[91][420],u_xpb_out[92][420],u_xpb_out[93][420],u_xpb_out[94][420],u_xpb_out[95][420],u_xpb_out[96][420],u_xpb_out[97][420],u_xpb_out[98][420],u_xpb_out[99][420],u_xpb_out[100][420],u_xpb_out[101][420],u_xpb_out[102][420],u_xpb_out[103][420],u_xpb_out[104][420],u_xpb_out[105][420]};

assign col_out_421 = {u_xpb_out[0][421],u_xpb_out[1][421],u_xpb_out[2][421],u_xpb_out[3][421],u_xpb_out[4][421],u_xpb_out[5][421],u_xpb_out[6][421],u_xpb_out[7][421],u_xpb_out[8][421],u_xpb_out[9][421],u_xpb_out[10][421],u_xpb_out[11][421],u_xpb_out[12][421],u_xpb_out[13][421],u_xpb_out[14][421],u_xpb_out[15][421],u_xpb_out[16][421],u_xpb_out[17][421],u_xpb_out[18][421],u_xpb_out[19][421],u_xpb_out[20][421],u_xpb_out[21][421],u_xpb_out[22][421],u_xpb_out[23][421],u_xpb_out[24][421],u_xpb_out[25][421],u_xpb_out[26][421],u_xpb_out[27][421],u_xpb_out[28][421],u_xpb_out[29][421],u_xpb_out[30][421],u_xpb_out[31][421],u_xpb_out[32][421],u_xpb_out[33][421],u_xpb_out[34][421],u_xpb_out[35][421],u_xpb_out[36][421],u_xpb_out[37][421],u_xpb_out[38][421],u_xpb_out[39][421],u_xpb_out[40][421],u_xpb_out[41][421],u_xpb_out[42][421],u_xpb_out[43][421],u_xpb_out[44][421],u_xpb_out[45][421],u_xpb_out[46][421],u_xpb_out[47][421],u_xpb_out[48][421],u_xpb_out[49][421],u_xpb_out[50][421],u_xpb_out[51][421],u_xpb_out[52][421],u_xpb_out[53][421],u_xpb_out[54][421],u_xpb_out[55][421],u_xpb_out[56][421],u_xpb_out[57][421],u_xpb_out[58][421],u_xpb_out[59][421],u_xpb_out[60][421],u_xpb_out[61][421],u_xpb_out[62][421],u_xpb_out[63][421],u_xpb_out[64][421],u_xpb_out[65][421],u_xpb_out[66][421],u_xpb_out[67][421],u_xpb_out[68][421],u_xpb_out[69][421],u_xpb_out[70][421],u_xpb_out[71][421],u_xpb_out[72][421],u_xpb_out[73][421],u_xpb_out[74][421],u_xpb_out[75][421],u_xpb_out[76][421],u_xpb_out[77][421],u_xpb_out[78][421],u_xpb_out[79][421],u_xpb_out[80][421],u_xpb_out[81][421],u_xpb_out[82][421],u_xpb_out[83][421],u_xpb_out[84][421],u_xpb_out[85][421],u_xpb_out[86][421],u_xpb_out[87][421],u_xpb_out[88][421],u_xpb_out[89][421],u_xpb_out[90][421],u_xpb_out[91][421],u_xpb_out[92][421],u_xpb_out[93][421],u_xpb_out[94][421],u_xpb_out[95][421],u_xpb_out[96][421],u_xpb_out[97][421],u_xpb_out[98][421],u_xpb_out[99][421],u_xpb_out[100][421],u_xpb_out[101][421],u_xpb_out[102][421],u_xpb_out[103][421],u_xpb_out[104][421],u_xpb_out[105][421]};

assign col_out_422 = {u_xpb_out[0][422],u_xpb_out[1][422],u_xpb_out[2][422],u_xpb_out[3][422],u_xpb_out[4][422],u_xpb_out[5][422],u_xpb_out[6][422],u_xpb_out[7][422],u_xpb_out[8][422],u_xpb_out[9][422],u_xpb_out[10][422],u_xpb_out[11][422],u_xpb_out[12][422],u_xpb_out[13][422],u_xpb_out[14][422],u_xpb_out[15][422],u_xpb_out[16][422],u_xpb_out[17][422],u_xpb_out[18][422],u_xpb_out[19][422],u_xpb_out[20][422],u_xpb_out[21][422],u_xpb_out[22][422],u_xpb_out[23][422],u_xpb_out[24][422],u_xpb_out[25][422],u_xpb_out[26][422],u_xpb_out[27][422],u_xpb_out[28][422],u_xpb_out[29][422],u_xpb_out[30][422],u_xpb_out[31][422],u_xpb_out[32][422],u_xpb_out[33][422],u_xpb_out[34][422],u_xpb_out[35][422],u_xpb_out[36][422],u_xpb_out[37][422],u_xpb_out[38][422],u_xpb_out[39][422],u_xpb_out[40][422],u_xpb_out[41][422],u_xpb_out[42][422],u_xpb_out[43][422],u_xpb_out[44][422],u_xpb_out[45][422],u_xpb_out[46][422],u_xpb_out[47][422],u_xpb_out[48][422],u_xpb_out[49][422],u_xpb_out[50][422],u_xpb_out[51][422],u_xpb_out[52][422],u_xpb_out[53][422],u_xpb_out[54][422],u_xpb_out[55][422],u_xpb_out[56][422],u_xpb_out[57][422],u_xpb_out[58][422],u_xpb_out[59][422],u_xpb_out[60][422],u_xpb_out[61][422],u_xpb_out[62][422],u_xpb_out[63][422],u_xpb_out[64][422],u_xpb_out[65][422],u_xpb_out[66][422],u_xpb_out[67][422],u_xpb_out[68][422],u_xpb_out[69][422],u_xpb_out[70][422],u_xpb_out[71][422],u_xpb_out[72][422],u_xpb_out[73][422],u_xpb_out[74][422],u_xpb_out[75][422],u_xpb_out[76][422],u_xpb_out[77][422],u_xpb_out[78][422],u_xpb_out[79][422],u_xpb_out[80][422],u_xpb_out[81][422],u_xpb_out[82][422],u_xpb_out[83][422],u_xpb_out[84][422],u_xpb_out[85][422],u_xpb_out[86][422],u_xpb_out[87][422],u_xpb_out[88][422],u_xpb_out[89][422],u_xpb_out[90][422],u_xpb_out[91][422],u_xpb_out[92][422],u_xpb_out[93][422],u_xpb_out[94][422],u_xpb_out[95][422],u_xpb_out[96][422],u_xpb_out[97][422],u_xpb_out[98][422],u_xpb_out[99][422],u_xpb_out[100][422],u_xpb_out[101][422],u_xpb_out[102][422],u_xpb_out[103][422],u_xpb_out[104][422],u_xpb_out[105][422]};

assign col_out_423 = {u_xpb_out[0][423],u_xpb_out[1][423],u_xpb_out[2][423],u_xpb_out[3][423],u_xpb_out[4][423],u_xpb_out[5][423],u_xpb_out[6][423],u_xpb_out[7][423],u_xpb_out[8][423],u_xpb_out[9][423],u_xpb_out[10][423],u_xpb_out[11][423],u_xpb_out[12][423],u_xpb_out[13][423],u_xpb_out[14][423],u_xpb_out[15][423],u_xpb_out[16][423],u_xpb_out[17][423],u_xpb_out[18][423],u_xpb_out[19][423],u_xpb_out[20][423],u_xpb_out[21][423],u_xpb_out[22][423],u_xpb_out[23][423],u_xpb_out[24][423],u_xpb_out[25][423],u_xpb_out[26][423],u_xpb_out[27][423],u_xpb_out[28][423],u_xpb_out[29][423],u_xpb_out[30][423],u_xpb_out[31][423],u_xpb_out[32][423],u_xpb_out[33][423],u_xpb_out[34][423],u_xpb_out[35][423],u_xpb_out[36][423],u_xpb_out[37][423],u_xpb_out[38][423],u_xpb_out[39][423],u_xpb_out[40][423],u_xpb_out[41][423],u_xpb_out[42][423],u_xpb_out[43][423],u_xpb_out[44][423],u_xpb_out[45][423],u_xpb_out[46][423],u_xpb_out[47][423],u_xpb_out[48][423],u_xpb_out[49][423],u_xpb_out[50][423],u_xpb_out[51][423],u_xpb_out[52][423],u_xpb_out[53][423],u_xpb_out[54][423],u_xpb_out[55][423],u_xpb_out[56][423],u_xpb_out[57][423],u_xpb_out[58][423],u_xpb_out[59][423],u_xpb_out[60][423],u_xpb_out[61][423],u_xpb_out[62][423],u_xpb_out[63][423],u_xpb_out[64][423],u_xpb_out[65][423],u_xpb_out[66][423],u_xpb_out[67][423],u_xpb_out[68][423],u_xpb_out[69][423],u_xpb_out[70][423],u_xpb_out[71][423],u_xpb_out[72][423],u_xpb_out[73][423],u_xpb_out[74][423],u_xpb_out[75][423],u_xpb_out[76][423],u_xpb_out[77][423],u_xpb_out[78][423],u_xpb_out[79][423],u_xpb_out[80][423],u_xpb_out[81][423],u_xpb_out[82][423],u_xpb_out[83][423],u_xpb_out[84][423],u_xpb_out[85][423],u_xpb_out[86][423],u_xpb_out[87][423],u_xpb_out[88][423],u_xpb_out[89][423],u_xpb_out[90][423],u_xpb_out[91][423],u_xpb_out[92][423],u_xpb_out[93][423],u_xpb_out[94][423],u_xpb_out[95][423],u_xpb_out[96][423],u_xpb_out[97][423],u_xpb_out[98][423],u_xpb_out[99][423],u_xpb_out[100][423],u_xpb_out[101][423],u_xpb_out[102][423],u_xpb_out[103][423],u_xpb_out[104][423],u_xpb_out[105][423]};

assign col_out_424 = {u_xpb_out[0][424],u_xpb_out[1][424],u_xpb_out[2][424],u_xpb_out[3][424],u_xpb_out[4][424],u_xpb_out[5][424],u_xpb_out[6][424],u_xpb_out[7][424],u_xpb_out[8][424],u_xpb_out[9][424],u_xpb_out[10][424],u_xpb_out[11][424],u_xpb_out[12][424],u_xpb_out[13][424],u_xpb_out[14][424],u_xpb_out[15][424],u_xpb_out[16][424],u_xpb_out[17][424],u_xpb_out[18][424],u_xpb_out[19][424],u_xpb_out[20][424],u_xpb_out[21][424],u_xpb_out[22][424],u_xpb_out[23][424],u_xpb_out[24][424],u_xpb_out[25][424],u_xpb_out[26][424],u_xpb_out[27][424],u_xpb_out[28][424],u_xpb_out[29][424],u_xpb_out[30][424],u_xpb_out[31][424],u_xpb_out[32][424],u_xpb_out[33][424],u_xpb_out[34][424],u_xpb_out[35][424],u_xpb_out[36][424],u_xpb_out[37][424],u_xpb_out[38][424],u_xpb_out[39][424],u_xpb_out[40][424],u_xpb_out[41][424],u_xpb_out[42][424],u_xpb_out[43][424],u_xpb_out[44][424],u_xpb_out[45][424],u_xpb_out[46][424],u_xpb_out[47][424],u_xpb_out[48][424],u_xpb_out[49][424],u_xpb_out[50][424],u_xpb_out[51][424],u_xpb_out[52][424],u_xpb_out[53][424],u_xpb_out[54][424],u_xpb_out[55][424],u_xpb_out[56][424],u_xpb_out[57][424],u_xpb_out[58][424],u_xpb_out[59][424],u_xpb_out[60][424],u_xpb_out[61][424],u_xpb_out[62][424],u_xpb_out[63][424],u_xpb_out[64][424],u_xpb_out[65][424],u_xpb_out[66][424],u_xpb_out[67][424],u_xpb_out[68][424],u_xpb_out[69][424],u_xpb_out[70][424],u_xpb_out[71][424],u_xpb_out[72][424],u_xpb_out[73][424],u_xpb_out[74][424],u_xpb_out[75][424],u_xpb_out[76][424],u_xpb_out[77][424],u_xpb_out[78][424],u_xpb_out[79][424],u_xpb_out[80][424],u_xpb_out[81][424],u_xpb_out[82][424],u_xpb_out[83][424],u_xpb_out[84][424],u_xpb_out[85][424],u_xpb_out[86][424],u_xpb_out[87][424],u_xpb_out[88][424],u_xpb_out[89][424],u_xpb_out[90][424],u_xpb_out[91][424],u_xpb_out[92][424],u_xpb_out[93][424],u_xpb_out[94][424],u_xpb_out[95][424],u_xpb_out[96][424],u_xpb_out[97][424],u_xpb_out[98][424],u_xpb_out[99][424],u_xpb_out[100][424],u_xpb_out[101][424],u_xpb_out[102][424],u_xpb_out[103][424],u_xpb_out[104][424],u_xpb_out[105][424]};

assign col_out_425 = {u_xpb_out[0][425],u_xpb_out[1][425],u_xpb_out[2][425],u_xpb_out[3][425],u_xpb_out[4][425],u_xpb_out[5][425],u_xpb_out[6][425],u_xpb_out[7][425],u_xpb_out[8][425],u_xpb_out[9][425],u_xpb_out[10][425],u_xpb_out[11][425],u_xpb_out[12][425],u_xpb_out[13][425],u_xpb_out[14][425],u_xpb_out[15][425],u_xpb_out[16][425],u_xpb_out[17][425],u_xpb_out[18][425],u_xpb_out[19][425],u_xpb_out[20][425],u_xpb_out[21][425],u_xpb_out[22][425],u_xpb_out[23][425],u_xpb_out[24][425],u_xpb_out[25][425],u_xpb_out[26][425],u_xpb_out[27][425],u_xpb_out[28][425],u_xpb_out[29][425],u_xpb_out[30][425],u_xpb_out[31][425],u_xpb_out[32][425],u_xpb_out[33][425],u_xpb_out[34][425],u_xpb_out[35][425],u_xpb_out[36][425],u_xpb_out[37][425],u_xpb_out[38][425],u_xpb_out[39][425],u_xpb_out[40][425],u_xpb_out[41][425],u_xpb_out[42][425],u_xpb_out[43][425],u_xpb_out[44][425],u_xpb_out[45][425],u_xpb_out[46][425],u_xpb_out[47][425],u_xpb_out[48][425],u_xpb_out[49][425],u_xpb_out[50][425],u_xpb_out[51][425],u_xpb_out[52][425],u_xpb_out[53][425],u_xpb_out[54][425],u_xpb_out[55][425],u_xpb_out[56][425],u_xpb_out[57][425],u_xpb_out[58][425],u_xpb_out[59][425],u_xpb_out[60][425],u_xpb_out[61][425],u_xpb_out[62][425],u_xpb_out[63][425],u_xpb_out[64][425],u_xpb_out[65][425],u_xpb_out[66][425],u_xpb_out[67][425],u_xpb_out[68][425],u_xpb_out[69][425],u_xpb_out[70][425],u_xpb_out[71][425],u_xpb_out[72][425],u_xpb_out[73][425],u_xpb_out[74][425],u_xpb_out[75][425],u_xpb_out[76][425],u_xpb_out[77][425],u_xpb_out[78][425],u_xpb_out[79][425],u_xpb_out[80][425],u_xpb_out[81][425],u_xpb_out[82][425],u_xpb_out[83][425],u_xpb_out[84][425],u_xpb_out[85][425],u_xpb_out[86][425],u_xpb_out[87][425],u_xpb_out[88][425],u_xpb_out[89][425],u_xpb_out[90][425],u_xpb_out[91][425],u_xpb_out[92][425],u_xpb_out[93][425],u_xpb_out[94][425],u_xpb_out[95][425],u_xpb_out[96][425],u_xpb_out[97][425],u_xpb_out[98][425],u_xpb_out[99][425],u_xpb_out[100][425],u_xpb_out[101][425],u_xpb_out[102][425],u_xpb_out[103][425],u_xpb_out[104][425],u_xpb_out[105][425]};

assign col_out_426 = {u_xpb_out[0][426],u_xpb_out[1][426],u_xpb_out[2][426],u_xpb_out[3][426],u_xpb_out[4][426],u_xpb_out[5][426],u_xpb_out[6][426],u_xpb_out[7][426],u_xpb_out[8][426],u_xpb_out[9][426],u_xpb_out[10][426],u_xpb_out[11][426],u_xpb_out[12][426],u_xpb_out[13][426],u_xpb_out[14][426],u_xpb_out[15][426],u_xpb_out[16][426],u_xpb_out[17][426],u_xpb_out[18][426],u_xpb_out[19][426],u_xpb_out[20][426],u_xpb_out[21][426],u_xpb_out[22][426],u_xpb_out[23][426],u_xpb_out[24][426],u_xpb_out[25][426],u_xpb_out[26][426],u_xpb_out[27][426],u_xpb_out[28][426],u_xpb_out[29][426],u_xpb_out[30][426],u_xpb_out[31][426],u_xpb_out[32][426],u_xpb_out[33][426],u_xpb_out[34][426],u_xpb_out[35][426],u_xpb_out[36][426],u_xpb_out[37][426],u_xpb_out[38][426],u_xpb_out[39][426],u_xpb_out[40][426],u_xpb_out[41][426],u_xpb_out[42][426],u_xpb_out[43][426],u_xpb_out[44][426],u_xpb_out[45][426],u_xpb_out[46][426],u_xpb_out[47][426],u_xpb_out[48][426],u_xpb_out[49][426],u_xpb_out[50][426],u_xpb_out[51][426],u_xpb_out[52][426],u_xpb_out[53][426],u_xpb_out[54][426],u_xpb_out[55][426],u_xpb_out[56][426],u_xpb_out[57][426],u_xpb_out[58][426],u_xpb_out[59][426],u_xpb_out[60][426],u_xpb_out[61][426],u_xpb_out[62][426],u_xpb_out[63][426],u_xpb_out[64][426],u_xpb_out[65][426],u_xpb_out[66][426],u_xpb_out[67][426],u_xpb_out[68][426],u_xpb_out[69][426],u_xpb_out[70][426],u_xpb_out[71][426],u_xpb_out[72][426],u_xpb_out[73][426],u_xpb_out[74][426],u_xpb_out[75][426],u_xpb_out[76][426],u_xpb_out[77][426],u_xpb_out[78][426],u_xpb_out[79][426],u_xpb_out[80][426],u_xpb_out[81][426],u_xpb_out[82][426],u_xpb_out[83][426],u_xpb_out[84][426],u_xpb_out[85][426],u_xpb_out[86][426],u_xpb_out[87][426],u_xpb_out[88][426],u_xpb_out[89][426],u_xpb_out[90][426],u_xpb_out[91][426],u_xpb_out[92][426],u_xpb_out[93][426],u_xpb_out[94][426],u_xpb_out[95][426],u_xpb_out[96][426],u_xpb_out[97][426],u_xpb_out[98][426],u_xpb_out[99][426],u_xpb_out[100][426],u_xpb_out[101][426],u_xpb_out[102][426],u_xpb_out[103][426],u_xpb_out[104][426],u_xpb_out[105][426]};

assign col_out_427 = {u_xpb_out[0][427],u_xpb_out[1][427],u_xpb_out[2][427],u_xpb_out[3][427],u_xpb_out[4][427],u_xpb_out[5][427],u_xpb_out[6][427],u_xpb_out[7][427],u_xpb_out[8][427],u_xpb_out[9][427],u_xpb_out[10][427],u_xpb_out[11][427],u_xpb_out[12][427],u_xpb_out[13][427],u_xpb_out[14][427],u_xpb_out[15][427],u_xpb_out[16][427],u_xpb_out[17][427],u_xpb_out[18][427],u_xpb_out[19][427],u_xpb_out[20][427],u_xpb_out[21][427],u_xpb_out[22][427],u_xpb_out[23][427],u_xpb_out[24][427],u_xpb_out[25][427],u_xpb_out[26][427],u_xpb_out[27][427],u_xpb_out[28][427],u_xpb_out[29][427],u_xpb_out[30][427],u_xpb_out[31][427],u_xpb_out[32][427],u_xpb_out[33][427],u_xpb_out[34][427],u_xpb_out[35][427],u_xpb_out[36][427],u_xpb_out[37][427],u_xpb_out[38][427],u_xpb_out[39][427],u_xpb_out[40][427],u_xpb_out[41][427],u_xpb_out[42][427],u_xpb_out[43][427],u_xpb_out[44][427],u_xpb_out[45][427],u_xpb_out[46][427],u_xpb_out[47][427],u_xpb_out[48][427],u_xpb_out[49][427],u_xpb_out[50][427],u_xpb_out[51][427],u_xpb_out[52][427],u_xpb_out[53][427],u_xpb_out[54][427],u_xpb_out[55][427],u_xpb_out[56][427],u_xpb_out[57][427],u_xpb_out[58][427],u_xpb_out[59][427],u_xpb_out[60][427],u_xpb_out[61][427],u_xpb_out[62][427],u_xpb_out[63][427],u_xpb_out[64][427],u_xpb_out[65][427],u_xpb_out[66][427],u_xpb_out[67][427],u_xpb_out[68][427],u_xpb_out[69][427],u_xpb_out[70][427],u_xpb_out[71][427],u_xpb_out[72][427],u_xpb_out[73][427],u_xpb_out[74][427],u_xpb_out[75][427],u_xpb_out[76][427],u_xpb_out[77][427],u_xpb_out[78][427],u_xpb_out[79][427],u_xpb_out[80][427],u_xpb_out[81][427],u_xpb_out[82][427],u_xpb_out[83][427],u_xpb_out[84][427],u_xpb_out[85][427],u_xpb_out[86][427],u_xpb_out[87][427],u_xpb_out[88][427],u_xpb_out[89][427],u_xpb_out[90][427],u_xpb_out[91][427],u_xpb_out[92][427],u_xpb_out[93][427],u_xpb_out[94][427],u_xpb_out[95][427],u_xpb_out[96][427],u_xpb_out[97][427],u_xpb_out[98][427],u_xpb_out[99][427],u_xpb_out[100][427],u_xpb_out[101][427],u_xpb_out[102][427],u_xpb_out[103][427],u_xpb_out[104][427],u_xpb_out[105][427]};

assign col_out_428 = {u_xpb_out[0][428],u_xpb_out[1][428],u_xpb_out[2][428],u_xpb_out[3][428],u_xpb_out[4][428],u_xpb_out[5][428],u_xpb_out[6][428],u_xpb_out[7][428],u_xpb_out[8][428],u_xpb_out[9][428],u_xpb_out[10][428],u_xpb_out[11][428],u_xpb_out[12][428],u_xpb_out[13][428],u_xpb_out[14][428],u_xpb_out[15][428],u_xpb_out[16][428],u_xpb_out[17][428],u_xpb_out[18][428],u_xpb_out[19][428],u_xpb_out[20][428],u_xpb_out[21][428],u_xpb_out[22][428],u_xpb_out[23][428],u_xpb_out[24][428],u_xpb_out[25][428],u_xpb_out[26][428],u_xpb_out[27][428],u_xpb_out[28][428],u_xpb_out[29][428],u_xpb_out[30][428],u_xpb_out[31][428],u_xpb_out[32][428],u_xpb_out[33][428],u_xpb_out[34][428],u_xpb_out[35][428],u_xpb_out[36][428],u_xpb_out[37][428],u_xpb_out[38][428],u_xpb_out[39][428],u_xpb_out[40][428],u_xpb_out[41][428],u_xpb_out[42][428],u_xpb_out[43][428],u_xpb_out[44][428],u_xpb_out[45][428],u_xpb_out[46][428],u_xpb_out[47][428],u_xpb_out[48][428],u_xpb_out[49][428],u_xpb_out[50][428],u_xpb_out[51][428],u_xpb_out[52][428],u_xpb_out[53][428],u_xpb_out[54][428],u_xpb_out[55][428],u_xpb_out[56][428],u_xpb_out[57][428],u_xpb_out[58][428],u_xpb_out[59][428],u_xpb_out[60][428],u_xpb_out[61][428],u_xpb_out[62][428],u_xpb_out[63][428],u_xpb_out[64][428],u_xpb_out[65][428],u_xpb_out[66][428],u_xpb_out[67][428],u_xpb_out[68][428],u_xpb_out[69][428],u_xpb_out[70][428],u_xpb_out[71][428],u_xpb_out[72][428],u_xpb_out[73][428],u_xpb_out[74][428],u_xpb_out[75][428],u_xpb_out[76][428],u_xpb_out[77][428],u_xpb_out[78][428],u_xpb_out[79][428],u_xpb_out[80][428],u_xpb_out[81][428],u_xpb_out[82][428],u_xpb_out[83][428],u_xpb_out[84][428],u_xpb_out[85][428],u_xpb_out[86][428],u_xpb_out[87][428],u_xpb_out[88][428],u_xpb_out[89][428],u_xpb_out[90][428],u_xpb_out[91][428],u_xpb_out[92][428],u_xpb_out[93][428],u_xpb_out[94][428],u_xpb_out[95][428],u_xpb_out[96][428],u_xpb_out[97][428],u_xpb_out[98][428],u_xpb_out[99][428],u_xpb_out[100][428],u_xpb_out[101][428],u_xpb_out[102][428],u_xpb_out[103][428],u_xpb_out[104][428],u_xpb_out[105][428]};

assign col_out_429 = {u_xpb_out[0][429],u_xpb_out[1][429],u_xpb_out[2][429],u_xpb_out[3][429],u_xpb_out[4][429],u_xpb_out[5][429],u_xpb_out[6][429],u_xpb_out[7][429],u_xpb_out[8][429],u_xpb_out[9][429],u_xpb_out[10][429],u_xpb_out[11][429],u_xpb_out[12][429],u_xpb_out[13][429],u_xpb_out[14][429],u_xpb_out[15][429],u_xpb_out[16][429],u_xpb_out[17][429],u_xpb_out[18][429],u_xpb_out[19][429],u_xpb_out[20][429],u_xpb_out[21][429],u_xpb_out[22][429],u_xpb_out[23][429],u_xpb_out[24][429],u_xpb_out[25][429],u_xpb_out[26][429],u_xpb_out[27][429],u_xpb_out[28][429],u_xpb_out[29][429],u_xpb_out[30][429],u_xpb_out[31][429],u_xpb_out[32][429],u_xpb_out[33][429],u_xpb_out[34][429],u_xpb_out[35][429],u_xpb_out[36][429],u_xpb_out[37][429],u_xpb_out[38][429],u_xpb_out[39][429],u_xpb_out[40][429],u_xpb_out[41][429],u_xpb_out[42][429],u_xpb_out[43][429],u_xpb_out[44][429],u_xpb_out[45][429],u_xpb_out[46][429],u_xpb_out[47][429],u_xpb_out[48][429],u_xpb_out[49][429],u_xpb_out[50][429],u_xpb_out[51][429],u_xpb_out[52][429],u_xpb_out[53][429],u_xpb_out[54][429],u_xpb_out[55][429],u_xpb_out[56][429],u_xpb_out[57][429],u_xpb_out[58][429],u_xpb_out[59][429],u_xpb_out[60][429],u_xpb_out[61][429],u_xpb_out[62][429],u_xpb_out[63][429],u_xpb_out[64][429],u_xpb_out[65][429],u_xpb_out[66][429],u_xpb_out[67][429],u_xpb_out[68][429],u_xpb_out[69][429],u_xpb_out[70][429],u_xpb_out[71][429],u_xpb_out[72][429],u_xpb_out[73][429],u_xpb_out[74][429],u_xpb_out[75][429],u_xpb_out[76][429],u_xpb_out[77][429],u_xpb_out[78][429],u_xpb_out[79][429],u_xpb_out[80][429],u_xpb_out[81][429],u_xpb_out[82][429],u_xpb_out[83][429],u_xpb_out[84][429],u_xpb_out[85][429],u_xpb_out[86][429],u_xpb_out[87][429],u_xpb_out[88][429],u_xpb_out[89][429],u_xpb_out[90][429],u_xpb_out[91][429],u_xpb_out[92][429],u_xpb_out[93][429],u_xpb_out[94][429],u_xpb_out[95][429],u_xpb_out[96][429],u_xpb_out[97][429],u_xpb_out[98][429],u_xpb_out[99][429],u_xpb_out[100][429],u_xpb_out[101][429],u_xpb_out[102][429],u_xpb_out[103][429],u_xpb_out[104][429],u_xpb_out[105][429]};

assign col_out_430 = {u_xpb_out[0][430],u_xpb_out[1][430],u_xpb_out[2][430],u_xpb_out[3][430],u_xpb_out[4][430],u_xpb_out[5][430],u_xpb_out[6][430],u_xpb_out[7][430],u_xpb_out[8][430],u_xpb_out[9][430],u_xpb_out[10][430],u_xpb_out[11][430],u_xpb_out[12][430],u_xpb_out[13][430],u_xpb_out[14][430],u_xpb_out[15][430],u_xpb_out[16][430],u_xpb_out[17][430],u_xpb_out[18][430],u_xpb_out[19][430],u_xpb_out[20][430],u_xpb_out[21][430],u_xpb_out[22][430],u_xpb_out[23][430],u_xpb_out[24][430],u_xpb_out[25][430],u_xpb_out[26][430],u_xpb_out[27][430],u_xpb_out[28][430],u_xpb_out[29][430],u_xpb_out[30][430],u_xpb_out[31][430],u_xpb_out[32][430],u_xpb_out[33][430],u_xpb_out[34][430],u_xpb_out[35][430],u_xpb_out[36][430],u_xpb_out[37][430],u_xpb_out[38][430],u_xpb_out[39][430],u_xpb_out[40][430],u_xpb_out[41][430],u_xpb_out[42][430],u_xpb_out[43][430],u_xpb_out[44][430],u_xpb_out[45][430],u_xpb_out[46][430],u_xpb_out[47][430],u_xpb_out[48][430],u_xpb_out[49][430],u_xpb_out[50][430],u_xpb_out[51][430],u_xpb_out[52][430],u_xpb_out[53][430],u_xpb_out[54][430],u_xpb_out[55][430],u_xpb_out[56][430],u_xpb_out[57][430],u_xpb_out[58][430],u_xpb_out[59][430],u_xpb_out[60][430],u_xpb_out[61][430],u_xpb_out[62][430],u_xpb_out[63][430],u_xpb_out[64][430],u_xpb_out[65][430],u_xpb_out[66][430],u_xpb_out[67][430],u_xpb_out[68][430],u_xpb_out[69][430],u_xpb_out[70][430],u_xpb_out[71][430],u_xpb_out[72][430],u_xpb_out[73][430],u_xpb_out[74][430],u_xpb_out[75][430],u_xpb_out[76][430],u_xpb_out[77][430],u_xpb_out[78][430],u_xpb_out[79][430],u_xpb_out[80][430],u_xpb_out[81][430],u_xpb_out[82][430],u_xpb_out[83][430],u_xpb_out[84][430],u_xpb_out[85][430],u_xpb_out[86][430],u_xpb_out[87][430],u_xpb_out[88][430],u_xpb_out[89][430],u_xpb_out[90][430],u_xpb_out[91][430],u_xpb_out[92][430],u_xpb_out[93][430],u_xpb_out[94][430],u_xpb_out[95][430],u_xpb_out[96][430],u_xpb_out[97][430],u_xpb_out[98][430],u_xpb_out[99][430],u_xpb_out[100][430],u_xpb_out[101][430],u_xpb_out[102][430],u_xpb_out[103][430],u_xpb_out[104][430],u_xpb_out[105][430]};

assign col_out_431 = {u_xpb_out[0][431],u_xpb_out[1][431],u_xpb_out[2][431],u_xpb_out[3][431],u_xpb_out[4][431],u_xpb_out[5][431],u_xpb_out[6][431],u_xpb_out[7][431],u_xpb_out[8][431],u_xpb_out[9][431],u_xpb_out[10][431],u_xpb_out[11][431],u_xpb_out[12][431],u_xpb_out[13][431],u_xpb_out[14][431],u_xpb_out[15][431],u_xpb_out[16][431],u_xpb_out[17][431],u_xpb_out[18][431],u_xpb_out[19][431],u_xpb_out[20][431],u_xpb_out[21][431],u_xpb_out[22][431],u_xpb_out[23][431],u_xpb_out[24][431],u_xpb_out[25][431],u_xpb_out[26][431],u_xpb_out[27][431],u_xpb_out[28][431],u_xpb_out[29][431],u_xpb_out[30][431],u_xpb_out[31][431],u_xpb_out[32][431],u_xpb_out[33][431],u_xpb_out[34][431],u_xpb_out[35][431],u_xpb_out[36][431],u_xpb_out[37][431],u_xpb_out[38][431],u_xpb_out[39][431],u_xpb_out[40][431],u_xpb_out[41][431],u_xpb_out[42][431],u_xpb_out[43][431],u_xpb_out[44][431],u_xpb_out[45][431],u_xpb_out[46][431],u_xpb_out[47][431],u_xpb_out[48][431],u_xpb_out[49][431],u_xpb_out[50][431],u_xpb_out[51][431],u_xpb_out[52][431],u_xpb_out[53][431],u_xpb_out[54][431],u_xpb_out[55][431],u_xpb_out[56][431],u_xpb_out[57][431],u_xpb_out[58][431],u_xpb_out[59][431],u_xpb_out[60][431],u_xpb_out[61][431],u_xpb_out[62][431],u_xpb_out[63][431],u_xpb_out[64][431],u_xpb_out[65][431],u_xpb_out[66][431],u_xpb_out[67][431],u_xpb_out[68][431],u_xpb_out[69][431],u_xpb_out[70][431],u_xpb_out[71][431],u_xpb_out[72][431],u_xpb_out[73][431],u_xpb_out[74][431],u_xpb_out[75][431],u_xpb_out[76][431],u_xpb_out[77][431],u_xpb_out[78][431],u_xpb_out[79][431],u_xpb_out[80][431],u_xpb_out[81][431],u_xpb_out[82][431],u_xpb_out[83][431],u_xpb_out[84][431],u_xpb_out[85][431],u_xpb_out[86][431],u_xpb_out[87][431],u_xpb_out[88][431],u_xpb_out[89][431],u_xpb_out[90][431],u_xpb_out[91][431],u_xpb_out[92][431],u_xpb_out[93][431],u_xpb_out[94][431],u_xpb_out[95][431],u_xpb_out[96][431],u_xpb_out[97][431],u_xpb_out[98][431],u_xpb_out[99][431],u_xpb_out[100][431],u_xpb_out[101][431],u_xpb_out[102][431],u_xpb_out[103][431],u_xpb_out[104][431],u_xpb_out[105][431]};

assign col_out_432 = {u_xpb_out[0][432],u_xpb_out[1][432],u_xpb_out[2][432],u_xpb_out[3][432],u_xpb_out[4][432],u_xpb_out[5][432],u_xpb_out[6][432],u_xpb_out[7][432],u_xpb_out[8][432],u_xpb_out[9][432],u_xpb_out[10][432],u_xpb_out[11][432],u_xpb_out[12][432],u_xpb_out[13][432],u_xpb_out[14][432],u_xpb_out[15][432],u_xpb_out[16][432],u_xpb_out[17][432],u_xpb_out[18][432],u_xpb_out[19][432],u_xpb_out[20][432],u_xpb_out[21][432],u_xpb_out[22][432],u_xpb_out[23][432],u_xpb_out[24][432],u_xpb_out[25][432],u_xpb_out[26][432],u_xpb_out[27][432],u_xpb_out[28][432],u_xpb_out[29][432],u_xpb_out[30][432],u_xpb_out[31][432],u_xpb_out[32][432],u_xpb_out[33][432],u_xpb_out[34][432],u_xpb_out[35][432],u_xpb_out[36][432],u_xpb_out[37][432],u_xpb_out[38][432],u_xpb_out[39][432],u_xpb_out[40][432],u_xpb_out[41][432],u_xpb_out[42][432],u_xpb_out[43][432],u_xpb_out[44][432],u_xpb_out[45][432],u_xpb_out[46][432],u_xpb_out[47][432],u_xpb_out[48][432],u_xpb_out[49][432],u_xpb_out[50][432],u_xpb_out[51][432],u_xpb_out[52][432],u_xpb_out[53][432],u_xpb_out[54][432],u_xpb_out[55][432],u_xpb_out[56][432],u_xpb_out[57][432],u_xpb_out[58][432],u_xpb_out[59][432],u_xpb_out[60][432],u_xpb_out[61][432],u_xpb_out[62][432],u_xpb_out[63][432],u_xpb_out[64][432],u_xpb_out[65][432],u_xpb_out[66][432],u_xpb_out[67][432],u_xpb_out[68][432],u_xpb_out[69][432],u_xpb_out[70][432],u_xpb_out[71][432],u_xpb_out[72][432],u_xpb_out[73][432],u_xpb_out[74][432],u_xpb_out[75][432],u_xpb_out[76][432],u_xpb_out[77][432],u_xpb_out[78][432],u_xpb_out[79][432],u_xpb_out[80][432],u_xpb_out[81][432],u_xpb_out[82][432],u_xpb_out[83][432],u_xpb_out[84][432],u_xpb_out[85][432],u_xpb_out[86][432],u_xpb_out[87][432],u_xpb_out[88][432],u_xpb_out[89][432],u_xpb_out[90][432],u_xpb_out[91][432],u_xpb_out[92][432],u_xpb_out[93][432],u_xpb_out[94][432],u_xpb_out[95][432],u_xpb_out[96][432],u_xpb_out[97][432],u_xpb_out[98][432],u_xpb_out[99][432],u_xpb_out[100][432],u_xpb_out[101][432],u_xpb_out[102][432],u_xpb_out[103][432],u_xpb_out[104][432],u_xpb_out[105][432]};

assign col_out_433 = {u_xpb_out[0][433],u_xpb_out[1][433],u_xpb_out[2][433],u_xpb_out[3][433],u_xpb_out[4][433],u_xpb_out[5][433],u_xpb_out[6][433],u_xpb_out[7][433],u_xpb_out[8][433],u_xpb_out[9][433],u_xpb_out[10][433],u_xpb_out[11][433],u_xpb_out[12][433],u_xpb_out[13][433],u_xpb_out[14][433],u_xpb_out[15][433],u_xpb_out[16][433],u_xpb_out[17][433],u_xpb_out[18][433],u_xpb_out[19][433],u_xpb_out[20][433],u_xpb_out[21][433],u_xpb_out[22][433],u_xpb_out[23][433],u_xpb_out[24][433],u_xpb_out[25][433],u_xpb_out[26][433],u_xpb_out[27][433],u_xpb_out[28][433],u_xpb_out[29][433],u_xpb_out[30][433],u_xpb_out[31][433],u_xpb_out[32][433],u_xpb_out[33][433],u_xpb_out[34][433],u_xpb_out[35][433],u_xpb_out[36][433],u_xpb_out[37][433],u_xpb_out[38][433],u_xpb_out[39][433],u_xpb_out[40][433],u_xpb_out[41][433],u_xpb_out[42][433],u_xpb_out[43][433],u_xpb_out[44][433],u_xpb_out[45][433],u_xpb_out[46][433],u_xpb_out[47][433],u_xpb_out[48][433],u_xpb_out[49][433],u_xpb_out[50][433],u_xpb_out[51][433],u_xpb_out[52][433],u_xpb_out[53][433],u_xpb_out[54][433],u_xpb_out[55][433],u_xpb_out[56][433],u_xpb_out[57][433],u_xpb_out[58][433],u_xpb_out[59][433],u_xpb_out[60][433],u_xpb_out[61][433],u_xpb_out[62][433],u_xpb_out[63][433],u_xpb_out[64][433],u_xpb_out[65][433],u_xpb_out[66][433],u_xpb_out[67][433],u_xpb_out[68][433],u_xpb_out[69][433],u_xpb_out[70][433],u_xpb_out[71][433],u_xpb_out[72][433],u_xpb_out[73][433],u_xpb_out[74][433],u_xpb_out[75][433],u_xpb_out[76][433],u_xpb_out[77][433],u_xpb_out[78][433],u_xpb_out[79][433],u_xpb_out[80][433],u_xpb_out[81][433],u_xpb_out[82][433],u_xpb_out[83][433],u_xpb_out[84][433],u_xpb_out[85][433],u_xpb_out[86][433],u_xpb_out[87][433],u_xpb_out[88][433],u_xpb_out[89][433],u_xpb_out[90][433],u_xpb_out[91][433],u_xpb_out[92][433],u_xpb_out[93][433],u_xpb_out[94][433],u_xpb_out[95][433],u_xpb_out[96][433],u_xpb_out[97][433],u_xpb_out[98][433],u_xpb_out[99][433],u_xpb_out[100][433],u_xpb_out[101][433],u_xpb_out[102][433],u_xpb_out[103][433],u_xpb_out[104][433],u_xpb_out[105][433]};

assign col_out_434 = {u_xpb_out[0][434],u_xpb_out[1][434],u_xpb_out[2][434],u_xpb_out[3][434],u_xpb_out[4][434],u_xpb_out[5][434],u_xpb_out[6][434],u_xpb_out[7][434],u_xpb_out[8][434],u_xpb_out[9][434],u_xpb_out[10][434],u_xpb_out[11][434],u_xpb_out[12][434],u_xpb_out[13][434],u_xpb_out[14][434],u_xpb_out[15][434],u_xpb_out[16][434],u_xpb_out[17][434],u_xpb_out[18][434],u_xpb_out[19][434],u_xpb_out[20][434],u_xpb_out[21][434],u_xpb_out[22][434],u_xpb_out[23][434],u_xpb_out[24][434],u_xpb_out[25][434],u_xpb_out[26][434],u_xpb_out[27][434],u_xpb_out[28][434],u_xpb_out[29][434],u_xpb_out[30][434],u_xpb_out[31][434],u_xpb_out[32][434],u_xpb_out[33][434],u_xpb_out[34][434],u_xpb_out[35][434],u_xpb_out[36][434],u_xpb_out[37][434],u_xpb_out[38][434],u_xpb_out[39][434],u_xpb_out[40][434],u_xpb_out[41][434],u_xpb_out[42][434],u_xpb_out[43][434],u_xpb_out[44][434],u_xpb_out[45][434],u_xpb_out[46][434],u_xpb_out[47][434],u_xpb_out[48][434],u_xpb_out[49][434],u_xpb_out[50][434],u_xpb_out[51][434],u_xpb_out[52][434],u_xpb_out[53][434],u_xpb_out[54][434],u_xpb_out[55][434],u_xpb_out[56][434],u_xpb_out[57][434],u_xpb_out[58][434],u_xpb_out[59][434],u_xpb_out[60][434],u_xpb_out[61][434],u_xpb_out[62][434],u_xpb_out[63][434],u_xpb_out[64][434],u_xpb_out[65][434],u_xpb_out[66][434],u_xpb_out[67][434],u_xpb_out[68][434],u_xpb_out[69][434],u_xpb_out[70][434],u_xpb_out[71][434],u_xpb_out[72][434],u_xpb_out[73][434],u_xpb_out[74][434],u_xpb_out[75][434],u_xpb_out[76][434],u_xpb_out[77][434],u_xpb_out[78][434],u_xpb_out[79][434],u_xpb_out[80][434],u_xpb_out[81][434],u_xpb_out[82][434],u_xpb_out[83][434],u_xpb_out[84][434],u_xpb_out[85][434],u_xpb_out[86][434],u_xpb_out[87][434],u_xpb_out[88][434],u_xpb_out[89][434],u_xpb_out[90][434],u_xpb_out[91][434],u_xpb_out[92][434],u_xpb_out[93][434],u_xpb_out[94][434],u_xpb_out[95][434],u_xpb_out[96][434],u_xpb_out[97][434],u_xpb_out[98][434],u_xpb_out[99][434],u_xpb_out[100][434],u_xpb_out[101][434],u_xpb_out[102][434],u_xpb_out[103][434],u_xpb_out[104][434],u_xpb_out[105][434]};

assign col_out_435 = {u_xpb_out[0][435],u_xpb_out[1][435],u_xpb_out[2][435],u_xpb_out[3][435],u_xpb_out[4][435],u_xpb_out[5][435],u_xpb_out[6][435],u_xpb_out[7][435],u_xpb_out[8][435],u_xpb_out[9][435],u_xpb_out[10][435],u_xpb_out[11][435],u_xpb_out[12][435],u_xpb_out[13][435],u_xpb_out[14][435],u_xpb_out[15][435],u_xpb_out[16][435],u_xpb_out[17][435],u_xpb_out[18][435],u_xpb_out[19][435],u_xpb_out[20][435],u_xpb_out[21][435],u_xpb_out[22][435],u_xpb_out[23][435],u_xpb_out[24][435],u_xpb_out[25][435],u_xpb_out[26][435],u_xpb_out[27][435],u_xpb_out[28][435],u_xpb_out[29][435],u_xpb_out[30][435],u_xpb_out[31][435],u_xpb_out[32][435],u_xpb_out[33][435],u_xpb_out[34][435],u_xpb_out[35][435],u_xpb_out[36][435],u_xpb_out[37][435],u_xpb_out[38][435],u_xpb_out[39][435],u_xpb_out[40][435],u_xpb_out[41][435],u_xpb_out[42][435],u_xpb_out[43][435],u_xpb_out[44][435],u_xpb_out[45][435],u_xpb_out[46][435],u_xpb_out[47][435],u_xpb_out[48][435],u_xpb_out[49][435],u_xpb_out[50][435],u_xpb_out[51][435],u_xpb_out[52][435],u_xpb_out[53][435],u_xpb_out[54][435],u_xpb_out[55][435],u_xpb_out[56][435],u_xpb_out[57][435],u_xpb_out[58][435],u_xpb_out[59][435],u_xpb_out[60][435],u_xpb_out[61][435],u_xpb_out[62][435],u_xpb_out[63][435],u_xpb_out[64][435],u_xpb_out[65][435],u_xpb_out[66][435],u_xpb_out[67][435],u_xpb_out[68][435],u_xpb_out[69][435],u_xpb_out[70][435],u_xpb_out[71][435],u_xpb_out[72][435],u_xpb_out[73][435],u_xpb_out[74][435],u_xpb_out[75][435],u_xpb_out[76][435],u_xpb_out[77][435],u_xpb_out[78][435],u_xpb_out[79][435],u_xpb_out[80][435],u_xpb_out[81][435],u_xpb_out[82][435],u_xpb_out[83][435],u_xpb_out[84][435],u_xpb_out[85][435],u_xpb_out[86][435],u_xpb_out[87][435],u_xpb_out[88][435],u_xpb_out[89][435],u_xpb_out[90][435],u_xpb_out[91][435],u_xpb_out[92][435],u_xpb_out[93][435],u_xpb_out[94][435],u_xpb_out[95][435],u_xpb_out[96][435],u_xpb_out[97][435],u_xpb_out[98][435],u_xpb_out[99][435],u_xpb_out[100][435],u_xpb_out[101][435],u_xpb_out[102][435],u_xpb_out[103][435],u_xpb_out[104][435],u_xpb_out[105][435]};

assign col_out_436 = {u_xpb_out[0][436],u_xpb_out[1][436],u_xpb_out[2][436],u_xpb_out[3][436],u_xpb_out[4][436],u_xpb_out[5][436],u_xpb_out[6][436],u_xpb_out[7][436],u_xpb_out[8][436],u_xpb_out[9][436],u_xpb_out[10][436],u_xpb_out[11][436],u_xpb_out[12][436],u_xpb_out[13][436],u_xpb_out[14][436],u_xpb_out[15][436],u_xpb_out[16][436],u_xpb_out[17][436],u_xpb_out[18][436],u_xpb_out[19][436],u_xpb_out[20][436],u_xpb_out[21][436],u_xpb_out[22][436],u_xpb_out[23][436],u_xpb_out[24][436],u_xpb_out[25][436],u_xpb_out[26][436],u_xpb_out[27][436],u_xpb_out[28][436],u_xpb_out[29][436],u_xpb_out[30][436],u_xpb_out[31][436],u_xpb_out[32][436],u_xpb_out[33][436],u_xpb_out[34][436],u_xpb_out[35][436],u_xpb_out[36][436],u_xpb_out[37][436],u_xpb_out[38][436],u_xpb_out[39][436],u_xpb_out[40][436],u_xpb_out[41][436],u_xpb_out[42][436],u_xpb_out[43][436],u_xpb_out[44][436],u_xpb_out[45][436],u_xpb_out[46][436],u_xpb_out[47][436],u_xpb_out[48][436],u_xpb_out[49][436],u_xpb_out[50][436],u_xpb_out[51][436],u_xpb_out[52][436],u_xpb_out[53][436],u_xpb_out[54][436],u_xpb_out[55][436],u_xpb_out[56][436],u_xpb_out[57][436],u_xpb_out[58][436],u_xpb_out[59][436],u_xpb_out[60][436],u_xpb_out[61][436],u_xpb_out[62][436],u_xpb_out[63][436],u_xpb_out[64][436],u_xpb_out[65][436],u_xpb_out[66][436],u_xpb_out[67][436],u_xpb_out[68][436],u_xpb_out[69][436],u_xpb_out[70][436],u_xpb_out[71][436],u_xpb_out[72][436],u_xpb_out[73][436],u_xpb_out[74][436],u_xpb_out[75][436],u_xpb_out[76][436],u_xpb_out[77][436],u_xpb_out[78][436],u_xpb_out[79][436],u_xpb_out[80][436],u_xpb_out[81][436],u_xpb_out[82][436],u_xpb_out[83][436],u_xpb_out[84][436],u_xpb_out[85][436],u_xpb_out[86][436],u_xpb_out[87][436],u_xpb_out[88][436],u_xpb_out[89][436],u_xpb_out[90][436],u_xpb_out[91][436],u_xpb_out[92][436],u_xpb_out[93][436],u_xpb_out[94][436],u_xpb_out[95][436],u_xpb_out[96][436],u_xpb_out[97][436],u_xpb_out[98][436],u_xpb_out[99][436],u_xpb_out[100][436],u_xpb_out[101][436],u_xpb_out[102][436],u_xpb_out[103][436],u_xpb_out[104][436],u_xpb_out[105][436]};

assign col_out_437 = {u_xpb_out[0][437],u_xpb_out[1][437],u_xpb_out[2][437],u_xpb_out[3][437],u_xpb_out[4][437],u_xpb_out[5][437],u_xpb_out[6][437],u_xpb_out[7][437],u_xpb_out[8][437],u_xpb_out[9][437],u_xpb_out[10][437],u_xpb_out[11][437],u_xpb_out[12][437],u_xpb_out[13][437],u_xpb_out[14][437],u_xpb_out[15][437],u_xpb_out[16][437],u_xpb_out[17][437],u_xpb_out[18][437],u_xpb_out[19][437],u_xpb_out[20][437],u_xpb_out[21][437],u_xpb_out[22][437],u_xpb_out[23][437],u_xpb_out[24][437],u_xpb_out[25][437],u_xpb_out[26][437],u_xpb_out[27][437],u_xpb_out[28][437],u_xpb_out[29][437],u_xpb_out[30][437],u_xpb_out[31][437],u_xpb_out[32][437],u_xpb_out[33][437],u_xpb_out[34][437],u_xpb_out[35][437],u_xpb_out[36][437],u_xpb_out[37][437],u_xpb_out[38][437],u_xpb_out[39][437],u_xpb_out[40][437],u_xpb_out[41][437],u_xpb_out[42][437],u_xpb_out[43][437],u_xpb_out[44][437],u_xpb_out[45][437],u_xpb_out[46][437],u_xpb_out[47][437],u_xpb_out[48][437],u_xpb_out[49][437],u_xpb_out[50][437],u_xpb_out[51][437],u_xpb_out[52][437],u_xpb_out[53][437],u_xpb_out[54][437],u_xpb_out[55][437],u_xpb_out[56][437],u_xpb_out[57][437],u_xpb_out[58][437],u_xpb_out[59][437],u_xpb_out[60][437],u_xpb_out[61][437],u_xpb_out[62][437],u_xpb_out[63][437],u_xpb_out[64][437],u_xpb_out[65][437],u_xpb_out[66][437],u_xpb_out[67][437],u_xpb_out[68][437],u_xpb_out[69][437],u_xpb_out[70][437],u_xpb_out[71][437],u_xpb_out[72][437],u_xpb_out[73][437],u_xpb_out[74][437],u_xpb_out[75][437],u_xpb_out[76][437],u_xpb_out[77][437],u_xpb_out[78][437],u_xpb_out[79][437],u_xpb_out[80][437],u_xpb_out[81][437],u_xpb_out[82][437],u_xpb_out[83][437],u_xpb_out[84][437],u_xpb_out[85][437],u_xpb_out[86][437],u_xpb_out[87][437],u_xpb_out[88][437],u_xpb_out[89][437],u_xpb_out[90][437],u_xpb_out[91][437],u_xpb_out[92][437],u_xpb_out[93][437],u_xpb_out[94][437],u_xpb_out[95][437],u_xpb_out[96][437],u_xpb_out[97][437],u_xpb_out[98][437],u_xpb_out[99][437],u_xpb_out[100][437],u_xpb_out[101][437],u_xpb_out[102][437],u_xpb_out[103][437],u_xpb_out[104][437],u_xpb_out[105][437]};

assign col_out_438 = {u_xpb_out[0][438],u_xpb_out[1][438],u_xpb_out[2][438],u_xpb_out[3][438],u_xpb_out[4][438],u_xpb_out[5][438],u_xpb_out[6][438],u_xpb_out[7][438],u_xpb_out[8][438],u_xpb_out[9][438],u_xpb_out[10][438],u_xpb_out[11][438],u_xpb_out[12][438],u_xpb_out[13][438],u_xpb_out[14][438],u_xpb_out[15][438],u_xpb_out[16][438],u_xpb_out[17][438],u_xpb_out[18][438],u_xpb_out[19][438],u_xpb_out[20][438],u_xpb_out[21][438],u_xpb_out[22][438],u_xpb_out[23][438],u_xpb_out[24][438],u_xpb_out[25][438],u_xpb_out[26][438],u_xpb_out[27][438],u_xpb_out[28][438],u_xpb_out[29][438],u_xpb_out[30][438],u_xpb_out[31][438],u_xpb_out[32][438],u_xpb_out[33][438],u_xpb_out[34][438],u_xpb_out[35][438],u_xpb_out[36][438],u_xpb_out[37][438],u_xpb_out[38][438],u_xpb_out[39][438],u_xpb_out[40][438],u_xpb_out[41][438],u_xpb_out[42][438],u_xpb_out[43][438],u_xpb_out[44][438],u_xpb_out[45][438],u_xpb_out[46][438],u_xpb_out[47][438],u_xpb_out[48][438],u_xpb_out[49][438],u_xpb_out[50][438],u_xpb_out[51][438],u_xpb_out[52][438],u_xpb_out[53][438],u_xpb_out[54][438],u_xpb_out[55][438],u_xpb_out[56][438],u_xpb_out[57][438],u_xpb_out[58][438],u_xpb_out[59][438],u_xpb_out[60][438],u_xpb_out[61][438],u_xpb_out[62][438],u_xpb_out[63][438],u_xpb_out[64][438],u_xpb_out[65][438],u_xpb_out[66][438],u_xpb_out[67][438],u_xpb_out[68][438],u_xpb_out[69][438],u_xpb_out[70][438],u_xpb_out[71][438],u_xpb_out[72][438],u_xpb_out[73][438],u_xpb_out[74][438],u_xpb_out[75][438],u_xpb_out[76][438],u_xpb_out[77][438],u_xpb_out[78][438],u_xpb_out[79][438],u_xpb_out[80][438],u_xpb_out[81][438],u_xpb_out[82][438],u_xpb_out[83][438],u_xpb_out[84][438],u_xpb_out[85][438],u_xpb_out[86][438],u_xpb_out[87][438],u_xpb_out[88][438],u_xpb_out[89][438],u_xpb_out[90][438],u_xpb_out[91][438],u_xpb_out[92][438],u_xpb_out[93][438],u_xpb_out[94][438],u_xpb_out[95][438],u_xpb_out[96][438],u_xpb_out[97][438],u_xpb_out[98][438],u_xpb_out[99][438],u_xpb_out[100][438],u_xpb_out[101][438],u_xpb_out[102][438],u_xpb_out[103][438],u_xpb_out[104][438],u_xpb_out[105][438]};

assign col_out_439 = {u_xpb_out[0][439],u_xpb_out[1][439],u_xpb_out[2][439],u_xpb_out[3][439],u_xpb_out[4][439],u_xpb_out[5][439],u_xpb_out[6][439],u_xpb_out[7][439],u_xpb_out[8][439],u_xpb_out[9][439],u_xpb_out[10][439],u_xpb_out[11][439],u_xpb_out[12][439],u_xpb_out[13][439],u_xpb_out[14][439],u_xpb_out[15][439],u_xpb_out[16][439],u_xpb_out[17][439],u_xpb_out[18][439],u_xpb_out[19][439],u_xpb_out[20][439],u_xpb_out[21][439],u_xpb_out[22][439],u_xpb_out[23][439],u_xpb_out[24][439],u_xpb_out[25][439],u_xpb_out[26][439],u_xpb_out[27][439],u_xpb_out[28][439],u_xpb_out[29][439],u_xpb_out[30][439],u_xpb_out[31][439],u_xpb_out[32][439],u_xpb_out[33][439],u_xpb_out[34][439],u_xpb_out[35][439],u_xpb_out[36][439],u_xpb_out[37][439],u_xpb_out[38][439],u_xpb_out[39][439],u_xpb_out[40][439],u_xpb_out[41][439],u_xpb_out[42][439],u_xpb_out[43][439],u_xpb_out[44][439],u_xpb_out[45][439],u_xpb_out[46][439],u_xpb_out[47][439],u_xpb_out[48][439],u_xpb_out[49][439],u_xpb_out[50][439],u_xpb_out[51][439],u_xpb_out[52][439],u_xpb_out[53][439],u_xpb_out[54][439],u_xpb_out[55][439],u_xpb_out[56][439],u_xpb_out[57][439],u_xpb_out[58][439],u_xpb_out[59][439],u_xpb_out[60][439],u_xpb_out[61][439],u_xpb_out[62][439],u_xpb_out[63][439],u_xpb_out[64][439],u_xpb_out[65][439],u_xpb_out[66][439],u_xpb_out[67][439],u_xpb_out[68][439],u_xpb_out[69][439],u_xpb_out[70][439],u_xpb_out[71][439],u_xpb_out[72][439],u_xpb_out[73][439],u_xpb_out[74][439],u_xpb_out[75][439],u_xpb_out[76][439],u_xpb_out[77][439],u_xpb_out[78][439],u_xpb_out[79][439],u_xpb_out[80][439],u_xpb_out[81][439],u_xpb_out[82][439],u_xpb_out[83][439],u_xpb_out[84][439],u_xpb_out[85][439],u_xpb_out[86][439],u_xpb_out[87][439],u_xpb_out[88][439],u_xpb_out[89][439],u_xpb_out[90][439],u_xpb_out[91][439],u_xpb_out[92][439],u_xpb_out[93][439],u_xpb_out[94][439],u_xpb_out[95][439],u_xpb_out[96][439],u_xpb_out[97][439],u_xpb_out[98][439],u_xpb_out[99][439],u_xpb_out[100][439],u_xpb_out[101][439],u_xpb_out[102][439],u_xpb_out[103][439],u_xpb_out[104][439],u_xpb_out[105][439]};

assign col_out_440 = {u_xpb_out[0][440],u_xpb_out[1][440],u_xpb_out[2][440],u_xpb_out[3][440],u_xpb_out[4][440],u_xpb_out[5][440],u_xpb_out[6][440],u_xpb_out[7][440],u_xpb_out[8][440],u_xpb_out[9][440],u_xpb_out[10][440],u_xpb_out[11][440],u_xpb_out[12][440],u_xpb_out[13][440],u_xpb_out[14][440],u_xpb_out[15][440],u_xpb_out[16][440],u_xpb_out[17][440],u_xpb_out[18][440],u_xpb_out[19][440],u_xpb_out[20][440],u_xpb_out[21][440],u_xpb_out[22][440],u_xpb_out[23][440],u_xpb_out[24][440],u_xpb_out[25][440],u_xpb_out[26][440],u_xpb_out[27][440],u_xpb_out[28][440],u_xpb_out[29][440],u_xpb_out[30][440],u_xpb_out[31][440],u_xpb_out[32][440],u_xpb_out[33][440],u_xpb_out[34][440],u_xpb_out[35][440],u_xpb_out[36][440],u_xpb_out[37][440],u_xpb_out[38][440],u_xpb_out[39][440],u_xpb_out[40][440],u_xpb_out[41][440],u_xpb_out[42][440],u_xpb_out[43][440],u_xpb_out[44][440],u_xpb_out[45][440],u_xpb_out[46][440],u_xpb_out[47][440],u_xpb_out[48][440],u_xpb_out[49][440],u_xpb_out[50][440],u_xpb_out[51][440],u_xpb_out[52][440],u_xpb_out[53][440],u_xpb_out[54][440],u_xpb_out[55][440],u_xpb_out[56][440],u_xpb_out[57][440],u_xpb_out[58][440],u_xpb_out[59][440],u_xpb_out[60][440],u_xpb_out[61][440],u_xpb_out[62][440],u_xpb_out[63][440],u_xpb_out[64][440],u_xpb_out[65][440],u_xpb_out[66][440],u_xpb_out[67][440],u_xpb_out[68][440],u_xpb_out[69][440],u_xpb_out[70][440],u_xpb_out[71][440],u_xpb_out[72][440],u_xpb_out[73][440],u_xpb_out[74][440],u_xpb_out[75][440],u_xpb_out[76][440],u_xpb_out[77][440],u_xpb_out[78][440],u_xpb_out[79][440],u_xpb_out[80][440],u_xpb_out[81][440],u_xpb_out[82][440],u_xpb_out[83][440],u_xpb_out[84][440],u_xpb_out[85][440],u_xpb_out[86][440],u_xpb_out[87][440],u_xpb_out[88][440],u_xpb_out[89][440],u_xpb_out[90][440],u_xpb_out[91][440],u_xpb_out[92][440],u_xpb_out[93][440],u_xpb_out[94][440],u_xpb_out[95][440],u_xpb_out[96][440],u_xpb_out[97][440],u_xpb_out[98][440],u_xpb_out[99][440],u_xpb_out[100][440],u_xpb_out[101][440],u_xpb_out[102][440],u_xpb_out[103][440],u_xpb_out[104][440],u_xpb_out[105][440]};

assign col_out_441 = {u_xpb_out[0][441],u_xpb_out[1][441],u_xpb_out[2][441],u_xpb_out[3][441],u_xpb_out[4][441],u_xpb_out[5][441],u_xpb_out[6][441],u_xpb_out[7][441],u_xpb_out[8][441],u_xpb_out[9][441],u_xpb_out[10][441],u_xpb_out[11][441],u_xpb_out[12][441],u_xpb_out[13][441],u_xpb_out[14][441],u_xpb_out[15][441],u_xpb_out[16][441],u_xpb_out[17][441],u_xpb_out[18][441],u_xpb_out[19][441],u_xpb_out[20][441],u_xpb_out[21][441],u_xpb_out[22][441],u_xpb_out[23][441],u_xpb_out[24][441],u_xpb_out[25][441],u_xpb_out[26][441],u_xpb_out[27][441],u_xpb_out[28][441],u_xpb_out[29][441],u_xpb_out[30][441],u_xpb_out[31][441],u_xpb_out[32][441],u_xpb_out[33][441],u_xpb_out[34][441],u_xpb_out[35][441],u_xpb_out[36][441],u_xpb_out[37][441],u_xpb_out[38][441],u_xpb_out[39][441],u_xpb_out[40][441],u_xpb_out[41][441],u_xpb_out[42][441],u_xpb_out[43][441],u_xpb_out[44][441],u_xpb_out[45][441],u_xpb_out[46][441],u_xpb_out[47][441],u_xpb_out[48][441],u_xpb_out[49][441],u_xpb_out[50][441],u_xpb_out[51][441],u_xpb_out[52][441],u_xpb_out[53][441],u_xpb_out[54][441],u_xpb_out[55][441],u_xpb_out[56][441],u_xpb_out[57][441],u_xpb_out[58][441],u_xpb_out[59][441],u_xpb_out[60][441],u_xpb_out[61][441],u_xpb_out[62][441],u_xpb_out[63][441],u_xpb_out[64][441],u_xpb_out[65][441],u_xpb_out[66][441],u_xpb_out[67][441],u_xpb_out[68][441],u_xpb_out[69][441],u_xpb_out[70][441],u_xpb_out[71][441],u_xpb_out[72][441],u_xpb_out[73][441],u_xpb_out[74][441],u_xpb_out[75][441],u_xpb_out[76][441],u_xpb_out[77][441],u_xpb_out[78][441],u_xpb_out[79][441],u_xpb_out[80][441],u_xpb_out[81][441],u_xpb_out[82][441],u_xpb_out[83][441],u_xpb_out[84][441],u_xpb_out[85][441],u_xpb_out[86][441],u_xpb_out[87][441],u_xpb_out[88][441],u_xpb_out[89][441],u_xpb_out[90][441],u_xpb_out[91][441],u_xpb_out[92][441],u_xpb_out[93][441],u_xpb_out[94][441],u_xpb_out[95][441],u_xpb_out[96][441],u_xpb_out[97][441],u_xpb_out[98][441],u_xpb_out[99][441],u_xpb_out[100][441],u_xpb_out[101][441],u_xpb_out[102][441],u_xpb_out[103][441],u_xpb_out[104][441],u_xpb_out[105][441]};

assign col_out_442 = {u_xpb_out[0][442],u_xpb_out[1][442],u_xpb_out[2][442],u_xpb_out[3][442],u_xpb_out[4][442],u_xpb_out[5][442],u_xpb_out[6][442],u_xpb_out[7][442],u_xpb_out[8][442],u_xpb_out[9][442],u_xpb_out[10][442],u_xpb_out[11][442],u_xpb_out[12][442],u_xpb_out[13][442],u_xpb_out[14][442],u_xpb_out[15][442],u_xpb_out[16][442],u_xpb_out[17][442],u_xpb_out[18][442],u_xpb_out[19][442],u_xpb_out[20][442],u_xpb_out[21][442],u_xpb_out[22][442],u_xpb_out[23][442],u_xpb_out[24][442],u_xpb_out[25][442],u_xpb_out[26][442],u_xpb_out[27][442],u_xpb_out[28][442],u_xpb_out[29][442],u_xpb_out[30][442],u_xpb_out[31][442],u_xpb_out[32][442],u_xpb_out[33][442],u_xpb_out[34][442],u_xpb_out[35][442],u_xpb_out[36][442],u_xpb_out[37][442],u_xpb_out[38][442],u_xpb_out[39][442],u_xpb_out[40][442],u_xpb_out[41][442],u_xpb_out[42][442],u_xpb_out[43][442],u_xpb_out[44][442],u_xpb_out[45][442],u_xpb_out[46][442],u_xpb_out[47][442],u_xpb_out[48][442],u_xpb_out[49][442],u_xpb_out[50][442],u_xpb_out[51][442],u_xpb_out[52][442],u_xpb_out[53][442],u_xpb_out[54][442],u_xpb_out[55][442],u_xpb_out[56][442],u_xpb_out[57][442],u_xpb_out[58][442],u_xpb_out[59][442],u_xpb_out[60][442],u_xpb_out[61][442],u_xpb_out[62][442],u_xpb_out[63][442],u_xpb_out[64][442],u_xpb_out[65][442],u_xpb_out[66][442],u_xpb_out[67][442],u_xpb_out[68][442],u_xpb_out[69][442],u_xpb_out[70][442],u_xpb_out[71][442],u_xpb_out[72][442],u_xpb_out[73][442],u_xpb_out[74][442],u_xpb_out[75][442],u_xpb_out[76][442],u_xpb_out[77][442],u_xpb_out[78][442],u_xpb_out[79][442],u_xpb_out[80][442],u_xpb_out[81][442],u_xpb_out[82][442],u_xpb_out[83][442],u_xpb_out[84][442],u_xpb_out[85][442],u_xpb_out[86][442],u_xpb_out[87][442],u_xpb_out[88][442],u_xpb_out[89][442],u_xpb_out[90][442],u_xpb_out[91][442],u_xpb_out[92][442],u_xpb_out[93][442],u_xpb_out[94][442],u_xpb_out[95][442],u_xpb_out[96][442],u_xpb_out[97][442],u_xpb_out[98][442],u_xpb_out[99][442],u_xpb_out[100][442],u_xpb_out[101][442],u_xpb_out[102][442],u_xpb_out[103][442],u_xpb_out[104][442],u_xpb_out[105][442]};

assign col_out_443 = {u_xpb_out[0][443],u_xpb_out[1][443],u_xpb_out[2][443],u_xpb_out[3][443],u_xpb_out[4][443],u_xpb_out[5][443],u_xpb_out[6][443],u_xpb_out[7][443],u_xpb_out[8][443],u_xpb_out[9][443],u_xpb_out[10][443],u_xpb_out[11][443],u_xpb_out[12][443],u_xpb_out[13][443],u_xpb_out[14][443],u_xpb_out[15][443],u_xpb_out[16][443],u_xpb_out[17][443],u_xpb_out[18][443],u_xpb_out[19][443],u_xpb_out[20][443],u_xpb_out[21][443],u_xpb_out[22][443],u_xpb_out[23][443],u_xpb_out[24][443],u_xpb_out[25][443],u_xpb_out[26][443],u_xpb_out[27][443],u_xpb_out[28][443],u_xpb_out[29][443],u_xpb_out[30][443],u_xpb_out[31][443],u_xpb_out[32][443],u_xpb_out[33][443],u_xpb_out[34][443],u_xpb_out[35][443],u_xpb_out[36][443],u_xpb_out[37][443],u_xpb_out[38][443],u_xpb_out[39][443],u_xpb_out[40][443],u_xpb_out[41][443],u_xpb_out[42][443],u_xpb_out[43][443],u_xpb_out[44][443],u_xpb_out[45][443],u_xpb_out[46][443],u_xpb_out[47][443],u_xpb_out[48][443],u_xpb_out[49][443],u_xpb_out[50][443],u_xpb_out[51][443],u_xpb_out[52][443],u_xpb_out[53][443],u_xpb_out[54][443],u_xpb_out[55][443],u_xpb_out[56][443],u_xpb_out[57][443],u_xpb_out[58][443],u_xpb_out[59][443],u_xpb_out[60][443],u_xpb_out[61][443],u_xpb_out[62][443],u_xpb_out[63][443],u_xpb_out[64][443],u_xpb_out[65][443],u_xpb_out[66][443],u_xpb_out[67][443],u_xpb_out[68][443],u_xpb_out[69][443],u_xpb_out[70][443],u_xpb_out[71][443],u_xpb_out[72][443],u_xpb_out[73][443],u_xpb_out[74][443],u_xpb_out[75][443],u_xpb_out[76][443],u_xpb_out[77][443],u_xpb_out[78][443],u_xpb_out[79][443],u_xpb_out[80][443],u_xpb_out[81][443],u_xpb_out[82][443],u_xpb_out[83][443],u_xpb_out[84][443],u_xpb_out[85][443],u_xpb_out[86][443],u_xpb_out[87][443],u_xpb_out[88][443],u_xpb_out[89][443],u_xpb_out[90][443],u_xpb_out[91][443],u_xpb_out[92][443],u_xpb_out[93][443],u_xpb_out[94][443],u_xpb_out[95][443],u_xpb_out[96][443],u_xpb_out[97][443],u_xpb_out[98][443],u_xpb_out[99][443],u_xpb_out[100][443],u_xpb_out[101][443],u_xpb_out[102][443],u_xpb_out[103][443],u_xpb_out[104][443],u_xpb_out[105][443]};

assign col_out_444 = {u_xpb_out[0][444],u_xpb_out[1][444],u_xpb_out[2][444],u_xpb_out[3][444],u_xpb_out[4][444],u_xpb_out[5][444],u_xpb_out[6][444],u_xpb_out[7][444],u_xpb_out[8][444],u_xpb_out[9][444],u_xpb_out[10][444],u_xpb_out[11][444],u_xpb_out[12][444],u_xpb_out[13][444],u_xpb_out[14][444],u_xpb_out[15][444],u_xpb_out[16][444],u_xpb_out[17][444],u_xpb_out[18][444],u_xpb_out[19][444],u_xpb_out[20][444],u_xpb_out[21][444],u_xpb_out[22][444],u_xpb_out[23][444],u_xpb_out[24][444],u_xpb_out[25][444],u_xpb_out[26][444],u_xpb_out[27][444],u_xpb_out[28][444],u_xpb_out[29][444],u_xpb_out[30][444],u_xpb_out[31][444],u_xpb_out[32][444],u_xpb_out[33][444],u_xpb_out[34][444],u_xpb_out[35][444],u_xpb_out[36][444],u_xpb_out[37][444],u_xpb_out[38][444],u_xpb_out[39][444],u_xpb_out[40][444],u_xpb_out[41][444],u_xpb_out[42][444],u_xpb_out[43][444],u_xpb_out[44][444],u_xpb_out[45][444],u_xpb_out[46][444],u_xpb_out[47][444],u_xpb_out[48][444],u_xpb_out[49][444],u_xpb_out[50][444],u_xpb_out[51][444],u_xpb_out[52][444],u_xpb_out[53][444],u_xpb_out[54][444],u_xpb_out[55][444],u_xpb_out[56][444],u_xpb_out[57][444],u_xpb_out[58][444],u_xpb_out[59][444],u_xpb_out[60][444],u_xpb_out[61][444],u_xpb_out[62][444],u_xpb_out[63][444],u_xpb_out[64][444],u_xpb_out[65][444],u_xpb_out[66][444],u_xpb_out[67][444],u_xpb_out[68][444],u_xpb_out[69][444],u_xpb_out[70][444],u_xpb_out[71][444],u_xpb_out[72][444],u_xpb_out[73][444],u_xpb_out[74][444],u_xpb_out[75][444],u_xpb_out[76][444],u_xpb_out[77][444],u_xpb_out[78][444],u_xpb_out[79][444],u_xpb_out[80][444],u_xpb_out[81][444],u_xpb_out[82][444],u_xpb_out[83][444],u_xpb_out[84][444],u_xpb_out[85][444],u_xpb_out[86][444],u_xpb_out[87][444],u_xpb_out[88][444],u_xpb_out[89][444],u_xpb_out[90][444],u_xpb_out[91][444],u_xpb_out[92][444],u_xpb_out[93][444],u_xpb_out[94][444],u_xpb_out[95][444],u_xpb_out[96][444],u_xpb_out[97][444],u_xpb_out[98][444],u_xpb_out[99][444],u_xpb_out[100][444],u_xpb_out[101][444],u_xpb_out[102][444],u_xpb_out[103][444],u_xpb_out[104][444],u_xpb_out[105][444]};

assign col_out_445 = {u_xpb_out[0][445],u_xpb_out[1][445],u_xpb_out[2][445],u_xpb_out[3][445],u_xpb_out[4][445],u_xpb_out[5][445],u_xpb_out[6][445],u_xpb_out[7][445],u_xpb_out[8][445],u_xpb_out[9][445],u_xpb_out[10][445],u_xpb_out[11][445],u_xpb_out[12][445],u_xpb_out[13][445],u_xpb_out[14][445],u_xpb_out[15][445],u_xpb_out[16][445],u_xpb_out[17][445],u_xpb_out[18][445],u_xpb_out[19][445],u_xpb_out[20][445],u_xpb_out[21][445],u_xpb_out[22][445],u_xpb_out[23][445],u_xpb_out[24][445],u_xpb_out[25][445],u_xpb_out[26][445],u_xpb_out[27][445],u_xpb_out[28][445],u_xpb_out[29][445],u_xpb_out[30][445],u_xpb_out[31][445],u_xpb_out[32][445],u_xpb_out[33][445],u_xpb_out[34][445],u_xpb_out[35][445],u_xpb_out[36][445],u_xpb_out[37][445],u_xpb_out[38][445],u_xpb_out[39][445],u_xpb_out[40][445],u_xpb_out[41][445],u_xpb_out[42][445],u_xpb_out[43][445],u_xpb_out[44][445],u_xpb_out[45][445],u_xpb_out[46][445],u_xpb_out[47][445],u_xpb_out[48][445],u_xpb_out[49][445],u_xpb_out[50][445],u_xpb_out[51][445],u_xpb_out[52][445],u_xpb_out[53][445],u_xpb_out[54][445],u_xpb_out[55][445],u_xpb_out[56][445],u_xpb_out[57][445],u_xpb_out[58][445],u_xpb_out[59][445],u_xpb_out[60][445],u_xpb_out[61][445],u_xpb_out[62][445],u_xpb_out[63][445],u_xpb_out[64][445],u_xpb_out[65][445],u_xpb_out[66][445],u_xpb_out[67][445],u_xpb_out[68][445],u_xpb_out[69][445],u_xpb_out[70][445],u_xpb_out[71][445],u_xpb_out[72][445],u_xpb_out[73][445],u_xpb_out[74][445],u_xpb_out[75][445],u_xpb_out[76][445],u_xpb_out[77][445],u_xpb_out[78][445],u_xpb_out[79][445],u_xpb_out[80][445],u_xpb_out[81][445],u_xpb_out[82][445],u_xpb_out[83][445],u_xpb_out[84][445],u_xpb_out[85][445],u_xpb_out[86][445],u_xpb_out[87][445],u_xpb_out[88][445],u_xpb_out[89][445],u_xpb_out[90][445],u_xpb_out[91][445],u_xpb_out[92][445],u_xpb_out[93][445],u_xpb_out[94][445],u_xpb_out[95][445],u_xpb_out[96][445],u_xpb_out[97][445],u_xpb_out[98][445],u_xpb_out[99][445],u_xpb_out[100][445],u_xpb_out[101][445],u_xpb_out[102][445],u_xpb_out[103][445],u_xpb_out[104][445],u_xpb_out[105][445]};

assign col_out_446 = {u_xpb_out[0][446],u_xpb_out[1][446],u_xpb_out[2][446],u_xpb_out[3][446],u_xpb_out[4][446],u_xpb_out[5][446],u_xpb_out[6][446],u_xpb_out[7][446],u_xpb_out[8][446],u_xpb_out[9][446],u_xpb_out[10][446],u_xpb_out[11][446],u_xpb_out[12][446],u_xpb_out[13][446],u_xpb_out[14][446],u_xpb_out[15][446],u_xpb_out[16][446],u_xpb_out[17][446],u_xpb_out[18][446],u_xpb_out[19][446],u_xpb_out[20][446],u_xpb_out[21][446],u_xpb_out[22][446],u_xpb_out[23][446],u_xpb_out[24][446],u_xpb_out[25][446],u_xpb_out[26][446],u_xpb_out[27][446],u_xpb_out[28][446],u_xpb_out[29][446],u_xpb_out[30][446],u_xpb_out[31][446],u_xpb_out[32][446],u_xpb_out[33][446],u_xpb_out[34][446],u_xpb_out[35][446],u_xpb_out[36][446],u_xpb_out[37][446],u_xpb_out[38][446],u_xpb_out[39][446],u_xpb_out[40][446],u_xpb_out[41][446],u_xpb_out[42][446],u_xpb_out[43][446],u_xpb_out[44][446],u_xpb_out[45][446],u_xpb_out[46][446],u_xpb_out[47][446],u_xpb_out[48][446],u_xpb_out[49][446],u_xpb_out[50][446],u_xpb_out[51][446],u_xpb_out[52][446],u_xpb_out[53][446],u_xpb_out[54][446],u_xpb_out[55][446],u_xpb_out[56][446],u_xpb_out[57][446],u_xpb_out[58][446],u_xpb_out[59][446],u_xpb_out[60][446],u_xpb_out[61][446],u_xpb_out[62][446],u_xpb_out[63][446],u_xpb_out[64][446],u_xpb_out[65][446],u_xpb_out[66][446],u_xpb_out[67][446],u_xpb_out[68][446],u_xpb_out[69][446],u_xpb_out[70][446],u_xpb_out[71][446],u_xpb_out[72][446],u_xpb_out[73][446],u_xpb_out[74][446],u_xpb_out[75][446],u_xpb_out[76][446],u_xpb_out[77][446],u_xpb_out[78][446],u_xpb_out[79][446],u_xpb_out[80][446],u_xpb_out[81][446],u_xpb_out[82][446],u_xpb_out[83][446],u_xpb_out[84][446],u_xpb_out[85][446],u_xpb_out[86][446],u_xpb_out[87][446],u_xpb_out[88][446],u_xpb_out[89][446],u_xpb_out[90][446],u_xpb_out[91][446],u_xpb_out[92][446],u_xpb_out[93][446],u_xpb_out[94][446],u_xpb_out[95][446],u_xpb_out[96][446],u_xpb_out[97][446],u_xpb_out[98][446],u_xpb_out[99][446],u_xpb_out[100][446],u_xpb_out[101][446],u_xpb_out[102][446],u_xpb_out[103][446],u_xpb_out[104][446],u_xpb_out[105][446]};

assign col_out_447 = {u_xpb_out[0][447],u_xpb_out[1][447],u_xpb_out[2][447],u_xpb_out[3][447],u_xpb_out[4][447],u_xpb_out[5][447],u_xpb_out[6][447],u_xpb_out[7][447],u_xpb_out[8][447],u_xpb_out[9][447],u_xpb_out[10][447],u_xpb_out[11][447],u_xpb_out[12][447],u_xpb_out[13][447],u_xpb_out[14][447],u_xpb_out[15][447],u_xpb_out[16][447],u_xpb_out[17][447],u_xpb_out[18][447],u_xpb_out[19][447],u_xpb_out[20][447],u_xpb_out[21][447],u_xpb_out[22][447],u_xpb_out[23][447],u_xpb_out[24][447],u_xpb_out[25][447],u_xpb_out[26][447],u_xpb_out[27][447],u_xpb_out[28][447],u_xpb_out[29][447],u_xpb_out[30][447],u_xpb_out[31][447],u_xpb_out[32][447],u_xpb_out[33][447],u_xpb_out[34][447],u_xpb_out[35][447],u_xpb_out[36][447],u_xpb_out[37][447],u_xpb_out[38][447],u_xpb_out[39][447],u_xpb_out[40][447],u_xpb_out[41][447],u_xpb_out[42][447],u_xpb_out[43][447],u_xpb_out[44][447],u_xpb_out[45][447],u_xpb_out[46][447],u_xpb_out[47][447],u_xpb_out[48][447],u_xpb_out[49][447],u_xpb_out[50][447],u_xpb_out[51][447],u_xpb_out[52][447],u_xpb_out[53][447],u_xpb_out[54][447],u_xpb_out[55][447],u_xpb_out[56][447],u_xpb_out[57][447],u_xpb_out[58][447],u_xpb_out[59][447],u_xpb_out[60][447],u_xpb_out[61][447],u_xpb_out[62][447],u_xpb_out[63][447],u_xpb_out[64][447],u_xpb_out[65][447],u_xpb_out[66][447],u_xpb_out[67][447],u_xpb_out[68][447],u_xpb_out[69][447],u_xpb_out[70][447],u_xpb_out[71][447],u_xpb_out[72][447],u_xpb_out[73][447],u_xpb_out[74][447],u_xpb_out[75][447],u_xpb_out[76][447],u_xpb_out[77][447],u_xpb_out[78][447],u_xpb_out[79][447],u_xpb_out[80][447],u_xpb_out[81][447],u_xpb_out[82][447],u_xpb_out[83][447],u_xpb_out[84][447],u_xpb_out[85][447],u_xpb_out[86][447],u_xpb_out[87][447],u_xpb_out[88][447],u_xpb_out[89][447],u_xpb_out[90][447],u_xpb_out[91][447],u_xpb_out[92][447],u_xpb_out[93][447],u_xpb_out[94][447],u_xpb_out[95][447],u_xpb_out[96][447],u_xpb_out[97][447],u_xpb_out[98][447],u_xpb_out[99][447],u_xpb_out[100][447],u_xpb_out[101][447],u_xpb_out[102][447],u_xpb_out[103][447],u_xpb_out[104][447],u_xpb_out[105][447]};

assign col_out_448 = {u_xpb_out[0][448],u_xpb_out[1][448],u_xpb_out[2][448],u_xpb_out[3][448],u_xpb_out[4][448],u_xpb_out[5][448],u_xpb_out[6][448],u_xpb_out[7][448],u_xpb_out[8][448],u_xpb_out[9][448],u_xpb_out[10][448],u_xpb_out[11][448],u_xpb_out[12][448],u_xpb_out[13][448],u_xpb_out[14][448],u_xpb_out[15][448],u_xpb_out[16][448],u_xpb_out[17][448],u_xpb_out[18][448],u_xpb_out[19][448],u_xpb_out[20][448],u_xpb_out[21][448],u_xpb_out[22][448],u_xpb_out[23][448],u_xpb_out[24][448],u_xpb_out[25][448],u_xpb_out[26][448],u_xpb_out[27][448],u_xpb_out[28][448],u_xpb_out[29][448],u_xpb_out[30][448],u_xpb_out[31][448],u_xpb_out[32][448],u_xpb_out[33][448],u_xpb_out[34][448],u_xpb_out[35][448],u_xpb_out[36][448],u_xpb_out[37][448],u_xpb_out[38][448],u_xpb_out[39][448],u_xpb_out[40][448],u_xpb_out[41][448],u_xpb_out[42][448],u_xpb_out[43][448],u_xpb_out[44][448],u_xpb_out[45][448],u_xpb_out[46][448],u_xpb_out[47][448],u_xpb_out[48][448],u_xpb_out[49][448],u_xpb_out[50][448],u_xpb_out[51][448],u_xpb_out[52][448],u_xpb_out[53][448],u_xpb_out[54][448],u_xpb_out[55][448],u_xpb_out[56][448],u_xpb_out[57][448],u_xpb_out[58][448],u_xpb_out[59][448],u_xpb_out[60][448],u_xpb_out[61][448],u_xpb_out[62][448],u_xpb_out[63][448],u_xpb_out[64][448],u_xpb_out[65][448],u_xpb_out[66][448],u_xpb_out[67][448],u_xpb_out[68][448],u_xpb_out[69][448],u_xpb_out[70][448],u_xpb_out[71][448],u_xpb_out[72][448],u_xpb_out[73][448],u_xpb_out[74][448],u_xpb_out[75][448],u_xpb_out[76][448],u_xpb_out[77][448],u_xpb_out[78][448],u_xpb_out[79][448],u_xpb_out[80][448],u_xpb_out[81][448],u_xpb_out[82][448],u_xpb_out[83][448],u_xpb_out[84][448],u_xpb_out[85][448],u_xpb_out[86][448],u_xpb_out[87][448],u_xpb_out[88][448],u_xpb_out[89][448],u_xpb_out[90][448],u_xpb_out[91][448],u_xpb_out[92][448],u_xpb_out[93][448],u_xpb_out[94][448],u_xpb_out[95][448],u_xpb_out[96][448],u_xpb_out[97][448],u_xpb_out[98][448],u_xpb_out[99][448],u_xpb_out[100][448],u_xpb_out[101][448],u_xpb_out[102][448],u_xpb_out[103][448],u_xpb_out[104][448],u_xpb_out[105][448]};

assign col_out_449 = {u_xpb_out[0][449],u_xpb_out[1][449],u_xpb_out[2][449],u_xpb_out[3][449],u_xpb_out[4][449],u_xpb_out[5][449],u_xpb_out[6][449],u_xpb_out[7][449],u_xpb_out[8][449],u_xpb_out[9][449],u_xpb_out[10][449],u_xpb_out[11][449],u_xpb_out[12][449],u_xpb_out[13][449],u_xpb_out[14][449],u_xpb_out[15][449],u_xpb_out[16][449],u_xpb_out[17][449],u_xpb_out[18][449],u_xpb_out[19][449],u_xpb_out[20][449],u_xpb_out[21][449],u_xpb_out[22][449],u_xpb_out[23][449],u_xpb_out[24][449],u_xpb_out[25][449],u_xpb_out[26][449],u_xpb_out[27][449],u_xpb_out[28][449],u_xpb_out[29][449],u_xpb_out[30][449],u_xpb_out[31][449],u_xpb_out[32][449],u_xpb_out[33][449],u_xpb_out[34][449],u_xpb_out[35][449],u_xpb_out[36][449],u_xpb_out[37][449],u_xpb_out[38][449],u_xpb_out[39][449],u_xpb_out[40][449],u_xpb_out[41][449],u_xpb_out[42][449],u_xpb_out[43][449],u_xpb_out[44][449],u_xpb_out[45][449],u_xpb_out[46][449],u_xpb_out[47][449],u_xpb_out[48][449],u_xpb_out[49][449],u_xpb_out[50][449],u_xpb_out[51][449],u_xpb_out[52][449],u_xpb_out[53][449],u_xpb_out[54][449],u_xpb_out[55][449],u_xpb_out[56][449],u_xpb_out[57][449],u_xpb_out[58][449],u_xpb_out[59][449],u_xpb_out[60][449],u_xpb_out[61][449],u_xpb_out[62][449],u_xpb_out[63][449],u_xpb_out[64][449],u_xpb_out[65][449],u_xpb_out[66][449],u_xpb_out[67][449],u_xpb_out[68][449],u_xpb_out[69][449],u_xpb_out[70][449],u_xpb_out[71][449],u_xpb_out[72][449],u_xpb_out[73][449],u_xpb_out[74][449],u_xpb_out[75][449],u_xpb_out[76][449],u_xpb_out[77][449],u_xpb_out[78][449],u_xpb_out[79][449],u_xpb_out[80][449],u_xpb_out[81][449],u_xpb_out[82][449],u_xpb_out[83][449],u_xpb_out[84][449],u_xpb_out[85][449],u_xpb_out[86][449],u_xpb_out[87][449],u_xpb_out[88][449],u_xpb_out[89][449],u_xpb_out[90][449],u_xpb_out[91][449],u_xpb_out[92][449],u_xpb_out[93][449],u_xpb_out[94][449],u_xpb_out[95][449],u_xpb_out[96][449],u_xpb_out[97][449],u_xpb_out[98][449],u_xpb_out[99][449],u_xpb_out[100][449],u_xpb_out[101][449],u_xpb_out[102][449],u_xpb_out[103][449],u_xpb_out[104][449],u_xpb_out[105][449]};

assign col_out_450 = {u_xpb_out[0][450],u_xpb_out[1][450],u_xpb_out[2][450],u_xpb_out[3][450],u_xpb_out[4][450],u_xpb_out[5][450],u_xpb_out[6][450],u_xpb_out[7][450],u_xpb_out[8][450],u_xpb_out[9][450],u_xpb_out[10][450],u_xpb_out[11][450],u_xpb_out[12][450],u_xpb_out[13][450],u_xpb_out[14][450],u_xpb_out[15][450],u_xpb_out[16][450],u_xpb_out[17][450],u_xpb_out[18][450],u_xpb_out[19][450],u_xpb_out[20][450],u_xpb_out[21][450],u_xpb_out[22][450],u_xpb_out[23][450],u_xpb_out[24][450],u_xpb_out[25][450],u_xpb_out[26][450],u_xpb_out[27][450],u_xpb_out[28][450],u_xpb_out[29][450],u_xpb_out[30][450],u_xpb_out[31][450],u_xpb_out[32][450],u_xpb_out[33][450],u_xpb_out[34][450],u_xpb_out[35][450],u_xpb_out[36][450],u_xpb_out[37][450],u_xpb_out[38][450],u_xpb_out[39][450],u_xpb_out[40][450],u_xpb_out[41][450],u_xpb_out[42][450],u_xpb_out[43][450],u_xpb_out[44][450],u_xpb_out[45][450],u_xpb_out[46][450],u_xpb_out[47][450],u_xpb_out[48][450],u_xpb_out[49][450],u_xpb_out[50][450],u_xpb_out[51][450],u_xpb_out[52][450],u_xpb_out[53][450],u_xpb_out[54][450],u_xpb_out[55][450],u_xpb_out[56][450],u_xpb_out[57][450],u_xpb_out[58][450],u_xpb_out[59][450],u_xpb_out[60][450],u_xpb_out[61][450],u_xpb_out[62][450],u_xpb_out[63][450],u_xpb_out[64][450],u_xpb_out[65][450],u_xpb_out[66][450],u_xpb_out[67][450],u_xpb_out[68][450],u_xpb_out[69][450],u_xpb_out[70][450],u_xpb_out[71][450],u_xpb_out[72][450],u_xpb_out[73][450],u_xpb_out[74][450],u_xpb_out[75][450],u_xpb_out[76][450],u_xpb_out[77][450],u_xpb_out[78][450],u_xpb_out[79][450],u_xpb_out[80][450],u_xpb_out[81][450],u_xpb_out[82][450],u_xpb_out[83][450],u_xpb_out[84][450],u_xpb_out[85][450],u_xpb_out[86][450],u_xpb_out[87][450],u_xpb_out[88][450],u_xpb_out[89][450],u_xpb_out[90][450],u_xpb_out[91][450],u_xpb_out[92][450],u_xpb_out[93][450],u_xpb_out[94][450],u_xpb_out[95][450],u_xpb_out[96][450],u_xpb_out[97][450],u_xpb_out[98][450],u_xpb_out[99][450],u_xpb_out[100][450],u_xpb_out[101][450],u_xpb_out[102][450],u_xpb_out[103][450],u_xpb_out[104][450],u_xpb_out[105][450]};

assign col_out_451 = {u_xpb_out[0][451],u_xpb_out[1][451],u_xpb_out[2][451],u_xpb_out[3][451],u_xpb_out[4][451],u_xpb_out[5][451],u_xpb_out[6][451],u_xpb_out[7][451],u_xpb_out[8][451],u_xpb_out[9][451],u_xpb_out[10][451],u_xpb_out[11][451],u_xpb_out[12][451],u_xpb_out[13][451],u_xpb_out[14][451],u_xpb_out[15][451],u_xpb_out[16][451],u_xpb_out[17][451],u_xpb_out[18][451],u_xpb_out[19][451],u_xpb_out[20][451],u_xpb_out[21][451],u_xpb_out[22][451],u_xpb_out[23][451],u_xpb_out[24][451],u_xpb_out[25][451],u_xpb_out[26][451],u_xpb_out[27][451],u_xpb_out[28][451],u_xpb_out[29][451],u_xpb_out[30][451],u_xpb_out[31][451],u_xpb_out[32][451],u_xpb_out[33][451],u_xpb_out[34][451],u_xpb_out[35][451],u_xpb_out[36][451],u_xpb_out[37][451],u_xpb_out[38][451],u_xpb_out[39][451],u_xpb_out[40][451],u_xpb_out[41][451],u_xpb_out[42][451],u_xpb_out[43][451],u_xpb_out[44][451],u_xpb_out[45][451],u_xpb_out[46][451],u_xpb_out[47][451],u_xpb_out[48][451],u_xpb_out[49][451],u_xpb_out[50][451],u_xpb_out[51][451],u_xpb_out[52][451],u_xpb_out[53][451],u_xpb_out[54][451],u_xpb_out[55][451],u_xpb_out[56][451],u_xpb_out[57][451],u_xpb_out[58][451],u_xpb_out[59][451],u_xpb_out[60][451],u_xpb_out[61][451],u_xpb_out[62][451],u_xpb_out[63][451],u_xpb_out[64][451],u_xpb_out[65][451],u_xpb_out[66][451],u_xpb_out[67][451],u_xpb_out[68][451],u_xpb_out[69][451],u_xpb_out[70][451],u_xpb_out[71][451],u_xpb_out[72][451],u_xpb_out[73][451],u_xpb_out[74][451],u_xpb_out[75][451],u_xpb_out[76][451],u_xpb_out[77][451],u_xpb_out[78][451],u_xpb_out[79][451],u_xpb_out[80][451],u_xpb_out[81][451],u_xpb_out[82][451],u_xpb_out[83][451],u_xpb_out[84][451],u_xpb_out[85][451],u_xpb_out[86][451],u_xpb_out[87][451],u_xpb_out[88][451],u_xpb_out[89][451],u_xpb_out[90][451],u_xpb_out[91][451],u_xpb_out[92][451],u_xpb_out[93][451],u_xpb_out[94][451],u_xpb_out[95][451],u_xpb_out[96][451],u_xpb_out[97][451],u_xpb_out[98][451],u_xpb_out[99][451],u_xpb_out[100][451],u_xpb_out[101][451],u_xpb_out[102][451],u_xpb_out[103][451],u_xpb_out[104][451],u_xpb_out[105][451]};

assign col_out_452 = {u_xpb_out[0][452],u_xpb_out[1][452],u_xpb_out[2][452],u_xpb_out[3][452],u_xpb_out[4][452],u_xpb_out[5][452],u_xpb_out[6][452],u_xpb_out[7][452],u_xpb_out[8][452],u_xpb_out[9][452],u_xpb_out[10][452],u_xpb_out[11][452],u_xpb_out[12][452],u_xpb_out[13][452],u_xpb_out[14][452],u_xpb_out[15][452],u_xpb_out[16][452],u_xpb_out[17][452],u_xpb_out[18][452],u_xpb_out[19][452],u_xpb_out[20][452],u_xpb_out[21][452],u_xpb_out[22][452],u_xpb_out[23][452],u_xpb_out[24][452],u_xpb_out[25][452],u_xpb_out[26][452],u_xpb_out[27][452],u_xpb_out[28][452],u_xpb_out[29][452],u_xpb_out[30][452],u_xpb_out[31][452],u_xpb_out[32][452],u_xpb_out[33][452],u_xpb_out[34][452],u_xpb_out[35][452],u_xpb_out[36][452],u_xpb_out[37][452],u_xpb_out[38][452],u_xpb_out[39][452],u_xpb_out[40][452],u_xpb_out[41][452],u_xpb_out[42][452],u_xpb_out[43][452],u_xpb_out[44][452],u_xpb_out[45][452],u_xpb_out[46][452],u_xpb_out[47][452],u_xpb_out[48][452],u_xpb_out[49][452],u_xpb_out[50][452],u_xpb_out[51][452],u_xpb_out[52][452],u_xpb_out[53][452],u_xpb_out[54][452],u_xpb_out[55][452],u_xpb_out[56][452],u_xpb_out[57][452],u_xpb_out[58][452],u_xpb_out[59][452],u_xpb_out[60][452],u_xpb_out[61][452],u_xpb_out[62][452],u_xpb_out[63][452],u_xpb_out[64][452],u_xpb_out[65][452],u_xpb_out[66][452],u_xpb_out[67][452],u_xpb_out[68][452],u_xpb_out[69][452],u_xpb_out[70][452],u_xpb_out[71][452],u_xpb_out[72][452],u_xpb_out[73][452],u_xpb_out[74][452],u_xpb_out[75][452],u_xpb_out[76][452],u_xpb_out[77][452],u_xpb_out[78][452],u_xpb_out[79][452],u_xpb_out[80][452],u_xpb_out[81][452],u_xpb_out[82][452],u_xpb_out[83][452],u_xpb_out[84][452],u_xpb_out[85][452],u_xpb_out[86][452],u_xpb_out[87][452],u_xpb_out[88][452],u_xpb_out[89][452],u_xpb_out[90][452],u_xpb_out[91][452],u_xpb_out[92][452],u_xpb_out[93][452],u_xpb_out[94][452],u_xpb_out[95][452],u_xpb_out[96][452],u_xpb_out[97][452],u_xpb_out[98][452],u_xpb_out[99][452],u_xpb_out[100][452],u_xpb_out[101][452],u_xpb_out[102][452],u_xpb_out[103][452],u_xpb_out[104][452],u_xpb_out[105][452]};

assign col_out_453 = {u_xpb_out[0][453],u_xpb_out[1][453],u_xpb_out[2][453],u_xpb_out[3][453],u_xpb_out[4][453],u_xpb_out[5][453],u_xpb_out[6][453],u_xpb_out[7][453],u_xpb_out[8][453],u_xpb_out[9][453],u_xpb_out[10][453],u_xpb_out[11][453],u_xpb_out[12][453],u_xpb_out[13][453],u_xpb_out[14][453],u_xpb_out[15][453],u_xpb_out[16][453],u_xpb_out[17][453],u_xpb_out[18][453],u_xpb_out[19][453],u_xpb_out[20][453],u_xpb_out[21][453],u_xpb_out[22][453],u_xpb_out[23][453],u_xpb_out[24][453],u_xpb_out[25][453],u_xpb_out[26][453],u_xpb_out[27][453],u_xpb_out[28][453],u_xpb_out[29][453],u_xpb_out[30][453],u_xpb_out[31][453],u_xpb_out[32][453],u_xpb_out[33][453],u_xpb_out[34][453],u_xpb_out[35][453],u_xpb_out[36][453],u_xpb_out[37][453],u_xpb_out[38][453],u_xpb_out[39][453],u_xpb_out[40][453],u_xpb_out[41][453],u_xpb_out[42][453],u_xpb_out[43][453],u_xpb_out[44][453],u_xpb_out[45][453],u_xpb_out[46][453],u_xpb_out[47][453],u_xpb_out[48][453],u_xpb_out[49][453],u_xpb_out[50][453],u_xpb_out[51][453],u_xpb_out[52][453],u_xpb_out[53][453],u_xpb_out[54][453],u_xpb_out[55][453],u_xpb_out[56][453],u_xpb_out[57][453],u_xpb_out[58][453],u_xpb_out[59][453],u_xpb_out[60][453],u_xpb_out[61][453],u_xpb_out[62][453],u_xpb_out[63][453],u_xpb_out[64][453],u_xpb_out[65][453],u_xpb_out[66][453],u_xpb_out[67][453],u_xpb_out[68][453],u_xpb_out[69][453],u_xpb_out[70][453],u_xpb_out[71][453],u_xpb_out[72][453],u_xpb_out[73][453],u_xpb_out[74][453],u_xpb_out[75][453],u_xpb_out[76][453],u_xpb_out[77][453],u_xpb_out[78][453],u_xpb_out[79][453],u_xpb_out[80][453],u_xpb_out[81][453],u_xpb_out[82][453],u_xpb_out[83][453],u_xpb_out[84][453],u_xpb_out[85][453],u_xpb_out[86][453],u_xpb_out[87][453],u_xpb_out[88][453],u_xpb_out[89][453],u_xpb_out[90][453],u_xpb_out[91][453],u_xpb_out[92][453],u_xpb_out[93][453],u_xpb_out[94][453],u_xpb_out[95][453],u_xpb_out[96][453],u_xpb_out[97][453],u_xpb_out[98][453],u_xpb_out[99][453],u_xpb_out[100][453],u_xpb_out[101][453],u_xpb_out[102][453],u_xpb_out[103][453],u_xpb_out[104][453],u_xpb_out[105][453]};

assign col_out_454 = {u_xpb_out[0][454],u_xpb_out[1][454],u_xpb_out[2][454],u_xpb_out[3][454],u_xpb_out[4][454],u_xpb_out[5][454],u_xpb_out[6][454],u_xpb_out[7][454],u_xpb_out[8][454],u_xpb_out[9][454],u_xpb_out[10][454],u_xpb_out[11][454],u_xpb_out[12][454],u_xpb_out[13][454],u_xpb_out[14][454],u_xpb_out[15][454],u_xpb_out[16][454],u_xpb_out[17][454],u_xpb_out[18][454],u_xpb_out[19][454],u_xpb_out[20][454],u_xpb_out[21][454],u_xpb_out[22][454],u_xpb_out[23][454],u_xpb_out[24][454],u_xpb_out[25][454],u_xpb_out[26][454],u_xpb_out[27][454],u_xpb_out[28][454],u_xpb_out[29][454],u_xpb_out[30][454],u_xpb_out[31][454],u_xpb_out[32][454],u_xpb_out[33][454],u_xpb_out[34][454],u_xpb_out[35][454],u_xpb_out[36][454],u_xpb_out[37][454],u_xpb_out[38][454],u_xpb_out[39][454],u_xpb_out[40][454],u_xpb_out[41][454],u_xpb_out[42][454],u_xpb_out[43][454],u_xpb_out[44][454],u_xpb_out[45][454],u_xpb_out[46][454],u_xpb_out[47][454],u_xpb_out[48][454],u_xpb_out[49][454],u_xpb_out[50][454],u_xpb_out[51][454],u_xpb_out[52][454],u_xpb_out[53][454],u_xpb_out[54][454],u_xpb_out[55][454],u_xpb_out[56][454],u_xpb_out[57][454],u_xpb_out[58][454],u_xpb_out[59][454],u_xpb_out[60][454],u_xpb_out[61][454],u_xpb_out[62][454],u_xpb_out[63][454],u_xpb_out[64][454],u_xpb_out[65][454],u_xpb_out[66][454],u_xpb_out[67][454],u_xpb_out[68][454],u_xpb_out[69][454],u_xpb_out[70][454],u_xpb_out[71][454],u_xpb_out[72][454],u_xpb_out[73][454],u_xpb_out[74][454],u_xpb_out[75][454],u_xpb_out[76][454],u_xpb_out[77][454],u_xpb_out[78][454],u_xpb_out[79][454],u_xpb_out[80][454],u_xpb_out[81][454],u_xpb_out[82][454],u_xpb_out[83][454],u_xpb_out[84][454],u_xpb_out[85][454],u_xpb_out[86][454],u_xpb_out[87][454],u_xpb_out[88][454],u_xpb_out[89][454],u_xpb_out[90][454],u_xpb_out[91][454],u_xpb_out[92][454],u_xpb_out[93][454],u_xpb_out[94][454],u_xpb_out[95][454],u_xpb_out[96][454],u_xpb_out[97][454],u_xpb_out[98][454],u_xpb_out[99][454],u_xpb_out[100][454],u_xpb_out[101][454],u_xpb_out[102][454],u_xpb_out[103][454],u_xpb_out[104][454],u_xpb_out[105][454]};

assign col_out_455 = {u_xpb_out[0][455],u_xpb_out[1][455],u_xpb_out[2][455],u_xpb_out[3][455],u_xpb_out[4][455],u_xpb_out[5][455],u_xpb_out[6][455],u_xpb_out[7][455],u_xpb_out[8][455],u_xpb_out[9][455],u_xpb_out[10][455],u_xpb_out[11][455],u_xpb_out[12][455],u_xpb_out[13][455],u_xpb_out[14][455],u_xpb_out[15][455],u_xpb_out[16][455],u_xpb_out[17][455],u_xpb_out[18][455],u_xpb_out[19][455],u_xpb_out[20][455],u_xpb_out[21][455],u_xpb_out[22][455],u_xpb_out[23][455],u_xpb_out[24][455],u_xpb_out[25][455],u_xpb_out[26][455],u_xpb_out[27][455],u_xpb_out[28][455],u_xpb_out[29][455],u_xpb_out[30][455],u_xpb_out[31][455],u_xpb_out[32][455],u_xpb_out[33][455],u_xpb_out[34][455],u_xpb_out[35][455],u_xpb_out[36][455],u_xpb_out[37][455],u_xpb_out[38][455],u_xpb_out[39][455],u_xpb_out[40][455],u_xpb_out[41][455],u_xpb_out[42][455],u_xpb_out[43][455],u_xpb_out[44][455],u_xpb_out[45][455],u_xpb_out[46][455],u_xpb_out[47][455],u_xpb_out[48][455],u_xpb_out[49][455],u_xpb_out[50][455],u_xpb_out[51][455],u_xpb_out[52][455],u_xpb_out[53][455],u_xpb_out[54][455],u_xpb_out[55][455],u_xpb_out[56][455],u_xpb_out[57][455],u_xpb_out[58][455],u_xpb_out[59][455],u_xpb_out[60][455],u_xpb_out[61][455],u_xpb_out[62][455],u_xpb_out[63][455],u_xpb_out[64][455],u_xpb_out[65][455],u_xpb_out[66][455],u_xpb_out[67][455],u_xpb_out[68][455],u_xpb_out[69][455],u_xpb_out[70][455],u_xpb_out[71][455],u_xpb_out[72][455],u_xpb_out[73][455],u_xpb_out[74][455],u_xpb_out[75][455],u_xpb_out[76][455],u_xpb_out[77][455],u_xpb_out[78][455],u_xpb_out[79][455],u_xpb_out[80][455],u_xpb_out[81][455],u_xpb_out[82][455],u_xpb_out[83][455],u_xpb_out[84][455],u_xpb_out[85][455],u_xpb_out[86][455],u_xpb_out[87][455],u_xpb_out[88][455],u_xpb_out[89][455],u_xpb_out[90][455],u_xpb_out[91][455],u_xpb_out[92][455],u_xpb_out[93][455],u_xpb_out[94][455],u_xpb_out[95][455],u_xpb_out[96][455],u_xpb_out[97][455],u_xpb_out[98][455],u_xpb_out[99][455],u_xpb_out[100][455],u_xpb_out[101][455],u_xpb_out[102][455],u_xpb_out[103][455],u_xpb_out[104][455],u_xpb_out[105][455]};

assign col_out_456 = {u_xpb_out[0][456],u_xpb_out[1][456],u_xpb_out[2][456],u_xpb_out[3][456],u_xpb_out[4][456],u_xpb_out[5][456],u_xpb_out[6][456],u_xpb_out[7][456],u_xpb_out[8][456],u_xpb_out[9][456],u_xpb_out[10][456],u_xpb_out[11][456],u_xpb_out[12][456],u_xpb_out[13][456],u_xpb_out[14][456],u_xpb_out[15][456],u_xpb_out[16][456],u_xpb_out[17][456],u_xpb_out[18][456],u_xpb_out[19][456],u_xpb_out[20][456],u_xpb_out[21][456],u_xpb_out[22][456],u_xpb_out[23][456],u_xpb_out[24][456],u_xpb_out[25][456],u_xpb_out[26][456],u_xpb_out[27][456],u_xpb_out[28][456],u_xpb_out[29][456],u_xpb_out[30][456],u_xpb_out[31][456],u_xpb_out[32][456],u_xpb_out[33][456],u_xpb_out[34][456],u_xpb_out[35][456],u_xpb_out[36][456],u_xpb_out[37][456],u_xpb_out[38][456],u_xpb_out[39][456],u_xpb_out[40][456],u_xpb_out[41][456],u_xpb_out[42][456],u_xpb_out[43][456],u_xpb_out[44][456],u_xpb_out[45][456],u_xpb_out[46][456],u_xpb_out[47][456],u_xpb_out[48][456],u_xpb_out[49][456],u_xpb_out[50][456],u_xpb_out[51][456],u_xpb_out[52][456],u_xpb_out[53][456],u_xpb_out[54][456],u_xpb_out[55][456],u_xpb_out[56][456],u_xpb_out[57][456],u_xpb_out[58][456],u_xpb_out[59][456],u_xpb_out[60][456],u_xpb_out[61][456],u_xpb_out[62][456],u_xpb_out[63][456],u_xpb_out[64][456],u_xpb_out[65][456],u_xpb_out[66][456],u_xpb_out[67][456],u_xpb_out[68][456],u_xpb_out[69][456],u_xpb_out[70][456],u_xpb_out[71][456],u_xpb_out[72][456],u_xpb_out[73][456],u_xpb_out[74][456],u_xpb_out[75][456],u_xpb_out[76][456],u_xpb_out[77][456],u_xpb_out[78][456],u_xpb_out[79][456],u_xpb_out[80][456],u_xpb_out[81][456],u_xpb_out[82][456],u_xpb_out[83][456],u_xpb_out[84][456],u_xpb_out[85][456],u_xpb_out[86][456],u_xpb_out[87][456],u_xpb_out[88][456],u_xpb_out[89][456],u_xpb_out[90][456],u_xpb_out[91][456],u_xpb_out[92][456],u_xpb_out[93][456],u_xpb_out[94][456],u_xpb_out[95][456],u_xpb_out[96][456],u_xpb_out[97][456],u_xpb_out[98][456],u_xpb_out[99][456],u_xpb_out[100][456],u_xpb_out[101][456],u_xpb_out[102][456],u_xpb_out[103][456],u_xpb_out[104][456],u_xpb_out[105][456]};

assign col_out_457 = {u_xpb_out[0][457],u_xpb_out[1][457],u_xpb_out[2][457],u_xpb_out[3][457],u_xpb_out[4][457],u_xpb_out[5][457],u_xpb_out[6][457],u_xpb_out[7][457],u_xpb_out[8][457],u_xpb_out[9][457],u_xpb_out[10][457],u_xpb_out[11][457],u_xpb_out[12][457],u_xpb_out[13][457],u_xpb_out[14][457],u_xpb_out[15][457],u_xpb_out[16][457],u_xpb_out[17][457],u_xpb_out[18][457],u_xpb_out[19][457],u_xpb_out[20][457],u_xpb_out[21][457],u_xpb_out[22][457],u_xpb_out[23][457],u_xpb_out[24][457],u_xpb_out[25][457],u_xpb_out[26][457],u_xpb_out[27][457],u_xpb_out[28][457],u_xpb_out[29][457],u_xpb_out[30][457],u_xpb_out[31][457],u_xpb_out[32][457],u_xpb_out[33][457],u_xpb_out[34][457],u_xpb_out[35][457],u_xpb_out[36][457],u_xpb_out[37][457],u_xpb_out[38][457],u_xpb_out[39][457],u_xpb_out[40][457],u_xpb_out[41][457],u_xpb_out[42][457],u_xpb_out[43][457],u_xpb_out[44][457],u_xpb_out[45][457],u_xpb_out[46][457],u_xpb_out[47][457],u_xpb_out[48][457],u_xpb_out[49][457],u_xpb_out[50][457],u_xpb_out[51][457],u_xpb_out[52][457],u_xpb_out[53][457],u_xpb_out[54][457],u_xpb_out[55][457],u_xpb_out[56][457],u_xpb_out[57][457],u_xpb_out[58][457],u_xpb_out[59][457],u_xpb_out[60][457],u_xpb_out[61][457],u_xpb_out[62][457],u_xpb_out[63][457],u_xpb_out[64][457],u_xpb_out[65][457],u_xpb_out[66][457],u_xpb_out[67][457],u_xpb_out[68][457],u_xpb_out[69][457],u_xpb_out[70][457],u_xpb_out[71][457],u_xpb_out[72][457],u_xpb_out[73][457],u_xpb_out[74][457],u_xpb_out[75][457],u_xpb_out[76][457],u_xpb_out[77][457],u_xpb_out[78][457],u_xpb_out[79][457],u_xpb_out[80][457],u_xpb_out[81][457],u_xpb_out[82][457],u_xpb_out[83][457],u_xpb_out[84][457],u_xpb_out[85][457],u_xpb_out[86][457],u_xpb_out[87][457],u_xpb_out[88][457],u_xpb_out[89][457],u_xpb_out[90][457],u_xpb_out[91][457],u_xpb_out[92][457],u_xpb_out[93][457],u_xpb_out[94][457],u_xpb_out[95][457],u_xpb_out[96][457],u_xpb_out[97][457],u_xpb_out[98][457],u_xpb_out[99][457],u_xpb_out[100][457],u_xpb_out[101][457],u_xpb_out[102][457],u_xpb_out[103][457],u_xpb_out[104][457],u_xpb_out[105][457]};

assign col_out_458 = {u_xpb_out[0][458],u_xpb_out[1][458],u_xpb_out[2][458],u_xpb_out[3][458],u_xpb_out[4][458],u_xpb_out[5][458],u_xpb_out[6][458],u_xpb_out[7][458],u_xpb_out[8][458],u_xpb_out[9][458],u_xpb_out[10][458],u_xpb_out[11][458],u_xpb_out[12][458],u_xpb_out[13][458],u_xpb_out[14][458],u_xpb_out[15][458],u_xpb_out[16][458],u_xpb_out[17][458],u_xpb_out[18][458],u_xpb_out[19][458],u_xpb_out[20][458],u_xpb_out[21][458],u_xpb_out[22][458],u_xpb_out[23][458],u_xpb_out[24][458],u_xpb_out[25][458],u_xpb_out[26][458],u_xpb_out[27][458],u_xpb_out[28][458],u_xpb_out[29][458],u_xpb_out[30][458],u_xpb_out[31][458],u_xpb_out[32][458],u_xpb_out[33][458],u_xpb_out[34][458],u_xpb_out[35][458],u_xpb_out[36][458],u_xpb_out[37][458],u_xpb_out[38][458],u_xpb_out[39][458],u_xpb_out[40][458],u_xpb_out[41][458],u_xpb_out[42][458],u_xpb_out[43][458],u_xpb_out[44][458],u_xpb_out[45][458],u_xpb_out[46][458],u_xpb_out[47][458],u_xpb_out[48][458],u_xpb_out[49][458],u_xpb_out[50][458],u_xpb_out[51][458],u_xpb_out[52][458],u_xpb_out[53][458],u_xpb_out[54][458],u_xpb_out[55][458],u_xpb_out[56][458],u_xpb_out[57][458],u_xpb_out[58][458],u_xpb_out[59][458],u_xpb_out[60][458],u_xpb_out[61][458],u_xpb_out[62][458],u_xpb_out[63][458],u_xpb_out[64][458],u_xpb_out[65][458],u_xpb_out[66][458],u_xpb_out[67][458],u_xpb_out[68][458],u_xpb_out[69][458],u_xpb_out[70][458],u_xpb_out[71][458],u_xpb_out[72][458],u_xpb_out[73][458],u_xpb_out[74][458],u_xpb_out[75][458],u_xpb_out[76][458],u_xpb_out[77][458],u_xpb_out[78][458],u_xpb_out[79][458],u_xpb_out[80][458],u_xpb_out[81][458],u_xpb_out[82][458],u_xpb_out[83][458],u_xpb_out[84][458],u_xpb_out[85][458],u_xpb_out[86][458],u_xpb_out[87][458],u_xpb_out[88][458],u_xpb_out[89][458],u_xpb_out[90][458],u_xpb_out[91][458],u_xpb_out[92][458],u_xpb_out[93][458],u_xpb_out[94][458],u_xpb_out[95][458],u_xpb_out[96][458],u_xpb_out[97][458],u_xpb_out[98][458],u_xpb_out[99][458],u_xpb_out[100][458],u_xpb_out[101][458],u_xpb_out[102][458],u_xpb_out[103][458],u_xpb_out[104][458],u_xpb_out[105][458]};

assign col_out_459 = {u_xpb_out[0][459],u_xpb_out[1][459],u_xpb_out[2][459],u_xpb_out[3][459],u_xpb_out[4][459],u_xpb_out[5][459],u_xpb_out[6][459],u_xpb_out[7][459],u_xpb_out[8][459],u_xpb_out[9][459],u_xpb_out[10][459],u_xpb_out[11][459],u_xpb_out[12][459],u_xpb_out[13][459],u_xpb_out[14][459],u_xpb_out[15][459],u_xpb_out[16][459],u_xpb_out[17][459],u_xpb_out[18][459],u_xpb_out[19][459],u_xpb_out[20][459],u_xpb_out[21][459],u_xpb_out[22][459],u_xpb_out[23][459],u_xpb_out[24][459],u_xpb_out[25][459],u_xpb_out[26][459],u_xpb_out[27][459],u_xpb_out[28][459],u_xpb_out[29][459],u_xpb_out[30][459],u_xpb_out[31][459],u_xpb_out[32][459],u_xpb_out[33][459],u_xpb_out[34][459],u_xpb_out[35][459],u_xpb_out[36][459],u_xpb_out[37][459],u_xpb_out[38][459],u_xpb_out[39][459],u_xpb_out[40][459],u_xpb_out[41][459],u_xpb_out[42][459],u_xpb_out[43][459],u_xpb_out[44][459],u_xpb_out[45][459],u_xpb_out[46][459],u_xpb_out[47][459],u_xpb_out[48][459],u_xpb_out[49][459],u_xpb_out[50][459],u_xpb_out[51][459],u_xpb_out[52][459],u_xpb_out[53][459],u_xpb_out[54][459],u_xpb_out[55][459],u_xpb_out[56][459],u_xpb_out[57][459],u_xpb_out[58][459],u_xpb_out[59][459],u_xpb_out[60][459],u_xpb_out[61][459],u_xpb_out[62][459],u_xpb_out[63][459],u_xpb_out[64][459],u_xpb_out[65][459],u_xpb_out[66][459],u_xpb_out[67][459],u_xpb_out[68][459],u_xpb_out[69][459],u_xpb_out[70][459],u_xpb_out[71][459],u_xpb_out[72][459],u_xpb_out[73][459],u_xpb_out[74][459],u_xpb_out[75][459],u_xpb_out[76][459],u_xpb_out[77][459],u_xpb_out[78][459],u_xpb_out[79][459],u_xpb_out[80][459],u_xpb_out[81][459],u_xpb_out[82][459],u_xpb_out[83][459],u_xpb_out[84][459],u_xpb_out[85][459],u_xpb_out[86][459],u_xpb_out[87][459],u_xpb_out[88][459],u_xpb_out[89][459],u_xpb_out[90][459],u_xpb_out[91][459],u_xpb_out[92][459],u_xpb_out[93][459],u_xpb_out[94][459],u_xpb_out[95][459],u_xpb_out[96][459],u_xpb_out[97][459],u_xpb_out[98][459],u_xpb_out[99][459],u_xpb_out[100][459],u_xpb_out[101][459],u_xpb_out[102][459],u_xpb_out[103][459],u_xpb_out[104][459],u_xpb_out[105][459]};

assign col_out_460 = {u_xpb_out[0][460],u_xpb_out[1][460],u_xpb_out[2][460],u_xpb_out[3][460],u_xpb_out[4][460],u_xpb_out[5][460],u_xpb_out[6][460],u_xpb_out[7][460],u_xpb_out[8][460],u_xpb_out[9][460],u_xpb_out[10][460],u_xpb_out[11][460],u_xpb_out[12][460],u_xpb_out[13][460],u_xpb_out[14][460],u_xpb_out[15][460],u_xpb_out[16][460],u_xpb_out[17][460],u_xpb_out[18][460],u_xpb_out[19][460],u_xpb_out[20][460],u_xpb_out[21][460],u_xpb_out[22][460],u_xpb_out[23][460],u_xpb_out[24][460],u_xpb_out[25][460],u_xpb_out[26][460],u_xpb_out[27][460],u_xpb_out[28][460],u_xpb_out[29][460],u_xpb_out[30][460],u_xpb_out[31][460],u_xpb_out[32][460],u_xpb_out[33][460],u_xpb_out[34][460],u_xpb_out[35][460],u_xpb_out[36][460],u_xpb_out[37][460],u_xpb_out[38][460],u_xpb_out[39][460],u_xpb_out[40][460],u_xpb_out[41][460],u_xpb_out[42][460],u_xpb_out[43][460],u_xpb_out[44][460],u_xpb_out[45][460],u_xpb_out[46][460],u_xpb_out[47][460],u_xpb_out[48][460],u_xpb_out[49][460],u_xpb_out[50][460],u_xpb_out[51][460],u_xpb_out[52][460],u_xpb_out[53][460],u_xpb_out[54][460],u_xpb_out[55][460],u_xpb_out[56][460],u_xpb_out[57][460],u_xpb_out[58][460],u_xpb_out[59][460],u_xpb_out[60][460],u_xpb_out[61][460],u_xpb_out[62][460],u_xpb_out[63][460],u_xpb_out[64][460],u_xpb_out[65][460],u_xpb_out[66][460],u_xpb_out[67][460],u_xpb_out[68][460],u_xpb_out[69][460],u_xpb_out[70][460],u_xpb_out[71][460],u_xpb_out[72][460],u_xpb_out[73][460],u_xpb_out[74][460],u_xpb_out[75][460],u_xpb_out[76][460],u_xpb_out[77][460],u_xpb_out[78][460],u_xpb_out[79][460],u_xpb_out[80][460],u_xpb_out[81][460],u_xpb_out[82][460],u_xpb_out[83][460],u_xpb_out[84][460],u_xpb_out[85][460],u_xpb_out[86][460],u_xpb_out[87][460],u_xpb_out[88][460],u_xpb_out[89][460],u_xpb_out[90][460],u_xpb_out[91][460],u_xpb_out[92][460],u_xpb_out[93][460],u_xpb_out[94][460],u_xpb_out[95][460],u_xpb_out[96][460],u_xpb_out[97][460],u_xpb_out[98][460],u_xpb_out[99][460],u_xpb_out[100][460],u_xpb_out[101][460],u_xpb_out[102][460],u_xpb_out[103][460],u_xpb_out[104][460],u_xpb_out[105][460]};

assign col_out_461 = {u_xpb_out[0][461],u_xpb_out[1][461],u_xpb_out[2][461],u_xpb_out[3][461],u_xpb_out[4][461],u_xpb_out[5][461],u_xpb_out[6][461],u_xpb_out[7][461],u_xpb_out[8][461],u_xpb_out[9][461],u_xpb_out[10][461],u_xpb_out[11][461],u_xpb_out[12][461],u_xpb_out[13][461],u_xpb_out[14][461],u_xpb_out[15][461],u_xpb_out[16][461],u_xpb_out[17][461],u_xpb_out[18][461],u_xpb_out[19][461],u_xpb_out[20][461],u_xpb_out[21][461],u_xpb_out[22][461],u_xpb_out[23][461],u_xpb_out[24][461],u_xpb_out[25][461],u_xpb_out[26][461],u_xpb_out[27][461],u_xpb_out[28][461],u_xpb_out[29][461],u_xpb_out[30][461],u_xpb_out[31][461],u_xpb_out[32][461],u_xpb_out[33][461],u_xpb_out[34][461],u_xpb_out[35][461],u_xpb_out[36][461],u_xpb_out[37][461],u_xpb_out[38][461],u_xpb_out[39][461],u_xpb_out[40][461],u_xpb_out[41][461],u_xpb_out[42][461],u_xpb_out[43][461],u_xpb_out[44][461],u_xpb_out[45][461],u_xpb_out[46][461],u_xpb_out[47][461],u_xpb_out[48][461],u_xpb_out[49][461],u_xpb_out[50][461],u_xpb_out[51][461],u_xpb_out[52][461],u_xpb_out[53][461],u_xpb_out[54][461],u_xpb_out[55][461],u_xpb_out[56][461],u_xpb_out[57][461],u_xpb_out[58][461],u_xpb_out[59][461],u_xpb_out[60][461],u_xpb_out[61][461],u_xpb_out[62][461],u_xpb_out[63][461],u_xpb_out[64][461],u_xpb_out[65][461],u_xpb_out[66][461],u_xpb_out[67][461],u_xpb_out[68][461],u_xpb_out[69][461],u_xpb_out[70][461],u_xpb_out[71][461],u_xpb_out[72][461],u_xpb_out[73][461],u_xpb_out[74][461],u_xpb_out[75][461],u_xpb_out[76][461],u_xpb_out[77][461],u_xpb_out[78][461],u_xpb_out[79][461],u_xpb_out[80][461],u_xpb_out[81][461],u_xpb_out[82][461],u_xpb_out[83][461],u_xpb_out[84][461],u_xpb_out[85][461],u_xpb_out[86][461],u_xpb_out[87][461],u_xpb_out[88][461],u_xpb_out[89][461],u_xpb_out[90][461],u_xpb_out[91][461],u_xpb_out[92][461],u_xpb_out[93][461],u_xpb_out[94][461],u_xpb_out[95][461],u_xpb_out[96][461],u_xpb_out[97][461],u_xpb_out[98][461],u_xpb_out[99][461],u_xpb_out[100][461],u_xpb_out[101][461],u_xpb_out[102][461],u_xpb_out[103][461],u_xpb_out[104][461],u_xpb_out[105][461]};

assign col_out_462 = {u_xpb_out[0][462],u_xpb_out[1][462],u_xpb_out[2][462],u_xpb_out[3][462],u_xpb_out[4][462],u_xpb_out[5][462],u_xpb_out[6][462],u_xpb_out[7][462],u_xpb_out[8][462],u_xpb_out[9][462],u_xpb_out[10][462],u_xpb_out[11][462],u_xpb_out[12][462],u_xpb_out[13][462],u_xpb_out[14][462],u_xpb_out[15][462],u_xpb_out[16][462],u_xpb_out[17][462],u_xpb_out[18][462],u_xpb_out[19][462],u_xpb_out[20][462],u_xpb_out[21][462],u_xpb_out[22][462],u_xpb_out[23][462],u_xpb_out[24][462],u_xpb_out[25][462],u_xpb_out[26][462],u_xpb_out[27][462],u_xpb_out[28][462],u_xpb_out[29][462],u_xpb_out[30][462],u_xpb_out[31][462],u_xpb_out[32][462],u_xpb_out[33][462],u_xpb_out[34][462],u_xpb_out[35][462],u_xpb_out[36][462],u_xpb_out[37][462],u_xpb_out[38][462],u_xpb_out[39][462],u_xpb_out[40][462],u_xpb_out[41][462],u_xpb_out[42][462],u_xpb_out[43][462],u_xpb_out[44][462],u_xpb_out[45][462],u_xpb_out[46][462],u_xpb_out[47][462],u_xpb_out[48][462],u_xpb_out[49][462],u_xpb_out[50][462],u_xpb_out[51][462],u_xpb_out[52][462],u_xpb_out[53][462],u_xpb_out[54][462],u_xpb_out[55][462],u_xpb_out[56][462],u_xpb_out[57][462],u_xpb_out[58][462],u_xpb_out[59][462],u_xpb_out[60][462],u_xpb_out[61][462],u_xpb_out[62][462],u_xpb_out[63][462],u_xpb_out[64][462],u_xpb_out[65][462],u_xpb_out[66][462],u_xpb_out[67][462],u_xpb_out[68][462],u_xpb_out[69][462],u_xpb_out[70][462],u_xpb_out[71][462],u_xpb_out[72][462],u_xpb_out[73][462],u_xpb_out[74][462],u_xpb_out[75][462],u_xpb_out[76][462],u_xpb_out[77][462],u_xpb_out[78][462],u_xpb_out[79][462],u_xpb_out[80][462],u_xpb_out[81][462],u_xpb_out[82][462],u_xpb_out[83][462],u_xpb_out[84][462],u_xpb_out[85][462],u_xpb_out[86][462],u_xpb_out[87][462],u_xpb_out[88][462],u_xpb_out[89][462],u_xpb_out[90][462],u_xpb_out[91][462],u_xpb_out[92][462],u_xpb_out[93][462],u_xpb_out[94][462],u_xpb_out[95][462],u_xpb_out[96][462],u_xpb_out[97][462],u_xpb_out[98][462],u_xpb_out[99][462],u_xpb_out[100][462],u_xpb_out[101][462],u_xpb_out[102][462],u_xpb_out[103][462],u_xpb_out[104][462],u_xpb_out[105][462]};

assign col_out_463 = {u_xpb_out[0][463],u_xpb_out[1][463],u_xpb_out[2][463],u_xpb_out[3][463],u_xpb_out[4][463],u_xpb_out[5][463],u_xpb_out[6][463],u_xpb_out[7][463],u_xpb_out[8][463],u_xpb_out[9][463],u_xpb_out[10][463],u_xpb_out[11][463],u_xpb_out[12][463],u_xpb_out[13][463],u_xpb_out[14][463],u_xpb_out[15][463],u_xpb_out[16][463],u_xpb_out[17][463],u_xpb_out[18][463],u_xpb_out[19][463],u_xpb_out[20][463],u_xpb_out[21][463],u_xpb_out[22][463],u_xpb_out[23][463],u_xpb_out[24][463],u_xpb_out[25][463],u_xpb_out[26][463],u_xpb_out[27][463],u_xpb_out[28][463],u_xpb_out[29][463],u_xpb_out[30][463],u_xpb_out[31][463],u_xpb_out[32][463],u_xpb_out[33][463],u_xpb_out[34][463],u_xpb_out[35][463],u_xpb_out[36][463],u_xpb_out[37][463],u_xpb_out[38][463],u_xpb_out[39][463],u_xpb_out[40][463],u_xpb_out[41][463],u_xpb_out[42][463],u_xpb_out[43][463],u_xpb_out[44][463],u_xpb_out[45][463],u_xpb_out[46][463],u_xpb_out[47][463],u_xpb_out[48][463],u_xpb_out[49][463],u_xpb_out[50][463],u_xpb_out[51][463],u_xpb_out[52][463],u_xpb_out[53][463],u_xpb_out[54][463],u_xpb_out[55][463],u_xpb_out[56][463],u_xpb_out[57][463],u_xpb_out[58][463],u_xpb_out[59][463],u_xpb_out[60][463],u_xpb_out[61][463],u_xpb_out[62][463],u_xpb_out[63][463],u_xpb_out[64][463],u_xpb_out[65][463],u_xpb_out[66][463],u_xpb_out[67][463],u_xpb_out[68][463],u_xpb_out[69][463],u_xpb_out[70][463],u_xpb_out[71][463],u_xpb_out[72][463],u_xpb_out[73][463],u_xpb_out[74][463],u_xpb_out[75][463],u_xpb_out[76][463],u_xpb_out[77][463],u_xpb_out[78][463],u_xpb_out[79][463],u_xpb_out[80][463],u_xpb_out[81][463],u_xpb_out[82][463],u_xpb_out[83][463],u_xpb_out[84][463],u_xpb_out[85][463],u_xpb_out[86][463],u_xpb_out[87][463],u_xpb_out[88][463],u_xpb_out[89][463],u_xpb_out[90][463],u_xpb_out[91][463],u_xpb_out[92][463],u_xpb_out[93][463],u_xpb_out[94][463],u_xpb_out[95][463],u_xpb_out[96][463],u_xpb_out[97][463],u_xpb_out[98][463],u_xpb_out[99][463],u_xpb_out[100][463],u_xpb_out[101][463],u_xpb_out[102][463],u_xpb_out[103][463],u_xpb_out[104][463],u_xpb_out[105][463]};

assign col_out_464 = {u_xpb_out[0][464],u_xpb_out[1][464],u_xpb_out[2][464],u_xpb_out[3][464],u_xpb_out[4][464],u_xpb_out[5][464],u_xpb_out[6][464],u_xpb_out[7][464],u_xpb_out[8][464],u_xpb_out[9][464],u_xpb_out[10][464],u_xpb_out[11][464],u_xpb_out[12][464],u_xpb_out[13][464],u_xpb_out[14][464],u_xpb_out[15][464],u_xpb_out[16][464],u_xpb_out[17][464],u_xpb_out[18][464],u_xpb_out[19][464],u_xpb_out[20][464],u_xpb_out[21][464],u_xpb_out[22][464],u_xpb_out[23][464],u_xpb_out[24][464],u_xpb_out[25][464],u_xpb_out[26][464],u_xpb_out[27][464],u_xpb_out[28][464],u_xpb_out[29][464],u_xpb_out[30][464],u_xpb_out[31][464],u_xpb_out[32][464],u_xpb_out[33][464],u_xpb_out[34][464],u_xpb_out[35][464],u_xpb_out[36][464],u_xpb_out[37][464],u_xpb_out[38][464],u_xpb_out[39][464],u_xpb_out[40][464],u_xpb_out[41][464],u_xpb_out[42][464],u_xpb_out[43][464],u_xpb_out[44][464],u_xpb_out[45][464],u_xpb_out[46][464],u_xpb_out[47][464],u_xpb_out[48][464],u_xpb_out[49][464],u_xpb_out[50][464],u_xpb_out[51][464],u_xpb_out[52][464],u_xpb_out[53][464],u_xpb_out[54][464],u_xpb_out[55][464],u_xpb_out[56][464],u_xpb_out[57][464],u_xpb_out[58][464],u_xpb_out[59][464],u_xpb_out[60][464],u_xpb_out[61][464],u_xpb_out[62][464],u_xpb_out[63][464],u_xpb_out[64][464],u_xpb_out[65][464],u_xpb_out[66][464],u_xpb_out[67][464],u_xpb_out[68][464],u_xpb_out[69][464],u_xpb_out[70][464],u_xpb_out[71][464],u_xpb_out[72][464],u_xpb_out[73][464],u_xpb_out[74][464],u_xpb_out[75][464],u_xpb_out[76][464],u_xpb_out[77][464],u_xpb_out[78][464],u_xpb_out[79][464],u_xpb_out[80][464],u_xpb_out[81][464],u_xpb_out[82][464],u_xpb_out[83][464],u_xpb_out[84][464],u_xpb_out[85][464],u_xpb_out[86][464],u_xpb_out[87][464],u_xpb_out[88][464],u_xpb_out[89][464],u_xpb_out[90][464],u_xpb_out[91][464],u_xpb_out[92][464],u_xpb_out[93][464],u_xpb_out[94][464],u_xpb_out[95][464],u_xpb_out[96][464],u_xpb_out[97][464],u_xpb_out[98][464],u_xpb_out[99][464],u_xpb_out[100][464],u_xpb_out[101][464],u_xpb_out[102][464],u_xpb_out[103][464],u_xpb_out[104][464],u_xpb_out[105][464]};

assign col_out_465 = {u_xpb_out[0][465],u_xpb_out[1][465],u_xpb_out[2][465],u_xpb_out[3][465],u_xpb_out[4][465],u_xpb_out[5][465],u_xpb_out[6][465],u_xpb_out[7][465],u_xpb_out[8][465],u_xpb_out[9][465],u_xpb_out[10][465],u_xpb_out[11][465],u_xpb_out[12][465],u_xpb_out[13][465],u_xpb_out[14][465],u_xpb_out[15][465],u_xpb_out[16][465],u_xpb_out[17][465],u_xpb_out[18][465],u_xpb_out[19][465],u_xpb_out[20][465],u_xpb_out[21][465],u_xpb_out[22][465],u_xpb_out[23][465],u_xpb_out[24][465],u_xpb_out[25][465],u_xpb_out[26][465],u_xpb_out[27][465],u_xpb_out[28][465],u_xpb_out[29][465],u_xpb_out[30][465],u_xpb_out[31][465],u_xpb_out[32][465],u_xpb_out[33][465],u_xpb_out[34][465],u_xpb_out[35][465],u_xpb_out[36][465],u_xpb_out[37][465],u_xpb_out[38][465],u_xpb_out[39][465],u_xpb_out[40][465],u_xpb_out[41][465],u_xpb_out[42][465],u_xpb_out[43][465],u_xpb_out[44][465],u_xpb_out[45][465],u_xpb_out[46][465],u_xpb_out[47][465],u_xpb_out[48][465],u_xpb_out[49][465],u_xpb_out[50][465],u_xpb_out[51][465],u_xpb_out[52][465],u_xpb_out[53][465],u_xpb_out[54][465],u_xpb_out[55][465],u_xpb_out[56][465],u_xpb_out[57][465],u_xpb_out[58][465],u_xpb_out[59][465],u_xpb_out[60][465],u_xpb_out[61][465],u_xpb_out[62][465],u_xpb_out[63][465],u_xpb_out[64][465],u_xpb_out[65][465],u_xpb_out[66][465],u_xpb_out[67][465],u_xpb_out[68][465],u_xpb_out[69][465],u_xpb_out[70][465],u_xpb_out[71][465],u_xpb_out[72][465],u_xpb_out[73][465],u_xpb_out[74][465],u_xpb_out[75][465],u_xpb_out[76][465],u_xpb_out[77][465],u_xpb_out[78][465],u_xpb_out[79][465],u_xpb_out[80][465],u_xpb_out[81][465],u_xpb_out[82][465],u_xpb_out[83][465],u_xpb_out[84][465],u_xpb_out[85][465],u_xpb_out[86][465],u_xpb_out[87][465],u_xpb_out[88][465],u_xpb_out[89][465],u_xpb_out[90][465],u_xpb_out[91][465],u_xpb_out[92][465],u_xpb_out[93][465],u_xpb_out[94][465],u_xpb_out[95][465],u_xpb_out[96][465],u_xpb_out[97][465],u_xpb_out[98][465],u_xpb_out[99][465],u_xpb_out[100][465],u_xpb_out[101][465],u_xpb_out[102][465],u_xpb_out[103][465],u_xpb_out[104][465],u_xpb_out[105][465]};

assign col_out_466 = {u_xpb_out[0][466],u_xpb_out[1][466],u_xpb_out[2][466],u_xpb_out[3][466],u_xpb_out[4][466],u_xpb_out[5][466],u_xpb_out[6][466],u_xpb_out[7][466],u_xpb_out[8][466],u_xpb_out[9][466],u_xpb_out[10][466],u_xpb_out[11][466],u_xpb_out[12][466],u_xpb_out[13][466],u_xpb_out[14][466],u_xpb_out[15][466],u_xpb_out[16][466],u_xpb_out[17][466],u_xpb_out[18][466],u_xpb_out[19][466],u_xpb_out[20][466],u_xpb_out[21][466],u_xpb_out[22][466],u_xpb_out[23][466],u_xpb_out[24][466],u_xpb_out[25][466],u_xpb_out[26][466],u_xpb_out[27][466],u_xpb_out[28][466],u_xpb_out[29][466],u_xpb_out[30][466],u_xpb_out[31][466],u_xpb_out[32][466],u_xpb_out[33][466],u_xpb_out[34][466],u_xpb_out[35][466],u_xpb_out[36][466],u_xpb_out[37][466],u_xpb_out[38][466],u_xpb_out[39][466],u_xpb_out[40][466],u_xpb_out[41][466],u_xpb_out[42][466],u_xpb_out[43][466],u_xpb_out[44][466],u_xpb_out[45][466],u_xpb_out[46][466],u_xpb_out[47][466],u_xpb_out[48][466],u_xpb_out[49][466],u_xpb_out[50][466],u_xpb_out[51][466],u_xpb_out[52][466],u_xpb_out[53][466],u_xpb_out[54][466],u_xpb_out[55][466],u_xpb_out[56][466],u_xpb_out[57][466],u_xpb_out[58][466],u_xpb_out[59][466],u_xpb_out[60][466],u_xpb_out[61][466],u_xpb_out[62][466],u_xpb_out[63][466],u_xpb_out[64][466],u_xpb_out[65][466],u_xpb_out[66][466],u_xpb_out[67][466],u_xpb_out[68][466],u_xpb_out[69][466],u_xpb_out[70][466],u_xpb_out[71][466],u_xpb_out[72][466],u_xpb_out[73][466],u_xpb_out[74][466],u_xpb_out[75][466],u_xpb_out[76][466],u_xpb_out[77][466],u_xpb_out[78][466],u_xpb_out[79][466],u_xpb_out[80][466],u_xpb_out[81][466],u_xpb_out[82][466],u_xpb_out[83][466],u_xpb_out[84][466],u_xpb_out[85][466],u_xpb_out[86][466],u_xpb_out[87][466],u_xpb_out[88][466],u_xpb_out[89][466],u_xpb_out[90][466],u_xpb_out[91][466],u_xpb_out[92][466],u_xpb_out[93][466],u_xpb_out[94][466],u_xpb_out[95][466],u_xpb_out[96][466],u_xpb_out[97][466],u_xpb_out[98][466],u_xpb_out[99][466],u_xpb_out[100][466],u_xpb_out[101][466],u_xpb_out[102][466],u_xpb_out[103][466],u_xpb_out[104][466],u_xpb_out[105][466]};

assign col_out_467 = {u_xpb_out[0][467],u_xpb_out[1][467],u_xpb_out[2][467],u_xpb_out[3][467],u_xpb_out[4][467],u_xpb_out[5][467],u_xpb_out[6][467],u_xpb_out[7][467],u_xpb_out[8][467],u_xpb_out[9][467],u_xpb_out[10][467],u_xpb_out[11][467],u_xpb_out[12][467],u_xpb_out[13][467],u_xpb_out[14][467],u_xpb_out[15][467],u_xpb_out[16][467],u_xpb_out[17][467],u_xpb_out[18][467],u_xpb_out[19][467],u_xpb_out[20][467],u_xpb_out[21][467],u_xpb_out[22][467],u_xpb_out[23][467],u_xpb_out[24][467],u_xpb_out[25][467],u_xpb_out[26][467],u_xpb_out[27][467],u_xpb_out[28][467],u_xpb_out[29][467],u_xpb_out[30][467],u_xpb_out[31][467],u_xpb_out[32][467],u_xpb_out[33][467],u_xpb_out[34][467],u_xpb_out[35][467],u_xpb_out[36][467],u_xpb_out[37][467],u_xpb_out[38][467],u_xpb_out[39][467],u_xpb_out[40][467],u_xpb_out[41][467],u_xpb_out[42][467],u_xpb_out[43][467],u_xpb_out[44][467],u_xpb_out[45][467],u_xpb_out[46][467],u_xpb_out[47][467],u_xpb_out[48][467],u_xpb_out[49][467],u_xpb_out[50][467],u_xpb_out[51][467],u_xpb_out[52][467],u_xpb_out[53][467],u_xpb_out[54][467],u_xpb_out[55][467],u_xpb_out[56][467],u_xpb_out[57][467],u_xpb_out[58][467],u_xpb_out[59][467],u_xpb_out[60][467],u_xpb_out[61][467],u_xpb_out[62][467],u_xpb_out[63][467],u_xpb_out[64][467],u_xpb_out[65][467],u_xpb_out[66][467],u_xpb_out[67][467],u_xpb_out[68][467],u_xpb_out[69][467],u_xpb_out[70][467],u_xpb_out[71][467],u_xpb_out[72][467],u_xpb_out[73][467],u_xpb_out[74][467],u_xpb_out[75][467],u_xpb_out[76][467],u_xpb_out[77][467],u_xpb_out[78][467],u_xpb_out[79][467],u_xpb_out[80][467],u_xpb_out[81][467],u_xpb_out[82][467],u_xpb_out[83][467],u_xpb_out[84][467],u_xpb_out[85][467],u_xpb_out[86][467],u_xpb_out[87][467],u_xpb_out[88][467],u_xpb_out[89][467],u_xpb_out[90][467],u_xpb_out[91][467],u_xpb_out[92][467],u_xpb_out[93][467],u_xpb_out[94][467],u_xpb_out[95][467],u_xpb_out[96][467],u_xpb_out[97][467],u_xpb_out[98][467],u_xpb_out[99][467],u_xpb_out[100][467],u_xpb_out[101][467],u_xpb_out[102][467],u_xpb_out[103][467],u_xpb_out[104][467],u_xpb_out[105][467]};

assign col_out_468 = {u_xpb_out[0][468],u_xpb_out[1][468],u_xpb_out[2][468],u_xpb_out[3][468],u_xpb_out[4][468],u_xpb_out[5][468],u_xpb_out[6][468],u_xpb_out[7][468],u_xpb_out[8][468],u_xpb_out[9][468],u_xpb_out[10][468],u_xpb_out[11][468],u_xpb_out[12][468],u_xpb_out[13][468],u_xpb_out[14][468],u_xpb_out[15][468],u_xpb_out[16][468],u_xpb_out[17][468],u_xpb_out[18][468],u_xpb_out[19][468],u_xpb_out[20][468],u_xpb_out[21][468],u_xpb_out[22][468],u_xpb_out[23][468],u_xpb_out[24][468],u_xpb_out[25][468],u_xpb_out[26][468],u_xpb_out[27][468],u_xpb_out[28][468],u_xpb_out[29][468],u_xpb_out[30][468],u_xpb_out[31][468],u_xpb_out[32][468],u_xpb_out[33][468],u_xpb_out[34][468],u_xpb_out[35][468],u_xpb_out[36][468],u_xpb_out[37][468],u_xpb_out[38][468],u_xpb_out[39][468],u_xpb_out[40][468],u_xpb_out[41][468],u_xpb_out[42][468],u_xpb_out[43][468],u_xpb_out[44][468],u_xpb_out[45][468],u_xpb_out[46][468],u_xpb_out[47][468],u_xpb_out[48][468],u_xpb_out[49][468],u_xpb_out[50][468],u_xpb_out[51][468],u_xpb_out[52][468],u_xpb_out[53][468],u_xpb_out[54][468],u_xpb_out[55][468],u_xpb_out[56][468],u_xpb_out[57][468],u_xpb_out[58][468],u_xpb_out[59][468],u_xpb_out[60][468],u_xpb_out[61][468],u_xpb_out[62][468],u_xpb_out[63][468],u_xpb_out[64][468],u_xpb_out[65][468],u_xpb_out[66][468],u_xpb_out[67][468],u_xpb_out[68][468],u_xpb_out[69][468],u_xpb_out[70][468],u_xpb_out[71][468],u_xpb_out[72][468],u_xpb_out[73][468],u_xpb_out[74][468],u_xpb_out[75][468],u_xpb_out[76][468],u_xpb_out[77][468],u_xpb_out[78][468],u_xpb_out[79][468],u_xpb_out[80][468],u_xpb_out[81][468],u_xpb_out[82][468],u_xpb_out[83][468],u_xpb_out[84][468],u_xpb_out[85][468],u_xpb_out[86][468],u_xpb_out[87][468],u_xpb_out[88][468],u_xpb_out[89][468],u_xpb_out[90][468],u_xpb_out[91][468],u_xpb_out[92][468],u_xpb_out[93][468],u_xpb_out[94][468],u_xpb_out[95][468],u_xpb_out[96][468],u_xpb_out[97][468],u_xpb_out[98][468],u_xpb_out[99][468],u_xpb_out[100][468],u_xpb_out[101][468],u_xpb_out[102][468],u_xpb_out[103][468],u_xpb_out[104][468],u_xpb_out[105][468]};

assign col_out_469 = {u_xpb_out[0][469],u_xpb_out[1][469],u_xpb_out[2][469],u_xpb_out[3][469],u_xpb_out[4][469],u_xpb_out[5][469],u_xpb_out[6][469],u_xpb_out[7][469],u_xpb_out[8][469],u_xpb_out[9][469],u_xpb_out[10][469],u_xpb_out[11][469],u_xpb_out[12][469],u_xpb_out[13][469],u_xpb_out[14][469],u_xpb_out[15][469],u_xpb_out[16][469],u_xpb_out[17][469],u_xpb_out[18][469],u_xpb_out[19][469],u_xpb_out[20][469],u_xpb_out[21][469],u_xpb_out[22][469],u_xpb_out[23][469],u_xpb_out[24][469],u_xpb_out[25][469],u_xpb_out[26][469],u_xpb_out[27][469],u_xpb_out[28][469],u_xpb_out[29][469],u_xpb_out[30][469],u_xpb_out[31][469],u_xpb_out[32][469],u_xpb_out[33][469],u_xpb_out[34][469],u_xpb_out[35][469],u_xpb_out[36][469],u_xpb_out[37][469],u_xpb_out[38][469],u_xpb_out[39][469],u_xpb_out[40][469],u_xpb_out[41][469],u_xpb_out[42][469],u_xpb_out[43][469],u_xpb_out[44][469],u_xpb_out[45][469],u_xpb_out[46][469],u_xpb_out[47][469],u_xpb_out[48][469],u_xpb_out[49][469],u_xpb_out[50][469],u_xpb_out[51][469],u_xpb_out[52][469],u_xpb_out[53][469],u_xpb_out[54][469],u_xpb_out[55][469],u_xpb_out[56][469],u_xpb_out[57][469],u_xpb_out[58][469],u_xpb_out[59][469],u_xpb_out[60][469],u_xpb_out[61][469],u_xpb_out[62][469],u_xpb_out[63][469],u_xpb_out[64][469],u_xpb_out[65][469],u_xpb_out[66][469],u_xpb_out[67][469],u_xpb_out[68][469],u_xpb_out[69][469],u_xpb_out[70][469],u_xpb_out[71][469],u_xpb_out[72][469],u_xpb_out[73][469],u_xpb_out[74][469],u_xpb_out[75][469],u_xpb_out[76][469],u_xpb_out[77][469],u_xpb_out[78][469],u_xpb_out[79][469],u_xpb_out[80][469],u_xpb_out[81][469],u_xpb_out[82][469],u_xpb_out[83][469],u_xpb_out[84][469],u_xpb_out[85][469],u_xpb_out[86][469],u_xpb_out[87][469],u_xpb_out[88][469],u_xpb_out[89][469],u_xpb_out[90][469],u_xpb_out[91][469],u_xpb_out[92][469],u_xpb_out[93][469],u_xpb_out[94][469],u_xpb_out[95][469],u_xpb_out[96][469],u_xpb_out[97][469],u_xpb_out[98][469],u_xpb_out[99][469],u_xpb_out[100][469],u_xpb_out[101][469],u_xpb_out[102][469],u_xpb_out[103][469],u_xpb_out[104][469],u_xpb_out[105][469]};

assign col_out_470 = {u_xpb_out[0][470],u_xpb_out[1][470],u_xpb_out[2][470],u_xpb_out[3][470],u_xpb_out[4][470],u_xpb_out[5][470],u_xpb_out[6][470],u_xpb_out[7][470],u_xpb_out[8][470],u_xpb_out[9][470],u_xpb_out[10][470],u_xpb_out[11][470],u_xpb_out[12][470],u_xpb_out[13][470],u_xpb_out[14][470],u_xpb_out[15][470],u_xpb_out[16][470],u_xpb_out[17][470],u_xpb_out[18][470],u_xpb_out[19][470],u_xpb_out[20][470],u_xpb_out[21][470],u_xpb_out[22][470],u_xpb_out[23][470],u_xpb_out[24][470],u_xpb_out[25][470],u_xpb_out[26][470],u_xpb_out[27][470],u_xpb_out[28][470],u_xpb_out[29][470],u_xpb_out[30][470],u_xpb_out[31][470],u_xpb_out[32][470],u_xpb_out[33][470],u_xpb_out[34][470],u_xpb_out[35][470],u_xpb_out[36][470],u_xpb_out[37][470],u_xpb_out[38][470],u_xpb_out[39][470],u_xpb_out[40][470],u_xpb_out[41][470],u_xpb_out[42][470],u_xpb_out[43][470],u_xpb_out[44][470],u_xpb_out[45][470],u_xpb_out[46][470],u_xpb_out[47][470],u_xpb_out[48][470],u_xpb_out[49][470],u_xpb_out[50][470],u_xpb_out[51][470],u_xpb_out[52][470],u_xpb_out[53][470],u_xpb_out[54][470],u_xpb_out[55][470],u_xpb_out[56][470],u_xpb_out[57][470],u_xpb_out[58][470],u_xpb_out[59][470],u_xpb_out[60][470],u_xpb_out[61][470],u_xpb_out[62][470],u_xpb_out[63][470],u_xpb_out[64][470],u_xpb_out[65][470],u_xpb_out[66][470],u_xpb_out[67][470],u_xpb_out[68][470],u_xpb_out[69][470],u_xpb_out[70][470],u_xpb_out[71][470],u_xpb_out[72][470],u_xpb_out[73][470],u_xpb_out[74][470],u_xpb_out[75][470],u_xpb_out[76][470],u_xpb_out[77][470],u_xpb_out[78][470],u_xpb_out[79][470],u_xpb_out[80][470],u_xpb_out[81][470],u_xpb_out[82][470],u_xpb_out[83][470],u_xpb_out[84][470],u_xpb_out[85][470],u_xpb_out[86][470],u_xpb_out[87][470],u_xpb_out[88][470],u_xpb_out[89][470],u_xpb_out[90][470],u_xpb_out[91][470],u_xpb_out[92][470],u_xpb_out[93][470],u_xpb_out[94][470],u_xpb_out[95][470],u_xpb_out[96][470],u_xpb_out[97][470],u_xpb_out[98][470],u_xpb_out[99][470],u_xpb_out[100][470],u_xpb_out[101][470],u_xpb_out[102][470],u_xpb_out[103][470],u_xpb_out[104][470],u_xpb_out[105][470]};

assign col_out_471 = {u_xpb_out[0][471],u_xpb_out[1][471],u_xpb_out[2][471],u_xpb_out[3][471],u_xpb_out[4][471],u_xpb_out[5][471],u_xpb_out[6][471],u_xpb_out[7][471],u_xpb_out[8][471],u_xpb_out[9][471],u_xpb_out[10][471],u_xpb_out[11][471],u_xpb_out[12][471],u_xpb_out[13][471],u_xpb_out[14][471],u_xpb_out[15][471],u_xpb_out[16][471],u_xpb_out[17][471],u_xpb_out[18][471],u_xpb_out[19][471],u_xpb_out[20][471],u_xpb_out[21][471],u_xpb_out[22][471],u_xpb_out[23][471],u_xpb_out[24][471],u_xpb_out[25][471],u_xpb_out[26][471],u_xpb_out[27][471],u_xpb_out[28][471],u_xpb_out[29][471],u_xpb_out[30][471],u_xpb_out[31][471],u_xpb_out[32][471],u_xpb_out[33][471],u_xpb_out[34][471],u_xpb_out[35][471],u_xpb_out[36][471],u_xpb_out[37][471],u_xpb_out[38][471],u_xpb_out[39][471],u_xpb_out[40][471],u_xpb_out[41][471],u_xpb_out[42][471],u_xpb_out[43][471],u_xpb_out[44][471],u_xpb_out[45][471],u_xpb_out[46][471],u_xpb_out[47][471],u_xpb_out[48][471],u_xpb_out[49][471],u_xpb_out[50][471],u_xpb_out[51][471],u_xpb_out[52][471],u_xpb_out[53][471],u_xpb_out[54][471],u_xpb_out[55][471],u_xpb_out[56][471],u_xpb_out[57][471],u_xpb_out[58][471],u_xpb_out[59][471],u_xpb_out[60][471],u_xpb_out[61][471],u_xpb_out[62][471],u_xpb_out[63][471],u_xpb_out[64][471],u_xpb_out[65][471],u_xpb_out[66][471],u_xpb_out[67][471],u_xpb_out[68][471],u_xpb_out[69][471],u_xpb_out[70][471],u_xpb_out[71][471],u_xpb_out[72][471],u_xpb_out[73][471],u_xpb_out[74][471],u_xpb_out[75][471],u_xpb_out[76][471],u_xpb_out[77][471],u_xpb_out[78][471],u_xpb_out[79][471],u_xpb_out[80][471],u_xpb_out[81][471],u_xpb_out[82][471],u_xpb_out[83][471],u_xpb_out[84][471],u_xpb_out[85][471],u_xpb_out[86][471],u_xpb_out[87][471],u_xpb_out[88][471],u_xpb_out[89][471],u_xpb_out[90][471],u_xpb_out[91][471],u_xpb_out[92][471],u_xpb_out[93][471],u_xpb_out[94][471],u_xpb_out[95][471],u_xpb_out[96][471],u_xpb_out[97][471],u_xpb_out[98][471],u_xpb_out[99][471],u_xpb_out[100][471],u_xpb_out[101][471],u_xpb_out[102][471],u_xpb_out[103][471],u_xpb_out[104][471],u_xpb_out[105][471]};

assign col_out_472 = {u_xpb_out[0][472],u_xpb_out[1][472],u_xpb_out[2][472],u_xpb_out[3][472],u_xpb_out[4][472],u_xpb_out[5][472],u_xpb_out[6][472],u_xpb_out[7][472],u_xpb_out[8][472],u_xpb_out[9][472],u_xpb_out[10][472],u_xpb_out[11][472],u_xpb_out[12][472],u_xpb_out[13][472],u_xpb_out[14][472],u_xpb_out[15][472],u_xpb_out[16][472],u_xpb_out[17][472],u_xpb_out[18][472],u_xpb_out[19][472],u_xpb_out[20][472],u_xpb_out[21][472],u_xpb_out[22][472],u_xpb_out[23][472],u_xpb_out[24][472],u_xpb_out[25][472],u_xpb_out[26][472],u_xpb_out[27][472],u_xpb_out[28][472],u_xpb_out[29][472],u_xpb_out[30][472],u_xpb_out[31][472],u_xpb_out[32][472],u_xpb_out[33][472],u_xpb_out[34][472],u_xpb_out[35][472],u_xpb_out[36][472],u_xpb_out[37][472],u_xpb_out[38][472],u_xpb_out[39][472],u_xpb_out[40][472],u_xpb_out[41][472],u_xpb_out[42][472],u_xpb_out[43][472],u_xpb_out[44][472],u_xpb_out[45][472],u_xpb_out[46][472],u_xpb_out[47][472],u_xpb_out[48][472],u_xpb_out[49][472],u_xpb_out[50][472],u_xpb_out[51][472],u_xpb_out[52][472],u_xpb_out[53][472],u_xpb_out[54][472],u_xpb_out[55][472],u_xpb_out[56][472],u_xpb_out[57][472],u_xpb_out[58][472],u_xpb_out[59][472],u_xpb_out[60][472],u_xpb_out[61][472],u_xpb_out[62][472],u_xpb_out[63][472],u_xpb_out[64][472],u_xpb_out[65][472],u_xpb_out[66][472],u_xpb_out[67][472],u_xpb_out[68][472],u_xpb_out[69][472],u_xpb_out[70][472],u_xpb_out[71][472],u_xpb_out[72][472],u_xpb_out[73][472],u_xpb_out[74][472],u_xpb_out[75][472],u_xpb_out[76][472],u_xpb_out[77][472],u_xpb_out[78][472],u_xpb_out[79][472],u_xpb_out[80][472],u_xpb_out[81][472],u_xpb_out[82][472],u_xpb_out[83][472],u_xpb_out[84][472],u_xpb_out[85][472],u_xpb_out[86][472],u_xpb_out[87][472],u_xpb_out[88][472],u_xpb_out[89][472],u_xpb_out[90][472],u_xpb_out[91][472],u_xpb_out[92][472],u_xpb_out[93][472],u_xpb_out[94][472],u_xpb_out[95][472],u_xpb_out[96][472],u_xpb_out[97][472],u_xpb_out[98][472],u_xpb_out[99][472],u_xpb_out[100][472],u_xpb_out[101][472],u_xpb_out[102][472],u_xpb_out[103][472],u_xpb_out[104][472],u_xpb_out[105][472]};

assign col_out_473 = {u_xpb_out[0][473],u_xpb_out[1][473],u_xpb_out[2][473],u_xpb_out[3][473],u_xpb_out[4][473],u_xpb_out[5][473],u_xpb_out[6][473],u_xpb_out[7][473],u_xpb_out[8][473],u_xpb_out[9][473],u_xpb_out[10][473],u_xpb_out[11][473],u_xpb_out[12][473],u_xpb_out[13][473],u_xpb_out[14][473],u_xpb_out[15][473],u_xpb_out[16][473],u_xpb_out[17][473],u_xpb_out[18][473],u_xpb_out[19][473],u_xpb_out[20][473],u_xpb_out[21][473],u_xpb_out[22][473],u_xpb_out[23][473],u_xpb_out[24][473],u_xpb_out[25][473],u_xpb_out[26][473],u_xpb_out[27][473],u_xpb_out[28][473],u_xpb_out[29][473],u_xpb_out[30][473],u_xpb_out[31][473],u_xpb_out[32][473],u_xpb_out[33][473],u_xpb_out[34][473],u_xpb_out[35][473],u_xpb_out[36][473],u_xpb_out[37][473],u_xpb_out[38][473],u_xpb_out[39][473],u_xpb_out[40][473],u_xpb_out[41][473],u_xpb_out[42][473],u_xpb_out[43][473],u_xpb_out[44][473],u_xpb_out[45][473],u_xpb_out[46][473],u_xpb_out[47][473],u_xpb_out[48][473],u_xpb_out[49][473],u_xpb_out[50][473],u_xpb_out[51][473],u_xpb_out[52][473],u_xpb_out[53][473],u_xpb_out[54][473],u_xpb_out[55][473],u_xpb_out[56][473],u_xpb_out[57][473],u_xpb_out[58][473],u_xpb_out[59][473],u_xpb_out[60][473],u_xpb_out[61][473],u_xpb_out[62][473],u_xpb_out[63][473],u_xpb_out[64][473],u_xpb_out[65][473],u_xpb_out[66][473],u_xpb_out[67][473],u_xpb_out[68][473],u_xpb_out[69][473],u_xpb_out[70][473],u_xpb_out[71][473],u_xpb_out[72][473],u_xpb_out[73][473],u_xpb_out[74][473],u_xpb_out[75][473],u_xpb_out[76][473],u_xpb_out[77][473],u_xpb_out[78][473],u_xpb_out[79][473],u_xpb_out[80][473],u_xpb_out[81][473],u_xpb_out[82][473],u_xpb_out[83][473],u_xpb_out[84][473],u_xpb_out[85][473],u_xpb_out[86][473],u_xpb_out[87][473],u_xpb_out[88][473],u_xpb_out[89][473],u_xpb_out[90][473],u_xpb_out[91][473],u_xpb_out[92][473],u_xpb_out[93][473],u_xpb_out[94][473],u_xpb_out[95][473],u_xpb_out[96][473],u_xpb_out[97][473],u_xpb_out[98][473],u_xpb_out[99][473],u_xpb_out[100][473],u_xpb_out[101][473],u_xpb_out[102][473],u_xpb_out[103][473],u_xpb_out[104][473],u_xpb_out[105][473]};

assign col_out_474 = {u_xpb_out[0][474],u_xpb_out[1][474],u_xpb_out[2][474],u_xpb_out[3][474],u_xpb_out[4][474],u_xpb_out[5][474],u_xpb_out[6][474],u_xpb_out[7][474],u_xpb_out[8][474],u_xpb_out[9][474],u_xpb_out[10][474],u_xpb_out[11][474],u_xpb_out[12][474],u_xpb_out[13][474],u_xpb_out[14][474],u_xpb_out[15][474],u_xpb_out[16][474],u_xpb_out[17][474],u_xpb_out[18][474],u_xpb_out[19][474],u_xpb_out[20][474],u_xpb_out[21][474],u_xpb_out[22][474],u_xpb_out[23][474],u_xpb_out[24][474],u_xpb_out[25][474],u_xpb_out[26][474],u_xpb_out[27][474],u_xpb_out[28][474],u_xpb_out[29][474],u_xpb_out[30][474],u_xpb_out[31][474],u_xpb_out[32][474],u_xpb_out[33][474],u_xpb_out[34][474],u_xpb_out[35][474],u_xpb_out[36][474],u_xpb_out[37][474],u_xpb_out[38][474],u_xpb_out[39][474],u_xpb_out[40][474],u_xpb_out[41][474],u_xpb_out[42][474],u_xpb_out[43][474],u_xpb_out[44][474],u_xpb_out[45][474],u_xpb_out[46][474],u_xpb_out[47][474],u_xpb_out[48][474],u_xpb_out[49][474],u_xpb_out[50][474],u_xpb_out[51][474],u_xpb_out[52][474],u_xpb_out[53][474],u_xpb_out[54][474],u_xpb_out[55][474],u_xpb_out[56][474],u_xpb_out[57][474],u_xpb_out[58][474],u_xpb_out[59][474],u_xpb_out[60][474],u_xpb_out[61][474],u_xpb_out[62][474],u_xpb_out[63][474],u_xpb_out[64][474],u_xpb_out[65][474],u_xpb_out[66][474],u_xpb_out[67][474],u_xpb_out[68][474],u_xpb_out[69][474],u_xpb_out[70][474],u_xpb_out[71][474],u_xpb_out[72][474],u_xpb_out[73][474],u_xpb_out[74][474],u_xpb_out[75][474],u_xpb_out[76][474],u_xpb_out[77][474],u_xpb_out[78][474],u_xpb_out[79][474],u_xpb_out[80][474],u_xpb_out[81][474],u_xpb_out[82][474],u_xpb_out[83][474],u_xpb_out[84][474],u_xpb_out[85][474],u_xpb_out[86][474],u_xpb_out[87][474],u_xpb_out[88][474],u_xpb_out[89][474],u_xpb_out[90][474],u_xpb_out[91][474],u_xpb_out[92][474],u_xpb_out[93][474],u_xpb_out[94][474],u_xpb_out[95][474],u_xpb_out[96][474],u_xpb_out[97][474],u_xpb_out[98][474],u_xpb_out[99][474],u_xpb_out[100][474],u_xpb_out[101][474],u_xpb_out[102][474],u_xpb_out[103][474],u_xpb_out[104][474],u_xpb_out[105][474]};

assign col_out_475 = {u_xpb_out[0][475],u_xpb_out[1][475],u_xpb_out[2][475],u_xpb_out[3][475],u_xpb_out[4][475],u_xpb_out[5][475],u_xpb_out[6][475],u_xpb_out[7][475],u_xpb_out[8][475],u_xpb_out[9][475],u_xpb_out[10][475],u_xpb_out[11][475],u_xpb_out[12][475],u_xpb_out[13][475],u_xpb_out[14][475],u_xpb_out[15][475],u_xpb_out[16][475],u_xpb_out[17][475],u_xpb_out[18][475],u_xpb_out[19][475],u_xpb_out[20][475],u_xpb_out[21][475],u_xpb_out[22][475],u_xpb_out[23][475],u_xpb_out[24][475],u_xpb_out[25][475],u_xpb_out[26][475],u_xpb_out[27][475],u_xpb_out[28][475],u_xpb_out[29][475],u_xpb_out[30][475],u_xpb_out[31][475],u_xpb_out[32][475],u_xpb_out[33][475],u_xpb_out[34][475],u_xpb_out[35][475],u_xpb_out[36][475],u_xpb_out[37][475],u_xpb_out[38][475],u_xpb_out[39][475],u_xpb_out[40][475],u_xpb_out[41][475],u_xpb_out[42][475],u_xpb_out[43][475],u_xpb_out[44][475],u_xpb_out[45][475],u_xpb_out[46][475],u_xpb_out[47][475],u_xpb_out[48][475],u_xpb_out[49][475],u_xpb_out[50][475],u_xpb_out[51][475],u_xpb_out[52][475],u_xpb_out[53][475],u_xpb_out[54][475],u_xpb_out[55][475],u_xpb_out[56][475],u_xpb_out[57][475],u_xpb_out[58][475],u_xpb_out[59][475],u_xpb_out[60][475],u_xpb_out[61][475],u_xpb_out[62][475],u_xpb_out[63][475],u_xpb_out[64][475],u_xpb_out[65][475],u_xpb_out[66][475],u_xpb_out[67][475],u_xpb_out[68][475],u_xpb_out[69][475],u_xpb_out[70][475],u_xpb_out[71][475],u_xpb_out[72][475],u_xpb_out[73][475],u_xpb_out[74][475],u_xpb_out[75][475],u_xpb_out[76][475],u_xpb_out[77][475],u_xpb_out[78][475],u_xpb_out[79][475],u_xpb_out[80][475],u_xpb_out[81][475],u_xpb_out[82][475],u_xpb_out[83][475],u_xpb_out[84][475],u_xpb_out[85][475],u_xpb_out[86][475],u_xpb_out[87][475],u_xpb_out[88][475],u_xpb_out[89][475],u_xpb_out[90][475],u_xpb_out[91][475],u_xpb_out[92][475],u_xpb_out[93][475],u_xpb_out[94][475],u_xpb_out[95][475],u_xpb_out[96][475],u_xpb_out[97][475],u_xpb_out[98][475],u_xpb_out[99][475],u_xpb_out[100][475],u_xpb_out[101][475],u_xpb_out[102][475],u_xpb_out[103][475],u_xpb_out[104][475],u_xpb_out[105][475]};

assign col_out_476 = {u_xpb_out[0][476],u_xpb_out[1][476],u_xpb_out[2][476],u_xpb_out[3][476],u_xpb_out[4][476],u_xpb_out[5][476],u_xpb_out[6][476],u_xpb_out[7][476],u_xpb_out[8][476],u_xpb_out[9][476],u_xpb_out[10][476],u_xpb_out[11][476],u_xpb_out[12][476],u_xpb_out[13][476],u_xpb_out[14][476],u_xpb_out[15][476],u_xpb_out[16][476],u_xpb_out[17][476],u_xpb_out[18][476],u_xpb_out[19][476],u_xpb_out[20][476],u_xpb_out[21][476],u_xpb_out[22][476],u_xpb_out[23][476],u_xpb_out[24][476],u_xpb_out[25][476],u_xpb_out[26][476],u_xpb_out[27][476],u_xpb_out[28][476],u_xpb_out[29][476],u_xpb_out[30][476],u_xpb_out[31][476],u_xpb_out[32][476],u_xpb_out[33][476],u_xpb_out[34][476],u_xpb_out[35][476],u_xpb_out[36][476],u_xpb_out[37][476],u_xpb_out[38][476],u_xpb_out[39][476],u_xpb_out[40][476],u_xpb_out[41][476],u_xpb_out[42][476],u_xpb_out[43][476],u_xpb_out[44][476],u_xpb_out[45][476],u_xpb_out[46][476],u_xpb_out[47][476],u_xpb_out[48][476],u_xpb_out[49][476],u_xpb_out[50][476],u_xpb_out[51][476],u_xpb_out[52][476],u_xpb_out[53][476],u_xpb_out[54][476],u_xpb_out[55][476],u_xpb_out[56][476],u_xpb_out[57][476],u_xpb_out[58][476],u_xpb_out[59][476],u_xpb_out[60][476],u_xpb_out[61][476],u_xpb_out[62][476],u_xpb_out[63][476],u_xpb_out[64][476],u_xpb_out[65][476],u_xpb_out[66][476],u_xpb_out[67][476],u_xpb_out[68][476],u_xpb_out[69][476],u_xpb_out[70][476],u_xpb_out[71][476],u_xpb_out[72][476],u_xpb_out[73][476],u_xpb_out[74][476],u_xpb_out[75][476],u_xpb_out[76][476],u_xpb_out[77][476],u_xpb_out[78][476],u_xpb_out[79][476],u_xpb_out[80][476],u_xpb_out[81][476],u_xpb_out[82][476],u_xpb_out[83][476],u_xpb_out[84][476],u_xpb_out[85][476],u_xpb_out[86][476],u_xpb_out[87][476],u_xpb_out[88][476],u_xpb_out[89][476],u_xpb_out[90][476],u_xpb_out[91][476],u_xpb_out[92][476],u_xpb_out[93][476],u_xpb_out[94][476],u_xpb_out[95][476],u_xpb_out[96][476],u_xpb_out[97][476],u_xpb_out[98][476],u_xpb_out[99][476],u_xpb_out[100][476],u_xpb_out[101][476],u_xpb_out[102][476],u_xpb_out[103][476],u_xpb_out[104][476],u_xpb_out[105][476]};

assign col_out_477 = {u_xpb_out[0][477],u_xpb_out[1][477],u_xpb_out[2][477],u_xpb_out[3][477],u_xpb_out[4][477],u_xpb_out[5][477],u_xpb_out[6][477],u_xpb_out[7][477],u_xpb_out[8][477],u_xpb_out[9][477],u_xpb_out[10][477],u_xpb_out[11][477],u_xpb_out[12][477],u_xpb_out[13][477],u_xpb_out[14][477],u_xpb_out[15][477],u_xpb_out[16][477],u_xpb_out[17][477],u_xpb_out[18][477],u_xpb_out[19][477],u_xpb_out[20][477],u_xpb_out[21][477],u_xpb_out[22][477],u_xpb_out[23][477],u_xpb_out[24][477],u_xpb_out[25][477],u_xpb_out[26][477],u_xpb_out[27][477],u_xpb_out[28][477],u_xpb_out[29][477],u_xpb_out[30][477],u_xpb_out[31][477],u_xpb_out[32][477],u_xpb_out[33][477],u_xpb_out[34][477],u_xpb_out[35][477],u_xpb_out[36][477],u_xpb_out[37][477],u_xpb_out[38][477],u_xpb_out[39][477],u_xpb_out[40][477],u_xpb_out[41][477],u_xpb_out[42][477],u_xpb_out[43][477],u_xpb_out[44][477],u_xpb_out[45][477],u_xpb_out[46][477],u_xpb_out[47][477],u_xpb_out[48][477],u_xpb_out[49][477],u_xpb_out[50][477],u_xpb_out[51][477],u_xpb_out[52][477],u_xpb_out[53][477],u_xpb_out[54][477],u_xpb_out[55][477],u_xpb_out[56][477],u_xpb_out[57][477],u_xpb_out[58][477],u_xpb_out[59][477],u_xpb_out[60][477],u_xpb_out[61][477],u_xpb_out[62][477],u_xpb_out[63][477],u_xpb_out[64][477],u_xpb_out[65][477],u_xpb_out[66][477],u_xpb_out[67][477],u_xpb_out[68][477],u_xpb_out[69][477],u_xpb_out[70][477],u_xpb_out[71][477],u_xpb_out[72][477],u_xpb_out[73][477],u_xpb_out[74][477],u_xpb_out[75][477],u_xpb_out[76][477],u_xpb_out[77][477],u_xpb_out[78][477],u_xpb_out[79][477],u_xpb_out[80][477],u_xpb_out[81][477],u_xpb_out[82][477],u_xpb_out[83][477],u_xpb_out[84][477],u_xpb_out[85][477],u_xpb_out[86][477],u_xpb_out[87][477],u_xpb_out[88][477],u_xpb_out[89][477],u_xpb_out[90][477],u_xpb_out[91][477],u_xpb_out[92][477],u_xpb_out[93][477],u_xpb_out[94][477],u_xpb_out[95][477],u_xpb_out[96][477],u_xpb_out[97][477],u_xpb_out[98][477],u_xpb_out[99][477],u_xpb_out[100][477],u_xpb_out[101][477],u_xpb_out[102][477],u_xpb_out[103][477],u_xpb_out[104][477],u_xpb_out[105][477]};

assign col_out_478 = {u_xpb_out[0][478],u_xpb_out[1][478],u_xpb_out[2][478],u_xpb_out[3][478],u_xpb_out[4][478],u_xpb_out[5][478],u_xpb_out[6][478],u_xpb_out[7][478],u_xpb_out[8][478],u_xpb_out[9][478],u_xpb_out[10][478],u_xpb_out[11][478],u_xpb_out[12][478],u_xpb_out[13][478],u_xpb_out[14][478],u_xpb_out[15][478],u_xpb_out[16][478],u_xpb_out[17][478],u_xpb_out[18][478],u_xpb_out[19][478],u_xpb_out[20][478],u_xpb_out[21][478],u_xpb_out[22][478],u_xpb_out[23][478],u_xpb_out[24][478],u_xpb_out[25][478],u_xpb_out[26][478],u_xpb_out[27][478],u_xpb_out[28][478],u_xpb_out[29][478],u_xpb_out[30][478],u_xpb_out[31][478],u_xpb_out[32][478],u_xpb_out[33][478],u_xpb_out[34][478],u_xpb_out[35][478],u_xpb_out[36][478],u_xpb_out[37][478],u_xpb_out[38][478],u_xpb_out[39][478],u_xpb_out[40][478],u_xpb_out[41][478],u_xpb_out[42][478],u_xpb_out[43][478],u_xpb_out[44][478],u_xpb_out[45][478],u_xpb_out[46][478],u_xpb_out[47][478],u_xpb_out[48][478],u_xpb_out[49][478],u_xpb_out[50][478],u_xpb_out[51][478],u_xpb_out[52][478],u_xpb_out[53][478],u_xpb_out[54][478],u_xpb_out[55][478],u_xpb_out[56][478],u_xpb_out[57][478],u_xpb_out[58][478],u_xpb_out[59][478],u_xpb_out[60][478],u_xpb_out[61][478],u_xpb_out[62][478],u_xpb_out[63][478],u_xpb_out[64][478],u_xpb_out[65][478],u_xpb_out[66][478],u_xpb_out[67][478],u_xpb_out[68][478],u_xpb_out[69][478],u_xpb_out[70][478],u_xpb_out[71][478],u_xpb_out[72][478],u_xpb_out[73][478],u_xpb_out[74][478],u_xpb_out[75][478],u_xpb_out[76][478],u_xpb_out[77][478],u_xpb_out[78][478],u_xpb_out[79][478],u_xpb_out[80][478],u_xpb_out[81][478],u_xpb_out[82][478],u_xpb_out[83][478],u_xpb_out[84][478],u_xpb_out[85][478],u_xpb_out[86][478],u_xpb_out[87][478],u_xpb_out[88][478],u_xpb_out[89][478],u_xpb_out[90][478],u_xpb_out[91][478],u_xpb_out[92][478],u_xpb_out[93][478],u_xpb_out[94][478],u_xpb_out[95][478],u_xpb_out[96][478],u_xpb_out[97][478],u_xpb_out[98][478],u_xpb_out[99][478],u_xpb_out[100][478],u_xpb_out[101][478],u_xpb_out[102][478],u_xpb_out[103][478],u_xpb_out[104][478],u_xpb_out[105][478]};

assign col_out_479 = {u_xpb_out[0][479],u_xpb_out[1][479],u_xpb_out[2][479],u_xpb_out[3][479],u_xpb_out[4][479],u_xpb_out[5][479],u_xpb_out[6][479],u_xpb_out[7][479],u_xpb_out[8][479],u_xpb_out[9][479],u_xpb_out[10][479],u_xpb_out[11][479],u_xpb_out[12][479],u_xpb_out[13][479],u_xpb_out[14][479],u_xpb_out[15][479],u_xpb_out[16][479],u_xpb_out[17][479],u_xpb_out[18][479],u_xpb_out[19][479],u_xpb_out[20][479],u_xpb_out[21][479],u_xpb_out[22][479],u_xpb_out[23][479],u_xpb_out[24][479],u_xpb_out[25][479],u_xpb_out[26][479],u_xpb_out[27][479],u_xpb_out[28][479],u_xpb_out[29][479],u_xpb_out[30][479],u_xpb_out[31][479],u_xpb_out[32][479],u_xpb_out[33][479],u_xpb_out[34][479],u_xpb_out[35][479],u_xpb_out[36][479],u_xpb_out[37][479],u_xpb_out[38][479],u_xpb_out[39][479],u_xpb_out[40][479],u_xpb_out[41][479],u_xpb_out[42][479],u_xpb_out[43][479],u_xpb_out[44][479],u_xpb_out[45][479],u_xpb_out[46][479],u_xpb_out[47][479],u_xpb_out[48][479],u_xpb_out[49][479],u_xpb_out[50][479],u_xpb_out[51][479],u_xpb_out[52][479],u_xpb_out[53][479],u_xpb_out[54][479],u_xpb_out[55][479],u_xpb_out[56][479],u_xpb_out[57][479],u_xpb_out[58][479],u_xpb_out[59][479],u_xpb_out[60][479],u_xpb_out[61][479],u_xpb_out[62][479],u_xpb_out[63][479],u_xpb_out[64][479],u_xpb_out[65][479],u_xpb_out[66][479],u_xpb_out[67][479],u_xpb_out[68][479],u_xpb_out[69][479],u_xpb_out[70][479],u_xpb_out[71][479],u_xpb_out[72][479],u_xpb_out[73][479],u_xpb_out[74][479],u_xpb_out[75][479],u_xpb_out[76][479],u_xpb_out[77][479],u_xpb_out[78][479],u_xpb_out[79][479],u_xpb_out[80][479],u_xpb_out[81][479],u_xpb_out[82][479],u_xpb_out[83][479],u_xpb_out[84][479],u_xpb_out[85][479],u_xpb_out[86][479],u_xpb_out[87][479],u_xpb_out[88][479],u_xpb_out[89][479],u_xpb_out[90][479],u_xpb_out[91][479],u_xpb_out[92][479],u_xpb_out[93][479],u_xpb_out[94][479],u_xpb_out[95][479],u_xpb_out[96][479],u_xpb_out[97][479],u_xpb_out[98][479],u_xpb_out[99][479],u_xpb_out[100][479],u_xpb_out[101][479],u_xpb_out[102][479],u_xpb_out[103][479],u_xpb_out[104][479],u_xpb_out[105][479]};

assign col_out_480 = {u_xpb_out[0][480],u_xpb_out[1][480],u_xpb_out[2][480],u_xpb_out[3][480],u_xpb_out[4][480],u_xpb_out[5][480],u_xpb_out[6][480],u_xpb_out[7][480],u_xpb_out[8][480],u_xpb_out[9][480],u_xpb_out[10][480],u_xpb_out[11][480],u_xpb_out[12][480],u_xpb_out[13][480],u_xpb_out[14][480],u_xpb_out[15][480],u_xpb_out[16][480],u_xpb_out[17][480],u_xpb_out[18][480],u_xpb_out[19][480],u_xpb_out[20][480],u_xpb_out[21][480],u_xpb_out[22][480],u_xpb_out[23][480],u_xpb_out[24][480],u_xpb_out[25][480],u_xpb_out[26][480],u_xpb_out[27][480],u_xpb_out[28][480],u_xpb_out[29][480],u_xpb_out[30][480],u_xpb_out[31][480],u_xpb_out[32][480],u_xpb_out[33][480],u_xpb_out[34][480],u_xpb_out[35][480],u_xpb_out[36][480],u_xpb_out[37][480],u_xpb_out[38][480],u_xpb_out[39][480],u_xpb_out[40][480],u_xpb_out[41][480],u_xpb_out[42][480],u_xpb_out[43][480],u_xpb_out[44][480],u_xpb_out[45][480],u_xpb_out[46][480],u_xpb_out[47][480],u_xpb_out[48][480],u_xpb_out[49][480],u_xpb_out[50][480],u_xpb_out[51][480],u_xpb_out[52][480],u_xpb_out[53][480],u_xpb_out[54][480],u_xpb_out[55][480],u_xpb_out[56][480],u_xpb_out[57][480],u_xpb_out[58][480],u_xpb_out[59][480],u_xpb_out[60][480],u_xpb_out[61][480],u_xpb_out[62][480],u_xpb_out[63][480],u_xpb_out[64][480],u_xpb_out[65][480],u_xpb_out[66][480],u_xpb_out[67][480],u_xpb_out[68][480],u_xpb_out[69][480],u_xpb_out[70][480],u_xpb_out[71][480],u_xpb_out[72][480],u_xpb_out[73][480],u_xpb_out[74][480],u_xpb_out[75][480],u_xpb_out[76][480],u_xpb_out[77][480],u_xpb_out[78][480],u_xpb_out[79][480],u_xpb_out[80][480],u_xpb_out[81][480],u_xpb_out[82][480],u_xpb_out[83][480],u_xpb_out[84][480],u_xpb_out[85][480],u_xpb_out[86][480],u_xpb_out[87][480],u_xpb_out[88][480],u_xpb_out[89][480],u_xpb_out[90][480],u_xpb_out[91][480],u_xpb_out[92][480],u_xpb_out[93][480],u_xpb_out[94][480],u_xpb_out[95][480],u_xpb_out[96][480],u_xpb_out[97][480],u_xpb_out[98][480],u_xpb_out[99][480],u_xpb_out[100][480],u_xpb_out[101][480],u_xpb_out[102][480],u_xpb_out[103][480],u_xpb_out[104][480],u_xpb_out[105][480]};

assign col_out_481 = {u_xpb_out[0][481],u_xpb_out[1][481],u_xpb_out[2][481],u_xpb_out[3][481],u_xpb_out[4][481],u_xpb_out[5][481],u_xpb_out[6][481],u_xpb_out[7][481],u_xpb_out[8][481],u_xpb_out[9][481],u_xpb_out[10][481],u_xpb_out[11][481],u_xpb_out[12][481],u_xpb_out[13][481],u_xpb_out[14][481],u_xpb_out[15][481],u_xpb_out[16][481],u_xpb_out[17][481],u_xpb_out[18][481],u_xpb_out[19][481],u_xpb_out[20][481],u_xpb_out[21][481],u_xpb_out[22][481],u_xpb_out[23][481],u_xpb_out[24][481],u_xpb_out[25][481],u_xpb_out[26][481],u_xpb_out[27][481],u_xpb_out[28][481],u_xpb_out[29][481],u_xpb_out[30][481],u_xpb_out[31][481],u_xpb_out[32][481],u_xpb_out[33][481],u_xpb_out[34][481],u_xpb_out[35][481],u_xpb_out[36][481],u_xpb_out[37][481],u_xpb_out[38][481],u_xpb_out[39][481],u_xpb_out[40][481],u_xpb_out[41][481],u_xpb_out[42][481],u_xpb_out[43][481],u_xpb_out[44][481],u_xpb_out[45][481],u_xpb_out[46][481],u_xpb_out[47][481],u_xpb_out[48][481],u_xpb_out[49][481],u_xpb_out[50][481],u_xpb_out[51][481],u_xpb_out[52][481],u_xpb_out[53][481],u_xpb_out[54][481],u_xpb_out[55][481],u_xpb_out[56][481],u_xpb_out[57][481],u_xpb_out[58][481],u_xpb_out[59][481],u_xpb_out[60][481],u_xpb_out[61][481],u_xpb_out[62][481],u_xpb_out[63][481],u_xpb_out[64][481],u_xpb_out[65][481],u_xpb_out[66][481],u_xpb_out[67][481],u_xpb_out[68][481],u_xpb_out[69][481],u_xpb_out[70][481],u_xpb_out[71][481],u_xpb_out[72][481],u_xpb_out[73][481],u_xpb_out[74][481],u_xpb_out[75][481],u_xpb_out[76][481],u_xpb_out[77][481],u_xpb_out[78][481],u_xpb_out[79][481],u_xpb_out[80][481],u_xpb_out[81][481],u_xpb_out[82][481],u_xpb_out[83][481],u_xpb_out[84][481],u_xpb_out[85][481],u_xpb_out[86][481],u_xpb_out[87][481],u_xpb_out[88][481],u_xpb_out[89][481],u_xpb_out[90][481],u_xpb_out[91][481],u_xpb_out[92][481],u_xpb_out[93][481],u_xpb_out[94][481],u_xpb_out[95][481],u_xpb_out[96][481],u_xpb_out[97][481],u_xpb_out[98][481],u_xpb_out[99][481],u_xpb_out[100][481],u_xpb_out[101][481],u_xpb_out[102][481],u_xpb_out[103][481],u_xpb_out[104][481],u_xpb_out[105][481]};

assign col_out_482 = {u_xpb_out[0][482],u_xpb_out[1][482],u_xpb_out[2][482],u_xpb_out[3][482],u_xpb_out[4][482],u_xpb_out[5][482],u_xpb_out[6][482],u_xpb_out[7][482],u_xpb_out[8][482],u_xpb_out[9][482],u_xpb_out[10][482],u_xpb_out[11][482],u_xpb_out[12][482],u_xpb_out[13][482],u_xpb_out[14][482],u_xpb_out[15][482],u_xpb_out[16][482],u_xpb_out[17][482],u_xpb_out[18][482],u_xpb_out[19][482],u_xpb_out[20][482],u_xpb_out[21][482],u_xpb_out[22][482],u_xpb_out[23][482],u_xpb_out[24][482],u_xpb_out[25][482],u_xpb_out[26][482],u_xpb_out[27][482],u_xpb_out[28][482],u_xpb_out[29][482],u_xpb_out[30][482],u_xpb_out[31][482],u_xpb_out[32][482],u_xpb_out[33][482],u_xpb_out[34][482],u_xpb_out[35][482],u_xpb_out[36][482],u_xpb_out[37][482],u_xpb_out[38][482],u_xpb_out[39][482],u_xpb_out[40][482],u_xpb_out[41][482],u_xpb_out[42][482],u_xpb_out[43][482],u_xpb_out[44][482],u_xpb_out[45][482],u_xpb_out[46][482],u_xpb_out[47][482],u_xpb_out[48][482],u_xpb_out[49][482],u_xpb_out[50][482],u_xpb_out[51][482],u_xpb_out[52][482],u_xpb_out[53][482],u_xpb_out[54][482],u_xpb_out[55][482],u_xpb_out[56][482],u_xpb_out[57][482],u_xpb_out[58][482],u_xpb_out[59][482],u_xpb_out[60][482],u_xpb_out[61][482],u_xpb_out[62][482],u_xpb_out[63][482],u_xpb_out[64][482],u_xpb_out[65][482],u_xpb_out[66][482],u_xpb_out[67][482],u_xpb_out[68][482],u_xpb_out[69][482],u_xpb_out[70][482],u_xpb_out[71][482],u_xpb_out[72][482],u_xpb_out[73][482],u_xpb_out[74][482],u_xpb_out[75][482],u_xpb_out[76][482],u_xpb_out[77][482],u_xpb_out[78][482],u_xpb_out[79][482],u_xpb_out[80][482],u_xpb_out[81][482],u_xpb_out[82][482],u_xpb_out[83][482],u_xpb_out[84][482],u_xpb_out[85][482],u_xpb_out[86][482],u_xpb_out[87][482],u_xpb_out[88][482],u_xpb_out[89][482],u_xpb_out[90][482],u_xpb_out[91][482],u_xpb_out[92][482],u_xpb_out[93][482],u_xpb_out[94][482],u_xpb_out[95][482],u_xpb_out[96][482],u_xpb_out[97][482],u_xpb_out[98][482],u_xpb_out[99][482],u_xpb_out[100][482],u_xpb_out[101][482],u_xpb_out[102][482],u_xpb_out[103][482],u_xpb_out[104][482],u_xpb_out[105][482]};

assign col_out_483 = {u_xpb_out[0][483],u_xpb_out[1][483],u_xpb_out[2][483],u_xpb_out[3][483],u_xpb_out[4][483],u_xpb_out[5][483],u_xpb_out[6][483],u_xpb_out[7][483],u_xpb_out[8][483],u_xpb_out[9][483],u_xpb_out[10][483],u_xpb_out[11][483],u_xpb_out[12][483],u_xpb_out[13][483],u_xpb_out[14][483],u_xpb_out[15][483],u_xpb_out[16][483],u_xpb_out[17][483],u_xpb_out[18][483],u_xpb_out[19][483],u_xpb_out[20][483],u_xpb_out[21][483],u_xpb_out[22][483],u_xpb_out[23][483],u_xpb_out[24][483],u_xpb_out[25][483],u_xpb_out[26][483],u_xpb_out[27][483],u_xpb_out[28][483],u_xpb_out[29][483],u_xpb_out[30][483],u_xpb_out[31][483],u_xpb_out[32][483],u_xpb_out[33][483],u_xpb_out[34][483],u_xpb_out[35][483],u_xpb_out[36][483],u_xpb_out[37][483],u_xpb_out[38][483],u_xpb_out[39][483],u_xpb_out[40][483],u_xpb_out[41][483],u_xpb_out[42][483],u_xpb_out[43][483],u_xpb_out[44][483],u_xpb_out[45][483],u_xpb_out[46][483],u_xpb_out[47][483],u_xpb_out[48][483],u_xpb_out[49][483],u_xpb_out[50][483],u_xpb_out[51][483],u_xpb_out[52][483],u_xpb_out[53][483],u_xpb_out[54][483],u_xpb_out[55][483],u_xpb_out[56][483],u_xpb_out[57][483],u_xpb_out[58][483],u_xpb_out[59][483],u_xpb_out[60][483],u_xpb_out[61][483],u_xpb_out[62][483],u_xpb_out[63][483],u_xpb_out[64][483],u_xpb_out[65][483],u_xpb_out[66][483],u_xpb_out[67][483],u_xpb_out[68][483],u_xpb_out[69][483],u_xpb_out[70][483],u_xpb_out[71][483],u_xpb_out[72][483],u_xpb_out[73][483],u_xpb_out[74][483],u_xpb_out[75][483],u_xpb_out[76][483],u_xpb_out[77][483],u_xpb_out[78][483],u_xpb_out[79][483],u_xpb_out[80][483],u_xpb_out[81][483],u_xpb_out[82][483],u_xpb_out[83][483],u_xpb_out[84][483],u_xpb_out[85][483],u_xpb_out[86][483],u_xpb_out[87][483],u_xpb_out[88][483],u_xpb_out[89][483],u_xpb_out[90][483],u_xpb_out[91][483],u_xpb_out[92][483],u_xpb_out[93][483],u_xpb_out[94][483],u_xpb_out[95][483],u_xpb_out[96][483],u_xpb_out[97][483],u_xpb_out[98][483],u_xpb_out[99][483],u_xpb_out[100][483],u_xpb_out[101][483],u_xpb_out[102][483],u_xpb_out[103][483],u_xpb_out[104][483],u_xpb_out[105][483]};

assign col_out_484 = {u_xpb_out[0][484],u_xpb_out[1][484],u_xpb_out[2][484],u_xpb_out[3][484],u_xpb_out[4][484],u_xpb_out[5][484],u_xpb_out[6][484],u_xpb_out[7][484],u_xpb_out[8][484],u_xpb_out[9][484],u_xpb_out[10][484],u_xpb_out[11][484],u_xpb_out[12][484],u_xpb_out[13][484],u_xpb_out[14][484],u_xpb_out[15][484],u_xpb_out[16][484],u_xpb_out[17][484],u_xpb_out[18][484],u_xpb_out[19][484],u_xpb_out[20][484],u_xpb_out[21][484],u_xpb_out[22][484],u_xpb_out[23][484],u_xpb_out[24][484],u_xpb_out[25][484],u_xpb_out[26][484],u_xpb_out[27][484],u_xpb_out[28][484],u_xpb_out[29][484],u_xpb_out[30][484],u_xpb_out[31][484],u_xpb_out[32][484],u_xpb_out[33][484],u_xpb_out[34][484],u_xpb_out[35][484],u_xpb_out[36][484],u_xpb_out[37][484],u_xpb_out[38][484],u_xpb_out[39][484],u_xpb_out[40][484],u_xpb_out[41][484],u_xpb_out[42][484],u_xpb_out[43][484],u_xpb_out[44][484],u_xpb_out[45][484],u_xpb_out[46][484],u_xpb_out[47][484],u_xpb_out[48][484],u_xpb_out[49][484],u_xpb_out[50][484],u_xpb_out[51][484],u_xpb_out[52][484],u_xpb_out[53][484],u_xpb_out[54][484],u_xpb_out[55][484],u_xpb_out[56][484],u_xpb_out[57][484],u_xpb_out[58][484],u_xpb_out[59][484],u_xpb_out[60][484],u_xpb_out[61][484],u_xpb_out[62][484],u_xpb_out[63][484],u_xpb_out[64][484],u_xpb_out[65][484],u_xpb_out[66][484],u_xpb_out[67][484],u_xpb_out[68][484],u_xpb_out[69][484],u_xpb_out[70][484],u_xpb_out[71][484],u_xpb_out[72][484],u_xpb_out[73][484],u_xpb_out[74][484],u_xpb_out[75][484],u_xpb_out[76][484],u_xpb_out[77][484],u_xpb_out[78][484],u_xpb_out[79][484],u_xpb_out[80][484],u_xpb_out[81][484],u_xpb_out[82][484],u_xpb_out[83][484],u_xpb_out[84][484],u_xpb_out[85][484],u_xpb_out[86][484],u_xpb_out[87][484],u_xpb_out[88][484],u_xpb_out[89][484],u_xpb_out[90][484],u_xpb_out[91][484],u_xpb_out[92][484],u_xpb_out[93][484],u_xpb_out[94][484],u_xpb_out[95][484],u_xpb_out[96][484],u_xpb_out[97][484],u_xpb_out[98][484],u_xpb_out[99][484],u_xpb_out[100][484],u_xpb_out[101][484],u_xpb_out[102][484],u_xpb_out[103][484],u_xpb_out[104][484],u_xpb_out[105][484]};

assign col_out_485 = {u_xpb_out[0][485],u_xpb_out[1][485],u_xpb_out[2][485],u_xpb_out[3][485],u_xpb_out[4][485],u_xpb_out[5][485],u_xpb_out[6][485],u_xpb_out[7][485],u_xpb_out[8][485],u_xpb_out[9][485],u_xpb_out[10][485],u_xpb_out[11][485],u_xpb_out[12][485],u_xpb_out[13][485],u_xpb_out[14][485],u_xpb_out[15][485],u_xpb_out[16][485],u_xpb_out[17][485],u_xpb_out[18][485],u_xpb_out[19][485],u_xpb_out[20][485],u_xpb_out[21][485],u_xpb_out[22][485],u_xpb_out[23][485],u_xpb_out[24][485],u_xpb_out[25][485],u_xpb_out[26][485],u_xpb_out[27][485],u_xpb_out[28][485],u_xpb_out[29][485],u_xpb_out[30][485],u_xpb_out[31][485],u_xpb_out[32][485],u_xpb_out[33][485],u_xpb_out[34][485],u_xpb_out[35][485],u_xpb_out[36][485],u_xpb_out[37][485],u_xpb_out[38][485],u_xpb_out[39][485],u_xpb_out[40][485],u_xpb_out[41][485],u_xpb_out[42][485],u_xpb_out[43][485],u_xpb_out[44][485],u_xpb_out[45][485],u_xpb_out[46][485],u_xpb_out[47][485],u_xpb_out[48][485],u_xpb_out[49][485],u_xpb_out[50][485],u_xpb_out[51][485],u_xpb_out[52][485],u_xpb_out[53][485],u_xpb_out[54][485],u_xpb_out[55][485],u_xpb_out[56][485],u_xpb_out[57][485],u_xpb_out[58][485],u_xpb_out[59][485],u_xpb_out[60][485],u_xpb_out[61][485],u_xpb_out[62][485],u_xpb_out[63][485],u_xpb_out[64][485],u_xpb_out[65][485],u_xpb_out[66][485],u_xpb_out[67][485],u_xpb_out[68][485],u_xpb_out[69][485],u_xpb_out[70][485],u_xpb_out[71][485],u_xpb_out[72][485],u_xpb_out[73][485],u_xpb_out[74][485],u_xpb_out[75][485],u_xpb_out[76][485],u_xpb_out[77][485],u_xpb_out[78][485],u_xpb_out[79][485],u_xpb_out[80][485],u_xpb_out[81][485],u_xpb_out[82][485],u_xpb_out[83][485],u_xpb_out[84][485],u_xpb_out[85][485],u_xpb_out[86][485],u_xpb_out[87][485],u_xpb_out[88][485],u_xpb_out[89][485],u_xpb_out[90][485],u_xpb_out[91][485],u_xpb_out[92][485],u_xpb_out[93][485],u_xpb_out[94][485],u_xpb_out[95][485],u_xpb_out[96][485],u_xpb_out[97][485],u_xpb_out[98][485],u_xpb_out[99][485],u_xpb_out[100][485],u_xpb_out[101][485],u_xpb_out[102][485],u_xpb_out[103][485],u_xpb_out[104][485],u_xpb_out[105][485]};

assign col_out_486 = {u_xpb_out[0][486],u_xpb_out[1][486],u_xpb_out[2][486],u_xpb_out[3][486],u_xpb_out[4][486],u_xpb_out[5][486],u_xpb_out[6][486],u_xpb_out[7][486],u_xpb_out[8][486],u_xpb_out[9][486],u_xpb_out[10][486],u_xpb_out[11][486],u_xpb_out[12][486],u_xpb_out[13][486],u_xpb_out[14][486],u_xpb_out[15][486],u_xpb_out[16][486],u_xpb_out[17][486],u_xpb_out[18][486],u_xpb_out[19][486],u_xpb_out[20][486],u_xpb_out[21][486],u_xpb_out[22][486],u_xpb_out[23][486],u_xpb_out[24][486],u_xpb_out[25][486],u_xpb_out[26][486],u_xpb_out[27][486],u_xpb_out[28][486],u_xpb_out[29][486],u_xpb_out[30][486],u_xpb_out[31][486],u_xpb_out[32][486],u_xpb_out[33][486],u_xpb_out[34][486],u_xpb_out[35][486],u_xpb_out[36][486],u_xpb_out[37][486],u_xpb_out[38][486],u_xpb_out[39][486],u_xpb_out[40][486],u_xpb_out[41][486],u_xpb_out[42][486],u_xpb_out[43][486],u_xpb_out[44][486],u_xpb_out[45][486],u_xpb_out[46][486],u_xpb_out[47][486],u_xpb_out[48][486],u_xpb_out[49][486],u_xpb_out[50][486],u_xpb_out[51][486],u_xpb_out[52][486],u_xpb_out[53][486],u_xpb_out[54][486],u_xpb_out[55][486],u_xpb_out[56][486],u_xpb_out[57][486],u_xpb_out[58][486],u_xpb_out[59][486],u_xpb_out[60][486],u_xpb_out[61][486],u_xpb_out[62][486],u_xpb_out[63][486],u_xpb_out[64][486],u_xpb_out[65][486],u_xpb_out[66][486],u_xpb_out[67][486],u_xpb_out[68][486],u_xpb_out[69][486],u_xpb_out[70][486],u_xpb_out[71][486],u_xpb_out[72][486],u_xpb_out[73][486],u_xpb_out[74][486],u_xpb_out[75][486],u_xpb_out[76][486],u_xpb_out[77][486],u_xpb_out[78][486],u_xpb_out[79][486],u_xpb_out[80][486],u_xpb_out[81][486],u_xpb_out[82][486],u_xpb_out[83][486],u_xpb_out[84][486],u_xpb_out[85][486],u_xpb_out[86][486],u_xpb_out[87][486],u_xpb_out[88][486],u_xpb_out[89][486],u_xpb_out[90][486],u_xpb_out[91][486],u_xpb_out[92][486],u_xpb_out[93][486],u_xpb_out[94][486],u_xpb_out[95][486],u_xpb_out[96][486],u_xpb_out[97][486],u_xpb_out[98][486],u_xpb_out[99][486],u_xpb_out[100][486],u_xpb_out[101][486],u_xpb_out[102][486],u_xpb_out[103][486],u_xpb_out[104][486],u_xpb_out[105][486]};

assign col_out_487 = {u_xpb_out[0][487],u_xpb_out[1][487],u_xpb_out[2][487],u_xpb_out[3][487],u_xpb_out[4][487],u_xpb_out[5][487],u_xpb_out[6][487],u_xpb_out[7][487],u_xpb_out[8][487],u_xpb_out[9][487],u_xpb_out[10][487],u_xpb_out[11][487],u_xpb_out[12][487],u_xpb_out[13][487],u_xpb_out[14][487],u_xpb_out[15][487],u_xpb_out[16][487],u_xpb_out[17][487],u_xpb_out[18][487],u_xpb_out[19][487],u_xpb_out[20][487],u_xpb_out[21][487],u_xpb_out[22][487],u_xpb_out[23][487],u_xpb_out[24][487],u_xpb_out[25][487],u_xpb_out[26][487],u_xpb_out[27][487],u_xpb_out[28][487],u_xpb_out[29][487],u_xpb_out[30][487],u_xpb_out[31][487],u_xpb_out[32][487],u_xpb_out[33][487],u_xpb_out[34][487],u_xpb_out[35][487],u_xpb_out[36][487],u_xpb_out[37][487],u_xpb_out[38][487],u_xpb_out[39][487],u_xpb_out[40][487],u_xpb_out[41][487],u_xpb_out[42][487],u_xpb_out[43][487],u_xpb_out[44][487],u_xpb_out[45][487],u_xpb_out[46][487],u_xpb_out[47][487],u_xpb_out[48][487],u_xpb_out[49][487],u_xpb_out[50][487],u_xpb_out[51][487],u_xpb_out[52][487],u_xpb_out[53][487],u_xpb_out[54][487],u_xpb_out[55][487],u_xpb_out[56][487],u_xpb_out[57][487],u_xpb_out[58][487],u_xpb_out[59][487],u_xpb_out[60][487],u_xpb_out[61][487],u_xpb_out[62][487],u_xpb_out[63][487],u_xpb_out[64][487],u_xpb_out[65][487],u_xpb_out[66][487],u_xpb_out[67][487],u_xpb_out[68][487],u_xpb_out[69][487],u_xpb_out[70][487],u_xpb_out[71][487],u_xpb_out[72][487],u_xpb_out[73][487],u_xpb_out[74][487],u_xpb_out[75][487],u_xpb_out[76][487],u_xpb_out[77][487],u_xpb_out[78][487],u_xpb_out[79][487],u_xpb_out[80][487],u_xpb_out[81][487],u_xpb_out[82][487],u_xpb_out[83][487],u_xpb_out[84][487],u_xpb_out[85][487],u_xpb_out[86][487],u_xpb_out[87][487],u_xpb_out[88][487],u_xpb_out[89][487],u_xpb_out[90][487],u_xpb_out[91][487],u_xpb_out[92][487],u_xpb_out[93][487],u_xpb_out[94][487],u_xpb_out[95][487],u_xpb_out[96][487],u_xpb_out[97][487],u_xpb_out[98][487],u_xpb_out[99][487],u_xpb_out[100][487],u_xpb_out[101][487],u_xpb_out[102][487],u_xpb_out[103][487],u_xpb_out[104][487],u_xpb_out[105][487]};

assign col_out_488 = {u_xpb_out[0][488],u_xpb_out[1][488],u_xpb_out[2][488],u_xpb_out[3][488],u_xpb_out[4][488],u_xpb_out[5][488],u_xpb_out[6][488],u_xpb_out[7][488],u_xpb_out[8][488],u_xpb_out[9][488],u_xpb_out[10][488],u_xpb_out[11][488],u_xpb_out[12][488],u_xpb_out[13][488],u_xpb_out[14][488],u_xpb_out[15][488],u_xpb_out[16][488],u_xpb_out[17][488],u_xpb_out[18][488],u_xpb_out[19][488],u_xpb_out[20][488],u_xpb_out[21][488],u_xpb_out[22][488],u_xpb_out[23][488],u_xpb_out[24][488],u_xpb_out[25][488],u_xpb_out[26][488],u_xpb_out[27][488],u_xpb_out[28][488],u_xpb_out[29][488],u_xpb_out[30][488],u_xpb_out[31][488],u_xpb_out[32][488],u_xpb_out[33][488],u_xpb_out[34][488],u_xpb_out[35][488],u_xpb_out[36][488],u_xpb_out[37][488],u_xpb_out[38][488],u_xpb_out[39][488],u_xpb_out[40][488],u_xpb_out[41][488],u_xpb_out[42][488],u_xpb_out[43][488],u_xpb_out[44][488],u_xpb_out[45][488],u_xpb_out[46][488],u_xpb_out[47][488],u_xpb_out[48][488],u_xpb_out[49][488],u_xpb_out[50][488],u_xpb_out[51][488],u_xpb_out[52][488],u_xpb_out[53][488],u_xpb_out[54][488],u_xpb_out[55][488],u_xpb_out[56][488],u_xpb_out[57][488],u_xpb_out[58][488],u_xpb_out[59][488],u_xpb_out[60][488],u_xpb_out[61][488],u_xpb_out[62][488],u_xpb_out[63][488],u_xpb_out[64][488],u_xpb_out[65][488],u_xpb_out[66][488],u_xpb_out[67][488],u_xpb_out[68][488],u_xpb_out[69][488],u_xpb_out[70][488],u_xpb_out[71][488],u_xpb_out[72][488],u_xpb_out[73][488],u_xpb_out[74][488],u_xpb_out[75][488],u_xpb_out[76][488],u_xpb_out[77][488],u_xpb_out[78][488],u_xpb_out[79][488],u_xpb_out[80][488],u_xpb_out[81][488],u_xpb_out[82][488],u_xpb_out[83][488],u_xpb_out[84][488],u_xpb_out[85][488],u_xpb_out[86][488],u_xpb_out[87][488],u_xpb_out[88][488],u_xpb_out[89][488],u_xpb_out[90][488],u_xpb_out[91][488],u_xpb_out[92][488],u_xpb_out[93][488],u_xpb_out[94][488],u_xpb_out[95][488],u_xpb_out[96][488],u_xpb_out[97][488],u_xpb_out[98][488],u_xpb_out[99][488],u_xpb_out[100][488],u_xpb_out[101][488],u_xpb_out[102][488],u_xpb_out[103][488],u_xpb_out[104][488],u_xpb_out[105][488]};

assign col_out_489 = {u_xpb_out[0][489],u_xpb_out[1][489],u_xpb_out[2][489],u_xpb_out[3][489],u_xpb_out[4][489],u_xpb_out[5][489],u_xpb_out[6][489],u_xpb_out[7][489],u_xpb_out[8][489],u_xpb_out[9][489],u_xpb_out[10][489],u_xpb_out[11][489],u_xpb_out[12][489],u_xpb_out[13][489],u_xpb_out[14][489],u_xpb_out[15][489],u_xpb_out[16][489],u_xpb_out[17][489],u_xpb_out[18][489],u_xpb_out[19][489],u_xpb_out[20][489],u_xpb_out[21][489],u_xpb_out[22][489],u_xpb_out[23][489],u_xpb_out[24][489],u_xpb_out[25][489],u_xpb_out[26][489],u_xpb_out[27][489],u_xpb_out[28][489],u_xpb_out[29][489],u_xpb_out[30][489],u_xpb_out[31][489],u_xpb_out[32][489],u_xpb_out[33][489],u_xpb_out[34][489],u_xpb_out[35][489],u_xpb_out[36][489],u_xpb_out[37][489],u_xpb_out[38][489],u_xpb_out[39][489],u_xpb_out[40][489],u_xpb_out[41][489],u_xpb_out[42][489],u_xpb_out[43][489],u_xpb_out[44][489],u_xpb_out[45][489],u_xpb_out[46][489],u_xpb_out[47][489],u_xpb_out[48][489],u_xpb_out[49][489],u_xpb_out[50][489],u_xpb_out[51][489],u_xpb_out[52][489],u_xpb_out[53][489],u_xpb_out[54][489],u_xpb_out[55][489],u_xpb_out[56][489],u_xpb_out[57][489],u_xpb_out[58][489],u_xpb_out[59][489],u_xpb_out[60][489],u_xpb_out[61][489],u_xpb_out[62][489],u_xpb_out[63][489],u_xpb_out[64][489],u_xpb_out[65][489],u_xpb_out[66][489],u_xpb_out[67][489],u_xpb_out[68][489],u_xpb_out[69][489],u_xpb_out[70][489],u_xpb_out[71][489],u_xpb_out[72][489],u_xpb_out[73][489],u_xpb_out[74][489],u_xpb_out[75][489],u_xpb_out[76][489],u_xpb_out[77][489],u_xpb_out[78][489],u_xpb_out[79][489],u_xpb_out[80][489],u_xpb_out[81][489],u_xpb_out[82][489],u_xpb_out[83][489],u_xpb_out[84][489],u_xpb_out[85][489],u_xpb_out[86][489],u_xpb_out[87][489],u_xpb_out[88][489],u_xpb_out[89][489],u_xpb_out[90][489],u_xpb_out[91][489],u_xpb_out[92][489],u_xpb_out[93][489],u_xpb_out[94][489],u_xpb_out[95][489],u_xpb_out[96][489],u_xpb_out[97][489],u_xpb_out[98][489],u_xpb_out[99][489],u_xpb_out[100][489],u_xpb_out[101][489],u_xpb_out[102][489],u_xpb_out[103][489],u_xpb_out[104][489],u_xpb_out[105][489]};

assign col_out_490 = {u_xpb_out[0][490],u_xpb_out[1][490],u_xpb_out[2][490],u_xpb_out[3][490],u_xpb_out[4][490],u_xpb_out[5][490],u_xpb_out[6][490],u_xpb_out[7][490],u_xpb_out[8][490],u_xpb_out[9][490],u_xpb_out[10][490],u_xpb_out[11][490],u_xpb_out[12][490],u_xpb_out[13][490],u_xpb_out[14][490],u_xpb_out[15][490],u_xpb_out[16][490],u_xpb_out[17][490],u_xpb_out[18][490],u_xpb_out[19][490],u_xpb_out[20][490],u_xpb_out[21][490],u_xpb_out[22][490],u_xpb_out[23][490],u_xpb_out[24][490],u_xpb_out[25][490],u_xpb_out[26][490],u_xpb_out[27][490],u_xpb_out[28][490],u_xpb_out[29][490],u_xpb_out[30][490],u_xpb_out[31][490],u_xpb_out[32][490],u_xpb_out[33][490],u_xpb_out[34][490],u_xpb_out[35][490],u_xpb_out[36][490],u_xpb_out[37][490],u_xpb_out[38][490],u_xpb_out[39][490],u_xpb_out[40][490],u_xpb_out[41][490],u_xpb_out[42][490],u_xpb_out[43][490],u_xpb_out[44][490],u_xpb_out[45][490],u_xpb_out[46][490],u_xpb_out[47][490],u_xpb_out[48][490],u_xpb_out[49][490],u_xpb_out[50][490],u_xpb_out[51][490],u_xpb_out[52][490],u_xpb_out[53][490],u_xpb_out[54][490],u_xpb_out[55][490],u_xpb_out[56][490],u_xpb_out[57][490],u_xpb_out[58][490],u_xpb_out[59][490],u_xpb_out[60][490],u_xpb_out[61][490],u_xpb_out[62][490],u_xpb_out[63][490],u_xpb_out[64][490],u_xpb_out[65][490],u_xpb_out[66][490],u_xpb_out[67][490],u_xpb_out[68][490],u_xpb_out[69][490],u_xpb_out[70][490],u_xpb_out[71][490],u_xpb_out[72][490],u_xpb_out[73][490],u_xpb_out[74][490],u_xpb_out[75][490],u_xpb_out[76][490],u_xpb_out[77][490],u_xpb_out[78][490],u_xpb_out[79][490],u_xpb_out[80][490],u_xpb_out[81][490],u_xpb_out[82][490],u_xpb_out[83][490],u_xpb_out[84][490],u_xpb_out[85][490],u_xpb_out[86][490],u_xpb_out[87][490],u_xpb_out[88][490],u_xpb_out[89][490],u_xpb_out[90][490],u_xpb_out[91][490],u_xpb_out[92][490],u_xpb_out[93][490],u_xpb_out[94][490],u_xpb_out[95][490],u_xpb_out[96][490],u_xpb_out[97][490],u_xpb_out[98][490],u_xpb_out[99][490],u_xpb_out[100][490],u_xpb_out[101][490],u_xpb_out[102][490],u_xpb_out[103][490],u_xpb_out[104][490],u_xpb_out[105][490]};

assign col_out_491 = {u_xpb_out[0][491],u_xpb_out[1][491],u_xpb_out[2][491],u_xpb_out[3][491],u_xpb_out[4][491],u_xpb_out[5][491],u_xpb_out[6][491],u_xpb_out[7][491],u_xpb_out[8][491],u_xpb_out[9][491],u_xpb_out[10][491],u_xpb_out[11][491],u_xpb_out[12][491],u_xpb_out[13][491],u_xpb_out[14][491],u_xpb_out[15][491],u_xpb_out[16][491],u_xpb_out[17][491],u_xpb_out[18][491],u_xpb_out[19][491],u_xpb_out[20][491],u_xpb_out[21][491],u_xpb_out[22][491],u_xpb_out[23][491],u_xpb_out[24][491],u_xpb_out[25][491],u_xpb_out[26][491],u_xpb_out[27][491],u_xpb_out[28][491],u_xpb_out[29][491],u_xpb_out[30][491],u_xpb_out[31][491],u_xpb_out[32][491],u_xpb_out[33][491],u_xpb_out[34][491],u_xpb_out[35][491],u_xpb_out[36][491],u_xpb_out[37][491],u_xpb_out[38][491],u_xpb_out[39][491],u_xpb_out[40][491],u_xpb_out[41][491],u_xpb_out[42][491],u_xpb_out[43][491],u_xpb_out[44][491],u_xpb_out[45][491],u_xpb_out[46][491],u_xpb_out[47][491],u_xpb_out[48][491],u_xpb_out[49][491],u_xpb_out[50][491],u_xpb_out[51][491],u_xpb_out[52][491],u_xpb_out[53][491],u_xpb_out[54][491],u_xpb_out[55][491],u_xpb_out[56][491],u_xpb_out[57][491],u_xpb_out[58][491],u_xpb_out[59][491],u_xpb_out[60][491],u_xpb_out[61][491],u_xpb_out[62][491],u_xpb_out[63][491],u_xpb_out[64][491],u_xpb_out[65][491],u_xpb_out[66][491],u_xpb_out[67][491],u_xpb_out[68][491],u_xpb_out[69][491],u_xpb_out[70][491],u_xpb_out[71][491],u_xpb_out[72][491],u_xpb_out[73][491],u_xpb_out[74][491],u_xpb_out[75][491],u_xpb_out[76][491],u_xpb_out[77][491],u_xpb_out[78][491],u_xpb_out[79][491],u_xpb_out[80][491],u_xpb_out[81][491],u_xpb_out[82][491],u_xpb_out[83][491],u_xpb_out[84][491],u_xpb_out[85][491],u_xpb_out[86][491],u_xpb_out[87][491],u_xpb_out[88][491],u_xpb_out[89][491],u_xpb_out[90][491],u_xpb_out[91][491],u_xpb_out[92][491],u_xpb_out[93][491],u_xpb_out[94][491],u_xpb_out[95][491],u_xpb_out[96][491],u_xpb_out[97][491],u_xpb_out[98][491],u_xpb_out[99][491],u_xpb_out[100][491],u_xpb_out[101][491],u_xpb_out[102][491],u_xpb_out[103][491],u_xpb_out[104][491],u_xpb_out[105][491]};

assign col_out_492 = {u_xpb_out[0][492],u_xpb_out[1][492],u_xpb_out[2][492],u_xpb_out[3][492],u_xpb_out[4][492],u_xpb_out[5][492],u_xpb_out[6][492],u_xpb_out[7][492],u_xpb_out[8][492],u_xpb_out[9][492],u_xpb_out[10][492],u_xpb_out[11][492],u_xpb_out[12][492],u_xpb_out[13][492],u_xpb_out[14][492],u_xpb_out[15][492],u_xpb_out[16][492],u_xpb_out[17][492],u_xpb_out[18][492],u_xpb_out[19][492],u_xpb_out[20][492],u_xpb_out[21][492],u_xpb_out[22][492],u_xpb_out[23][492],u_xpb_out[24][492],u_xpb_out[25][492],u_xpb_out[26][492],u_xpb_out[27][492],u_xpb_out[28][492],u_xpb_out[29][492],u_xpb_out[30][492],u_xpb_out[31][492],u_xpb_out[32][492],u_xpb_out[33][492],u_xpb_out[34][492],u_xpb_out[35][492],u_xpb_out[36][492],u_xpb_out[37][492],u_xpb_out[38][492],u_xpb_out[39][492],u_xpb_out[40][492],u_xpb_out[41][492],u_xpb_out[42][492],u_xpb_out[43][492],u_xpb_out[44][492],u_xpb_out[45][492],u_xpb_out[46][492],u_xpb_out[47][492],u_xpb_out[48][492],u_xpb_out[49][492],u_xpb_out[50][492],u_xpb_out[51][492],u_xpb_out[52][492],u_xpb_out[53][492],u_xpb_out[54][492],u_xpb_out[55][492],u_xpb_out[56][492],u_xpb_out[57][492],u_xpb_out[58][492],u_xpb_out[59][492],u_xpb_out[60][492],u_xpb_out[61][492],u_xpb_out[62][492],u_xpb_out[63][492],u_xpb_out[64][492],u_xpb_out[65][492],u_xpb_out[66][492],u_xpb_out[67][492],u_xpb_out[68][492],u_xpb_out[69][492],u_xpb_out[70][492],u_xpb_out[71][492],u_xpb_out[72][492],u_xpb_out[73][492],u_xpb_out[74][492],u_xpb_out[75][492],u_xpb_out[76][492],u_xpb_out[77][492],u_xpb_out[78][492],u_xpb_out[79][492],u_xpb_out[80][492],u_xpb_out[81][492],u_xpb_out[82][492],u_xpb_out[83][492],u_xpb_out[84][492],u_xpb_out[85][492],u_xpb_out[86][492],u_xpb_out[87][492],u_xpb_out[88][492],u_xpb_out[89][492],u_xpb_out[90][492],u_xpb_out[91][492],u_xpb_out[92][492],u_xpb_out[93][492],u_xpb_out[94][492],u_xpb_out[95][492],u_xpb_out[96][492],u_xpb_out[97][492],u_xpb_out[98][492],u_xpb_out[99][492],u_xpb_out[100][492],u_xpb_out[101][492],u_xpb_out[102][492],u_xpb_out[103][492],u_xpb_out[104][492],u_xpb_out[105][492]};

assign col_out_493 = {u_xpb_out[0][493],u_xpb_out[1][493],u_xpb_out[2][493],u_xpb_out[3][493],u_xpb_out[4][493],u_xpb_out[5][493],u_xpb_out[6][493],u_xpb_out[7][493],u_xpb_out[8][493],u_xpb_out[9][493],u_xpb_out[10][493],u_xpb_out[11][493],u_xpb_out[12][493],u_xpb_out[13][493],u_xpb_out[14][493],u_xpb_out[15][493],u_xpb_out[16][493],u_xpb_out[17][493],u_xpb_out[18][493],u_xpb_out[19][493],u_xpb_out[20][493],u_xpb_out[21][493],u_xpb_out[22][493],u_xpb_out[23][493],u_xpb_out[24][493],u_xpb_out[25][493],u_xpb_out[26][493],u_xpb_out[27][493],u_xpb_out[28][493],u_xpb_out[29][493],u_xpb_out[30][493],u_xpb_out[31][493],u_xpb_out[32][493],u_xpb_out[33][493],u_xpb_out[34][493],u_xpb_out[35][493],u_xpb_out[36][493],u_xpb_out[37][493],u_xpb_out[38][493],u_xpb_out[39][493],u_xpb_out[40][493],u_xpb_out[41][493],u_xpb_out[42][493],u_xpb_out[43][493],u_xpb_out[44][493],u_xpb_out[45][493],u_xpb_out[46][493],u_xpb_out[47][493],u_xpb_out[48][493],u_xpb_out[49][493],u_xpb_out[50][493],u_xpb_out[51][493],u_xpb_out[52][493],u_xpb_out[53][493],u_xpb_out[54][493],u_xpb_out[55][493],u_xpb_out[56][493],u_xpb_out[57][493],u_xpb_out[58][493],u_xpb_out[59][493],u_xpb_out[60][493],u_xpb_out[61][493],u_xpb_out[62][493],u_xpb_out[63][493],u_xpb_out[64][493],u_xpb_out[65][493],u_xpb_out[66][493],u_xpb_out[67][493],u_xpb_out[68][493],u_xpb_out[69][493],u_xpb_out[70][493],u_xpb_out[71][493],u_xpb_out[72][493],u_xpb_out[73][493],u_xpb_out[74][493],u_xpb_out[75][493],u_xpb_out[76][493],u_xpb_out[77][493],u_xpb_out[78][493],u_xpb_out[79][493],u_xpb_out[80][493],u_xpb_out[81][493],u_xpb_out[82][493],u_xpb_out[83][493],u_xpb_out[84][493],u_xpb_out[85][493],u_xpb_out[86][493],u_xpb_out[87][493],u_xpb_out[88][493],u_xpb_out[89][493],u_xpb_out[90][493],u_xpb_out[91][493],u_xpb_out[92][493],u_xpb_out[93][493],u_xpb_out[94][493],u_xpb_out[95][493],u_xpb_out[96][493],u_xpb_out[97][493],u_xpb_out[98][493],u_xpb_out[99][493],u_xpb_out[100][493],u_xpb_out[101][493],u_xpb_out[102][493],u_xpb_out[103][493],u_xpb_out[104][493],u_xpb_out[105][493]};

assign col_out_494 = {u_xpb_out[0][494],u_xpb_out[1][494],u_xpb_out[2][494],u_xpb_out[3][494],u_xpb_out[4][494],u_xpb_out[5][494],u_xpb_out[6][494],u_xpb_out[7][494],u_xpb_out[8][494],u_xpb_out[9][494],u_xpb_out[10][494],u_xpb_out[11][494],u_xpb_out[12][494],u_xpb_out[13][494],u_xpb_out[14][494],u_xpb_out[15][494],u_xpb_out[16][494],u_xpb_out[17][494],u_xpb_out[18][494],u_xpb_out[19][494],u_xpb_out[20][494],u_xpb_out[21][494],u_xpb_out[22][494],u_xpb_out[23][494],u_xpb_out[24][494],u_xpb_out[25][494],u_xpb_out[26][494],u_xpb_out[27][494],u_xpb_out[28][494],u_xpb_out[29][494],u_xpb_out[30][494],u_xpb_out[31][494],u_xpb_out[32][494],u_xpb_out[33][494],u_xpb_out[34][494],u_xpb_out[35][494],u_xpb_out[36][494],u_xpb_out[37][494],u_xpb_out[38][494],u_xpb_out[39][494],u_xpb_out[40][494],u_xpb_out[41][494],u_xpb_out[42][494],u_xpb_out[43][494],u_xpb_out[44][494],u_xpb_out[45][494],u_xpb_out[46][494],u_xpb_out[47][494],u_xpb_out[48][494],u_xpb_out[49][494],u_xpb_out[50][494],u_xpb_out[51][494],u_xpb_out[52][494],u_xpb_out[53][494],u_xpb_out[54][494],u_xpb_out[55][494],u_xpb_out[56][494],u_xpb_out[57][494],u_xpb_out[58][494],u_xpb_out[59][494],u_xpb_out[60][494],u_xpb_out[61][494],u_xpb_out[62][494],u_xpb_out[63][494],u_xpb_out[64][494],u_xpb_out[65][494],u_xpb_out[66][494],u_xpb_out[67][494],u_xpb_out[68][494],u_xpb_out[69][494],u_xpb_out[70][494],u_xpb_out[71][494],u_xpb_out[72][494],u_xpb_out[73][494],u_xpb_out[74][494],u_xpb_out[75][494],u_xpb_out[76][494],u_xpb_out[77][494],u_xpb_out[78][494],u_xpb_out[79][494],u_xpb_out[80][494],u_xpb_out[81][494],u_xpb_out[82][494],u_xpb_out[83][494],u_xpb_out[84][494],u_xpb_out[85][494],u_xpb_out[86][494],u_xpb_out[87][494],u_xpb_out[88][494],u_xpb_out[89][494],u_xpb_out[90][494],u_xpb_out[91][494],u_xpb_out[92][494],u_xpb_out[93][494],u_xpb_out[94][494],u_xpb_out[95][494],u_xpb_out[96][494],u_xpb_out[97][494],u_xpb_out[98][494],u_xpb_out[99][494],u_xpb_out[100][494],u_xpb_out[101][494],u_xpb_out[102][494],u_xpb_out[103][494],u_xpb_out[104][494],u_xpb_out[105][494]};

assign col_out_495 = {u_xpb_out[0][495],u_xpb_out[1][495],u_xpb_out[2][495],u_xpb_out[3][495],u_xpb_out[4][495],u_xpb_out[5][495],u_xpb_out[6][495],u_xpb_out[7][495],u_xpb_out[8][495],u_xpb_out[9][495],u_xpb_out[10][495],u_xpb_out[11][495],u_xpb_out[12][495],u_xpb_out[13][495],u_xpb_out[14][495],u_xpb_out[15][495],u_xpb_out[16][495],u_xpb_out[17][495],u_xpb_out[18][495],u_xpb_out[19][495],u_xpb_out[20][495],u_xpb_out[21][495],u_xpb_out[22][495],u_xpb_out[23][495],u_xpb_out[24][495],u_xpb_out[25][495],u_xpb_out[26][495],u_xpb_out[27][495],u_xpb_out[28][495],u_xpb_out[29][495],u_xpb_out[30][495],u_xpb_out[31][495],u_xpb_out[32][495],u_xpb_out[33][495],u_xpb_out[34][495],u_xpb_out[35][495],u_xpb_out[36][495],u_xpb_out[37][495],u_xpb_out[38][495],u_xpb_out[39][495],u_xpb_out[40][495],u_xpb_out[41][495],u_xpb_out[42][495],u_xpb_out[43][495],u_xpb_out[44][495],u_xpb_out[45][495],u_xpb_out[46][495],u_xpb_out[47][495],u_xpb_out[48][495],u_xpb_out[49][495],u_xpb_out[50][495],u_xpb_out[51][495],u_xpb_out[52][495],u_xpb_out[53][495],u_xpb_out[54][495],u_xpb_out[55][495],u_xpb_out[56][495],u_xpb_out[57][495],u_xpb_out[58][495],u_xpb_out[59][495],u_xpb_out[60][495],u_xpb_out[61][495],u_xpb_out[62][495],u_xpb_out[63][495],u_xpb_out[64][495],u_xpb_out[65][495],u_xpb_out[66][495],u_xpb_out[67][495],u_xpb_out[68][495],u_xpb_out[69][495],u_xpb_out[70][495],u_xpb_out[71][495],u_xpb_out[72][495],u_xpb_out[73][495],u_xpb_out[74][495],u_xpb_out[75][495],u_xpb_out[76][495],u_xpb_out[77][495],u_xpb_out[78][495],u_xpb_out[79][495],u_xpb_out[80][495],u_xpb_out[81][495],u_xpb_out[82][495],u_xpb_out[83][495],u_xpb_out[84][495],u_xpb_out[85][495],u_xpb_out[86][495],u_xpb_out[87][495],u_xpb_out[88][495],u_xpb_out[89][495],u_xpb_out[90][495],u_xpb_out[91][495],u_xpb_out[92][495],u_xpb_out[93][495],u_xpb_out[94][495],u_xpb_out[95][495],u_xpb_out[96][495],u_xpb_out[97][495],u_xpb_out[98][495],u_xpb_out[99][495],u_xpb_out[100][495],u_xpb_out[101][495],u_xpb_out[102][495],u_xpb_out[103][495],u_xpb_out[104][495],u_xpb_out[105][495]};

assign col_out_496 = {u_xpb_out[0][496],u_xpb_out[1][496],u_xpb_out[2][496],u_xpb_out[3][496],u_xpb_out[4][496],u_xpb_out[5][496],u_xpb_out[6][496],u_xpb_out[7][496],u_xpb_out[8][496],u_xpb_out[9][496],u_xpb_out[10][496],u_xpb_out[11][496],u_xpb_out[12][496],u_xpb_out[13][496],u_xpb_out[14][496],u_xpb_out[15][496],u_xpb_out[16][496],u_xpb_out[17][496],u_xpb_out[18][496],u_xpb_out[19][496],u_xpb_out[20][496],u_xpb_out[21][496],u_xpb_out[22][496],u_xpb_out[23][496],u_xpb_out[24][496],u_xpb_out[25][496],u_xpb_out[26][496],u_xpb_out[27][496],u_xpb_out[28][496],u_xpb_out[29][496],u_xpb_out[30][496],u_xpb_out[31][496],u_xpb_out[32][496],u_xpb_out[33][496],u_xpb_out[34][496],u_xpb_out[35][496],u_xpb_out[36][496],u_xpb_out[37][496],u_xpb_out[38][496],u_xpb_out[39][496],u_xpb_out[40][496],u_xpb_out[41][496],u_xpb_out[42][496],u_xpb_out[43][496],u_xpb_out[44][496],u_xpb_out[45][496],u_xpb_out[46][496],u_xpb_out[47][496],u_xpb_out[48][496],u_xpb_out[49][496],u_xpb_out[50][496],u_xpb_out[51][496],u_xpb_out[52][496],u_xpb_out[53][496],u_xpb_out[54][496],u_xpb_out[55][496],u_xpb_out[56][496],u_xpb_out[57][496],u_xpb_out[58][496],u_xpb_out[59][496],u_xpb_out[60][496],u_xpb_out[61][496],u_xpb_out[62][496],u_xpb_out[63][496],u_xpb_out[64][496],u_xpb_out[65][496],u_xpb_out[66][496],u_xpb_out[67][496],u_xpb_out[68][496],u_xpb_out[69][496],u_xpb_out[70][496],u_xpb_out[71][496],u_xpb_out[72][496],u_xpb_out[73][496],u_xpb_out[74][496],u_xpb_out[75][496],u_xpb_out[76][496],u_xpb_out[77][496],u_xpb_out[78][496],u_xpb_out[79][496],u_xpb_out[80][496],u_xpb_out[81][496],u_xpb_out[82][496],u_xpb_out[83][496],u_xpb_out[84][496],u_xpb_out[85][496],u_xpb_out[86][496],u_xpb_out[87][496],u_xpb_out[88][496],u_xpb_out[89][496],u_xpb_out[90][496],u_xpb_out[91][496],u_xpb_out[92][496],u_xpb_out[93][496],u_xpb_out[94][496],u_xpb_out[95][496],u_xpb_out[96][496],u_xpb_out[97][496],u_xpb_out[98][496],u_xpb_out[99][496],u_xpb_out[100][496],u_xpb_out[101][496],u_xpb_out[102][496],u_xpb_out[103][496],u_xpb_out[104][496],u_xpb_out[105][496]};

assign col_out_497 = {u_xpb_out[0][497],u_xpb_out[1][497],u_xpb_out[2][497],u_xpb_out[3][497],u_xpb_out[4][497],u_xpb_out[5][497],u_xpb_out[6][497],u_xpb_out[7][497],u_xpb_out[8][497],u_xpb_out[9][497],u_xpb_out[10][497],u_xpb_out[11][497],u_xpb_out[12][497],u_xpb_out[13][497],u_xpb_out[14][497],u_xpb_out[15][497],u_xpb_out[16][497],u_xpb_out[17][497],u_xpb_out[18][497],u_xpb_out[19][497],u_xpb_out[20][497],u_xpb_out[21][497],u_xpb_out[22][497],u_xpb_out[23][497],u_xpb_out[24][497],u_xpb_out[25][497],u_xpb_out[26][497],u_xpb_out[27][497],u_xpb_out[28][497],u_xpb_out[29][497],u_xpb_out[30][497],u_xpb_out[31][497],u_xpb_out[32][497],u_xpb_out[33][497],u_xpb_out[34][497],u_xpb_out[35][497],u_xpb_out[36][497],u_xpb_out[37][497],u_xpb_out[38][497],u_xpb_out[39][497],u_xpb_out[40][497],u_xpb_out[41][497],u_xpb_out[42][497],u_xpb_out[43][497],u_xpb_out[44][497],u_xpb_out[45][497],u_xpb_out[46][497],u_xpb_out[47][497],u_xpb_out[48][497],u_xpb_out[49][497],u_xpb_out[50][497],u_xpb_out[51][497],u_xpb_out[52][497],u_xpb_out[53][497],u_xpb_out[54][497],u_xpb_out[55][497],u_xpb_out[56][497],u_xpb_out[57][497],u_xpb_out[58][497],u_xpb_out[59][497],u_xpb_out[60][497],u_xpb_out[61][497],u_xpb_out[62][497],u_xpb_out[63][497],u_xpb_out[64][497],u_xpb_out[65][497],u_xpb_out[66][497],u_xpb_out[67][497],u_xpb_out[68][497],u_xpb_out[69][497],u_xpb_out[70][497],u_xpb_out[71][497],u_xpb_out[72][497],u_xpb_out[73][497],u_xpb_out[74][497],u_xpb_out[75][497],u_xpb_out[76][497],u_xpb_out[77][497],u_xpb_out[78][497],u_xpb_out[79][497],u_xpb_out[80][497],u_xpb_out[81][497],u_xpb_out[82][497],u_xpb_out[83][497],u_xpb_out[84][497],u_xpb_out[85][497],u_xpb_out[86][497],u_xpb_out[87][497],u_xpb_out[88][497],u_xpb_out[89][497],u_xpb_out[90][497],u_xpb_out[91][497],u_xpb_out[92][497],u_xpb_out[93][497],u_xpb_out[94][497],u_xpb_out[95][497],u_xpb_out[96][497],u_xpb_out[97][497],u_xpb_out[98][497],u_xpb_out[99][497],u_xpb_out[100][497],u_xpb_out[101][497],u_xpb_out[102][497],u_xpb_out[103][497],u_xpb_out[104][497],u_xpb_out[105][497]};

assign col_out_498 = {u_xpb_out[0][498],u_xpb_out[1][498],u_xpb_out[2][498],u_xpb_out[3][498],u_xpb_out[4][498],u_xpb_out[5][498],u_xpb_out[6][498],u_xpb_out[7][498],u_xpb_out[8][498],u_xpb_out[9][498],u_xpb_out[10][498],u_xpb_out[11][498],u_xpb_out[12][498],u_xpb_out[13][498],u_xpb_out[14][498],u_xpb_out[15][498],u_xpb_out[16][498],u_xpb_out[17][498],u_xpb_out[18][498],u_xpb_out[19][498],u_xpb_out[20][498],u_xpb_out[21][498],u_xpb_out[22][498],u_xpb_out[23][498],u_xpb_out[24][498],u_xpb_out[25][498],u_xpb_out[26][498],u_xpb_out[27][498],u_xpb_out[28][498],u_xpb_out[29][498],u_xpb_out[30][498],u_xpb_out[31][498],u_xpb_out[32][498],u_xpb_out[33][498],u_xpb_out[34][498],u_xpb_out[35][498],u_xpb_out[36][498],u_xpb_out[37][498],u_xpb_out[38][498],u_xpb_out[39][498],u_xpb_out[40][498],u_xpb_out[41][498],u_xpb_out[42][498],u_xpb_out[43][498],u_xpb_out[44][498],u_xpb_out[45][498],u_xpb_out[46][498],u_xpb_out[47][498],u_xpb_out[48][498],u_xpb_out[49][498],u_xpb_out[50][498],u_xpb_out[51][498],u_xpb_out[52][498],u_xpb_out[53][498],u_xpb_out[54][498],u_xpb_out[55][498],u_xpb_out[56][498],u_xpb_out[57][498],u_xpb_out[58][498],u_xpb_out[59][498],u_xpb_out[60][498],u_xpb_out[61][498],u_xpb_out[62][498],u_xpb_out[63][498],u_xpb_out[64][498],u_xpb_out[65][498],u_xpb_out[66][498],u_xpb_out[67][498],u_xpb_out[68][498],u_xpb_out[69][498],u_xpb_out[70][498],u_xpb_out[71][498],u_xpb_out[72][498],u_xpb_out[73][498],u_xpb_out[74][498],u_xpb_out[75][498],u_xpb_out[76][498],u_xpb_out[77][498],u_xpb_out[78][498],u_xpb_out[79][498],u_xpb_out[80][498],u_xpb_out[81][498],u_xpb_out[82][498],u_xpb_out[83][498],u_xpb_out[84][498],u_xpb_out[85][498],u_xpb_out[86][498],u_xpb_out[87][498],u_xpb_out[88][498],u_xpb_out[89][498],u_xpb_out[90][498],u_xpb_out[91][498],u_xpb_out[92][498],u_xpb_out[93][498],u_xpb_out[94][498],u_xpb_out[95][498],u_xpb_out[96][498],u_xpb_out[97][498],u_xpb_out[98][498],u_xpb_out[99][498],u_xpb_out[100][498],u_xpb_out[101][498],u_xpb_out[102][498],u_xpb_out[103][498],u_xpb_out[104][498],u_xpb_out[105][498]};

assign col_out_499 = {u_xpb_out[0][499],u_xpb_out[1][499],u_xpb_out[2][499],u_xpb_out[3][499],u_xpb_out[4][499],u_xpb_out[5][499],u_xpb_out[6][499],u_xpb_out[7][499],u_xpb_out[8][499],u_xpb_out[9][499],u_xpb_out[10][499],u_xpb_out[11][499],u_xpb_out[12][499],u_xpb_out[13][499],u_xpb_out[14][499],u_xpb_out[15][499],u_xpb_out[16][499],u_xpb_out[17][499],u_xpb_out[18][499],u_xpb_out[19][499],u_xpb_out[20][499],u_xpb_out[21][499],u_xpb_out[22][499],u_xpb_out[23][499],u_xpb_out[24][499],u_xpb_out[25][499],u_xpb_out[26][499],u_xpb_out[27][499],u_xpb_out[28][499],u_xpb_out[29][499],u_xpb_out[30][499],u_xpb_out[31][499],u_xpb_out[32][499],u_xpb_out[33][499],u_xpb_out[34][499],u_xpb_out[35][499],u_xpb_out[36][499],u_xpb_out[37][499],u_xpb_out[38][499],u_xpb_out[39][499],u_xpb_out[40][499],u_xpb_out[41][499],u_xpb_out[42][499],u_xpb_out[43][499],u_xpb_out[44][499],u_xpb_out[45][499],u_xpb_out[46][499],u_xpb_out[47][499],u_xpb_out[48][499],u_xpb_out[49][499],u_xpb_out[50][499],u_xpb_out[51][499],u_xpb_out[52][499],u_xpb_out[53][499],u_xpb_out[54][499],u_xpb_out[55][499],u_xpb_out[56][499],u_xpb_out[57][499],u_xpb_out[58][499],u_xpb_out[59][499],u_xpb_out[60][499],u_xpb_out[61][499],u_xpb_out[62][499],u_xpb_out[63][499],u_xpb_out[64][499],u_xpb_out[65][499],u_xpb_out[66][499],u_xpb_out[67][499],u_xpb_out[68][499],u_xpb_out[69][499],u_xpb_out[70][499],u_xpb_out[71][499],u_xpb_out[72][499],u_xpb_out[73][499],u_xpb_out[74][499],u_xpb_out[75][499],u_xpb_out[76][499],u_xpb_out[77][499],u_xpb_out[78][499],u_xpb_out[79][499],u_xpb_out[80][499],u_xpb_out[81][499],u_xpb_out[82][499],u_xpb_out[83][499],u_xpb_out[84][499],u_xpb_out[85][499],u_xpb_out[86][499],u_xpb_out[87][499],u_xpb_out[88][499],u_xpb_out[89][499],u_xpb_out[90][499],u_xpb_out[91][499],u_xpb_out[92][499],u_xpb_out[93][499],u_xpb_out[94][499],u_xpb_out[95][499],u_xpb_out[96][499],u_xpb_out[97][499],u_xpb_out[98][499],u_xpb_out[99][499],u_xpb_out[100][499],u_xpb_out[101][499],u_xpb_out[102][499],u_xpb_out[103][499],u_xpb_out[104][499],u_xpb_out[105][499]};

assign col_out_500 = {u_xpb_out[0][500],u_xpb_out[1][500],u_xpb_out[2][500],u_xpb_out[3][500],u_xpb_out[4][500],u_xpb_out[5][500],u_xpb_out[6][500],u_xpb_out[7][500],u_xpb_out[8][500],u_xpb_out[9][500],u_xpb_out[10][500],u_xpb_out[11][500],u_xpb_out[12][500],u_xpb_out[13][500],u_xpb_out[14][500],u_xpb_out[15][500],u_xpb_out[16][500],u_xpb_out[17][500],u_xpb_out[18][500],u_xpb_out[19][500],u_xpb_out[20][500],u_xpb_out[21][500],u_xpb_out[22][500],u_xpb_out[23][500],u_xpb_out[24][500],u_xpb_out[25][500],u_xpb_out[26][500],u_xpb_out[27][500],u_xpb_out[28][500],u_xpb_out[29][500],u_xpb_out[30][500],u_xpb_out[31][500],u_xpb_out[32][500],u_xpb_out[33][500],u_xpb_out[34][500],u_xpb_out[35][500],u_xpb_out[36][500],u_xpb_out[37][500],u_xpb_out[38][500],u_xpb_out[39][500],u_xpb_out[40][500],u_xpb_out[41][500],u_xpb_out[42][500],u_xpb_out[43][500],u_xpb_out[44][500],u_xpb_out[45][500],u_xpb_out[46][500],u_xpb_out[47][500],u_xpb_out[48][500],u_xpb_out[49][500],u_xpb_out[50][500],u_xpb_out[51][500],u_xpb_out[52][500],u_xpb_out[53][500],u_xpb_out[54][500],u_xpb_out[55][500],u_xpb_out[56][500],u_xpb_out[57][500],u_xpb_out[58][500],u_xpb_out[59][500],u_xpb_out[60][500],u_xpb_out[61][500],u_xpb_out[62][500],u_xpb_out[63][500],u_xpb_out[64][500],u_xpb_out[65][500],u_xpb_out[66][500],u_xpb_out[67][500],u_xpb_out[68][500],u_xpb_out[69][500],u_xpb_out[70][500],u_xpb_out[71][500],u_xpb_out[72][500],u_xpb_out[73][500],u_xpb_out[74][500],u_xpb_out[75][500],u_xpb_out[76][500],u_xpb_out[77][500],u_xpb_out[78][500],u_xpb_out[79][500],u_xpb_out[80][500],u_xpb_out[81][500],u_xpb_out[82][500],u_xpb_out[83][500],u_xpb_out[84][500],u_xpb_out[85][500],u_xpb_out[86][500],u_xpb_out[87][500],u_xpb_out[88][500],u_xpb_out[89][500],u_xpb_out[90][500],u_xpb_out[91][500],u_xpb_out[92][500],u_xpb_out[93][500],u_xpb_out[94][500],u_xpb_out[95][500],u_xpb_out[96][500],u_xpb_out[97][500],u_xpb_out[98][500],u_xpb_out[99][500],u_xpb_out[100][500],u_xpb_out[101][500],u_xpb_out[102][500],u_xpb_out[103][500],u_xpb_out[104][500],u_xpb_out[105][500]};

assign col_out_501 = {u_xpb_out[0][501],u_xpb_out[1][501],u_xpb_out[2][501],u_xpb_out[3][501],u_xpb_out[4][501],u_xpb_out[5][501],u_xpb_out[6][501],u_xpb_out[7][501],u_xpb_out[8][501],u_xpb_out[9][501],u_xpb_out[10][501],u_xpb_out[11][501],u_xpb_out[12][501],u_xpb_out[13][501],u_xpb_out[14][501],u_xpb_out[15][501],u_xpb_out[16][501],u_xpb_out[17][501],u_xpb_out[18][501],u_xpb_out[19][501],u_xpb_out[20][501],u_xpb_out[21][501],u_xpb_out[22][501],u_xpb_out[23][501],u_xpb_out[24][501],u_xpb_out[25][501],u_xpb_out[26][501],u_xpb_out[27][501],u_xpb_out[28][501],u_xpb_out[29][501],u_xpb_out[30][501],u_xpb_out[31][501],u_xpb_out[32][501],u_xpb_out[33][501],u_xpb_out[34][501],u_xpb_out[35][501],u_xpb_out[36][501],u_xpb_out[37][501],u_xpb_out[38][501],u_xpb_out[39][501],u_xpb_out[40][501],u_xpb_out[41][501],u_xpb_out[42][501],u_xpb_out[43][501],u_xpb_out[44][501],u_xpb_out[45][501],u_xpb_out[46][501],u_xpb_out[47][501],u_xpb_out[48][501],u_xpb_out[49][501],u_xpb_out[50][501],u_xpb_out[51][501],u_xpb_out[52][501],u_xpb_out[53][501],u_xpb_out[54][501],u_xpb_out[55][501],u_xpb_out[56][501],u_xpb_out[57][501],u_xpb_out[58][501],u_xpb_out[59][501],u_xpb_out[60][501],u_xpb_out[61][501],u_xpb_out[62][501],u_xpb_out[63][501],u_xpb_out[64][501],u_xpb_out[65][501],u_xpb_out[66][501],u_xpb_out[67][501],u_xpb_out[68][501],u_xpb_out[69][501],u_xpb_out[70][501],u_xpb_out[71][501],u_xpb_out[72][501],u_xpb_out[73][501],u_xpb_out[74][501],u_xpb_out[75][501],u_xpb_out[76][501],u_xpb_out[77][501],u_xpb_out[78][501],u_xpb_out[79][501],u_xpb_out[80][501],u_xpb_out[81][501],u_xpb_out[82][501],u_xpb_out[83][501],u_xpb_out[84][501],u_xpb_out[85][501],u_xpb_out[86][501],u_xpb_out[87][501],u_xpb_out[88][501],u_xpb_out[89][501],u_xpb_out[90][501],u_xpb_out[91][501],u_xpb_out[92][501],u_xpb_out[93][501],u_xpb_out[94][501],u_xpb_out[95][501],u_xpb_out[96][501],u_xpb_out[97][501],u_xpb_out[98][501],u_xpb_out[99][501],u_xpb_out[100][501],u_xpb_out[101][501],u_xpb_out[102][501],u_xpb_out[103][501],u_xpb_out[104][501],u_xpb_out[105][501]};

assign col_out_502 = {u_xpb_out[0][502],u_xpb_out[1][502],u_xpb_out[2][502],u_xpb_out[3][502],u_xpb_out[4][502],u_xpb_out[5][502],u_xpb_out[6][502],u_xpb_out[7][502],u_xpb_out[8][502],u_xpb_out[9][502],u_xpb_out[10][502],u_xpb_out[11][502],u_xpb_out[12][502],u_xpb_out[13][502],u_xpb_out[14][502],u_xpb_out[15][502],u_xpb_out[16][502],u_xpb_out[17][502],u_xpb_out[18][502],u_xpb_out[19][502],u_xpb_out[20][502],u_xpb_out[21][502],u_xpb_out[22][502],u_xpb_out[23][502],u_xpb_out[24][502],u_xpb_out[25][502],u_xpb_out[26][502],u_xpb_out[27][502],u_xpb_out[28][502],u_xpb_out[29][502],u_xpb_out[30][502],u_xpb_out[31][502],u_xpb_out[32][502],u_xpb_out[33][502],u_xpb_out[34][502],u_xpb_out[35][502],u_xpb_out[36][502],u_xpb_out[37][502],u_xpb_out[38][502],u_xpb_out[39][502],u_xpb_out[40][502],u_xpb_out[41][502],u_xpb_out[42][502],u_xpb_out[43][502],u_xpb_out[44][502],u_xpb_out[45][502],u_xpb_out[46][502],u_xpb_out[47][502],u_xpb_out[48][502],u_xpb_out[49][502],u_xpb_out[50][502],u_xpb_out[51][502],u_xpb_out[52][502],u_xpb_out[53][502],u_xpb_out[54][502],u_xpb_out[55][502],u_xpb_out[56][502],u_xpb_out[57][502],u_xpb_out[58][502],u_xpb_out[59][502],u_xpb_out[60][502],u_xpb_out[61][502],u_xpb_out[62][502],u_xpb_out[63][502],u_xpb_out[64][502],u_xpb_out[65][502],u_xpb_out[66][502],u_xpb_out[67][502],u_xpb_out[68][502],u_xpb_out[69][502],u_xpb_out[70][502],u_xpb_out[71][502],u_xpb_out[72][502],u_xpb_out[73][502],u_xpb_out[74][502],u_xpb_out[75][502],u_xpb_out[76][502],u_xpb_out[77][502],u_xpb_out[78][502],u_xpb_out[79][502],u_xpb_out[80][502],u_xpb_out[81][502],u_xpb_out[82][502],u_xpb_out[83][502],u_xpb_out[84][502],u_xpb_out[85][502],u_xpb_out[86][502],u_xpb_out[87][502],u_xpb_out[88][502],u_xpb_out[89][502],u_xpb_out[90][502],u_xpb_out[91][502],u_xpb_out[92][502],u_xpb_out[93][502],u_xpb_out[94][502],u_xpb_out[95][502],u_xpb_out[96][502],u_xpb_out[97][502],u_xpb_out[98][502],u_xpb_out[99][502],u_xpb_out[100][502],u_xpb_out[101][502],u_xpb_out[102][502],u_xpb_out[103][502],u_xpb_out[104][502],u_xpb_out[105][502]};

assign col_out_503 = {u_xpb_out[0][503],u_xpb_out[1][503],u_xpb_out[2][503],u_xpb_out[3][503],u_xpb_out[4][503],u_xpb_out[5][503],u_xpb_out[6][503],u_xpb_out[7][503],u_xpb_out[8][503],u_xpb_out[9][503],u_xpb_out[10][503],u_xpb_out[11][503],u_xpb_out[12][503],u_xpb_out[13][503],u_xpb_out[14][503],u_xpb_out[15][503],u_xpb_out[16][503],u_xpb_out[17][503],u_xpb_out[18][503],u_xpb_out[19][503],u_xpb_out[20][503],u_xpb_out[21][503],u_xpb_out[22][503],u_xpb_out[23][503],u_xpb_out[24][503],u_xpb_out[25][503],u_xpb_out[26][503],u_xpb_out[27][503],u_xpb_out[28][503],u_xpb_out[29][503],u_xpb_out[30][503],u_xpb_out[31][503],u_xpb_out[32][503],u_xpb_out[33][503],u_xpb_out[34][503],u_xpb_out[35][503],u_xpb_out[36][503],u_xpb_out[37][503],u_xpb_out[38][503],u_xpb_out[39][503],u_xpb_out[40][503],u_xpb_out[41][503],u_xpb_out[42][503],u_xpb_out[43][503],u_xpb_out[44][503],u_xpb_out[45][503],u_xpb_out[46][503],u_xpb_out[47][503],u_xpb_out[48][503],u_xpb_out[49][503],u_xpb_out[50][503],u_xpb_out[51][503],u_xpb_out[52][503],u_xpb_out[53][503],u_xpb_out[54][503],u_xpb_out[55][503],u_xpb_out[56][503],u_xpb_out[57][503],u_xpb_out[58][503],u_xpb_out[59][503],u_xpb_out[60][503],u_xpb_out[61][503],u_xpb_out[62][503],u_xpb_out[63][503],u_xpb_out[64][503],u_xpb_out[65][503],u_xpb_out[66][503],u_xpb_out[67][503],u_xpb_out[68][503],u_xpb_out[69][503],u_xpb_out[70][503],u_xpb_out[71][503],u_xpb_out[72][503],u_xpb_out[73][503],u_xpb_out[74][503],u_xpb_out[75][503],u_xpb_out[76][503],u_xpb_out[77][503],u_xpb_out[78][503],u_xpb_out[79][503],u_xpb_out[80][503],u_xpb_out[81][503],u_xpb_out[82][503],u_xpb_out[83][503],u_xpb_out[84][503],u_xpb_out[85][503],u_xpb_out[86][503],u_xpb_out[87][503],u_xpb_out[88][503],u_xpb_out[89][503],u_xpb_out[90][503],u_xpb_out[91][503],u_xpb_out[92][503],u_xpb_out[93][503],u_xpb_out[94][503],u_xpb_out[95][503],u_xpb_out[96][503],u_xpb_out[97][503],u_xpb_out[98][503],u_xpb_out[99][503],u_xpb_out[100][503],u_xpb_out[101][503],u_xpb_out[102][503],u_xpb_out[103][503],u_xpb_out[104][503],u_xpb_out[105][503]};

assign col_out_504 = {u_xpb_out[0][504],u_xpb_out[1][504],u_xpb_out[2][504],u_xpb_out[3][504],u_xpb_out[4][504],u_xpb_out[5][504],u_xpb_out[6][504],u_xpb_out[7][504],u_xpb_out[8][504],u_xpb_out[9][504],u_xpb_out[10][504],u_xpb_out[11][504],u_xpb_out[12][504],u_xpb_out[13][504],u_xpb_out[14][504],u_xpb_out[15][504],u_xpb_out[16][504],u_xpb_out[17][504],u_xpb_out[18][504],u_xpb_out[19][504],u_xpb_out[20][504],u_xpb_out[21][504],u_xpb_out[22][504],u_xpb_out[23][504],u_xpb_out[24][504],u_xpb_out[25][504],u_xpb_out[26][504],u_xpb_out[27][504],u_xpb_out[28][504],u_xpb_out[29][504],u_xpb_out[30][504],u_xpb_out[31][504],u_xpb_out[32][504],u_xpb_out[33][504],u_xpb_out[34][504],u_xpb_out[35][504],u_xpb_out[36][504],u_xpb_out[37][504],u_xpb_out[38][504],u_xpb_out[39][504],u_xpb_out[40][504],u_xpb_out[41][504],u_xpb_out[42][504],u_xpb_out[43][504],u_xpb_out[44][504],u_xpb_out[45][504],u_xpb_out[46][504],u_xpb_out[47][504],u_xpb_out[48][504],u_xpb_out[49][504],u_xpb_out[50][504],u_xpb_out[51][504],u_xpb_out[52][504],u_xpb_out[53][504],u_xpb_out[54][504],u_xpb_out[55][504],u_xpb_out[56][504],u_xpb_out[57][504],u_xpb_out[58][504],u_xpb_out[59][504],u_xpb_out[60][504],u_xpb_out[61][504],u_xpb_out[62][504],u_xpb_out[63][504],u_xpb_out[64][504],u_xpb_out[65][504],u_xpb_out[66][504],u_xpb_out[67][504],u_xpb_out[68][504],u_xpb_out[69][504],u_xpb_out[70][504],u_xpb_out[71][504],u_xpb_out[72][504],u_xpb_out[73][504],u_xpb_out[74][504],u_xpb_out[75][504],u_xpb_out[76][504],u_xpb_out[77][504],u_xpb_out[78][504],u_xpb_out[79][504],u_xpb_out[80][504],u_xpb_out[81][504],u_xpb_out[82][504],u_xpb_out[83][504],u_xpb_out[84][504],u_xpb_out[85][504],u_xpb_out[86][504],u_xpb_out[87][504],u_xpb_out[88][504],u_xpb_out[89][504],u_xpb_out[90][504],u_xpb_out[91][504],u_xpb_out[92][504],u_xpb_out[93][504],u_xpb_out[94][504],u_xpb_out[95][504],u_xpb_out[96][504],u_xpb_out[97][504],u_xpb_out[98][504],u_xpb_out[99][504],u_xpb_out[100][504],u_xpb_out[101][504],u_xpb_out[102][504],u_xpb_out[103][504],u_xpb_out[104][504],u_xpb_out[105][504]};

assign col_out_505 = {u_xpb_out[0][505],u_xpb_out[1][505],u_xpb_out[2][505],u_xpb_out[3][505],u_xpb_out[4][505],u_xpb_out[5][505],u_xpb_out[6][505],u_xpb_out[7][505],u_xpb_out[8][505],u_xpb_out[9][505],u_xpb_out[10][505],u_xpb_out[11][505],u_xpb_out[12][505],u_xpb_out[13][505],u_xpb_out[14][505],u_xpb_out[15][505],u_xpb_out[16][505],u_xpb_out[17][505],u_xpb_out[18][505],u_xpb_out[19][505],u_xpb_out[20][505],u_xpb_out[21][505],u_xpb_out[22][505],u_xpb_out[23][505],u_xpb_out[24][505],u_xpb_out[25][505],u_xpb_out[26][505],u_xpb_out[27][505],u_xpb_out[28][505],u_xpb_out[29][505],u_xpb_out[30][505],u_xpb_out[31][505],u_xpb_out[32][505],u_xpb_out[33][505],u_xpb_out[34][505],u_xpb_out[35][505],u_xpb_out[36][505],u_xpb_out[37][505],u_xpb_out[38][505],u_xpb_out[39][505],u_xpb_out[40][505],u_xpb_out[41][505],u_xpb_out[42][505],u_xpb_out[43][505],u_xpb_out[44][505],u_xpb_out[45][505],u_xpb_out[46][505],u_xpb_out[47][505],u_xpb_out[48][505],u_xpb_out[49][505],u_xpb_out[50][505],u_xpb_out[51][505],u_xpb_out[52][505],u_xpb_out[53][505],u_xpb_out[54][505],u_xpb_out[55][505],u_xpb_out[56][505],u_xpb_out[57][505],u_xpb_out[58][505],u_xpb_out[59][505],u_xpb_out[60][505],u_xpb_out[61][505],u_xpb_out[62][505],u_xpb_out[63][505],u_xpb_out[64][505],u_xpb_out[65][505],u_xpb_out[66][505],u_xpb_out[67][505],u_xpb_out[68][505],u_xpb_out[69][505],u_xpb_out[70][505],u_xpb_out[71][505],u_xpb_out[72][505],u_xpb_out[73][505],u_xpb_out[74][505],u_xpb_out[75][505],u_xpb_out[76][505],u_xpb_out[77][505],u_xpb_out[78][505],u_xpb_out[79][505],u_xpb_out[80][505],u_xpb_out[81][505],u_xpb_out[82][505],u_xpb_out[83][505],u_xpb_out[84][505],u_xpb_out[85][505],u_xpb_out[86][505],u_xpb_out[87][505],u_xpb_out[88][505],u_xpb_out[89][505],u_xpb_out[90][505],u_xpb_out[91][505],u_xpb_out[92][505],u_xpb_out[93][505],u_xpb_out[94][505],u_xpb_out[95][505],u_xpb_out[96][505],u_xpb_out[97][505],u_xpb_out[98][505],u_xpb_out[99][505],u_xpb_out[100][505],u_xpb_out[101][505],u_xpb_out[102][505],u_xpb_out[103][505],u_xpb_out[104][505],u_xpb_out[105][505]};

assign col_out_506 = {u_xpb_out[0][506],u_xpb_out[1][506],u_xpb_out[2][506],u_xpb_out[3][506],u_xpb_out[4][506],u_xpb_out[5][506],u_xpb_out[6][506],u_xpb_out[7][506],u_xpb_out[8][506],u_xpb_out[9][506],u_xpb_out[10][506],u_xpb_out[11][506],u_xpb_out[12][506],u_xpb_out[13][506],u_xpb_out[14][506],u_xpb_out[15][506],u_xpb_out[16][506],u_xpb_out[17][506],u_xpb_out[18][506],u_xpb_out[19][506],u_xpb_out[20][506],u_xpb_out[21][506],u_xpb_out[22][506],u_xpb_out[23][506],u_xpb_out[24][506],u_xpb_out[25][506],u_xpb_out[26][506],u_xpb_out[27][506],u_xpb_out[28][506],u_xpb_out[29][506],u_xpb_out[30][506],u_xpb_out[31][506],u_xpb_out[32][506],u_xpb_out[33][506],u_xpb_out[34][506],u_xpb_out[35][506],u_xpb_out[36][506],u_xpb_out[37][506],u_xpb_out[38][506],u_xpb_out[39][506],u_xpb_out[40][506],u_xpb_out[41][506],u_xpb_out[42][506],u_xpb_out[43][506],u_xpb_out[44][506],u_xpb_out[45][506],u_xpb_out[46][506],u_xpb_out[47][506],u_xpb_out[48][506],u_xpb_out[49][506],u_xpb_out[50][506],u_xpb_out[51][506],u_xpb_out[52][506],u_xpb_out[53][506],u_xpb_out[54][506],u_xpb_out[55][506],u_xpb_out[56][506],u_xpb_out[57][506],u_xpb_out[58][506],u_xpb_out[59][506],u_xpb_out[60][506],u_xpb_out[61][506],u_xpb_out[62][506],u_xpb_out[63][506],u_xpb_out[64][506],u_xpb_out[65][506],u_xpb_out[66][506],u_xpb_out[67][506],u_xpb_out[68][506],u_xpb_out[69][506],u_xpb_out[70][506],u_xpb_out[71][506],u_xpb_out[72][506],u_xpb_out[73][506],u_xpb_out[74][506],u_xpb_out[75][506],u_xpb_out[76][506],u_xpb_out[77][506],u_xpb_out[78][506],u_xpb_out[79][506],u_xpb_out[80][506],u_xpb_out[81][506],u_xpb_out[82][506],u_xpb_out[83][506],u_xpb_out[84][506],u_xpb_out[85][506],u_xpb_out[86][506],u_xpb_out[87][506],u_xpb_out[88][506],u_xpb_out[89][506],u_xpb_out[90][506],u_xpb_out[91][506],u_xpb_out[92][506],u_xpb_out[93][506],u_xpb_out[94][506],u_xpb_out[95][506],u_xpb_out[96][506],u_xpb_out[97][506],u_xpb_out[98][506],u_xpb_out[99][506],u_xpb_out[100][506],u_xpb_out[101][506],u_xpb_out[102][506],u_xpb_out[103][506],u_xpb_out[104][506],u_xpb_out[105][506]};

assign col_out_507 = {u_xpb_out[0][507],u_xpb_out[1][507],u_xpb_out[2][507],u_xpb_out[3][507],u_xpb_out[4][507],u_xpb_out[5][507],u_xpb_out[6][507],u_xpb_out[7][507],u_xpb_out[8][507],u_xpb_out[9][507],u_xpb_out[10][507],u_xpb_out[11][507],u_xpb_out[12][507],u_xpb_out[13][507],u_xpb_out[14][507],u_xpb_out[15][507],u_xpb_out[16][507],u_xpb_out[17][507],u_xpb_out[18][507],u_xpb_out[19][507],u_xpb_out[20][507],u_xpb_out[21][507],u_xpb_out[22][507],u_xpb_out[23][507],u_xpb_out[24][507],u_xpb_out[25][507],u_xpb_out[26][507],u_xpb_out[27][507],u_xpb_out[28][507],u_xpb_out[29][507],u_xpb_out[30][507],u_xpb_out[31][507],u_xpb_out[32][507],u_xpb_out[33][507],u_xpb_out[34][507],u_xpb_out[35][507],u_xpb_out[36][507],u_xpb_out[37][507],u_xpb_out[38][507],u_xpb_out[39][507],u_xpb_out[40][507],u_xpb_out[41][507],u_xpb_out[42][507],u_xpb_out[43][507],u_xpb_out[44][507],u_xpb_out[45][507],u_xpb_out[46][507],u_xpb_out[47][507],u_xpb_out[48][507],u_xpb_out[49][507],u_xpb_out[50][507],u_xpb_out[51][507],u_xpb_out[52][507],u_xpb_out[53][507],u_xpb_out[54][507],u_xpb_out[55][507],u_xpb_out[56][507],u_xpb_out[57][507],u_xpb_out[58][507],u_xpb_out[59][507],u_xpb_out[60][507],u_xpb_out[61][507],u_xpb_out[62][507],u_xpb_out[63][507],u_xpb_out[64][507],u_xpb_out[65][507],u_xpb_out[66][507],u_xpb_out[67][507],u_xpb_out[68][507],u_xpb_out[69][507],u_xpb_out[70][507],u_xpb_out[71][507],u_xpb_out[72][507],u_xpb_out[73][507],u_xpb_out[74][507],u_xpb_out[75][507],u_xpb_out[76][507],u_xpb_out[77][507],u_xpb_out[78][507],u_xpb_out[79][507],u_xpb_out[80][507],u_xpb_out[81][507],u_xpb_out[82][507],u_xpb_out[83][507],u_xpb_out[84][507],u_xpb_out[85][507],u_xpb_out[86][507],u_xpb_out[87][507],u_xpb_out[88][507],u_xpb_out[89][507],u_xpb_out[90][507],u_xpb_out[91][507],u_xpb_out[92][507],u_xpb_out[93][507],u_xpb_out[94][507],u_xpb_out[95][507],u_xpb_out[96][507],u_xpb_out[97][507],u_xpb_out[98][507],u_xpb_out[99][507],u_xpb_out[100][507],u_xpb_out[101][507],u_xpb_out[102][507],u_xpb_out[103][507],u_xpb_out[104][507],u_xpb_out[105][507]};

assign col_out_508 = {u_xpb_out[0][508],u_xpb_out[1][508],u_xpb_out[2][508],u_xpb_out[3][508],u_xpb_out[4][508],u_xpb_out[5][508],u_xpb_out[6][508],u_xpb_out[7][508],u_xpb_out[8][508],u_xpb_out[9][508],u_xpb_out[10][508],u_xpb_out[11][508],u_xpb_out[12][508],u_xpb_out[13][508],u_xpb_out[14][508],u_xpb_out[15][508],u_xpb_out[16][508],u_xpb_out[17][508],u_xpb_out[18][508],u_xpb_out[19][508],u_xpb_out[20][508],u_xpb_out[21][508],u_xpb_out[22][508],u_xpb_out[23][508],u_xpb_out[24][508],u_xpb_out[25][508],u_xpb_out[26][508],u_xpb_out[27][508],u_xpb_out[28][508],u_xpb_out[29][508],u_xpb_out[30][508],u_xpb_out[31][508],u_xpb_out[32][508],u_xpb_out[33][508],u_xpb_out[34][508],u_xpb_out[35][508],u_xpb_out[36][508],u_xpb_out[37][508],u_xpb_out[38][508],u_xpb_out[39][508],u_xpb_out[40][508],u_xpb_out[41][508],u_xpb_out[42][508],u_xpb_out[43][508],u_xpb_out[44][508],u_xpb_out[45][508],u_xpb_out[46][508],u_xpb_out[47][508],u_xpb_out[48][508],u_xpb_out[49][508],u_xpb_out[50][508],u_xpb_out[51][508],u_xpb_out[52][508],u_xpb_out[53][508],u_xpb_out[54][508],u_xpb_out[55][508],u_xpb_out[56][508],u_xpb_out[57][508],u_xpb_out[58][508],u_xpb_out[59][508],u_xpb_out[60][508],u_xpb_out[61][508],u_xpb_out[62][508],u_xpb_out[63][508],u_xpb_out[64][508],u_xpb_out[65][508],u_xpb_out[66][508],u_xpb_out[67][508],u_xpb_out[68][508],u_xpb_out[69][508],u_xpb_out[70][508],u_xpb_out[71][508],u_xpb_out[72][508],u_xpb_out[73][508],u_xpb_out[74][508],u_xpb_out[75][508],u_xpb_out[76][508],u_xpb_out[77][508],u_xpb_out[78][508],u_xpb_out[79][508],u_xpb_out[80][508],u_xpb_out[81][508],u_xpb_out[82][508],u_xpb_out[83][508],u_xpb_out[84][508],u_xpb_out[85][508],u_xpb_out[86][508],u_xpb_out[87][508],u_xpb_out[88][508],u_xpb_out[89][508],u_xpb_out[90][508],u_xpb_out[91][508],u_xpb_out[92][508],u_xpb_out[93][508],u_xpb_out[94][508],u_xpb_out[95][508],u_xpb_out[96][508],u_xpb_out[97][508],u_xpb_out[98][508],u_xpb_out[99][508],u_xpb_out[100][508],u_xpb_out[101][508],u_xpb_out[102][508],u_xpb_out[103][508],u_xpb_out[104][508],u_xpb_out[105][508]};

assign col_out_509 = {u_xpb_out[0][509],u_xpb_out[1][509],u_xpb_out[2][509],u_xpb_out[3][509],u_xpb_out[4][509],u_xpb_out[5][509],u_xpb_out[6][509],u_xpb_out[7][509],u_xpb_out[8][509],u_xpb_out[9][509],u_xpb_out[10][509],u_xpb_out[11][509],u_xpb_out[12][509],u_xpb_out[13][509],u_xpb_out[14][509],u_xpb_out[15][509],u_xpb_out[16][509],u_xpb_out[17][509],u_xpb_out[18][509],u_xpb_out[19][509],u_xpb_out[20][509],u_xpb_out[21][509],u_xpb_out[22][509],u_xpb_out[23][509],u_xpb_out[24][509],u_xpb_out[25][509],u_xpb_out[26][509],u_xpb_out[27][509],u_xpb_out[28][509],u_xpb_out[29][509],u_xpb_out[30][509],u_xpb_out[31][509],u_xpb_out[32][509],u_xpb_out[33][509],u_xpb_out[34][509],u_xpb_out[35][509],u_xpb_out[36][509],u_xpb_out[37][509],u_xpb_out[38][509],u_xpb_out[39][509],u_xpb_out[40][509],u_xpb_out[41][509],u_xpb_out[42][509],u_xpb_out[43][509],u_xpb_out[44][509],u_xpb_out[45][509],u_xpb_out[46][509],u_xpb_out[47][509],u_xpb_out[48][509],u_xpb_out[49][509],u_xpb_out[50][509],u_xpb_out[51][509],u_xpb_out[52][509],u_xpb_out[53][509],u_xpb_out[54][509],u_xpb_out[55][509],u_xpb_out[56][509],u_xpb_out[57][509],u_xpb_out[58][509],u_xpb_out[59][509],u_xpb_out[60][509],u_xpb_out[61][509],u_xpb_out[62][509],u_xpb_out[63][509],u_xpb_out[64][509],u_xpb_out[65][509],u_xpb_out[66][509],u_xpb_out[67][509],u_xpb_out[68][509],u_xpb_out[69][509],u_xpb_out[70][509],u_xpb_out[71][509],u_xpb_out[72][509],u_xpb_out[73][509],u_xpb_out[74][509],u_xpb_out[75][509],u_xpb_out[76][509],u_xpb_out[77][509],u_xpb_out[78][509],u_xpb_out[79][509],u_xpb_out[80][509],u_xpb_out[81][509],u_xpb_out[82][509],u_xpb_out[83][509],u_xpb_out[84][509],u_xpb_out[85][509],u_xpb_out[86][509],u_xpb_out[87][509],u_xpb_out[88][509],u_xpb_out[89][509],u_xpb_out[90][509],u_xpb_out[91][509],u_xpb_out[92][509],u_xpb_out[93][509],u_xpb_out[94][509],u_xpb_out[95][509],u_xpb_out[96][509],u_xpb_out[97][509],u_xpb_out[98][509],u_xpb_out[99][509],u_xpb_out[100][509],u_xpb_out[101][509],u_xpb_out[102][509],u_xpb_out[103][509],u_xpb_out[104][509],u_xpb_out[105][509]};

assign col_out_510 = {u_xpb_out[0][510],u_xpb_out[1][510],u_xpb_out[2][510],u_xpb_out[3][510],u_xpb_out[4][510],u_xpb_out[5][510],u_xpb_out[6][510],u_xpb_out[7][510],u_xpb_out[8][510],u_xpb_out[9][510],u_xpb_out[10][510],u_xpb_out[11][510],u_xpb_out[12][510],u_xpb_out[13][510],u_xpb_out[14][510],u_xpb_out[15][510],u_xpb_out[16][510],u_xpb_out[17][510],u_xpb_out[18][510],u_xpb_out[19][510],u_xpb_out[20][510],u_xpb_out[21][510],u_xpb_out[22][510],u_xpb_out[23][510],u_xpb_out[24][510],u_xpb_out[25][510],u_xpb_out[26][510],u_xpb_out[27][510],u_xpb_out[28][510],u_xpb_out[29][510],u_xpb_out[30][510],u_xpb_out[31][510],u_xpb_out[32][510],u_xpb_out[33][510],u_xpb_out[34][510],u_xpb_out[35][510],u_xpb_out[36][510],u_xpb_out[37][510],u_xpb_out[38][510],u_xpb_out[39][510],u_xpb_out[40][510],u_xpb_out[41][510],u_xpb_out[42][510],u_xpb_out[43][510],u_xpb_out[44][510],u_xpb_out[45][510],u_xpb_out[46][510],u_xpb_out[47][510],u_xpb_out[48][510],u_xpb_out[49][510],u_xpb_out[50][510],u_xpb_out[51][510],u_xpb_out[52][510],u_xpb_out[53][510],u_xpb_out[54][510],u_xpb_out[55][510],u_xpb_out[56][510],u_xpb_out[57][510],u_xpb_out[58][510],u_xpb_out[59][510],u_xpb_out[60][510],u_xpb_out[61][510],u_xpb_out[62][510],u_xpb_out[63][510],u_xpb_out[64][510],u_xpb_out[65][510],u_xpb_out[66][510],u_xpb_out[67][510],u_xpb_out[68][510],u_xpb_out[69][510],u_xpb_out[70][510],u_xpb_out[71][510],u_xpb_out[72][510],u_xpb_out[73][510],u_xpb_out[74][510],u_xpb_out[75][510],u_xpb_out[76][510],u_xpb_out[77][510],u_xpb_out[78][510],u_xpb_out[79][510],u_xpb_out[80][510],u_xpb_out[81][510],u_xpb_out[82][510],u_xpb_out[83][510],u_xpb_out[84][510],u_xpb_out[85][510],u_xpb_out[86][510],u_xpb_out[87][510],u_xpb_out[88][510],u_xpb_out[89][510],u_xpb_out[90][510],u_xpb_out[91][510],u_xpb_out[92][510],u_xpb_out[93][510],u_xpb_out[94][510],u_xpb_out[95][510],u_xpb_out[96][510],u_xpb_out[97][510],u_xpb_out[98][510],u_xpb_out[99][510],u_xpb_out[100][510],u_xpb_out[101][510],u_xpb_out[102][510],u_xpb_out[103][510],u_xpb_out[104][510],u_xpb_out[105][510]};

assign col_out_511 = {u_xpb_out[0][511],u_xpb_out[1][511],u_xpb_out[2][511],u_xpb_out[3][511],u_xpb_out[4][511],u_xpb_out[5][511],u_xpb_out[6][511],u_xpb_out[7][511],u_xpb_out[8][511],u_xpb_out[9][511],u_xpb_out[10][511],u_xpb_out[11][511],u_xpb_out[12][511],u_xpb_out[13][511],u_xpb_out[14][511],u_xpb_out[15][511],u_xpb_out[16][511],u_xpb_out[17][511],u_xpb_out[18][511],u_xpb_out[19][511],u_xpb_out[20][511],u_xpb_out[21][511],u_xpb_out[22][511],u_xpb_out[23][511],u_xpb_out[24][511],u_xpb_out[25][511],u_xpb_out[26][511],u_xpb_out[27][511],u_xpb_out[28][511],u_xpb_out[29][511],u_xpb_out[30][511],u_xpb_out[31][511],u_xpb_out[32][511],u_xpb_out[33][511],u_xpb_out[34][511],u_xpb_out[35][511],u_xpb_out[36][511],u_xpb_out[37][511],u_xpb_out[38][511],u_xpb_out[39][511],u_xpb_out[40][511],u_xpb_out[41][511],u_xpb_out[42][511],u_xpb_out[43][511],u_xpb_out[44][511],u_xpb_out[45][511],u_xpb_out[46][511],u_xpb_out[47][511],u_xpb_out[48][511],u_xpb_out[49][511],u_xpb_out[50][511],u_xpb_out[51][511],u_xpb_out[52][511],u_xpb_out[53][511],u_xpb_out[54][511],u_xpb_out[55][511],u_xpb_out[56][511],u_xpb_out[57][511],u_xpb_out[58][511],u_xpb_out[59][511],u_xpb_out[60][511],u_xpb_out[61][511],u_xpb_out[62][511],u_xpb_out[63][511],u_xpb_out[64][511],u_xpb_out[65][511],u_xpb_out[66][511],u_xpb_out[67][511],u_xpb_out[68][511],u_xpb_out[69][511],u_xpb_out[70][511],u_xpb_out[71][511],u_xpb_out[72][511],u_xpb_out[73][511],u_xpb_out[74][511],u_xpb_out[75][511],u_xpb_out[76][511],u_xpb_out[77][511],u_xpb_out[78][511],u_xpb_out[79][511],u_xpb_out[80][511],u_xpb_out[81][511],u_xpb_out[82][511],u_xpb_out[83][511],u_xpb_out[84][511],u_xpb_out[85][511],u_xpb_out[86][511],u_xpb_out[87][511],u_xpb_out[88][511],u_xpb_out[89][511],u_xpb_out[90][511],u_xpb_out[91][511],u_xpb_out[92][511],u_xpb_out[93][511],u_xpb_out[94][511],u_xpb_out[95][511],u_xpb_out[96][511],u_xpb_out[97][511],u_xpb_out[98][511],u_xpb_out[99][511],u_xpb_out[100][511],u_xpb_out[101][511],u_xpb_out[102][511],u_xpb_out[103][511],u_xpb_out[104][511],u_xpb_out[105][511]};

assign col_out_512 = {u_xpb_out[0][512],u_xpb_out[1][512],u_xpb_out[2][512],u_xpb_out[3][512],u_xpb_out[4][512],u_xpb_out[5][512],u_xpb_out[6][512],u_xpb_out[7][512],u_xpb_out[8][512],u_xpb_out[9][512],u_xpb_out[10][512],u_xpb_out[11][512],u_xpb_out[12][512],u_xpb_out[13][512],u_xpb_out[14][512],u_xpb_out[15][512],u_xpb_out[16][512],u_xpb_out[17][512],u_xpb_out[18][512],u_xpb_out[19][512],u_xpb_out[20][512],u_xpb_out[21][512],u_xpb_out[22][512],u_xpb_out[23][512],u_xpb_out[24][512],u_xpb_out[25][512],u_xpb_out[26][512],u_xpb_out[27][512],u_xpb_out[28][512],u_xpb_out[29][512],u_xpb_out[30][512],u_xpb_out[31][512],u_xpb_out[32][512],u_xpb_out[33][512],u_xpb_out[34][512],u_xpb_out[35][512],u_xpb_out[36][512],u_xpb_out[37][512],u_xpb_out[38][512],u_xpb_out[39][512],u_xpb_out[40][512],u_xpb_out[41][512],u_xpb_out[42][512],u_xpb_out[43][512],u_xpb_out[44][512],u_xpb_out[45][512],u_xpb_out[46][512],u_xpb_out[47][512],u_xpb_out[48][512],u_xpb_out[49][512],u_xpb_out[50][512],u_xpb_out[51][512],u_xpb_out[52][512],u_xpb_out[53][512],u_xpb_out[54][512],u_xpb_out[55][512],u_xpb_out[56][512],u_xpb_out[57][512],u_xpb_out[58][512],u_xpb_out[59][512],u_xpb_out[60][512],u_xpb_out[61][512],u_xpb_out[62][512],u_xpb_out[63][512],u_xpb_out[64][512],u_xpb_out[65][512],u_xpb_out[66][512],u_xpb_out[67][512],u_xpb_out[68][512],u_xpb_out[69][512],u_xpb_out[70][512],u_xpb_out[71][512],u_xpb_out[72][512],u_xpb_out[73][512],u_xpb_out[74][512],u_xpb_out[75][512],u_xpb_out[76][512],u_xpb_out[77][512],u_xpb_out[78][512],u_xpb_out[79][512],u_xpb_out[80][512],u_xpb_out[81][512],u_xpb_out[82][512],u_xpb_out[83][512],u_xpb_out[84][512],u_xpb_out[85][512],u_xpb_out[86][512],u_xpb_out[87][512],u_xpb_out[88][512],u_xpb_out[89][512],u_xpb_out[90][512],u_xpb_out[91][512],u_xpb_out[92][512],u_xpb_out[93][512],u_xpb_out[94][512],u_xpb_out[95][512],u_xpb_out[96][512],u_xpb_out[97][512],u_xpb_out[98][512],u_xpb_out[99][512],u_xpb_out[100][512],u_xpb_out[101][512],u_xpb_out[102][512],u_xpb_out[103][512],u_xpb_out[104][512],u_xpb_out[105][512]};

assign col_out_513 = {u_xpb_out[0][513],u_xpb_out[1][513],u_xpb_out[2][513],u_xpb_out[3][513],u_xpb_out[4][513],u_xpb_out[5][513],u_xpb_out[6][513],u_xpb_out[7][513],u_xpb_out[8][513],u_xpb_out[9][513],u_xpb_out[10][513],u_xpb_out[11][513],u_xpb_out[12][513],u_xpb_out[13][513],u_xpb_out[14][513],u_xpb_out[15][513],u_xpb_out[16][513],u_xpb_out[17][513],u_xpb_out[18][513],u_xpb_out[19][513],u_xpb_out[20][513],u_xpb_out[21][513],u_xpb_out[22][513],u_xpb_out[23][513],u_xpb_out[24][513],u_xpb_out[25][513],u_xpb_out[26][513],u_xpb_out[27][513],u_xpb_out[28][513],u_xpb_out[29][513],u_xpb_out[30][513],u_xpb_out[31][513],u_xpb_out[32][513],u_xpb_out[33][513],u_xpb_out[34][513],u_xpb_out[35][513],u_xpb_out[36][513],u_xpb_out[37][513],u_xpb_out[38][513],u_xpb_out[39][513],u_xpb_out[40][513],u_xpb_out[41][513],u_xpb_out[42][513],u_xpb_out[43][513],u_xpb_out[44][513],u_xpb_out[45][513],u_xpb_out[46][513],u_xpb_out[47][513],u_xpb_out[48][513],u_xpb_out[49][513],u_xpb_out[50][513],u_xpb_out[51][513],u_xpb_out[52][513],u_xpb_out[53][513],u_xpb_out[54][513],u_xpb_out[55][513],u_xpb_out[56][513],u_xpb_out[57][513],u_xpb_out[58][513],u_xpb_out[59][513],u_xpb_out[60][513],u_xpb_out[61][513],u_xpb_out[62][513],u_xpb_out[63][513],u_xpb_out[64][513],u_xpb_out[65][513],u_xpb_out[66][513],u_xpb_out[67][513],u_xpb_out[68][513],u_xpb_out[69][513],u_xpb_out[70][513],u_xpb_out[71][513],u_xpb_out[72][513],u_xpb_out[73][513],u_xpb_out[74][513],u_xpb_out[75][513],u_xpb_out[76][513],u_xpb_out[77][513],u_xpb_out[78][513],u_xpb_out[79][513],u_xpb_out[80][513],u_xpb_out[81][513],u_xpb_out[82][513],u_xpb_out[83][513],u_xpb_out[84][513],u_xpb_out[85][513],u_xpb_out[86][513],u_xpb_out[87][513],u_xpb_out[88][513],u_xpb_out[89][513],u_xpb_out[90][513],u_xpb_out[91][513],u_xpb_out[92][513],u_xpb_out[93][513],u_xpb_out[94][513],u_xpb_out[95][513],u_xpb_out[96][513],u_xpb_out[97][513],u_xpb_out[98][513],u_xpb_out[99][513],u_xpb_out[100][513],u_xpb_out[101][513],u_xpb_out[102][513],u_xpb_out[103][513],u_xpb_out[104][513],u_xpb_out[105][513]};

assign col_out_514 = {u_xpb_out[0][514],u_xpb_out[1][514],u_xpb_out[2][514],u_xpb_out[3][514],u_xpb_out[4][514],u_xpb_out[5][514],u_xpb_out[6][514],u_xpb_out[7][514],u_xpb_out[8][514],u_xpb_out[9][514],u_xpb_out[10][514],u_xpb_out[11][514],u_xpb_out[12][514],u_xpb_out[13][514],u_xpb_out[14][514],u_xpb_out[15][514],u_xpb_out[16][514],u_xpb_out[17][514],u_xpb_out[18][514],u_xpb_out[19][514],u_xpb_out[20][514],u_xpb_out[21][514],u_xpb_out[22][514],u_xpb_out[23][514],u_xpb_out[24][514],u_xpb_out[25][514],u_xpb_out[26][514],u_xpb_out[27][514],u_xpb_out[28][514],u_xpb_out[29][514],u_xpb_out[30][514],u_xpb_out[31][514],u_xpb_out[32][514],u_xpb_out[33][514],u_xpb_out[34][514],u_xpb_out[35][514],u_xpb_out[36][514],u_xpb_out[37][514],u_xpb_out[38][514],u_xpb_out[39][514],u_xpb_out[40][514],u_xpb_out[41][514],u_xpb_out[42][514],u_xpb_out[43][514],u_xpb_out[44][514],u_xpb_out[45][514],u_xpb_out[46][514],u_xpb_out[47][514],u_xpb_out[48][514],u_xpb_out[49][514],u_xpb_out[50][514],u_xpb_out[51][514],u_xpb_out[52][514],u_xpb_out[53][514],u_xpb_out[54][514],u_xpb_out[55][514],u_xpb_out[56][514],u_xpb_out[57][514],u_xpb_out[58][514],u_xpb_out[59][514],u_xpb_out[60][514],u_xpb_out[61][514],u_xpb_out[62][514],u_xpb_out[63][514],u_xpb_out[64][514],u_xpb_out[65][514],u_xpb_out[66][514],u_xpb_out[67][514],u_xpb_out[68][514],u_xpb_out[69][514],u_xpb_out[70][514],u_xpb_out[71][514],u_xpb_out[72][514],u_xpb_out[73][514],u_xpb_out[74][514],u_xpb_out[75][514],u_xpb_out[76][514],u_xpb_out[77][514],u_xpb_out[78][514],u_xpb_out[79][514],u_xpb_out[80][514],u_xpb_out[81][514],u_xpb_out[82][514],u_xpb_out[83][514],u_xpb_out[84][514],u_xpb_out[85][514],u_xpb_out[86][514],u_xpb_out[87][514],u_xpb_out[88][514],u_xpb_out[89][514],u_xpb_out[90][514],u_xpb_out[91][514],u_xpb_out[92][514],u_xpb_out[93][514],u_xpb_out[94][514],u_xpb_out[95][514],u_xpb_out[96][514],u_xpb_out[97][514],u_xpb_out[98][514],u_xpb_out[99][514],u_xpb_out[100][514],u_xpb_out[101][514],u_xpb_out[102][514],u_xpb_out[103][514],u_xpb_out[104][514],u_xpb_out[105][514]};

assign col_out_515 = {u_xpb_out[0][515],u_xpb_out[1][515],u_xpb_out[2][515],u_xpb_out[3][515],u_xpb_out[4][515],u_xpb_out[5][515],u_xpb_out[6][515],u_xpb_out[7][515],u_xpb_out[8][515],u_xpb_out[9][515],u_xpb_out[10][515],u_xpb_out[11][515],u_xpb_out[12][515],u_xpb_out[13][515],u_xpb_out[14][515],u_xpb_out[15][515],u_xpb_out[16][515],u_xpb_out[17][515],u_xpb_out[18][515],u_xpb_out[19][515],u_xpb_out[20][515],u_xpb_out[21][515],u_xpb_out[22][515],u_xpb_out[23][515],u_xpb_out[24][515],u_xpb_out[25][515],u_xpb_out[26][515],u_xpb_out[27][515],u_xpb_out[28][515],u_xpb_out[29][515],u_xpb_out[30][515],u_xpb_out[31][515],u_xpb_out[32][515],u_xpb_out[33][515],u_xpb_out[34][515],u_xpb_out[35][515],u_xpb_out[36][515],u_xpb_out[37][515],u_xpb_out[38][515],u_xpb_out[39][515],u_xpb_out[40][515],u_xpb_out[41][515],u_xpb_out[42][515],u_xpb_out[43][515],u_xpb_out[44][515],u_xpb_out[45][515],u_xpb_out[46][515],u_xpb_out[47][515],u_xpb_out[48][515],u_xpb_out[49][515],u_xpb_out[50][515],u_xpb_out[51][515],u_xpb_out[52][515],u_xpb_out[53][515],u_xpb_out[54][515],u_xpb_out[55][515],u_xpb_out[56][515],u_xpb_out[57][515],u_xpb_out[58][515],u_xpb_out[59][515],u_xpb_out[60][515],u_xpb_out[61][515],u_xpb_out[62][515],u_xpb_out[63][515],u_xpb_out[64][515],u_xpb_out[65][515],u_xpb_out[66][515],u_xpb_out[67][515],u_xpb_out[68][515],u_xpb_out[69][515],u_xpb_out[70][515],u_xpb_out[71][515],u_xpb_out[72][515],u_xpb_out[73][515],u_xpb_out[74][515],u_xpb_out[75][515],u_xpb_out[76][515],u_xpb_out[77][515],u_xpb_out[78][515],u_xpb_out[79][515],u_xpb_out[80][515],u_xpb_out[81][515],u_xpb_out[82][515],u_xpb_out[83][515],u_xpb_out[84][515],u_xpb_out[85][515],u_xpb_out[86][515],u_xpb_out[87][515],u_xpb_out[88][515],u_xpb_out[89][515],u_xpb_out[90][515],u_xpb_out[91][515],u_xpb_out[92][515],u_xpb_out[93][515],u_xpb_out[94][515],u_xpb_out[95][515],u_xpb_out[96][515],u_xpb_out[97][515],u_xpb_out[98][515],u_xpb_out[99][515],u_xpb_out[100][515],u_xpb_out[101][515],u_xpb_out[102][515],u_xpb_out[103][515],u_xpb_out[104][515],u_xpb_out[105][515]};

assign col_out_516 = {u_xpb_out[0][516],u_xpb_out[1][516],u_xpb_out[2][516],u_xpb_out[3][516],u_xpb_out[4][516],u_xpb_out[5][516],u_xpb_out[6][516],u_xpb_out[7][516],u_xpb_out[8][516],u_xpb_out[9][516],u_xpb_out[10][516],u_xpb_out[11][516],u_xpb_out[12][516],u_xpb_out[13][516],u_xpb_out[14][516],u_xpb_out[15][516],u_xpb_out[16][516],u_xpb_out[17][516],u_xpb_out[18][516],u_xpb_out[19][516],u_xpb_out[20][516],u_xpb_out[21][516],u_xpb_out[22][516],u_xpb_out[23][516],u_xpb_out[24][516],u_xpb_out[25][516],u_xpb_out[26][516],u_xpb_out[27][516],u_xpb_out[28][516],u_xpb_out[29][516],u_xpb_out[30][516],u_xpb_out[31][516],u_xpb_out[32][516],u_xpb_out[33][516],u_xpb_out[34][516],u_xpb_out[35][516],u_xpb_out[36][516],u_xpb_out[37][516],u_xpb_out[38][516],u_xpb_out[39][516],u_xpb_out[40][516],u_xpb_out[41][516],u_xpb_out[42][516],u_xpb_out[43][516],u_xpb_out[44][516],u_xpb_out[45][516],u_xpb_out[46][516],u_xpb_out[47][516],u_xpb_out[48][516],u_xpb_out[49][516],u_xpb_out[50][516],u_xpb_out[51][516],u_xpb_out[52][516],u_xpb_out[53][516],u_xpb_out[54][516],u_xpb_out[55][516],u_xpb_out[56][516],u_xpb_out[57][516],u_xpb_out[58][516],u_xpb_out[59][516],u_xpb_out[60][516],u_xpb_out[61][516],u_xpb_out[62][516],u_xpb_out[63][516],u_xpb_out[64][516],u_xpb_out[65][516],u_xpb_out[66][516],u_xpb_out[67][516],u_xpb_out[68][516],u_xpb_out[69][516],u_xpb_out[70][516],u_xpb_out[71][516],u_xpb_out[72][516],u_xpb_out[73][516],u_xpb_out[74][516],u_xpb_out[75][516],u_xpb_out[76][516],u_xpb_out[77][516],u_xpb_out[78][516],u_xpb_out[79][516],u_xpb_out[80][516],u_xpb_out[81][516],u_xpb_out[82][516],u_xpb_out[83][516],u_xpb_out[84][516],u_xpb_out[85][516],u_xpb_out[86][516],u_xpb_out[87][516],u_xpb_out[88][516],u_xpb_out[89][516],u_xpb_out[90][516],u_xpb_out[91][516],u_xpb_out[92][516],u_xpb_out[93][516],u_xpb_out[94][516],u_xpb_out[95][516],u_xpb_out[96][516],u_xpb_out[97][516],u_xpb_out[98][516],u_xpb_out[99][516],u_xpb_out[100][516],u_xpb_out[101][516],u_xpb_out[102][516],u_xpb_out[103][516],u_xpb_out[104][516],u_xpb_out[105][516]};

assign col_out_517 = {u_xpb_out[0][517],u_xpb_out[1][517],u_xpb_out[2][517],u_xpb_out[3][517],u_xpb_out[4][517],u_xpb_out[5][517],u_xpb_out[6][517],u_xpb_out[7][517],u_xpb_out[8][517],u_xpb_out[9][517],u_xpb_out[10][517],u_xpb_out[11][517],u_xpb_out[12][517],u_xpb_out[13][517],u_xpb_out[14][517],u_xpb_out[15][517],u_xpb_out[16][517],u_xpb_out[17][517],u_xpb_out[18][517],u_xpb_out[19][517],u_xpb_out[20][517],u_xpb_out[21][517],u_xpb_out[22][517],u_xpb_out[23][517],u_xpb_out[24][517],u_xpb_out[25][517],u_xpb_out[26][517],u_xpb_out[27][517],u_xpb_out[28][517],u_xpb_out[29][517],u_xpb_out[30][517],u_xpb_out[31][517],u_xpb_out[32][517],u_xpb_out[33][517],u_xpb_out[34][517],u_xpb_out[35][517],u_xpb_out[36][517],u_xpb_out[37][517],u_xpb_out[38][517],u_xpb_out[39][517],u_xpb_out[40][517],u_xpb_out[41][517],u_xpb_out[42][517],u_xpb_out[43][517],u_xpb_out[44][517],u_xpb_out[45][517],u_xpb_out[46][517],u_xpb_out[47][517],u_xpb_out[48][517],u_xpb_out[49][517],u_xpb_out[50][517],u_xpb_out[51][517],u_xpb_out[52][517],u_xpb_out[53][517],u_xpb_out[54][517],u_xpb_out[55][517],u_xpb_out[56][517],u_xpb_out[57][517],u_xpb_out[58][517],u_xpb_out[59][517],u_xpb_out[60][517],u_xpb_out[61][517],u_xpb_out[62][517],u_xpb_out[63][517],u_xpb_out[64][517],u_xpb_out[65][517],u_xpb_out[66][517],u_xpb_out[67][517],u_xpb_out[68][517],u_xpb_out[69][517],u_xpb_out[70][517],u_xpb_out[71][517],u_xpb_out[72][517],u_xpb_out[73][517],u_xpb_out[74][517],u_xpb_out[75][517],u_xpb_out[76][517],u_xpb_out[77][517],u_xpb_out[78][517],u_xpb_out[79][517],u_xpb_out[80][517],u_xpb_out[81][517],u_xpb_out[82][517],u_xpb_out[83][517],u_xpb_out[84][517],u_xpb_out[85][517],u_xpb_out[86][517],u_xpb_out[87][517],u_xpb_out[88][517],u_xpb_out[89][517],u_xpb_out[90][517],u_xpb_out[91][517],u_xpb_out[92][517],u_xpb_out[93][517],u_xpb_out[94][517],u_xpb_out[95][517],u_xpb_out[96][517],u_xpb_out[97][517],u_xpb_out[98][517],u_xpb_out[99][517],u_xpb_out[100][517],u_xpb_out[101][517],u_xpb_out[102][517],u_xpb_out[103][517],u_xpb_out[104][517],u_xpb_out[105][517]};

assign col_out_518 = {u_xpb_out[0][518],u_xpb_out[1][518],u_xpb_out[2][518],u_xpb_out[3][518],u_xpb_out[4][518],u_xpb_out[5][518],u_xpb_out[6][518],u_xpb_out[7][518],u_xpb_out[8][518],u_xpb_out[9][518],u_xpb_out[10][518],u_xpb_out[11][518],u_xpb_out[12][518],u_xpb_out[13][518],u_xpb_out[14][518],u_xpb_out[15][518],u_xpb_out[16][518],u_xpb_out[17][518],u_xpb_out[18][518],u_xpb_out[19][518],u_xpb_out[20][518],u_xpb_out[21][518],u_xpb_out[22][518],u_xpb_out[23][518],u_xpb_out[24][518],u_xpb_out[25][518],u_xpb_out[26][518],u_xpb_out[27][518],u_xpb_out[28][518],u_xpb_out[29][518],u_xpb_out[30][518],u_xpb_out[31][518],u_xpb_out[32][518],u_xpb_out[33][518],u_xpb_out[34][518],u_xpb_out[35][518],u_xpb_out[36][518],u_xpb_out[37][518],u_xpb_out[38][518],u_xpb_out[39][518],u_xpb_out[40][518],u_xpb_out[41][518],u_xpb_out[42][518],u_xpb_out[43][518],u_xpb_out[44][518],u_xpb_out[45][518],u_xpb_out[46][518],u_xpb_out[47][518],u_xpb_out[48][518],u_xpb_out[49][518],u_xpb_out[50][518],u_xpb_out[51][518],u_xpb_out[52][518],u_xpb_out[53][518],u_xpb_out[54][518],u_xpb_out[55][518],u_xpb_out[56][518],u_xpb_out[57][518],u_xpb_out[58][518],u_xpb_out[59][518],u_xpb_out[60][518],u_xpb_out[61][518],u_xpb_out[62][518],u_xpb_out[63][518],u_xpb_out[64][518],u_xpb_out[65][518],u_xpb_out[66][518],u_xpb_out[67][518],u_xpb_out[68][518],u_xpb_out[69][518],u_xpb_out[70][518],u_xpb_out[71][518],u_xpb_out[72][518],u_xpb_out[73][518],u_xpb_out[74][518],u_xpb_out[75][518],u_xpb_out[76][518],u_xpb_out[77][518],u_xpb_out[78][518],u_xpb_out[79][518],u_xpb_out[80][518],u_xpb_out[81][518],u_xpb_out[82][518],u_xpb_out[83][518],u_xpb_out[84][518],u_xpb_out[85][518],u_xpb_out[86][518],u_xpb_out[87][518],u_xpb_out[88][518],u_xpb_out[89][518],u_xpb_out[90][518],u_xpb_out[91][518],u_xpb_out[92][518],u_xpb_out[93][518],u_xpb_out[94][518],u_xpb_out[95][518],u_xpb_out[96][518],u_xpb_out[97][518],u_xpb_out[98][518],u_xpb_out[99][518],u_xpb_out[100][518],u_xpb_out[101][518],u_xpb_out[102][518],u_xpb_out[103][518],u_xpb_out[104][518],u_xpb_out[105][518]};

assign col_out_519 = {u_xpb_out[0][519],u_xpb_out[1][519],u_xpb_out[2][519],u_xpb_out[3][519],u_xpb_out[4][519],u_xpb_out[5][519],u_xpb_out[6][519],u_xpb_out[7][519],u_xpb_out[8][519],u_xpb_out[9][519],u_xpb_out[10][519],u_xpb_out[11][519],u_xpb_out[12][519],u_xpb_out[13][519],u_xpb_out[14][519],u_xpb_out[15][519],u_xpb_out[16][519],u_xpb_out[17][519],u_xpb_out[18][519],u_xpb_out[19][519],u_xpb_out[20][519],u_xpb_out[21][519],u_xpb_out[22][519],u_xpb_out[23][519],u_xpb_out[24][519],u_xpb_out[25][519],u_xpb_out[26][519],u_xpb_out[27][519],u_xpb_out[28][519],u_xpb_out[29][519],u_xpb_out[30][519],u_xpb_out[31][519],u_xpb_out[32][519],u_xpb_out[33][519],u_xpb_out[34][519],u_xpb_out[35][519],u_xpb_out[36][519],u_xpb_out[37][519],u_xpb_out[38][519],u_xpb_out[39][519],u_xpb_out[40][519],u_xpb_out[41][519],u_xpb_out[42][519],u_xpb_out[43][519],u_xpb_out[44][519],u_xpb_out[45][519],u_xpb_out[46][519],u_xpb_out[47][519],u_xpb_out[48][519],u_xpb_out[49][519],u_xpb_out[50][519],u_xpb_out[51][519],u_xpb_out[52][519],u_xpb_out[53][519],u_xpb_out[54][519],u_xpb_out[55][519],u_xpb_out[56][519],u_xpb_out[57][519],u_xpb_out[58][519],u_xpb_out[59][519],u_xpb_out[60][519],u_xpb_out[61][519],u_xpb_out[62][519],u_xpb_out[63][519],u_xpb_out[64][519],u_xpb_out[65][519],u_xpb_out[66][519],u_xpb_out[67][519],u_xpb_out[68][519],u_xpb_out[69][519],u_xpb_out[70][519],u_xpb_out[71][519],u_xpb_out[72][519],u_xpb_out[73][519],u_xpb_out[74][519],u_xpb_out[75][519],u_xpb_out[76][519],u_xpb_out[77][519],u_xpb_out[78][519],u_xpb_out[79][519],u_xpb_out[80][519],u_xpb_out[81][519],u_xpb_out[82][519],u_xpb_out[83][519],u_xpb_out[84][519],u_xpb_out[85][519],u_xpb_out[86][519],u_xpb_out[87][519],u_xpb_out[88][519],u_xpb_out[89][519],u_xpb_out[90][519],u_xpb_out[91][519],u_xpb_out[92][519],u_xpb_out[93][519],u_xpb_out[94][519],u_xpb_out[95][519],u_xpb_out[96][519],u_xpb_out[97][519],u_xpb_out[98][519],u_xpb_out[99][519],u_xpb_out[100][519],u_xpb_out[101][519],u_xpb_out[102][519],u_xpb_out[103][519],u_xpb_out[104][519],u_xpb_out[105][519]};

assign col_out_520 = {u_xpb_out[0][520],u_xpb_out[1][520],u_xpb_out[2][520],u_xpb_out[3][520],u_xpb_out[4][520],u_xpb_out[5][520],u_xpb_out[6][520],u_xpb_out[7][520],u_xpb_out[8][520],u_xpb_out[9][520],u_xpb_out[10][520],u_xpb_out[11][520],u_xpb_out[12][520],u_xpb_out[13][520],u_xpb_out[14][520],u_xpb_out[15][520],u_xpb_out[16][520],u_xpb_out[17][520],u_xpb_out[18][520],u_xpb_out[19][520],u_xpb_out[20][520],u_xpb_out[21][520],u_xpb_out[22][520],u_xpb_out[23][520],u_xpb_out[24][520],u_xpb_out[25][520],u_xpb_out[26][520],u_xpb_out[27][520],u_xpb_out[28][520],u_xpb_out[29][520],u_xpb_out[30][520],u_xpb_out[31][520],u_xpb_out[32][520],u_xpb_out[33][520],u_xpb_out[34][520],u_xpb_out[35][520],u_xpb_out[36][520],u_xpb_out[37][520],u_xpb_out[38][520],u_xpb_out[39][520],u_xpb_out[40][520],u_xpb_out[41][520],u_xpb_out[42][520],u_xpb_out[43][520],u_xpb_out[44][520],u_xpb_out[45][520],u_xpb_out[46][520],u_xpb_out[47][520],u_xpb_out[48][520],u_xpb_out[49][520],u_xpb_out[50][520],u_xpb_out[51][520],u_xpb_out[52][520],u_xpb_out[53][520],u_xpb_out[54][520],u_xpb_out[55][520],u_xpb_out[56][520],u_xpb_out[57][520],u_xpb_out[58][520],u_xpb_out[59][520],u_xpb_out[60][520],u_xpb_out[61][520],u_xpb_out[62][520],u_xpb_out[63][520],u_xpb_out[64][520],u_xpb_out[65][520],u_xpb_out[66][520],u_xpb_out[67][520],u_xpb_out[68][520],u_xpb_out[69][520],u_xpb_out[70][520],u_xpb_out[71][520],u_xpb_out[72][520],u_xpb_out[73][520],u_xpb_out[74][520],u_xpb_out[75][520],u_xpb_out[76][520],u_xpb_out[77][520],u_xpb_out[78][520],u_xpb_out[79][520],u_xpb_out[80][520],u_xpb_out[81][520],u_xpb_out[82][520],u_xpb_out[83][520],u_xpb_out[84][520],u_xpb_out[85][520],u_xpb_out[86][520],u_xpb_out[87][520],u_xpb_out[88][520],u_xpb_out[89][520],u_xpb_out[90][520],u_xpb_out[91][520],u_xpb_out[92][520],u_xpb_out[93][520],u_xpb_out[94][520],u_xpb_out[95][520],u_xpb_out[96][520],u_xpb_out[97][520],u_xpb_out[98][520],u_xpb_out[99][520],u_xpb_out[100][520],u_xpb_out[101][520],u_xpb_out[102][520],u_xpb_out[103][520],u_xpb_out[104][520],u_xpb_out[105][520]};

assign col_out_521 = {u_xpb_out[0][521],u_xpb_out[1][521],u_xpb_out[2][521],u_xpb_out[3][521],u_xpb_out[4][521],u_xpb_out[5][521],u_xpb_out[6][521],u_xpb_out[7][521],u_xpb_out[8][521],u_xpb_out[9][521],u_xpb_out[10][521],u_xpb_out[11][521],u_xpb_out[12][521],u_xpb_out[13][521],u_xpb_out[14][521],u_xpb_out[15][521],u_xpb_out[16][521],u_xpb_out[17][521],u_xpb_out[18][521],u_xpb_out[19][521],u_xpb_out[20][521],u_xpb_out[21][521],u_xpb_out[22][521],u_xpb_out[23][521],u_xpb_out[24][521],u_xpb_out[25][521],u_xpb_out[26][521],u_xpb_out[27][521],u_xpb_out[28][521],u_xpb_out[29][521],u_xpb_out[30][521],u_xpb_out[31][521],u_xpb_out[32][521],u_xpb_out[33][521],u_xpb_out[34][521],u_xpb_out[35][521],u_xpb_out[36][521],u_xpb_out[37][521],u_xpb_out[38][521],u_xpb_out[39][521],u_xpb_out[40][521],u_xpb_out[41][521],u_xpb_out[42][521],u_xpb_out[43][521],u_xpb_out[44][521],u_xpb_out[45][521],u_xpb_out[46][521],u_xpb_out[47][521],u_xpb_out[48][521],u_xpb_out[49][521],u_xpb_out[50][521],u_xpb_out[51][521],u_xpb_out[52][521],u_xpb_out[53][521],u_xpb_out[54][521],u_xpb_out[55][521],u_xpb_out[56][521],u_xpb_out[57][521],u_xpb_out[58][521],u_xpb_out[59][521],u_xpb_out[60][521],u_xpb_out[61][521],u_xpb_out[62][521],u_xpb_out[63][521],u_xpb_out[64][521],u_xpb_out[65][521],u_xpb_out[66][521],u_xpb_out[67][521],u_xpb_out[68][521],u_xpb_out[69][521],u_xpb_out[70][521],u_xpb_out[71][521],u_xpb_out[72][521],u_xpb_out[73][521],u_xpb_out[74][521],u_xpb_out[75][521],u_xpb_out[76][521],u_xpb_out[77][521],u_xpb_out[78][521],u_xpb_out[79][521],u_xpb_out[80][521],u_xpb_out[81][521],u_xpb_out[82][521],u_xpb_out[83][521],u_xpb_out[84][521],u_xpb_out[85][521],u_xpb_out[86][521],u_xpb_out[87][521],u_xpb_out[88][521],u_xpb_out[89][521],u_xpb_out[90][521],u_xpb_out[91][521],u_xpb_out[92][521],u_xpb_out[93][521],u_xpb_out[94][521],u_xpb_out[95][521],u_xpb_out[96][521],u_xpb_out[97][521],u_xpb_out[98][521],u_xpb_out[99][521],u_xpb_out[100][521],u_xpb_out[101][521],u_xpb_out[102][521],u_xpb_out[103][521],u_xpb_out[104][521],u_xpb_out[105][521]};

assign col_out_522 = {u_xpb_out[0][522],u_xpb_out[1][522],u_xpb_out[2][522],u_xpb_out[3][522],u_xpb_out[4][522],u_xpb_out[5][522],u_xpb_out[6][522],u_xpb_out[7][522],u_xpb_out[8][522],u_xpb_out[9][522],u_xpb_out[10][522],u_xpb_out[11][522],u_xpb_out[12][522],u_xpb_out[13][522],u_xpb_out[14][522],u_xpb_out[15][522],u_xpb_out[16][522],u_xpb_out[17][522],u_xpb_out[18][522],u_xpb_out[19][522],u_xpb_out[20][522],u_xpb_out[21][522],u_xpb_out[22][522],u_xpb_out[23][522],u_xpb_out[24][522],u_xpb_out[25][522],u_xpb_out[26][522],u_xpb_out[27][522],u_xpb_out[28][522],u_xpb_out[29][522],u_xpb_out[30][522],u_xpb_out[31][522],u_xpb_out[32][522],u_xpb_out[33][522],u_xpb_out[34][522],u_xpb_out[35][522],u_xpb_out[36][522],u_xpb_out[37][522],u_xpb_out[38][522],u_xpb_out[39][522],u_xpb_out[40][522],u_xpb_out[41][522],u_xpb_out[42][522],u_xpb_out[43][522],u_xpb_out[44][522],u_xpb_out[45][522],u_xpb_out[46][522],u_xpb_out[47][522],u_xpb_out[48][522],u_xpb_out[49][522],u_xpb_out[50][522],u_xpb_out[51][522],u_xpb_out[52][522],u_xpb_out[53][522],u_xpb_out[54][522],u_xpb_out[55][522],u_xpb_out[56][522],u_xpb_out[57][522],u_xpb_out[58][522],u_xpb_out[59][522],u_xpb_out[60][522],u_xpb_out[61][522],u_xpb_out[62][522],u_xpb_out[63][522],u_xpb_out[64][522],u_xpb_out[65][522],u_xpb_out[66][522],u_xpb_out[67][522],u_xpb_out[68][522],u_xpb_out[69][522],u_xpb_out[70][522],u_xpb_out[71][522],u_xpb_out[72][522],u_xpb_out[73][522],u_xpb_out[74][522],u_xpb_out[75][522],u_xpb_out[76][522],u_xpb_out[77][522],u_xpb_out[78][522],u_xpb_out[79][522],u_xpb_out[80][522],u_xpb_out[81][522],u_xpb_out[82][522],u_xpb_out[83][522],u_xpb_out[84][522],u_xpb_out[85][522],u_xpb_out[86][522],u_xpb_out[87][522],u_xpb_out[88][522],u_xpb_out[89][522],u_xpb_out[90][522],u_xpb_out[91][522],u_xpb_out[92][522],u_xpb_out[93][522],u_xpb_out[94][522],u_xpb_out[95][522],u_xpb_out[96][522],u_xpb_out[97][522],u_xpb_out[98][522],u_xpb_out[99][522],u_xpb_out[100][522],u_xpb_out[101][522],u_xpb_out[102][522],u_xpb_out[103][522],u_xpb_out[104][522],u_xpb_out[105][522]};

assign col_out_523 = {u_xpb_out[0][523],u_xpb_out[1][523],u_xpb_out[2][523],u_xpb_out[3][523],u_xpb_out[4][523],u_xpb_out[5][523],u_xpb_out[6][523],u_xpb_out[7][523],u_xpb_out[8][523],u_xpb_out[9][523],u_xpb_out[10][523],u_xpb_out[11][523],u_xpb_out[12][523],u_xpb_out[13][523],u_xpb_out[14][523],u_xpb_out[15][523],u_xpb_out[16][523],u_xpb_out[17][523],u_xpb_out[18][523],u_xpb_out[19][523],u_xpb_out[20][523],u_xpb_out[21][523],u_xpb_out[22][523],u_xpb_out[23][523],u_xpb_out[24][523],u_xpb_out[25][523],u_xpb_out[26][523],u_xpb_out[27][523],u_xpb_out[28][523],u_xpb_out[29][523],u_xpb_out[30][523],u_xpb_out[31][523],u_xpb_out[32][523],u_xpb_out[33][523],u_xpb_out[34][523],u_xpb_out[35][523],u_xpb_out[36][523],u_xpb_out[37][523],u_xpb_out[38][523],u_xpb_out[39][523],u_xpb_out[40][523],u_xpb_out[41][523],u_xpb_out[42][523],u_xpb_out[43][523],u_xpb_out[44][523],u_xpb_out[45][523],u_xpb_out[46][523],u_xpb_out[47][523],u_xpb_out[48][523],u_xpb_out[49][523],u_xpb_out[50][523],u_xpb_out[51][523],u_xpb_out[52][523],u_xpb_out[53][523],u_xpb_out[54][523],u_xpb_out[55][523],u_xpb_out[56][523],u_xpb_out[57][523],u_xpb_out[58][523],u_xpb_out[59][523],u_xpb_out[60][523],u_xpb_out[61][523],u_xpb_out[62][523],u_xpb_out[63][523],u_xpb_out[64][523],u_xpb_out[65][523],u_xpb_out[66][523],u_xpb_out[67][523],u_xpb_out[68][523],u_xpb_out[69][523],u_xpb_out[70][523],u_xpb_out[71][523],u_xpb_out[72][523],u_xpb_out[73][523],u_xpb_out[74][523],u_xpb_out[75][523],u_xpb_out[76][523],u_xpb_out[77][523],u_xpb_out[78][523],u_xpb_out[79][523],u_xpb_out[80][523],u_xpb_out[81][523],u_xpb_out[82][523],u_xpb_out[83][523],u_xpb_out[84][523],u_xpb_out[85][523],u_xpb_out[86][523],u_xpb_out[87][523],u_xpb_out[88][523],u_xpb_out[89][523],u_xpb_out[90][523],u_xpb_out[91][523],u_xpb_out[92][523],u_xpb_out[93][523],u_xpb_out[94][523],u_xpb_out[95][523],u_xpb_out[96][523],u_xpb_out[97][523],u_xpb_out[98][523],u_xpb_out[99][523],u_xpb_out[100][523],u_xpb_out[101][523],u_xpb_out[102][523],u_xpb_out[103][523],u_xpb_out[104][523],u_xpb_out[105][523]};

assign col_out_524 = {u_xpb_out[0][524],u_xpb_out[1][524],u_xpb_out[2][524],u_xpb_out[3][524],u_xpb_out[4][524],u_xpb_out[5][524],u_xpb_out[6][524],u_xpb_out[7][524],u_xpb_out[8][524],u_xpb_out[9][524],u_xpb_out[10][524],u_xpb_out[11][524],u_xpb_out[12][524],u_xpb_out[13][524],u_xpb_out[14][524],u_xpb_out[15][524],u_xpb_out[16][524],u_xpb_out[17][524],u_xpb_out[18][524],u_xpb_out[19][524],u_xpb_out[20][524],u_xpb_out[21][524],u_xpb_out[22][524],u_xpb_out[23][524],u_xpb_out[24][524],u_xpb_out[25][524],u_xpb_out[26][524],u_xpb_out[27][524],u_xpb_out[28][524],u_xpb_out[29][524],u_xpb_out[30][524],u_xpb_out[31][524],u_xpb_out[32][524],u_xpb_out[33][524],u_xpb_out[34][524],u_xpb_out[35][524],u_xpb_out[36][524],u_xpb_out[37][524],u_xpb_out[38][524],u_xpb_out[39][524],u_xpb_out[40][524],u_xpb_out[41][524],u_xpb_out[42][524],u_xpb_out[43][524],u_xpb_out[44][524],u_xpb_out[45][524],u_xpb_out[46][524],u_xpb_out[47][524],u_xpb_out[48][524],u_xpb_out[49][524],u_xpb_out[50][524],u_xpb_out[51][524],u_xpb_out[52][524],u_xpb_out[53][524],u_xpb_out[54][524],u_xpb_out[55][524],u_xpb_out[56][524],u_xpb_out[57][524],u_xpb_out[58][524],u_xpb_out[59][524],u_xpb_out[60][524],u_xpb_out[61][524],u_xpb_out[62][524],u_xpb_out[63][524],u_xpb_out[64][524],u_xpb_out[65][524],u_xpb_out[66][524],u_xpb_out[67][524],u_xpb_out[68][524],u_xpb_out[69][524],u_xpb_out[70][524],u_xpb_out[71][524],u_xpb_out[72][524],u_xpb_out[73][524],u_xpb_out[74][524],u_xpb_out[75][524],u_xpb_out[76][524],u_xpb_out[77][524],u_xpb_out[78][524],u_xpb_out[79][524],u_xpb_out[80][524],u_xpb_out[81][524],u_xpb_out[82][524],u_xpb_out[83][524],u_xpb_out[84][524],u_xpb_out[85][524],u_xpb_out[86][524],u_xpb_out[87][524],u_xpb_out[88][524],u_xpb_out[89][524],u_xpb_out[90][524],u_xpb_out[91][524],u_xpb_out[92][524],u_xpb_out[93][524],u_xpb_out[94][524],u_xpb_out[95][524],u_xpb_out[96][524],u_xpb_out[97][524],u_xpb_out[98][524],u_xpb_out[99][524],u_xpb_out[100][524],u_xpb_out[101][524],u_xpb_out[102][524],u_xpb_out[103][524],u_xpb_out[104][524],u_xpb_out[105][524]};

assign col_out_525 = {u_xpb_out[0][525],u_xpb_out[1][525],u_xpb_out[2][525],u_xpb_out[3][525],u_xpb_out[4][525],u_xpb_out[5][525],u_xpb_out[6][525],u_xpb_out[7][525],u_xpb_out[8][525],u_xpb_out[9][525],u_xpb_out[10][525],u_xpb_out[11][525],u_xpb_out[12][525],u_xpb_out[13][525],u_xpb_out[14][525],u_xpb_out[15][525],u_xpb_out[16][525],u_xpb_out[17][525],u_xpb_out[18][525],u_xpb_out[19][525],u_xpb_out[20][525],u_xpb_out[21][525],u_xpb_out[22][525],u_xpb_out[23][525],u_xpb_out[24][525],u_xpb_out[25][525],u_xpb_out[26][525],u_xpb_out[27][525],u_xpb_out[28][525],u_xpb_out[29][525],u_xpb_out[30][525],u_xpb_out[31][525],u_xpb_out[32][525],u_xpb_out[33][525],u_xpb_out[34][525],u_xpb_out[35][525],u_xpb_out[36][525],u_xpb_out[37][525],u_xpb_out[38][525],u_xpb_out[39][525],u_xpb_out[40][525],u_xpb_out[41][525],u_xpb_out[42][525],u_xpb_out[43][525],u_xpb_out[44][525],u_xpb_out[45][525],u_xpb_out[46][525],u_xpb_out[47][525],u_xpb_out[48][525],u_xpb_out[49][525],u_xpb_out[50][525],u_xpb_out[51][525],u_xpb_out[52][525],u_xpb_out[53][525],u_xpb_out[54][525],u_xpb_out[55][525],u_xpb_out[56][525],u_xpb_out[57][525],u_xpb_out[58][525],u_xpb_out[59][525],u_xpb_out[60][525],u_xpb_out[61][525],u_xpb_out[62][525],u_xpb_out[63][525],u_xpb_out[64][525],u_xpb_out[65][525],u_xpb_out[66][525],u_xpb_out[67][525],u_xpb_out[68][525],u_xpb_out[69][525],u_xpb_out[70][525],u_xpb_out[71][525],u_xpb_out[72][525],u_xpb_out[73][525],u_xpb_out[74][525],u_xpb_out[75][525],u_xpb_out[76][525],u_xpb_out[77][525],u_xpb_out[78][525],u_xpb_out[79][525],u_xpb_out[80][525],u_xpb_out[81][525],u_xpb_out[82][525],u_xpb_out[83][525],u_xpb_out[84][525],u_xpb_out[85][525],u_xpb_out[86][525],u_xpb_out[87][525],u_xpb_out[88][525],u_xpb_out[89][525],u_xpb_out[90][525],u_xpb_out[91][525],u_xpb_out[92][525],u_xpb_out[93][525],u_xpb_out[94][525],u_xpb_out[95][525],u_xpb_out[96][525],u_xpb_out[97][525],u_xpb_out[98][525],u_xpb_out[99][525],u_xpb_out[100][525],u_xpb_out[101][525],u_xpb_out[102][525],u_xpb_out[103][525],u_xpb_out[104][525],u_xpb_out[105][525]};

assign col_out_526 = {u_xpb_out[0][526],u_xpb_out[1][526],u_xpb_out[2][526],u_xpb_out[3][526],u_xpb_out[4][526],u_xpb_out[5][526],u_xpb_out[6][526],u_xpb_out[7][526],u_xpb_out[8][526],u_xpb_out[9][526],u_xpb_out[10][526],u_xpb_out[11][526],u_xpb_out[12][526],u_xpb_out[13][526],u_xpb_out[14][526],u_xpb_out[15][526],u_xpb_out[16][526],u_xpb_out[17][526],u_xpb_out[18][526],u_xpb_out[19][526],u_xpb_out[20][526],u_xpb_out[21][526],u_xpb_out[22][526],u_xpb_out[23][526],u_xpb_out[24][526],u_xpb_out[25][526],u_xpb_out[26][526],u_xpb_out[27][526],u_xpb_out[28][526],u_xpb_out[29][526],u_xpb_out[30][526],u_xpb_out[31][526],u_xpb_out[32][526],u_xpb_out[33][526],u_xpb_out[34][526],u_xpb_out[35][526],u_xpb_out[36][526],u_xpb_out[37][526],u_xpb_out[38][526],u_xpb_out[39][526],u_xpb_out[40][526],u_xpb_out[41][526],u_xpb_out[42][526],u_xpb_out[43][526],u_xpb_out[44][526],u_xpb_out[45][526],u_xpb_out[46][526],u_xpb_out[47][526],u_xpb_out[48][526],u_xpb_out[49][526],u_xpb_out[50][526],u_xpb_out[51][526],u_xpb_out[52][526],u_xpb_out[53][526],u_xpb_out[54][526],u_xpb_out[55][526],u_xpb_out[56][526],u_xpb_out[57][526],u_xpb_out[58][526],u_xpb_out[59][526],u_xpb_out[60][526],u_xpb_out[61][526],u_xpb_out[62][526],u_xpb_out[63][526],u_xpb_out[64][526],u_xpb_out[65][526],u_xpb_out[66][526],u_xpb_out[67][526],u_xpb_out[68][526],u_xpb_out[69][526],u_xpb_out[70][526],u_xpb_out[71][526],u_xpb_out[72][526],u_xpb_out[73][526],u_xpb_out[74][526],u_xpb_out[75][526],u_xpb_out[76][526],u_xpb_out[77][526],u_xpb_out[78][526],u_xpb_out[79][526],u_xpb_out[80][526],u_xpb_out[81][526],u_xpb_out[82][526],u_xpb_out[83][526],u_xpb_out[84][526],u_xpb_out[85][526],u_xpb_out[86][526],u_xpb_out[87][526],u_xpb_out[88][526],u_xpb_out[89][526],u_xpb_out[90][526],u_xpb_out[91][526],u_xpb_out[92][526],u_xpb_out[93][526],u_xpb_out[94][526],u_xpb_out[95][526],u_xpb_out[96][526],u_xpb_out[97][526],u_xpb_out[98][526],u_xpb_out[99][526],u_xpb_out[100][526],u_xpb_out[101][526],u_xpb_out[102][526],u_xpb_out[103][526],u_xpb_out[104][526],u_xpb_out[105][526]};

assign col_out_527 = {u_xpb_out[0][527],u_xpb_out[1][527],u_xpb_out[2][527],u_xpb_out[3][527],u_xpb_out[4][527],u_xpb_out[5][527],u_xpb_out[6][527],u_xpb_out[7][527],u_xpb_out[8][527],u_xpb_out[9][527],u_xpb_out[10][527],u_xpb_out[11][527],u_xpb_out[12][527],u_xpb_out[13][527],u_xpb_out[14][527],u_xpb_out[15][527],u_xpb_out[16][527],u_xpb_out[17][527],u_xpb_out[18][527],u_xpb_out[19][527],u_xpb_out[20][527],u_xpb_out[21][527],u_xpb_out[22][527],u_xpb_out[23][527],u_xpb_out[24][527],u_xpb_out[25][527],u_xpb_out[26][527],u_xpb_out[27][527],u_xpb_out[28][527],u_xpb_out[29][527],u_xpb_out[30][527],u_xpb_out[31][527],u_xpb_out[32][527],u_xpb_out[33][527],u_xpb_out[34][527],u_xpb_out[35][527],u_xpb_out[36][527],u_xpb_out[37][527],u_xpb_out[38][527],u_xpb_out[39][527],u_xpb_out[40][527],u_xpb_out[41][527],u_xpb_out[42][527],u_xpb_out[43][527],u_xpb_out[44][527],u_xpb_out[45][527],u_xpb_out[46][527],u_xpb_out[47][527],u_xpb_out[48][527],u_xpb_out[49][527],u_xpb_out[50][527],u_xpb_out[51][527],u_xpb_out[52][527],u_xpb_out[53][527],u_xpb_out[54][527],u_xpb_out[55][527],u_xpb_out[56][527],u_xpb_out[57][527],u_xpb_out[58][527],u_xpb_out[59][527],u_xpb_out[60][527],u_xpb_out[61][527],u_xpb_out[62][527],u_xpb_out[63][527],u_xpb_out[64][527],u_xpb_out[65][527],u_xpb_out[66][527],u_xpb_out[67][527],u_xpb_out[68][527],u_xpb_out[69][527],u_xpb_out[70][527],u_xpb_out[71][527],u_xpb_out[72][527],u_xpb_out[73][527],u_xpb_out[74][527],u_xpb_out[75][527],u_xpb_out[76][527],u_xpb_out[77][527],u_xpb_out[78][527],u_xpb_out[79][527],u_xpb_out[80][527],u_xpb_out[81][527],u_xpb_out[82][527],u_xpb_out[83][527],u_xpb_out[84][527],u_xpb_out[85][527],u_xpb_out[86][527],u_xpb_out[87][527],u_xpb_out[88][527],u_xpb_out[89][527],u_xpb_out[90][527],u_xpb_out[91][527],u_xpb_out[92][527],u_xpb_out[93][527],u_xpb_out[94][527],u_xpb_out[95][527],u_xpb_out[96][527],u_xpb_out[97][527],u_xpb_out[98][527],u_xpb_out[99][527],u_xpb_out[100][527],u_xpb_out[101][527],u_xpb_out[102][527],u_xpb_out[103][527],u_xpb_out[104][527],u_xpb_out[105][527]};

assign col_out_528 = {u_xpb_out[0][528],u_xpb_out[1][528],u_xpb_out[2][528],u_xpb_out[3][528],u_xpb_out[4][528],u_xpb_out[5][528],u_xpb_out[6][528],u_xpb_out[7][528],u_xpb_out[8][528],u_xpb_out[9][528],u_xpb_out[10][528],u_xpb_out[11][528],u_xpb_out[12][528],u_xpb_out[13][528],u_xpb_out[14][528],u_xpb_out[15][528],u_xpb_out[16][528],u_xpb_out[17][528],u_xpb_out[18][528],u_xpb_out[19][528],u_xpb_out[20][528],u_xpb_out[21][528],u_xpb_out[22][528],u_xpb_out[23][528],u_xpb_out[24][528],u_xpb_out[25][528],u_xpb_out[26][528],u_xpb_out[27][528],u_xpb_out[28][528],u_xpb_out[29][528],u_xpb_out[30][528],u_xpb_out[31][528],u_xpb_out[32][528],u_xpb_out[33][528],u_xpb_out[34][528],u_xpb_out[35][528],u_xpb_out[36][528],u_xpb_out[37][528],u_xpb_out[38][528],u_xpb_out[39][528],u_xpb_out[40][528],u_xpb_out[41][528],u_xpb_out[42][528],u_xpb_out[43][528],u_xpb_out[44][528],u_xpb_out[45][528],u_xpb_out[46][528],u_xpb_out[47][528],u_xpb_out[48][528],u_xpb_out[49][528],u_xpb_out[50][528],u_xpb_out[51][528],u_xpb_out[52][528],u_xpb_out[53][528],u_xpb_out[54][528],u_xpb_out[55][528],u_xpb_out[56][528],u_xpb_out[57][528],u_xpb_out[58][528],u_xpb_out[59][528],u_xpb_out[60][528],u_xpb_out[61][528],u_xpb_out[62][528],u_xpb_out[63][528],u_xpb_out[64][528],u_xpb_out[65][528],u_xpb_out[66][528],u_xpb_out[67][528],u_xpb_out[68][528],u_xpb_out[69][528],u_xpb_out[70][528],u_xpb_out[71][528],u_xpb_out[72][528],u_xpb_out[73][528],u_xpb_out[74][528],u_xpb_out[75][528],u_xpb_out[76][528],u_xpb_out[77][528],u_xpb_out[78][528],u_xpb_out[79][528],u_xpb_out[80][528],u_xpb_out[81][528],u_xpb_out[82][528],u_xpb_out[83][528],u_xpb_out[84][528],u_xpb_out[85][528],u_xpb_out[86][528],u_xpb_out[87][528],u_xpb_out[88][528],u_xpb_out[89][528],u_xpb_out[90][528],u_xpb_out[91][528],u_xpb_out[92][528],u_xpb_out[93][528],u_xpb_out[94][528],u_xpb_out[95][528],u_xpb_out[96][528],u_xpb_out[97][528],u_xpb_out[98][528],u_xpb_out[99][528],u_xpb_out[100][528],u_xpb_out[101][528],u_xpb_out[102][528],u_xpb_out[103][528],u_xpb_out[104][528],u_xpb_out[105][528]};

assign col_out_529 = {u_xpb_out[0][529],u_xpb_out[1][529],u_xpb_out[2][529],u_xpb_out[3][529],u_xpb_out[4][529],u_xpb_out[5][529],u_xpb_out[6][529],u_xpb_out[7][529],u_xpb_out[8][529],u_xpb_out[9][529],u_xpb_out[10][529],u_xpb_out[11][529],u_xpb_out[12][529],u_xpb_out[13][529],u_xpb_out[14][529],u_xpb_out[15][529],u_xpb_out[16][529],u_xpb_out[17][529],u_xpb_out[18][529],u_xpb_out[19][529],u_xpb_out[20][529],u_xpb_out[21][529],u_xpb_out[22][529],u_xpb_out[23][529],u_xpb_out[24][529],u_xpb_out[25][529],u_xpb_out[26][529],u_xpb_out[27][529],u_xpb_out[28][529],u_xpb_out[29][529],u_xpb_out[30][529],u_xpb_out[31][529],u_xpb_out[32][529],u_xpb_out[33][529],u_xpb_out[34][529],u_xpb_out[35][529],u_xpb_out[36][529],u_xpb_out[37][529],u_xpb_out[38][529],u_xpb_out[39][529],u_xpb_out[40][529],u_xpb_out[41][529],u_xpb_out[42][529],u_xpb_out[43][529],u_xpb_out[44][529],u_xpb_out[45][529],u_xpb_out[46][529],u_xpb_out[47][529],u_xpb_out[48][529],u_xpb_out[49][529],u_xpb_out[50][529],u_xpb_out[51][529],u_xpb_out[52][529],u_xpb_out[53][529],u_xpb_out[54][529],u_xpb_out[55][529],u_xpb_out[56][529],u_xpb_out[57][529],u_xpb_out[58][529],u_xpb_out[59][529],u_xpb_out[60][529],u_xpb_out[61][529],u_xpb_out[62][529],u_xpb_out[63][529],u_xpb_out[64][529],u_xpb_out[65][529],u_xpb_out[66][529],u_xpb_out[67][529],u_xpb_out[68][529],u_xpb_out[69][529],u_xpb_out[70][529],u_xpb_out[71][529],u_xpb_out[72][529],u_xpb_out[73][529],u_xpb_out[74][529],u_xpb_out[75][529],u_xpb_out[76][529],u_xpb_out[77][529],u_xpb_out[78][529],u_xpb_out[79][529],u_xpb_out[80][529],u_xpb_out[81][529],u_xpb_out[82][529],u_xpb_out[83][529],u_xpb_out[84][529],u_xpb_out[85][529],u_xpb_out[86][529],u_xpb_out[87][529],u_xpb_out[88][529],u_xpb_out[89][529],u_xpb_out[90][529],u_xpb_out[91][529],u_xpb_out[92][529],u_xpb_out[93][529],u_xpb_out[94][529],u_xpb_out[95][529],u_xpb_out[96][529],u_xpb_out[97][529],u_xpb_out[98][529],u_xpb_out[99][529],u_xpb_out[100][529],u_xpb_out[101][529],u_xpb_out[102][529],u_xpb_out[103][529],u_xpb_out[104][529],u_xpb_out[105][529]};

assign col_out_530 = {u_xpb_out[0][530],u_xpb_out[1][530],u_xpb_out[2][530],u_xpb_out[3][530],u_xpb_out[4][530],u_xpb_out[5][530],u_xpb_out[6][530],u_xpb_out[7][530],u_xpb_out[8][530],u_xpb_out[9][530],u_xpb_out[10][530],u_xpb_out[11][530],u_xpb_out[12][530],u_xpb_out[13][530],u_xpb_out[14][530],u_xpb_out[15][530],u_xpb_out[16][530],u_xpb_out[17][530],u_xpb_out[18][530],u_xpb_out[19][530],u_xpb_out[20][530],u_xpb_out[21][530],u_xpb_out[22][530],u_xpb_out[23][530],u_xpb_out[24][530],u_xpb_out[25][530],u_xpb_out[26][530],u_xpb_out[27][530],u_xpb_out[28][530],u_xpb_out[29][530],u_xpb_out[30][530],u_xpb_out[31][530],u_xpb_out[32][530],u_xpb_out[33][530],u_xpb_out[34][530],u_xpb_out[35][530],u_xpb_out[36][530],u_xpb_out[37][530],u_xpb_out[38][530],u_xpb_out[39][530],u_xpb_out[40][530],u_xpb_out[41][530],u_xpb_out[42][530],u_xpb_out[43][530],u_xpb_out[44][530],u_xpb_out[45][530],u_xpb_out[46][530],u_xpb_out[47][530],u_xpb_out[48][530],u_xpb_out[49][530],u_xpb_out[50][530],u_xpb_out[51][530],u_xpb_out[52][530],u_xpb_out[53][530],u_xpb_out[54][530],u_xpb_out[55][530],u_xpb_out[56][530],u_xpb_out[57][530],u_xpb_out[58][530],u_xpb_out[59][530],u_xpb_out[60][530],u_xpb_out[61][530],u_xpb_out[62][530],u_xpb_out[63][530],u_xpb_out[64][530],u_xpb_out[65][530],u_xpb_out[66][530],u_xpb_out[67][530],u_xpb_out[68][530],u_xpb_out[69][530],u_xpb_out[70][530],u_xpb_out[71][530],u_xpb_out[72][530],u_xpb_out[73][530],u_xpb_out[74][530],u_xpb_out[75][530],u_xpb_out[76][530],u_xpb_out[77][530],u_xpb_out[78][530],u_xpb_out[79][530],u_xpb_out[80][530],u_xpb_out[81][530],u_xpb_out[82][530],u_xpb_out[83][530],u_xpb_out[84][530],u_xpb_out[85][530],u_xpb_out[86][530],u_xpb_out[87][530],u_xpb_out[88][530],u_xpb_out[89][530],u_xpb_out[90][530],u_xpb_out[91][530],u_xpb_out[92][530],u_xpb_out[93][530],u_xpb_out[94][530],u_xpb_out[95][530],u_xpb_out[96][530],u_xpb_out[97][530],u_xpb_out[98][530],u_xpb_out[99][530],u_xpb_out[100][530],u_xpb_out[101][530],u_xpb_out[102][530],u_xpb_out[103][530],u_xpb_out[104][530],u_xpb_out[105][530]};

assign col_out_531 = {u_xpb_out[0][531],u_xpb_out[1][531],u_xpb_out[2][531],u_xpb_out[3][531],u_xpb_out[4][531],u_xpb_out[5][531],u_xpb_out[6][531],u_xpb_out[7][531],u_xpb_out[8][531],u_xpb_out[9][531],u_xpb_out[10][531],u_xpb_out[11][531],u_xpb_out[12][531],u_xpb_out[13][531],u_xpb_out[14][531],u_xpb_out[15][531],u_xpb_out[16][531],u_xpb_out[17][531],u_xpb_out[18][531],u_xpb_out[19][531],u_xpb_out[20][531],u_xpb_out[21][531],u_xpb_out[22][531],u_xpb_out[23][531],u_xpb_out[24][531],u_xpb_out[25][531],u_xpb_out[26][531],u_xpb_out[27][531],u_xpb_out[28][531],u_xpb_out[29][531],u_xpb_out[30][531],u_xpb_out[31][531],u_xpb_out[32][531],u_xpb_out[33][531],u_xpb_out[34][531],u_xpb_out[35][531],u_xpb_out[36][531],u_xpb_out[37][531],u_xpb_out[38][531],u_xpb_out[39][531],u_xpb_out[40][531],u_xpb_out[41][531],u_xpb_out[42][531],u_xpb_out[43][531],u_xpb_out[44][531],u_xpb_out[45][531],u_xpb_out[46][531],u_xpb_out[47][531],u_xpb_out[48][531],u_xpb_out[49][531],u_xpb_out[50][531],u_xpb_out[51][531],u_xpb_out[52][531],u_xpb_out[53][531],u_xpb_out[54][531],u_xpb_out[55][531],u_xpb_out[56][531],u_xpb_out[57][531],u_xpb_out[58][531],u_xpb_out[59][531],u_xpb_out[60][531],u_xpb_out[61][531],u_xpb_out[62][531],u_xpb_out[63][531],u_xpb_out[64][531],u_xpb_out[65][531],u_xpb_out[66][531],u_xpb_out[67][531],u_xpb_out[68][531],u_xpb_out[69][531],u_xpb_out[70][531],u_xpb_out[71][531],u_xpb_out[72][531],u_xpb_out[73][531],u_xpb_out[74][531],u_xpb_out[75][531],u_xpb_out[76][531],u_xpb_out[77][531],u_xpb_out[78][531],u_xpb_out[79][531],u_xpb_out[80][531],u_xpb_out[81][531],u_xpb_out[82][531],u_xpb_out[83][531],u_xpb_out[84][531],u_xpb_out[85][531],u_xpb_out[86][531],u_xpb_out[87][531],u_xpb_out[88][531],u_xpb_out[89][531],u_xpb_out[90][531],u_xpb_out[91][531],u_xpb_out[92][531],u_xpb_out[93][531],u_xpb_out[94][531],u_xpb_out[95][531],u_xpb_out[96][531],u_xpb_out[97][531],u_xpb_out[98][531],u_xpb_out[99][531],u_xpb_out[100][531],u_xpb_out[101][531],u_xpb_out[102][531],u_xpb_out[103][531],u_xpb_out[104][531],u_xpb_out[105][531]};

assign col_out_532 = {u_xpb_out[0][532],u_xpb_out[1][532],u_xpb_out[2][532],u_xpb_out[3][532],u_xpb_out[4][532],u_xpb_out[5][532],u_xpb_out[6][532],u_xpb_out[7][532],u_xpb_out[8][532],u_xpb_out[9][532],u_xpb_out[10][532],u_xpb_out[11][532],u_xpb_out[12][532],u_xpb_out[13][532],u_xpb_out[14][532],u_xpb_out[15][532],u_xpb_out[16][532],u_xpb_out[17][532],u_xpb_out[18][532],u_xpb_out[19][532],u_xpb_out[20][532],u_xpb_out[21][532],u_xpb_out[22][532],u_xpb_out[23][532],u_xpb_out[24][532],u_xpb_out[25][532],u_xpb_out[26][532],u_xpb_out[27][532],u_xpb_out[28][532],u_xpb_out[29][532],u_xpb_out[30][532],u_xpb_out[31][532],u_xpb_out[32][532],u_xpb_out[33][532],u_xpb_out[34][532],u_xpb_out[35][532],u_xpb_out[36][532],u_xpb_out[37][532],u_xpb_out[38][532],u_xpb_out[39][532],u_xpb_out[40][532],u_xpb_out[41][532],u_xpb_out[42][532],u_xpb_out[43][532],u_xpb_out[44][532],u_xpb_out[45][532],u_xpb_out[46][532],u_xpb_out[47][532],u_xpb_out[48][532],u_xpb_out[49][532],u_xpb_out[50][532],u_xpb_out[51][532],u_xpb_out[52][532],u_xpb_out[53][532],u_xpb_out[54][532],u_xpb_out[55][532],u_xpb_out[56][532],u_xpb_out[57][532],u_xpb_out[58][532],u_xpb_out[59][532],u_xpb_out[60][532],u_xpb_out[61][532],u_xpb_out[62][532],u_xpb_out[63][532],u_xpb_out[64][532],u_xpb_out[65][532],u_xpb_out[66][532],u_xpb_out[67][532],u_xpb_out[68][532],u_xpb_out[69][532],u_xpb_out[70][532],u_xpb_out[71][532],u_xpb_out[72][532],u_xpb_out[73][532],u_xpb_out[74][532],u_xpb_out[75][532],u_xpb_out[76][532],u_xpb_out[77][532],u_xpb_out[78][532],u_xpb_out[79][532],u_xpb_out[80][532],u_xpb_out[81][532],u_xpb_out[82][532],u_xpb_out[83][532],u_xpb_out[84][532],u_xpb_out[85][532],u_xpb_out[86][532],u_xpb_out[87][532],u_xpb_out[88][532],u_xpb_out[89][532],u_xpb_out[90][532],u_xpb_out[91][532],u_xpb_out[92][532],u_xpb_out[93][532],u_xpb_out[94][532],u_xpb_out[95][532],u_xpb_out[96][532],u_xpb_out[97][532],u_xpb_out[98][532],u_xpb_out[99][532],u_xpb_out[100][532],u_xpb_out[101][532],u_xpb_out[102][532],u_xpb_out[103][532],u_xpb_out[104][532],u_xpb_out[105][532]};

assign col_out_533 = {u_xpb_out[0][533],u_xpb_out[1][533],u_xpb_out[2][533],u_xpb_out[3][533],u_xpb_out[4][533],u_xpb_out[5][533],u_xpb_out[6][533],u_xpb_out[7][533],u_xpb_out[8][533],u_xpb_out[9][533],u_xpb_out[10][533],u_xpb_out[11][533],u_xpb_out[12][533],u_xpb_out[13][533],u_xpb_out[14][533],u_xpb_out[15][533],u_xpb_out[16][533],u_xpb_out[17][533],u_xpb_out[18][533],u_xpb_out[19][533],u_xpb_out[20][533],u_xpb_out[21][533],u_xpb_out[22][533],u_xpb_out[23][533],u_xpb_out[24][533],u_xpb_out[25][533],u_xpb_out[26][533],u_xpb_out[27][533],u_xpb_out[28][533],u_xpb_out[29][533],u_xpb_out[30][533],u_xpb_out[31][533],u_xpb_out[32][533],u_xpb_out[33][533],u_xpb_out[34][533],u_xpb_out[35][533],u_xpb_out[36][533],u_xpb_out[37][533],u_xpb_out[38][533],u_xpb_out[39][533],u_xpb_out[40][533],u_xpb_out[41][533],u_xpb_out[42][533],u_xpb_out[43][533],u_xpb_out[44][533],u_xpb_out[45][533],u_xpb_out[46][533],u_xpb_out[47][533],u_xpb_out[48][533],u_xpb_out[49][533],u_xpb_out[50][533],u_xpb_out[51][533],u_xpb_out[52][533],u_xpb_out[53][533],u_xpb_out[54][533],u_xpb_out[55][533],u_xpb_out[56][533],u_xpb_out[57][533],u_xpb_out[58][533],u_xpb_out[59][533],u_xpb_out[60][533],u_xpb_out[61][533],u_xpb_out[62][533],u_xpb_out[63][533],u_xpb_out[64][533],u_xpb_out[65][533],u_xpb_out[66][533],u_xpb_out[67][533],u_xpb_out[68][533],u_xpb_out[69][533],u_xpb_out[70][533],u_xpb_out[71][533],u_xpb_out[72][533],u_xpb_out[73][533],u_xpb_out[74][533],u_xpb_out[75][533],u_xpb_out[76][533],u_xpb_out[77][533],u_xpb_out[78][533],u_xpb_out[79][533],u_xpb_out[80][533],u_xpb_out[81][533],u_xpb_out[82][533],u_xpb_out[83][533],u_xpb_out[84][533],u_xpb_out[85][533],u_xpb_out[86][533],u_xpb_out[87][533],u_xpb_out[88][533],u_xpb_out[89][533],u_xpb_out[90][533],u_xpb_out[91][533],u_xpb_out[92][533],u_xpb_out[93][533],u_xpb_out[94][533],u_xpb_out[95][533],u_xpb_out[96][533],u_xpb_out[97][533],u_xpb_out[98][533],u_xpb_out[99][533],u_xpb_out[100][533],u_xpb_out[101][533],u_xpb_out[102][533],u_xpb_out[103][533],u_xpb_out[104][533],u_xpb_out[105][533]};

assign col_out_534 = {u_xpb_out[0][534],u_xpb_out[1][534],u_xpb_out[2][534],u_xpb_out[3][534],u_xpb_out[4][534],u_xpb_out[5][534],u_xpb_out[6][534],u_xpb_out[7][534],u_xpb_out[8][534],u_xpb_out[9][534],u_xpb_out[10][534],u_xpb_out[11][534],u_xpb_out[12][534],u_xpb_out[13][534],u_xpb_out[14][534],u_xpb_out[15][534],u_xpb_out[16][534],u_xpb_out[17][534],u_xpb_out[18][534],u_xpb_out[19][534],u_xpb_out[20][534],u_xpb_out[21][534],u_xpb_out[22][534],u_xpb_out[23][534],u_xpb_out[24][534],u_xpb_out[25][534],u_xpb_out[26][534],u_xpb_out[27][534],u_xpb_out[28][534],u_xpb_out[29][534],u_xpb_out[30][534],u_xpb_out[31][534],u_xpb_out[32][534],u_xpb_out[33][534],u_xpb_out[34][534],u_xpb_out[35][534],u_xpb_out[36][534],u_xpb_out[37][534],u_xpb_out[38][534],u_xpb_out[39][534],u_xpb_out[40][534],u_xpb_out[41][534],u_xpb_out[42][534],u_xpb_out[43][534],u_xpb_out[44][534],u_xpb_out[45][534],u_xpb_out[46][534],u_xpb_out[47][534],u_xpb_out[48][534],u_xpb_out[49][534],u_xpb_out[50][534],u_xpb_out[51][534],u_xpb_out[52][534],u_xpb_out[53][534],u_xpb_out[54][534],u_xpb_out[55][534],u_xpb_out[56][534],u_xpb_out[57][534],u_xpb_out[58][534],u_xpb_out[59][534],u_xpb_out[60][534],u_xpb_out[61][534],u_xpb_out[62][534],u_xpb_out[63][534],u_xpb_out[64][534],u_xpb_out[65][534],u_xpb_out[66][534],u_xpb_out[67][534],u_xpb_out[68][534],u_xpb_out[69][534],u_xpb_out[70][534],u_xpb_out[71][534],u_xpb_out[72][534],u_xpb_out[73][534],u_xpb_out[74][534],u_xpb_out[75][534],u_xpb_out[76][534],u_xpb_out[77][534],u_xpb_out[78][534],u_xpb_out[79][534],u_xpb_out[80][534],u_xpb_out[81][534],u_xpb_out[82][534],u_xpb_out[83][534],u_xpb_out[84][534],u_xpb_out[85][534],u_xpb_out[86][534],u_xpb_out[87][534],u_xpb_out[88][534],u_xpb_out[89][534],u_xpb_out[90][534],u_xpb_out[91][534],u_xpb_out[92][534],u_xpb_out[93][534],u_xpb_out[94][534],u_xpb_out[95][534],u_xpb_out[96][534],u_xpb_out[97][534],u_xpb_out[98][534],u_xpb_out[99][534],u_xpb_out[100][534],u_xpb_out[101][534],u_xpb_out[102][534],u_xpb_out[103][534],u_xpb_out[104][534],u_xpb_out[105][534]};

assign col_out_535 = {u_xpb_out[0][535],u_xpb_out[1][535],u_xpb_out[2][535],u_xpb_out[3][535],u_xpb_out[4][535],u_xpb_out[5][535],u_xpb_out[6][535],u_xpb_out[7][535],u_xpb_out[8][535],u_xpb_out[9][535],u_xpb_out[10][535],u_xpb_out[11][535],u_xpb_out[12][535],u_xpb_out[13][535],u_xpb_out[14][535],u_xpb_out[15][535],u_xpb_out[16][535],u_xpb_out[17][535],u_xpb_out[18][535],u_xpb_out[19][535],u_xpb_out[20][535],u_xpb_out[21][535],u_xpb_out[22][535],u_xpb_out[23][535],u_xpb_out[24][535],u_xpb_out[25][535],u_xpb_out[26][535],u_xpb_out[27][535],u_xpb_out[28][535],u_xpb_out[29][535],u_xpb_out[30][535],u_xpb_out[31][535],u_xpb_out[32][535],u_xpb_out[33][535],u_xpb_out[34][535],u_xpb_out[35][535],u_xpb_out[36][535],u_xpb_out[37][535],u_xpb_out[38][535],u_xpb_out[39][535],u_xpb_out[40][535],u_xpb_out[41][535],u_xpb_out[42][535],u_xpb_out[43][535],u_xpb_out[44][535],u_xpb_out[45][535],u_xpb_out[46][535],u_xpb_out[47][535],u_xpb_out[48][535],u_xpb_out[49][535],u_xpb_out[50][535],u_xpb_out[51][535],u_xpb_out[52][535],u_xpb_out[53][535],u_xpb_out[54][535],u_xpb_out[55][535],u_xpb_out[56][535],u_xpb_out[57][535],u_xpb_out[58][535],u_xpb_out[59][535],u_xpb_out[60][535],u_xpb_out[61][535],u_xpb_out[62][535],u_xpb_out[63][535],u_xpb_out[64][535],u_xpb_out[65][535],u_xpb_out[66][535],u_xpb_out[67][535],u_xpb_out[68][535],u_xpb_out[69][535],u_xpb_out[70][535],u_xpb_out[71][535],u_xpb_out[72][535],u_xpb_out[73][535],u_xpb_out[74][535],u_xpb_out[75][535],u_xpb_out[76][535],u_xpb_out[77][535],u_xpb_out[78][535],u_xpb_out[79][535],u_xpb_out[80][535],u_xpb_out[81][535],u_xpb_out[82][535],u_xpb_out[83][535],u_xpb_out[84][535],u_xpb_out[85][535],u_xpb_out[86][535],u_xpb_out[87][535],u_xpb_out[88][535],u_xpb_out[89][535],u_xpb_out[90][535],u_xpb_out[91][535],u_xpb_out[92][535],u_xpb_out[93][535],u_xpb_out[94][535],u_xpb_out[95][535],u_xpb_out[96][535],u_xpb_out[97][535],u_xpb_out[98][535],u_xpb_out[99][535],u_xpb_out[100][535],u_xpb_out[101][535],u_xpb_out[102][535],u_xpb_out[103][535],u_xpb_out[104][535],u_xpb_out[105][535]};

assign col_out_536 = {u_xpb_out[0][536],u_xpb_out[1][536],u_xpb_out[2][536],u_xpb_out[3][536],u_xpb_out[4][536],u_xpb_out[5][536],u_xpb_out[6][536],u_xpb_out[7][536],u_xpb_out[8][536],u_xpb_out[9][536],u_xpb_out[10][536],u_xpb_out[11][536],u_xpb_out[12][536],u_xpb_out[13][536],u_xpb_out[14][536],u_xpb_out[15][536],u_xpb_out[16][536],u_xpb_out[17][536],u_xpb_out[18][536],u_xpb_out[19][536],u_xpb_out[20][536],u_xpb_out[21][536],u_xpb_out[22][536],u_xpb_out[23][536],u_xpb_out[24][536],u_xpb_out[25][536],u_xpb_out[26][536],u_xpb_out[27][536],u_xpb_out[28][536],u_xpb_out[29][536],u_xpb_out[30][536],u_xpb_out[31][536],u_xpb_out[32][536],u_xpb_out[33][536],u_xpb_out[34][536],u_xpb_out[35][536],u_xpb_out[36][536],u_xpb_out[37][536],u_xpb_out[38][536],u_xpb_out[39][536],u_xpb_out[40][536],u_xpb_out[41][536],u_xpb_out[42][536],u_xpb_out[43][536],u_xpb_out[44][536],u_xpb_out[45][536],u_xpb_out[46][536],u_xpb_out[47][536],u_xpb_out[48][536],u_xpb_out[49][536],u_xpb_out[50][536],u_xpb_out[51][536],u_xpb_out[52][536],u_xpb_out[53][536],u_xpb_out[54][536],u_xpb_out[55][536],u_xpb_out[56][536],u_xpb_out[57][536],u_xpb_out[58][536],u_xpb_out[59][536],u_xpb_out[60][536],u_xpb_out[61][536],u_xpb_out[62][536],u_xpb_out[63][536],u_xpb_out[64][536],u_xpb_out[65][536],u_xpb_out[66][536],u_xpb_out[67][536],u_xpb_out[68][536],u_xpb_out[69][536],u_xpb_out[70][536],u_xpb_out[71][536],u_xpb_out[72][536],u_xpb_out[73][536],u_xpb_out[74][536],u_xpb_out[75][536],u_xpb_out[76][536],u_xpb_out[77][536],u_xpb_out[78][536],u_xpb_out[79][536],u_xpb_out[80][536],u_xpb_out[81][536],u_xpb_out[82][536],u_xpb_out[83][536],u_xpb_out[84][536],u_xpb_out[85][536],u_xpb_out[86][536],u_xpb_out[87][536],u_xpb_out[88][536],u_xpb_out[89][536],u_xpb_out[90][536],u_xpb_out[91][536],u_xpb_out[92][536],u_xpb_out[93][536],u_xpb_out[94][536],u_xpb_out[95][536],u_xpb_out[96][536],u_xpb_out[97][536],u_xpb_out[98][536],u_xpb_out[99][536],u_xpb_out[100][536],u_xpb_out[101][536],u_xpb_out[102][536],u_xpb_out[103][536],u_xpb_out[104][536],u_xpb_out[105][536]};

assign col_out_537 = {u_xpb_out[0][537],u_xpb_out[1][537],u_xpb_out[2][537],u_xpb_out[3][537],u_xpb_out[4][537],u_xpb_out[5][537],u_xpb_out[6][537],u_xpb_out[7][537],u_xpb_out[8][537],u_xpb_out[9][537],u_xpb_out[10][537],u_xpb_out[11][537],u_xpb_out[12][537],u_xpb_out[13][537],u_xpb_out[14][537],u_xpb_out[15][537],u_xpb_out[16][537],u_xpb_out[17][537],u_xpb_out[18][537],u_xpb_out[19][537],u_xpb_out[20][537],u_xpb_out[21][537],u_xpb_out[22][537],u_xpb_out[23][537],u_xpb_out[24][537],u_xpb_out[25][537],u_xpb_out[26][537],u_xpb_out[27][537],u_xpb_out[28][537],u_xpb_out[29][537],u_xpb_out[30][537],u_xpb_out[31][537],u_xpb_out[32][537],u_xpb_out[33][537],u_xpb_out[34][537],u_xpb_out[35][537],u_xpb_out[36][537],u_xpb_out[37][537],u_xpb_out[38][537],u_xpb_out[39][537],u_xpb_out[40][537],u_xpb_out[41][537],u_xpb_out[42][537],u_xpb_out[43][537],u_xpb_out[44][537],u_xpb_out[45][537],u_xpb_out[46][537],u_xpb_out[47][537],u_xpb_out[48][537],u_xpb_out[49][537],u_xpb_out[50][537],u_xpb_out[51][537],u_xpb_out[52][537],u_xpb_out[53][537],u_xpb_out[54][537],u_xpb_out[55][537],u_xpb_out[56][537],u_xpb_out[57][537],u_xpb_out[58][537],u_xpb_out[59][537],u_xpb_out[60][537],u_xpb_out[61][537],u_xpb_out[62][537],u_xpb_out[63][537],u_xpb_out[64][537],u_xpb_out[65][537],u_xpb_out[66][537],u_xpb_out[67][537],u_xpb_out[68][537],u_xpb_out[69][537],u_xpb_out[70][537],u_xpb_out[71][537],u_xpb_out[72][537],u_xpb_out[73][537],u_xpb_out[74][537],u_xpb_out[75][537],u_xpb_out[76][537],u_xpb_out[77][537],u_xpb_out[78][537],u_xpb_out[79][537],u_xpb_out[80][537],u_xpb_out[81][537],u_xpb_out[82][537],u_xpb_out[83][537],u_xpb_out[84][537],u_xpb_out[85][537],u_xpb_out[86][537],u_xpb_out[87][537],u_xpb_out[88][537],u_xpb_out[89][537],u_xpb_out[90][537],u_xpb_out[91][537],u_xpb_out[92][537],u_xpb_out[93][537],u_xpb_out[94][537],u_xpb_out[95][537],u_xpb_out[96][537],u_xpb_out[97][537],u_xpb_out[98][537],u_xpb_out[99][537],u_xpb_out[100][537],u_xpb_out[101][537],u_xpb_out[102][537],u_xpb_out[103][537],u_xpb_out[104][537],u_xpb_out[105][537]};

assign col_out_538 = {u_xpb_out[0][538],u_xpb_out[1][538],u_xpb_out[2][538],u_xpb_out[3][538],u_xpb_out[4][538],u_xpb_out[5][538],u_xpb_out[6][538],u_xpb_out[7][538],u_xpb_out[8][538],u_xpb_out[9][538],u_xpb_out[10][538],u_xpb_out[11][538],u_xpb_out[12][538],u_xpb_out[13][538],u_xpb_out[14][538],u_xpb_out[15][538],u_xpb_out[16][538],u_xpb_out[17][538],u_xpb_out[18][538],u_xpb_out[19][538],u_xpb_out[20][538],u_xpb_out[21][538],u_xpb_out[22][538],u_xpb_out[23][538],u_xpb_out[24][538],u_xpb_out[25][538],u_xpb_out[26][538],u_xpb_out[27][538],u_xpb_out[28][538],u_xpb_out[29][538],u_xpb_out[30][538],u_xpb_out[31][538],u_xpb_out[32][538],u_xpb_out[33][538],u_xpb_out[34][538],u_xpb_out[35][538],u_xpb_out[36][538],u_xpb_out[37][538],u_xpb_out[38][538],u_xpb_out[39][538],u_xpb_out[40][538],u_xpb_out[41][538],u_xpb_out[42][538],u_xpb_out[43][538],u_xpb_out[44][538],u_xpb_out[45][538],u_xpb_out[46][538],u_xpb_out[47][538],u_xpb_out[48][538],u_xpb_out[49][538],u_xpb_out[50][538],u_xpb_out[51][538],u_xpb_out[52][538],u_xpb_out[53][538],u_xpb_out[54][538],u_xpb_out[55][538],u_xpb_out[56][538],u_xpb_out[57][538],u_xpb_out[58][538],u_xpb_out[59][538],u_xpb_out[60][538],u_xpb_out[61][538],u_xpb_out[62][538],u_xpb_out[63][538],u_xpb_out[64][538],u_xpb_out[65][538],u_xpb_out[66][538],u_xpb_out[67][538],u_xpb_out[68][538],u_xpb_out[69][538],u_xpb_out[70][538],u_xpb_out[71][538],u_xpb_out[72][538],u_xpb_out[73][538],u_xpb_out[74][538],u_xpb_out[75][538],u_xpb_out[76][538],u_xpb_out[77][538],u_xpb_out[78][538],u_xpb_out[79][538],u_xpb_out[80][538],u_xpb_out[81][538],u_xpb_out[82][538],u_xpb_out[83][538],u_xpb_out[84][538],u_xpb_out[85][538],u_xpb_out[86][538],u_xpb_out[87][538],u_xpb_out[88][538],u_xpb_out[89][538],u_xpb_out[90][538],u_xpb_out[91][538],u_xpb_out[92][538],u_xpb_out[93][538],u_xpb_out[94][538],u_xpb_out[95][538],u_xpb_out[96][538],u_xpb_out[97][538],u_xpb_out[98][538],u_xpb_out[99][538],u_xpb_out[100][538],u_xpb_out[101][538],u_xpb_out[102][538],u_xpb_out[103][538],u_xpb_out[104][538],u_xpb_out[105][538]};

assign col_out_539 = {u_xpb_out[0][539],u_xpb_out[1][539],u_xpb_out[2][539],u_xpb_out[3][539],u_xpb_out[4][539],u_xpb_out[5][539],u_xpb_out[6][539],u_xpb_out[7][539],u_xpb_out[8][539],u_xpb_out[9][539],u_xpb_out[10][539],u_xpb_out[11][539],u_xpb_out[12][539],u_xpb_out[13][539],u_xpb_out[14][539],u_xpb_out[15][539],u_xpb_out[16][539],u_xpb_out[17][539],u_xpb_out[18][539],u_xpb_out[19][539],u_xpb_out[20][539],u_xpb_out[21][539],u_xpb_out[22][539],u_xpb_out[23][539],u_xpb_out[24][539],u_xpb_out[25][539],u_xpb_out[26][539],u_xpb_out[27][539],u_xpb_out[28][539],u_xpb_out[29][539],u_xpb_out[30][539],u_xpb_out[31][539],u_xpb_out[32][539],u_xpb_out[33][539],u_xpb_out[34][539],u_xpb_out[35][539],u_xpb_out[36][539],u_xpb_out[37][539],u_xpb_out[38][539],u_xpb_out[39][539],u_xpb_out[40][539],u_xpb_out[41][539],u_xpb_out[42][539],u_xpb_out[43][539],u_xpb_out[44][539],u_xpb_out[45][539],u_xpb_out[46][539],u_xpb_out[47][539],u_xpb_out[48][539],u_xpb_out[49][539],u_xpb_out[50][539],u_xpb_out[51][539],u_xpb_out[52][539],u_xpb_out[53][539],u_xpb_out[54][539],u_xpb_out[55][539],u_xpb_out[56][539],u_xpb_out[57][539],u_xpb_out[58][539],u_xpb_out[59][539],u_xpb_out[60][539],u_xpb_out[61][539],u_xpb_out[62][539],u_xpb_out[63][539],u_xpb_out[64][539],u_xpb_out[65][539],u_xpb_out[66][539],u_xpb_out[67][539],u_xpb_out[68][539],u_xpb_out[69][539],u_xpb_out[70][539],u_xpb_out[71][539],u_xpb_out[72][539],u_xpb_out[73][539],u_xpb_out[74][539],u_xpb_out[75][539],u_xpb_out[76][539],u_xpb_out[77][539],u_xpb_out[78][539],u_xpb_out[79][539],u_xpb_out[80][539],u_xpb_out[81][539],u_xpb_out[82][539],u_xpb_out[83][539],u_xpb_out[84][539],u_xpb_out[85][539],u_xpb_out[86][539],u_xpb_out[87][539],u_xpb_out[88][539],u_xpb_out[89][539],u_xpb_out[90][539],u_xpb_out[91][539],u_xpb_out[92][539],u_xpb_out[93][539],u_xpb_out[94][539],u_xpb_out[95][539],u_xpb_out[96][539],u_xpb_out[97][539],u_xpb_out[98][539],u_xpb_out[99][539],u_xpb_out[100][539],u_xpb_out[101][539],u_xpb_out[102][539],u_xpb_out[103][539],u_xpb_out[104][539],u_xpb_out[105][539]};

assign col_out_540 = {u_xpb_out[0][540],u_xpb_out[1][540],u_xpb_out[2][540],u_xpb_out[3][540],u_xpb_out[4][540],u_xpb_out[5][540],u_xpb_out[6][540],u_xpb_out[7][540],u_xpb_out[8][540],u_xpb_out[9][540],u_xpb_out[10][540],u_xpb_out[11][540],u_xpb_out[12][540],u_xpb_out[13][540],u_xpb_out[14][540],u_xpb_out[15][540],u_xpb_out[16][540],u_xpb_out[17][540],u_xpb_out[18][540],u_xpb_out[19][540],u_xpb_out[20][540],u_xpb_out[21][540],u_xpb_out[22][540],u_xpb_out[23][540],u_xpb_out[24][540],u_xpb_out[25][540],u_xpb_out[26][540],u_xpb_out[27][540],u_xpb_out[28][540],u_xpb_out[29][540],u_xpb_out[30][540],u_xpb_out[31][540],u_xpb_out[32][540],u_xpb_out[33][540],u_xpb_out[34][540],u_xpb_out[35][540],u_xpb_out[36][540],u_xpb_out[37][540],u_xpb_out[38][540],u_xpb_out[39][540],u_xpb_out[40][540],u_xpb_out[41][540],u_xpb_out[42][540],u_xpb_out[43][540],u_xpb_out[44][540],u_xpb_out[45][540],u_xpb_out[46][540],u_xpb_out[47][540],u_xpb_out[48][540],u_xpb_out[49][540],u_xpb_out[50][540],u_xpb_out[51][540],u_xpb_out[52][540],u_xpb_out[53][540],u_xpb_out[54][540],u_xpb_out[55][540],u_xpb_out[56][540],u_xpb_out[57][540],u_xpb_out[58][540],u_xpb_out[59][540],u_xpb_out[60][540],u_xpb_out[61][540],u_xpb_out[62][540],u_xpb_out[63][540],u_xpb_out[64][540],u_xpb_out[65][540],u_xpb_out[66][540],u_xpb_out[67][540],u_xpb_out[68][540],u_xpb_out[69][540],u_xpb_out[70][540],u_xpb_out[71][540],u_xpb_out[72][540],u_xpb_out[73][540],u_xpb_out[74][540],u_xpb_out[75][540],u_xpb_out[76][540],u_xpb_out[77][540],u_xpb_out[78][540],u_xpb_out[79][540],u_xpb_out[80][540],u_xpb_out[81][540],u_xpb_out[82][540],u_xpb_out[83][540],u_xpb_out[84][540],u_xpb_out[85][540],u_xpb_out[86][540],u_xpb_out[87][540],u_xpb_out[88][540],u_xpb_out[89][540],u_xpb_out[90][540],u_xpb_out[91][540],u_xpb_out[92][540],u_xpb_out[93][540],u_xpb_out[94][540],u_xpb_out[95][540],u_xpb_out[96][540],u_xpb_out[97][540],u_xpb_out[98][540],u_xpb_out[99][540],u_xpb_out[100][540],u_xpb_out[101][540],u_xpb_out[102][540],u_xpb_out[103][540],u_xpb_out[104][540],u_xpb_out[105][540]};

assign col_out_541 = {u_xpb_out[0][541],u_xpb_out[1][541],u_xpb_out[2][541],u_xpb_out[3][541],u_xpb_out[4][541],u_xpb_out[5][541],u_xpb_out[6][541],u_xpb_out[7][541],u_xpb_out[8][541],u_xpb_out[9][541],u_xpb_out[10][541],u_xpb_out[11][541],u_xpb_out[12][541],u_xpb_out[13][541],u_xpb_out[14][541],u_xpb_out[15][541],u_xpb_out[16][541],u_xpb_out[17][541],u_xpb_out[18][541],u_xpb_out[19][541],u_xpb_out[20][541],u_xpb_out[21][541],u_xpb_out[22][541],u_xpb_out[23][541],u_xpb_out[24][541],u_xpb_out[25][541],u_xpb_out[26][541],u_xpb_out[27][541],u_xpb_out[28][541],u_xpb_out[29][541],u_xpb_out[30][541],u_xpb_out[31][541],u_xpb_out[32][541],u_xpb_out[33][541],u_xpb_out[34][541],u_xpb_out[35][541],u_xpb_out[36][541],u_xpb_out[37][541],u_xpb_out[38][541],u_xpb_out[39][541],u_xpb_out[40][541],u_xpb_out[41][541],u_xpb_out[42][541],u_xpb_out[43][541],u_xpb_out[44][541],u_xpb_out[45][541],u_xpb_out[46][541],u_xpb_out[47][541],u_xpb_out[48][541],u_xpb_out[49][541],u_xpb_out[50][541],u_xpb_out[51][541],u_xpb_out[52][541],u_xpb_out[53][541],u_xpb_out[54][541],u_xpb_out[55][541],u_xpb_out[56][541],u_xpb_out[57][541],u_xpb_out[58][541],u_xpb_out[59][541],u_xpb_out[60][541],u_xpb_out[61][541],u_xpb_out[62][541],u_xpb_out[63][541],u_xpb_out[64][541],u_xpb_out[65][541],u_xpb_out[66][541],u_xpb_out[67][541],u_xpb_out[68][541],u_xpb_out[69][541],u_xpb_out[70][541],u_xpb_out[71][541],u_xpb_out[72][541],u_xpb_out[73][541],u_xpb_out[74][541],u_xpb_out[75][541],u_xpb_out[76][541],u_xpb_out[77][541],u_xpb_out[78][541],u_xpb_out[79][541],u_xpb_out[80][541],u_xpb_out[81][541],u_xpb_out[82][541],u_xpb_out[83][541],u_xpb_out[84][541],u_xpb_out[85][541],u_xpb_out[86][541],u_xpb_out[87][541],u_xpb_out[88][541],u_xpb_out[89][541],u_xpb_out[90][541],u_xpb_out[91][541],u_xpb_out[92][541],u_xpb_out[93][541],u_xpb_out[94][541],u_xpb_out[95][541],u_xpb_out[96][541],u_xpb_out[97][541],u_xpb_out[98][541],u_xpb_out[99][541],u_xpb_out[100][541],u_xpb_out[101][541],u_xpb_out[102][541],u_xpb_out[103][541],u_xpb_out[104][541],u_xpb_out[105][541]};

assign col_out_542 = {u_xpb_out[0][542],u_xpb_out[1][542],u_xpb_out[2][542],u_xpb_out[3][542],u_xpb_out[4][542],u_xpb_out[5][542],u_xpb_out[6][542],u_xpb_out[7][542],u_xpb_out[8][542],u_xpb_out[9][542],u_xpb_out[10][542],u_xpb_out[11][542],u_xpb_out[12][542],u_xpb_out[13][542],u_xpb_out[14][542],u_xpb_out[15][542],u_xpb_out[16][542],u_xpb_out[17][542],u_xpb_out[18][542],u_xpb_out[19][542],u_xpb_out[20][542],u_xpb_out[21][542],u_xpb_out[22][542],u_xpb_out[23][542],u_xpb_out[24][542],u_xpb_out[25][542],u_xpb_out[26][542],u_xpb_out[27][542],u_xpb_out[28][542],u_xpb_out[29][542],u_xpb_out[30][542],u_xpb_out[31][542],u_xpb_out[32][542],u_xpb_out[33][542],u_xpb_out[34][542],u_xpb_out[35][542],u_xpb_out[36][542],u_xpb_out[37][542],u_xpb_out[38][542],u_xpb_out[39][542],u_xpb_out[40][542],u_xpb_out[41][542],u_xpb_out[42][542],u_xpb_out[43][542],u_xpb_out[44][542],u_xpb_out[45][542],u_xpb_out[46][542],u_xpb_out[47][542],u_xpb_out[48][542],u_xpb_out[49][542],u_xpb_out[50][542],u_xpb_out[51][542],u_xpb_out[52][542],u_xpb_out[53][542],u_xpb_out[54][542],u_xpb_out[55][542],u_xpb_out[56][542],u_xpb_out[57][542],u_xpb_out[58][542],u_xpb_out[59][542],u_xpb_out[60][542],u_xpb_out[61][542],u_xpb_out[62][542],u_xpb_out[63][542],u_xpb_out[64][542],u_xpb_out[65][542],u_xpb_out[66][542],u_xpb_out[67][542],u_xpb_out[68][542],u_xpb_out[69][542],u_xpb_out[70][542],u_xpb_out[71][542],u_xpb_out[72][542],u_xpb_out[73][542],u_xpb_out[74][542],u_xpb_out[75][542],u_xpb_out[76][542],u_xpb_out[77][542],u_xpb_out[78][542],u_xpb_out[79][542],u_xpb_out[80][542],u_xpb_out[81][542],u_xpb_out[82][542],u_xpb_out[83][542],u_xpb_out[84][542],u_xpb_out[85][542],u_xpb_out[86][542],u_xpb_out[87][542],u_xpb_out[88][542],u_xpb_out[89][542],u_xpb_out[90][542],u_xpb_out[91][542],u_xpb_out[92][542],u_xpb_out[93][542],u_xpb_out[94][542],u_xpb_out[95][542],u_xpb_out[96][542],u_xpb_out[97][542],u_xpb_out[98][542],u_xpb_out[99][542],u_xpb_out[100][542],u_xpb_out[101][542],u_xpb_out[102][542],u_xpb_out[103][542],u_xpb_out[104][542],u_xpb_out[105][542]};

assign col_out_543 = {u_xpb_out[0][543],u_xpb_out[1][543],u_xpb_out[2][543],u_xpb_out[3][543],u_xpb_out[4][543],u_xpb_out[5][543],u_xpb_out[6][543],u_xpb_out[7][543],u_xpb_out[8][543],u_xpb_out[9][543],u_xpb_out[10][543],u_xpb_out[11][543],u_xpb_out[12][543],u_xpb_out[13][543],u_xpb_out[14][543],u_xpb_out[15][543],u_xpb_out[16][543],u_xpb_out[17][543],u_xpb_out[18][543],u_xpb_out[19][543],u_xpb_out[20][543],u_xpb_out[21][543],u_xpb_out[22][543],u_xpb_out[23][543],u_xpb_out[24][543],u_xpb_out[25][543],u_xpb_out[26][543],u_xpb_out[27][543],u_xpb_out[28][543],u_xpb_out[29][543],u_xpb_out[30][543],u_xpb_out[31][543],u_xpb_out[32][543],u_xpb_out[33][543],u_xpb_out[34][543],u_xpb_out[35][543],u_xpb_out[36][543],u_xpb_out[37][543],u_xpb_out[38][543],u_xpb_out[39][543],u_xpb_out[40][543],u_xpb_out[41][543],u_xpb_out[42][543],u_xpb_out[43][543],u_xpb_out[44][543],u_xpb_out[45][543],u_xpb_out[46][543],u_xpb_out[47][543],u_xpb_out[48][543],u_xpb_out[49][543],u_xpb_out[50][543],u_xpb_out[51][543],u_xpb_out[52][543],u_xpb_out[53][543],u_xpb_out[54][543],u_xpb_out[55][543],u_xpb_out[56][543],u_xpb_out[57][543],u_xpb_out[58][543],u_xpb_out[59][543],u_xpb_out[60][543],u_xpb_out[61][543],u_xpb_out[62][543],u_xpb_out[63][543],u_xpb_out[64][543],u_xpb_out[65][543],u_xpb_out[66][543],u_xpb_out[67][543],u_xpb_out[68][543],u_xpb_out[69][543],u_xpb_out[70][543],u_xpb_out[71][543],u_xpb_out[72][543],u_xpb_out[73][543],u_xpb_out[74][543],u_xpb_out[75][543],u_xpb_out[76][543],u_xpb_out[77][543],u_xpb_out[78][543],u_xpb_out[79][543],u_xpb_out[80][543],u_xpb_out[81][543],u_xpb_out[82][543],u_xpb_out[83][543],u_xpb_out[84][543],u_xpb_out[85][543],u_xpb_out[86][543],u_xpb_out[87][543],u_xpb_out[88][543],u_xpb_out[89][543],u_xpb_out[90][543],u_xpb_out[91][543],u_xpb_out[92][543],u_xpb_out[93][543],u_xpb_out[94][543],u_xpb_out[95][543],u_xpb_out[96][543],u_xpb_out[97][543],u_xpb_out[98][543],u_xpb_out[99][543],u_xpb_out[100][543],u_xpb_out[101][543],u_xpb_out[102][543],u_xpb_out[103][543],u_xpb_out[104][543],u_xpb_out[105][543]};

assign col_out_544 = {u_xpb_out[0][544],u_xpb_out[1][544],u_xpb_out[2][544],u_xpb_out[3][544],u_xpb_out[4][544],u_xpb_out[5][544],u_xpb_out[6][544],u_xpb_out[7][544],u_xpb_out[8][544],u_xpb_out[9][544],u_xpb_out[10][544],u_xpb_out[11][544],u_xpb_out[12][544],u_xpb_out[13][544],u_xpb_out[14][544],u_xpb_out[15][544],u_xpb_out[16][544],u_xpb_out[17][544],u_xpb_out[18][544],u_xpb_out[19][544],u_xpb_out[20][544],u_xpb_out[21][544],u_xpb_out[22][544],u_xpb_out[23][544],u_xpb_out[24][544],u_xpb_out[25][544],u_xpb_out[26][544],u_xpb_out[27][544],u_xpb_out[28][544],u_xpb_out[29][544],u_xpb_out[30][544],u_xpb_out[31][544],u_xpb_out[32][544],u_xpb_out[33][544],u_xpb_out[34][544],u_xpb_out[35][544],u_xpb_out[36][544],u_xpb_out[37][544],u_xpb_out[38][544],u_xpb_out[39][544],u_xpb_out[40][544],u_xpb_out[41][544],u_xpb_out[42][544],u_xpb_out[43][544],u_xpb_out[44][544],u_xpb_out[45][544],u_xpb_out[46][544],u_xpb_out[47][544],u_xpb_out[48][544],u_xpb_out[49][544],u_xpb_out[50][544],u_xpb_out[51][544],u_xpb_out[52][544],u_xpb_out[53][544],u_xpb_out[54][544],u_xpb_out[55][544],u_xpb_out[56][544],u_xpb_out[57][544],u_xpb_out[58][544],u_xpb_out[59][544],u_xpb_out[60][544],u_xpb_out[61][544],u_xpb_out[62][544],u_xpb_out[63][544],u_xpb_out[64][544],u_xpb_out[65][544],u_xpb_out[66][544],u_xpb_out[67][544],u_xpb_out[68][544],u_xpb_out[69][544],u_xpb_out[70][544],u_xpb_out[71][544],u_xpb_out[72][544],u_xpb_out[73][544],u_xpb_out[74][544],u_xpb_out[75][544],u_xpb_out[76][544],u_xpb_out[77][544],u_xpb_out[78][544],u_xpb_out[79][544],u_xpb_out[80][544],u_xpb_out[81][544],u_xpb_out[82][544],u_xpb_out[83][544],u_xpb_out[84][544],u_xpb_out[85][544],u_xpb_out[86][544],u_xpb_out[87][544],u_xpb_out[88][544],u_xpb_out[89][544],u_xpb_out[90][544],u_xpb_out[91][544],u_xpb_out[92][544],u_xpb_out[93][544],u_xpb_out[94][544],u_xpb_out[95][544],u_xpb_out[96][544],u_xpb_out[97][544],u_xpb_out[98][544],u_xpb_out[99][544],u_xpb_out[100][544],u_xpb_out[101][544],u_xpb_out[102][544],u_xpb_out[103][544],u_xpb_out[104][544],u_xpb_out[105][544]};

assign col_out_545 = {u_xpb_out[0][545],u_xpb_out[1][545],u_xpb_out[2][545],u_xpb_out[3][545],u_xpb_out[4][545],u_xpb_out[5][545],u_xpb_out[6][545],u_xpb_out[7][545],u_xpb_out[8][545],u_xpb_out[9][545],u_xpb_out[10][545],u_xpb_out[11][545],u_xpb_out[12][545],u_xpb_out[13][545],u_xpb_out[14][545],u_xpb_out[15][545],u_xpb_out[16][545],u_xpb_out[17][545],u_xpb_out[18][545],u_xpb_out[19][545],u_xpb_out[20][545],u_xpb_out[21][545],u_xpb_out[22][545],u_xpb_out[23][545],u_xpb_out[24][545],u_xpb_out[25][545],u_xpb_out[26][545],u_xpb_out[27][545],u_xpb_out[28][545],u_xpb_out[29][545],u_xpb_out[30][545],u_xpb_out[31][545],u_xpb_out[32][545],u_xpb_out[33][545],u_xpb_out[34][545],u_xpb_out[35][545],u_xpb_out[36][545],u_xpb_out[37][545],u_xpb_out[38][545],u_xpb_out[39][545],u_xpb_out[40][545],u_xpb_out[41][545],u_xpb_out[42][545],u_xpb_out[43][545],u_xpb_out[44][545],u_xpb_out[45][545],u_xpb_out[46][545],u_xpb_out[47][545],u_xpb_out[48][545],u_xpb_out[49][545],u_xpb_out[50][545],u_xpb_out[51][545],u_xpb_out[52][545],u_xpb_out[53][545],u_xpb_out[54][545],u_xpb_out[55][545],u_xpb_out[56][545],u_xpb_out[57][545],u_xpb_out[58][545],u_xpb_out[59][545],u_xpb_out[60][545],u_xpb_out[61][545],u_xpb_out[62][545],u_xpb_out[63][545],u_xpb_out[64][545],u_xpb_out[65][545],u_xpb_out[66][545],u_xpb_out[67][545],u_xpb_out[68][545],u_xpb_out[69][545],u_xpb_out[70][545],u_xpb_out[71][545],u_xpb_out[72][545],u_xpb_out[73][545],u_xpb_out[74][545],u_xpb_out[75][545],u_xpb_out[76][545],u_xpb_out[77][545],u_xpb_out[78][545],u_xpb_out[79][545],u_xpb_out[80][545],u_xpb_out[81][545],u_xpb_out[82][545],u_xpb_out[83][545],u_xpb_out[84][545],u_xpb_out[85][545],u_xpb_out[86][545],u_xpb_out[87][545],u_xpb_out[88][545],u_xpb_out[89][545],u_xpb_out[90][545],u_xpb_out[91][545],u_xpb_out[92][545],u_xpb_out[93][545],u_xpb_out[94][545],u_xpb_out[95][545],u_xpb_out[96][545],u_xpb_out[97][545],u_xpb_out[98][545],u_xpb_out[99][545],u_xpb_out[100][545],u_xpb_out[101][545],u_xpb_out[102][545],u_xpb_out[103][545],u_xpb_out[104][545],u_xpb_out[105][545]};

assign col_out_546 = {u_xpb_out[0][546],u_xpb_out[1][546],u_xpb_out[2][546],u_xpb_out[3][546],u_xpb_out[4][546],u_xpb_out[5][546],u_xpb_out[6][546],u_xpb_out[7][546],u_xpb_out[8][546],u_xpb_out[9][546],u_xpb_out[10][546],u_xpb_out[11][546],u_xpb_out[12][546],u_xpb_out[13][546],u_xpb_out[14][546],u_xpb_out[15][546],u_xpb_out[16][546],u_xpb_out[17][546],u_xpb_out[18][546],u_xpb_out[19][546],u_xpb_out[20][546],u_xpb_out[21][546],u_xpb_out[22][546],u_xpb_out[23][546],u_xpb_out[24][546],u_xpb_out[25][546],u_xpb_out[26][546],u_xpb_out[27][546],u_xpb_out[28][546],u_xpb_out[29][546],u_xpb_out[30][546],u_xpb_out[31][546],u_xpb_out[32][546],u_xpb_out[33][546],u_xpb_out[34][546],u_xpb_out[35][546],u_xpb_out[36][546],u_xpb_out[37][546],u_xpb_out[38][546],u_xpb_out[39][546],u_xpb_out[40][546],u_xpb_out[41][546],u_xpb_out[42][546],u_xpb_out[43][546],u_xpb_out[44][546],u_xpb_out[45][546],u_xpb_out[46][546],u_xpb_out[47][546],u_xpb_out[48][546],u_xpb_out[49][546],u_xpb_out[50][546],u_xpb_out[51][546],u_xpb_out[52][546],u_xpb_out[53][546],u_xpb_out[54][546],u_xpb_out[55][546],u_xpb_out[56][546],u_xpb_out[57][546],u_xpb_out[58][546],u_xpb_out[59][546],u_xpb_out[60][546],u_xpb_out[61][546],u_xpb_out[62][546],u_xpb_out[63][546],u_xpb_out[64][546],u_xpb_out[65][546],u_xpb_out[66][546],u_xpb_out[67][546],u_xpb_out[68][546],u_xpb_out[69][546],u_xpb_out[70][546],u_xpb_out[71][546],u_xpb_out[72][546],u_xpb_out[73][546],u_xpb_out[74][546],u_xpb_out[75][546],u_xpb_out[76][546],u_xpb_out[77][546],u_xpb_out[78][546],u_xpb_out[79][546],u_xpb_out[80][546],u_xpb_out[81][546],u_xpb_out[82][546],u_xpb_out[83][546],u_xpb_out[84][546],u_xpb_out[85][546],u_xpb_out[86][546],u_xpb_out[87][546],u_xpb_out[88][546],u_xpb_out[89][546],u_xpb_out[90][546],u_xpb_out[91][546],u_xpb_out[92][546],u_xpb_out[93][546],u_xpb_out[94][546],u_xpb_out[95][546],u_xpb_out[96][546],u_xpb_out[97][546],u_xpb_out[98][546],u_xpb_out[99][546],u_xpb_out[100][546],u_xpb_out[101][546],u_xpb_out[102][546],u_xpb_out[103][546],u_xpb_out[104][546],u_xpb_out[105][546]};

assign col_out_547 = {u_xpb_out[0][547],u_xpb_out[1][547],u_xpb_out[2][547],u_xpb_out[3][547],u_xpb_out[4][547],u_xpb_out[5][547],u_xpb_out[6][547],u_xpb_out[7][547],u_xpb_out[8][547],u_xpb_out[9][547],u_xpb_out[10][547],u_xpb_out[11][547],u_xpb_out[12][547],u_xpb_out[13][547],u_xpb_out[14][547],u_xpb_out[15][547],u_xpb_out[16][547],u_xpb_out[17][547],u_xpb_out[18][547],u_xpb_out[19][547],u_xpb_out[20][547],u_xpb_out[21][547],u_xpb_out[22][547],u_xpb_out[23][547],u_xpb_out[24][547],u_xpb_out[25][547],u_xpb_out[26][547],u_xpb_out[27][547],u_xpb_out[28][547],u_xpb_out[29][547],u_xpb_out[30][547],u_xpb_out[31][547],u_xpb_out[32][547],u_xpb_out[33][547],u_xpb_out[34][547],u_xpb_out[35][547],u_xpb_out[36][547],u_xpb_out[37][547],u_xpb_out[38][547],u_xpb_out[39][547],u_xpb_out[40][547],u_xpb_out[41][547],u_xpb_out[42][547],u_xpb_out[43][547],u_xpb_out[44][547],u_xpb_out[45][547],u_xpb_out[46][547],u_xpb_out[47][547],u_xpb_out[48][547],u_xpb_out[49][547],u_xpb_out[50][547],u_xpb_out[51][547],u_xpb_out[52][547],u_xpb_out[53][547],u_xpb_out[54][547],u_xpb_out[55][547],u_xpb_out[56][547],u_xpb_out[57][547],u_xpb_out[58][547],u_xpb_out[59][547],u_xpb_out[60][547],u_xpb_out[61][547],u_xpb_out[62][547],u_xpb_out[63][547],u_xpb_out[64][547],u_xpb_out[65][547],u_xpb_out[66][547],u_xpb_out[67][547],u_xpb_out[68][547],u_xpb_out[69][547],u_xpb_out[70][547],u_xpb_out[71][547],u_xpb_out[72][547],u_xpb_out[73][547],u_xpb_out[74][547],u_xpb_out[75][547],u_xpb_out[76][547],u_xpb_out[77][547],u_xpb_out[78][547],u_xpb_out[79][547],u_xpb_out[80][547],u_xpb_out[81][547],u_xpb_out[82][547],u_xpb_out[83][547],u_xpb_out[84][547],u_xpb_out[85][547],u_xpb_out[86][547],u_xpb_out[87][547],u_xpb_out[88][547],u_xpb_out[89][547],u_xpb_out[90][547],u_xpb_out[91][547],u_xpb_out[92][547],u_xpb_out[93][547],u_xpb_out[94][547],u_xpb_out[95][547],u_xpb_out[96][547],u_xpb_out[97][547],u_xpb_out[98][547],u_xpb_out[99][547],u_xpb_out[100][547],u_xpb_out[101][547],u_xpb_out[102][547],u_xpb_out[103][547],u_xpb_out[104][547],u_xpb_out[105][547]};

assign col_out_548 = {u_xpb_out[0][548],u_xpb_out[1][548],u_xpb_out[2][548],u_xpb_out[3][548],u_xpb_out[4][548],u_xpb_out[5][548],u_xpb_out[6][548],u_xpb_out[7][548],u_xpb_out[8][548],u_xpb_out[9][548],u_xpb_out[10][548],u_xpb_out[11][548],u_xpb_out[12][548],u_xpb_out[13][548],u_xpb_out[14][548],u_xpb_out[15][548],u_xpb_out[16][548],u_xpb_out[17][548],u_xpb_out[18][548],u_xpb_out[19][548],u_xpb_out[20][548],u_xpb_out[21][548],u_xpb_out[22][548],u_xpb_out[23][548],u_xpb_out[24][548],u_xpb_out[25][548],u_xpb_out[26][548],u_xpb_out[27][548],u_xpb_out[28][548],u_xpb_out[29][548],u_xpb_out[30][548],u_xpb_out[31][548],u_xpb_out[32][548],u_xpb_out[33][548],u_xpb_out[34][548],u_xpb_out[35][548],u_xpb_out[36][548],u_xpb_out[37][548],u_xpb_out[38][548],u_xpb_out[39][548],u_xpb_out[40][548],u_xpb_out[41][548],u_xpb_out[42][548],u_xpb_out[43][548],u_xpb_out[44][548],u_xpb_out[45][548],u_xpb_out[46][548],u_xpb_out[47][548],u_xpb_out[48][548],u_xpb_out[49][548],u_xpb_out[50][548],u_xpb_out[51][548],u_xpb_out[52][548],u_xpb_out[53][548],u_xpb_out[54][548],u_xpb_out[55][548],u_xpb_out[56][548],u_xpb_out[57][548],u_xpb_out[58][548],u_xpb_out[59][548],u_xpb_out[60][548],u_xpb_out[61][548],u_xpb_out[62][548],u_xpb_out[63][548],u_xpb_out[64][548],u_xpb_out[65][548],u_xpb_out[66][548],u_xpb_out[67][548],u_xpb_out[68][548],u_xpb_out[69][548],u_xpb_out[70][548],u_xpb_out[71][548],u_xpb_out[72][548],u_xpb_out[73][548],u_xpb_out[74][548],u_xpb_out[75][548],u_xpb_out[76][548],u_xpb_out[77][548],u_xpb_out[78][548],u_xpb_out[79][548],u_xpb_out[80][548],u_xpb_out[81][548],u_xpb_out[82][548],u_xpb_out[83][548],u_xpb_out[84][548],u_xpb_out[85][548],u_xpb_out[86][548],u_xpb_out[87][548],u_xpb_out[88][548],u_xpb_out[89][548],u_xpb_out[90][548],u_xpb_out[91][548],u_xpb_out[92][548],u_xpb_out[93][548],u_xpb_out[94][548],u_xpb_out[95][548],u_xpb_out[96][548],u_xpb_out[97][548],u_xpb_out[98][548],u_xpb_out[99][548],u_xpb_out[100][548],u_xpb_out[101][548],u_xpb_out[102][548],u_xpb_out[103][548],u_xpb_out[104][548],u_xpb_out[105][548]};

assign col_out_549 = {u_xpb_out[0][549],u_xpb_out[1][549],u_xpb_out[2][549],u_xpb_out[3][549],u_xpb_out[4][549],u_xpb_out[5][549],u_xpb_out[6][549],u_xpb_out[7][549],u_xpb_out[8][549],u_xpb_out[9][549],u_xpb_out[10][549],u_xpb_out[11][549],u_xpb_out[12][549],u_xpb_out[13][549],u_xpb_out[14][549],u_xpb_out[15][549],u_xpb_out[16][549],u_xpb_out[17][549],u_xpb_out[18][549],u_xpb_out[19][549],u_xpb_out[20][549],u_xpb_out[21][549],u_xpb_out[22][549],u_xpb_out[23][549],u_xpb_out[24][549],u_xpb_out[25][549],u_xpb_out[26][549],u_xpb_out[27][549],u_xpb_out[28][549],u_xpb_out[29][549],u_xpb_out[30][549],u_xpb_out[31][549],u_xpb_out[32][549],u_xpb_out[33][549],u_xpb_out[34][549],u_xpb_out[35][549],u_xpb_out[36][549],u_xpb_out[37][549],u_xpb_out[38][549],u_xpb_out[39][549],u_xpb_out[40][549],u_xpb_out[41][549],u_xpb_out[42][549],u_xpb_out[43][549],u_xpb_out[44][549],u_xpb_out[45][549],u_xpb_out[46][549],u_xpb_out[47][549],u_xpb_out[48][549],u_xpb_out[49][549],u_xpb_out[50][549],u_xpb_out[51][549],u_xpb_out[52][549],u_xpb_out[53][549],u_xpb_out[54][549],u_xpb_out[55][549],u_xpb_out[56][549],u_xpb_out[57][549],u_xpb_out[58][549],u_xpb_out[59][549],u_xpb_out[60][549],u_xpb_out[61][549],u_xpb_out[62][549],u_xpb_out[63][549],u_xpb_out[64][549],u_xpb_out[65][549],u_xpb_out[66][549],u_xpb_out[67][549],u_xpb_out[68][549],u_xpb_out[69][549],u_xpb_out[70][549],u_xpb_out[71][549],u_xpb_out[72][549],u_xpb_out[73][549],u_xpb_out[74][549],u_xpb_out[75][549],u_xpb_out[76][549],u_xpb_out[77][549],u_xpb_out[78][549],u_xpb_out[79][549],u_xpb_out[80][549],u_xpb_out[81][549],u_xpb_out[82][549],u_xpb_out[83][549],u_xpb_out[84][549],u_xpb_out[85][549],u_xpb_out[86][549],u_xpb_out[87][549],u_xpb_out[88][549],u_xpb_out[89][549],u_xpb_out[90][549],u_xpb_out[91][549],u_xpb_out[92][549],u_xpb_out[93][549],u_xpb_out[94][549],u_xpb_out[95][549],u_xpb_out[96][549],u_xpb_out[97][549],u_xpb_out[98][549],u_xpb_out[99][549],u_xpb_out[100][549],u_xpb_out[101][549],u_xpb_out[102][549],u_xpb_out[103][549],u_xpb_out[104][549],u_xpb_out[105][549]};

assign col_out_550 = {u_xpb_out[0][550],u_xpb_out[1][550],u_xpb_out[2][550],u_xpb_out[3][550],u_xpb_out[4][550],u_xpb_out[5][550],u_xpb_out[6][550],u_xpb_out[7][550],u_xpb_out[8][550],u_xpb_out[9][550],u_xpb_out[10][550],u_xpb_out[11][550],u_xpb_out[12][550],u_xpb_out[13][550],u_xpb_out[14][550],u_xpb_out[15][550],u_xpb_out[16][550],u_xpb_out[17][550],u_xpb_out[18][550],u_xpb_out[19][550],u_xpb_out[20][550],u_xpb_out[21][550],u_xpb_out[22][550],u_xpb_out[23][550],u_xpb_out[24][550],u_xpb_out[25][550],u_xpb_out[26][550],u_xpb_out[27][550],u_xpb_out[28][550],u_xpb_out[29][550],u_xpb_out[30][550],u_xpb_out[31][550],u_xpb_out[32][550],u_xpb_out[33][550],u_xpb_out[34][550],u_xpb_out[35][550],u_xpb_out[36][550],u_xpb_out[37][550],u_xpb_out[38][550],u_xpb_out[39][550],u_xpb_out[40][550],u_xpb_out[41][550],u_xpb_out[42][550],u_xpb_out[43][550],u_xpb_out[44][550],u_xpb_out[45][550],u_xpb_out[46][550],u_xpb_out[47][550],u_xpb_out[48][550],u_xpb_out[49][550],u_xpb_out[50][550],u_xpb_out[51][550],u_xpb_out[52][550],u_xpb_out[53][550],u_xpb_out[54][550],u_xpb_out[55][550],u_xpb_out[56][550],u_xpb_out[57][550],u_xpb_out[58][550],u_xpb_out[59][550],u_xpb_out[60][550],u_xpb_out[61][550],u_xpb_out[62][550],u_xpb_out[63][550],u_xpb_out[64][550],u_xpb_out[65][550],u_xpb_out[66][550],u_xpb_out[67][550],u_xpb_out[68][550],u_xpb_out[69][550],u_xpb_out[70][550],u_xpb_out[71][550],u_xpb_out[72][550],u_xpb_out[73][550],u_xpb_out[74][550],u_xpb_out[75][550],u_xpb_out[76][550],u_xpb_out[77][550],u_xpb_out[78][550],u_xpb_out[79][550],u_xpb_out[80][550],u_xpb_out[81][550],u_xpb_out[82][550],u_xpb_out[83][550],u_xpb_out[84][550],u_xpb_out[85][550],u_xpb_out[86][550],u_xpb_out[87][550],u_xpb_out[88][550],u_xpb_out[89][550],u_xpb_out[90][550],u_xpb_out[91][550],u_xpb_out[92][550],u_xpb_out[93][550],u_xpb_out[94][550],u_xpb_out[95][550],u_xpb_out[96][550],u_xpb_out[97][550],u_xpb_out[98][550],u_xpb_out[99][550],u_xpb_out[100][550],u_xpb_out[101][550],u_xpb_out[102][550],u_xpb_out[103][550],u_xpb_out[104][550],u_xpb_out[105][550]};

assign col_out_551 = {u_xpb_out[0][551],u_xpb_out[1][551],u_xpb_out[2][551],u_xpb_out[3][551],u_xpb_out[4][551],u_xpb_out[5][551],u_xpb_out[6][551],u_xpb_out[7][551],u_xpb_out[8][551],u_xpb_out[9][551],u_xpb_out[10][551],u_xpb_out[11][551],u_xpb_out[12][551],u_xpb_out[13][551],u_xpb_out[14][551],u_xpb_out[15][551],u_xpb_out[16][551],u_xpb_out[17][551],u_xpb_out[18][551],u_xpb_out[19][551],u_xpb_out[20][551],u_xpb_out[21][551],u_xpb_out[22][551],u_xpb_out[23][551],u_xpb_out[24][551],u_xpb_out[25][551],u_xpb_out[26][551],u_xpb_out[27][551],u_xpb_out[28][551],u_xpb_out[29][551],u_xpb_out[30][551],u_xpb_out[31][551],u_xpb_out[32][551],u_xpb_out[33][551],u_xpb_out[34][551],u_xpb_out[35][551],u_xpb_out[36][551],u_xpb_out[37][551],u_xpb_out[38][551],u_xpb_out[39][551],u_xpb_out[40][551],u_xpb_out[41][551],u_xpb_out[42][551],u_xpb_out[43][551],u_xpb_out[44][551],u_xpb_out[45][551],u_xpb_out[46][551],u_xpb_out[47][551],u_xpb_out[48][551],u_xpb_out[49][551],u_xpb_out[50][551],u_xpb_out[51][551],u_xpb_out[52][551],u_xpb_out[53][551],u_xpb_out[54][551],u_xpb_out[55][551],u_xpb_out[56][551],u_xpb_out[57][551],u_xpb_out[58][551],u_xpb_out[59][551],u_xpb_out[60][551],u_xpb_out[61][551],u_xpb_out[62][551],u_xpb_out[63][551],u_xpb_out[64][551],u_xpb_out[65][551],u_xpb_out[66][551],u_xpb_out[67][551],u_xpb_out[68][551],u_xpb_out[69][551],u_xpb_out[70][551],u_xpb_out[71][551],u_xpb_out[72][551],u_xpb_out[73][551],u_xpb_out[74][551],u_xpb_out[75][551],u_xpb_out[76][551],u_xpb_out[77][551],u_xpb_out[78][551],u_xpb_out[79][551],u_xpb_out[80][551],u_xpb_out[81][551],u_xpb_out[82][551],u_xpb_out[83][551],u_xpb_out[84][551],u_xpb_out[85][551],u_xpb_out[86][551],u_xpb_out[87][551],u_xpb_out[88][551],u_xpb_out[89][551],u_xpb_out[90][551],u_xpb_out[91][551],u_xpb_out[92][551],u_xpb_out[93][551],u_xpb_out[94][551],u_xpb_out[95][551],u_xpb_out[96][551],u_xpb_out[97][551],u_xpb_out[98][551],u_xpb_out[99][551],u_xpb_out[100][551],u_xpb_out[101][551],u_xpb_out[102][551],u_xpb_out[103][551],u_xpb_out[104][551],u_xpb_out[105][551]};

assign col_out_552 = {u_xpb_out[0][552],u_xpb_out[1][552],u_xpb_out[2][552],u_xpb_out[3][552],u_xpb_out[4][552],u_xpb_out[5][552],u_xpb_out[6][552],u_xpb_out[7][552],u_xpb_out[8][552],u_xpb_out[9][552],u_xpb_out[10][552],u_xpb_out[11][552],u_xpb_out[12][552],u_xpb_out[13][552],u_xpb_out[14][552],u_xpb_out[15][552],u_xpb_out[16][552],u_xpb_out[17][552],u_xpb_out[18][552],u_xpb_out[19][552],u_xpb_out[20][552],u_xpb_out[21][552],u_xpb_out[22][552],u_xpb_out[23][552],u_xpb_out[24][552],u_xpb_out[25][552],u_xpb_out[26][552],u_xpb_out[27][552],u_xpb_out[28][552],u_xpb_out[29][552],u_xpb_out[30][552],u_xpb_out[31][552],u_xpb_out[32][552],u_xpb_out[33][552],u_xpb_out[34][552],u_xpb_out[35][552],u_xpb_out[36][552],u_xpb_out[37][552],u_xpb_out[38][552],u_xpb_out[39][552],u_xpb_out[40][552],u_xpb_out[41][552],u_xpb_out[42][552],u_xpb_out[43][552],u_xpb_out[44][552],u_xpb_out[45][552],u_xpb_out[46][552],u_xpb_out[47][552],u_xpb_out[48][552],u_xpb_out[49][552],u_xpb_out[50][552],u_xpb_out[51][552],u_xpb_out[52][552],u_xpb_out[53][552],u_xpb_out[54][552],u_xpb_out[55][552],u_xpb_out[56][552],u_xpb_out[57][552],u_xpb_out[58][552],u_xpb_out[59][552],u_xpb_out[60][552],u_xpb_out[61][552],u_xpb_out[62][552],u_xpb_out[63][552],u_xpb_out[64][552],u_xpb_out[65][552],u_xpb_out[66][552],u_xpb_out[67][552],u_xpb_out[68][552],u_xpb_out[69][552],u_xpb_out[70][552],u_xpb_out[71][552],u_xpb_out[72][552],u_xpb_out[73][552],u_xpb_out[74][552],u_xpb_out[75][552],u_xpb_out[76][552],u_xpb_out[77][552],u_xpb_out[78][552],u_xpb_out[79][552],u_xpb_out[80][552],u_xpb_out[81][552],u_xpb_out[82][552],u_xpb_out[83][552],u_xpb_out[84][552],u_xpb_out[85][552],u_xpb_out[86][552],u_xpb_out[87][552],u_xpb_out[88][552],u_xpb_out[89][552],u_xpb_out[90][552],u_xpb_out[91][552],u_xpb_out[92][552],u_xpb_out[93][552],u_xpb_out[94][552],u_xpb_out[95][552],u_xpb_out[96][552],u_xpb_out[97][552],u_xpb_out[98][552],u_xpb_out[99][552],u_xpb_out[100][552],u_xpb_out[101][552],u_xpb_out[102][552],u_xpb_out[103][552],u_xpb_out[104][552],u_xpb_out[105][552]};

assign col_out_553 = {u_xpb_out[0][553],u_xpb_out[1][553],u_xpb_out[2][553],u_xpb_out[3][553],u_xpb_out[4][553],u_xpb_out[5][553],u_xpb_out[6][553],u_xpb_out[7][553],u_xpb_out[8][553],u_xpb_out[9][553],u_xpb_out[10][553],u_xpb_out[11][553],u_xpb_out[12][553],u_xpb_out[13][553],u_xpb_out[14][553],u_xpb_out[15][553],u_xpb_out[16][553],u_xpb_out[17][553],u_xpb_out[18][553],u_xpb_out[19][553],u_xpb_out[20][553],u_xpb_out[21][553],u_xpb_out[22][553],u_xpb_out[23][553],u_xpb_out[24][553],u_xpb_out[25][553],u_xpb_out[26][553],u_xpb_out[27][553],u_xpb_out[28][553],u_xpb_out[29][553],u_xpb_out[30][553],u_xpb_out[31][553],u_xpb_out[32][553],u_xpb_out[33][553],u_xpb_out[34][553],u_xpb_out[35][553],u_xpb_out[36][553],u_xpb_out[37][553],u_xpb_out[38][553],u_xpb_out[39][553],u_xpb_out[40][553],u_xpb_out[41][553],u_xpb_out[42][553],u_xpb_out[43][553],u_xpb_out[44][553],u_xpb_out[45][553],u_xpb_out[46][553],u_xpb_out[47][553],u_xpb_out[48][553],u_xpb_out[49][553],u_xpb_out[50][553],u_xpb_out[51][553],u_xpb_out[52][553],u_xpb_out[53][553],u_xpb_out[54][553],u_xpb_out[55][553],u_xpb_out[56][553],u_xpb_out[57][553],u_xpb_out[58][553],u_xpb_out[59][553],u_xpb_out[60][553],u_xpb_out[61][553],u_xpb_out[62][553],u_xpb_out[63][553],u_xpb_out[64][553],u_xpb_out[65][553],u_xpb_out[66][553],u_xpb_out[67][553],u_xpb_out[68][553],u_xpb_out[69][553],u_xpb_out[70][553],u_xpb_out[71][553],u_xpb_out[72][553],u_xpb_out[73][553],u_xpb_out[74][553],u_xpb_out[75][553],u_xpb_out[76][553],u_xpb_out[77][553],u_xpb_out[78][553],u_xpb_out[79][553],u_xpb_out[80][553],u_xpb_out[81][553],u_xpb_out[82][553],u_xpb_out[83][553],u_xpb_out[84][553],u_xpb_out[85][553],u_xpb_out[86][553],u_xpb_out[87][553],u_xpb_out[88][553],u_xpb_out[89][553],u_xpb_out[90][553],u_xpb_out[91][553],u_xpb_out[92][553],u_xpb_out[93][553],u_xpb_out[94][553],u_xpb_out[95][553],u_xpb_out[96][553],u_xpb_out[97][553],u_xpb_out[98][553],u_xpb_out[99][553],u_xpb_out[100][553],u_xpb_out[101][553],u_xpb_out[102][553],u_xpb_out[103][553],u_xpb_out[104][553],u_xpb_out[105][553]};

assign col_out_554 = {u_xpb_out[0][554],u_xpb_out[1][554],u_xpb_out[2][554],u_xpb_out[3][554],u_xpb_out[4][554],u_xpb_out[5][554],u_xpb_out[6][554],u_xpb_out[7][554],u_xpb_out[8][554],u_xpb_out[9][554],u_xpb_out[10][554],u_xpb_out[11][554],u_xpb_out[12][554],u_xpb_out[13][554],u_xpb_out[14][554],u_xpb_out[15][554],u_xpb_out[16][554],u_xpb_out[17][554],u_xpb_out[18][554],u_xpb_out[19][554],u_xpb_out[20][554],u_xpb_out[21][554],u_xpb_out[22][554],u_xpb_out[23][554],u_xpb_out[24][554],u_xpb_out[25][554],u_xpb_out[26][554],u_xpb_out[27][554],u_xpb_out[28][554],u_xpb_out[29][554],u_xpb_out[30][554],u_xpb_out[31][554],u_xpb_out[32][554],u_xpb_out[33][554],u_xpb_out[34][554],u_xpb_out[35][554],u_xpb_out[36][554],u_xpb_out[37][554],u_xpb_out[38][554],u_xpb_out[39][554],u_xpb_out[40][554],u_xpb_out[41][554],u_xpb_out[42][554],u_xpb_out[43][554],u_xpb_out[44][554],u_xpb_out[45][554],u_xpb_out[46][554],u_xpb_out[47][554],u_xpb_out[48][554],u_xpb_out[49][554],u_xpb_out[50][554],u_xpb_out[51][554],u_xpb_out[52][554],u_xpb_out[53][554],u_xpb_out[54][554],u_xpb_out[55][554],u_xpb_out[56][554],u_xpb_out[57][554],u_xpb_out[58][554],u_xpb_out[59][554],u_xpb_out[60][554],u_xpb_out[61][554],u_xpb_out[62][554],u_xpb_out[63][554],u_xpb_out[64][554],u_xpb_out[65][554],u_xpb_out[66][554],u_xpb_out[67][554],u_xpb_out[68][554],u_xpb_out[69][554],u_xpb_out[70][554],u_xpb_out[71][554],u_xpb_out[72][554],u_xpb_out[73][554],u_xpb_out[74][554],u_xpb_out[75][554],u_xpb_out[76][554],u_xpb_out[77][554],u_xpb_out[78][554],u_xpb_out[79][554],u_xpb_out[80][554],u_xpb_out[81][554],u_xpb_out[82][554],u_xpb_out[83][554],u_xpb_out[84][554],u_xpb_out[85][554],u_xpb_out[86][554],u_xpb_out[87][554],u_xpb_out[88][554],u_xpb_out[89][554],u_xpb_out[90][554],u_xpb_out[91][554],u_xpb_out[92][554],u_xpb_out[93][554],u_xpb_out[94][554],u_xpb_out[95][554],u_xpb_out[96][554],u_xpb_out[97][554],u_xpb_out[98][554],u_xpb_out[99][554],u_xpb_out[100][554],u_xpb_out[101][554],u_xpb_out[102][554],u_xpb_out[103][554],u_xpb_out[104][554],u_xpb_out[105][554]};

assign col_out_555 = {u_xpb_out[0][555],u_xpb_out[1][555],u_xpb_out[2][555],u_xpb_out[3][555],u_xpb_out[4][555],u_xpb_out[5][555],u_xpb_out[6][555],u_xpb_out[7][555],u_xpb_out[8][555],u_xpb_out[9][555],u_xpb_out[10][555],u_xpb_out[11][555],u_xpb_out[12][555],u_xpb_out[13][555],u_xpb_out[14][555],u_xpb_out[15][555],u_xpb_out[16][555],u_xpb_out[17][555],u_xpb_out[18][555],u_xpb_out[19][555],u_xpb_out[20][555],u_xpb_out[21][555],u_xpb_out[22][555],u_xpb_out[23][555],u_xpb_out[24][555],u_xpb_out[25][555],u_xpb_out[26][555],u_xpb_out[27][555],u_xpb_out[28][555],u_xpb_out[29][555],u_xpb_out[30][555],u_xpb_out[31][555],u_xpb_out[32][555],u_xpb_out[33][555],u_xpb_out[34][555],u_xpb_out[35][555],u_xpb_out[36][555],u_xpb_out[37][555],u_xpb_out[38][555],u_xpb_out[39][555],u_xpb_out[40][555],u_xpb_out[41][555],u_xpb_out[42][555],u_xpb_out[43][555],u_xpb_out[44][555],u_xpb_out[45][555],u_xpb_out[46][555],u_xpb_out[47][555],u_xpb_out[48][555],u_xpb_out[49][555],u_xpb_out[50][555],u_xpb_out[51][555],u_xpb_out[52][555],u_xpb_out[53][555],u_xpb_out[54][555],u_xpb_out[55][555],u_xpb_out[56][555],u_xpb_out[57][555],u_xpb_out[58][555],u_xpb_out[59][555],u_xpb_out[60][555],u_xpb_out[61][555],u_xpb_out[62][555],u_xpb_out[63][555],u_xpb_out[64][555],u_xpb_out[65][555],u_xpb_out[66][555],u_xpb_out[67][555],u_xpb_out[68][555],u_xpb_out[69][555],u_xpb_out[70][555],u_xpb_out[71][555],u_xpb_out[72][555],u_xpb_out[73][555],u_xpb_out[74][555],u_xpb_out[75][555],u_xpb_out[76][555],u_xpb_out[77][555],u_xpb_out[78][555],u_xpb_out[79][555],u_xpb_out[80][555],u_xpb_out[81][555],u_xpb_out[82][555],u_xpb_out[83][555],u_xpb_out[84][555],u_xpb_out[85][555],u_xpb_out[86][555],u_xpb_out[87][555],u_xpb_out[88][555],u_xpb_out[89][555],u_xpb_out[90][555],u_xpb_out[91][555],u_xpb_out[92][555],u_xpb_out[93][555],u_xpb_out[94][555],u_xpb_out[95][555],u_xpb_out[96][555],u_xpb_out[97][555],u_xpb_out[98][555],u_xpb_out[99][555],u_xpb_out[100][555],u_xpb_out[101][555],u_xpb_out[102][555],u_xpb_out[103][555],u_xpb_out[104][555],u_xpb_out[105][555]};

assign col_out_556 = {u_xpb_out[0][556],u_xpb_out[1][556],u_xpb_out[2][556],u_xpb_out[3][556],u_xpb_out[4][556],u_xpb_out[5][556],u_xpb_out[6][556],u_xpb_out[7][556],u_xpb_out[8][556],u_xpb_out[9][556],u_xpb_out[10][556],u_xpb_out[11][556],u_xpb_out[12][556],u_xpb_out[13][556],u_xpb_out[14][556],u_xpb_out[15][556],u_xpb_out[16][556],u_xpb_out[17][556],u_xpb_out[18][556],u_xpb_out[19][556],u_xpb_out[20][556],u_xpb_out[21][556],u_xpb_out[22][556],u_xpb_out[23][556],u_xpb_out[24][556],u_xpb_out[25][556],u_xpb_out[26][556],u_xpb_out[27][556],u_xpb_out[28][556],u_xpb_out[29][556],u_xpb_out[30][556],u_xpb_out[31][556],u_xpb_out[32][556],u_xpb_out[33][556],u_xpb_out[34][556],u_xpb_out[35][556],u_xpb_out[36][556],u_xpb_out[37][556],u_xpb_out[38][556],u_xpb_out[39][556],u_xpb_out[40][556],u_xpb_out[41][556],u_xpb_out[42][556],u_xpb_out[43][556],u_xpb_out[44][556],u_xpb_out[45][556],u_xpb_out[46][556],u_xpb_out[47][556],u_xpb_out[48][556],u_xpb_out[49][556],u_xpb_out[50][556],u_xpb_out[51][556],u_xpb_out[52][556],u_xpb_out[53][556],u_xpb_out[54][556],u_xpb_out[55][556],u_xpb_out[56][556],u_xpb_out[57][556],u_xpb_out[58][556],u_xpb_out[59][556],u_xpb_out[60][556],u_xpb_out[61][556],u_xpb_out[62][556],u_xpb_out[63][556],u_xpb_out[64][556],u_xpb_out[65][556],u_xpb_out[66][556],u_xpb_out[67][556],u_xpb_out[68][556],u_xpb_out[69][556],u_xpb_out[70][556],u_xpb_out[71][556],u_xpb_out[72][556],u_xpb_out[73][556],u_xpb_out[74][556],u_xpb_out[75][556],u_xpb_out[76][556],u_xpb_out[77][556],u_xpb_out[78][556],u_xpb_out[79][556],u_xpb_out[80][556],u_xpb_out[81][556],u_xpb_out[82][556],u_xpb_out[83][556],u_xpb_out[84][556],u_xpb_out[85][556],u_xpb_out[86][556],u_xpb_out[87][556],u_xpb_out[88][556],u_xpb_out[89][556],u_xpb_out[90][556],u_xpb_out[91][556],u_xpb_out[92][556],u_xpb_out[93][556],u_xpb_out[94][556],u_xpb_out[95][556],u_xpb_out[96][556],u_xpb_out[97][556],u_xpb_out[98][556],u_xpb_out[99][556],u_xpb_out[100][556],u_xpb_out[101][556],u_xpb_out[102][556],u_xpb_out[103][556],u_xpb_out[104][556],u_xpb_out[105][556]};

assign col_out_557 = {u_xpb_out[0][557],u_xpb_out[1][557],u_xpb_out[2][557],u_xpb_out[3][557],u_xpb_out[4][557],u_xpb_out[5][557],u_xpb_out[6][557],u_xpb_out[7][557],u_xpb_out[8][557],u_xpb_out[9][557],u_xpb_out[10][557],u_xpb_out[11][557],u_xpb_out[12][557],u_xpb_out[13][557],u_xpb_out[14][557],u_xpb_out[15][557],u_xpb_out[16][557],u_xpb_out[17][557],u_xpb_out[18][557],u_xpb_out[19][557],u_xpb_out[20][557],u_xpb_out[21][557],u_xpb_out[22][557],u_xpb_out[23][557],u_xpb_out[24][557],u_xpb_out[25][557],u_xpb_out[26][557],u_xpb_out[27][557],u_xpb_out[28][557],u_xpb_out[29][557],u_xpb_out[30][557],u_xpb_out[31][557],u_xpb_out[32][557],u_xpb_out[33][557],u_xpb_out[34][557],u_xpb_out[35][557],u_xpb_out[36][557],u_xpb_out[37][557],u_xpb_out[38][557],u_xpb_out[39][557],u_xpb_out[40][557],u_xpb_out[41][557],u_xpb_out[42][557],u_xpb_out[43][557],u_xpb_out[44][557],u_xpb_out[45][557],u_xpb_out[46][557],u_xpb_out[47][557],u_xpb_out[48][557],u_xpb_out[49][557],u_xpb_out[50][557],u_xpb_out[51][557],u_xpb_out[52][557],u_xpb_out[53][557],u_xpb_out[54][557],u_xpb_out[55][557],u_xpb_out[56][557],u_xpb_out[57][557],u_xpb_out[58][557],u_xpb_out[59][557],u_xpb_out[60][557],u_xpb_out[61][557],u_xpb_out[62][557],u_xpb_out[63][557],u_xpb_out[64][557],u_xpb_out[65][557],u_xpb_out[66][557],u_xpb_out[67][557],u_xpb_out[68][557],u_xpb_out[69][557],u_xpb_out[70][557],u_xpb_out[71][557],u_xpb_out[72][557],u_xpb_out[73][557],u_xpb_out[74][557],u_xpb_out[75][557],u_xpb_out[76][557],u_xpb_out[77][557],u_xpb_out[78][557],u_xpb_out[79][557],u_xpb_out[80][557],u_xpb_out[81][557],u_xpb_out[82][557],u_xpb_out[83][557],u_xpb_out[84][557],u_xpb_out[85][557],u_xpb_out[86][557],u_xpb_out[87][557],u_xpb_out[88][557],u_xpb_out[89][557],u_xpb_out[90][557],u_xpb_out[91][557],u_xpb_out[92][557],u_xpb_out[93][557],u_xpb_out[94][557],u_xpb_out[95][557],u_xpb_out[96][557],u_xpb_out[97][557],u_xpb_out[98][557],u_xpb_out[99][557],u_xpb_out[100][557],u_xpb_out[101][557],u_xpb_out[102][557],u_xpb_out[103][557],u_xpb_out[104][557],u_xpb_out[105][557]};

assign col_out_558 = {u_xpb_out[0][558],u_xpb_out[1][558],u_xpb_out[2][558],u_xpb_out[3][558],u_xpb_out[4][558],u_xpb_out[5][558],u_xpb_out[6][558],u_xpb_out[7][558],u_xpb_out[8][558],u_xpb_out[9][558],u_xpb_out[10][558],u_xpb_out[11][558],u_xpb_out[12][558],u_xpb_out[13][558],u_xpb_out[14][558],u_xpb_out[15][558],u_xpb_out[16][558],u_xpb_out[17][558],u_xpb_out[18][558],u_xpb_out[19][558],u_xpb_out[20][558],u_xpb_out[21][558],u_xpb_out[22][558],u_xpb_out[23][558],u_xpb_out[24][558],u_xpb_out[25][558],u_xpb_out[26][558],u_xpb_out[27][558],u_xpb_out[28][558],u_xpb_out[29][558],u_xpb_out[30][558],u_xpb_out[31][558],u_xpb_out[32][558],u_xpb_out[33][558],u_xpb_out[34][558],u_xpb_out[35][558],u_xpb_out[36][558],u_xpb_out[37][558],u_xpb_out[38][558],u_xpb_out[39][558],u_xpb_out[40][558],u_xpb_out[41][558],u_xpb_out[42][558],u_xpb_out[43][558],u_xpb_out[44][558],u_xpb_out[45][558],u_xpb_out[46][558],u_xpb_out[47][558],u_xpb_out[48][558],u_xpb_out[49][558],u_xpb_out[50][558],u_xpb_out[51][558],u_xpb_out[52][558],u_xpb_out[53][558],u_xpb_out[54][558],u_xpb_out[55][558],u_xpb_out[56][558],u_xpb_out[57][558],u_xpb_out[58][558],u_xpb_out[59][558],u_xpb_out[60][558],u_xpb_out[61][558],u_xpb_out[62][558],u_xpb_out[63][558],u_xpb_out[64][558],u_xpb_out[65][558],u_xpb_out[66][558],u_xpb_out[67][558],u_xpb_out[68][558],u_xpb_out[69][558],u_xpb_out[70][558],u_xpb_out[71][558],u_xpb_out[72][558],u_xpb_out[73][558],u_xpb_out[74][558],u_xpb_out[75][558],u_xpb_out[76][558],u_xpb_out[77][558],u_xpb_out[78][558],u_xpb_out[79][558],u_xpb_out[80][558],u_xpb_out[81][558],u_xpb_out[82][558],u_xpb_out[83][558],u_xpb_out[84][558],u_xpb_out[85][558],u_xpb_out[86][558],u_xpb_out[87][558],u_xpb_out[88][558],u_xpb_out[89][558],u_xpb_out[90][558],u_xpb_out[91][558],u_xpb_out[92][558],u_xpb_out[93][558],u_xpb_out[94][558],u_xpb_out[95][558],u_xpb_out[96][558],u_xpb_out[97][558],u_xpb_out[98][558],u_xpb_out[99][558],u_xpb_out[100][558],u_xpb_out[101][558],u_xpb_out[102][558],u_xpb_out[103][558],u_xpb_out[104][558],u_xpb_out[105][558]};

assign col_out_559 = {u_xpb_out[0][559],u_xpb_out[1][559],u_xpb_out[2][559],u_xpb_out[3][559],u_xpb_out[4][559],u_xpb_out[5][559],u_xpb_out[6][559],u_xpb_out[7][559],u_xpb_out[8][559],u_xpb_out[9][559],u_xpb_out[10][559],u_xpb_out[11][559],u_xpb_out[12][559],u_xpb_out[13][559],u_xpb_out[14][559],u_xpb_out[15][559],u_xpb_out[16][559],u_xpb_out[17][559],u_xpb_out[18][559],u_xpb_out[19][559],u_xpb_out[20][559],u_xpb_out[21][559],u_xpb_out[22][559],u_xpb_out[23][559],u_xpb_out[24][559],u_xpb_out[25][559],u_xpb_out[26][559],u_xpb_out[27][559],u_xpb_out[28][559],u_xpb_out[29][559],u_xpb_out[30][559],u_xpb_out[31][559],u_xpb_out[32][559],u_xpb_out[33][559],u_xpb_out[34][559],u_xpb_out[35][559],u_xpb_out[36][559],u_xpb_out[37][559],u_xpb_out[38][559],u_xpb_out[39][559],u_xpb_out[40][559],u_xpb_out[41][559],u_xpb_out[42][559],u_xpb_out[43][559],u_xpb_out[44][559],u_xpb_out[45][559],u_xpb_out[46][559],u_xpb_out[47][559],u_xpb_out[48][559],u_xpb_out[49][559],u_xpb_out[50][559],u_xpb_out[51][559],u_xpb_out[52][559],u_xpb_out[53][559],u_xpb_out[54][559],u_xpb_out[55][559],u_xpb_out[56][559],u_xpb_out[57][559],u_xpb_out[58][559],u_xpb_out[59][559],u_xpb_out[60][559],u_xpb_out[61][559],u_xpb_out[62][559],u_xpb_out[63][559],u_xpb_out[64][559],u_xpb_out[65][559],u_xpb_out[66][559],u_xpb_out[67][559],u_xpb_out[68][559],u_xpb_out[69][559],u_xpb_out[70][559],u_xpb_out[71][559],u_xpb_out[72][559],u_xpb_out[73][559],u_xpb_out[74][559],u_xpb_out[75][559],u_xpb_out[76][559],u_xpb_out[77][559],u_xpb_out[78][559],u_xpb_out[79][559],u_xpb_out[80][559],u_xpb_out[81][559],u_xpb_out[82][559],u_xpb_out[83][559],u_xpb_out[84][559],u_xpb_out[85][559],u_xpb_out[86][559],u_xpb_out[87][559],u_xpb_out[88][559],u_xpb_out[89][559],u_xpb_out[90][559],u_xpb_out[91][559],u_xpb_out[92][559],u_xpb_out[93][559],u_xpb_out[94][559],u_xpb_out[95][559],u_xpb_out[96][559],u_xpb_out[97][559],u_xpb_out[98][559],u_xpb_out[99][559],u_xpb_out[100][559],u_xpb_out[101][559],u_xpb_out[102][559],u_xpb_out[103][559],u_xpb_out[104][559],u_xpb_out[105][559]};

assign col_out_560 = {u_xpb_out[0][560],u_xpb_out[1][560],u_xpb_out[2][560],u_xpb_out[3][560],u_xpb_out[4][560],u_xpb_out[5][560],u_xpb_out[6][560],u_xpb_out[7][560],u_xpb_out[8][560],u_xpb_out[9][560],u_xpb_out[10][560],u_xpb_out[11][560],u_xpb_out[12][560],u_xpb_out[13][560],u_xpb_out[14][560],u_xpb_out[15][560],u_xpb_out[16][560],u_xpb_out[17][560],u_xpb_out[18][560],u_xpb_out[19][560],u_xpb_out[20][560],u_xpb_out[21][560],u_xpb_out[22][560],u_xpb_out[23][560],u_xpb_out[24][560],u_xpb_out[25][560],u_xpb_out[26][560],u_xpb_out[27][560],u_xpb_out[28][560],u_xpb_out[29][560],u_xpb_out[30][560],u_xpb_out[31][560],u_xpb_out[32][560],u_xpb_out[33][560],u_xpb_out[34][560],u_xpb_out[35][560],u_xpb_out[36][560],u_xpb_out[37][560],u_xpb_out[38][560],u_xpb_out[39][560],u_xpb_out[40][560],u_xpb_out[41][560],u_xpb_out[42][560],u_xpb_out[43][560],u_xpb_out[44][560],u_xpb_out[45][560],u_xpb_out[46][560],u_xpb_out[47][560],u_xpb_out[48][560],u_xpb_out[49][560],u_xpb_out[50][560],u_xpb_out[51][560],u_xpb_out[52][560],u_xpb_out[53][560],u_xpb_out[54][560],u_xpb_out[55][560],u_xpb_out[56][560],u_xpb_out[57][560],u_xpb_out[58][560],u_xpb_out[59][560],u_xpb_out[60][560],u_xpb_out[61][560],u_xpb_out[62][560],u_xpb_out[63][560],u_xpb_out[64][560],u_xpb_out[65][560],u_xpb_out[66][560],u_xpb_out[67][560],u_xpb_out[68][560],u_xpb_out[69][560],u_xpb_out[70][560],u_xpb_out[71][560],u_xpb_out[72][560],u_xpb_out[73][560],u_xpb_out[74][560],u_xpb_out[75][560],u_xpb_out[76][560],u_xpb_out[77][560],u_xpb_out[78][560],u_xpb_out[79][560],u_xpb_out[80][560],u_xpb_out[81][560],u_xpb_out[82][560],u_xpb_out[83][560],u_xpb_out[84][560],u_xpb_out[85][560],u_xpb_out[86][560],u_xpb_out[87][560],u_xpb_out[88][560],u_xpb_out[89][560],u_xpb_out[90][560],u_xpb_out[91][560],u_xpb_out[92][560],u_xpb_out[93][560],u_xpb_out[94][560],u_xpb_out[95][560],u_xpb_out[96][560],u_xpb_out[97][560],u_xpb_out[98][560],u_xpb_out[99][560],u_xpb_out[100][560],u_xpb_out[101][560],u_xpb_out[102][560],u_xpb_out[103][560],u_xpb_out[104][560],u_xpb_out[105][560]};

assign col_out_561 = {u_xpb_out[0][561],u_xpb_out[1][561],u_xpb_out[2][561],u_xpb_out[3][561],u_xpb_out[4][561],u_xpb_out[5][561],u_xpb_out[6][561],u_xpb_out[7][561],u_xpb_out[8][561],u_xpb_out[9][561],u_xpb_out[10][561],u_xpb_out[11][561],u_xpb_out[12][561],u_xpb_out[13][561],u_xpb_out[14][561],u_xpb_out[15][561],u_xpb_out[16][561],u_xpb_out[17][561],u_xpb_out[18][561],u_xpb_out[19][561],u_xpb_out[20][561],u_xpb_out[21][561],u_xpb_out[22][561],u_xpb_out[23][561],u_xpb_out[24][561],u_xpb_out[25][561],u_xpb_out[26][561],u_xpb_out[27][561],u_xpb_out[28][561],u_xpb_out[29][561],u_xpb_out[30][561],u_xpb_out[31][561],u_xpb_out[32][561],u_xpb_out[33][561],u_xpb_out[34][561],u_xpb_out[35][561],u_xpb_out[36][561],u_xpb_out[37][561],u_xpb_out[38][561],u_xpb_out[39][561],u_xpb_out[40][561],u_xpb_out[41][561],u_xpb_out[42][561],u_xpb_out[43][561],u_xpb_out[44][561],u_xpb_out[45][561],u_xpb_out[46][561],u_xpb_out[47][561],u_xpb_out[48][561],u_xpb_out[49][561],u_xpb_out[50][561],u_xpb_out[51][561],u_xpb_out[52][561],u_xpb_out[53][561],u_xpb_out[54][561],u_xpb_out[55][561],u_xpb_out[56][561],u_xpb_out[57][561],u_xpb_out[58][561],u_xpb_out[59][561],u_xpb_out[60][561],u_xpb_out[61][561],u_xpb_out[62][561],u_xpb_out[63][561],u_xpb_out[64][561],u_xpb_out[65][561],u_xpb_out[66][561],u_xpb_out[67][561],u_xpb_out[68][561],u_xpb_out[69][561],u_xpb_out[70][561],u_xpb_out[71][561],u_xpb_out[72][561],u_xpb_out[73][561],u_xpb_out[74][561],u_xpb_out[75][561],u_xpb_out[76][561],u_xpb_out[77][561],u_xpb_out[78][561],u_xpb_out[79][561],u_xpb_out[80][561],u_xpb_out[81][561],u_xpb_out[82][561],u_xpb_out[83][561],u_xpb_out[84][561],u_xpb_out[85][561],u_xpb_out[86][561],u_xpb_out[87][561],u_xpb_out[88][561],u_xpb_out[89][561],u_xpb_out[90][561],u_xpb_out[91][561],u_xpb_out[92][561],u_xpb_out[93][561],u_xpb_out[94][561],u_xpb_out[95][561],u_xpb_out[96][561],u_xpb_out[97][561],u_xpb_out[98][561],u_xpb_out[99][561],u_xpb_out[100][561],u_xpb_out[101][561],u_xpb_out[102][561],u_xpb_out[103][561],u_xpb_out[104][561],u_xpb_out[105][561]};

assign col_out_562 = {u_xpb_out[0][562],u_xpb_out[1][562],u_xpb_out[2][562],u_xpb_out[3][562],u_xpb_out[4][562],u_xpb_out[5][562],u_xpb_out[6][562],u_xpb_out[7][562],u_xpb_out[8][562],u_xpb_out[9][562],u_xpb_out[10][562],u_xpb_out[11][562],u_xpb_out[12][562],u_xpb_out[13][562],u_xpb_out[14][562],u_xpb_out[15][562],u_xpb_out[16][562],u_xpb_out[17][562],u_xpb_out[18][562],u_xpb_out[19][562],u_xpb_out[20][562],u_xpb_out[21][562],u_xpb_out[22][562],u_xpb_out[23][562],u_xpb_out[24][562],u_xpb_out[25][562],u_xpb_out[26][562],u_xpb_out[27][562],u_xpb_out[28][562],u_xpb_out[29][562],u_xpb_out[30][562],u_xpb_out[31][562],u_xpb_out[32][562],u_xpb_out[33][562],u_xpb_out[34][562],u_xpb_out[35][562],u_xpb_out[36][562],u_xpb_out[37][562],u_xpb_out[38][562],u_xpb_out[39][562],u_xpb_out[40][562],u_xpb_out[41][562],u_xpb_out[42][562],u_xpb_out[43][562],u_xpb_out[44][562],u_xpb_out[45][562],u_xpb_out[46][562],u_xpb_out[47][562],u_xpb_out[48][562],u_xpb_out[49][562],u_xpb_out[50][562],u_xpb_out[51][562],u_xpb_out[52][562],u_xpb_out[53][562],u_xpb_out[54][562],u_xpb_out[55][562],u_xpb_out[56][562],u_xpb_out[57][562],u_xpb_out[58][562],u_xpb_out[59][562],u_xpb_out[60][562],u_xpb_out[61][562],u_xpb_out[62][562],u_xpb_out[63][562],u_xpb_out[64][562],u_xpb_out[65][562],u_xpb_out[66][562],u_xpb_out[67][562],u_xpb_out[68][562],u_xpb_out[69][562],u_xpb_out[70][562],u_xpb_out[71][562],u_xpb_out[72][562],u_xpb_out[73][562],u_xpb_out[74][562],u_xpb_out[75][562],u_xpb_out[76][562],u_xpb_out[77][562],u_xpb_out[78][562],u_xpb_out[79][562],u_xpb_out[80][562],u_xpb_out[81][562],u_xpb_out[82][562],u_xpb_out[83][562],u_xpb_out[84][562],u_xpb_out[85][562],u_xpb_out[86][562],u_xpb_out[87][562],u_xpb_out[88][562],u_xpb_out[89][562],u_xpb_out[90][562],u_xpb_out[91][562],u_xpb_out[92][562],u_xpb_out[93][562],u_xpb_out[94][562],u_xpb_out[95][562],u_xpb_out[96][562],u_xpb_out[97][562],u_xpb_out[98][562],u_xpb_out[99][562],u_xpb_out[100][562],u_xpb_out[101][562],u_xpb_out[102][562],u_xpb_out[103][562],u_xpb_out[104][562],u_xpb_out[105][562]};

assign col_out_563 = {u_xpb_out[0][563],u_xpb_out[1][563],u_xpb_out[2][563],u_xpb_out[3][563],u_xpb_out[4][563],u_xpb_out[5][563],u_xpb_out[6][563],u_xpb_out[7][563],u_xpb_out[8][563],u_xpb_out[9][563],u_xpb_out[10][563],u_xpb_out[11][563],u_xpb_out[12][563],u_xpb_out[13][563],u_xpb_out[14][563],u_xpb_out[15][563],u_xpb_out[16][563],u_xpb_out[17][563],u_xpb_out[18][563],u_xpb_out[19][563],u_xpb_out[20][563],u_xpb_out[21][563],u_xpb_out[22][563],u_xpb_out[23][563],u_xpb_out[24][563],u_xpb_out[25][563],u_xpb_out[26][563],u_xpb_out[27][563],u_xpb_out[28][563],u_xpb_out[29][563],u_xpb_out[30][563],u_xpb_out[31][563],u_xpb_out[32][563],u_xpb_out[33][563],u_xpb_out[34][563],u_xpb_out[35][563],u_xpb_out[36][563],u_xpb_out[37][563],u_xpb_out[38][563],u_xpb_out[39][563],u_xpb_out[40][563],u_xpb_out[41][563],u_xpb_out[42][563],u_xpb_out[43][563],u_xpb_out[44][563],u_xpb_out[45][563],u_xpb_out[46][563],u_xpb_out[47][563],u_xpb_out[48][563],u_xpb_out[49][563],u_xpb_out[50][563],u_xpb_out[51][563],u_xpb_out[52][563],u_xpb_out[53][563],u_xpb_out[54][563],u_xpb_out[55][563],u_xpb_out[56][563],u_xpb_out[57][563],u_xpb_out[58][563],u_xpb_out[59][563],u_xpb_out[60][563],u_xpb_out[61][563],u_xpb_out[62][563],u_xpb_out[63][563],u_xpb_out[64][563],u_xpb_out[65][563],u_xpb_out[66][563],u_xpb_out[67][563],u_xpb_out[68][563],u_xpb_out[69][563],u_xpb_out[70][563],u_xpb_out[71][563],u_xpb_out[72][563],u_xpb_out[73][563],u_xpb_out[74][563],u_xpb_out[75][563],u_xpb_out[76][563],u_xpb_out[77][563],u_xpb_out[78][563],u_xpb_out[79][563],u_xpb_out[80][563],u_xpb_out[81][563],u_xpb_out[82][563],u_xpb_out[83][563],u_xpb_out[84][563],u_xpb_out[85][563],u_xpb_out[86][563],u_xpb_out[87][563],u_xpb_out[88][563],u_xpb_out[89][563],u_xpb_out[90][563],u_xpb_out[91][563],u_xpb_out[92][563],u_xpb_out[93][563],u_xpb_out[94][563],u_xpb_out[95][563],u_xpb_out[96][563],u_xpb_out[97][563],u_xpb_out[98][563],u_xpb_out[99][563],u_xpb_out[100][563],u_xpb_out[101][563],u_xpb_out[102][563],u_xpb_out[103][563],u_xpb_out[104][563],u_xpb_out[105][563]};

assign col_out_564 = {u_xpb_out[0][564],u_xpb_out[1][564],u_xpb_out[2][564],u_xpb_out[3][564],u_xpb_out[4][564],u_xpb_out[5][564],u_xpb_out[6][564],u_xpb_out[7][564],u_xpb_out[8][564],u_xpb_out[9][564],u_xpb_out[10][564],u_xpb_out[11][564],u_xpb_out[12][564],u_xpb_out[13][564],u_xpb_out[14][564],u_xpb_out[15][564],u_xpb_out[16][564],u_xpb_out[17][564],u_xpb_out[18][564],u_xpb_out[19][564],u_xpb_out[20][564],u_xpb_out[21][564],u_xpb_out[22][564],u_xpb_out[23][564],u_xpb_out[24][564],u_xpb_out[25][564],u_xpb_out[26][564],u_xpb_out[27][564],u_xpb_out[28][564],u_xpb_out[29][564],u_xpb_out[30][564],u_xpb_out[31][564],u_xpb_out[32][564],u_xpb_out[33][564],u_xpb_out[34][564],u_xpb_out[35][564],u_xpb_out[36][564],u_xpb_out[37][564],u_xpb_out[38][564],u_xpb_out[39][564],u_xpb_out[40][564],u_xpb_out[41][564],u_xpb_out[42][564],u_xpb_out[43][564],u_xpb_out[44][564],u_xpb_out[45][564],u_xpb_out[46][564],u_xpb_out[47][564],u_xpb_out[48][564],u_xpb_out[49][564],u_xpb_out[50][564],u_xpb_out[51][564],u_xpb_out[52][564],u_xpb_out[53][564],u_xpb_out[54][564],u_xpb_out[55][564],u_xpb_out[56][564],u_xpb_out[57][564],u_xpb_out[58][564],u_xpb_out[59][564],u_xpb_out[60][564],u_xpb_out[61][564],u_xpb_out[62][564],u_xpb_out[63][564],u_xpb_out[64][564],u_xpb_out[65][564],u_xpb_out[66][564],u_xpb_out[67][564],u_xpb_out[68][564],u_xpb_out[69][564],u_xpb_out[70][564],u_xpb_out[71][564],u_xpb_out[72][564],u_xpb_out[73][564],u_xpb_out[74][564],u_xpb_out[75][564],u_xpb_out[76][564],u_xpb_out[77][564],u_xpb_out[78][564],u_xpb_out[79][564],u_xpb_out[80][564],u_xpb_out[81][564],u_xpb_out[82][564],u_xpb_out[83][564],u_xpb_out[84][564],u_xpb_out[85][564],u_xpb_out[86][564],u_xpb_out[87][564],u_xpb_out[88][564],u_xpb_out[89][564],u_xpb_out[90][564],u_xpb_out[91][564],u_xpb_out[92][564],u_xpb_out[93][564],u_xpb_out[94][564],u_xpb_out[95][564],u_xpb_out[96][564],u_xpb_out[97][564],u_xpb_out[98][564],u_xpb_out[99][564],u_xpb_out[100][564],u_xpb_out[101][564],u_xpb_out[102][564],u_xpb_out[103][564],u_xpb_out[104][564],u_xpb_out[105][564]};

assign col_out_565 = {u_xpb_out[0][565],u_xpb_out[1][565],u_xpb_out[2][565],u_xpb_out[3][565],u_xpb_out[4][565],u_xpb_out[5][565],u_xpb_out[6][565],u_xpb_out[7][565],u_xpb_out[8][565],u_xpb_out[9][565],u_xpb_out[10][565],u_xpb_out[11][565],u_xpb_out[12][565],u_xpb_out[13][565],u_xpb_out[14][565],u_xpb_out[15][565],u_xpb_out[16][565],u_xpb_out[17][565],u_xpb_out[18][565],u_xpb_out[19][565],u_xpb_out[20][565],u_xpb_out[21][565],u_xpb_out[22][565],u_xpb_out[23][565],u_xpb_out[24][565],u_xpb_out[25][565],u_xpb_out[26][565],u_xpb_out[27][565],u_xpb_out[28][565],u_xpb_out[29][565],u_xpb_out[30][565],u_xpb_out[31][565],u_xpb_out[32][565],u_xpb_out[33][565],u_xpb_out[34][565],u_xpb_out[35][565],u_xpb_out[36][565],u_xpb_out[37][565],u_xpb_out[38][565],u_xpb_out[39][565],u_xpb_out[40][565],u_xpb_out[41][565],u_xpb_out[42][565],u_xpb_out[43][565],u_xpb_out[44][565],u_xpb_out[45][565],u_xpb_out[46][565],u_xpb_out[47][565],u_xpb_out[48][565],u_xpb_out[49][565],u_xpb_out[50][565],u_xpb_out[51][565],u_xpb_out[52][565],u_xpb_out[53][565],u_xpb_out[54][565],u_xpb_out[55][565],u_xpb_out[56][565],u_xpb_out[57][565],u_xpb_out[58][565],u_xpb_out[59][565],u_xpb_out[60][565],u_xpb_out[61][565],u_xpb_out[62][565],u_xpb_out[63][565],u_xpb_out[64][565],u_xpb_out[65][565],u_xpb_out[66][565],u_xpb_out[67][565],u_xpb_out[68][565],u_xpb_out[69][565],u_xpb_out[70][565],u_xpb_out[71][565],u_xpb_out[72][565],u_xpb_out[73][565],u_xpb_out[74][565],u_xpb_out[75][565],u_xpb_out[76][565],u_xpb_out[77][565],u_xpb_out[78][565],u_xpb_out[79][565],u_xpb_out[80][565],u_xpb_out[81][565],u_xpb_out[82][565],u_xpb_out[83][565],u_xpb_out[84][565],u_xpb_out[85][565],u_xpb_out[86][565],u_xpb_out[87][565],u_xpb_out[88][565],u_xpb_out[89][565],u_xpb_out[90][565],u_xpb_out[91][565],u_xpb_out[92][565],u_xpb_out[93][565],u_xpb_out[94][565],u_xpb_out[95][565],u_xpb_out[96][565],u_xpb_out[97][565],u_xpb_out[98][565],u_xpb_out[99][565],u_xpb_out[100][565],u_xpb_out[101][565],u_xpb_out[102][565],u_xpb_out[103][565],u_xpb_out[104][565],u_xpb_out[105][565]};

assign col_out_566 = {u_xpb_out[0][566],u_xpb_out[1][566],u_xpb_out[2][566],u_xpb_out[3][566],u_xpb_out[4][566],u_xpb_out[5][566],u_xpb_out[6][566],u_xpb_out[7][566],u_xpb_out[8][566],u_xpb_out[9][566],u_xpb_out[10][566],u_xpb_out[11][566],u_xpb_out[12][566],u_xpb_out[13][566],u_xpb_out[14][566],u_xpb_out[15][566],u_xpb_out[16][566],u_xpb_out[17][566],u_xpb_out[18][566],u_xpb_out[19][566],u_xpb_out[20][566],u_xpb_out[21][566],u_xpb_out[22][566],u_xpb_out[23][566],u_xpb_out[24][566],u_xpb_out[25][566],u_xpb_out[26][566],u_xpb_out[27][566],u_xpb_out[28][566],u_xpb_out[29][566],u_xpb_out[30][566],u_xpb_out[31][566],u_xpb_out[32][566],u_xpb_out[33][566],u_xpb_out[34][566],u_xpb_out[35][566],u_xpb_out[36][566],u_xpb_out[37][566],u_xpb_out[38][566],u_xpb_out[39][566],u_xpb_out[40][566],u_xpb_out[41][566],u_xpb_out[42][566],u_xpb_out[43][566],u_xpb_out[44][566],u_xpb_out[45][566],u_xpb_out[46][566],u_xpb_out[47][566],u_xpb_out[48][566],u_xpb_out[49][566],u_xpb_out[50][566],u_xpb_out[51][566],u_xpb_out[52][566],u_xpb_out[53][566],u_xpb_out[54][566],u_xpb_out[55][566],u_xpb_out[56][566],u_xpb_out[57][566],u_xpb_out[58][566],u_xpb_out[59][566],u_xpb_out[60][566],u_xpb_out[61][566],u_xpb_out[62][566],u_xpb_out[63][566],u_xpb_out[64][566],u_xpb_out[65][566],u_xpb_out[66][566],u_xpb_out[67][566],u_xpb_out[68][566],u_xpb_out[69][566],u_xpb_out[70][566],u_xpb_out[71][566],u_xpb_out[72][566],u_xpb_out[73][566],u_xpb_out[74][566],u_xpb_out[75][566],u_xpb_out[76][566],u_xpb_out[77][566],u_xpb_out[78][566],u_xpb_out[79][566],u_xpb_out[80][566],u_xpb_out[81][566],u_xpb_out[82][566],u_xpb_out[83][566],u_xpb_out[84][566],u_xpb_out[85][566],u_xpb_out[86][566],u_xpb_out[87][566],u_xpb_out[88][566],u_xpb_out[89][566],u_xpb_out[90][566],u_xpb_out[91][566],u_xpb_out[92][566],u_xpb_out[93][566],u_xpb_out[94][566],u_xpb_out[95][566],u_xpb_out[96][566],u_xpb_out[97][566],u_xpb_out[98][566],u_xpb_out[99][566],u_xpb_out[100][566],u_xpb_out[101][566],u_xpb_out[102][566],u_xpb_out[103][566],u_xpb_out[104][566],u_xpb_out[105][566]};

assign col_out_567 = {u_xpb_out[0][567],u_xpb_out[1][567],u_xpb_out[2][567],u_xpb_out[3][567],u_xpb_out[4][567],u_xpb_out[5][567],u_xpb_out[6][567],u_xpb_out[7][567],u_xpb_out[8][567],u_xpb_out[9][567],u_xpb_out[10][567],u_xpb_out[11][567],u_xpb_out[12][567],u_xpb_out[13][567],u_xpb_out[14][567],u_xpb_out[15][567],u_xpb_out[16][567],u_xpb_out[17][567],u_xpb_out[18][567],u_xpb_out[19][567],u_xpb_out[20][567],u_xpb_out[21][567],u_xpb_out[22][567],u_xpb_out[23][567],u_xpb_out[24][567],u_xpb_out[25][567],u_xpb_out[26][567],u_xpb_out[27][567],u_xpb_out[28][567],u_xpb_out[29][567],u_xpb_out[30][567],u_xpb_out[31][567],u_xpb_out[32][567],u_xpb_out[33][567],u_xpb_out[34][567],u_xpb_out[35][567],u_xpb_out[36][567],u_xpb_out[37][567],u_xpb_out[38][567],u_xpb_out[39][567],u_xpb_out[40][567],u_xpb_out[41][567],u_xpb_out[42][567],u_xpb_out[43][567],u_xpb_out[44][567],u_xpb_out[45][567],u_xpb_out[46][567],u_xpb_out[47][567],u_xpb_out[48][567],u_xpb_out[49][567],u_xpb_out[50][567],u_xpb_out[51][567],u_xpb_out[52][567],u_xpb_out[53][567],u_xpb_out[54][567],u_xpb_out[55][567],u_xpb_out[56][567],u_xpb_out[57][567],u_xpb_out[58][567],u_xpb_out[59][567],u_xpb_out[60][567],u_xpb_out[61][567],u_xpb_out[62][567],u_xpb_out[63][567],u_xpb_out[64][567],u_xpb_out[65][567],u_xpb_out[66][567],u_xpb_out[67][567],u_xpb_out[68][567],u_xpb_out[69][567],u_xpb_out[70][567],u_xpb_out[71][567],u_xpb_out[72][567],u_xpb_out[73][567],u_xpb_out[74][567],u_xpb_out[75][567],u_xpb_out[76][567],u_xpb_out[77][567],u_xpb_out[78][567],u_xpb_out[79][567],u_xpb_out[80][567],u_xpb_out[81][567],u_xpb_out[82][567],u_xpb_out[83][567],u_xpb_out[84][567],u_xpb_out[85][567],u_xpb_out[86][567],u_xpb_out[87][567],u_xpb_out[88][567],u_xpb_out[89][567],u_xpb_out[90][567],u_xpb_out[91][567],u_xpb_out[92][567],u_xpb_out[93][567],u_xpb_out[94][567],u_xpb_out[95][567],u_xpb_out[96][567],u_xpb_out[97][567],u_xpb_out[98][567],u_xpb_out[99][567],u_xpb_out[100][567],u_xpb_out[101][567],u_xpb_out[102][567],u_xpb_out[103][567],u_xpb_out[104][567],u_xpb_out[105][567]};

assign col_out_568 = {u_xpb_out[0][568],u_xpb_out[1][568],u_xpb_out[2][568],u_xpb_out[3][568],u_xpb_out[4][568],u_xpb_out[5][568],u_xpb_out[6][568],u_xpb_out[7][568],u_xpb_out[8][568],u_xpb_out[9][568],u_xpb_out[10][568],u_xpb_out[11][568],u_xpb_out[12][568],u_xpb_out[13][568],u_xpb_out[14][568],u_xpb_out[15][568],u_xpb_out[16][568],u_xpb_out[17][568],u_xpb_out[18][568],u_xpb_out[19][568],u_xpb_out[20][568],u_xpb_out[21][568],u_xpb_out[22][568],u_xpb_out[23][568],u_xpb_out[24][568],u_xpb_out[25][568],u_xpb_out[26][568],u_xpb_out[27][568],u_xpb_out[28][568],u_xpb_out[29][568],u_xpb_out[30][568],u_xpb_out[31][568],u_xpb_out[32][568],u_xpb_out[33][568],u_xpb_out[34][568],u_xpb_out[35][568],u_xpb_out[36][568],u_xpb_out[37][568],u_xpb_out[38][568],u_xpb_out[39][568],u_xpb_out[40][568],u_xpb_out[41][568],u_xpb_out[42][568],u_xpb_out[43][568],u_xpb_out[44][568],u_xpb_out[45][568],u_xpb_out[46][568],u_xpb_out[47][568],u_xpb_out[48][568],u_xpb_out[49][568],u_xpb_out[50][568],u_xpb_out[51][568],u_xpb_out[52][568],u_xpb_out[53][568],u_xpb_out[54][568],u_xpb_out[55][568],u_xpb_out[56][568],u_xpb_out[57][568],u_xpb_out[58][568],u_xpb_out[59][568],u_xpb_out[60][568],u_xpb_out[61][568],u_xpb_out[62][568],u_xpb_out[63][568],u_xpb_out[64][568],u_xpb_out[65][568],u_xpb_out[66][568],u_xpb_out[67][568],u_xpb_out[68][568],u_xpb_out[69][568],u_xpb_out[70][568],u_xpb_out[71][568],u_xpb_out[72][568],u_xpb_out[73][568],u_xpb_out[74][568],u_xpb_out[75][568],u_xpb_out[76][568],u_xpb_out[77][568],u_xpb_out[78][568],u_xpb_out[79][568],u_xpb_out[80][568],u_xpb_out[81][568],u_xpb_out[82][568],u_xpb_out[83][568],u_xpb_out[84][568],u_xpb_out[85][568],u_xpb_out[86][568],u_xpb_out[87][568],u_xpb_out[88][568],u_xpb_out[89][568],u_xpb_out[90][568],u_xpb_out[91][568],u_xpb_out[92][568],u_xpb_out[93][568],u_xpb_out[94][568],u_xpb_out[95][568],u_xpb_out[96][568],u_xpb_out[97][568],u_xpb_out[98][568],u_xpb_out[99][568],u_xpb_out[100][568],u_xpb_out[101][568],u_xpb_out[102][568],u_xpb_out[103][568],u_xpb_out[104][568],u_xpb_out[105][568]};

assign col_out_569 = {u_xpb_out[0][569],u_xpb_out[1][569],u_xpb_out[2][569],u_xpb_out[3][569],u_xpb_out[4][569],u_xpb_out[5][569],u_xpb_out[6][569],u_xpb_out[7][569],u_xpb_out[8][569],u_xpb_out[9][569],u_xpb_out[10][569],u_xpb_out[11][569],u_xpb_out[12][569],u_xpb_out[13][569],u_xpb_out[14][569],u_xpb_out[15][569],u_xpb_out[16][569],u_xpb_out[17][569],u_xpb_out[18][569],u_xpb_out[19][569],u_xpb_out[20][569],u_xpb_out[21][569],u_xpb_out[22][569],u_xpb_out[23][569],u_xpb_out[24][569],u_xpb_out[25][569],u_xpb_out[26][569],u_xpb_out[27][569],u_xpb_out[28][569],u_xpb_out[29][569],u_xpb_out[30][569],u_xpb_out[31][569],u_xpb_out[32][569],u_xpb_out[33][569],u_xpb_out[34][569],u_xpb_out[35][569],u_xpb_out[36][569],u_xpb_out[37][569],u_xpb_out[38][569],u_xpb_out[39][569],u_xpb_out[40][569],u_xpb_out[41][569],u_xpb_out[42][569],u_xpb_out[43][569],u_xpb_out[44][569],u_xpb_out[45][569],u_xpb_out[46][569],u_xpb_out[47][569],u_xpb_out[48][569],u_xpb_out[49][569],u_xpb_out[50][569],u_xpb_out[51][569],u_xpb_out[52][569],u_xpb_out[53][569],u_xpb_out[54][569],u_xpb_out[55][569],u_xpb_out[56][569],u_xpb_out[57][569],u_xpb_out[58][569],u_xpb_out[59][569],u_xpb_out[60][569],u_xpb_out[61][569],u_xpb_out[62][569],u_xpb_out[63][569],u_xpb_out[64][569],u_xpb_out[65][569],u_xpb_out[66][569],u_xpb_out[67][569],u_xpb_out[68][569],u_xpb_out[69][569],u_xpb_out[70][569],u_xpb_out[71][569],u_xpb_out[72][569],u_xpb_out[73][569],u_xpb_out[74][569],u_xpb_out[75][569],u_xpb_out[76][569],u_xpb_out[77][569],u_xpb_out[78][569],u_xpb_out[79][569],u_xpb_out[80][569],u_xpb_out[81][569],u_xpb_out[82][569],u_xpb_out[83][569],u_xpb_out[84][569],u_xpb_out[85][569],u_xpb_out[86][569],u_xpb_out[87][569],u_xpb_out[88][569],u_xpb_out[89][569],u_xpb_out[90][569],u_xpb_out[91][569],u_xpb_out[92][569],u_xpb_out[93][569],u_xpb_out[94][569],u_xpb_out[95][569],u_xpb_out[96][569],u_xpb_out[97][569],u_xpb_out[98][569],u_xpb_out[99][569],u_xpb_out[100][569],u_xpb_out[101][569],u_xpb_out[102][569],u_xpb_out[103][569],u_xpb_out[104][569],u_xpb_out[105][569]};

assign col_out_570 = {u_xpb_out[0][570],u_xpb_out[1][570],u_xpb_out[2][570],u_xpb_out[3][570],u_xpb_out[4][570],u_xpb_out[5][570],u_xpb_out[6][570],u_xpb_out[7][570],u_xpb_out[8][570],u_xpb_out[9][570],u_xpb_out[10][570],u_xpb_out[11][570],u_xpb_out[12][570],u_xpb_out[13][570],u_xpb_out[14][570],u_xpb_out[15][570],u_xpb_out[16][570],u_xpb_out[17][570],u_xpb_out[18][570],u_xpb_out[19][570],u_xpb_out[20][570],u_xpb_out[21][570],u_xpb_out[22][570],u_xpb_out[23][570],u_xpb_out[24][570],u_xpb_out[25][570],u_xpb_out[26][570],u_xpb_out[27][570],u_xpb_out[28][570],u_xpb_out[29][570],u_xpb_out[30][570],u_xpb_out[31][570],u_xpb_out[32][570],u_xpb_out[33][570],u_xpb_out[34][570],u_xpb_out[35][570],u_xpb_out[36][570],u_xpb_out[37][570],u_xpb_out[38][570],u_xpb_out[39][570],u_xpb_out[40][570],u_xpb_out[41][570],u_xpb_out[42][570],u_xpb_out[43][570],u_xpb_out[44][570],u_xpb_out[45][570],u_xpb_out[46][570],u_xpb_out[47][570],u_xpb_out[48][570],u_xpb_out[49][570],u_xpb_out[50][570],u_xpb_out[51][570],u_xpb_out[52][570],u_xpb_out[53][570],u_xpb_out[54][570],u_xpb_out[55][570],u_xpb_out[56][570],u_xpb_out[57][570],u_xpb_out[58][570],u_xpb_out[59][570],u_xpb_out[60][570],u_xpb_out[61][570],u_xpb_out[62][570],u_xpb_out[63][570],u_xpb_out[64][570],u_xpb_out[65][570],u_xpb_out[66][570],u_xpb_out[67][570],u_xpb_out[68][570],u_xpb_out[69][570],u_xpb_out[70][570],u_xpb_out[71][570],u_xpb_out[72][570],u_xpb_out[73][570],u_xpb_out[74][570],u_xpb_out[75][570],u_xpb_out[76][570],u_xpb_out[77][570],u_xpb_out[78][570],u_xpb_out[79][570],u_xpb_out[80][570],u_xpb_out[81][570],u_xpb_out[82][570],u_xpb_out[83][570],u_xpb_out[84][570],u_xpb_out[85][570],u_xpb_out[86][570],u_xpb_out[87][570],u_xpb_out[88][570],u_xpb_out[89][570],u_xpb_out[90][570],u_xpb_out[91][570],u_xpb_out[92][570],u_xpb_out[93][570],u_xpb_out[94][570],u_xpb_out[95][570],u_xpb_out[96][570],u_xpb_out[97][570],u_xpb_out[98][570],u_xpb_out[99][570],u_xpb_out[100][570],u_xpb_out[101][570],u_xpb_out[102][570],u_xpb_out[103][570],u_xpb_out[104][570],u_xpb_out[105][570]};

assign col_out_571 = {u_xpb_out[0][571],u_xpb_out[1][571],u_xpb_out[2][571],u_xpb_out[3][571],u_xpb_out[4][571],u_xpb_out[5][571],u_xpb_out[6][571],u_xpb_out[7][571],u_xpb_out[8][571],u_xpb_out[9][571],u_xpb_out[10][571],u_xpb_out[11][571],u_xpb_out[12][571],u_xpb_out[13][571],u_xpb_out[14][571],u_xpb_out[15][571],u_xpb_out[16][571],u_xpb_out[17][571],u_xpb_out[18][571],u_xpb_out[19][571],u_xpb_out[20][571],u_xpb_out[21][571],u_xpb_out[22][571],u_xpb_out[23][571],u_xpb_out[24][571],u_xpb_out[25][571],u_xpb_out[26][571],u_xpb_out[27][571],u_xpb_out[28][571],u_xpb_out[29][571],u_xpb_out[30][571],u_xpb_out[31][571],u_xpb_out[32][571],u_xpb_out[33][571],u_xpb_out[34][571],u_xpb_out[35][571],u_xpb_out[36][571],u_xpb_out[37][571],u_xpb_out[38][571],u_xpb_out[39][571],u_xpb_out[40][571],u_xpb_out[41][571],u_xpb_out[42][571],u_xpb_out[43][571],u_xpb_out[44][571],u_xpb_out[45][571],u_xpb_out[46][571],u_xpb_out[47][571],u_xpb_out[48][571],u_xpb_out[49][571],u_xpb_out[50][571],u_xpb_out[51][571],u_xpb_out[52][571],u_xpb_out[53][571],u_xpb_out[54][571],u_xpb_out[55][571],u_xpb_out[56][571],u_xpb_out[57][571],u_xpb_out[58][571],u_xpb_out[59][571],u_xpb_out[60][571],u_xpb_out[61][571],u_xpb_out[62][571],u_xpb_out[63][571],u_xpb_out[64][571],u_xpb_out[65][571],u_xpb_out[66][571],u_xpb_out[67][571],u_xpb_out[68][571],u_xpb_out[69][571],u_xpb_out[70][571],u_xpb_out[71][571],u_xpb_out[72][571],u_xpb_out[73][571],u_xpb_out[74][571],u_xpb_out[75][571],u_xpb_out[76][571],u_xpb_out[77][571],u_xpb_out[78][571],u_xpb_out[79][571],u_xpb_out[80][571],u_xpb_out[81][571],u_xpb_out[82][571],u_xpb_out[83][571],u_xpb_out[84][571],u_xpb_out[85][571],u_xpb_out[86][571],u_xpb_out[87][571],u_xpb_out[88][571],u_xpb_out[89][571],u_xpb_out[90][571],u_xpb_out[91][571],u_xpb_out[92][571],u_xpb_out[93][571],u_xpb_out[94][571],u_xpb_out[95][571],u_xpb_out[96][571],u_xpb_out[97][571],u_xpb_out[98][571],u_xpb_out[99][571],u_xpb_out[100][571],u_xpb_out[101][571],u_xpb_out[102][571],u_xpb_out[103][571],u_xpb_out[104][571],u_xpb_out[105][571]};

assign col_out_572 = {u_xpb_out[0][572],u_xpb_out[1][572],u_xpb_out[2][572],u_xpb_out[3][572],u_xpb_out[4][572],u_xpb_out[5][572],u_xpb_out[6][572],u_xpb_out[7][572],u_xpb_out[8][572],u_xpb_out[9][572],u_xpb_out[10][572],u_xpb_out[11][572],u_xpb_out[12][572],u_xpb_out[13][572],u_xpb_out[14][572],u_xpb_out[15][572],u_xpb_out[16][572],u_xpb_out[17][572],u_xpb_out[18][572],u_xpb_out[19][572],u_xpb_out[20][572],u_xpb_out[21][572],u_xpb_out[22][572],u_xpb_out[23][572],u_xpb_out[24][572],u_xpb_out[25][572],u_xpb_out[26][572],u_xpb_out[27][572],u_xpb_out[28][572],u_xpb_out[29][572],u_xpb_out[30][572],u_xpb_out[31][572],u_xpb_out[32][572],u_xpb_out[33][572],u_xpb_out[34][572],u_xpb_out[35][572],u_xpb_out[36][572],u_xpb_out[37][572],u_xpb_out[38][572],u_xpb_out[39][572],u_xpb_out[40][572],u_xpb_out[41][572],u_xpb_out[42][572],u_xpb_out[43][572],u_xpb_out[44][572],u_xpb_out[45][572],u_xpb_out[46][572],u_xpb_out[47][572],u_xpb_out[48][572],u_xpb_out[49][572],u_xpb_out[50][572],u_xpb_out[51][572],u_xpb_out[52][572],u_xpb_out[53][572],u_xpb_out[54][572],u_xpb_out[55][572],u_xpb_out[56][572],u_xpb_out[57][572],u_xpb_out[58][572],u_xpb_out[59][572],u_xpb_out[60][572],u_xpb_out[61][572],u_xpb_out[62][572],u_xpb_out[63][572],u_xpb_out[64][572],u_xpb_out[65][572],u_xpb_out[66][572],u_xpb_out[67][572],u_xpb_out[68][572],u_xpb_out[69][572],u_xpb_out[70][572],u_xpb_out[71][572],u_xpb_out[72][572],u_xpb_out[73][572],u_xpb_out[74][572],u_xpb_out[75][572],u_xpb_out[76][572],u_xpb_out[77][572],u_xpb_out[78][572],u_xpb_out[79][572],u_xpb_out[80][572],u_xpb_out[81][572],u_xpb_out[82][572],u_xpb_out[83][572],u_xpb_out[84][572],u_xpb_out[85][572],u_xpb_out[86][572],u_xpb_out[87][572],u_xpb_out[88][572],u_xpb_out[89][572],u_xpb_out[90][572],u_xpb_out[91][572],u_xpb_out[92][572],u_xpb_out[93][572],u_xpb_out[94][572],u_xpb_out[95][572],u_xpb_out[96][572],u_xpb_out[97][572],u_xpb_out[98][572],u_xpb_out[99][572],u_xpb_out[100][572],u_xpb_out[101][572],u_xpb_out[102][572],u_xpb_out[103][572],u_xpb_out[104][572],u_xpb_out[105][572]};

assign col_out_573 = {u_xpb_out[0][573],u_xpb_out[1][573],u_xpb_out[2][573],u_xpb_out[3][573],u_xpb_out[4][573],u_xpb_out[5][573],u_xpb_out[6][573],u_xpb_out[7][573],u_xpb_out[8][573],u_xpb_out[9][573],u_xpb_out[10][573],u_xpb_out[11][573],u_xpb_out[12][573],u_xpb_out[13][573],u_xpb_out[14][573],u_xpb_out[15][573],u_xpb_out[16][573],u_xpb_out[17][573],u_xpb_out[18][573],u_xpb_out[19][573],u_xpb_out[20][573],u_xpb_out[21][573],u_xpb_out[22][573],u_xpb_out[23][573],u_xpb_out[24][573],u_xpb_out[25][573],u_xpb_out[26][573],u_xpb_out[27][573],u_xpb_out[28][573],u_xpb_out[29][573],u_xpb_out[30][573],u_xpb_out[31][573],u_xpb_out[32][573],u_xpb_out[33][573],u_xpb_out[34][573],u_xpb_out[35][573],u_xpb_out[36][573],u_xpb_out[37][573],u_xpb_out[38][573],u_xpb_out[39][573],u_xpb_out[40][573],u_xpb_out[41][573],u_xpb_out[42][573],u_xpb_out[43][573],u_xpb_out[44][573],u_xpb_out[45][573],u_xpb_out[46][573],u_xpb_out[47][573],u_xpb_out[48][573],u_xpb_out[49][573],u_xpb_out[50][573],u_xpb_out[51][573],u_xpb_out[52][573],u_xpb_out[53][573],u_xpb_out[54][573],u_xpb_out[55][573],u_xpb_out[56][573],u_xpb_out[57][573],u_xpb_out[58][573],u_xpb_out[59][573],u_xpb_out[60][573],u_xpb_out[61][573],u_xpb_out[62][573],u_xpb_out[63][573],u_xpb_out[64][573],u_xpb_out[65][573],u_xpb_out[66][573],u_xpb_out[67][573],u_xpb_out[68][573],u_xpb_out[69][573],u_xpb_out[70][573],u_xpb_out[71][573],u_xpb_out[72][573],u_xpb_out[73][573],u_xpb_out[74][573],u_xpb_out[75][573],u_xpb_out[76][573],u_xpb_out[77][573],u_xpb_out[78][573],u_xpb_out[79][573],u_xpb_out[80][573],u_xpb_out[81][573],u_xpb_out[82][573],u_xpb_out[83][573],u_xpb_out[84][573],u_xpb_out[85][573],u_xpb_out[86][573],u_xpb_out[87][573],u_xpb_out[88][573],u_xpb_out[89][573],u_xpb_out[90][573],u_xpb_out[91][573],u_xpb_out[92][573],u_xpb_out[93][573],u_xpb_out[94][573],u_xpb_out[95][573],u_xpb_out[96][573],u_xpb_out[97][573],u_xpb_out[98][573],u_xpb_out[99][573],u_xpb_out[100][573],u_xpb_out[101][573],u_xpb_out[102][573],u_xpb_out[103][573],u_xpb_out[104][573],u_xpb_out[105][573]};

assign col_out_574 = {u_xpb_out[0][574],u_xpb_out[1][574],u_xpb_out[2][574],u_xpb_out[3][574],u_xpb_out[4][574],u_xpb_out[5][574],u_xpb_out[6][574],u_xpb_out[7][574],u_xpb_out[8][574],u_xpb_out[9][574],u_xpb_out[10][574],u_xpb_out[11][574],u_xpb_out[12][574],u_xpb_out[13][574],u_xpb_out[14][574],u_xpb_out[15][574],u_xpb_out[16][574],u_xpb_out[17][574],u_xpb_out[18][574],u_xpb_out[19][574],u_xpb_out[20][574],u_xpb_out[21][574],u_xpb_out[22][574],u_xpb_out[23][574],u_xpb_out[24][574],u_xpb_out[25][574],u_xpb_out[26][574],u_xpb_out[27][574],u_xpb_out[28][574],u_xpb_out[29][574],u_xpb_out[30][574],u_xpb_out[31][574],u_xpb_out[32][574],u_xpb_out[33][574],u_xpb_out[34][574],u_xpb_out[35][574],u_xpb_out[36][574],u_xpb_out[37][574],u_xpb_out[38][574],u_xpb_out[39][574],u_xpb_out[40][574],u_xpb_out[41][574],u_xpb_out[42][574],u_xpb_out[43][574],u_xpb_out[44][574],u_xpb_out[45][574],u_xpb_out[46][574],u_xpb_out[47][574],u_xpb_out[48][574],u_xpb_out[49][574],u_xpb_out[50][574],u_xpb_out[51][574],u_xpb_out[52][574],u_xpb_out[53][574],u_xpb_out[54][574],u_xpb_out[55][574],u_xpb_out[56][574],u_xpb_out[57][574],u_xpb_out[58][574],u_xpb_out[59][574],u_xpb_out[60][574],u_xpb_out[61][574],u_xpb_out[62][574],u_xpb_out[63][574],u_xpb_out[64][574],u_xpb_out[65][574],u_xpb_out[66][574],u_xpb_out[67][574],u_xpb_out[68][574],u_xpb_out[69][574],u_xpb_out[70][574],u_xpb_out[71][574],u_xpb_out[72][574],u_xpb_out[73][574],u_xpb_out[74][574],u_xpb_out[75][574],u_xpb_out[76][574],u_xpb_out[77][574],u_xpb_out[78][574],u_xpb_out[79][574],u_xpb_out[80][574],u_xpb_out[81][574],u_xpb_out[82][574],u_xpb_out[83][574],u_xpb_out[84][574],u_xpb_out[85][574],u_xpb_out[86][574],u_xpb_out[87][574],u_xpb_out[88][574],u_xpb_out[89][574],u_xpb_out[90][574],u_xpb_out[91][574],u_xpb_out[92][574],u_xpb_out[93][574],u_xpb_out[94][574],u_xpb_out[95][574],u_xpb_out[96][574],u_xpb_out[97][574],u_xpb_out[98][574],u_xpb_out[99][574],u_xpb_out[100][574],u_xpb_out[101][574],u_xpb_out[102][574],u_xpb_out[103][574],u_xpb_out[104][574],u_xpb_out[105][574]};

assign col_out_575 = {u_xpb_out[0][575],u_xpb_out[1][575],u_xpb_out[2][575],u_xpb_out[3][575],u_xpb_out[4][575],u_xpb_out[5][575],u_xpb_out[6][575],u_xpb_out[7][575],u_xpb_out[8][575],u_xpb_out[9][575],u_xpb_out[10][575],u_xpb_out[11][575],u_xpb_out[12][575],u_xpb_out[13][575],u_xpb_out[14][575],u_xpb_out[15][575],u_xpb_out[16][575],u_xpb_out[17][575],u_xpb_out[18][575],u_xpb_out[19][575],u_xpb_out[20][575],u_xpb_out[21][575],u_xpb_out[22][575],u_xpb_out[23][575],u_xpb_out[24][575],u_xpb_out[25][575],u_xpb_out[26][575],u_xpb_out[27][575],u_xpb_out[28][575],u_xpb_out[29][575],u_xpb_out[30][575],u_xpb_out[31][575],u_xpb_out[32][575],u_xpb_out[33][575],u_xpb_out[34][575],u_xpb_out[35][575],u_xpb_out[36][575],u_xpb_out[37][575],u_xpb_out[38][575],u_xpb_out[39][575],u_xpb_out[40][575],u_xpb_out[41][575],u_xpb_out[42][575],u_xpb_out[43][575],u_xpb_out[44][575],u_xpb_out[45][575],u_xpb_out[46][575],u_xpb_out[47][575],u_xpb_out[48][575],u_xpb_out[49][575],u_xpb_out[50][575],u_xpb_out[51][575],u_xpb_out[52][575],u_xpb_out[53][575],u_xpb_out[54][575],u_xpb_out[55][575],u_xpb_out[56][575],u_xpb_out[57][575],u_xpb_out[58][575],u_xpb_out[59][575],u_xpb_out[60][575],u_xpb_out[61][575],u_xpb_out[62][575],u_xpb_out[63][575],u_xpb_out[64][575],u_xpb_out[65][575],u_xpb_out[66][575],u_xpb_out[67][575],u_xpb_out[68][575],u_xpb_out[69][575],u_xpb_out[70][575],u_xpb_out[71][575],u_xpb_out[72][575],u_xpb_out[73][575],u_xpb_out[74][575],u_xpb_out[75][575],u_xpb_out[76][575],u_xpb_out[77][575],u_xpb_out[78][575],u_xpb_out[79][575],u_xpb_out[80][575],u_xpb_out[81][575],u_xpb_out[82][575],u_xpb_out[83][575],u_xpb_out[84][575],u_xpb_out[85][575],u_xpb_out[86][575],u_xpb_out[87][575],u_xpb_out[88][575],u_xpb_out[89][575],u_xpb_out[90][575],u_xpb_out[91][575],u_xpb_out[92][575],u_xpb_out[93][575],u_xpb_out[94][575],u_xpb_out[95][575],u_xpb_out[96][575],u_xpb_out[97][575],u_xpb_out[98][575],u_xpb_out[99][575],u_xpb_out[100][575],u_xpb_out[101][575],u_xpb_out[102][575],u_xpb_out[103][575],u_xpb_out[104][575],u_xpb_out[105][575]};

assign col_out_576 = {u_xpb_out[0][576],u_xpb_out[1][576],u_xpb_out[2][576],u_xpb_out[3][576],u_xpb_out[4][576],u_xpb_out[5][576],u_xpb_out[6][576],u_xpb_out[7][576],u_xpb_out[8][576],u_xpb_out[9][576],u_xpb_out[10][576],u_xpb_out[11][576],u_xpb_out[12][576],u_xpb_out[13][576],u_xpb_out[14][576],u_xpb_out[15][576],u_xpb_out[16][576],u_xpb_out[17][576],u_xpb_out[18][576],u_xpb_out[19][576],u_xpb_out[20][576],u_xpb_out[21][576],u_xpb_out[22][576],u_xpb_out[23][576],u_xpb_out[24][576],u_xpb_out[25][576],u_xpb_out[26][576],u_xpb_out[27][576],u_xpb_out[28][576],u_xpb_out[29][576],u_xpb_out[30][576],u_xpb_out[31][576],u_xpb_out[32][576],u_xpb_out[33][576],u_xpb_out[34][576],u_xpb_out[35][576],u_xpb_out[36][576],u_xpb_out[37][576],u_xpb_out[38][576],u_xpb_out[39][576],u_xpb_out[40][576],u_xpb_out[41][576],u_xpb_out[42][576],u_xpb_out[43][576],u_xpb_out[44][576],u_xpb_out[45][576],u_xpb_out[46][576],u_xpb_out[47][576],u_xpb_out[48][576],u_xpb_out[49][576],u_xpb_out[50][576],u_xpb_out[51][576],u_xpb_out[52][576],u_xpb_out[53][576],u_xpb_out[54][576],u_xpb_out[55][576],u_xpb_out[56][576],u_xpb_out[57][576],u_xpb_out[58][576],u_xpb_out[59][576],u_xpb_out[60][576],u_xpb_out[61][576],u_xpb_out[62][576],u_xpb_out[63][576],u_xpb_out[64][576],u_xpb_out[65][576],u_xpb_out[66][576],u_xpb_out[67][576],u_xpb_out[68][576],u_xpb_out[69][576],u_xpb_out[70][576],u_xpb_out[71][576],u_xpb_out[72][576],u_xpb_out[73][576],u_xpb_out[74][576],u_xpb_out[75][576],u_xpb_out[76][576],u_xpb_out[77][576],u_xpb_out[78][576],u_xpb_out[79][576],u_xpb_out[80][576],u_xpb_out[81][576],u_xpb_out[82][576],u_xpb_out[83][576],u_xpb_out[84][576],u_xpb_out[85][576],u_xpb_out[86][576],u_xpb_out[87][576],u_xpb_out[88][576],u_xpb_out[89][576],u_xpb_out[90][576],u_xpb_out[91][576],u_xpb_out[92][576],u_xpb_out[93][576],u_xpb_out[94][576],u_xpb_out[95][576],u_xpb_out[96][576],u_xpb_out[97][576],u_xpb_out[98][576],u_xpb_out[99][576],u_xpb_out[100][576],u_xpb_out[101][576],u_xpb_out[102][576],u_xpb_out[103][576],u_xpb_out[104][576],u_xpb_out[105][576]};

assign col_out_577 = {u_xpb_out[0][577],u_xpb_out[1][577],u_xpb_out[2][577],u_xpb_out[3][577],u_xpb_out[4][577],u_xpb_out[5][577],u_xpb_out[6][577],u_xpb_out[7][577],u_xpb_out[8][577],u_xpb_out[9][577],u_xpb_out[10][577],u_xpb_out[11][577],u_xpb_out[12][577],u_xpb_out[13][577],u_xpb_out[14][577],u_xpb_out[15][577],u_xpb_out[16][577],u_xpb_out[17][577],u_xpb_out[18][577],u_xpb_out[19][577],u_xpb_out[20][577],u_xpb_out[21][577],u_xpb_out[22][577],u_xpb_out[23][577],u_xpb_out[24][577],u_xpb_out[25][577],u_xpb_out[26][577],u_xpb_out[27][577],u_xpb_out[28][577],u_xpb_out[29][577],u_xpb_out[30][577],u_xpb_out[31][577],u_xpb_out[32][577],u_xpb_out[33][577],u_xpb_out[34][577],u_xpb_out[35][577],u_xpb_out[36][577],u_xpb_out[37][577],u_xpb_out[38][577],u_xpb_out[39][577],u_xpb_out[40][577],u_xpb_out[41][577],u_xpb_out[42][577],u_xpb_out[43][577],u_xpb_out[44][577],u_xpb_out[45][577],u_xpb_out[46][577],u_xpb_out[47][577],u_xpb_out[48][577],u_xpb_out[49][577],u_xpb_out[50][577],u_xpb_out[51][577],u_xpb_out[52][577],u_xpb_out[53][577],u_xpb_out[54][577],u_xpb_out[55][577],u_xpb_out[56][577],u_xpb_out[57][577],u_xpb_out[58][577],u_xpb_out[59][577],u_xpb_out[60][577],u_xpb_out[61][577],u_xpb_out[62][577],u_xpb_out[63][577],u_xpb_out[64][577],u_xpb_out[65][577],u_xpb_out[66][577],u_xpb_out[67][577],u_xpb_out[68][577],u_xpb_out[69][577],u_xpb_out[70][577],u_xpb_out[71][577],u_xpb_out[72][577],u_xpb_out[73][577],u_xpb_out[74][577],u_xpb_out[75][577],u_xpb_out[76][577],u_xpb_out[77][577],u_xpb_out[78][577],u_xpb_out[79][577],u_xpb_out[80][577],u_xpb_out[81][577],u_xpb_out[82][577],u_xpb_out[83][577],u_xpb_out[84][577],u_xpb_out[85][577],u_xpb_out[86][577],u_xpb_out[87][577],u_xpb_out[88][577],u_xpb_out[89][577],u_xpb_out[90][577],u_xpb_out[91][577],u_xpb_out[92][577],u_xpb_out[93][577],u_xpb_out[94][577],u_xpb_out[95][577],u_xpb_out[96][577],u_xpb_out[97][577],u_xpb_out[98][577],u_xpb_out[99][577],u_xpb_out[100][577],u_xpb_out[101][577],u_xpb_out[102][577],u_xpb_out[103][577],u_xpb_out[104][577],u_xpb_out[105][577]};

assign col_out_578 = {u_xpb_out[0][578],u_xpb_out[1][578],u_xpb_out[2][578],u_xpb_out[3][578],u_xpb_out[4][578],u_xpb_out[5][578],u_xpb_out[6][578],u_xpb_out[7][578],u_xpb_out[8][578],u_xpb_out[9][578],u_xpb_out[10][578],u_xpb_out[11][578],u_xpb_out[12][578],u_xpb_out[13][578],u_xpb_out[14][578],u_xpb_out[15][578],u_xpb_out[16][578],u_xpb_out[17][578],u_xpb_out[18][578],u_xpb_out[19][578],u_xpb_out[20][578],u_xpb_out[21][578],u_xpb_out[22][578],u_xpb_out[23][578],u_xpb_out[24][578],u_xpb_out[25][578],u_xpb_out[26][578],u_xpb_out[27][578],u_xpb_out[28][578],u_xpb_out[29][578],u_xpb_out[30][578],u_xpb_out[31][578],u_xpb_out[32][578],u_xpb_out[33][578],u_xpb_out[34][578],u_xpb_out[35][578],u_xpb_out[36][578],u_xpb_out[37][578],u_xpb_out[38][578],u_xpb_out[39][578],u_xpb_out[40][578],u_xpb_out[41][578],u_xpb_out[42][578],u_xpb_out[43][578],u_xpb_out[44][578],u_xpb_out[45][578],u_xpb_out[46][578],u_xpb_out[47][578],u_xpb_out[48][578],u_xpb_out[49][578],u_xpb_out[50][578],u_xpb_out[51][578],u_xpb_out[52][578],u_xpb_out[53][578],u_xpb_out[54][578],u_xpb_out[55][578],u_xpb_out[56][578],u_xpb_out[57][578],u_xpb_out[58][578],u_xpb_out[59][578],u_xpb_out[60][578],u_xpb_out[61][578],u_xpb_out[62][578],u_xpb_out[63][578],u_xpb_out[64][578],u_xpb_out[65][578],u_xpb_out[66][578],u_xpb_out[67][578],u_xpb_out[68][578],u_xpb_out[69][578],u_xpb_out[70][578],u_xpb_out[71][578],u_xpb_out[72][578],u_xpb_out[73][578],u_xpb_out[74][578],u_xpb_out[75][578],u_xpb_out[76][578],u_xpb_out[77][578],u_xpb_out[78][578],u_xpb_out[79][578],u_xpb_out[80][578],u_xpb_out[81][578],u_xpb_out[82][578],u_xpb_out[83][578],u_xpb_out[84][578],u_xpb_out[85][578],u_xpb_out[86][578],u_xpb_out[87][578],u_xpb_out[88][578],u_xpb_out[89][578],u_xpb_out[90][578],u_xpb_out[91][578],u_xpb_out[92][578],u_xpb_out[93][578],u_xpb_out[94][578],u_xpb_out[95][578],u_xpb_out[96][578],u_xpb_out[97][578],u_xpb_out[98][578],u_xpb_out[99][578],u_xpb_out[100][578],u_xpb_out[101][578],u_xpb_out[102][578],u_xpb_out[103][578],u_xpb_out[104][578],u_xpb_out[105][578]};

assign col_out_579 = {u_xpb_out[0][579],u_xpb_out[1][579],u_xpb_out[2][579],u_xpb_out[3][579],u_xpb_out[4][579],u_xpb_out[5][579],u_xpb_out[6][579],u_xpb_out[7][579],u_xpb_out[8][579],u_xpb_out[9][579],u_xpb_out[10][579],u_xpb_out[11][579],u_xpb_out[12][579],u_xpb_out[13][579],u_xpb_out[14][579],u_xpb_out[15][579],u_xpb_out[16][579],u_xpb_out[17][579],u_xpb_out[18][579],u_xpb_out[19][579],u_xpb_out[20][579],u_xpb_out[21][579],u_xpb_out[22][579],u_xpb_out[23][579],u_xpb_out[24][579],u_xpb_out[25][579],u_xpb_out[26][579],u_xpb_out[27][579],u_xpb_out[28][579],u_xpb_out[29][579],u_xpb_out[30][579],u_xpb_out[31][579],u_xpb_out[32][579],u_xpb_out[33][579],u_xpb_out[34][579],u_xpb_out[35][579],u_xpb_out[36][579],u_xpb_out[37][579],u_xpb_out[38][579],u_xpb_out[39][579],u_xpb_out[40][579],u_xpb_out[41][579],u_xpb_out[42][579],u_xpb_out[43][579],u_xpb_out[44][579],u_xpb_out[45][579],u_xpb_out[46][579],u_xpb_out[47][579],u_xpb_out[48][579],u_xpb_out[49][579],u_xpb_out[50][579],u_xpb_out[51][579],u_xpb_out[52][579],u_xpb_out[53][579],u_xpb_out[54][579],u_xpb_out[55][579],u_xpb_out[56][579],u_xpb_out[57][579],u_xpb_out[58][579],u_xpb_out[59][579],u_xpb_out[60][579],u_xpb_out[61][579],u_xpb_out[62][579],u_xpb_out[63][579],u_xpb_out[64][579],u_xpb_out[65][579],u_xpb_out[66][579],u_xpb_out[67][579],u_xpb_out[68][579],u_xpb_out[69][579],u_xpb_out[70][579],u_xpb_out[71][579],u_xpb_out[72][579],u_xpb_out[73][579],u_xpb_out[74][579],u_xpb_out[75][579],u_xpb_out[76][579],u_xpb_out[77][579],u_xpb_out[78][579],u_xpb_out[79][579],u_xpb_out[80][579],u_xpb_out[81][579],u_xpb_out[82][579],u_xpb_out[83][579],u_xpb_out[84][579],u_xpb_out[85][579],u_xpb_out[86][579],u_xpb_out[87][579],u_xpb_out[88][579],u_xpb_out[89][579],u_xpb_out[90][579],u_xpb_out[91][579],u_xpb_out[92][579],u_xpb_out[93][579],u_xpb_out[94][579],u_xpb_out[95][579],u_xpb_out[96][579],u_xpb_out[97][579],u_xpb_out[98][579],u_xpb_out[99][579],u_xpb_out[100][579],u_xpb_out[101][579],u_xpb_out[102][579],u_xpb_out[103][579],u_xpb_out[104][579],u_xpb_out[105][579]};

assign col_out_580 = {u_xpb_out[0][580],u_xpb_out[1][580],u_xpb_out[2][580],u_xpb_out[3][580],u_xpb_out[4][580],u_xpb_out[5][580],u_xpb_out[6][580],u_xpb_out[7][580],u_xpb_out[8][580],u_xpb_out[9][580],u_xpb_out[10][580],u_xpb_out[11][580],u_xpb_out[12][580],u_xpb_out[13][580],u_xpb_out[14][580],u_xpb_out[15][580],u_xpb_out[16][580],u_xpb_out[17][580],u_xpb_out[18][580],u_xpb_out[19][580],u_xpb_out[20][580],u_xpb_out[21][580],u_xpb_out[22][580],u_xpb_out[23][580],u_xpb_out[24][580],u_xpb_out[25][580],u_xpb_out[26][580],u_xpb_out[27][580],u_xpb_out[28][580],u_xpb_out[29][580],u_xpb_out[30][580],u_xpb_out[31][580],u_xpb_out[32][580],u_xpb_out[33][580],u_xpb_out[34][580],u_xpb_out[35][580],u_xpb_out[36][580],u_xpb_out[37][580],u_xpb_out[38][580],u_xpb_out[39][580],u_xpb_out[40][580],u_xpb_out[41][580],u_xpb_out[42][580],u_xpb_out[43][580],u_xpb_out[44][580],u_xpb_out[45][580],u_xpb_out[46][580],u_xpb_out[47][580],u_xpb_out[48][580],u_xpb_out[49][580],u_xpb_out[50][580],u_xpb_out[51][580],u_xpb_out[52][580],u_xpb_out[53][580],u_xpb_out[54][580],u_xpb_out[55][580],u_xpb_out[56][580],u_xpb_out[57][580],u_xpb_out[58][580],u_xpb_out[59][580],u_xpb_out[60][580],u_xpb_out[61][580],u_xpb_out[62][580],u_xpb_out[63][580],u_xpb_out[64][580],u_xpb_out[65][580],u_xpb_out[66][580],u_xpb_out[67][580],u_xpb_out[68][580],u_xpb_out[69][580],u_xpb_out[70][580],u_xpb_out[71][580],u_xpb_out[72][580],u_xpb_out[73][580],u_xpb_out[74][580],u_xpb_out[75][580],u_xpb_out[76][580],u_xpb_out[77][580],u_xpb_out[78][580],u_xpb_out[79][580],u_xpb_out[80][580],u_xpb_out[81][580],u_xpb_out[82][580],u_xpb_out[83][580],u_xpb_out[84][580],u_xpb_out[85][580],u_xpb_out[86][580],u_xpb_out[87][580],u_xpb_out[88][580],u_xpb_out[89][580],u_xpb_out[90][580],u_xpb_out[91][580],u_xpb_out[92][580],u_xpb_out[93][580],u_xpb_out[94][580],u_xpb_out[95][580],u_xpb_out[96][580],u_xpb_out[97][580],u_xpb_out[98][580],u_xpb_out[99][580],u_xpb_out[100][580],u_xpb_out[101][580],u_xpb_out[102][580],u_xpb_out[103][580],u_xpb_out[104][580],u_xpb_out[105][580]};

assign col_out_581 = {u_xpb_out[0][581],u_xpb_out[1][581],u_xpb_out[2][581],u_xpb_out[3][581],u_xpb_out[4][581],u_xpb_out[5][581],u_xpb_out[6][581],u_xpb_out[7][581],u_xpb_out[8][581],u_xpb_out[9][581],u_xpb_out[10][581],u_xpb_out[11][581],u_xpb_out[12][581],u_xpb_out[13][581],u_xpb_out[14][581],u_xpb_out[15][581],u_xpb_out[16][581],u_xpb_out[17][581],u_xpb_out[18][581],u_xpb_out[19][581],u_xpb_out[20][581],u_xpb_out[21][581],u_xpb_out[22][581],u_xpb_out[23][581],u_xpb_out[24][581],u_xpb_out[25][581],u_xpb_out[26][581],u_xpb_out[27][581],u_xpb_out[28][581],u_xpb_out[29][581],u_xpb_out[30][581],u_xpb_out[31][581],u_xpb_out[32][581],u_xpb_out[33][581],u_xpb_out[34][581],u_xpb_out[35][581],u_xpb_out[36][581],u_xpb_out[37][581],u_xpb_out[38][581],u_xpb_out[39][581],u_xpb_out[40][581],u_xpb_out[41][581],u_xpb_out[42][581],u_xpb_out[43][581],u_xpb_out[44][581],u_xpb_out[45][581],u_xpb_out[46][581],u_xpb_out[47][581],u_xpb_out[48][581],u_xpb_out[49][581],u_xpb_out[50][581],u_xpb_out[51][581],u_xpb_out[52][581],u_xpb_out[53][581],u_xpb_out[54][581],u_xpb_out[55][581],u_xpb_out[56][581],u_xpb_out[57][581],u_xpb_out[58][581],u_xpb_out[59][581],u_xpb_out[60][581],u_xpb_out[61][581],u_xpb_out[62][581],u_xpb_out[63][581],u_xpb_out[64][581],u_xpb_out[65][581],u_xpb_out[66][581],u_xpb_out[67][581],u_xpb_out[68][581],u_xpb_out[69][581],u_xpb_out[70][581],u_xpb_out[71][581],u_xpb_out[72][581],u_xpb_out[73][581],u_xpb_out[74][581],u_xpb_out[75][581],u_xpb_out[76][581],u_xpb_out[77][581],u_xpb_out[78][581],u_xpb_out[79][581],u_xpb_out[80][581],u_xpb_out[81][581],u_xpb_out[82][581],u_xpb_out[83][581],u_xpb_out[84][581],u_xpb_out[85][581],u_xpb_out[86][581],u_xpb_out[87][581],u_xpb_out[88][581],u_xpb_out[89][581],u_xpb_out[90][581],u_xpb_out[91][581],u_xpb_out[92][581],u_xpb_out[93][581],u_xpb_out[94][581],u_xpb_out[95][581],u_xpb_out[96][581],u_xpb_out[97][581],u_xpb_out[98][581],u_xpb_out[99][581],u_xpb_out[100][581],u_xpb_out[101][581],u_xpb_out[102][581],u_xpb_out[103][581],u_xpb_out[104][581],u_xpb_out[105][581]};

assign col_out_582 = {u_xpb_out[0][582],u_xpb_out[1][582],u_xpb_out[2][582],u_xpb_out[3][582],u_xpb_out[4][582],u_xpb_out[5][582],u_xpb_out[6][582],u_xpb_out[7][582],u_xpb_out[8][582],u_xpb_out[9][582],u_xpb_out[10][582],u_xpb_out[11][582],u_xpb_out[12][582],u_xpb_out[13][582],u_xpb_out[14][582],u_xpb_out[15][582],u_xpb_out[16][582],u_xpb_out[17][582],u_xpb_out[18][582],u_xpb_out[19][582],u_xpb_out[20][582],u_xpb_out[21][582],u_xpb_out[22][582],u_xpb_out[23][582],u_xpb_out[24][582],u_xpb_out[25][582],u_xpb_out[26][582],u_xpb_out[27][582],u_xpb_out[28][582],u_xpb_out[29][582],u_xpb_out[30][582],u_xpb_out[31][582],u_xpb_out[32][582],u_xpb_out[33][582],u_xpb_out[34][582],u_xpb_out[35][582],u_xpb_out[36][582],u_xpb_out[37][582],u_xpb_out[38][582],u_xpb_out[39][582],u_xpb_out[40][582],u_xpb_out[41][582],u_xpb_out[42][582],u_xpb_out[43][582],u_xpb_out[44][582],u_xpb_out[45][582],u_xpb_out[46][582],u_xpb_out[47][582],u_xpb_out[48][582],u_xpb_out[49][582],u_xpb_out[50][582],u_xpb_out[51][582],u_xpb_out[52][582],u_xpb_out[53][582],u_xpb_out[54][582],u_xpb_out[55][582],u_xpb_out[56][582],u_xpb_out[57][582],u_xpb_out[58][582],u_xpb_out[59][582],u_xpb_out[60][582],u_xpb_out[61][582],u_xpb_out[62][582],u_xpb_out[63][582],u_xpb_out[64][582],u_xpb_out[65][582],u_xpb_out[66][582],u_xpb_out[67][582],u_xpb_out[68][582],u_xpb_out[69][582],u_xpb_out[70][582],u_xpb_out[71][582],u_xpb_out[72][582],u_xpb_out[73][582],u_xpb_out[74][582],u_xpb_out[75][582],u_xpb_out[76][582],u_xpb_out[77][582],u_xpb_out[78][582],u_xpb_out[79][582],u_xpb_out[80][582],u_xpb_out[81][582],u_xpb_out[82][582],u_xpb_out[83][582],u_xpb_out[84][582],u_xpb_out[85][582],u_xpb_out[86][582],u_xpb_out[87][582],u_xpb_out[88][582],u_xpb_out[89][582],u_xpb_out[90][582],u_xpb_out[91][582],u_xpb_out[92][582],u_xpb_out[93][582],u_xpb_out[94][582],u_xpb_out[95][582],u_xpb_out[96][582],u_xpb_out[97][582],u_xpb_out[98][582],u_xpb_out[99][582],u_xpb_out[100][582],u_xpb_out[101][582],u_xpb_out[102][582],u_xpb_out[103][582],u_xpb_out[104][582],u_xpb_out[105][582]};

assign col_out_583 = {u_xpb_out[0][583],u_xpb_out[1][583],u_xpb_out[2][583],u_xpb_out[3][583],u_xpb_out[4][583],u_xpb_out[5][583],u_xpb_out[6][583],u_xpb_out[7][583],u_xpb_out[8][583],u_xpb_out[9][583],u_xpb_out[10][583],u_xpb_out[11][583],u_xpb_out[12][583],u_xpb_out[13][583],u_xpb_out[14][583],u_xpb_out[15][583],u_xpb_out[16][583],u_xpb_out[17][583],u_xpb_out[18][583],u_xpb_out[19][583],u_xpb_out[20][583],u_xpb_out[21][583],u_xpb_out[22][583],u_xpb_out[23][583],u_xpb_out[24][583],u_xpb_out[25][583],u_xpb_out[26][583],u_xpb_out[27][583],u_xpb_out[28][583],u_xpb_out[29][583],u_xpb_out[30][583],u_xpb_out[31][583],u_xpb_out[32][583],u_xpb_out[33][583],u_xpb_out[34][583],u_xpb_out[35][583],u_xpb_out[36][583],u_xpb_out[37][583],u_xpb_out[38][583],u_xpb_out[39][583],u_xpb_out[40][583],u_xpb_out[41][583],u_xpb_out[42][583],u_xpb_out[43][583],u_xpb_out[44][583],u_xpb_out[45][583],u_xpb_out[46][583],u_xpb_out[47][583],u_xpb_out[48][583],u_xpb_out[49][583],u_xpb_out[50][583],u_xpb_out[51][583],u_xpb_out[52][583],u_xpb_out[53][583],u_xpb_out[54][583],u_xpb_out[55][583],u_xpb_out[56][583],u_xpb_out[57][583],u_xpb_out[58][583],u_xpb_out[59][583],u_xpb_out[60][583],u_xpb_out[61][583],u_xpb_out[62][583],u_xpb_out[63][583],u_xpb_out[64][583],u_xpb_out[65][583],u_xpb_out[66][583],u_xpb_out[67][583],u_xpb_out[68][583],u_xpb_out[69][583],u_xpb_out[70][583],u_xpb_out[71][583],u_xpb_out[72][583],u_xpb_out[73][583],u_xpb_out[74][583],u_xpb_out[75][583],u_xpb_out[76][583],u_xpb_out[77][583],u_xpb_out[78][583],u_xpb_out[79][583],u_xpb_out[80][583],u_xpb_out[81][583],u_xpb_out[82][583],u_xpb_out[83][583],u_xpb_out[84][583],u_xpb_out[85][583],u_xpb_out[86][583],u_xpb_out[87][583],u_xpb_out[88][583],u_xpb_out[89][583],u_xpb_out[90][583],u_xpb_out[91][583],u_xpb_out[92][583],u_xpb_out[93][583],u_xpb_out[94][583],u_xpb_out[95][583],u_xpb_out[96][583],u_xpb_out[97][583],u_xpb_out[98][583],u_xpb_out[99][583],u_xpb_out[100][583],u_xpb_out[101][583],u_xpb_out[102][583],u_xpb_out[103][583],u_xpb_out[104][583],u_xpb_out[105][583]};

assign col_out_584 = {u_xpb_out[0][584],u_xpb_out[1][584],u_xpb_out[2][584],u_xpb_out[3][584],u_xpb_out[4][584],u_xpb_out[5][584],u_xpb_out[6][584],u_xpb_out[7][584],u_xpb_out[8][584],u_xpb_out[9][584],u_xpb_out[10][584],u_xpb_out[11][584],u_xpb_out[12][584],u_xpb_out[13][584],u_xpb_out[14][584],u_xpb_out[15][584],u_xpb_out[16][584],u_xpb_out[17][584],u_xpb_out[18][584],u_xpb_out[19][584],u_xpb_out[20][584],u_xpb_out[21][584],u_xpb_out[22][584],u_xpb_out[23][584],u_xpb_out[24][584],u_xpb_out[25][584],u_xpb_out[26][584],u_xpb_out[27][584],u_xpb_out[28][584],u_xpb_out[29][584],u_xpb_out[30][584],u_xpb_out[31][584],u_xpb_out[32][584],u_xpb_out[33][584],u_xpb_out[34][584],u_xpb_out[35][584],u_xpb_out[36][584],u_xpb_out[37][584],u_xpb_out[38][584],u_xpb_out[39][584],u_xpb_out[40][584],u_xpb_out[41][584],u_xpb_out[42][584],u_xpb_out[43][584],u_xpb_out[44][584],u_xpb_out[45][584],u_xpb_out[46][584],u_xpb_out[47][584],u_xpb_out[48][584],u_xpb_out[49][584],u_xpb_out[50][584],u_xpb_out[51][584],u_xpb_out[52][584],u_xpb_out[53][584],u_xpb_out[54][584],u_xpb_out[55][584],u_xpb_out[56][584],u_xpb_out[57][584],u_xpb_out[58][584],u_xpb_out[59][584],u_xpb_out[60][584],u_xpb_out[61][584],u_xpb_out[62][584],u_xpb_out[63][584],u_xpb_out[64][584],u_xpb_out[65][584],u_xpb_out[66][584],u_xpb_out[67][584],u_xpb_out[68][584],u_xpb_out[69][584],u_xpb_out[70][584],u_xpb_out[71][584],u_xpb_out[72][584],u_xpb_out[73][584],u_xpb_out[74][584],u_xpb_out[75][584],u_xpb_out[76][584],u_xpb_out[77][584],u_xpb_out[78][584],u_xpb_out[79][584],u_xpb_out[80][584],u_xpb_out[81][584],u_xpb_out[82][584],u_xpb_out[83][584],u_xpb_out[84][584],u_xpb_out[85][584],u_xpb_out[86][584],u_xpb_out[87][584],u_xpb_out[88][584],u_xpb_out[89][584],u_xpb_out[90][584],u_xpb_out[91][584],u_xpb_out[92][584],u_xpb_out[93][584],u_xpb_out[94][584],u_xpb_out[95][584],u_xpb_out[96][584],u_xpb_out[97][584],u_xpb_out[98][584],u_xpb_out[99][584],u_xpb_out[100][584],u_xpb_out[101][584],u_xpb_out[102][584],u_xpb_out[103][584],u_xpb_out[104][584],u_xpb_out[105][584]};

assign col_out_585 = {u_xpb_out[0][585],u_xpb_out[1][585],u_xpb_out[2][585],u_xpb_out[3][585],u_xpb_out[4][585],u_xpb_out[5][585],u_xpb_out[6][585],u_xpb_out[7][585],u_xpb_out[8][585],u_xpb_out[9][585],u_xpb_out[10][585],u_xpb_out[11][585],u_xpb_out[12][585],u_xpb_out[13][585],u_xpb_out[14][585],u_xpb_out[15][585],u_xpb_out[16][585],u_xpb_out[17][585],u_xpb_out[18][585],u_xpb_out[19][585],u_xpb_out[20][585],u_xpb_out[21][585],u_xpb_out[22][585],u_xpb_out[23][585],u_xpb_out[24][585],u_xpb_out[25][585],u_xpb_out[26][585],u_xpb_out[27][585],u_xpb_out[28][585],u_xpb_out[29][585],u_xpb_out[30][585],u_xpb_out[31][585],u_xpb_out[32][585],u_xpb_out[33][585],u_xpb_out[34][585],u_xpb_out[35][585],u_xpb_out[36][585],u_xpb_out[37][585],u_xpb_out[38][585],u_xpb_out[39][585],u_xpb_out[40][585],u_xpb_out[41][585],u_xpb_out[42][585],u_xpb_out[43][585],u_xpb_out[44][585],u_xpb_out[45][585],u_xpb_out[46][585],u_xpb_out[47][585],u_xpb_out[48][585],u_xpb_out[49][585],u_xpb_out[50][585],u_xpb_out[51][585],u_xpb_out[52][585],u_xpb_out[53][585],u_xpb_out[54][585],u_xpb_out[55][585],u_xpb_out[56][585],u_xpb_out[57][585],u_xpb_out[58][585],u_xpb_out[59][585],u_xpb_out[60][585],u_xpb_out[61][585],u_xpb_out[62][585],u_xpb_out[63][585],u_xpb_out[64][585],u_xpb_out[65][585],u_xpb_out[66][585],u_xpb_out[67][585],u_xpb_out[68][585],u_xpb_out[69][585],u_xpb_out[70][585],u_xpb_out[71][585],u_xpb_out[72][585],u_xpb_out[73][585],u_xpb_out[74][585],u_xpb_out[75][585],u_xpb_out[76][585],u_xpb_out[77][585],u_xpb_out[78][585],u_xpb_out[79][585],u_xpb_out[80][585],u_xpb_out[81][585],u_xpb_out[82][585],u_xpb_out[83][585],u_xpb_out[84][585],u_xpb_out[85][585],u_xpb_out[86][585],u_xpb_out[87][585],u_xpb_out[88][585],u_xpb_out[89][585],u_xpb_out[90][585],u_xpb_out[91][585],u_xpb_out[92][585],u_xpb_out[93][585],u_xpb_out[94][585],u_xpb_out[95][585],u_xpb_out[96][585],u_xpb_out[97][585],u_xpb_out[98][585],u_xpb_out[99][585],u_xpb_out[100][585],u_xpb_out[101][585],u_xpb_out[102][585],u_xpb_out[103][585],u_xpb_out[104][585],u_xpb_out[105][585]};

assign col_out_586 = {u_xpb_out[0][586],u_xpb_out[1][586],u_xpb_out[2][586],u_xpb_out[3][586],u_xpb_out[4][586],u_xpb_out[5][586],u_xpb_out[6][586],u_xpb_out[7][586],u_xpb_out[8][586],u_xpb_out[9][586],u_xpb_out[10][586],u_xpb_out[11][586],u_xpb_out[12][586],u_xpb_out[13][586],u_xpb_out[14][586],u_xpb_out[15][586],u_xpb_out[16][586],u_xpb_out[17][586],u_xpb_out[18][586],u_xpb_out[19][586],u_xpb_out[20][586],u_xpb_out[21][586],u_xpb_out[22][586],u_xpb_out[23][586],u_xpb_out[24][586],u_xpb_out[25][586],u_xpb_out[26][586],u_xpb_out[27][586],u_xpb_out[28][586],u_xpb_out[29][586],u_xpb_out[30][586],u_xpb_out[31][586],u_xpb_out[32][586],u_xpb_out[33][586],u_xpb_out[34][586],u_xpb_out[35][586],u_xpb_out[36][586],u_xpb_out[37][586],u_xpb_out[38][586],u_xpb_out[39][586],u_xpb_out[40][586],u_xpb_out[41][586],u_xpb_out[42][586],u_xpb_out[43][586],u_xpb_out[44][586],u_xpb_out[45][586],u_xpb_out[46][586],u_xpb_out[47][586],u_xpb_out[48][586],u_xpb_out[49][586],u_xpb_out[50][586],u_xpb_out[51][586],u_xpb_out[52][586],u_xpb_out[53][586],u_xpb_out[54][586],u_xpb_out[55][586],u_xpb_out[56][586],u_xpb_out[57][586],u_xpb_out[58][586],u_xpb_out[59][586],u_xpb_out[60][586],u_xpb_out[61][586],u_xpb_out[62][586],u_xpb_out[63][586],u_xpb_out[64][586],u_xpb_out[65][586],u_xpb_out[66][586],u_xpb_out[67][586],u_xpb_out[68][586],u_xpb_out[69][586],u_xpb_out[70][586],u_xpb_out[71][586],u_xpb_out[72][586],u_xpb_out[73][586],u_xpb_out[74][586],u_xpb_out[75][586],u_xpb_out[76][586],u_xpb_out[77][586],u_xpb_out[78][586],u_xpb_out[79][586],u_xpb_out[80][586],u_xpb_out[81][586],u_xpb_out[82][586],u_xpb_out[83][586],u_xpb_out[84][586],u_xpb_out[85][586],u_xpb_out[86][586],u_xpb_out[87][586],u_xpb_out[88][586],u_xpb_out[89][586],u_xpb_out[90][586],u_xpb_out[91][586],u_xpb_out[92][586],u_xpb_out[93][586],u_xpb_out[94][586],u_xpb_out[95][586],u_xpb_out[96][586],u_xpb_out[97][586],u_xpb_out[98][586],u_xpb_out[99][586],u_xpb_out[100][586],u_xpb_out[101][586],u_xpb_out[102][586],u_xpb_out[103][586],u_xpb_out[104][586],u_xpb_out[105][586]};

assign col_out_587 = {u_xpb_out[0][587],u_xpb_out[1][587],u_xpb_out[2][587],u_xpb_out[3][587],u_xpb_out[4][587],u_xpb_out[5][587],u_xpb_out[6][587],u_xpb_out[7][587],u_xpb_out[8][587],u_xpb_out[9][587],u_xpb_out[10][587],u_xpb_out[11][587],u_xpb_out[12][587],u_xpb_out[13][587],u_xpb_out[14][587],u_xpb_out[15][587],u_xpb_out[16][587],u_xpb_out[17][587],u_xpb_out[18][587],u_xpb_out[19][587],u_xpb_out[20][587],u_xpb_out[21][587],u_xpb_out[22][587],u_xpb_out[23][587],u_xpb_out[24][587],u_xpb_out[25][587],u_xpb_out[26][587],u_xpb_out[27][587],u_xpb_out[28][587],u_xpb_out[29][587],u_xpb_out[30][587],u_xpb_out[31][587],u_xpb_out[32][587],u_xpb_out[33][587],u_xpb_out[34][587],u_xpb_out[35][587],u_xpb_out[36][587],u_xpb_out[37][587],u_xpb_out[38][587],u_xpb_out[39][587],u_xpb_out[40][587],u_xpb_out[41][587],u_xpb_out[42][587],u_xpb_out[43][587],u_xpb_out[44][587],u_xpb_out[45][587],u_xpb_out[46][587],u_xpb_out[47][587],u_xpb_out[48][587],u_xpb_out[49][587],u_xpb_out[50][587],u_xpb_out[51][587],u_xpb_out[52][587],u_xpb_out[53][587],u_xpb_out[54][587],u_xpb_out[55][587],u_xpb_out[56][587],u_xpb_out[57][587],u_xpb_out[58][587],u_xpb_out[59][587],u_xpb_out[60][587],u_xpb_out[61][587],u_xpb_out[62][587],u_xpb_out[63][587],u_xpb_out[64][587],u_xpb_out[65][587],u_xpb_out[66][587],u_xpb_out[67][587],u_xpb_out[68][587],u_xpb_out[69][587],u_xpb_out[70][587],u_xpb_out[71][587],u_xpb_out[72][587],u_xpb_out[73][587],u_xpb_out[74][587],u_xpb_out[75][587],u_xpb_out[76][587],u_xpb_out[77][587],u_xpb_out[78][587],u_xpb_out[79][587],u_xpb_out[80][587],u_xpb_out[81][587],u_xpb_out[82][587],u_xpb_out[83][587],u_xpb_out[84][587],u_xpb_out[85][587],u_xpb_out[86][587],u_xpb_out[87][587],u_xpb_out[88][587],u_xpb_out[89][587],u_xpb_out[90][587],u_xpb_out[91][587],u_xpb_out[92][587],u_xpb_out[93][587],u_xpb_out[94][587],u_xpb_out[95][587],u_xpb_out[96][587],u_xpb_out[97][587],u_xpb_out[98][587],u_xpb_out[99][587],u_xpb_out[100][587],u_xpb_out[101][587],u_xpb_out[102][587],u_xpb_out[103][587],u_xpb_out[104][587],u_xpb_out[105][587]};

assign col_out_588 = {u_xpb_out[0][588],u_xpb_out[1][588],u_xpb_out[2][588],u_xpb_out[3][588],u_xpb_out[4][588],u_xpb_out[5][588],u_xpb_out[6][588],u_xpb_out[7][588],u_xpb_out[8][588],u_xpb_out[9][588],u_xpb_out[10][588],u_xpb_out[11][588],u_xpb_out[12][588],u_xpb_out[13][588],u_xpb_out[14][588],u_xpb_out[15][588],u_xpb_out[16][588],u_xpb_out[17][588],u_xpb_out[18][588],u_xpb_out[19][588],u_xpb_out[20][588],u_xpb_out[21][588],u_xpb_out[22][588],u_xpb_out[23][588],u_xpb_out[24][588],u_xpb_out[25][588],u_xpb_out[26][588],u_xpb_out[27][588],u_xpb_out[28][588],u_xpb_out[29][588],u_xpb_out[30][588],u_xpb_out[31][588],u_xpb_out[32][588],u_xpb_out[33][588],u_xpb_out[34][588],u_xpb_out[35][588],u_xpb_out[36][588],u_xpb_out[37][588],u_xpb_out[38][588],u_xpb_out[39][588],u_xpb_out[40][588],u_xpb_out[41][588],u_xpb_out[42][588],u_xpb_out[43][588],u_xpb_out[44][588],u_xpb_out[45][588],u_xpb_out[46][588],u_xpb_out[47][588],u_xpb_out[48][588],u_xpb_out[49][588],u_xpb_out[50][588],u_xpb_out[51][588],u_xpb_out[52][588],u_xpb_out[53][588],u_xpb_out[54][588],u_xpb_out[55][588],u_xpb_out[56][588],u_xpb_out[57][588],u_xpb_out[58][588],u_xpb_out[59][588],u_xpb_out[60][588],u_xpb_out[61][588],u_xpb_out[62][588],u_xpb_out[63][588],u_xpb_out[64][588],u_xpb_out[65][588],u_xpb_out[66][588],u_xpb_out[67][588],u_xpb_out[68][588],u_xpb_out[69][588],u_xpb_out[70][588],u_xpb_out[71][588],u_xpb_out[72][588],u_xpb_out[73][588],u_xpb_out[74][588],u_xpb_out[75][588],u_xpb_out[76][588],u_xpb_out[77][588],u_xpb_out[78][588],u_xpb_out[79][588],u_xpb_out[80][588],u_xpb_out[81][588],u_xpb_out[82][588],u_xpb_out[83][588],u_xpb_out[84][588],u_xpb_out[85][588],u_xpb_out[86][588],u_xpb_out[87][588],u_xpb_out[88][588],u_xpb_out[89][588],u_xpb_out[90][588],u_xpb_out[91][588],u_xpb_out[92][588],u_xpb_out[93][588],u_xpb_out[94][588],u_xpb_out[95][588],u_xpb_out[96][588],u_xpb_out[97][588],u_xpb_out[98][588],u_xpb_out[99][588],u_xpb_out[100][588],u_xpb_out[101][588],u_xpb_out[102][588],u_xpb_out[103][588],u_xpb_out[104][588],u_xpb_out[105][588]};

assign col_out_589 = {u_xpb_out[0][589],u_xpb_out[1][589],u_xpb_out[2][589],u_xpb_out[3][589],u_xpb_out[4][589],u_xpb_out[5][589],u_xpb_out[6][589],u_xpb_out[7][589],u_xpb_out[8][589],u_xpb_out[9][589],u_xpb_out[10][589],u_xpb_out[11][589],u_xpb_out[12][589],u_xpb_out[13][589],u_xpb_out[14][589],u_xpb_out[15][589],u_xpb_out[16][589],u_xpb_out[17][589],u_xpb_out[18][589],u_xpb_out[19][589],u_xpb_out[20][589],u_xpb_out[21][589],u_xpb_out[22][589],u_xpb_out[23][589],u_xpb_out[24][589],u_xpb_out[25][589],u_xpb_out[26][589],u_xpb_out[27][589],u_xpb_out[28][589],u_xpb_out[29][589],u_xpb_out[30][589],u_xpb_out[31][589],u_xpb_out[32][589],u_xpb_out[33][589],u_xpb_out[34][589],u_xpb_out[35][589],u_xpb_out[36][589],u_xpb_out[37][589],u_xpb_out[38][589],u_xpb_out[39][589],u_xpb_out[40][589],u_xpb_out[41][589],u_xpb_out[42][589],u_xpb_out[43][589],u_xpb_out[44][589],u_xpb_out[45][589],u_xpb_out[46][589],u_xpb_out[47][589],u_xpb_out[48][589],u_xpb_out[49][589],u_xpb_out[50][589],u_xpb_out[51][589],u_xpb_out[52][589],u_xpb_out[53][589],u_xpb_out[54][589],u_xpb_out[55][589],u_xpb_out[56][589],u_xpb_out[57][589],u_xpb_out[58][589],u_xpb_out[59][589],u_xpb_out[60][589],u_xpb_out[61][589],u_xpb_out[62][589],u_xpb_out[63][589],u_xpb_out[64][589],u_xpb_out[65][589],u_xpb_out[66][589],u_xpb_out[67][589],u_xpb_out[68][589],u_xpb_out[69][589],u_xpb_out[70][589],u_xpb_out[71][589],u_xpb_out[72][589],u_xpb_out[73][589],u_xpb_out[74][589],u_xpb_out[75][589],u_xpb_out[76][589],u_xpb_out[77][589],u_xpb_out[78][589],u_xpb_out[79][589],u_xpb_out[80][589],u_xpb_out[81][589],u_xpb_out[82][589],u_xpb_out[83][589],u_xpb_out[84][589],u_xpb_out[85][589],u_xpb_out[86][589],u_xpb_out[87][589],u_xpb_out[88][589],u_xpb_out[89][589],u_xpb_out[90][589],u_xpb_out[91][589],u_xpb_out[92][589],u_xpb_out[93][589],u_xpb_out[94][589],u_xpb_out[95][589],u_xpb_out[96][589],u_xpb_out[97][589],u_xpb_out[98][589],u_xpb_out[99][589],u_xpb_out[100][589],u_xpb_out[101][589],u_xpb_out[102][589],u_xpb_out[103][589],u_xpb_out[104][589],u_xpb_out[105][589]};

assign col_out_590 = {u_xpb_out[0][590],u_xpb_out[1][590],u_xpb_out[2][590],u_xpb_out[3][590],u_xpb_out[4][590],u_xpb_out[5][590],u_xpb_out[6][590],u_xpb_out[7][590],u_xpb_out[8][590],u_xpb_out[9][590],u_xpb_out[10][590],u_xpb_out[11][590],u_xpb_out[12][590],u_xpb_out[13][590],u_xpb_out[14][590],u_xpb_out[15][590],u_xpb_out[16][590],u_xpb_out[17][590],u_xpb_out[18][590],u_xpb_out[19][590],u_xpb_out[20][590],u_xpb_out[21][590],u_xpb_out[22][590],u_xpb_out[23][590],u_xpb_out[24][590],u_xpb_out[25][590],u_xpb_out[26][590],u_xpb_out[27][590],u_xpb_out[28][590],u_xpb_out[29][590],u_xpb_out[30][590],u_xpb_out[31][590],u_xpb_out[32][590],u_xpb_out[33][590],u_xpb_out[34][590],u_xpb_out[35][590],u_xpb_out[36][590],u_xpb_out[37][590],u_xpb_out[38][590],u_xpb_out[39][590],u_xpb_out[40][590],u_xpb_out[41][590],u_xpb_out[42][590],u_xpb_out[43][590],u_xpb_out[44][590],u_xpb_out[45][590],u_xpb_out[46][590],u_xpb_out[47][590],u_xpb_out[48][590],u_xpb_out[49][590],u_xpb_out[50][590],u_xpb_out[51][590],u_xpb_out[52][590],u_xpb_out[53][590],u_xpb_out[54][590],u_xpb_out[55][590],u_xpb_out[56][590],u_xpb_out[57][590],u_xpb_out[58][590],u_xpb_out[59][590],u_xpb_out[60][590],u_xpb_out[61][590],u_xpb_out[62][590],u_xpb_out[63][590],u_xpb_out[64][590],u_xpb_out[65][590],u_xpb_out[66][590],u_xpb_out[67][590],u_xpb_out[68][590],u_xpb_out[69][590],u_xpb_out[70][590],u_xpb_out[71][590],u_xpb_out[72][590],u_xpb_out[73][590],u_xpb_out[74][590],u_xpb_out[75][590],u_xpb_out[76][590],u_xpb_out[77][590],u_xpb_out[78][590],u_xpb_out[79][590],u_xpb_out[80][590],u_xpb_out[81][590],u_xpb_out[82][590],u_xpb_out[83][590],u_xpb_out[84][590],u_xpb_out[85][590],u_xpb_out[86][590],u_xpb_out[87][590],u_xpb_out[88][590],u_xpb_out[89][590],u_xpb_out[90][590],u_xpb_out[91][590],u_xpb_out[92][590],u_xpb_out[93][590],u_xpb_out[94][590],u_xpb_out[95][590],u_xpb_out[96][590],u_xpb_out[97][590],u_xpb_out[98][590],u_xpb_out[99][590],u_xpb_out[100][590],u_xpb_out[101][590],u_xpb_out[102][590],u_xpb_out[103][590],u_xpb_out[104][590],u_xpb_out[105][590]};

assign col_out_591 = {u_xpb_out[0][591],u_xpb_out[1][591],u_xpb_out[2][591],u_xpb_out[3][591],u_xpb_out[4][591],u_xpb_out[5][591],u_xpb_out[6][591],u_xpb_out[7][591],u_xpb_out[8][591],u_xpb_out[9][591],u_xpb_out[10][591],u_xpb_out[11][591],u_xpb_out[12][591],u_xpb_out[13][591],u_xpb_out[14][591],u_xpb_out[15][591],u_xpb_out[16][591],u_xpb_out[17][591],u_xpb_out[18][591],u_xpb_out[19][591],u_xpb_out[20][591],u_xpb_out[21][591],u_xpb_out[22][591],u_xpb_out[23][591],u_xpb_out[24][591],u_xpb_out[25][591],u_xpb_out[26][591],u_xpb_out[27][591],u_xpb_out[28][591],u_xpb_out[29][591],u_xpb_out[30][591],u_xpb_out[31][591],u_xpb_out[32][591],u_xpb_out[33][591],u_xpb_out[34][591],u_xpb_out[35][591],u_xpb_out[36][591],u_xpb_out[37][591],u_xpb_out[38][591],u_xpb_out[39][591],u_xpb_out[40][591],u_xpb_out[41][591],u_xpb_out[42][591],u_xpb_out[43][591],u_xpb_out[44][591],u_xpb_out[45][591],u_xpb_out[46][591],u_xpb_out[47][591],u_xpb_out[48][591],u_xpb_out[49][591],u_xpb_out[50][591],u_xpb_out[51][591],u_xpb_out[52][591],u_xpb_out[53][591],u_xpb_out[54][591],u_xpb_out[55][591],u_xpb_out[56][591],u_xpb_out[57][591],u_xpb_out[58][591],u_xpb_out[59][591],u_xpb_out[60][591],u_xpb_out[61][591],u_xpb_out[62][591],u_xpb_out[63][591],u_xpb_out[64][591],u_xpb_out[65][591],u_xpb_out[66][591],u_xpb_out[67][591],u_xpb_out[68][591],u_xpb_out[69][591],u_xpb_out[70][591],u_xpb_out[71][591],u_xpb_out[72][591],u_xpb_out[73][591],u_xpb_out[74][591],u_xpb_out[75][591],u_xpb_out[76][591],u_xpb_out[77][591],u_xpb_out[78][591],u_xpb_out[79][591],u_xpb_out[80][591],u_xpb_out[81][591],u_xpb_out[82][591],u_xpb_out[83][591],u_xpb_out[84][591],u_xpb_out[85][591],u_xpb_out[86][591],u_xpb_out[87][591],u_xpb_out[88][591],u_xpb_out[89][591],u_xpb_out[90][591],u_xpb_out[91][591],u_xpb_out[92][591],u_xpb_out[93][591],u_xpb_out[94][591],u_xpb_out[95][591],u_xpb_out[96][591],u_xpb_out[97][591],u_xpb_out[98][591],u_xpb_out[99][591],u_xpb_out[100][591],u_xpb_out[101][591],u_xpb_out[102][591],u_xpb_out[103][591],u_xpb_out[104][591],u_xpb_out[105][591]};

assign col_out_592 = {u_xpb_out[0][592],u_xpb_out[1][592],u_xpb_out[2][592],u_xpb_out[3][592],u_xpb_out[4][592],u_xpb_out[5][592],u_xpb_out[6][592],u_xpb_out[7][592],u_xpb_out[8][592],u_xpb_out[9][592],u_xpb_out[10][592],u_xpb_out[11][592],u_xpb_out[12][592],u_xpb_out[13][592],u_xpb_out[14][592],u_xpb_out[15][592],u_xpb_out[16][592],u_xpb_out[17][592],u_xpb_out[18][592],u_xpb_out[19][592],u_xpb_out[20][592],u_xpb_out[21][592],u_xpb_out[22][592],u_xpb_out[23][592],u_xpb_out[24][592],u_xpb_out[25][592],u_xpb_out[26][592],u_xpb_out[27][592],u_xpb_out[28][592],u_xpb_out[29][592],u_xpb_out[30][592],u_xpb_out[31][592],u_xpb_out[32][592],u_xpb_out[33][592],u_xpb_out[34][592],u_xpb_out[35][592],u_xpb_out[36][592],u_xpb_out[37][592],u_xpb_out[38][592],u_xpb_out[39][592],u_xpb_out[40][592],u_xpb_out[41][592],u_xpb_out[42][592],u_xpb_out[43][592],u_xpb_out[44][592],u_xpb_out[45][592],u_xpb_out[46][592],u_xpb_out[47][592],u_xpb_out[48][592],u_xpb_out[49][592],u_xpb_out[50][592],u_xpb_out[51][592],u_xpb_out[52][592],u_xpb_out[53][592],u_xpb_out[54][592],u_xpb_out[55][592],u_xpb_out[56][592],u_xpb_out[57][592],u_xpb_out[58][592],u_xpb_out[59][592],u_xpb_out[60][592],u_xpb_out[61][592],u_xpb_out[62][592],u_xpb_out[63][592],u_xpb_out[64][592],u_xpb_out[65][592],u_xpb_out[66][592],u_xpb_out[67][592],u_xpb_out[68][592],u_xpb_out[69][592],u_xpb_out[70][592],u_xpb_out[71][592],u_xpb_out[72][592],u_xpb_out[73][592],u_xpb_out[74][592],u_xpb_out[75][592],u_xpb_out[76][592],u_xpb_out[77][592],u_xpb_out[78][592],u_xpb_out[79][592],u_xpb_out[80][592],u_xpb_out[81][592],u_xpb_out[82][592],u_xpb_out[83][592],u_xpb_out[84][592],u_xpb_out[85][592],u_xpb_out[86][592],u_xpb_out[87][592],u_xpb_out[88][592],u_xpb_out[89][592],u_xpb_out[90][592],u_xpb_out[91][592],u_xpb_out[92][592],u_xpb_out[93][592],u_xpb_out[94][592],u_xpb_out[95][592],u_xpb_out[96][592],u_xpb_out[97][592],u_xpb_out[98][592],u_xpb_out[99][592],u_xpb_out[100][592],u_xpb_out[101][592],u_xpb_out[102][592],u_xpb_out[103][592],u_xpb_out[104][592],u_xpb_out[105][592]};

assign col_out_593 = {u_xpb_out[0][593],u_xpb_out[1][593],u_xpb_out[2][593],u_xpb_out[3][593],u_xpb_out[4][593],u_xpb_out[5][593],u_xpb_out[6][593],u_xpb_out[7][593],u_xpb_out[8][593],u_xpb_out[9][593],u_xpb_out[10][593],u_xpb_out[11][593],u_xpb_out[12][593],u_xpb_out[13][593],u_xpb_out[14][593],u_xpb_out[15][593],u_xpb_out[16][593],u_xpb_out[17][593],u_xpb_out[18][593],u_xpb_out[19][593],u_xpb_out[20][593],u_xpb_out[21][593],u_xpb_out[22][593],u_xpb_out[23][593],u_xpb_out[24][593],u_xpb_out[25][593],u_xpb_out[26][593],u_xpb_out[27][593],u_xpb_out[28][593],u_xpb_out[29][593],u_xpb_out[30][593],u_xpb_out[31][593],u_xpb_out[32][593],u_xpb_out[33][593],u_xpb_out[34][593],u_xpb_out[35][593],u_xpb_out[36][593],u_xpb_out[37][593],u_xpb_out[38][593],u_xpb_out[39][593],u_xpb_out[40][593],u_xpb_out[41][593],u_xpb_out[42][593],u_xpb_out[43][593],u_xpb_out[44][593],u_xpb_out[45][593],u_xpb_out[46][593],u_xpb_out[47][593],u_xpb_out[48][593],u_xpb_out[49][593],u_xpb_out[50][593],u_xpb_out[51][593],u_xpb_out[52][593],u_xpb_out[53][593],u_xpb_out[54][593],u_xpb_out[55][593],u_xpb_out[56][593],u_xpb_out[57][593],u_xpb_out[58][593],u_xpb_out[59][593],u_xpb_out[60][593],u_xpb_out[61][593],u_xpb_out[62][593],u_xpb_out[63][593],u_xpb_out[64][593],u_xpb_out[65][593],u_xpb_out[66][593],u_xpb_out[67][593],u_xpb_out[68][593],u_xpb_out[69][593],u_xpb_out[70][593],u_xpb_out[71][593],u_xpb_out[72][593],u_xpb_out[73][593],u_xpb_out[74][593],u_xpb_out[75][593],u_xpb_out[76][593],u_xpb_out[77][593],u_xpb_out[78][593],u_xpb_out[79][593],u_xpb_out[80][593],u_xpb_out[81][593],u_xpb_out[82][593],u_xpb_out[83][593],u_xpb_out[84][593],u_xpb_out[85][593],u_xpb_out[86][593],u_xpb_out[87][593],u_xpb_out[88][593],u_xpb_out[89][593],u_xpb_out[90][593],u_xpb_out[91][593],u_xpb_out[92][593],u_xpb_out[93][593],u_xpb_out[94][593],u_xpb_out[95][593],u_xpb_out[96][593],u_xpb_out[97][593],u_xpb_out[98][593],u_xpb_out[99][593],u_xpb_out[100][593],u_xpb_out[101][593],u_xpb_out[102][593],u_xpb_out[103][593],u_xpb_out[104][593],u_xpb_out[105][593]};

assign col_out_594 = {u_xpb_out[0][594],u_xpb_out[1][594],u_xpb_out[2][594],u_xpb_out[3][594],u_xpb_out[4][594],u_xpb_out[5][594],u_xpb_out[6][594],u_xpb_out[7][594],u_xpb_out[8][594],u_xpb_out[9][594],u_xpb_out[10][594],u_xpb_out[11][594],u_xpb_out[12][594],u_xpb_out[13][594],u_xpb_out[14][594],u_xpb_out[15][594],u_xpb_out[16][594],u_xpb_out[17][594],u_xpb_out[18][594],u_xpb_out[19][594],u_xpb_out[20][594],u_xpb_out[21][594],u_xpb_out[22][594],u_xpb_out[23][594],u_xpb_out[24][594],u_xpb_out[25][594],u_xpb_out[26][594],u_xpb_out[27][594],u_xpb_out[28][594],u_xpb_out[29][594],u_xpb_out[30][594],u_xpb_out[31][594],u_xpb_out[32][594],u_xpb_out[33][594],u_xpb_out[34][594],u_xpb_out[35][594],u_xpb_out[36][594],u_xpb_out[37][594],u_xpb_out[38][594],u_xpb_out[39][594],u_xpb_out[40][594],u_xpb_out[41][594],u_xpb_out[42][594],u_xpb_out[43][594],u_xpb_out[44][594],u_xpb_out[45][594],u_xpb_out[46][594],u_xpb_out[47][594],u_xpb_out[48][594],u_xpb_out[49][594],u_xpb_out[50][594],u_xpb_out[51][594],u_xpb_out[52][594],u_xpb_out[53][594],u_xpb_out[54][594],u_xpb_out[55][594],u_xpb_out[56][594],u_xpb_out[57][594],u_xpb_out[58][594],u_xpb_out[59][594],u_xpb_out[60][594],u_xpb_out[61][594],u_xpb_out[62][594],u_xpb_out[63][594],u_xpb_out[64][594],u_xpb_out[65][594],u_xpb_out[66][594],u_xpb_out[67][594],u_xpb_out[68][594],u_xpb_out[69][594],u_xpb_out[70][594],u_xpb_out[71][594],u_xpb_out[72][594],u_xpb_out[73][594],u_xpb_out[74][594],u_xpb_out[75][594],u_xpb_out[76][594],u_xpb_out[77][594],u_xpb_out[78][594],u_xpb_out[79][594],u_xpb_out[80][594],u_xpb_out[81][594],u_xpb_out[82][594],u_xpb_out[83][594],u_xpb_out[84][594],u_xpb_out[85][594],u_xpb_out[86][594],u_xpb_out[87][594],u_xpb_out[88][594],u_xpb_out[89][594],u_xpb_out[90][594],u_xpb_out[91][594],u_xpb_out[92][594],u_xpb_out[93][594],u_xpb_out[94][594],u_xpb_out[95][594],u_xpb_out[96][594],u_xpb_out[97][594],u_xpb_out[98][594],u_xpb_out[99][594],u_xpb_out[100][594],u_xpb_out[101][594],u_xpb_out[102][594],u_xpb_out[103][594],u_xpb_out[104][594],u_xpb_out[105][594]};

assign col_out_595 = {u_xpb_out[0][595],u_xpb_out[1][595],u_xpb_out[2][595],u_xpb_out[3][595],u_xpb_out[4][595],u_xpb_out[5][595],u_xpb_out[6][595],u_xpb_out[7][595],u_xpb_out[8][595],u_xpb_out[9][595],u_xpb_out[10][595],u_xpb_out[11][595],u_xpb_out[12][595],u_xpb_out[13][595],u_xpb_out[14][595],u_xpb_out[15][595],u_xpb_out[16][595],u_xpb_out[17][595],u_xpb_out[18][595],u_xpb_out[19][595],u_xpb_out[20][595],u_xpb_out[21][595],u_xpb_out[22][595],u_xpb_out[23][595],u_xpb_out[24][595],u_xpb_out[25][595],u_xpb_out[26][595],u_xpb_out[27][595],u_xpb_out[28][595],u_xpb_out[29][595],u_xpb_out[30][595],u_xpb_out[31][595],u_xpb_out[32][595],u_xpb_out[33][595],u_xpb_out[34][595],u_xpb_out[35][595],u_xpb_out[36][595],u_xpb_out[37][595],u_xpb_out[38][595],u_xpb_out[39][595],u_xpb_out[40][595],u_xpb_out[41][595],u_xpb_out[42][595],u_xpb_out[43][595],u_xpb_out[44][595],u_xpb_out[45][595],u_xpb_out[46][595],u_xpb_out[47][595],u_xpb_out[48][595],u_xpb_out[49][595],u_xpb_out[50][595],u_xpb_out[51][595],u_xpb_out[52][595],u_xpb_out[53][595],u_xpb_out[54][595],u_xpb_out[55][595],u_xpb_out[56][595],u_xpb_out[57][595],u_xpb_out[58][595],u_xpb_out[59][595],u_xpb_out[60][595],u_xpb_out[61][595],u_xpb_out[62][595],u_xpb_out[63][595],u_xpb_out[64][595],u_xpb_out[65][595],u_xpb_out[66][595],u_xpb_out[67][595],u_xpb_out[68][595],u_xpb_out[69][595],u_xpb_out[70][595],u_xpb_out[71][595],u_xpb_out[72][595],u_xpb_out[73][595],u_xpb_out[74][595],u_xpb_out[75][595],u_xpb_out[76][595],u_xpb_out[77][595],u_xpb_out[78][595],u_xpb_out[79][595],u_xpb_out[80][595],u_xpb_out[81][595],u_xpb_out[82][595],u_xpb_out[83][595],u_xpb_out[84][595],u_xpb_out[85][595],u_xpb_out[86][595],u_xpb_out[87][595],u_xpb_out[88][595],u_xpb_out[89][595],u_xpb_out[90][595],u_xpb_out[91][595],u_xpb_out[92][595],u_xpb_out[93][595],u_xpb_out[94][595],u_xpb_out[95][595],u_xpb_out[96][595],u_xpb_out[97][595],u_xpb_out[98][595],u_xpb_out[99][595],u_xpb_out[100][595],u_xpb_out[101][595],u_xpb_out[102][595],u_xpb_out[103][595],u_xpb_out[104][595],u_xpb_out[105][595]};

assign col_out_596 = {u_xpb_out[0][596],u_xpb_out[1][596],u_xpb_out[2][596],u_xpb_out[3][596],u_xpb_out[4][596],u_xpb_out[5][596],u_xpb_out[6][596],u_xpb_out[7][596],u_xpb_out[8][596],u_xpb_out[9][596],u_xpb_out[10][596],u_xpb_out[11][596],u_xpb_out[12][596],u_xpb_out[13][596],u_xpb_out[14][596],u_xpb_out[15][596],u_xpb_out[16][596],u_xpb_out[17][596],u_xpb_out[18][596],u_xpb_out[19][596],u_xpb_out[20][596],u_xpb_out[21][596],u_xpb_out[22][596],u_xpb_out[23][596],u_xpb_out[24][596],u_xpb_out[25][596],u_xpb_out[26][596],u_xpb_out[27][596],u_xpb_out[28][596],u_xpb_out[29][596],u_xpb_out[30][596],u_xpb_out[31][596],u_xpb_out[32][596],u_xpb_out[33][596],u_xpb_out[34][596],u_xpb_out[35][596],u_xpb_out[36][596],u_xpb_out[37][596],u_xpb_out[38][596],u_xpb_out[39][596],u_xpb_out[40][596],u_xpb_out[41][596],u_xpb_out[42][596],u_xpb_out[43][596],u_xpb_out[44][596],u_xpb_out[45][596],u_xpb_out[46][596],u_xpb_out[47][596],u_xpb_out[48][596],u_xpb_out[49][596],u_xpb_out[50][596],u_xpb_out[51][596],u_xpb_out[52][596],u_xpb_out[53][596],u_xpb_out[54][596],u_xpb_out[55][596],u_xpb_out[56][596],u_xpb_out[57][596],u_xpb_out[58][596],u_xpb_out[59][596],u_xpb_out[60][596],u_xpb_out[61][596],u_xpb_out[62][596],u_xpb_out[63][596],u_xpb_out[64][596],u_xpb_out[65][596],u_xpb_out[66][596],u_xpb_out[67][596],u_xpb_out[68][596],u_xpb_out[69][596],u_xpb_out[70][596],u_xpb_out[71][596],u_xpb_out[72][596],u_xpb_out[73][596],u_xpb_out[74][596],u_xpb_out[75][596],u_xpb_out[76][596],u_xpb_out[77][596],u_xpb_out[78][596],u_xpb_out[79][596],u_xpb_out[80][596],u_xpb_out[81][596],u_xpb_out[82][596],u_xpb_out[83][596],u_xpb_out[84][596],u_xpb_out[85][596],u_xpb_out[86][596],u_xpb_out[87][596],u_xpb_out[88][596],u_xpb_out[89][596],u_xpb_out[90][596],u_xpb_out[91][596],u_xpb_out[92][596],u_xpb_out[93][596],u_xpb_out[94][596],u_xpb_out[95][596],u_xpb_out[96][596],u_xpb_out[97][596],u_xpb_out[98][596],u_xpb_out[99][596],u_xpb_out[100][596],u_xpb_out[101][596],u_xpb_out[102][596],u_xpb_out[103][596],u_xpb_out[104][596],u_xpb_out[105][596]};

assign col_out_597 = {u_xpb_out[0][597],u_xpb_out[1][597],u_xpb_out[2][597],u_xpb_out[3][597],u_xpb_out[4][597],u_xpb_out[5][597],u_xpb_out[6][597],u_xpb_out[7][597],u_xpb_out[8][597],u_xpb_out[9][597],u_xpb_out[10][597],u_xpb_out[11][597],u_xpb_out[12][597],u_xpb_out[13][597],u_xpb_out[14][597],u_xpb_out[15][597],u_xpb_out[16][597],u_xpb_out[17][597],u_xpb_out[18][597],u_xpb_out[19][597],u_xpb_out[20][597],u_xpb_out[21][597],u_xpb_out[22][597],u_xpb_out[23][597],u_xpb_out[24][597],u_xpb_out[25][597],u_xpb_out[26][597],u_xpb_out[27][597],u_xpb_out[28][597],u_xpb_out[29][597],u_xpb_out[30][597],u_xpb_out[31][597],u_xpb_out[32][597],u_xpb_out[33][597],u_xpb_out[34][597],u_xpb_out[35][597],u_xpb_out[36][597],u_xpb_out[37][597],u_xpb_out[38][597],u_xpb_out[39][597],u_xpb_out[40][597],u_xpb_out[41][597],u_xpb_out[42][597],u_xpb_out[43][597],u_xpb_out[44][597],u_xpb_out[45][597],u_xpb_out[46][597],u_xpb_out[47][597],u_xpb_out[48][597],u_xpb_out[49][597],u_xpb_out[50][597],u_xpb_out[51][597],u_xpb_out[52][597],u_xpb_out[53][597],u_xpb_out[54][597],u_xpb_out[55][597],u_xpb_out[56][597],u_xpb_out[57][597],u_xpb_out[58][597],u_xpb_out[59][597],u_xpb_out[60][597],u_xpb_out[61][597],u_xpb_out[62][597],u_xpb_out[63][597],u_xpb_out[64][597],u_xpb_out[65][597],u_xpb_out[66][597],u_xpb_out[67][597],u_xpb_out[68][597],u_xpb_out[69][597],u_xpb_out[70][597],u_xpb_out[71][597],u_xpb_out[72][597],u_xpb_out[73][597],u_xpb_out[74][597],u_xpb_out[75][597],u_xpb_out[76][597],u_xpb_out[77][597],u_xpb_out[78][597],u_xpb_out[79][597],u_xpb_out[80][597],u_xpb_out[81][597],u_xpb_out[82][597],u_xpb_out[83][597],u_xpb_out[84][597],u_xpb_out[85][597],u_xpb_out[86][597],u_xpb_out[87][597],u_xpb_out[88][597],u_xpb_out[89][597],u_xpb_out[90][597],u_xpb_out[91][597],u_xpb_out[92][597],u_xpb_out[93][597],u_xpb_out[94][597],u_xpb_out[95][597],u_xpb_out[96][597],u_xpb_out[97][597],u_xpb_out[98][597],u_xpb_out[99][597],u_xpb_out[100][597],u_xpb_out[101][597],u_xpb_out[102][597],u_xpb_out[103][597],u_xpb_out[104][597],u_xpb_out[105][597]};

assign col_out_598 = {u_xpb_out[0][598],u_xpb_out[1][598],u_xpb_out[2][598],u_xpb_out[3][598],u_xpb_out[4][598],u_xpb_out[5][598],u_xpb_out[6][598],u_xpb_out[7][598],u_xpb_out[8][598],u_xpb_out[9][598],u_xpb_out[10][598],u_xpb_out[11][598],u_xpb_out[12][598],u_xpb_out[13][598],u_xpb_out[14][598],u_xpb_out[15][598],u_xpb_out[16][598],u_xpb_out[17][598],u_xpb_out[18][598],u_xpb_out[19][598],u_xpb_out[20][598],u_xpb_out[21][598],u_xpb_out[22][598],u_xpb_out[23][598],u_xpb_out[24][598],u_xpb_out[25][598],u_xpb_out[26][598],u_xpb_out[27][598],u_xpb_out[28][598],u_xpb_out[29][598],u_xpb_out[30][598],u_xpb_out[31][598],u_xpb_out[32][598],u_xpb_out[33][598],u_xpb_out[34][598],u_xpb_out[35][598],u_xpb_out[36][598],u_xpb_out[37][598],u_xpb_out[38][598],u_xpb_out[39][598],u_xpb_out[40][598],u_xpb_out[41][598],u_xpb_out[42][598],u_xpb_out[43][598],u_xpb_out[44][598],u_xpb_out[45][598],u_xpb_out[46][598],u_xpb_out[47][598],u_xpb_out[48][598],u_xpb_out[49][598],u_xpb_out[50][598],u_xpb_out[51][598],u_xpb_out[52][598],u_xpb_out[53][598],u_xpb_out[54][598],u_xpb_out[55][598],u_xpb_out[56][598],u_xpb_out[57][598],u_xpb_out[58][598],u_xpb_out[59][598],u_xpb_out[60][598],u_xpb_out[61][598],u_xpb_out[62][598],u_xpb_out[63][598],u_xpb_out[64][598],u_xpb_out[65][598],u_xpb_out[66][598],u_xpb_out[67][598],u_xpb_out[68][598],u_xpb_out[69][598],u_xpb_out[70][598],u_xpb_out[71][598],u_xpb_out[72][598],u_xpb_out[73][598],u_xpb_out[74][598],u_xpb_out[75][598],u_xpb_out[76][598],u_xpb_out[77][598],u_xpb_out[78][598],u_xpb_out[79][598],u_xpb_out[80][598],u_xpb_out[81][598],u_xpb_out[82][598],u_xpb_out[83][598],u_xpb_out[84][598],u_xpb_out[85][598],u_xpb_out[86][598],u_xpb_out[87][598],u_xpb_out[88][598],u_xpb_out[89][598],u_xpb_out[90][598],u_xpb_out[91][598],u_xpb_out[92][598],u_xpb_out[93][598],u_xpb_out[94][598],u_xpb_out[95][598],u_xpb_out[96][598],u_xpb_out[97][598],u_xpb_out[98][598],u_xpb_out[99][598],u_xpb_out[100][598],u_xpb_out[101][598],u_xpb_out[102][598],u_xpb_out[103][598],u_xpb_out[104][598],u_xpb_out[105][598]};

assign col_out_599 = {u_xpb_out[0][599],u_xpb_out[1][599],u_xpb_out[2][599],u_xpb_out[3][599],u_xpb_out[4][599],u_xpb_out[5][599],u_xpb_out[6][599],u_xpb_out[7][599],u_xpb_out[8][599],u_xpb_out[9][599],u_xpb_out[10][599],u_xpb_out[11][599],u_xpb_out[12][599],u_xpb_out[13][599],u_xpb_out[14][599],u_xpb_out[15][599],u_xpb_out[16][599],u_xpb_out[17][599],u_xpb_out[18][599],u_xpb_out[19][599],u_xpb_out[20][599],u_xpb_out[21][599],u_xpb_out[22][599],u_xpb_out[23][599],u_xpb_out[24][599],u_xpb_out[25][599],u_xpb_out[26][599],u_xpb_out[27][599],u_xpb_out[28][599],u_xpb_out[29][599],u_xpb_out[30][599],u_xpb_out[31][599],u_xpb_out[32][599],u_xpb_out[33][599],u_xpb_out[34][599],u_xpb_out[35][599],u_xpb_out[36][599],u_xpb_out[37][599],u_xpb_out[38][599],u_xpb_out[39][599],u_xpb_out[40][599],u_xpb_out[41][599],u_xpb_out[42][599],u_xpb_out[43][599],u_xpb_out[44][599],u_xpb_out[45][599],u_xpb_out[46][599],u_xpb_out[47][599],u_xpb_out[48][599],u_xpb_out[49][599],u_xpb_out[50][599],u_xpb_out[51][599],u_xpb_out[52][599],u_xpb_out[53][599],u_xpb_out[54][599],u_xpb_out[55][599],u_xpb_out[56][599],u_xpb_out[57][599],u_xpb_out[58][599],u_xpb_out[59][599],u_xpb_out[60][599],u_xpb_out[61][599],u_xpb_out[62][599],u_xpb_out[63][599],u_xpb_out[64][599],u_xpb_out[65][599],u_xpb_out[66][599],u_xpb_out[67][599],u_xpb_out[68][599],u_xpb_out[69][599],u_xpb_out[70][599],u_xpb_out[71][599],u_xpb_out[72][599],u_xpb_out[73][599],u_xpb_out[74][599],u_xpb_out[75][599],u_xpb_out[76][599],u_xpb_out[77][599],u_xpb_out[78][599],u_xpb_out[79][599],u_xpb_out[80][599],u_xpb_out[81][599],u_xpb_out[82][599],u_xpb_out[83][599],u_xpb_out[84][599],u_xpb_out[85][599],u_xpb_out[86][599],u_xpb_out[87][599],u_xpb_out[88][599],u_xpb_out[89][599],u_xpb_out[90][599],u_xpb_out[91][599],u_xpb_out[92][599],u_xpb_out[93][599],u_xpb_out[94][599],u_xpb_out[95][599],u_xpb_out[96][599],u_xpb_out[97][599],u_xpb_out[98][599],u_xpb_out[99][599],u_xpb_out[100][599],u_xpb_out[101][599],u_xpb_out[102][599],u_xpb_out[103][599],u_xpb_out[104][599],u_xpb_out[105][599]};

assign col_out_600 = {u_xpb_out[0][600],u_xpb_out[1][600],u_xpb_out[2][600],u_xpb_out[3][600],u_xpb_out[4][600],u_xpb_out[5][600],u_xpb_out[6][600],u_xpb_out[7][600],u_xpb_out[8][600],u_xpb_out[9][600],u_xpb_out[10][600],u_xpb_out[11][600],u_xpb_out[12][600],u_xpb_out[13][600],u_xpb_out[14][600],u_xpb_out[15][600],u_xpb_out[16][600],u_xpb_out[17][600],u_xpb_out[18][600],u_xpb_out[19][600],u_xpb_out[20][600],u_xpb_out[21][600],u_xpb_out[22][600],u_xpb_out[23][600],u_xpb_out[24][600],u_xpb_out[25][600],u_xpb_out[26][600],u_xpb_out[27][600],u_xpb_out[28][600],u_xpb_out[29][600],u_xpb_out[30][600],u_xpb_out[31][600],u_xpb_out[32][600],u_xpb_out[33][600],u_xpb_out[34][600],u_xpb_out[35][600],u_xpb_out[36][600],u_xpb_out[37][600],u_xpb_out[38][600],u_xpb_out[39][600],u_xpb_out[40][600],u_xpb_out[41][600],u_xpb_out[42][600],u_xpb_out[43][600],u_xpb_out[44][600],u_xpb_out[45][600],u_xpb_out[46][600],u_xpb_out[47][600],u_xpb_out[48][600],u_xpb_out[49][600],u_xpb_out[50][600],u_xpb_out[51][600],u_xpb_out[52][600],u_xpb_out[53][600],u_xpb_out[54][600],u_xpb_out[55][600],u_xpb_out[56][600],u_xpb_out[57][600],u_xpb_out[58][600],u_xpb_out[59][600],u_xpb_out[60][600],u_xpb_out[61][600],u_xpb_out[62][600],u_xpb_out[63][600],u_xpb_out[64][600],u_xpb_out[65][600],u_xpb_out[66][600],u_xpb_out[67][600],u_xpb_out[68][600],u_xpb_out[69][600],u_xpb_out[70][600],u_xpb_out[71][600],u_xpb_out[72][600],u_xpb_out[73][600],u_xpb_out[74][600],u_xpb_out[75][600],u_xpb_out[76][600],u_xpb_out[77][600],u_xpb_out[78][600],u_xpb_out[79][600],u_xpb_out[80][600],u_xpb_out[81][600],u_xpb_out[82][600],u_xpb_out[83][600],u_xpb_out[84][600],u_xpb_out[85][600],u_xpb_out[86][600],u_xpb_out[87][600],u_xpb_out[88][600],u_xpb_out[89][600],u_xpb_out[90][600],u_xpb_out[91][600],u_xpb_out[92][600],u_xpb_out[93][600],u_xpb_out[94][600],u_xpb_out[95][600],u_xpb_out[96][600],u_xpb_out[97][600],u_xpb_out[98][600],u_xpb_out[99][600],u_xpb_out[100][600],u_xpb_out[101][600],u_xpb_out[102][600],u_xpb_out[103][600],u_xpb_out[104][600],u_xpb_out[105][600]};

assign col_out_601 = {u_xpb_out[0][601],u_xpb_out[1][601],u_xpb_out[2][601],u_xpb_out[3][601],u_xpb_out[4][601],u_xpb_out[5][601],u_xpb_out[6][601],u_xpb_out[7][601],u_xpb_out[8][601],u_xpb_out[9][601],u_xpb_out[10][601],u_xpb_out[11][601],u_xpb_out[12][601],u_xpb_out[13][601],u_xpb_out[14][601],u_xpb_out[15][601],u_xpb_out[16][601],u_xpb_out[17][601],u_xpb_out[18][601],u_xpb_out[19][601],u_xpb_out[20][601],u_xpb_out[21][601],u_xpb_out[22][601],u_xpb_out[23][601],u_xpb_out[24][601],u_xpb_out[25][601],u_xpb_out[26][601],u_xpb_out[27][601],u_xpb_out[28][601],u_xpb_out[29][601],u_xpb_out[30][601],u_xpb_out[31][601],u_xpb_out[32][601],u_xpb_out[33][601],u_xpb_out[34][601],u_xpb_out[35][601],u_xpb_out[36][601],u_xpb_out[37][601],u_xpb_out[38][601],u_xpb_out[39][601],u_xpb_out[40][601],u_xpb_out[41][601],u_xpb_out[42][601],u_xpb_out[43][601],u_xpb_out[44][601],u_xpb_out[45][601],u_xpb_out[46][601],u_xpb_out[47][601],u_xpb_out[48][601],u_xpb_out[49][601],u_xpb_out[50][601],u_xpb_out[51][601],u_xpb_out[52][601],u_xpb_out[53][601],u_xpb_out[54][601],u_xpb_out[55][601],u_xpb_out[56][601],u_xpb_out[57][601],u_xpb_out[58][601],u_xpb_out[59][601],u_xpb_out[60][601],u_xpb_out[61][601],u_xpb_out[62][601],u_xpb_out[63][601],u_xpb_out[64][601],u_xpb_out[65][601],u_xpb_out[66][601],u_xpb_out[67][601],u_xpb_out[68][601],u_xpb_out[69][601],u_xpb_out[70][601],u_xpb_out[71][601],u_xpb_out[72][601],u_xpb_out[73][601],u_xpb_out[74][601],u_xpb_out[75][601],u_xpb_out[76][601],u_xpb_out[77][601],u_xpb_out[78][601],u_xpb_out[79][601],u_xpb_out[80][601],u_xpb_out[81][601],u_xpb_out[82][601],u_xpb_out[83][601],u_xpb_out[84][601],u_xpb_out[85][601],u_xpb_out[86][601],u_xpb_out[87][601],u_xpb_out[88][601],u_xpb_out[89][601],u_xpb_out[90][601],u_xpb_out[91][601],u_xpb_out[92][601],u_xpb_out[93][601],u_xpb_out[94][601],u_xpb_out[95][601],u_xpb_out[96][601],u_xpb_out[97][601],u_xpb_out[98][601],u_xpb_out[99][601],u_xpb_out[100][601],u_xpb_out[101][601],u_xpb_out[102][601],u_xpb_out[103][601],u_xpb_out[104][601],u_xpb_out[105][601]};

assign col_out_602 = {u_xpb_out[0][602],u_xpb_out[1][602],u_xpb_out[2][602],u_xpb_out[3][602],u_xpb_out[4][602],u_xpb_out[5][602],u_xpb_out[6][602],u_xpb_out[7][602],u_xpb_out[8][602],u_xpb_out[9][602],u_xpb_out[10][602],u_xpb_out[11][602],u_xpb_out[12][602],u_xpb_out[13][602],u_xpb_out[14][602],u_xpb_out[15][602],u_xpb_out[16][602],u_xpb_out[17][602],u_xpb_out[18][602],u_xpb_out[19][602],u_xpb_out[20][602],u_xpb_out[21][602],u_xpb_out[22][602],u_xpb_out[23][602],u_xpb_out[24][602],u_xpb_out[25][602],u_xpb_out[26][602],u_xpb_out[27][602],u_xpb_out[28][602],u_xpb_out[29][602],u_xpb_out[30][602],u_xpb_out[31][602],u_xpb_out[32][602],u_xpb_out[33][602],u_xpb_out[34][602],u_xpb_out[35][602],u_xpb_out[36][602],u_xpb_out[37][602],u_xpb_out[38][602],u_xpb_out[39][602],u_xpb_out[40][602],u_xpb_out[41][602],u_xpb_out[42][602],u_xpb_out[43][602],u_xpb_out[44][602],u_xpb_out[45][602],u_xpb_out[46][602],u_xpb_out[47][602],u_xpb_out[48][602],u_xpb_out[49][602],u_xpb_out[50][602],u_xpb_out[51][602],u_xpb_out[52][602],u_xpb_out[53][602],u_xpb_out[54][602],u_xpb_out[55][602],u_xpb_out[56][602],u_xpb_out[57][602],u_xpb_out[58][602],u_xpb_out[59][602],u_xpb_out[60][602],u_xpb_out[61][602],u_xpb_out[62][602],u_xpb_out[63][602],u_xpb_out[64][602],u_xpb_out[65][602],u_xpb_out[66][602],u_xpb_out[67][602],u_xpb_out[68][602],u_xpb_out[69][602],u_xpb_out[70][602],u_xpb_out[71][602],u_xpb_out[72][602],u_xpb_out[73][602],u_xpb_out[74][602],u_xpb_out[75][602],u_xpb_out[76][602],u_xpb_out[77][602],u_xpb_out[78][602],u_xpb_out[79][602],u_xpb_out[80][602],u_xpb_out[81][602],u_xpb_out[82][602],u_xpb_out[83][602],u_xpb_out[84][602],u_xpb_out[85][602],u_xpb_out[86][602],u_xpb_out[87][602],u_xpb_out[88][602],u_xpb_out[89][602],u_xpb_out[90][602],u_xpb_out[91][602],u_xpb_out[92][602],u_xpb_out[93][602],u_xpb_out[94][602],u_xpb_out[95][602],u_xpb_out[96][602],u_xpb_out[97][602],u_xpb_out[98][602],u_xpb_out[99][602],u_xpb_out[100][602],u_xpb_out[101][602],u_xpb_out[102][602],u_xpb_out[103][602],u_xpb_out[104][602],u_xpb_out[105][602]};

assign col_out_603 = {u_xpb_out[0][603],u_xpb_out[1][603],u_xpb_out[2][603],u_xpb_out[3][603],u_xpb_out[4][603],u_xpb_out[5][603],u_xpb_out[6][603],u_xpb_out[7][603],u_xpb_out[8][603],u_xpb_out[9][603],u_xpb_out[10][603],u_xpb_out[11][603],u_xpb_out[12][603],u_xpb_out[13][603],u_xpb_out[14][603],u_xpb_out[15][603],u_xpb_out[16][603],u_xpb_out[17][603],u_xpb_out[18][603],u_xpb_out[19][603],u_xpb_out[20][603],u_xpb_out[21][603],u_xpb_out[22][603],u_xpb_out[23][603],u_xpb_out[24][603],u_xpb_out[25][603],u_xpb_out[26][603],u_xpb_out[27][603],u_xpb_out[28][603],u_xpb_out[29][603],u_xpb_out[30][603],u_xpb_out[31][603],u_xpb_out[32][603],u_xpb_out[33][603],u_xpb_out[34][603],u_xpb_out[35][603],u_xpb_out[36][603],u_xpb_out[37][603],u_xpb_out[38][603],u_xpb_out[39][603],u_xpb_out[40][603],u_xpb_out[41][603],u_xpb_out[42][603],u_xpb_out[43][603],u_xpb_out[44][603],u_xpb_out[45][603],u_xpb_out[46][603],u_xpb_out[47][603],u_xpb_out[48][603],u_xpb_out[49][603],u_xpb_out[50][603],u_xpb_out[51][603],u_xpb_out[52][603],u_xpb_out[53][603],u_xpb_out[54][603],u_xpb_out[55][603],u_xpb_out[56][603],u_xpb_out[57][603],u_xpb_out[58][603],u_xpb_out[59][603],u_xpb_out[60][603],u_xpb_out[61][603],u_xpb_out[62][603],u_xpb_out[63][603],u_xpb_out[64][603],u_xpb_out[65][603],u_xpb_out[66][603],u_xpb_out[67][603],u_xpb_out[68][603],u_xpb_out[69][603],u_xpb_out[70][603],u_xpb_out[71][603],u_xpb_out[72][603],u_xpb_out[73][603],u_xpb_out[74][603],u_xpb_out[75][603],u_xpb_out[76][603],u_xpb_out[77][603],u_xpb_out[78][603],u_xpb_out[79][603],u_xpb_out[80][603],u_xpb_out[81][603],u_xpb_out[82][603],u_xpb_out[83][603],u_xpb_out[84][603],u_xpb_out[85][603],u_xpb_out[86][603],u_xpb_out[87][603],u_xpb_out[88][603],u_xpb_out[89][603],u_xpb_out[90][603],u_xpb_out[91][603],u_xpb_out[92][603],u_xpb_out[93][603],u_xpb_out[94][603],u_xpb_out[95][603],u_xpb_out[96][603],u_xpb_out[97][603],u_xpb_out[98][603],u_xpb_out[99][603],u_xpb_out[100][603],u_xpb_out[101][603],u_xpb_out[102][603],u_xpb_out[103][603],u_xpb_out[104][603],u_xpb_out[105][603]};

assign col_out_604 = {u_xpb_out[0][604],u_xpb_out[1][604],u_xpb_out[2][604],u_xpb_out[3][604],u_xpb_out[4][604],u_xpb_out[5][604],u_xpb_out[6][604],u_xpb_out[7][604],u_xpb_out[8][604],u_xpb_out[9][604],u_xpb_out[10][604],u_xpb_out[11][604],u_xpb_out[12][604],u_xpb_out[13][604],u_xpb_out[14][604],u_xpb_out[15][604],u_xpb_out[16][604],u_xpb_out[17][604],u_xpb_out[18][604],u_xpb_out[19][604],u_xpb_out[20][604],u_xpb_out[21][604],u_xpb_out[22][604],u_xpb_out[23][604],u_xpb_out[24][604],u_xpb_out[25][604],u_xpb_out[26][604],u_xpb_out[27][604],u_xpb_out[28][604],u_xpb_out[29][604],u_xpb_out[30][604],u_xpb_out[31][604],u_xpb_out[32][604],u_xpb_out[33][604],u_xpb_out[34][604],u_xpb_out[35][604],u_xpb_out[36][604],u_xpb_out[37][604],u_xpb_out[38][604],u_xpb_out[39][604],u_xpb_out[40][604],u_xpb_out[41][604],u_xpb_out[42][604],u_xpb_out[43][604],u_xpb_out[44][604],u_xpb_out[45][604],u_xpb_out[46][604],u_xpb_out[47][604],u_xpb_out[48][604],u_xpb_out[49][604],u_xpb_out[50][604],u_xpb_out[51][604],u_xpb_out[52][604],u_xpb_out[53][604],u_xpb_out[54][604],u_xpb_out[55][604],u_xpb_out[56][604],u_xpb_out[57][604],u_xpb_out[58][604],u_xpb_out[59][604],u_xpb_out[60][604],u_xpb_out[61][604],u_xpb_out[62][604],u_xpb_out[63][604],u_xpb_out[64][604],u_xpb_out[65][604],u_xpb_out[66][604],u_xpb_out[67][604],u_xpb_out[68][604],u_xpb_out[69][604],u_xpb_out[70][604],u_xpb_out[71][604],u_xpb_out[72][604],u_xpb_out[73][604],u_xpb_out[74][604],u_xpb_out[75][604],u_xpb_out[76][604],u_xpb_out[77][604],u_xpb_out[78][604],u_xpb_out[79][604],u_xpb_out[80][604],u_xpb_out[81][604],u_xpb_out[82][604],u_xpb_out[83][604],u_xpb_out[84][604],u_xpb_out[85][604],u_xpb_out[86][604],u_xpb_out[87][604],u_xpb_out[88][604],u_xpb_out[89][604],u_xpb_out[90][604],u_xpb_out[91][604],u_xpb_out[92][604],u_xpb_out[93][604],u_xpb_out[94][604],u_xpb_out[95][604],u_xpb_out[96][604],u_xpb_out[97][604],u_xpb_out[98][604],u_xpb_out[99][604],u_xpb_out[100][604],u_xpb_out[101][604],u_xpb_out[102][604],u_xpb_out[103][604],u_xpb_out[104][604],u_xpb_out[105][604]};

assign col_out_605 = {u_xpb_out[0][605],u_xpb_out[1][605],u_xpb_out[2][605],u_xpb_out[3][605],u_xpb_out[4][605],u_xpb_out[5][605],u_xpb_out[6][605],u_xpb_out[7][605],u_xpb_out[8][605],u_xpb_out[9][605],u_xpb_out[10][605],u_xpb_out[11][605],u_xpb_out[12][605],u_xpb_out[13][605],u_xpb_out[14][605],u_xpb_out[15][605],u_xpb_out[16][605],u_xpb_out[17][605],u_xpb_out[18][605],u_xpb_out[19][605],u_xpb_out[20][605],u_xpb_out[21][605],u_xpb_out[22][605],u_xpb_out[23][605],u_xpb_out[24][605],u_xpb_out[25][605],u_xpb_out[26][605],u_xpb_out[27][605],u_xpb_out[28][605],u_xpb_out[29][605],u_xpb_out[30][605],u_xpb_out[31][605],u_xpb_out[32][605],u_xpb_out[33][605],u_xpb_out[34][605],u_xpb_out[35][605],u_xpb_out[36][605],u_xpb_out[37][605],u_xpb_out[38][605],u_xpb_out[39][605],u_xpb_out[40][605],u_xpb_out[41][605],u_xpb_out[42][605],u_xpb_out[43][605],u_xpb_out[44][605],u_xpb_out[45][605],u_xpb_out[46][605],u_xpb_out[47][605],u_xpb_out[48][605],u_xpb_out[49][605],u_xpb_out[50][605],u_xpb_out[51][605],u_xpb_out[52][605],u_xpb_out[53][605],u_xpb_out[54][605],u_xpb_out[55][605],u_xpb_out[56][605],u_xpb_out[57][605],u_xpb_out[58][605],u_xpb_out[59][605],u_xpb_out[60][605],u_xpb_out[61][605],u_xpb_out[62][605],u_xpb_out[63][605],u_xpb_out[64][605],u_xpb_out[65][605],u_xpb_out[66][605],u_xpb_out[67][605],u_xpb_out[68][605],u_xpb_out[69][605],u_xpb_out[70][605],u_xpb_out[71][605],u_xpb_out[72][605],u_xpb_out[73][605],u_xpb_out[74][605],u_xpb_out[75][605],u_xpb_out[76][605],u_xpb_out[77][605],u_xpb_out[78][605],u_xpb_out[79][605],u_xpb_out[80][605],u_xpb_out[81][605],u_xpb_out[82][605],u_xpb_out[83][605],u_xpb_out[84][605],u_xpb_out[85][605],u_xpb_out[86][605],u_xpb_out[87][605],u_xpb_out[88][605],u_xpb_out[89][605],u_xpb_out[90][605],u_xpb_out[91][605],u_xpb_out[92][605],u_xpb_out[93][605],u_xpb_out[94][605],u_xpb_out[95][605],u_xpb_out[96][605],u_xpb_out[97][605],u_xpb_out[98][605],u_xpb_out[99][605],u_xpb_out[100][605],u_xpb_out[101][605],u_xpb_out[102][605],u_xpb_out[103][605],u_xpb_out[104][605],u_xpb_out[105][605]};

assign col_out_606 = {u_xpb_out[0][606],u_xpb_out[1][606],u_xpb_out[2][606],u_xpb_out[3][606],u_xpb_out[4][606],u_xpb_out[5][606],u_xpb_out[6][606],u_xpb_out[7][606],u_xpb_out[8][606],u_xpb_out[9][606],u_xpb_out[10][606],u_xpb_out[11][606],u_xpb_out[12][606],u_xpb_out[13][606],u_xpb_out[14][606],u_xpb_out[15][606],u_xpb_out[16][606],u_xpb_out[17][606],u_xpb_out[18][606],u_xpb_out[19][606],u_xpb_out[20][606],u_xpb_out[21][606],u_xpb_out[22][606],u_xpb_out[23][606],u_xpb_out[24][606],u_xpb_out[25][606],u_xpb_out[26][606],u_xpb_out[27][606],u_xpb_out[28][606],u_xpb_out[29][606],u_xpb_out[30][606],u_xpb_out[31][606],u_xpb_out[32][606],u_xpb_out[33][606],u_xpb_out[34][606],u_xpb_out[35][606],u_xpb_out[36][606],u_xpb_out[37][606],u_xpb_out[38][606],u_xpb_out[39][606],u_xpb_out[40][606],u_xpb_out[41][606],u_xpb_out[42][606],u_xpb_out[43][606],u_xpb_out[44][606],u_xpb_out[45][606],u_xpb_out[46][606],u_xpb_out[47][606],u_xpb_out[48][606],u_xpb_out[49][606],u_xpb_out[50][606],u_xpb_out[51][606],u_xpb_out[52][606],u_xpb_out[53][606],u_xpb_out[54][606],u_xpb_out[55][606],u_xpb_out[56][606],u_xpb_out[57][606],u_xpb_out[58][606],u_xpb_out[59][606],u_xpb_out[60][606],u_xpb_out[61][606],u_xpb_out[62][606],u_xpb_out[63][606],u_xpb_out[64][606],u_xpb_out[65][606],u_xpb_out[66][606],u_xpb_out[67][606],u_xpb_out[68][606],u_xpb_out[69][606],u_xpb_out[70][606],u_xpb_out[71][606],u_xpb_out[72][606],u_xpb_out[73][606],u_xpb_out[74][606],u_xpb_out[75][606],u_xpb_out[76][606],u_xpb_out[77][606],u_xpb_out[78][606],u_xpb_out[79][606],u_xpb_out[80][606],u_xpb_out[81][606],u_xpb_out[82][606],u_xpb_out[83][606],u_xpb_out[84][606],u_xpb_out[85][606],u_xpb_out[86][606],u_xpb_out[87][606],u_xpb_out[88][606],u_xpb_out[89][606],u_xpb_out[90][606],u_xpb_out[91][606],u_xpb_out[92][606],u_xpb_out[93][606],u_xpb_out[94][606],u_xpb_out[95][606],u_xpb_out[96][606],u_xpb_out[97][606],u_xpb_out[98][606],u_xpb_out[99][606],u_xpb_out[100][606],u_xpb_out[101][606],u_xpb_out[102][606],u_xpb_out[103][606],u_xpb_out[104][606],u_xpb_out[105][606]};

assign col_out_607 = {u_xpb_out[0][607],u_xpb_out[1][607],u_xpb_out[2][607],u_xpb_out[3][607],u_xpb_out[4][607],u_xpb_out[5][607],u_xpb_out[6][607],u_xpb_out[7][607],u_xpb_out[8][607],u_xpb_out[9][607],u_xpb_out[10][607],u_xpb_out[11][607],u_xpb_out[12][607],u_xpb_out[13][607],u_xpb_out[14][607],u_xpb_out[15][607],u_xpb_out[16][607],u_xpb_out[17][607],u_xpb_out[18][607],u_xpb_out[19][607],u_xpb_out[20][607],u_xpb_out[21][607],u_xpb_out[22][607],u_xpb_out[23][607],u_xpb_out[24][607],u_xpb_out[25][607],u_xpb_out[26][607],u_xpb_out[27][607],u_xpb_out[28][607],u_xpb_out[29][607],u_xpb_out[30][607],u_xpb_out[31][607],u_xpb_out[32][607],u_xpb_out[33][607],u_xpb_out[34][607],u_xpb_out[35][607],u_xpb_out[36][607],u_xpb_out[37][607],u_xpb_out[38][607],u_xpb_out[39][607],u_xpb_out[40][607],u_xpb_out[41][607],u_xpb_out[42][607],u_xpb_out[43][607],u_xpb_out[44][607],u_xpb_out[45][607],u_xpb_out[46][607],u_xpb_out[47][607],u_xpb_out[48][607],u_xpb_out[49][607],u_xpb_out[50][607],u_xpb_out[51][607],u_xpb_out[52][607],u_xpb_out[53][607],u_xpb_out[54][607],u_xpb_out[55][607],u_xpb_out[56][607],u_xpb_out[57][607],u_xpb_out[58][607],u_xpb_out[59][607],u_xpb_out[60][607],u_xpb_out[61][607],u_xpb_out[62][607],u_xpb_out[63][607],u_xpb_out[64][607],u_xpb_out[65][607],u_xpb_out[66][607],u_xpb_out[67][607],u_xpb_out[68][607],u_xpb_out[69][607],u_xpb_out[70][607],u_xpb_out[71][607],u_xpb_out[72][607],u_xpb_out[73][607],u_xpb_out[74][607],u_xpb_out[75][607],u_xpb_out[76][607],u_xpb_out[77][607],u_xpb_out[78][607],u_xpb_out[79][607],u_xpb_out[80][607],u_xpb_out[81][607],u_xpb_out[82][607],u_xpb_out[83][607],u_xpb_out[84][607],u_xpb_out[85][607],u_xpb_out[86][607],u_xpb_out[87][607],u_xpb_out[88][607],u_xpb_out[89][607],u_xpb_out[90][607],u_xpb_out[91][607],u_xpb_out[92][607],u_xpb_out[93][607],u_xpb_out[94][607],u_xpb_out[95][607],u_xpb_out[96][607],u_xpb_out[97][607],u_xpb_out[98][607],u_xpb_out[99][607],u_xpb_out[100][607],u_xpb_out[101][607],u_xpb_out[102][607],u_xpb_out[103][607],u_xpb_out[104][607],u_xpb_out[105][607]};

assign col_out_608 = {u_xpb_out[0][608],u_xpb_out[1][608],u_xpb_out[2][608],u_xpb_out[3][608],u_xpb_out[4][608],u_xpb_out[5][608],u_xpb_out[6][608],u_xpb_out[7][608],u_xpb_out[8][608],u_xpb_out[9][608],u_xpb_out[10][608],u_xpb_out[11][608],u_xpb_out[12][608],u_xpb_out[13][608],u_xpb_out[14][608],u_xpb_out[15][608],u_xpb_out[16][608],u_xpb_out[17][608],u_xpb_out[18][608],u_xpb_out[19][608],u_xpb_out[20][608],u_xpb_out[21][608],u_xpb_out[22][608],u_xpb_out[23][608],u_xpb_out[24][608],u_xpb_out[25][608],u_xpb_out[26][608],u_xpb_out[27][608],u_xpb_out[28][608],u_xpb_out[29][608],u_xpb_out[30][608],u_xpb_out[31][608],u_xpb_out[32][608],u_xpb_out[33][608],u_xpb_out[34][608],u_xpb_out[35][608],u_xpb_out[36][608],u_xpb_out[37][608],u_xpb_out[38][608],u_xpb_out[39][608],u_xpb_out[40][608],u_xpb_out[41][608],u_xpb_out[42][608],u_xpb_out[43][608],u_xpb_out[44][608],u_xpb_out[45][608],u_xpb_out[46][608],u_xpb_out[47][608],u_xpb_out[48][608],u_xpb_out[49][608],u_xpb_out[50][608],u_xpb_out[51][608],u_xpb_out[52][608],u_xpb_out[53][608],u_xpb_out[54][608],u_xpb_out[55][608],u_xpb_out[56][608],u_xpb_out[57][608],u_xpb_out[58][608],u_xpb_out[59][608],u_xpb_out[60][608],u_xpb_out[61][608],u_xpb_out[62][608],u_xpb_out[63][608],u_xpb_out[64][608],u_xpb_out[65][608],u_xpb_out[66][608],u_xpb_out[67][608],u_xpb_out[68][608],u_xpb_out[69][608],u_xpb_out[70][608],u_xpb_out[71][608],u_xpb_out[72][608],u_xpb_out[73][608],u_xpb_out[74][608],u_xpb_out[75][608],u_xpb_out[76][608],u_xpb_out[77][608],u_xpb_out[78][608],u_xpb_out[79][608],u_xpb_out[80][608],u_xpb_out[81][608],u_xpb_out[82][608],u_xpb_out[83][608],u_xpb_out[84][608],u_xpb_out[85][608],u_xpb_out[86][608],u_xpb_out[87][608],u_xpb_out[88][608],u_xpb_out[89][608],u_xpb_out[90][608],u_xpb_out[91][608],u_xpb_out[92][608],u_xpb_out[93][608],u_xpb_out[94][608],u_xpb_out[95][608],u_xpb_out[96][608],u_xpb_out[97][608],u_xpb_out[98][608],u_xpb_out[99][608],u_xpb_out[100][608],u_xpb_out[101][608],u_xpb_out[102][608],u_xpb_out[103][608],u_xpb_out[104][608],u_xpb_out[105][608]};

assign col_out_609 = {u_xpb_out[0][609],u_xpb_out[1][609],u_xpb_out[2][609],u_xpb_out[3][609],u_xpb_out[4][609],u_xpb_out[5][609],u_xpb_out[6][609],u_xpb_out[7][609],u_xpb_out[8][609],u_xpb_out[9][609],u_xpb_out[10][609],u_xpb_out[11][609],u_xpb_out[12][609],u_xpb_out[13][609],u_xpb_out[14][609],u_xpb_out[15][609],u_xpb_out[16][609],u_xpb_out[17][609],u_xpb_out[18][609],u_xpb_out[19][609],u_xpb_out[20][609],u_xpb_out[21][609],u_xpb_out[22][609],u_xpb_out[23][609],u_xpb_out[24][609],u_xpb_out[25][609],u_xpb_out[26][609],u_xpb_out[27][609],u_xpb_out[28][609],u_xpb_out[29][609],u_xpb_out[30][609],u_xpb_out[31][609],u_xpb_out[32][609],u_xpb_out[33][609],u_xpb_out[34][609],u_xpb_out[35][609],u_xpb_out[36][609],u_xpb_out[37][609],u_xpb_out[38][609],u_xpb_out[39][609],u_xpb_out[40][609],u_xpb_out[41][609],u_xpb_out[42][609],u_xpb_out[43][609],u_xpb_out[44][609],u_xpb_out[45][609],u_xpb_out[46][609],u_xpb_out[47][609],u_xpb_out[48][609],u_xpb_out[49][609],u_xpb_out[50][609],u_xpb_out[51][609],u_xpb_out[52][609],u_xpb_out[53][609],u_xpb_out[54][609],u_xpb_out[55][609],u_xpb_out[56][609],u_xpb_out[57][609],u_xpb_out[58][609],u_xpb_out[59][609],u_xpb_out[60][609],u_xpb_out[61][609],u_xpb_out[62][609],u_xpb_out[63][609],u_xpb_out[64][609],u_xpb_out[65][609],u_xpb_out[66][609],u_xpb_out[67][609],u_xpb_out[68][609],u_xpb_out[69][609],u_xpb_out[70][609],u_xpb_out[71][609],u_xpb_out[72][609],u_xpb_out[73][609],u_xpb_out[74][609],u_xpb_out[75][609],u_xpb_out[76][609],u_xpb_out[77][609],u_xpb_out[78][609],u_xpb_out[79][609],u_xpb_out[80][609],u_xpb_out[81][609],u_xpb_out[82][609],u_xpb_out[83][609],u_xpb_out[84][609],u_xpb_out[85][609],u_xpb_out[86][609],u_xpb_out[87][609],u_xpb_out[88][609],u_xpb_out[89][609],u_xpb_out[90][609],u_xpb_out[91][609],u_xpb_out[92][609],u_xpb_out[93][609],u_xpb_out[94][609],u_xpb_out[95][609],u_xpb_out[96][609],u_xpb_out[97][609],u_xpb_out[98][609],u_xpb_out[99][609],u_xpb_out[100][609],u_xpb_out[101][609],u_xpb_out[102][609],u_xpb_out[103][609],u_xpb_out[104][609],u_xpb_out[105][609]};

assign col_out_610 = {u_xpb_out[0][610],u_xpb_out[1][610],u_xpb_out[2][610],u_xpb_out[3][610],u_xpb_out[4][610],u_xpb_out[5][610],u_xpb_out[6][610],u_xpb_out[7][610],u_xpb_out[8][610],u_xpb_out[9][610],u_xpb_out[10][610],u_xpb_out[11][610],u_xpb_out[12][610],u_xpb_out[13][610],u_xpb_out[14][610],u_xpb_out[15][610],u_xpb_out[16][610],u_xpb_out[17][610],u_xpb_out[18][610],u_xpb_out[19][610],u_xpb_out[20][610],u_xpb_out[21][610],u_xpb_out[22][610],u_xpb_out[23][610],u_xpb_out[24][610],u_xpb_out[25][610],u_xpb_out[26][610],u_xpb_out[27][610],u_xpb_out[28][610],u_xpb_out[29][610],u_xpb_out[30][610],u_xpb_out[31][610],u_xpb_out[32][610],u_xpb_out[33][610],u_xpb_out[34][610],u_xpb_out[35][610],u_xpb_out[36][610],u_xpb_out[37][610],u_xpb_out[38][610],u_xpb_out[39][610],u_xpb_out[40][610],u_xpb_out[41][610],u_xpb_out[42][610],u_xpb_out[43][610],u_xpb_out[44][610],u_xpb_out[45][610],u_xpb_out[46][610],u_xpb_out[47][610],u_xpb_out[48][610],u_xpb_out[49][610],u_xpb_out[50][610],u_xpb_out[51][610],u_xpb_out[52][610],u_xpb_out[53][610],u_xpb_out[54][610],u_xpb_out[55][610],u_xpb_out[56][610],u_xpb_out[57][610],u_xpb_out[58][610],u_xpb_out[59][610],u_xpb_out[60][610],u_xpb_out[61][610],u_xpb_out[62][610],u_xpb_out[63][610],u_xpb_out[64][610],u_xpb_out[65][610],u_xpb_out[66][610],u_xpb_out[67][610],u_xpb_out[68][610],u_xpb_out[69][610],u_xpb_out[70][610],u_xpb_out[71][610],u_xpb_out[72][610],u_xpb_out[73][610],u_xpb_out[74][610],u_xpb_out[75][610],u_xpb_out[76][610],u_xpb_out[77][610],u_xpb_out[78][610],u_xpb_out[79][610],u_xpb_out[80][610],u_xpb_out[81][610],u_xpb_out[82][610],u_xpb_out[83][610],u_xpb_out[84][610],u_xpb_out[85][610],u_xpb_out[86][610],u_xpb_out[87][610],u_xpb_out[88][610],u_xpb_out[89][610],u_xpb_out[90][610],u_xpb_out[91][610],u_xpb_out[92][610],u_xpb_out[93][610],u_xpb_out[94][610],u_xpb_out[95][610],u_xpb_out[96][610],u_xpb_out[97][610],u_xpb_out[98][610],u_xpb_out[99][610],u_xpb_out[100][610],u_xpb_out[101][610],u_xpb_out[102][610],u_xpb_out[103][610],u_xpb_out[104][610],u_xpb_out[105][610]};

assign col_out_611 = {u_xpb_out[0][611],u_xpb_out[1][611],u_xpb_out[2][611],u_xpb_out[3][611],u_xpb_out[4][611],u_xpb_out[5][611],u_xpb_out[6][611],u_xpb_out[7][611],u_xpb_out[8][611],u_xpb_out[9][611],u_xpb_out[10][611],u_xpb_out[11][611],u_xpb_out[12][611],u_xpb_out[13][611],u_xpb_out[14][611],u_xpb_out[15][611],u_xpb_out[16][611],u_xpb_out[17][611],u_xpb_out[18][611],u_xpb_out[19][611],u_xpb_out[20][611],u_xpb_out[21][611],u_xpb_out[22][611],u_xpb_out[23][611],u_xpb_out[24][611],u_xpb_out[25][611],u_xpb_out[26][611],u_xpb_out[27][611],u_xpb_out[28][611],u_xpb_out[29][611],u_xpb_out[30][611],u_xpb_out[31][611],u_xpb_out[32][611],u_xpb_out[33][611],u_xpb_out[34][611],u_xpb_out[35][611],u_xpb_out[36][611],u_xpb_out[37][611],u_xpb_out[38][611],u_xpb_out[39][611],u_xpb_out[40][611],u_xpb_out[41][611],u_xpb_out[42][611],u_xpb_out[43][611],u_xpb_out[44][611],u_xpb_out[45][611],u_xpb_out[46][611],u_xpb_out[47][611],u_xpb_out[48][611],u_xpb_out[49][611],u_xpb_out[50][611],u_xpb_out[51][611],u_xpb_out[52][611],u_xpb_out[53][611],u_xpb_out[54][611],u_xpb_out[55][611],u_xpb_out[56][611],u_xpb_out[57][611],u_xpb_out[58][611],u_xpb_out[59][611],u_xpb_out[60][611],u_xpb_out[61][611],u_xpb_out[62][611],u_xpb_out[63][611],u_xpb_out[64][611],u_xpb_out[65][611],u_xpb_out[66][611],u_xpb_out[67][611],u_xpb_out[68][611],u_xpb_out[69][611],u_xpb_out[70][611],u_xpb_out[71][611],u_xpb_out[72][611],u_xpb_out[73][611],u_xpb_out[74][611],u_xpb_out[75][611],u_xpb_out[76][611],u_xpb_out[77][611],u_xpb_out[78][611],u_xpb_out[79][611],u_xpb_out[80][611],u_xpb_out[81][611],u_xpb_out[82][611],u_xpb_out[83][611],u_xpb_out[84][611],u_xpb_out[85][611],u_xpb_out[86][611],u_xpb_out[87][611],u_xpb_out[88][611],u_xpb_out[89][611],u_xpb_out[90][611],u_xpb_out[91][611],u_xpb_out[92][611],u_xpb_out[93][611],u_xpb_out[94][611],u_xpb_out[95][611],u_xpb_out[96][611],u_xpb_out[97][611],u_xpb_out[98][611],u_xpb_out[99][611],u_xpb_out[100][611],u_xpb_out[101][611],u_xpb_out[102][611],u_xpb_out[103][611],u_xpb_out[104][611],u_xpb_out[105][611]};

assign col_out_612 = {u_xpb_out[0][612],u_xpb_out[1][612],u_xpb_out[2][612],u_xpb_out[3][612],u_xpb_out[4][612],u_xpb_out[5][612],u_xpb_out[6][612],u_xpb_out[7][612],u_xpb_out[8][612],u_xpb_out[9][612],u_xpb_out[10][612],u_xpb_out[11][612],u_xpb_out[12][612],u_xpb_out[13][612],u_xpb_out[14][612],u_xpb_out[15][612],u_xpb_out[16][612],u_xpb_out[17][612],u_xpb_out[18][612],u_xpb_out[19][612],u_xpb_out[20][612],u_xpb_out[21][612],u_xpb_out[22][612],u_xpb_out[23][612],u_xpb_out[24][612],u_xpb_out[25][612],u_xpb_out[26][612],u_xpb_out[27][612],u_xpb_out[28][612],u_xpb_out[29][612],u_xpb_out[30][612],u_xpb_out[31][612],u_xpb_out[32][612],u_xpb_out[33][612],u_xpb_out[34][612],u_xpb_out[35][612],u_xpb_out[36][612],u_xpb_out[37][612],u_xpb_out[38][612],u_xpb_out[39][612],u_xpb_out[40][612],u_xpb_out[41][612],u_xpb_out[42][612],u_xpb_out[43][612],u_xpb_out[44][612],u_xpb_out[45][612],u_xpb_out[46][612],u_xpb_out[47][612],u_xpb_out[48][612],u_xpb_out[49][612],u_xpb_out[50][612],u_xpb_out[51][612],u_xpb_out[52][612],u_xpb_out[53][612],u_xpb_out[54][612],u_xpb_out[55][612],u_xpb_out[56][612],u_xpb_out[57][612],u_xpb_out[58][612],u_xpb_out[59][612],u_xpb_out[60][612],u_xpb_out[61][612],u_xpb_out[62][612],u_xpb_out[63][612],u_xpb_out[64][612],u_xpb_out[65][612],u_xpb_out[66][612],u_xpb_out[67][612],u_xpb_out[68][612],u_xpb_out[69][612],u_xpb_out[70][612],u_xpb_out[71][612],u_xpb_out[72][612],u_xpb_out[73][612],u_xpb_out[74][612],u_xpb_out[75][612],u_xpb_out[76][612],u_xpb_out[77][612],u_xpb_out[78][612],u_xpb_out[79][612],u_xpb_out[80][612],u_xpb_out[81][612],u_xpb_out[82][612],u_xpb_out[83][612],u_xpb_out[84][612],u_xpb_out[85][612],u_xpb_out[86][612],u_xpb_out[87][612],u_xpb_out[88][612],u_xpb_out[89][612],u_xpb_out[90][612],u_xpb_out[91][612],u_xpb_out[92][612],u_xpb_out[93][612],u_xpb_out[94][612],u_xpb_out[95][612],u_xpb_out[96][612],u_xpb_out[97][612],u_xpb_out[98][612],u_xpb_out[99][612],u_xpb_out[100][612],u_xpb_out[101][612],u_xpb_out[102][612],u_xpb_out[103][612],u_xpb_out[104][612],u_xpb_out[105][612]};

assign col_out_613 = {u_xpb_out[0][613],u_xpb_out[1][613],u_xpb_out[2][613],u_xpb_out[3][613],u_xpb_out[4][613],u_xpb_out[5][613],u_xpb_out[6][613],u_xpb_out[7][613],u_xpb_out[8][613],u_xpb_out[9][613],u_xpb_out[10][613],u_xpb_out[11][613],u_xpb_out[12][613],u_xpb_out[13][613],u_xpb_out[14][613],u_xpb_out[15][613],u_xpb_out[16][613],u_xpb_out[17][613],u_xpb_out[18][613],u_xpb_out[19][613],u_xpb_out[20][613],u_xpb_out[21][613],u_xpb_out[22][613],u_xpb_out[23][613],u_xpb_out[24][613],u_xpb_out[25][613],u_xpb_out[26][613],u_xpb_out[27][613],u_xpb_out[28][613],u_xpb_out[29][613],u_xpb_out[30][613],u_xpb_out[31][613],u_xpb_out[32][613],u_xpb_out[33][613],u_xpb_out[34][613],u_xpb_out[35][613],u_xpb_out[36][613],u_xpb_out[37][613],u_xpb_out[38][613],u_xpb_out[39][613],u_xpb_out[40][613],u_xpb_out[41][613],u_xpb_out[42][613],u_xpb_out[43][613],u_xpb_out[44][613],u_xpb_out[45][613],u_xpb_out[46][613],u_xpb_out[47][613],u_xpb_out[48][613],u_xpb_out[49][613],u_xpb_out[50][613],u_xpb_out[51][613],u_xpb_out[52][613],u_xpb_out[53][613],u_xpb_out[54][613],u_xpb_out[55][613],u_xpb_out[56][613],u_xpb_out[57][613],u_xpb_out[58][613],u_xpb_out[59][613],u_xpb_out[60][613],u_xpb_out[61][613],u_xpb_out[62][613],u_xpb_out[63][613],u_xpb_out[64][613],u_xpb_out[65][613],u_xpb_out[66][613],u_xpb_out[67][613],u_xpb_out[68][613],u_xpb_out[69][613],u_xpb_out[70][613],u_xpb_out[71][613],u_xpb_out[72][613],u_xpb_out[73][613],u_xpb_out[74][613],u_xpb_out[75][613],u_xpb_out[76][613],u_xpb_out[77][613],u_xpb_out[78][613],u_xpb_out[79][613],u_xpb_out[80][613],u_xpb_out[81][613],u_xpb_out[82][613],u_xpb_out[83][613],u_xpb_out[84][613],u_xpb_out[85][613],u_xpb_out[86][613],u_xpb_out[87][613],u_xpb_out[88][613],u_xpb_out[89][613],u_xpb_out[90][613],u_xpb_out[91][613],u_xpb_out[92][613],u_xpb_out[93][613],u_xpb_out[94][613],u_xpb_out[95][613],u_xpb_out[96][613],u_xpb_out[97][613],u_xpb_out[98][613],u_xpb_out[99][613],u_xpb_out[100][613],u_xpb_out[101][613],u_xpb_out[102][613],u_xpb_out[103][613],u_xpb_out[104][613],u_xpb_out[105][613]};

assign col_out_614 = {u_xpb_out[0][614],u_xpb_out[1][614],u_xpb_out[2][614],u_xpb_out[3][614],u_xpb_out[4][614],u_xpb_out[5][614],u_xpb_out[6][614],u_xpb_out[7][614],u_xpb_out[8][614],u_xpb_out[9][614],u_xpb_out[10][614],u_xpb_out[11][614],u_xpb_out[12][614],u_xpb_out[13][614],u_xpb_out[14][614],u_xpb_out[15][614],u_xpb_out[16][614],u_xpb_out[17][614],u_xpb_out[18][614],u_xpb_out[19][614],u_xpb_out[20][614],u_xpb_out[21][614],u_xpb_out[22][614],u_xpb_out[23][614],u_xpb_out[24][614],u_xpb_out[25][614],u_xpb_out[26][614],u_xpb_out[27][614],u_xpb_out[28][614],u_xpb_out[29][614],u_xpb_out[30][614],u_xpb_out[31][614],u_xpb_out[32][614],u_xpb_out[33][614],u_xpb_out[34][614],u_xpb_out[35][614],u_xpb_out[36][614],u_xpb_out[37][614],u_xpb_out[38][614],u_xpb_out[39][614],u_xpb_out[40][614],u_xpb_out[41][614],u_xpb_out[42][614],u_xpb_out[43][614],u_xpb_out[44][614],u_xpb_out[45][614],u_xpb_out[46][614],u_xpb_out[47][614],u_xpb_out[48][614],u_xpb_out[49][614],u_xpb_out[50][614],u_xpb_out[51][614],u_xpb_out[52][614],u_xpb_out[53][614],u_xpb_out[54][614],u_xpb_out[55][614],u_xpb_out[56][614],u_xpb_out[57][614],u_xpb_out[58][614],u_xpb_out[59][614],u_xpb_out[60][614],u_xpb_out[61][614],u_xpb_out[62][614],u_xpb_out[63][614],u_xpb_out[64][614],u_xpb_out[65][614],u_xpb_out[66][614],u_xpb_out[67][614],u_xpb_out[68][614],u_xpb_out[69][614],u_xpb_out[70][614],u_xpb_out[71][614],u_xpb_out[72][614],u_xpb_out[73][614],u_xpb_out[74][614],u_xpb_out[75][614],u_xpb_out[76][614],u_xpb_out[77][614],u_xpb_out[78][614],u_xpb_out[79][614],u_xpb_out[80][614],u_xpb_out[81][614],u_xpb_out[82][614],u_xpb_out[83][614],u_xpb_out[84][614],u_xpb_out[85][614],u_xpb_out[86][614],u_xpb_out[87][614],u_xpb_out[88][614],u_xpb_out[89][614],u_xpb_out[90][614],u_xpb_out[91][614],u_xpb_out[92][614],u_xpb_out[93][614],u_xpb_out[94][614],u_xpb_out[95][614],u_xpb_out[96][614],u_xpb_out[97][614],u_xpb_out[98][614],u_xpb_out[99][614],u_xpb_out[100][614],u_xpb_out[101][614],u_xpb_out[102][614],u_xpb_out[103][614],u_xpb_out[104][614],u_xpb_out[105][614]};

assign col_out_615 = {u_xpb_out[0][615],u_xpb_out[1][615],u_xpb_out[2][615],u_xpb_out[3][615],u_xpb_out[4][615],u_xpb_out[5][615],u_xpb_out[6][615],u_xpb_out[7][615],u_xpb_out[8][615],u_xpb_out[9][615],u_xpb_out[10][615],u_xpb_out[11][615],u_xpb_out[12][615],u_xpb_out[13][615],u_xpb_out[14][615],u_xpb_out[15][615],u_xpb_out[16][615],u_xpb_out[17][615],u_xpb_out[18][615],u_xpb_out[19][615],u_xpb_out[20][615],u_xpb_out[21][615],u_xpb_out[22][615],u_xpb_out[23][615],u_xpb_out[24][615],u_xpb_out[25][615],u_xpb_out[26][615],u_xpb_out[27][615],u_xpb_out[28][615],u_xpb_out[29][615],u_xpb_out[30][615],u_xpb_out[31][615],u_xpb_out[32][615],u_xpb_out[33][615],u_xpb_out[34][615],u_xpb_out[35][615],u_xpb_out[36][615],u_xpb_out[37][615],u_xpb_out[38][615],u_xpb_out[39][615],u_xpb_out[40][615],u_xpb_out[41][615],u_xpb_out[42][615],u_xpb_out[43][615],u_xpb_out[44][615],u_xpb_out[45][615],u_xpb_out[46][615],u_xpb_out[47][615],u_xpb_out[48][615],u_xpb_out[49][615],u_xpb_out[50][615],u_xpb_out[51][615],u_xpb_out[52][615],u_xpb_out[53][615],u_xpb_out[54][615],u_xpb_out[55][615],u_xpb_out[56][615],u_xpb_out[57][615],u_xpb_out[58][615],u_xpb_out[59][615],u_xpb_out[60][615],u_xpb_out[61][615],u_xpb_out[62][615],u_xpb_out[63][615],u_xpb_out[64][615],u_xpb_out[65][615],u_xpb_out[66][615],u_xpb_out[67][615],u_xpb_out[68][615],u_xpb_out[69][615],u_xpb_out[70][615],u_xpb_out[71][615],u_xpb_out[72][615],u_xpb_out[73][615],u_xpb_out[74][615],u_xpb_out[75][615],u_xpb_out[76][615],u_xpb_out[77][615],u_xpb_out[78][615],u_xpb_out[79][615],u_xpb_out[80][615],u_xpb_out[81][615],u_xpb_out[82][615],u_xpb_out[83][615],u_xpb_out[84][615],u_xpb_out[85][615],u_xpb_out[86][615],u_xpb_out[87][615],u_xpb_out[88][615],u_xpb_out[89][615],u_xpb_out[90][615],u_xpb_out[91][615],u_xpb_out[92][615],u_xpb_out[93][615],u_xpb_out[94][615],u_xpb_out[95][615],u_xpb_out[96][615],u_xpb_out[97][615],u_xpb_out[98][615],u_xpb_out[99][615],u_xpb_out[100][615],u_xpb_out[101][615],u_xpb_out[102][615],u_xpb_out[103][615],u_xpb_out[104][615],u_xpb_out[105][615]};

assign col_out_616 = {u_xpb_out[0][616],u_xpb_out[1][616],u_xpb_out[2][616],u_xpb_out[3][616],u_xpb_out[4][616],u_xpb_out[5][616],u_xpb_out[6][616],u_xpb_out[7][616],u_xpb_out[8][616],u_xpb_out[9][616],u_xpb_out[10][616],u_xpb_out[11][616],u_xpb_out[12][616],u_xpb_out[13][616],u_xpb_out[14][616],u_xpb_out[15][616],u_xpb_out[16][616],u_xpb_out[17][616],u_xpb_out[18][616],u_xpb_out[19][616],u_xpb_out[20][616],u_xpb_out[21][616],u_xpb_out[22][616],u_xpb_out[23][616],u_xpb_out[24][616],u_xpb_out[25][616],u_xpb_out[26][616],u_xpb_out[27][616],u_xpb_out[28][616],u_xpb_out[29][616],u_xpb_out[30][616],u_xpb_out[31][616],u_xpb_out[32][616],u_xpb_out[33][616],u_xpb_out[34][616],u_xpb_out[35][616],u_xpb_out[36][616],u_xpb_out[37][616],u_xpb_out[38][616],u_xpb_out[39][616],u_xpb_out[40][616],u_xpb_out[41][616],u_xpb_out[42][616],u_xpb_out[43][616],u_xpb_out[44][616],u_xpb_out[45][616],u_xpb_out[46][616],u_xpb_out[47][616],u_xpb_out[48][616],u_xpb_out[49][616],u_xpb_out[50][616],u_xpb_out[51][616],u_xpb_out[52][616],u_xpb_out[53][616],u_xpb_out[54][616],u_xpb_out[55][616],u_xpb_out[56][616],u_xpb_out[57][616],u_xpb_out[58][616],u_xpb_out[59][616],u_xpb_out[60][616],u_xpb_out[61][616],u_xpb_out[62][616],u_xpb_out[63][616],u_xpb_out[64][616],u_xpb_out[65][616],u_xpb_out[66][616],u_xpb_out[67][616],u_xpb_out[68][616],u_xpb_out[69][616],u_xpb_out[70][616],u_xpb_out[71][616],u_xpb_out[72][616],u_xpb_out[73][616],u_xpb_out[74][616],u_xpb_out[75][616],u_xpb_out[76][616],u_xpb_out[77][616],u_xpb_out[78][616],u_xpb_out[79][616],u_xpb_out[80][616],u_xpb_out[81][616],u_xpb_out[82][616],u_xpb_out[83][616],u_xpb_out[84][616],u_xpb_out[85][616],u_xpb_out[86][616],u_xpb_out[87][616],u_xpb_out[88][616],u_xpb_out[89][616],u_xpb_out[90][616],u_xpb_out[91][616],u_xpb_out[92][616],u_xpb_out[93][616],u_xpb_out[94][616],u_xpb_out[95][616],u_xpb_out[96][616],u_xpb_out[97][616],u_xpb_out[98][616],u_xpb_out[99][616],u_xpb_out[100][616],u_xpb_out[101][616],u_xpb_out[102][616],u_xpb_out[103][616],u_xpb_out[104][616],u_xpb_out[105][616]};

assign col_out_617 = {u_xpb_out[0][617],u_xpb_out[1][617],u_xpb_out[2][617],u_xpb_out[3][617],u_xpb_out[4][617],u_xpb_out[5][617],u_xpb_out[6][617],u_xpb_out[7][617],u_xpb_out[8][617],u_xpb_out[9][617],u_xpb_out[10][617],u_xpb_out[11][617],u_xpb_out[12][617],u_xpb_out[13][617],u_xpb_out[14][617],u_xpb_out[15][617],u_xpb_out[16][617],u_xpb_out[17][617],u_xpb_out[18][617],u_xpb_out[19][617],u_xpb_out[20][617],u_xpb_out[21][617],u_xpb_out[22][617],u_xpb_out[23][617],u_xpb_out[24][617],u_xpb_out[25][617],u_xpb_out[26][617],u_xpb_out[27][617],u_xpb_out[28][617],u_xpb_out[29][617],u_xpb_out[30][617],u_xpb_out[31][617],u_xpb_out[32][617],u_xpb_out[33][617],u_xpb_out[34][617],u_xpb_out[35][617],u_xpb_out[36][617],u_xpb_out[37][617],u_xpb_out[38][617],u_xpb_out[39][617],u_xpb_out[40][617],u_xpb_out[41][617],u_xpb_out[42][617],u_xpb_out[43][617],u_xpb_out[44][617],u_xpb_out[45][617],u_xpb_out[46][617],u_xpb_out[47][617],u_xpb_out[48][617],u_xpb_out[49][617],u_xpb_out[50][617],u_xpb_out[51][617],u_xpb_out[52][617],u_xpb_out[53][617],u_xpb_out[54][617],u_xpb_out[55][617],u_xpb_out[56][617],u_xpb_out[57][617],u_xpb_out[58][617],u_xpb_out[59][617],u_xpb_out[60][617],u_xpb_out[61][617],u_xpb_out[62][617],u_xpb_out[63][617],u_xpb_out[64][617],u_xpb_out[65][617],u_xpb_out[66][617],u_xpb_out[67][617],u_xpb_out[68][617],u_xpb_out[69][617],u_xpb_out[70][617],u_xpb_out[71][617],u_xpb_out[72][617],u_xpb_out[73][617],u_xpb_out[74][617],u_xpb_out[75][617],u_xpb_out[76][617],u_xpb_out[77][617],u_xpb_out[78][617],u_xpb_out[79][617],u_xpb_out[80][617],u_xpb_out[81][617],u_xpb_out[82][617],u_xpb_out[83][617],u_xpb_out[84][617],u_xpb_out[85][617],u_xpb_out[86][617],u_xpb_out[87][617],u_xpb_out[88][617],u_xpb_out[89][617],u_xpb_out[90][617],u_xpb_out[91][617],u_xpb_out[92][617],u_xpb_out[93][617],u_xpb_out[94][617],u_xpb_out[95][617],u_xpb_out[96][617],u_xpb_out[97][617],u_xpb_out[98][617],u_xpb_out[99][617],u_xpb_out[100][617],u_xpb_out[101][617],u_xpb_out[102][617],u_xpb_out[103][617],u_xpb_out[104][617],u_xpb_out[105][617]};

assign col_out_618 = {u_xpb_out[0][618],u_xpb_out[1][618],u_xpb_out[2][618],u_xpb_out[3][618],u_xpb_out[4][618],u_xpb_out[5][618],u_xpb_out[6][618],u_xpb_out[7][618],u_xpb_out[8][618],u_xpb_out[9][618],u_xpb_out[10][618],u_xpb_out[11][618],u_xpb_out[12][618],u_xpb_out[13][618],u_xpb_out[14][618],u_xpb_out[15][618],u_xpb_out[16][618],u_xpb_out[17][618],u_xpb_out[18][618],u_xpb_out[19][618],u_xpb_out[20][618],u_xpb_out[21][618],u_xpb_out[22][618],u_xpb_out[23][618],u_xpb_out[24][618],u_xpb_out[25][618],u_xpb_out[26][618],u_xpb_out[27][618],u_xpb_out[28][618],u_xpb_out[29][618],u_xpb_out[30][618],u_xpb_out[31][618],u_xpb_out[32][618],u_xpb_out[33][618],u_xpb_out[34][618],u_xpb_out[35][618],u_xpb_out[36][618],u_xpb_out[37][618],u_xpb_out[38][618],u_xpb_out[39][618],u_xpb_out[40][618],u_xpb_out[41][618],u_xpb_out[42][618],u_xpb_out[43][618],u_xpb_out[44][618],u_xpb_out[45][618],u_xpb_out[46][618],u_xpb_out[47][618],u_xpb_out[48][618],u_xpb_out[49][618],u_xpb_out[50][618],u_xpb_out[51][618],u_xpb_out[52][618],u_xpb_out[53][618],u_xpb_out[54][618],u_xpb_out[55][618],u_xpb_out[56][618],u_xpb_out[57][618],u_xpb_out[58][618],u_xpb_out[59][618],u_xpb_out[60][618],u_xpb_out[61][618],u_xpb_out[62][618],u_xpb_out[63][618],u_xpb_out[64][618],u_xpb_out[65][618],u_xpb_out[66][618],u_xpb_out[67][618],u_xpb_out[68][618],u_xpb_out[69][618],u_xpb_out[70][618],u_xpb_out[71][618],u_xpb_out[72][618],u_xpb_out[73][618],u_xpb_out[74][618],u_xpb_out[75][618],u_xpb_out[76][618],u_xpb_out[77][618],u_xpb_out[78][618],u_xpb_out[79][618],u_xpb_out[80][618],u_xpb_out[81][618],u_xpb_out[82][618],u_xpb_out[83][618],u_xpb_out[84][618],u_xpb_out[85][618],u_xpb_out[86][618],u_xpb_out[87][618],u_xpb_out[88][618],u_xpb_out[89][618],u_xpb_out[90][618],u_xpb_out[91][618],u_xpb_out[92][618],u_xpb_out[93][618],u_xpb_out[94][618],u_xpb_out[95][618],u_xpb_out[96][618],u_xpb_out[97][618],u_xpb_out[98][618],u_xpb_out[99][618],u_xpb_out[100][618],u_xpb_out[101][618],u_xpb_out[102][618],u_xpb_out[103][618],u_xpb_out[104][618],u_xpb_out[105][618]};

assign col_out_619 = {u_xpb_out[0][619],u_xpb_out[1][619],u_xpb_out[2][619],u_xpb_out[3][619],u_xpb_out[4][619],u_xpb_out[5][619],u_xpb_out[6][619],u_xpb_out[7][619],u_xpb_out[8][619],u_xpb_out[9][619],u_xpb_out[10][619],u_xpb_out[11][619],u_xpb_out[12][619],u_xpb_out[13][619],u_xpb_out[14][619],u_xpb_out[15][619],u_xpb_out[16][619],u_xpb_out[17][619],u_xpb_out[18][619],u_xpb_out[19][619],u_xpb_out[20][619],u_xpb_out[21][619],u_xpb_out[22][619],u_xpb_out[23][619],u_xpb_out[24][619],u_xpb_out[25][619],u_xpb_out[26][619],u_xpb_out[27][619],u_xpb_out[28][619],u_xpb_out[29][619],u_xpb_out[30][619],u_xpb_out[31][619],u_xpb_out[32][619],u_xpb_out[33][619],u_xpb_out[34][619],u_xpb_out[35][619],u_xpb_out[36][619],u_xpb_out[37][619],u_xpb_out[38][619],u_xpb_out[39][619],u_xpb_out[40][619],u_xpb_out[41][619],u_xpb_out[42][619],u_xpb_out[43][619],u_xpb_out[44][619],u_xpb_out[45][619],u_xpb_out[46][619],u_xpb_out[47][619],u_xpb_out[48][619],u_xpb_out[49][619],u_xpb_out[50][619],u_xpb_out[51][619],u_xpb_out[52][619],u_xpb_out[53][619],u_xpb_out[54][619],u_xpb_out[55][619],u_xpb_out[56][619],u_xpb_out[57][619],u_xpb_out[58][619],u_xpb_out[59][619],u_xpb_out[60][619],u_xpb_out[61][619],u_xpb_out[62][619],u_xpb_out[63][619],u_xpb_out[64][619],u_xpb_out[65][619],u_xpb_out[66][619],u_xpb_out[67][619],u_xpb_out[68][619],u_xpb_out[69][619],u_xpb_out[70][619],u_xpb_out[71][619],u_xpb_out[72][619],u_xpb_out[73][619],u_xpb_out[74][619],u_xpb_out[75][619],u_xpb_out[76][619],u_xpb_out[77][619],u_xpb_out[78][619],u_xpb_out[79][619],u_xpb_out[80][619],u_xpb_out[81][619],u_xpb_out[82][619],u_xpb_out[83][619],u_xpb_out[84][619],u_xpb_out[85][619],u_xpb_out[86][619],u_xpb_out[87][619],u_xpb_out[88][619],u_xpb_out[89][619],u_xpb_out[90][619],u_xpb_out[91][619],u_xpb_out[92][619],u_xpb_out[93][619],u_xpb_out[94][619],u_xpb_out[95][619],u_xpb_out[96][619],u_xpb_out[97][619],u_xpb_out[98][619],u_xpb_out[99][619],u_xpb_out[100][619],u_xpb_out[101][619],u_xpb_out[102][619],u_xpb_out[103][619],u_xpb_out[104][619],u_xpb_out[105][619]};

assign col_out_620 = {u_xpb_out[0][620],u_xpb_out[1][620],u_xpb_out[2][620],u_xpb_out[3][620],u_xpb_out[4][620],u_xpb_out[5][620],u_xpb_out[6][620],u_xpb_out[7][620],u_xpb_out[8][620],u_xpb_out[9][620],u_xpb_out[10][620],u_xpb_out[11][620],u_xpb_out[12][620],u_xpb_out[13][620],u_xpb_out[14][620],u_xpb_out[15][620],u_xpb_out[16][620],u_xpb_out[17][620],u_xpb_out[18][620],u_xpb_out[19][620],u_xpb_out[20][620],u_xpb_out[21][620],u_xpb_out[22][620],u_xpb_out[23][620],u_xpb_out[24][620],u_xpb_out[25][620],u_xpb_out[26][620],u_xpb_out[27][620],u_xpb_out[28][620],u_xpb_out[29][620],u_xpb_out[30][620],u_xpb_out[31][620],u_xpb_out[32][620],u_xpb_out[33][620],u_xpb_out[34][620],u_xpb_out[35][620],u_xpb_out[36][620],u_xpb_out[37][620],u_xpb_out[38][620],u_xpb_out[39][620],u_xpb_out[40][620],u_xpb_out[41][620],u_xpb_out[42][620],u_xpb_out[43][620],u_xpb_out[44][620],u_xpb_out[45][620],u_xpb_out[46][620],u_xpb_out[47][620],u_xpb_out[48][620],u_xpb_out[49][620],u_xpb_out[50][620],u_xpb_out[51][620],u_xpb_out[52][620],u_xpb_out[53][620],u_xpb_out[54][620],u_xpb_out[55][620],u_xpb_out[56][620],u_xpb_out[57][620],u_xpb_out[58][620],u_xpb_out[59][620],u_xpb_out[60][620],u_xpb_out[61][620],u_xpb_out[62][620],u_xpb_out[63][620],u_xpb_out[64][620],u_xpb_out[65][620],u_xpb_out[66][620],u_xpb_out[67][620],u_xpb_out[68][620],u_xpb_out[69][620],u_xpb_out[70][620],u_xpb_out[71][620],u_xpb_out[72][620],u_xpb_out[73][620],u_xpb_out[74][620],u_xpb_out[75][620],u_xpb_out[76][620],u_xpb_out[77][620],u_xpb_out[78][620],u_xpb_out[79][620],u_xpb_out[80][620],u_xpb_out[81][620],u_xpb_out[82][620],u_xpb_out[83][620],u_xpb_out[84][620],u_xpb_out[85][620],u_xpb_out[86][620],u_xpb_out[87][620],u_xpb_out[88][620],u_xpb_out[89][620],u_xpb_out[90][620],u_xpb_out[91][620],u_xpb_out[92][620],u_xpb_out[93][620],u_xpb_out[94][620],u_xpb_out[95][620],u_xpb_out[96][620],u_xpb_out[97][620],u_xpb_out[98][620],u_xpb_out[99][620],u_xpb_out[100][620],u_xpb_out[101][620],u_xpb_out[102][620],u_xpb_out[103][620],u_xpb_out[104][620],u_xpb_out[105][620]};

assign col_out_621 = {u_xpb_out[0][621],u_xpb_out[1][621],u_xpb_out[2][621],u_xpb_out[3][621],u_xpb_out[4][621],u_xpb_out[5][621],u_xpb_out[6][621],u_xpb_out[7][621],u_xpb_out[8][621],u_xpb_out[9][621],u_xpb_out[10][621],u_xpb_out[11][621],u_xpb_out[12][621],u_xpb_out[13][621],u_xpb_out[14][621],u_xpb_out[15][621],u_xpb_out[16][621],u_xpb_out[17][621],u_xpb_out[18][621],u_xpb_out[19][621],u_xpb_out[20][621],u_xpb_out[21][621],u_xpb_out[22][621],u_xpb_out[23][621],u_xpb_out[24][621],u_xpb_out[25][621],u_xpb_out[26][621],u_xpb_out[27][621],u_xpb_out[28][621],u_xpb_out[29][621],u_xpb_out[30][621],u_xpb_out[31][621],u_xpb_out[32][621],u_xpb_out[33][621],u_xpb_out[34][621],u_xpb_out[35][621],u_xpb_out[36][621],u_xpb_out[37][621],u_xpb_out[38][621],u_xpb_out[39][621],u_xpb_out[40][621],u_xpb_out[41][621],u_xpb_out[42][621],u_xpb_out[43][621],u_xpb_out[44][621],u_xpb_out[45][621],u_xpb_out[46][621],u_xpb_out[47][621],u_xpb_out[48][621],u_xpb_out[49][621],u_xpb_out[50][621],u_xpb_out[51][621],u_xpb_out[52][621],u_xpb_out[53][621],u_xpb_out[54][621],u_xpb_out[55][621],u_xpb_out[56][621],u_xpb_out[57][621],u_xpb_out[58][621],u_xpb_out[59][621],u_xpb_out[60][621],u_xpb_out[61][621],u_xpb_out[62][621],u_xpb_out[63][621],u_xpb_out[64][621],u_xpb_out[65][621],u_xpb_out[66][621],u_xpb_out[67][621],u_xpb_out[68][621],u_xpb_out[69][621],u_xpb_out[70][621],u_xpb_out[71][621],u_xpb_out[72][621],u_xpb_out[73][621],u_xpb_out[74][621],u_xpb_out[75][621],u_xpb_out[76][621],u_xpb_out[77][621],u_xpb_out[78][621],u_xpb_out[79][621],u_xpb_out[80][621],u_xpb_out[81][621],u_xpb_out[82][621],u_xpb_out[83][621],u_xpb_out[84][621],u_xpb_out[85][621],u_xpb_out[86][621],u_xpb_out[87][621],u_xpb_out[88][621],u_xpb_out[89][621],u_xpb_out[90][621],u_xpb_out[91][621],u_xpb_out[92][621],u_xpb_out[93][621],u_xpb_out[94][621],u_xpb_out[95][621],u_xpb_out[96][621],u_xpb_out[97][621],u_xpb_out[98][621],u_xpb_out[99][621],u_xpb_out[100][621],u_xpb_out[101][621],u_xpb_out[102][621],u_xpb_out[103][621],u_xpb_out[104][621],u_xpb_out[105][621]};

assign col_out_622 = {u_xpb_out[0][622],u_xpb_out[1][622],u_xpb_out[2][622],u_xpb_out[3][622],u_xpb_out[4][622],u_xpb_out[5][622],u_xpb_out[6][622],u_xpb_out[7][622],u_xpb_out[8][622],u_xpb_out[9][622],u_xpb_out[10][622],u_xpb_out[11][622],u_xpb_out[12][622],u_xpb_out[13][622],u_xpb_out[14][622],u_xpb_out[15][622],u_xpb_out[16][622],u_xpb_out[17][622],u_xpb_out[18][622],u_xpb_out[19][622],u_xpb_out[20][622],u_xpb_out[21][622],u_xpb_out[22][622],u_xpb_out[23][622],u_xpb_out[24][622],u_xpb_out[25][622],u_xpb_out[26][622],u_xpb_out[27][622],u_xpb_out[28][622],u_xpb_out[29][622],u_xpb_out[30][622],u_xpb_out[31][622],u_xpb_out[32][622],u_xpb_out[33][622],u_xpb_out[34][622],u_xpb_out[35][622],u_xpb_out[36][622],u_xpb_out[37][622],u_xpb_out[38][622],u_xpb_out[39][622],u_xpb_out[40][622],u_xpb_out[41][622],u_xpb_out[42][622],u_xpb_out[43][622],u_xpb_out[44][622],u_xpb_out[45][622],u_xpb_out[46][622],u_xpb_out[47][622],u_xpb_out[48][622],u_xpb_out[49][622],u_xpb_out[50][622],u_xpb_out[51][622],u_xpb_out[52][622],u_xpb_out[53][622],u_xpb_out[54][622],u_xpb_out[55][622],u_xpb_out[56][622],u_xpb_out[57][622],u_xpb_out[58][622],u_xpb_out[59][622],u_xpb_out[60][622],u_xpb_out[61][622],u_xpb_out[62][622],u_xpb_out[63][622],u_xpb_out[64][622],u_xpb_out[65][622],u_xpb_out[66][622],u_xpb_out[67][622],u_xpb_out[68][622],u_xpb_out[69][622],u_xpb_out[70][622],u_xpb_out[71][622],u_xpb_out[72][622],u_xpb_out[73][622],u_xpb_out[74][622],u_xpb_out[75][622],u_xpb_out[76][622],u_xpb_out[77][622],u_xpb_out[78][622],u_xpb_out[79][622],u_xpb_out[80][622],u_xpb_out[81][622],u_xpb_out[82][622],u_xpb_out[83][622],u_xpb_out[84][622],u_xpb_out[85][622],u_xpb_out[86][622],u_xpb_out[87][622],u_xpb_out[88][622],u_xpb_out[89][622],u_xpb_out[90][622],u_xpb_out[91][622],u_xpb_out[92][622],u_xpb_out[93][622],u_xpb_out[94][622],u_xpb_out[95][622],u_xpb_out[96][622],u_xpb_out[97][622],u_xpb_out[98][622],u_xpb_out[99][622],u_xpb_out[100][622],u_xpb_out[101][622],u_xpb_out[102][622],u_xpb_out[103][622],u_xpb_out[104][622],u_xpb_out[105][622]};

assign col_out_623 = {u_xpb_out[0][623],u_xpb_out[1][623],u_xpb_out[2][623],u_xpb_out[3][623],u_xpb_out[4][623],u_xpb_out[5][623],u_xpb_out[6][623],u_xpb_out[7][623],u_xpb_out[8][623],u_xpb_out[9][623],u_xpb_out[10][623],u_xpb_out[11][623],u_xpb_out[12][623],u_xpb_out[13][623],u_xpb_out[14][623],u_xpb_out[15][623],u_xpb_out[16][623],u_xpb_out[17][623],u_xpb_out[18][623],u_xpb_out[19][623],u_xpb_out[20][623],u_xpb_out[21][623],u_xpb_out[22][623],u_xpb_out[23][623],u_xpb_out[24][623],u_xpb_out[25][623],u_xpb_out[26][623],u_xpb_out[27][623],u_xpb_out[28][623],u_xpb_out[29][623],u_xpb_out[30][623],u_xpb_out[31][623],u_xpb_out[32][623],u_xpb_out[33][623],u_xpb_out[34][623],u_xpb_out[35][623],u_xpb_out[36][623],u_xpb_out[37][623],u_xpb_out[38][623],u_xpb_out[39][623],u_xpb_out[40][623],u_xpb_out[41][623],u_xpb_out[42][623],u_xpb_out[43][623],u_xpb_out[44][623],u_xpb_out[45][623],u_xpb_out[46][623],u_xpb_out[47][623],u_xpb_out[48][623],u_xpb_out[49][623],u_xpb_out[50][623],u_xpb_out[51][623],u_xpb_out[52][623],u_xpb_out[53][623],u_xpb_out[54][623],u_xpb_out[55][623],u_xpb_out[56][623],u_xpb_out[57][623],u_xpb_out[58][623],u_xpb_out[59][623],u_xpb_out[60][623],u_xpb_out[61][623],u_xpb_out[62][623],u_xpb_out[63][623],u_xpb_out[64][623],u_xpb_out[65][623],u_xpb_out[66][623],u_xpb_out[67][623],u_xpb_out[68][623],u_xpb_out[69][623],u_xpb_out[70][623],u_xpb_out[71][623],u_xpb_out[72][623],u_xpb_out[73][623],u_xpb_out[74][623],u_xpb_out[75][623],u_xpb_out[76][623],u_xpb_out[77][623],u_xpb_out[78][623],u_xpb_out[79][623],u_xpb_out[80][623],u_xpb_out[81][623],u_xpb_out[82][623],u_xpb_out[83][623],u_xpb_out[84][623],u_xpb_out[85][623],u_xpb_out[86][623],u_xpb_out[87][623],u_xpb_out[88][623],u_xpb_out[89][623],u_xpb_out[90][623],u_xpb_out[91][623],u_xpb_out[92][623],u_xpb_out[93][623],u_xpb_out[94][623],u_xpb_out[95][623],u_xpb_out[96][623],u_xpb_out[97][623],u_xpb_out[98][623],u_xpb_out[99][623],u_xpb_out[100][623],u_xpb_out[101][623],u_xpb_out[102][623],u_xpb_out[103][623],u_xpb_out[104][623],u_xpb_out[105][623]};

assign col_out_624 = {u_xpb_out[0][624],u_xpb_out[1][624],u_xpb_out[2][624],u_xpb_out[3][624],u_xpb_out[4][624],u_xpb_out[5][624],u_xpb_out[6][624],u_xpb_out[7][624],u_xpb_out[8][624],u_xpb_out[9][624],u_xpb_out[10][624],u_xpb_out[11][624],u_xpb_out[12][624],u_xpb_out[13][624],u_xpb_out[14][624],u_xpb_out[15][624],u_xpb_out[16][624],u_xpb_out[17][624],u_xpb_out[18][624],u_xpb_out[19][624],u_xpb_out[20][624],u_xpb_out[21][624],u_xpb_out[22][624],u_xpb_out[23][624],u_xpb_out[24][624],u_xpb_out[25][624],u_xpb_out[26][624],u_xpb_out[27][624],u_xpb_out[28][624],u_xpb_out[29][624],u_xpb_out[30][624],u_xpb_out[31][624],u_xpb_out[32][624],u_xpb_out[33][624],u_xpb_out[34][624],u_xpb_out[35][624],u_xpb_out[36][624],u_xpb_out[37][624],u_xpb_out[38][624],u_xpb_out[39][624],u_xpb_out[40][624],u_xpb_out[41][624],u_xpb_out[42][624],u_xpb_out[43][624],u_xpb_out[44][624],u_xpb_out[45][624],u_xpb_out[46][624],u_xpb_out[47][624],u_xpb_out[48][624],u_xpb_out[49][624],u_xpb_out[50][624],u_xpb_out[51][624],u_xpb_out[52][624],u_xpb_out[53][624],u_xpb_out[54][624],u_xpb_out[55][624],u_xpb_out[56][624],u_xpb_out[57][624],u_xpb_out[58][624],u_xpb_out[59][624],u_xpb_out[60][624],u_xpb_out[61][624],u_xpb_out[62][624],u_xpb_out[63][624],u_xpb_out[64][624],u_xpb_out[65][624],u_xpb_out[66][624],u_xpb_out[67][624],u_xpb_out[68][624],u_xpb_out[69][624],u_xpb_out[70][624],u_xpb_out[71][624],u_xpb_out[72][624],u_xpb_out[73][624],u_xpb_out[74][624],u_xpb_out[75][624],u_xpb_out[76][624],u_xpb_out[77][624],u_xpb_out[78][624],u_xpb_out[79][624],u_xpb_out[80][624],u_xpb_out[81][624],u_xpb_out[82][624],u_xpb_out[83][624],u_xpb_out[84][624],u_xpb_out[85][624],u_xpb_out[86][624],u_xpb_out[87][624],u_xpb_out[88][624],u_xpb_out[89][624],u_xpb_out[90][624],u_xpb_out[91][624],u_xpb_out[92][624],u_xpb_out[93][624],u_xpb_out[94][624],u_xpb_out[95][624],u_xpb_out[96][624],u_xpb_out[97][624],u_xpb_out[98][624],u_xpb_out[99][624],u_xpb_out[100][624],u_xpb_out[101][624],u_xpb_out[102][624],u_xpb_out[103][624],u_xpb_out[104][624],u_xpb_out[105][624]};

assign col_out_625 = {u_xpb_out[0][625],u_xpb_out[1][625],u_xpb_out[2][625],u_xpb_out[3][625],u_xpb_out[4][625],u_xpb_out[5][625],u_xpb_out[6][625],u_xpb_out[7][625],u_xpb_out[8][625],u_xpb_out[9][625],u_xpb_out[10][625],u_xpb_out[11][625],u_xpb_out[12][625],u_xpb_out[13][625],u_xpb_out[14][625],u_xpb_out[15][625],u_xpb_out[16][625],u_xpb_out[17][625],u_xpb_out[18][625],u_xpb_out[19][625],u_xpb_out[20][625],u_xpb_out[21][625],u_xpb_out[22][625],u_xpb_out[23][625],u_xpb_out[24][625],u_xpb_out[25][625],u_xpb_out[26][625],u_xpb_out[27][625],u_xpb_out[28][625],u_xpb_out[29][625],u_xpb_out[30][625],u_xpb_out[31][625],u_xpb_out[32][625],u_xpb_out[33][625],u_xpb_out[34][625],u_xpb_out[35][625],u_xpb_out[36][625],u_xpb_out[37][625],u_xpb_out[38][625],u_xpb_out[39][625],u_xpb_out[40][625],u_xpb_out[41][625],u_xpb_out[42][625],u_xpb_out[43][625],u_xpb_out[44][625],u_xpb_out[45][625],u_xpb_out[46][625],u_xpb_out[47][625],u_xpb_out[48][625],u_xpb_out[49][625],u_xpb_out[50][625],u_xpb_out[51][625],u_xpb_out[52][625],u_xpb_out[53][625],u_xpb_out[54][625],u_xpb_out[55][625],u_xpb_out[56][625],u_xpb_out[57][625],u_xpb_out[58][625],u_xpb_out[59][625],u_xpb_out[60][625],u_xpb_out[61][625],u_xpb_out[62][625],u_xpb_out[63][625],u_xpb_out[64][625],u_xpb_out[65][625],u_xpb_out[66][625],u_xpb_out[67][625],u_xpb_out[68][625],u_xpb_out[69][625],u_xpb_out[70][625],u_xpb_out[71][625],u_xpb_out[72][625],u_xpb_out[73][625],u_xpb_out[74][625],u_xpb_out[75][625],u_xpb_out[76][625],u_xpb_out[77][625],u_xpb_out[78][625],u_xpb_out[79][625],u_xpb_out[80][625],u_xpb_out[81][625],u_xpb_out[82][625],u_xpb_out[83][625],u_xpb_out[84][625],u_xpb_out[85][625],u_xpb_out[86][625],u_xpb_out[87][625],u_xpb_out[88][625],u_xpb_out[89][625],u_xpb_out[90][625],u_xpb_out[91][625],u_xpb_out[92][625],u_xpb_out[93][625],u_xpb_out[94][625],u_xpb_out[95][625],u_xpb_out[96][625],u_xpb_out[97][625],u_xpb_out[98][625],u_xpb_out[99][625],u_xpb_out[100][625],u_xpb_out[101][625],u_xpb_out[102][625],u_xpb_out[103][625],u_xpb_out[104][625],u_xpb_out[105][625]};

assign col_out_626 = {u_xpb_out[0][626],u_xpb_out[1][626],u_xpb_out[2][626],u_xpb_out[3][626],u_xpb_out[4][626],u_xpb_out[5][626],u_xpb_out[6][626],u_xpb_out[7][626],u_xpb_out[8][626],u_xpb_out[9][626],u_xpb_out[10][626],u_xpb_out[11][626],u_xpb_out[12][626],u_xpb_out[13][626],u_xpb_out[14][626],u_xpb_out[15][626],u_xpb_out[16][626],u_xpb_out[17][626],u_xpb_out[18][626],u_xpb_out[19][626],u_xpb_out[20][626],u_xpb_out[21][626],u_xpb_out[22][626],u_xpb_out[23][626],u_xpb_out[24][626],u_xpb_out[25][626],u_xpb_out[26][626],u_xpb_out[27][626],u_xpb_out[28][626],u_xpb_out[29][626],u_xpb_out[30][626],u_xpb_out[31][626],u_xpb_out[32][626],u_xpb_out[33][626],u_xpb_out[34][626],u_xpb_out[35][626],u_xpb_out[36][626],u_xpb_out[37][626],u_xpb_out[38][626],u_xpb_out[39][626],u_xpb_out[40][626],u_xpb_out[41][626],u_xpb_out[42][626],u_xpb_out[43][626],u_xpb_out[44][626],u_xpb_out[45][626],u_xpb_out[46][626],u_xpb_out[47][626],u_xpb_out[48][626],u_xpb_out[49][626],u_xpb_out[50][626],u_xpb_out[51][626],u_xpb_out[52][626],u_xpb_out[53][626],u_xpb_out[54][626],u_xpb_out[55][626],u_xpb_out[56][626],u_xpb_out[57][626],u_xpb_out[58][626],u_xpb_out[59][626],u_xpb_out[60][626],u_xpb_out[61][626],u_xpb_out[62][626],u_xpb_out[63][626],u_xpb_out[64][626],u_xpb_out[65][626],u_xpb_out[66][626],u_xpb_out[67][626],u_xpb_out[68][626],u_xpb_out[69][626],u_xpb_out[70][626],u_xpb_out[71][626],u_xpb_out[72][626],u_xpb_out[73][626],u_xpb_out[74][626],u_xpb_out[75][626],u_xpb_out[76][626],u_xpb_out[77][626],u_xpb_out[78][626],u_xpb_out[79][626],u_xpb_out[80][626],u_xpb_out[81][626],u_xpb_out[82][626],u_xpb_out[83][626],u_xpb_out[84][626],u_xpb_out[85][626],u_xpb_out[86][626],u_xpb_out[87][626],u_xpb_out[88][626],u_xpb_out[89][626],u_xpb_out[90][626],u_xpb_out[91][626],u_xpb_out[92][626],u_xpb_out[93][626],u_xpb_out[94][626],u_xpb_out[95][626],u_xpb_out[96][626],u_xpb_out[97][626],u_xpb_out[98][626],u_xpb_out[99][626],u_xpb_out[100][626],u_xpb_out[101][626],u_xpb_out[102][626],u_xpb_out[103][626],u_xpb_out[104][626],u_xpb_out[105][626]};

assign col_out_627 = {u_xpb_out[0][627],u_xpb_out[1][627],u_xpb_out[2][627],u_xpb_out[3][627],u_xpb_out[4][627],u_xpb_out[5][627],u_xpb_out[6][627],u_xpb_out[7][627],u_xpb_out[8][627],u_xpb_out[9][627],u_xpb_out[10][627],u_xpb_out[11][627],u_xpb_out[12][627],u_xpb_out[13][627],u_xpb_out[14][627],u_xpb_out[15][627],u_xpb_out[16][627],u_xpb_out[17][627],u_xpb_out[18][627],u_xpb_out[19][627],u_xpb_out[20][627],u_xpb_out[21][627],u_xpb_out[22][627],u_xpb_out[23][627],u_xpb_out[24][627],u_xpb_out[25][627],u_xpb_out[26][627],u_xpb_out[27][627],u_xpb_out[28][627],u_xpb_out[29][627],u_xpb_out[30][627],u_xpb_out[31][627],u_xpb_out[32][627],u_xpb_out[33][627],u_xpb_out[34][627],u_xpb_out[35][627],u_xpb_out[36][627],u_xpb_out[37][627],u_xpb_out[38][627],u_xpb_out[39][627],u_xpb_out[40][627],u_xpb_out[41][627],u_xpb_out[42][627],u_xpb_out[43][627],u_xpb_out[44][627],u_xpb_out[45][627],u_xpb_out[46][627],u_xpb_out[47][627],u_xpb_out[48][627],u_xpb_out[49][627],u_xpb_out[50][627],u_xpb_out[51][627],u_xpb_out[52][627],u_xpb_out[53][627],u_xpb_out[54][627],u_xpb_out[55][627],u_xpb_out[56][627],u_xpb_out[57][627],u_xpb_out[58][627],u_xpb_out[59][627],u_xpb_out[60][627],u_xpb_out[61][627],u_xpb_out[62][627],u_xpb_out[63][627],u_xpb_out[64][627],u_xpb_out[65][627],u_xpb_out[66][627],u_xpb_out[67][627],u_xpb_out[68][627],u_xpb_out[69][627],u_xpb_out[70][627],u_xpb_out[71][627],u_xpb_out[72][627],u_xpb_out[73][627],u_xpb_out[74][627],u_xpb_out[75][627],u_xpb_out[76][627],u_xpb_out[77][627],u_xpb_out[78][627],u_xpb_out[79][627],u_xpb_out[80][627],u_xpb_out[81][627],u_xpb_out[82][627],u_xpb_out[83][627],u_xpb_out[84][627],u_xpb_out[85][627],u_xpb_out[86][627],u_xpb_out[87][627],u_xpb_out[88][627],u_xpb_out[89][627],u_xpb_out[90][627],u_xpb_out[91][627],u_xpb_out[92][627],u_xpb_out[93][627],u_xpb_out[94][627],u_xpb_out[95][627],u_xpb_out[96][627],u_xpb_out[97][627],u_xpb_out[98][627],u_xpb_out[99][627],u_xpb_out[100][627],u_xpb_out[101][627],u_xpb_out[102][627],u_xpb_out[103][627],u_xpb_out[104][627],u_xpb_out[105][627]};

assign col_out_628 = {u_xpb_out[0][628],u_xpb_out[1][628],u_xpb_out[2][628],u_xpb_out[3][628],u_xpb_out[4][628],u_xpb_out[5][628],u_xpb_out[6][628],u_xpb_out[7][628],u_xpb_out[8][628],u_xpb_out[9][628],u_xpb_out[10][628],u_xpb_out[11][628],u_xpb_out[12][628],u_xpb_out[13][628],u_xpb_out[14][628],u_xpb_out[15][628],u_xpb_out[16][628],u_xpb_out[17][628],u_xpb_out[18][628],u_xpb_out[19][628],u_xpb_out[20][628],u_xpb_out[21][628],u_xpb_out[22][628],u_xpb_out[23][628],u_xpb_out[24][628],u_xpb_out[25][628],u_xpb_out[26][628],u_xpb_out[27][628],u_xpb_out[28][628],u_xpb_out[29][628],u_xpb_out[30][628],u_xpb_out[31][628],u_xpb_out[32][628],u_xpb_out[33][628],u_xpb_out[34][628],u_xpb_out[35][628],u_xpb_out[36][628],u_xpb_out[37][628],u_xpb_out[38][628],u_xpb_out[39][628],u_xpb_out[40][628],u_xpb_out[41][628],u_xpb_out[42][628],u_xpb_out[43][628],u_xpb_out[44][628],u_xpb_out[45][628],u_xpb_out[46][628],u_xpb_out[47][628],u_xpb_out[48][628],u_xpb_out[49][628],u_xpb_out[50][628],u_xpb_out[51][628],u_xpb_out[52][628],u_xpb_out[53][628],u_xpb_out[54][628],u_xpb_out[55][628],u_xpb_out[56][628],u_xpb_out[57][628],u_xpb_out[58][628],u_xpb_out[59][628],u_xpb_out[60][628],u_xpb_out[61][628],u_xpb_out[62][628],u_xpb_out[63][628],u_xpb_out[64][628],u_xpb_out[65][628],u_xpb_out[66][628],u_xpb_out[67][628],u_xpb_out[68][628],u_xpb_out[69][628],u_xpb_out[70][628],u_xpb_out[71][628],u_xpb_out[72][628],u_xpb_out[73][628],u_xpb_out[74][628],u_xpb_out[75][628],u_xpb_out[76][628],u_xpb_out[77][628],u_xpb_out[78][628],u_xpb_out[79][628],u_xpb_out[80][628],u_xpb_out[81][628],u_xpb_out[82][628],u_xpb_out[83][628],u_xpb_out[84][628],u_xpb_out[85][628],u_xpb_out[86][628],u_xpb_out[87][628],u_xpb_out[88][628],u_xpb_out[89][628],u_xpb_out[90][628],u_xpb_out[91][628],u_xpb_out[92][628],u_xpb_out[93][628],u_xpb_out[94][628],u_xpb_out[95][628],u_xpb_out[96][628],u_xpb_out[97][628],u_xpb_out[98][628],u_xpb_out[99][628],u_xpb_out[100][628],u_xpb_out[101][628],u_xpb_out[102][628],u_xpb_out[103][628],u_xpb_out[104][628],u_xpb_out[105][628]};

assign col_out_629 = {u_xpb_out[0][629],u_xpb_out[1][629],u_xpb_out[2][629],u_xpb_out[3][629],u_xpb_out[4][629],u_xpb_out[5][629],u_xpb_out[6][629],u_xpb_out[7][629],u_xpb_out[8][629],u_xpb_out[9][629],u_xpb_out[10][629],u_xpb_out[11][629],u_xpb_out[12][629],u_xpb_out[13][629],u_xpb_out[14][629],u_xpb_out[15][629],u_xpb_out[16][629],u_xpb_out[17][629],u_xpb_out[18][629],u_xpb_out[19][629],u_xpb_out[20][629],u_xpb_out[21][629],u_xpb_out[22][629],u_xpb_out[23][629],u_xpb_out[24][629],u_xpb_out[25][629],u_xpb_out[26][629],u_xpb_out[27][629],u_xpb_out[28][629],u_xpb_out[29][629],u_xpb_out[30][629],u_xpb_out[31][629],u_xpb_out[32][629],u_xpb_out[33][629],u_xpb_out[34][629],u_xpb_out[35][629],u_xpb_out[36][629],u_xpb_out[37][629],u_xpb_out[38][629],u_xpb_out[39][629],u_xpb_out[40][629],u_xpb_out[41][629],u_xpb_out[42][629],u_xpb_out[43][629],u_xpb_out[44][629],u_xpb_out[45][629],u_xpb_out[46][629],u_xpb_out[47][629],u_xpb_out[48][629],u_xpb_out[49][629],u_xpb_out[50][629],u_xpb_out[51][629],u_xpb_out[52][629],u_xpb_out[53][629],u_xpb_out[54][629],u_xpb_out[55][629],u_xpb_out[56][629],u_xpb_out[57][629],u_xpb_out[58][629],u_xpb_out[59][629],u_xpb_out[60][629],u_xpb_out[61][629],u_xpb_out[62][629],u_xpb_out[63][629],u_xpb_out[64][629],u_xpb_out[65][629],u_xpb_out[66][629],u_xpb_out[67][629],u_xpb_out[68][629],u_xpb_out[69][629],u_xpb_out[70][629],u_xpb_out[71][629],u_xpb_out[72][629],u_xpb_out[73][629],u_xpb_out[74][629],u_xpb_out[75][629],u_xpb_out[76][629],u_xpb_out[77][629],u_xpb_out[78][629],u_xpb_out[79][629],u_xpb_out[80][629],u_xpb_out[81][629],u_xpb_out[82][629],u_xpb_out[83][629],u_xpb_out[84][629],u_xpb_out[85][629],u_xpb_out[86][629],u_xpb_out[87][629],u_xpb_out[88][629],u_xpb_out[89][629],u_xpb_out[90][629],u_xpb_out[91][629],u_xpb_out[92][629],u_xpb_out[93][629],u_xpb_out[94][629],u_xpb_out[95][629],u_xpb_out[96][629],u_xpb_out[97][629],u_xpb_out[98][629],u_xpb_out[99][629],u_xpb_out[100][629],u_xpb_out[101][629],u_xpb_out[102][629],u_xpb_out[103][629],u_xpb_out[104][629],u_xpb_out[105][629]};

assign col_out_630 = {u_xpb_out[0][630],u_xpb_out[1][630],u_xpb_out[2][630],u_xpb_out[3][630],u_xpb_out[4][630],u_xpb_out[5][630],u_xpb_out[6][630],u_xpb_out[7][630],u_xpb_out[8][630],u_xpb_out[9][630],u_xpb_out[10][630],u_xpb_out[11][630],u_xpb_out[12][630],u_xpb_out[13][630],u_xpb_out[14][630],u_xpb_out[15][630],u_xpb_out[16][630],u_xpb_out[17][630],u_xpb_out[18][630],u_xpb_out[19][630],u_xpb_out[20][630],u_xpb_out[21][630],u_xpb_out[22][630],u_xpb_out[23][630],u_xpb_out[24][630],u_xpb_out[25][630],u_xpb_out[26][630],u_xpb_out[27][630],u_xpb_out[28][630],u_xpb_out[29][630],u_xpb_out[30][630],u_xpb_out[31][630],u_xpb_out[32][630],u_xpb_out[33][630],u_xpb_out[34][630],u_xpb_out[35][630],u_xpb_out[36][630],u_xpb_out[37][630],u_xpb_out[38][630],u_xpb_out[39][630],u_xpb_out[40][630],u_xpb_out[41][630],u_xpb_out[42][630],u_xpb_out[43][630],u_xpb_out[44][630],u_xpb_out[45][630],u_xpb_out[46][630],u_xpb_out[47][630],u_xpb_out[48][630],u_xpb_out[49][630],u_xpb_out[50][630],u_xpb_out[51][630],u_xpb_out[52][630],u_xpb_out[53][630],u_xpb_out[54][630],u_xpb_out[55][630],u_xpb_out[56][630],u_xpb_out[57][630],u_xpb_out[58][630],u_xpb_out[59][630],u_xpb_out[60][630],u_xpb_out[61][630],u_xpb_out[62][630],u_xpb_out[63][630],u_xpb_out[64][630],u_xpb_out[65][630],u_xpb_out[66][630],u_xpb_out[67][630],u_xpb_out[68][630],u_xpb_out[69][630],u_xpb_out[70][630],u_xpb_out[71][630],u_xpb_out[72][630],u_xpb_out[73][630],u_xpb_out[74][630],u_xpb_out[75][630],u_xpb_out[76][630],u_xpb_out[77][630],u_xpb_out[78][630],u_xpb_out[79][630],u_xpb_out[80][630],u_xpb_out[81][630],u_xpb_out[82][630],u_xpb_out[83][630],u_xpb_out[84][630],u_xpb_out[85][630],u_xpb_out[86][630],u_xpb_out[87][630],u_xpb_out[88][630],u_xpb_out[89][630],u_xpb_out[90][630],u_xpb_out[91][630],u_xpb_out[92][630],u_xpb_out[93][630],u_xpb_out[94][630],u_xpb_out[95][630],u_xpb_out[96][630],u_xpb_out[97][630],u_xpb_out[98][630],u_xpb_out[99][630],u_xpb_out[100][630],u_xpb_out[101][630],u_xpb_out[102][630],u_xpb_out[103][630],u_xpb_out[104][630],u_xpb_out[105][630]};

assign col_out_631 = {u_xpb_out[0][631],u_xpb_out[1][631],u_xpb_out[2][631],u_xpb_out[3][631],u_xpb_out[4][631],u_xpb_out[5][631],u_xpb_out[6][631],u_xpb_out[7][631],u_xpb_out[8][631],u_xpb_out[9][631],u_xpb_out[10][631],u_xpb_out[11][631],u_xpb_out[12][631],u_xpb_out[13][631],u_xpb_out[14][631],u_xpb_out[15][631],u_xpb_out[16][631],u_xpb_out[17][631],u_xpb_out[18][631],u_xpb_out[19][631],u_xpb_out[20][631],u_xpb_out[21][631],u_xpb_out[22][631],u_xpb_out[23][631],u_xpb_out[24][631],u_xpb_out[25][631],u_xpb_out[26][631],u_xpb_out[27][631],u_xpb_out[28][631],u_xpb_out[29][631],u_xpb_out[30][631],u_xpb_out[31][631],u_xpb_out[32][631],u_xpb_out[33][631],u_xpb_out[34][631],u_xpb_out[35][631],u_xpb_out[36][631],u_xpb_out[37][631],u_xpb_out[38][631],u_xpb_out[39][631],u_xpb_out[40][631],u_xpb_out[41][631],u_xpb_out[42][631],u_xpb_out[43][631],u_xpb_out[44][631],u_xpb_out[45][631],u_xpb_out[46][631],u_xpb_out[47][631],u_xpb_out[48][631],u_xpb_out[49][631],u_xpb_out[50][631],u_xpb_out[51][631],u_xpb_out[52][631],u_xpb_out[53][631],u_xpb_out[54][631],u_xpb_out[55][631],u_xpb_out[56][631],u_xpb_out[57][631],u_xpb_out[58][631],u_xpb_out[59][631],u_xpb_out[60][631],u_xpb_out[61][631],u_xpb_out[62][631],u_xpb_out[63][631],u_xpb_out[64][631],u_xpb_out[65][631],u_xpb_out[66][631],u_xpb_out[67][631],u_xpb_out[68][631],u_xpb_out[69][631],u_xpb_out[70][631],u_xpb_out[71][631],u_xpb_out[72][631],u_xpb_out[73][631],u_xpb_out[74][631],u_xpb_out[75][631],u_xpb_out[76][631],u_xpb_out[77][631],u_xpb_out[78][631],u_xpb_out[79][631],u_xpb_out[80][631],u_xpb_out[81][631],u_xpb_out[82][631],u_xpb_out[83][631],u_xpb_out[84][631],u_xpb_out[85][631],u_xpb_out[86][631],u_xpb_out[87][631],u_xpb_out[88][631],u_xpb_out[89][631],u_xpb_out[90][631],u_xpb_out[91][631],u_xpb_out[92][631],u_xpb_out[93][631],u_xpb_out[94][631],u_xpb_out[95][631],u_xpb_out[96][631],u_xpb_out[97][631],u_xpb_out[98][631],u_xpb_out[99][631],u_xpb_out[100][631],u_xpb_out[101][631],u_xpb_out[102][631],u_xpb_out[103][631],u_xpb_out[104][631],u_xpb_out[105][631]};

assign col_out_632 = {u_xpb_out[0][632],u_xpb_out[1][632],u_xpb_out[2][632],u_xpb_out[3][632],u_xpb_out[4][632],u_xpb_out[5][632],u_xpb_out[6][632],u_xpb_out[7][632],u_xpb_out[8][632],u_xpb_out[9][632],u_xpb_out[10][632],u_xpb_out[11][632],u_xpb_out[12][632],u_xpb_out[13][632],u_xpb_out[14][632],u_xpb_out[15][632],u_xpb_out[16][632],u_xpb_out[17][632],u_xpb_out[18][632],u_xpb_out[19][632],u_xpb_out[20][632],u_xpb_out[21][632],u_xpb_out[22][632],u_xpb_out[23][632],u_xpb_out[24][632],u_xpb_out[25][632],u_xpb_out[26][632],u_xpb_out[27][632],u_xpb_out[28][632],u_xpb_out[29][632],u_xpb_out[30][632],u_xpb_out[31][632],u_xpb_out[32][632],u_xpb_out[33][632],u_xpb_out[34][632],u_xpb_out[35][632],u_xpb_out[36][632],u_xpb_out[37][632],u_xpb_out[38][632],u_xpb_out[39][632],u_xpb_out[40][632],u_xpb_out[41][632],u_xpb_out[42][632],u_xpb_out[43][632],u_xpb_out[44][632],u_xpb_out[45][632],u_xpb_out[46][632],u_xpb_out[47][632],u_xpb_out[48][632],u_xpb_out[49][632],u_xpb_out[50][632],u_xpb_out[51][632],u_xpb_out[52][632],u_xpb_out[53][632],u_xpb_out[54][632],u_xpb_out[55][632],u_xpb_out[56][632],u_xpb_out[57][632],u_xpb_out[58][632],u_xpb_out[59][632],u_xpb_out[60][632],u_xpb_out[61][632],u_xpb_out[62][632],u_xpb_out[63][632],u_xpb_out[64][632],u_xpb_out[65][632],u_xpb_out[66][632],u_xpb_out[67][632],u_xpb_out[68][632],u_xpb_out[69][632],u_xpb_out[70][632],u_xpb_out[71][632],u_xpb_out[72][632],u_xpb_out[73][632],u_xpb_out[74][632],u_xpb_out[75][632],u_xpb_out[76][632],u_xpb_out[77][632],u_xpb_out[78][632],u_xpb_out[79][632],u_xpb_out[80][632],u_xpb_out[81][632],u_xpb_out[82][632],u_xpb_out[83][632],u_xpb_out[84][632],u_xpb_out[85][632],u_xpb_out[86][632],u_xpb_out[87][632],u_xpb_out[88][632],u_xpb_out[89][632],u_xpb_out[90][632],u_xpb_out[91][632],u_xpb_out[92][632],u_xpb_out[93][632],u_xpb_out[94][632],u_xpb_out[95][632],u_xpb_out[96][632],u_xpb_out[97][632],u_xpb_out[98][632],u_xpb_out[99][632],u_xpb_out[100][632],u_xpb_out[101][632],u_xpb_out[102][632],u_xpb_out[103][632],u_xpb_out[104][632],u_xpb_out[105][632]};

assign col_out_633 = {u_xpb_out[0][633],u_xpb_out[1][633],u_xpb_out[2][633],u_xpb_out[3][633],u_xpb_out[4][633],u_xpb_out[5][633],u_xpb_out[6][633],u_xpb_out[7][633],u_xpb_out[8][633],u_xpb_out[9][633],u_xpb_out[10][633],u_xpb_out[11][633],u_xpb_out[12][633],u_xpb_out[13][633],u_xpb_out[14][633],u_xpb_out[15][633],u_xpb_out[16][633],u_xpb_out[17][633],u_xpb_out[18][633],u_xpb_out[19][633],u_xpb_out[20][633],u_xpb_out[21][633],u_xpb_out[22][633],u_xpb_out[23][633],u_xpb_out[24][633],u_xpb_out[25][633],u_xpb_out[26][633],u_xpb_out[27][633],u_xpb_out[28][633],u_xpb_out[29][633],u_xpb_out[30][633],u_xpb_out[31][633],u_xpb_out[32][633],u_xpb_out[33][633],u_xpb_out[34][633],u_xpb_out[35][633],u_xpb_out[36][633],u_xpb_out[37][633],u_xpb_out[38][633],u_xpb_out[39][633],u_xpb_out[40][633],u_xpb_out[41][633],u_xpb_out[42][633],u_xpb_out[43][633],u_xpb_out[44][633],u_xpb_out[45][633],u_xpb_out[46][633],u_xpb_out[47][633],u_xpb_out[48][633],u_xpb_out[49][633],u_xpb_out[50][633],u_xpb_out[51][633],u_xpb_out[52][633],u_xpb_out[53][633],u_xpb_out[54][633],u_xpb_out[55][633],u_xpb_out[56][633],u_xpb_out[57][633],u_xpb_out[58][633],u_xpb_out[59][633],u_xpb_out[60][633],u_xpb_out[61][633],u_xpb_out[62][633],u_xpb_out[63][633],u_xpb_out[64][633],u_xpb_out[65][633],u_xpb_out[66][633],u_xpb_out[67][633],u_xpb_out[68][633],u_xpb_out[69][633],u_xpb_out[70][633],u_xpb_out[71][633],u_xpb_out[72][633],u_xpb_out[73][633],u_xpb_out[74][633],u_xpb_out[75][633],u_xpb_out[76][633],u_xpb_out[77][633],u_xpb_out[78][633],u_xpb_out[79][633],u_xpb_out[80][633],u_xpb_out[81][633],u_xpb_out[82][633],u_xpb_out[83][633],u_xpb_out[84][633],u_xpb_out[85][633],u_xpb_out[86][633],u_xpb_out[87][633],u_xpb_out[88][633],u_xpb_out[89][633],u_xpb_out[90][633],u_xpb_out[91][633],u_xpb_out[92][633],u_xpb_out[93][633],u_xpb_out[94][633],u_xpb_out[95][633],u_xpb_out[96][633],u_xpb_out[97][633],u_xpb_out[98][633],u_xpb_out[99][633],u_xpb_out[100][633],u_xpb_out[101][633],u_xpb_out[102][633],u_xpb_out[103][633],u_xpb_out[104][633],u_xpb_out[105][633]};

assign col_out_634 = {u_xpb_out[0][634],u_xpb_out[1][634],u_xpb_out[2][634],u_xpb_out[3][634],u_xpb_out[4][634],u_xpb_out[5][634],u_xpb_out[6][634],u_xpb_out[7][634],u_xpb_out[8][634],u_xpb_out[9][634],u_xpb_out[10][634],u_xpb_out[11][634],u_xpb_out[12][634],u_xpb_out[13][634],u_xpb_out[14][634],u_xpb_out[15][634],u_xpb_out[16][634],u_xpb_out[17][634],u_xpb_out[18][634],u_xpb_out[19][634],u_xpb_out[20][634],u_xpb_out[21][634],u_xpb_out[22][634],u_xpb_out[23][634],u_xpb_out[24][634],u_xpb_out[25][634],u_xpb_out[26][634],u_xpb_out[27][634],u_xpb_out[28][634],u_xpb_out[29][634],u_xpb_out[30][634],u_xpb_out[31][634],u_xpb_out[32][634],u_xpb_out[33][634],u_xpb_out[34][634],u_xpb_out[35][634],u_xpb_out[36][634],u_xpb_out[37][634],u_xpb_out[38][634],u_xpb_out[39][634],u_xpb_out[40][634],u_xpb_out[41][634],u_xpb_out[42][634],u_xpb_out[43][634],u_xpb_out[44][634],u_xpb_out[45][634],u_xpb_out[46][634],u_xpb_out[47][634],u_xpb_out[48][634],u_xpb_out[49][634],u_xpb_out[50][634],u_xpb_out[51][634],u_xpb_out[52][634],u_xpb_out[53][634],u_xpb_out[54][634],u_xpb_out[55][634],u_xpb_out[56][634],u_xpb_out[57][634],u_xpb_out[58][634],u_xpb_out[59][634],u_xpb_out[60][634],u_xpb_out[61][634],u_xpb_out[62][634],u_xpb_out[63][634],u_xpb_out[64][634],u_xpb_out[65][634],u_xpb_out[66][634],u_xpb_out[67][634],u_xpb_out[68][634],u_xpb_out[69][634],u_xpb_out[70][634],u_xpb_out[71][634],u_xpb_out[72][634],u_xpb_out[73][634],u_xpb_out[74][634],u_xpb_out[75][634],u_xpb_out[76][634],u_xpb_out[77][634],u_xpb_out[78][634],u_xpb_out[79][634],u_xpb_out[80][634],u_xpb_out[81][634],u_xpb_out[82][634],u_xpb_out[83][634],u_xpb_out[84][634],u_xpb_out[85][634],u_xpb_out[86][634],u_xpb_out[87][634],u_xpb_out[88][634],u_xpb_out[89][634],u_xpb_out[90][634],u_xpb_out[91][634],u_xpb_out[92][634],u_xpb_out[93][634],u_xpb_out[94][634],u_xpb_out[95][634],u_xpb_out[96][634],u_xpb_out[97][634],u_xpb_out[98][634],u_xpb_out[99][634],u_xpb_out[100][634],u_xpb_out[101][634],u_xpb_out[102][634],u_xpb_out[103][634],u_xpb_out[104][634],u_xpb_out[105][634]};

assign col_out_635 = {u_xpb_out[0][635],u_xpb_out[1][635],u_xpb_out[2][635],u_xpb_out[3][635],u_xpb_out[4][635],u_xpb_out[5][635],u_xpb_out[6][635],u_xpb_out[7][635],u_xpb_out[8][635],u_xpb_out[9][635],u_xpb_out[10][635],u_xpb_out[11][635],u_xpb_out[12][635],u_xpb_out[13][635],u_xpb_out[14][635],u_xpb_out[15][635],u_xpb_out[16][635],u_xpb_out[17][635],u_xpb_out[18][635],u_xpb_out[19][635],u_xpb_out[20][635],u_xpb_out[21][635],u_xpb_out[22][635],u_xpb_out[23][635],u_xpb_out[24][635],u_xpb_out[25][635],u_xpb_out[26][635],u_xpb_out[27][635],u_xpb_out[28][635],u_xpb_out[29][635],u_xpb_out[30][635],u_xpb_out[31][635],u_xpb_out[32][635],u_xpb_out[33][635],u_xpb_out[34][635],u_xpb_out[35][635],u_xpb_out[36][635],u_xpb_out[37][635],u_xpb_out[38][635],u_xpb_out[39][635],u_xpb_out[40][635],u_xpb_out[41][635],u_xpb_out[42][635],u_xpb_out[43][635],u_xpb_out[44][635],u_xpb_out[45][635],u_xpb_out[46][635],u_xpb_out[47][635],u_xpb_out[48][635],u_xpb_out[49][635],u_xpb_out[50][635],u_xpb_out[51][635],u_xpb_out[52][635],u_xpb_out[53][635],u_xpb_out[54][635],u_xpb_out[55][635],u_xpb_out[56][635],u_xpb_out[57][635],u_xpb_out[58][635],u_xpb_out[59][635],u_xpb_out[60][635],u_xpb_out[61][635],u_xpb_out[62][635],u_xpb_out[63][635],u_xpb_out[64][635],u_xpb_out[65][635],u_xpb_out[66][635],u_xpb_out[67][635],u_xpb_out[68][635],u_xpb_out[69][635],u_xpb_out[70][635],u_xpb_out[71][635],u_xpb_out[72][635],u_xpb_out[73][635],u_xpb_out[74][635],u_xpb_out[75][635],u_xpb_out[76][635],u_xpb_out[77][635],u_xpb_out[78][635],u_xpb_out[79][635],u_xpb_out[80][635],u_xpb_out[81][635],u_xpb_out[82][635],u_xpb_out[83][635],u_xpb_out[84][635],u_xpb_out[85][635],u_xpb_out[86][635],u_xpb_out[87][635],u_xpb_out[88][635],u_xpb_out[89][635],u_xpb_out[90][635],u_xpb_out[91][635],u_xpb_out[92][635],u_xpb_out[93][635],u_xpb_out[94][635],u_xpb_out[95][635],u_xpb_out[96][635],u_xpb_out[97][635],u_xpb_out[98][635],u_xpb_out[99][635],u_xpb_out[100][635],u_xpb_out[101][635],u_xpb_out[102][635],u_xpb_out[103][635],u_xpb_out[104][635],u_xpb_out[105][635]};

assign col_out_636 = {u_xpb_out[0][636],u_xpb_out[1][636],u_xpb_out[2][636],u_xpb_out[3][636],u_xpb_out[4][636],u_xpb_out[5][636],u_xpb_out[6][636],u_xpb_out[7][636],u_xpb_out[8][636],u_xpb_out[9][636],u_xpb_out[10][636],u_xpb_out[11][636],u_xpb_out[12][636],u_xpb_out[13][636],u_xpb_out[14][636],u_xpb_out[15][636],u_xpb_out[16][636],u_xpb_out[17][636],u_xpb_out[18][636],u_xpb_out[19][636],u_xpb_out[20][636],u_xpb_out[21][636],u_xpb_out[22][636],u_xpb_out[23][636],u_xpb_out[24][636],u_xpb_out[25][636],u_xpb_out[26][636],u_xpb_out[27][636],u_xpb_out[28][636],u_xpb_out[29][636],u_xpb_out[30][636],u_xpb_out[31][636],u_xpb_out[32][636],u_xpb_out[33][636],u_xpb_out[34][636],u_xpb_out[35][636],u_xpb_out[36][636],u_xpb_out[37][636],u_xpb_out[38][636],u_xpb_out[39][636],u_xpb_out[40][636],u_xpb_out[41][636],u_xpb_out[42][636],u_xpb_out[43][636],u_xpb_out[44][636],u_xpb_out[45][636],u_xpb_out[46][636],u_xpb_out[47][636],u_xpb_out[48][636],u_xpb_out[49][636],u_xpb_out[50][636],u_xpb_out[51][636],u_xpb_out[52][636],u_xpb_out[53][636],u_xpb_out[54][636],u_xpb_out[55][636],u_xpb_out[56][636],u_xpb_out[57][636],u_xpb_out[58][636],u_xpb_out[59][636],u_xpb_out[60][636],u_xpb_out[61][636],u_xpb_out[62][636],u_xpb_out[63][636],u_xpb_out[64][636],u_xpb_out[65][636],u_xpb_out[66][636],u_xpb_out[67][636],u_xpb_out[68][636],u_xpb_out[69][636],u_xpb_out[70][636],u_xpb_out[71][636],u_xpb_out[72][636],u_xpb_out[73][636],u_xpb_out[74][636],u_xpb_out[75][636],u_xpb_out[76][636],u_xpb_out[77][636],u_xpb_out[78][636],u_xpb_out[79][636],u_xpb_out[80][636],u_xpb_out[81][636],u_xpb_out[82][636],u_xpb_out[83][636],u_xpb_out[84][636],u_xpb_out[85][636],u_xpb_out[86][636],u_xpb_out[87][636],u_xpb_out[88][636],u_xpb_out[89][636],u_xpb_out[90][636],u_xpb_out[91][636],u_xpb_out[92][636],u_xpb_out[93][636],u_xpb_out[94][636],u_xpb_out[95][636],u_xpb_out[96][636],u_xpb_out[97][636],u_xpb_out[98][636],u_xpb_out[99][636],u_xpb_out[100][636],u_xpb_out[101][636],u_xpb_out[102][636],u_xpb_out[103][636],u_xpb_out[104][636],u_xpb_out[105][636]};

assign col_out_637 = {u_xpb_out[0][637],u_xpb_out[1][637],u_xpb_out[2][637],u_xpb_out[3][637],u_xpb_out[4][637],u_xpb_out[5][637],u_xpb_out[6][637],u_xpb_out[7][637],u_xpb_out[8][637],u_xpb_out[9][637],u_xpb_out[10][637],u_xpb_out[11][637],u_xpb_out[12][637],u_xpb_out[13][637],u_xpb_out[14][637],u_xpb_out[15][637],u_xpb_out[16][637],u_xpb_out[17][637],u_xpb_out[18][637],u_xpb_out[19][637],u_xpb_out[20][637],u_xpb_out[21][637],u_xpb_out[22][637],u_xpb_out[23][637],u_xpb_out[24][637],u_xpb_out[25][637],u_xpb_out[26][637],u_xpb_out[27][637],u_xpb_out[28][637],u_xpb_out[29][637],u_xpb_out[30][637],u_xpb_out[31][637],u_xpb_out[32][637],u_xpb_out[33][637],u_xpb_out[34][637],u_xpb_out[35][637],u_xpb_out[36][637],u_xpb_out[37][637],u_xpb_out[38][637],u_xpb_out[39][637],u_xpb_out[40][637],u_xpb_out[41][637],u_xpb_out[42][637],u_xpb_out[43][637],u_xpb_out[44][637],u_xpb_out[45][637],u_xpb_out[46][637],u_xpb_out[47][637],u_xpb_out[48][637],u_xpb_out[49][637],u_xpb_out[50][637],u_xpb_out[51][637],u_xpb_out[52][637],u_xpb_out[53][637],u_xpb_out[54][637],u_xpb_out[55][637],u_xpb_out[56][637],u_xpb_out[57][637],u_xpb_out[58][637],u_xpb_out[59][637],u_xpb_out[60][637],u_xpb_out[61][637],u_xpb_out[62][637],u_xpb_out[63][637],u_xpb_out[64][637],u_xpb_out[65][637],u_xpb_out[66][637],u_xpb_out[67][637],u_xpb_out[68][637],u_xpb_out[69][637],u_xpb_out[70][637],u_xpb_out[71][637],u_xpb_out[72][637],u_xpb_out[73][637],u_xpb_out[74][637],u_xpb_out[75][637],u_xpb_out[76][637],u_xpb_out[77][637],u_xpb_out[78][637],u_xpb_out[79][637],u_xpb_out[80][637],u_xpb_out[81][637],u_xpb_out[82][637],u_xpb_out[83][637],u_xpb_out[84][637],u_xpb_out[85][637],u_xpb_out[86][637],u_xpb_out[87][637],u_xpb_out[88][637],u_xpb_out[89][637],u_xpb_out[90][637],u_xpb_out[91][637],u_xpb_out[92][637],u_xpb_out[93][637],u_xpb_out[94][637],u_xpb_out[95][637],u_xpb_out[96][637],u_xpb_out[97][637],u_xpb_out[98][637],u_xpb_out[99][637],u_xpb_out[100][637],u_xpb_out[101][637],u_xpb_out[102][637],u_xpb_out[103][637],u_xpb_out[104][637],u_xpb_out[105][637]};

assign col_out_638 = {u_xpb_out[0][638],u_xpb_out[1][638],u_xpb_out[2][638],u_xpb_out[3][638],u_xpb_out[4][638],u_xpb_out[5][638],u_xpb_out[6][638],u_xpb_out[7][638],u_xpb_out[8][638],u_xpb_out[9][638],u_xpb_out[10][638],u_xpb_out[11][638],u_xpb_out[12][638],u_xpb_out[13][638],u_xpb_out[14][638],u_xpb_out[15][638],u_xpb_out[16][638],u_xpb_out[17][638],u_xpb_out[18][638],u_xpb_out[19][638],u_xpb_out[20][638],u_xpb_out[21][638],u_xpb_out[22][638],u_xpb_out[23][638],u_xpb_out[24][638],u_xpb_out[25][638],u_xpb_out[26][638],u_xpb_out[27][638],u_xpb_out[28][638],u_xpb_out[29][638],u_xpb_out[30][638],u_xpb_out[31][638],u_xpb_out[32][638],u_xpb_out[33][638],u_xpb_out[34][638],u_xpb_out[35][638],u_xpb_out[36][638],u_xpb_out[37][638],u_xpb_out[38][638],u_xpb_out[39][638],u_xpb_out[40][638],u_xpb_out[41][638],u_xpb_out[42][638],u_xpb_out[43][638],u_xpb_out[44][638],u_xpb_out[45][638],u_xpb_out[46][638],u_xpb_out[47][638],u_xpb_out[48][638],u_xpb_out[49][638],u_xpb_out[50][638],u_xpb_out[51][638],u_xpb_out[52][638],u_xpb_out[53][638],u_xpb_out[54][638],u_xpb_out[55][638],u_xpb_out[56][638],u_xpb_out[57][638],u_xpb_out[58][638],u_xpb_out[59][638],u_xpb_out[60][638],u_xpb_out[61][638],u_xpb_out[62][638],u_xpb_out[63][638],u_xpb_out[64][638],u_xpb_out[65][638],u_xpb_out[66][638],u_xpb_out[67][638],u_xpb_out[68][638],u_xpb_out[69][638],u_xpb_out[70][638],u_xpb_out[71][638],u_xpb_out[72][638],u_xpb_out[73][638],u_xpb_out[74][638],u_xpb_out[75][638],u_xpb_out[76][638],u_xpb_out[77][638],u_xpb_out[78][638],u_xpb_out[79][638],u_xpb_out[80][638],u_xpb_out[81][638],u_xpb_out[82][638],u_xpb_out[83][638],u_xpb_out[84][638],u_xpb_out[85][638],u_xpb_out[86][638],u_xpb_out[87][638],u_xpb_out[88][638],u_xpb_out[89][638],u_xpb_out[90][638],u_xpb_out[91][638],u_xpb_out[92][638],u_xpb_out[93][638],u_xpb_out[94][638],u_xpb_out[95][638],u_xpb_out[96][638],u_xpb_out[97][638],u_xpb_out[98][638],u_xpb_out[99][638],u_xpb_out[100][638],u_xpb_out[101][638],u_xpb_out[102][638],u_xpb_out[103][638],u_xpb_out[104][638],u_xpb_out[105][638]};

assign col_out_639 = {u_xpb_out[0][639],u_xpb_out[1][639],u_xpb_out[2][639],u_xpb_out[3][639],u_xpb_out[4][639],u_xpb_out[5][639],u_xpb_out[6][639],u_xpb_out[7][639],u_xpb_out[8][639],u_xpb_out[9][639],u_xpb_out[10][639],u_xpb_out[11][639],u_xpb_out[12][639],u_xpb_out[13][639],u_xpb_out[14][639],u_xpb_out[15][639],u_xpb_out[16][639],u_xpb_out[17][639],u_xpb_out[18][639],u_xpb_out[19][639],u_xpb_out[20][639],u_xpb_out[21][639],u_xpb_out[22][639],u_xpb_out[23][639],u_xpb_out[24][639],u_xpb_out[25][639],u_xpb_out[26][639],u_xpb_out[27][639],u_xpb_out[28][639],u_xpb_out[29][639],u_xpb_out[30][639],u_xpb_out[31][639],u_xpb_out[32][639],u_xpb_out[33][639],u_xpb_out[34][639],u_xpb_out[35][639],u_xpb_out[36][639],u_xpb_out[37][639],u_xpb_out[38][639],u_xpb_out[39][639],u_xpb_out[40][639],u_xpb_out[41][639],u_xpb_out[42][639],u_xpb_out[43][639],u_xpb_out[44][639],u_xpb_out[45][639],u_xpb_out[46][639],u_xpb_out[47][639],u_xpb_out[48][639],u_xpb_out[49][639],u_xpb_out[50][639],u_xpb_out[51][639],u_xpb_out[52][639],u_xpb_out[53][639],u_xpb_out[54][639],u_xpb_out[55][639],u_xpb_out[56][639],u_xpb_out[57][639],u_xpb_out[58][639],u_xpb_out[59][639],u_xpb_out[60][639],u_xpb_out[61][639],u_xpb_out[62][639],u_xpb_out[63][639],u_xpb_out[64][639],u_xpb_out[65][639],u_xpb_out[66][639],u_xpb_out[67][639],u_xpb_out[68][639],u_xpb_out[69][639],u_xpb_out[70][639],u_xpb_out[71][639],u_xpb_out[72][639],u_xpb_out[73][639],u_xpb_out[74][639],u_xpb_out[75][639],u_xpb_out[76][639],u_xpb_out[77][639],u_xpb_out[78][639],u_xpb_out[79][639],u_xpb_out[80][639],u_xpb_out[81][639],u_xpb_out[82][639],u_xpb_out[83][639],u_xpb_out[84][639],u_xpb_out[85][639],u_xpb_out[86][639],u_xpb_out[87][639],u_xpb_out[88][639],u_xpb_out[89][639],u_xpb_out[90][639],u_xpb_out[91][639],u_xpb_out[92][639],u_xpb_out[93][639],u_xpb_out[94][639],u_xpb_out[95][639],u_xpb_out[96][639],u_xpb_out[97][639],u_xpb_out[98][639],u_xpb_out[99][639],u_xpb_out[100][639],u_xpb_out[101][639],u_xpb_out[102][639],u_xpb_out[103][639],u_xpb_out[104][639],u_xpb_out[105][639]};

assign col_out_640 = {u_xpb_out[0][640],u_xpb_out[1][640],u_xpb_out[2][640],u_xpb_out[3][640],u_xpb_out[4][640],u_xpb_out[5][640],u_xpb_out[6][640],u_xpb_out[7][640],u_xpb_out[8][640],u_xpb_out[9][640],u_xpb_out[10][640],u_xpb_out[11][640],u_xpb_out[12][640],u_xpb_out[13][640],u_xpb_out[14][640],u_xpb_out[15][640],u_xpb_out[16][640],u_xpb_out[17][640],u_xpb_out[18][640],u_xpb_out[19][640],u_xpb_out[20][640],u_xpb_out[21][640],u_xpb_out[22][640],u_xpb_out[23][640],u_xpb_out[24][640],u_xpb_out[25][640],u_xpb_out[26][640],u_xpb_out[27][640],u_xpb_out[28][640],u_xpb_out[29][640],u_xpb_out[30][640],u_xpb_out[31][640],u_xpb_out[32][640],u_xpb_out[33][640],u_xpb_out[34][640],u_xpb_out[35][640],u_xpb_out[36][640],u_xpb_out[37][640],u_xpb_out[38][640],u_xpb_out[39][640],u_xpb_out[40][640],u_xpb_out[41][640],u_xpb_out[42][640],u_xpb_out[43][640],u_xpb_out[44][640],u_xpb_out[45][640],u_xpb_out[46][640],u_xpb_out[47][640],u_xpb_out[48][640],u_xpb_out[49][640],u_xpb_out[50][640],u_xpb_out[51][640],u_xpb_out[52][640],u_xpb_out[53][640],u_xpb_out[54][640],u_xpb_out[55][640],u_xpb_out[56][640],u_xpb_out[57][640],u_xpb_out[58][640],u_xpb_out[59][640],u_xpb_out[60][640],u_xpb_out[61][640],u_xpb_out[62][640],u_xpb_out[63][640],u_xpb_out[64][640],u_xpb_out[65][640],u_xpb_out[66][640],u_xpb_out[67][640],u_xpb_out[68][640],u_xpb_out[69][640],u_xpb_out[70][640],u_xpb_out[71][640],u_xpb_out[72][640],u_xpb_out[73][640],u_xpb_out[74][640],u_xpb_out[75][640],u_xpb_out[76][640],u_xpb_out[77][640],u_xpb_out[78][640],u_xpb_out[79][640],u_xpb_out[80][640],u_xpb_out[81][640],u_xpb_out[82][640],u_xpb_out[83][640],u_xpb_out[84][640],u_xpb_out[85][640],u_xpb_out[86][640],u_xpb_out[87][640],u_xpb_out[88][640],u_xpb_out[89][640],u_xpb_out[90][640],u_xpb_out[91][640],u_xpb_out[92][640],u_xpb_out[93][640],u_xpb_out[94][640],u_xpb_out[95][640],u_xpb_out[96][640],u_xpb_out[97][640],u_xpb_out[98][640],u_xpb_out[99][640],u_xpb_out[100][640],u_xpb_out[101][640],u_xpb_out[102][640],u_xpb_out[103][640],u_xpb_out[104][640],u_xpb_out[105][640]};

assign col_out_641 = {u_xpb_out[0][641],u_xpb_out[1][641],u_xpb_out[2][641],u_xpb_out[3][641],u_xpb_out[4][641],u_xpb_out[5][641],u_xpb_out[6][641],u_xpb_out[7][641],u_xpb_out[8][641],u_xpb_out[9][641],u_xpb_out[10][641],u_xpb_out[11][641],u_xpb_out[12][641],u_xpb_out[13][641],u_xpb_out[14][641],u_xpb_out[15][641],u_xpb_out[16][641],u_xpb_out[17][641],u_xpb_out[18][641],u_xpb_out[19][641],u_xpb_out[20][641],u_xpb_out[21][641],u_xpb_out[22][641],u_xpb_out[23][641],u_xpb_out[24][641],u_xpb_out[25][641],u_xpb_out[26][641],u_xpb_out[27][641],u_xpb_out[28][641],u_xpb_out[29][641],u_xpb_out[30][641],u_xpb_out[31][641],u_xpb_out[32][641],u_xpb_out[33][641],u_xpb_out[34][641],u_xpb_out[35][641],u_xpb_out[36][641],u_xpb_out[37][641],u_xpb_out[38][641],u_xpb_out[39][641],u_xpb_out[40][641],u_xpb_out[41][641],u_xpb_out[42][641],u_xpb_out[43][641],u_xpb_out[44][641],u_xpb_out[45][641],u_xpb_out[46][641],u_xpb_out[47][641],u_xpb_out[48][641],u_xpb_out[49][641],u_xpb_out[50][641],u_xpb_out[51][641],u_xpb_out[52][641],u_xpb_out[53][641],u_xpb_out[54][641],u_xpb_out[55][641],u_xpb_out[56][641],u_xpb_out[57][641],u_xpb_out[58][641],u_xpb_out[59][641],u_xpb_out[60][641],u_xpb_out[61][641],u_xpb_out[62][641],u_xpb_out[63][641],u_xpb_out[64][641],u_xpb_out[65][641],u_xpb_out[66][641],u_xpb_out[67][641],u_xpb_out[68][641],u_xpb_out[69][641],u_xpb_out[70][641],u_xpb_out[71][641],u_xpb_out[72][641],u_xpb_out[73][641],u_xpb_out[74][641],u_xpb_out[75][641],u_xpb_out[76][641],u_xpb_out[77][641],u_xpb_out[78][641],u_xpb_out[79][641],u_xpb_out[80][641],u_xpb_out[81][641],u_xpb_out[82][641],u_xpb_out[83][641],u_xpb_out[84][641],u_xpb_out[85][641],u_xpb_out[86][641],u_xpb_out[87][641],u_xpb_out[88][641],u_xpb_out[89][641],u_xpb_out[90][641],u_xpb_out[91][641],u_xpb_out[92][641],u_xpb_out[93][641],u_xpb_out[94][641],u_xpb_out[95][641],u_xpb_out[96][641],u_xpb_out[97][641],u_xpb_out[98][641],u_xpb_out[99][641],u_xpb_out[100][641],u_xpb_out[101][641],u_xpb_out[102][641],u_xpb_out[103][641],u_xpb_out[104][641],u_xpb_out[105][641]};

assign col_out_642 = {u_xpb_out[0][642],u_xpb_out[1][642],u_xpb_out[2][642],u_xpb_out[3][642],u_xpb_out[4][642],u_xpb_out[5][642],u_xpb_out[6][642],u_xpb_out[7][642],u_xpb_out[8][642],u_xpb_out[9][642],u_xpb_out[10][642],u_xpb_out[11][642],u_xpb_out[12][642],u_xpb_out[13][642],u_xpb_out[14][642],u_xpb_out[15][642],u_xpb_out[16][642],u_xpb_out[17][642],u_xpb_out[18][642],u_xpb_out[19][642],u_xpb_out[20][642],u_xpb_out[21][642],u_xpb_out[22][642],u_xpb_out[23][642],u_xpb_out[24][642],u_xpb_out[25][642],u_xpb_out[26][642],u_xpb_out[27][642],u_xpb_out[28][642],u_xpb_out[29][642],u_xpb_out[30][642],u_xpb_out[31][642],u_xpb_out[32][642],u_xpb_out[33][642],u_xpb_out[34][642],u_xpb_out[35][642],u_xpb_out[36][642],u_xpb_out[37][642],u_xpb_out[38][642],u_xpb_out[39][642],u_xpb_out[40][642],u_xpb_out[41][642],u_xpb_out[42][642],u_xpb_out[43][642],u_xpb_out[44][642],u_xpb_out[45][642],u_xpb_out[46][642],u_xpb_out[47][642],u_xpb_out[48][642],u_xpb_out[49][642],u_xpb_out[50][642],u_xpb_out[51][642],u_xpb_out[52][642],u_xpb_out[53][642],u_xpb_out[54][642],u_xpb_out[55][642],u_xpb_out[56][642],u_xpb_out[57][642],u_xpb_out[58][642],u_xpb_out[59][642],u_xpb_out[60][642],u_xpb_out[61][642],u_xpb_out[62][642],u_xpb_out[63][642],u_xpb_out[64][642],u_xpb_out[65][642],u_xpb_out[66][642],u_xpb_out[67][642],u_xpb_out[68][642],u_xpb_out[69][642],u_xpb_out[70][642],u_xpb_out[71][642],u_xpb_out[72][642],u_xpb_out[73][642],u_xpb_out[74][642],u_xpb_out[75][642],u_xpb_out[76][642],u_xpb_out[77][642],u_xpb_out[78][642],u_xpb_out[79][642],u_xpb_out[80][642],u_xpb_out[81][642],u_xpb_out[82][642],u_xpb_out[83][642],u_xpb_out[84][642],u_xpb_out[85][642],u_xpb_out[86][642],u_xpb_out[87][642],u_xpb_out[88][642],u_xpb_out[89][642],u_xpb_out[90][642],u_xpb_out[91][642],u_xpb_out[92][642],u_xpb_out[93][642],u_xpb_out[94][642],u_xpb_out[95][642],u_xpb_out[96][642],u_xpb_out[97][642],u_xpb_out[98][642],u_xpb_out[99][642],u_xpb_out[100][642],u_xpb_out[101][642],u_xpb_out[102][642],u_xpb_out[103][642],u_xpb_out[104][642],u_xpb_out[105][642]};

assign col_out_643 = {u_xpb_out[0][643],u_xpb_out[1][643],u_xpb_out[2][643],u_xpb_out[3][643],u_xpb_out[4][643],u_xpb_out[5][643],u_xpb_out[6][643],u_xpb_out[7][643],u_xpb_out[8][643],u_xpb_out[9][643],u_xpb_out[10][643],u_xpb_out[11][643],u_xpb_out[12][643],u_xpb_out[13][643],u_xpb_out[14][643],u_xpb_out[15][643],u_xpb_out[16][643],u_xpb_out[17][643],u_xpb_out[18][643],u_xpb_out[19][643],u_xpb_out[20][643],u_xpb_out[21][643],u_xpb_out[22][643],u_xpb_out[23][643],u_xpb_out[24][643],u_xpb_out[25][643],u_xpb_out[26][643],u_xpb_out[27][643],u_xpb_out[28][643],u_xpb_out[29][643],u_xpb_out[30][643],u_xpb_out[31][643],u_xpb_out[32][643],u_xpb_out[33][643],u_xpb_out[34][643],u_xpb_out[35][643],u_xpb_out[36][643],u_xpb_out[37][643],u_xpb_out[38][643],u_xpb_out[39][643],u_xpb_out[40][643],u_xpb_out[41][643],u_xpb_out[42][643],u_xpb_out[43][643],u_xpb_out[44][643],u_xpb_out[45][643],u_xpb_out[46][643],u_xpb_out[47][643],u_xpb_out[48][643],u_xpb_out[49][643],u_xpb_out[50][643],u_xpb_out[51][643],u_xpb_out[52][643],u_xpb_out[53][643],u_xpb_out[54][643],u_xpb_out[55][643],u_xpb_out[56][643],u_xpb_out[57][643],u_xpb_out[58][643],u_xpb_out[59][643],u_xpb_out[60][643],u_xpb_out[61][643],u_xpb_out[62][643],u_xpb_out[63][643],u_xpb_out[64][643],u_xpb_out[65][643],u_xpb_out[66][643],u_xpb_out[67][643],u_xpb_out[68][643],u_xpb_out[69][643],u_xpb_out[70][643],u_xpb_out[71][643],u_xpb_out[72][643],u_xpb_out[73][643],u_xpb_out[74][643],u_xpb_out[75][643],u_xpb_out[76][643],u_xpb_out[77][643],u_xpb_out[78][643],u_xpb_out[79][643],u_xpb_out[80][643],u_xpb_out[81][643],u_xpb_out[82][643],u_xpb_out[83][643],u_xpb_out[84][643],u_xpb_out[85][643],u_xpb_out[86][643],u_xpb_out[87][643],u_xpb_out[88][643],u_xpb_out[89][643],u_xpb_out[90][643],u_xpb_out[91][643],u_xpb_out[92][643],u_xpb_out[93][643],u_xpb_out[94][643],u_xpb_out[95][643],u_xpb_out[96][643],u_xpb_out[97][643],u_xpb_out[98][643],u_xpb_out[99][643],u_xpb_out[100][643],u_xpb_out[101][643],u_xpb_out[102][643],u_xpb_out[103][643],u_xpb_out[104][643],u_xpb_out[105][643]};

assign col_out_644 = {u_xpb_out[0][644],u_xpb_out[1][644],u_xpb_out[2][644],u_xpb_out[3][644],u_xpb_out[4][644],u_xpb_out[5][644],u_xpb_out[6][644],u_xpb_out[7][644],u_xpb_out[8][644],u_xpb_out[9][644],u_xpb_out[10][644],u_xpb_out[11][644],u_xpb_out[12][644],u_xpb_out[13][644],u_xpb_out[14][644],u_xpb_out[15][644],u_xpb_out[16][644],u_xpb_out[17][644],u_xpb_out[18][644],u_xpb_out[19][644],u_xpb_out[20][644],u_xpb_out[21][644],u_xpb_out[22][644],u_xpb_out[23][644],u_xpb_out[24][644],u_xpb_out[25][644],u_xpb_out[26][644],u_xpb_out[27][644],u_xpb_out[28][644],u_xpb_out[29][644],u_xpb_out[30][644],u_xpb_out[31][644],u_xpb_out[32][644],u_xpb_out[33][644],u_xpb_out[34][644],u_xpb_out[35][644],u_xpb_out[36][644],u_xpb_out[37][644],u_xpb_out[38][644],u_xpb_out[39][644],u_xpb_out[40][644],u_xpb_out[41][644],u_xpb_out[42][644],u_xpb_out[43][644],u_xpb_out[44][644],u_xpb_out[45][644],u_xpb_out[46][644],u_xpb_out[47][644],u_xpb_out[48][644],u_xpb_out[49][644],u_xpb_out[50][644],u_xpb_out[51][644],u_xpb_out[52][644],u_xpb_out[53][644],u_xpb_out[54][644],u_xpb_out[55][644],u_xpb_out[56][644],u_xpb_out[57][644],u_xpb_out[58][644],u_xpb_out[59][644],u_xpb_out[60][644],u_xpb_out[61][644],u_xpb_out[62][644],u_xpb_out[63][644],u_xpb_out[64][644],u_xpb_out[65][644],u_xpb_out[66][644],u_xpb_out[67][644],u_xpb_out[68][644],u_xpb_out[69][644],u_xpb_out[70][644],u_xpb_out[71][644],u_xpb_out[72][644],u_xpb_out[73][644],u_xpb_out[74][644],u_xpb_out[75][644],u_xpb_out[76][644],u_xpb_out[77][644],u_xpb_out[78][644],u_xpb_out[79][644],u_xpb_out[80][644],u_xpb_out[81][644],u_xpb_out[82][644],u_xpb_out[83][644],u_xpb_out[84][644],u_xpb_out[85][644],u_xpb_out[86][644],u_xpb_out[87][644],u_xpb_out[88][644],u_xpb_out[89][644],u_xpb_out[90][644],u_xpb_out[91][644],u_xpb_out[92][644],u_xpb_out[93][644],u_xpb_out[94][644],u_xpb_out[95][644],u_xpb_out[96][644],u_xpb_out[97][644],u_xpb_out[98][644],u_xpb_out[99][644],u_xpb_out[100][644],u_xpb_out[101][644],u_xpb_out[102][644],u_xpb_out[103][644],u_xpb_out[104][644],u_xpb_out[105][644]};

assign col_out_645 = {u_xpb_out[0][645],u_xpb_out[1][645],u_xpb_out[2][645],u_xpb_out[3][645],u_xpb_out[4][645],u_xpb_out[5][645],u_xpb_out[6][645],u_xpb_out[7][645],u_xpb_out[8][645],u_xpb_out[9][645],u_xpb_out[10][645],u_xpb_out[11][645],u_xpb_out[12][645],u_xpb_out[13][645],u_xpb_out[14][645],u_xpb_out[15][645],u_xpb_out[16][645],u_xpb_out[17][645],u_xpb_out[18][645],u_xpb_out[19][645],u_xpb_out[20][645],u_xpb_out[21][645],u_xpb_out[22][645],u_xpb_out[23][645],u_xpb_out[24][645],u_xpb_out[25][645],u_xpb_out[26][645],u_xpb_out[27][645],u_xpb_out[28][645],u_xpb_out[29][645],u_xpb_out[30][645],u_xpb_out[31][645],u_xpb_out[32][645],u_xpb_out[33][645],u_xpb_out[34][645],u_xpb_out[35][645],u_xpb_out[36][645],u_xpb_out[37][645],u_xpb_out[38][645],u_xpb_out[39][645],u_xpb_out[40][645],u_xpb_out[41][645],u_xpb_out[42][645],u_xpb_out[43][645],u_xpb_out[44][645],u_xpb_out[45][645],u_xpb_out[46][645],u_xpb_out[47][645],u_xpb_out[48][645],u_xpb_out[49][645],u_xpb_out[50][645],u_xpb_out[51][645],u_xpb_out[52][645],u_xpb_out[53][645],u_xpb_out[54][645],u_xpb_out[55][645],u_xpb_out[56][645],u_xpb_out[57][645],u_xpb_out[58][645],u_xpb_out[59][645],u_xpb_out[60][645],u_xpb_out[61][645],u_xpb_out[62][645],u_xpb_out[63][645],u_xpb_out[64][645],u_xpb_out[65][645],u_xpb_out[66][645],u_xpb_out[67][645],u_xpb_out[68][645],u_xpb_out[69][645],u_xpb_out[70][645],u_xpb_out[71][645],u_xpb_out[72][645],u_xpb_out[73][645],u_xpb_out[74][645],u_xpb_out[75][645],u_xpb_out[76][645],u_xpb_out[77][645],u_xpb_out[78][645],u_xpb_out[79][645],u_xpb_out[80][645],u_xpb_out[81][645],u_xpb_out[82][645],u_xpb_out[83][645],u_xpb_out[84][645],u_xpb_out[85][645],u_xpb_out[86][645],u_xpb_out[87][645],u_xpb_out[88][645],u_xpb_out[89][645],u_xpb_out[90][645],u_xpb_out[91][645],u_xpb_out[92][645],u_xpb_out[93][645],u_xpb_out[94][645],u_xpb_out[95][645],u_xpb_out[96][645],u_xpb_out[97][645],u_xpb_out[98][645],u_xpb_out[99][645],u_xpb_out[100][645],u_xpb_out[101][645],u_xpb_out[102][645],u_xpb_out[103][645],u_xpb_out[104][645],u_xpb_out[105][645]};

assign col_out_646 = {u_xpb_out[0][646],u_xpb_out[1][646],u_xpb_out[2][646],u_xpb_out[3][646],u_xpb_out[4][646],u_xpb_out[5][646],u_xpb_out[6][646],u_xpb_out[7][646],u_xpb_out[8][646],u_xpb_out[9][646],u_xpb_out[10][646],u_xpb_out[11][646],u_xpb_out[12][646],u_xpb_out[13][646],u_xpb_out[14][646],u_xpb_out[15][646],u_xpb_out[16][646],u_xpb_out[17][646],u_xpb_out[18][646],u_xpb_out[19][646],u_xpb_out[20][646],u_xpb_out[21][646],u_xpb_out[22][646],u_xpb_out[23][646],u_xpb_out[24][646],u_xpb_out[25][646],u_xpb_out[26][646],u_xpb_out[27][646],u_xpb_out[28][646],u_xpb_out[29][646],u_xpb_out[30][646],u_xpb_out[31][646],u_xpb_out[32][646],u_xpb_out[33][646],u_xpb_out[34][646],u_xpb_out[35][646],u_xpb_out[36][646],u_xpb_out[37][646],u_xpb_out[38][646],u_xpb_out[39][646],u_xpb_out[40][646],u_xpb_out[41][646],u_xpb_out[42][646],u_xpb_out[43][646],u_xpb_out[44][646],u_xpb_out[45][646],u_xpb_out[46][646],u_xpb_out[47][646],u_xpb_out[48][646],u_xpb_out[49][646],u_xpb_out[50][646],u_xpb_out[51][646],u_xpb_out[52][646],u_xpb_out[53][646],u_xpb_out[54][646],u_xpb_out[55][646],u_xpb_out[56][646],u_xpb_out[57][646],u_xpb_out[58][646],u_xpb_out[59][646],u_xpb_out[60][646],u_xpb_out[61][646],u_xpb_out[62][646],u_xpb_out[63][646],u_xpb_out[64][646],u_xpb_out[65][646],u_xpb_out[66][646],u_xpb_out[67][646],u_xpb_out[68][646],u_xpb_out[69][646],u_xpb_out[70][646],u_xpb_out[71][646],u_xpb_out[72][646],u_xpb_out[73][646],u_xpb_out[74][646],u_xpb_out[75][646],u_xpb_out[76][646],u_xpb_out[77][646],u_xpb_out[78][646],u_xpb_out[79][646],u_xpb_out[80][646],u_xpb_out[81][646],u_xpb_out[82][646],u_xpb_out[83][646],u_xpb_out[84][646],u_xpb_out[85][646],u_xpb_out[86][646],u_xpb_out[87][646],u_xpb_out[88][646],u_xpb_out[89][646],u_xpb_out[90][646],u_xpb_out[91][646],u_xpb_out[92][646],u_xpb_out[93][646],u_xpb_out[94][646],u_xpb_out[95][646],u_xpb_out[96][646],u_xpb_out[97][646],u_xpb_out[98][646],u_xpb_out[99][646],u_xpb_out[100][646],u_xpb_out[101][646],u_xpb_out[102][646],u_xpb_out[103][646],u_xpb_out[104][646],u_xpb_out[105][646]};

assign col_out_647 = {u_xpb_out[0][647],u_xpb_out[1][647],u_xpb_out[2][647],u_xpb_out[3][647],u_xpb_out[4][647],u_xpb_out[5][647],u_xpb_out[6][647],u_xpb_out[7][647],u_xpb_out[8][647],u_xpb_out[9][647],u_xpb_out[10][647],u_xpb_out[11][647],u_xpb_out[12][647],u_xpb_out[13][647],u_xpb_out[14][647],u_xpb_out[15][647],u_xpb_out[16][647],u_xpb_out[17][647],u_xpb_out[18][647],u_xpb_out[19][647],u_xpb_out[20][647],u_xpb_out[21][647],u_xpb_out[22][647],u_xpb_out[23][647],u_xpb_out[24][647],u_xpb_out[25][647],u_xpb_out[26][647],u_xpb_out[27][647],u_xpb_out[28][647],u_xpb_out[29][647],u_xpb_out[30][647],u_xpb_out[31][647],u_xpb_out[32][647],u_xpb_out[33][647],u_xpb_out[34][647],u_xpb_out[35][647],u_xpb_out[36][647],u_xpb_out[37][647],u_xpb_out[38][647],u_xpb_out[39][647],u_xpb_out[40][647],u_xpb_out[41][647],u_xpb_out[42][647],u_xpb_out[43][647],u_xpb_out[44][647],u_xpb_out[45][647],u_xpb_out[46][647],u_xpb_out[47][647],u_xpb_out[48][647],u_xpb_out[49][647],u_xpb_out[50][647],u_xpb_out[51][647],u_xpb_out[52][647],u_xpb_out[53][647],u_xpb_out[54][647],u_xpb_out[55][647],u_xpb_out[56][647],u_xpb_out[57][647],u_xpb_out[58][647],u_xpb_out[59][647],u_xpb_out[60][647],u_xpb_out[61][647],u_xpb_out[62][647],u_xpb_out[63][647],u_xpb_out[64][647],u_xpb_out[65][647],u_xpb_out[66][647],u_xpb_out[67][647],u_xpb_out[68][647],u_xpb_out[69][647],u_xpb_out[70][647],u_xpb_out[71][647],u_xpb_out[72][647],u_xpb_out[73][647],u_xpb_out[74][647],u_xpb_out[75][647],u_xpb_out[76][647],u_xpb_out[77][647],u_xpb_out[78][647],u_xpb_out[79][647],u_xpb_out[80][647],u_xpb_out[81][647],u_xpb_out[82][647],u_xpb_out[83][647],u_xpb_out[84][647],u_xpb_out[85][647],u_xpb_out[86][647],u_xpb_out[87][647],u_xpb_out[88][647],u_xpb_out[89][647],u_xpb_out[90][647],u_xpb_out[91][647],u_xpb_out[92][647],u_xpb_out[93][647],u_xpb_out[94][647],u_xpb_out[95][647],u_xpb_out[96][647],u_xpb_out[97][647],u_xpb_out[98][647],u_xpb_out[99][647],u_xpb_out[100][647],u_xpb_out[101][647],u_xpb_out[102][647],u_xpb_out[103][647],u_xpb_out[104][647],u_xpb_out[105][647]};

assign col_out_648 = {u_xpb_out[0][648],u_xpb_out[1][648],u_xpb_out[2][648],u_xpb_out[3][648],u_xpb_out[4][648],u_xpb_out[5][648],u_xpb_out[6][648],u_xpb_out[7][648],u_xpb_out[8][648],u_xpb_out[9][648],u_xpb_out[10][648],u_xpb_out[11][648],u_xpb_out[12][648],u_xpb_out[13][648],u_xpb_out[14][648],u_xpb_out[15][648],u_xpb_out[16][648],u_xpb_out[17][648],u_xpb_out[18][648],u_xpb_out[19][648],u_xpb_out[20][648],u_xpb_out[21][648],u_xpb_out[22][648],u_xpb_out[23][648],u_xpb_out[24][648],u_xpb_out[25][648],u_xpb_out[26][648],u_xpb_out[27][648],u_xpb_out[28][648],u_xpb_out[29][648],u_xpb_out[30][648],u_xpb_out[31][648],u_xpb_out[32][648],u_xpb_out[33][648],u_xpb_out[34][648],u_xpb_out[35][648],u_xpb_out[36][648],u_xpb_out[37][648],u_xpb_out[38][648],u_xpb_out[39][648],u_xpb_out[40][648],u_xpb_out[41][648],u_xpb_out[42][648],u_xpb_out[43][648],u_xpb_out[44][648],u_xpb_out[45][648],u_xpb_out[46][648],u_xpb_out[47][648],u_xpb_out[48][648],u_xpb_out[49][648],u_xpb_out[50][648],u_xpb_out[51][648],u_xpb_out[52][648],u_xpb_out[53][648],u_xpb_out[54][648],u_xpb_out[55][648],u_xpb_out[56][648],u_xpb_out[57][648],u_xpb_out[58][648],u_xpb_out[59][648],u_xpb_out[60][648],u_xpb_out[61][648],u_xpb_out[62][648],u_xpb_out[63][648],u_xpb_out[64][648],u_xpb_out[65][648],u_xpb_out[66][648],u_xpb_out[67][648],u_xpb_out[68][648],u_xpb_out[69][648],u_xpb_out[70][648],u_xpb_out[71][648],u_xpb_out[72][648],u_xpb_out[73][648],u_xpb_out[74][648],u_xpb_out[75][648],u_xpb_out[76][648],u_xpb_out[77][648],u_xpb_out[78][648],u_xpb_out[79][648],u_xpb_out[80][648],u_xpb_out[81][648],u_xpb_out[82][648],u_xpb_out[83][648],u_xpb_out[84][648],u_xpb_out[85][648],u_xpb_out[86][648],u_xpb_out[87][648],u_xpb_out[88][648],u_xpb_out[89][648],u_xpb_out[90][648],u_xpb_out[91][648],u_xpb_out[92][648],u_xpb_out[93][648],u_xpb_out[94][648],u_xpb_out[95][648],u_xpb_out[96][648],u_xpb_out[97][648],u_xpb_out[98][648],u_xpb_out[99][648],u_xpb_out[100][648],u_xpb_out[101][648],u_xpb_out[102][648],u_xpb_out[103][648],u_xpb_out[104][648],u_xpb_out[105][648]};

assign col_out_649 = {u_xpb_out[0][649],u_xpb_out[1][649],u_xpb_out[2][649],u_xpb_out[3][649],u_xpb_out[4][649],u_xpb_out[5][649],u_xpb_out[6][649],u_xpb_out[7][649],u_xpb_out[8][649],u_xpb_out[9][649],u_xpb_out[10][649],u_xpb_out[11][649],u_xpb_out[12][649],u_xpb_out[13][649],u_xpb_out[14][649],u_xpb_out[15][649],u_xpb_out[16][649],u_xpb_out[17][649],u_xpb_out[18][649],u_xpb_out[19][649],u_xpb_out[20][649],u_xpb_out[21][649],u_xpb_out[22][649],u_xpb_out[23][649],u_xpb_out[24][649],u_xpb_out[25][649],u_xpb_out[26][649],u_xpb_out[27][649],u_xpb_out[28][649],u_xpb_out[29][649],u_xpb_out[30][649],u_xpb_out[31][649],u_xpb_out[32][649],u_xpb_out[33][649],u_xpb_out[34][649],u_xpb_out[35][649],u_xpb_out[36][649],u_xpb_out[37][649],u_xpb_out[38][649],u_xpb_out[39][649],u_xpb_out[40][649],u_xpb_out[41][649],u_xpb_out[42][649],u_xpb_out[43][649],u_xpb_out[44][649],u_xpb_out[45][649],u_xpb_out[46][649],u_xpb_out[47][649],u_xpb_out[48][649],u_xpb_out[49][649],u_xpb_out[50][649],u_xpb_out[51][649],u_xpb_out[52][649],u_xpb_out[53][649],u_xpb_out[54][649],u_xpb_out[55][649],u_xpb_out[56][649],u_xpb_out[57][649],u_xpb_out[58][649],u_xpb_out[59][649],u_xpb_out[60][649],u_xpb_out[61][649],u_xpb_out[62][649],u_xpb_out[63][649],u_xpb_out[64][649],u_xpb_out[65][649],u_xpb_out[66][649],u_xpb_out[67][649],u_xpb_out[68][649],u_xpb_out[69][649],u_xpb_out[70][649],u_xpb_out[71][649],u_xpb_out[72][649],u_xpb_out[73][649],u_xpb_out[74][649],u_xpb_out[75][649],u_xpb_out[76][649],u_xpb_out[77][649],u_xpb_out[78][649],u_xpb_out[79][649],u_xpb_out[80][649],u_xpb_out[81][649],u_xpb_out[82][649],u_xpb_out[83][649],u_xpb_out[84][649],u_xpb_out[85][649],u_xpb_out[86][649],u_xpb_out[87][649],u_xpb_out[88][649],u_xpb_out[89][649],u_xpb_out[90][649],u_xpb_out[91][649],u_xpb_out[92][649],u_xpb_out[93][649],u_xpb_out[94][649],u_xpb_out[95][649],u_xpb_out[96][649],u_xpb_out[97][649],u_xpb_out[98][649],u_xpb_out[99][649],u_xpb_out[100][649],u_xpb_out[101][649],u_xpb_out[102][649],u_xpb_out[103][649],u_xpb_out[104][649],u_xpb_out[105][649]};

assign col_out_650 = {u_xpb_out[0][650],u_xpb_out[1][650],u_xpb_out[2][650],u_xpb_out[3][650],u_xpb_out[4][650],u_xpb_out[5][650],u_xpb_out[6][650],u_xpb_out[7][650],u_xpb_out[8][650],u_xpb_out[9][650],u_xpb_out[10][650],u_xpb_out[11][650],u_xpb_out[12][650],u_xpb_out[13][650],u_xpb_out[14][650],u_xpb_out[15][650],u_xpb_out[16][650],u_xpb_out[17][650],u_xpb_out[18][650],u_xpb_out[19][650],u_xpb_out[20][650],u_xpb_out[21][650],u_xpb_out[22][650],u_xpb_out[23][650],u_xpb_out[24][650],u_xpb_out[25][650],u_xpb_out[26][650],u_xpb_out[27][650],u_xpb_out[28][650],u_xpb_out[29][650],u_xpb_out[30][650],u_xpb_out[31][650],u_xpb_out[32][650],u_xpb_out[33][650],u_xpb_out[34][650],u_xpb_out[35][650],u_xpb_out[36][650],u_xpb_out[37][650],u_xpb_out[38][650],u_xpb_out[39][650],u_xpb_out[40][650],u_xpb_out[41][650],u_xpb_out[42][650],u_xpb_out[43][650],u_xpb_out[44][650],u_xpb_out[45][650],u_xpb_out[46][650],u_xpb_out[47][650],u_xpb_out[48][650],u_xpb_out[49][650],u_xpb_out[50][650],u_xpb_out[51][650],u_xpb_out[52][650],u_xpb_out[53][650],u_xpb_out[54][650],u_xpb_out[55][650],u_xpb_out[56][650],u_xpb_out[57][650],u_xpb_out[58][650],u_xpb_out[59][650],u_xpb_out[60][650],u_xpb_out[61][650],u_xpb_out[62][650],u_xpb_out[63][650],u_xpb_out[64][650],u_xpb_out[65][650],u_xpb_out[66][650],u_xpb_out[67][650],u_xpb_out[68][650],u_xpb_out[69][650],u_xpb_out[70][650],u_xpb_out[71][650],u_xpb_out[72][650],u_xpb_out[73][650],u_xpb_out[74][650],u_xpb_out[75][650],u_xpb_out[76][650],u_xpb_out[77][650],u_xpb_out[78][650],u_xpb_out[79][650],u_xpb_out[80][650],u_xpb_out[81][650],u_xpb_out[82][650],u_xpb_out[83][650],u_xpb_out[84][650],u_xpb_out[85][650],u_xpb_out[86][650],u_xpb_out[87][650],u_xpb_out[88][650],u_xpb_out[89][650],u_xpb_out[90][650],u_xpb_out[91][650],u_xpb_out[92][650],u_xpb_out[93][650],u_xpb_out[94][650],u_xpb_out[95][650],u_xpb_out[96][650],u_xpb_out[97][650],u_xpb_out[98][650],u_xpb_out[99][650],u_xpb_out[100][650],u_xpb_out[101][650],u_xpb_out[102][650],u_xpb_out[103][650],u_xpb_out[104][650],u_xpb_out[105][650]};

assign col_out_651 = {u_xpb_out[0][651],u_xpb_out[1][651],u_xpb_out[2][651],u_xpb_out[3][651],u_xpb_out[4][651],u_xpb_out[5][651],u_xpb_out[6][651],u_xpb_out[7][651],u_xpb_out[8][651],u_xpb_out[9][651],u_xpb_out[10][651],u_xpb_out[11][651],u_xpb_out[12][651],u_xpb_out[13][651],u_xpb_out[14][651],u_xpb_out[15][651],u_xpb_out[16][651],u_xpb_out[17][651],u_xpb_out[18][651],u_xpb_out[19][651],u_xpb_out[20][651],u_xpb_out[21][651],u_xpb_out[22][651],u_xpb_out[23][651],u_xpb_out[24][651],u_xpb_out[25][651],u_xpb_out[26][651],u_xpb_out[27][651],u_xpb_out[28][651],u_xpb_out[29][651],u_xpb_out[30][651],u_xpb_out[31][651],u_xpb_out[32][651],u_xpb_out[33][651],u_xpb_out[34][651],u_xpb_out[35][651],u_xpb_out[36][651],u_xpb_out[37][651],u_xpb_out[38][651],u_xpb_out[39][651],u_xpb_out[40][651],u_xpb_out[41][651],u_xpb_out[42][651],u_xpb_out[43][651],u_xpb_out[44][651],u_xpb_out[45][651],u_xpb_out[46][651],u_xpb_out[47][651],u_xpb_out[48][651],u_xpb_out[49][651],u_xpb_out[50][651],u_xpb_out[51][651],u_xpb_out[52][651],u_xpb_out[53][651],u_xpb_out[54][651],u_xpb_out[55][651],u_xpb_out[56][651],u_xpb_out[57][651],u_xpb_out[58][651],u_xpb_out[59][651],u_xpb_out[60][651],u_xpb_out[61][651],u_xpb_out[62][651],u_xpb_out[63][651],u_xpb_out[64][651],u_xpb_out[65][651],u_xpb_out[66][651],u_xpb_out[67][651],u_xpb_out[68][651],u_xpb_out[69][651],u_xpb_out[70][651],u_xpb_out[71][651],u_xpb_out[72][651],u_xpb_out[73][651],u_xpb_out[74][651],u_xpb_out[75][651],u_xpb_out[76][651],u_xpb_out[77][651],u_xpb_out[78][651],u_xpb_out[79][651],u_xpb_out[80][651],u_xpb_out[81][651],u_xpb_out[82][651],u_xpb_out[83][651],u_xpb_out[84][651],u_xpb_out[85][651],u_xpb_out[86][651],u_xpb_out[87][651],u_xpb_out[88][651],u_xpb_out[89][651],u_xpb_out[90][651],u_xpb_out[91][651],u_xpb_out[92][651],u_xpb_out[93][651],u_xpb_out[94][651],u_xpb_out[95][651],u_xpb_out[96][651],u_xpb_out[97][651],u_xpb_out[98][651],u_xpb_out[99][651],u_xpb_out[100][651],u_xpb_out[101][651],u_xpb_out[102][651],u_xpb_out[103][651],u_xpb_out[104][651],u_xpb_out[105][651]};

assign col_out_652 = {u_xpb_out[0][652],u_xpb_out[1][652],u_xpb_out[2][652],u_xpb_out[3][652],u_xpb_out[4][652],u_xpb_out[5][652],u_xpb_out[6][652],u_xpb_out[7][652],u_xpb_out[8][652],u_xpb_out[9][652],u_xpb_out[10][652],u_xpb_out[11][652],u_xpb_out[12][652],u_xpb_out[13][652],u_xpb_out[14][652],u_xpb_out[15][652],u_xpb_out[16][652],u_xpb_out[17][652],u_xpb_out[18][652],u_xpb_out[19][652],u_xpb_out[20][652],u_xpb_out[21][652],u_xpb_out[22][652],u_xpb_out[23][652],u_xpb_out[24][652],u_xpb_out[25][652],u_xpb_out[26][652],u_xpb_out[27][652],u_xpb_out[28][652],u_xpb_out[29][652],u_xpb_out[30][652],u_xpb_out[31][652],u_xpb_out[32][652],u_xpb_out[33][652],u_xpb_out[34][652],u_xpb_out[35][652],u_xpb_out[36][652],u_xpb_out[37][652],u_xpb_out[38][652],u_xpb_out[39][652],u_xpb_out[40][652],u_xpb_out[41][652],u_xpb_out[42][652],u_xpb_out[43][652],u_xpb_out[44][652],u_xpb_out[45][652],u_xpb_out[46][652],u_xpb_out[47][652],u_xpb_out[48][652],u_xpb_out[49][652],u_xpb_out[50][652],u_xpb_out[51][652],u_xpb_out[52][652],u_xpb_out[53][652],u_xpb_out[54][652],u_xpb_out[55][652],u_xpb_out[56][652],u_xpb_out[57][652],u_xpb_out[58][652],u_xpb_out[59][652],u_xpb_out[60][652],u_xpb_out[61][652],u_xpb_out[62][652],u_xpb_out[63][652],u_xpb_out[64][652],u_xpb_out[65][652],u_xpb_out[66][652],u_xpb_out[67][652],u_xpb_out[68][652],u_xpb_out[69][652],u_xpb_out[70][652],u_xpb_out[71][652],u_xpb_out[72][652],u_xpb_out[73][652],u_xpb_out[74][652],u_xpb_out[75][652],u_xpb_out[76][652],u_xpb_out[77][652],u_xpb_out[78][652],u_xpb_out[79][652],u_xpb_out[80][652],u_xpb_out[81][652],u_xpb_out[82][652],u_xpb_out[83][652],u_xpb_out[84][652],u_xpb_out[85][652],u_xpb_out[86][652],u_xpb_out[87][652],u_xpb_out[88][652],u_xpb_out[89][652],u_xpb_out[90][652],u_xpb_out[91][652],u_xpb_out[92][652],u_xpb_out[93][652],u_xpb_out[94][652],u_xpb_out[95][652],u_xpb_out[96][652],u_xpb_out[97][652],u_xpb_out[98][652],u_xpb_out[99][652],u_xpb_out[100][652],u_xpb_out[101][652],u_xpb_out[102][652],u_xpb_out[103][652],u_xpb_out[104][652],u_xpb_out[105][652]};

assign col_out_653 = {u_xpb_out[0][653],u_xpb_out[1][653],u_xpb_out[2][653],u_xpb_out[3][653],u_xpb_out[4][653],u_xpb_out[5][653],u_xpb_out[6][653],u_xpb_out[7][653],u_xpb_out[8][653],u_xpb_out[9][653],u_xpb_out[10][653],u_xpb_out[11][653],u_xpb_out[12][653],u_xpb_out[13][653],u_xpb_out[14][653],u_xpb_out[15][653],u_xpb_out[16][653],u_xpb_out[17][653],u_xpb_out[18][653],u_xpb_out[19][653],u_xpb_out[20][653],u_xpb_out[21][653],u_xpb_out[22][653],u_xpb_out[23][653],u_xpb_out[24][653],u_xpb_out[25][653],u_xpb_out[26][653],u_xpb_out[27][653],u_xpb_out[28][653],u_xpb_out[29][653],u_xpb_out[30][653],u_xpb_out[31][653],u_xpb_out[32][653],u_xpb_out[33][653],u_xpb_out[34][653],u_xpb_out[35][653],u_xpb_out[36][653],u_xpb_out[37][653],u_xpb_out[38][653],u_xpb_out[39][653],u_xpb_out[40][653],u_xpb_out[41][653],u_xpb_out[42][653],u_xpb_out[43][653],u_xpb_out[44][653],u_xpb_out[45][653],u_xpb_out[46][653],u_xpb_out[47][653],u_xpb_out[48][653],u_xpb_out[49][653],u_xpb_out[50][653],u_xpb_out[51][653],u_xpb_out[52][653],u_xpb_out[53][653],u_xpb_out[54][653],u_xpb_out[55][653],u_xpb_out[56][653],u_xpb_out[57][653],u_xpb_out[58][653],u_xpb_out[59][653],u_xpb_out[60][653],u_xpb_out[61][653],u_xpb_out[62][653],u_xpb_out[63][653],u_xpb_out[64][653],u_xpb_out[65][653],u_xpb_out[66][653],u_xpb_out[67][653],u_xpb_out[68][653],u_xpb_out[69][653],u_xpb_out[70][653],u_xpb_out[71][653],u_xpb_out[72][653],u_xpb_out[73][653],u_xpb_out[74][653],u_xpb_out[75][653],u_xpb_out[76][653],u_xpb_out[77][653],u_xpb_out[78][653],u_xpb_out[79][653],u_xpb_out[80][653],u_xpb_out[81][653],u_xpb_out[82][653],u_xpb_out[83][653],u_xpb_out[84][653],u_xpb_out[85][653],u_xpb_out[86][653],u_xpb_out[87][653],u_xpb_out[88][653],u_xpb_out[89][653],u_xpb_out[90][653],u_xpb_out[91][653],u_xpb_out[92][653],u_xpb_out[93][653],u_xpb_out[94][653],u_xpb_out[95][653],u_xpb_out[96][653],u_xpb_out[97][653],u_xpb_out[98][653],u_xpb_out[99][653],u_xpb_out[100][653],u_xpb_out[101][653],u_xpb_out[102][653],u_xpb_out[103][653],u_xpb_out[104][653],u_xpb_out[105][653]};

assign col_out_654 = {u_xpb_out[0][654],u_xpb_out[1][654],u_xpb_out[2][654],u_xpb_out[3][654],u_xpb_out[4][654],u_xpb_out[5][654],u_xpb_out[6][654],u_xpb_out[7][654],u_xpb_out[8][654],u_xpb_out[9][654],u_xpb_out[10][654],u_xpb_out[11][654],u_xpb_out[12][654],u_xpb_out[13][654],u_xpb_out[14][654],u_xpb_out[15][654],u_xpb_out[16][654],u_xpb_out[17][654],u_xpb_out[18][654],u_xpb_out[19][654],u_xpb_out[20][654],u_xpb_out[21][654],u_xpb_out[22][654],u_xpb_out[23][654],u_xpb_out[24][654],u_xpb_out[25][654],u_xpb_out[26][654],u_xpb_out[27][654],u_xpb_out[28][654],u_xpb_out[29][654],u_xpb_out[30][654],u_xpb_out[31][654],u_xpb_out[32][654],u_xpb_out[33][654],u_xpb_out[34][654],u_xpb_out[35][654],u_xpb_out[36][654],u_xpb_out[37][654],u_xpb_out[38][654],u_xpb_out[39][654],u_xpb_out[40][654],u_xpb_out[41][654],u_xpb_out[42][654],u_xpb_out[43][654],u_xpb_out[44][654],u_xpb_out[45][654],u_xpb_out[46][654],u_xpb_out[47][654],u_xpb_out[48][654],u_xpb_out[49][654],u_xpb_out[50][654],u_xpb_out[51][654],u_xpb_out[52][654],u_xpb_out[53][654],u_xpb_out[54][654],u_xpb_out[55][654],u_xpb_out[56][654],u_xpb_out[57][654],u_xpb_out[58][654],u_xpb_out[59][654],u_xpb_out[60][654],u_xpb_out[61][654],u_xpb_out[62][654],u_xpb_out[63][654],u_xpb_out[64][654],u_xpb_out[65][654],u_xpb_out[66][654],u_xpb_out[67][654],u_xpb_out[68][654],u_xpb_out[69][654],u_xpb_out[70][654],u_xpb_out[71][654],u_xpb_out[72][654],u_xpb_out[73][654],u_xpb_out[74][654],u_xpb_out[75][654],u_xpb_out[76][654],u_xpb_out[77][654],u_xpb_out[78][654],u_xpb_out[79][654],u_xpb_out[80][654],u_xpb_out[81][654],u_xpb_out[82][654],u_xpb_out[83][654],u_xpb_out[84][654],u_xpb_out[85][654],u_xpb_out[86][654],u_xpb_out[87][654],u_xpb_out[88][654],u_xpb_out[89][654],u_xpb_out[90][654],u_xpb_out[91][654],u_xpb_out[92][654],u_xpb_out[93][654],u_xpb_out[94][654],u_xpb_out[95][654],u_xpb_out[96][654],u_xpb_out[97][654],u_xpb_out[98][654],u_xpb_out[99][654],u_xpb_out[100][654],u_xpb_out[101][654],u_xpb_out[102][654],u_xpb_out[103][654],u_xpb_out[104][654],u_xpb_out[105][654]};

assign col_out_655 = {u_xpb_out[0][655],u_xpb_out[1][655],u_xpb_out[2][655],u_xpb_out[3][655],u_xpb_out[4][655],u_xpb_out[5][655],u_xpb_out[6][655],u_xpb_out[7][655],u_xpb_out[8][655],u_xpb_out[9][655],u_xpb_out[10][655],u_xpb_out[11][655],u_xpb_out[12][655],u_xpb_out[13][655],u_xpb_out[14][655],u_xpb_out[15][655],u_xpb_out[16][655],u_xpb_out[17][655],u_xpb_out[18][655],u_xpb_out[19][655],u_xpb_out[20][655],u_xpb_out[21][655],u_xpb_out[22][655],u_xpb_out[23][655],u_xpb_out[24][655],u_xpb_out[25][655],u_xpb_out[26][655],u_xpb_out[27][655],u_xpb_out[28][655],u_xpb_out[29][655],u_xpb_out[30][655],u_xpb_out[31][655],u_xpb_out[32][655],u_xpb_out[33][655],u_xpb_out[34][655],u_xpb_out[35][655],u_xpb_out[36][655],u_xpb_out[37][655],u_xpb_out[38][655],u_xpb_out[39][655],u_xpb_out[40][655],u_xpb_out[41][655],u_xpb_out[42][655],u_xpb_out[43][655],u_xpb_out[44][655],u_xpb_out[45][655],u_xpb_out[46][655],u_xpb_out[47][655],u_xpb_out[48][655],u_xpb_out[49][655],u_xpb_out[50][655],u_xpb_out[51][655],u_xpb_out[52][655],u_xpb_out[53][655],u_xpb_out[54][655],u_xpb_out[55][655],u_xpb_out[56][655],u_xpb_out[57][655],u_xpb_out[58][655],u_xpb_out[59][655],u_xpb_out[60][655],u_xpb_out[61][655],u_xpb_out[62][655],u_xpb_out[63][655],u_xpb_out[64][655],u_xpb_out[65][655],u_xpb_out[66][655],u_xpb_out[67][655],u_xpb_out[68][655],u_xpb_out[69][655],u_xpb_out[70][655],u_xpb_out[71][655],u_xpb_out[72][655],u_xpb_out[73][655],u_xpb_out[74][655],u_xpb_out[75][655],u_xpb_out[76][655],u_xpb_out[77][655],u_xpb_out[78][655],u_xpb_out[79][655],u_xpb_out[80][655],u_xpb_out[81][655],u_xpb_out[82][655],u_xpb_out[83][655],u_xpb_out[84][655],u_xpb_out[85][655],u_xpb_out[86][655],u_xpb_out[87][655],u_xpb_out[88][655],u_xpb_out[89][655],u_xpb_out[90][655],u_xpb_out[91][655],u_xpb_out[92][655],u_xpb_out[93][655],u_xpb_out[94][655],u_xpb_out[95][655],u_xpb_out[96][655],u_xpb_out[97][655],u_xpb_out[98][655],u_xpb_out[99][655],u_xpb_out[100][655],u_xpb_out[101][655],u_xpb_out[102][655],u_xpb_out[103][655],u_xpb_out[104][655],u_xpb_out[105][655]};

assign col_out_656 = {u_xpb_out[0][656],u_xpb_out[1][656],u_xpb_out[2][656],u_xpb_out[3][656],u_xpb_out[4][656],u_xpb_out[5][656],u_xpb_out[6][656],u_xpb_out[7][656],u_xpb_out[8][656],u_xpb_out[9][656],u_xpb_out[10][656],u_xpb_out[11][656],u_xpb_out[12][656],u_xpb_out[13][656],u_xpb_out[14][656],u_xpb_out[15][656],u_xpb_out[16][656],u_xpb_out[17][656],u_xpb_out[18][656],u_xpb_out[19][656],u_xpb_out[20][656],u_xpb_out[21][656],u_xpb_out[22][656],u_xpb_out[23][656],u_xpb_out[24][656],u_xpb_out[25][656],u_xpb_out[26][656],u_xpb_out[27][656],u_xpb_out[28][656],u_xpb_out[29][656],u_xpb_out[30][656],u_xpb_out[31][656],u_xpb_out[32][656],u_xpb_out[33][656],u_xpb_out[34][656],u_xpb_out[35][656],u_xpb_out[36][656],u_xpb_out[37][656],u_xpb_out[38][656],u_xpb_out[39][656],u_xpb_out[40][656],u_xpb_out[41][656],u_xpb_out[42][656],u_xpb_out[43][656],u_xpb_out[44][656],u_xpb_out[45][656],u_xpb_out[46][656],u_xpb_out[47][656],u_xpb_out[48][656],u_xpb_out[49][656],u_xpb_out[50][656],u_xpb_out[51][656],u_xpb_out[52][656],u_xpb_out[53][656],u_xpb_out[54][656],u_xpb_out[55][656],u_xpb_out[56][656],u_xpb_out[57][656],u_xpb_out[58][656],u_xpb_out[59][656],u_xpb_out[60][656],u_xpb_out[61][656],u_xpb_out[62][656],u_xpb_out[63][656],u_xpb_out[64][656],u_xpb_out[65][656],u_xpb_out[66][656],u_xpb_out[67][656],u_xpb_out[68][656],u_xpb_out[69][656],u_xpb_out[70][656],u_xpb_out[71][656],u_xpb_out[72][656],u_xpb_out[73][656],u_xpb_out[74][656],u_xpb_out[75][656],u_xpb_out[76][656],u_xpb_out[77][656],u_xpb_out[78][656],u_xpb_out[79][656],u_xpb_out[80][656],u_xpb_out[81][656],u_xpb_out[82][656],u_xpb_out[83][656],u_xpb_out[84][656],u_xpb_out[85][656],u_xpb_out[86][656],u_xpb_out[87][656],u_xpb_out[88][656],u_xpb_out[89][656],u_xpb_out[90][656],u_xpb_out[91][656],u_xpb_out[92][656],u_xpb_out[93][656],u_xpb_out[94][656],u_xpb_out[95][656],u_xpb_out[96][656],u_xpb_out[97][656],u_xpb_out[98][656],u_xpb_out[99][656],u_xpb_out[100][656],u_xpb_out[101][656],u_xpb_out[102][656],u_xpb_out[103][656],u_xpb_out[104][656],u_xpb_out[105][656]};

assign col_out_657 = {u_xpb_out[0][657],u_xpb_out[1][657],u_xpb_out[2][657],u_xpb_out[3][657],u_xpb_out[4][657],u_xpb_out[5][657],u_xpb_out[6][657],u_xpb_out[7][657],u_xpb_out[8][657],u_xpb_out[9][657],u_xpb_out[10][657],u_xpb_out[11][657],u_xpb_out[12][657],u_xpb_out[13][657],u_xpb_out[14][657],u_xpb_out[15][657],u_xpb_out[16][657],u_xpb_out[17][657],u_xpb_out[18][657],u_xpb_out[19][657],u_xpb_out[20][657],u_xpb_out[21][657],u_xpb_out[22][657],u_xpb_out[23][657],u_xpb_out[24][657],u_xpb_out[25][657],u_xpb_out[26][657],u_xpb_out[27][657],u_xpb_out[28][657],u_xpb_out[29][657],u_xpb_out[30][657],u_xpb_out[31][657],u_xpb_out[32][657],u_xpb_out[33][657],u_xpb_out[34][657],u_xpb_out[35][657],u_xpb_out[36][657],u_xpb_out[37][657],u_xpb_out[38][657],u_xpb_out[39][657],u_xpb_out[40][657],u_xpb_out[41][657],u_xpb_out[42][657],u_xpb_out[43][657],u_xpb_out[44][657],u_xpb_out[45][657],u_xpb_out[46][657],u_xpb_out[47][657],u_xpb_out[48][657],u_xpb_out[49][657],u_xpb_out[50][657],u_xpb_out[51][657],u_xpb_out[52][657],u_xpb_out[53][657],u_xpb_out[54][657],u_xpb_out[55][657],u_xpb_out[56][657],u_xpb_out[57][657],u_xpb_out[58][657],u_xpb_out[59][657],u_xpb_out[60][657],u_xpb_out[61][657],u_xpb_out[62][657],u_xpb_out[63][657],u_xpb_out[64][657],u_xpb_out[65][657],u_xpb_out[66][657],u_xpb_out[67][657],u_xpb_out[68][657],u_xpb_out[69][657],u_xpb_out[70][657],u_xpb_out[71][657],u_xpb_out[72][657],u_xpb_out[73][657],u_xpb_out[74][657],u_xpb_out[75][657],u_xpb_out[76][657],u_xpb_out[77][657],u_xpb_out[78][657],u_xpb_out[79][657],u_xpb_out[80][657],u_xpb_out[81][657],u_xpb_out[82][657],u_xpb_out[83][657],u_xpb_out[84][657],u_xpb_out[85][657],u_xpb_out[86][657],u_xpb_out[87][657],u_xpb_out[88][657],u_xpb_out[89][657],u_xpb_out[90][657],u_xpb_out[91][657],u_xpb_out[92][657],u_xpb_out[93][657],u_xpb_out[94][657],u_xpb_out[95][657],u_xpb_out[96][657],u_xpb_out[97][657],u_xpb_out[98][657],u_xpb_out[99][657],u_xpb_out[100][657],u_xpb_out[101][657],u_xpb_out[102][657],u_xpb_out[103][657],u_xpb_out[104][657],u_xpb_out[105][657]};

assign col_out_658 = {u_xpb_out[0][658],u_xpb_out[1][658],u_xpb_out[2][658],u_xpb_out[3][658],u_xpb_out[4][658],u_xpb_out[5][658],u_xpb_out[6][658],u_xpb_out[7][658],u_xpb_out[8][658],u_xpb_out[9][658],u_xpb_out[10][658],u_xpb_out[11][658],u_xpb_out[12][658],u_xpb_out[13][658],u_xpb_out[14][658],u_xpb_out[15][658],u_xpb_out[16][658],u_xpb_out[17][658],u_xpb_out[18][658],u_xpb_out[19][658],u_xpb_out[20][658],u_xpb_out[21][658],u_xpb_out[22][658],u_xpb_out[23][658],u_xpb_out[24][658],u_xpb_out[25][658],u_xpb_out[26][658],u_xpb_out[27][658],u_xpb_out[28][658],u_xpb_out[29][658],u_xpb_out[30][658],u_xpb_out[31][658],u_xpb_out[32][658],u_xpb_out[33][658],u_xpb_out[34][658],u_xpb_out[35][658],u_xpb_out[36][658],u_xpb_out[37][658],u_xpb_out[38][658],u_xpb_out[39][658],u_xpb_out[40][658],u_xpb_out[41][658],u_xpb_out[42][658],u_xpb_out[43][658],u_xpb_out[44][658],u_xpb_out[45][658],u_xpb_out[46][658],u_xpb_out[47][658],u_xpb_out[48][658],u_xpb_out[49][658],u_xpb_out[50][658],u_xpb_out[51][658],u_xpb_out[52][658],u_xpb_out[53][658],u_xpb_out[54][658],u_xpb_out[55][658],u_xpb_out[56][658],u_xpb_out[57][658],u_xpb_out[58][658],u_xpb_out[59][658],u_xpb_out[60][658],u_xpb_out[61][658],u_xpb_out[62][658],u_xpb_out[63][658],u_xpb_out[64][658],u_xpb_out[65][658],u_xpb_out[66][658],u_xpb_out[67][658],u_xpb_out[68][658],u_xpb_out[69][658],u_xpb_out[70][658],u_xpb_out[71][658],u_xpb_out[72][658],u_xpb_out[73][658],u_xpb_out[74][658],u_xpb_out[75][658],u_xpb_out[76][658],u_xpb_out[77][658],u_xpb_out[78][658],u_xpb_out[79][658],u_xpb_out[80][658],u_xpb_out[81][658],u_xpb_out[82][658],u_xpb_out[83][658],u_xpb_out[84][658],u_xpb_out[85][658],u_xpb_out[86][658],u_xpb_out[87][658],u_xpb_out[88][658],u_xpb_out[89][658],u_xpb_out[90][658],u_xpb_out[91][658],u_xpb_out[92][658],u_xpb_out[93][658],u_xpb_out[94][658],u_xpb_out[95][658],u_xpb_out[96][658],u_xpb_out[97][658],u_xpb_out[98][658],u_xpb_out[99][658],u_xpb_out[100][658],u_xpb_out[101][658],u_xpb_out[102][658],u_xpb_out[103][658],u_xpb_out[104][658],u_xpb_out[105][658]};

assign col_out_659 = {u_xpb_out[0][659],u_xpb_out[1][659],u_xpb_out[2][659],u_xpb_out[3][659],u_xpb_out[4][659],u_xpb_out[5][659],u_xpb_out[6][659],u_xpb_out[7][659],u_xpb_out[8][659],u_xpb_out[9][659],u_xpb_out[10][659],u_xpb_out[11][659],u_xpb_out[12][659],u_xpb_out[13][659],u_xpb_out[14][659],u_xpb_out[15][659],u_xpb_out[16][659],u_xpb_out[17][659],u_xpb_out[18][659],u_xpb_out[19][659],u_xpb_out[20][659],u_xpb_out[21][659],u_xpb_out[22][659],u_xpb_out[23][659],u_xpb_out[24][659],u_xpb_out[25][659],u_xpb_out[26][659],u_xpb_out[27][659],u_xpb_out[28][659],u_xpb_out[29][659],u_xpb_out[30][659],u_xpb_out[31][659],u_xpb_out[32][659],u_xpb_out[33][659],u_xpb_out[34][659],u_xpb_out[35][659],u_xpb_out[36][659],u_xpb_out[37][659],u_xpb_out[38][659],u_xpb_out[39][659],u_xpb_out[40][659],u_xpb_out[41][659],u_xpb_out[42][659],u_xpb_out[43][659],u_xpb_out[44][659],u_xpb_out[45][659],u_xpb_out[46][659],u_xpb_out[47][659],u_xpb_out[48][659],u_xpb_out[49][659],u_xpb_out[50][659],u_xpb_out[51][659],u_xpb_out[52][659],u_xpb_out[53][659],u_xpb_out[54][659],u_xpb_out[55][659],u_xpb_out[56][659],u_xpb_out[57][659],u_xpb_out[58][659],u_xpb_out[59][659],u_xpb_out[60][659],u_xpb_out[61][659],u_xpb_out[62][659],u_xpb_out[63][659],u_xpb_out[64][659],u_xpb_out[65][659],u_xpb_out[66][659],u_xpb_out[67][659],u_xpb_out[68][659],u_xpb_out[69][659],u_xpb_out[70][659],u_xpb_out[71][659],u_xpb_out[72][659],u_xpb_out[73][659],u_xpb_out[74][659],u_xpb_out[75][659],u_xpb_out[76][659],u_xpb_out[77][659],u_xpb_out[78][659],u_xpb_out[79][659],u_xpb_out[80][659],u_xpb_out[81][659],u_xpb_out[82][659],u_xpb_out[83][659],u_xpb_out[84][659],u_xpb_out[85][659],u_xpb_out[86][659],u_xpb_out[87][659],u_xpb_out[88][659],u_xpb_out[89][659],u_xpb_out[90][659],u_xpb_out[91][659],u_xpb_out[92][659],u_xpb_out[93][659],u_xpb_out[94][659],u_xpb_out[95][659],u_xpb_out[96][659],u_xpb_out[97][659],u_xpb_out[98][659],u_xpb_out[99][659],u_xpb_out[100][659],u_xpb_out[101][659],u_xpb_out[102][659],u_xpb_out[103][659],u_xpb_out[104][659],u_xpb_out[105][659]};

assign col_out_660 = {u_xpb_out[0][660],u_xpb_out[1][660],u_xpb_out[2][660],u_xpb_out[3][660],u_xpb_out[4][660],u_xpb_out[5][660],u_xpb_out[6][660],u_xpb_out[7][660],u_xpb_out[8][660],u_xpb_out[9][660],u_xpb_out[10][660],u_xpb_out[11][660],u_xpb_out[12][660],u_xpb_out[13][660],u_xpb_out[14][660],u_xpb_out[15][660],u_xpb_out[16][660],u_xpb_out[17][660],u_xpb_out[18][660],u_xpb_out[19][660],u_xpb_out[20][660],u_xpb_out[21][660],u_xpb_out[22][660],u_xpb_out[23][660],u_xpb_out[24][660],u_xpb_out[25][660],u_xpb_out[26][660],u_xpb_out[27][660],u_xpb_out[28][660],u_xpb_out[29][660],u_xpb_out[30][660],u_xpb_out[31][660],u_xpb_out[32][660],u_xpb_out[33][660],u_xpb_out[34][660],u_xpb_out[35][660],u_xpb_out[36][660],u_xpb_out[37][660],u_xpb_out[38][660],u_xpb_out[39][660],u_xpb_out[40][660],u_xpb_out[41][660],u_xpb_out[42][660],u_xpb_out[43][660],u_xpb_out[44][660],u_xpb_out[45][660],u_xpb_out[46][660],u_xpb_out[47][660],u_xpb_out[48][660],u_xpb_out[49][660],u_xpb_out[50][660],u_xpb_out[51][660],u_xpb_out[52][660],u_xpb_out[53][660],u_xpb_out[54][660],u_xpb_out[55][660],u_xpb_out[56][660],u_xpb_out[57][660],u_xpb_out[58][660],u_xpb_out[59][660],u_xpb_out[60][660],u_xpb_out[61][660],u_xpb_out[62][660],u_xpb_out[63][660],u_xpb_out[64][660],u_xpb_out[65][660],u_xpb_out[66][660],u_xpb_out[67][660],u_xpb_out[68][660],u_xpb_out[69][660],u_xpb_out[70][660],u_xpb_out[71][660],u_xpb_out[72][660],u_xpb_out[73][660],u_xpb_out[74][660],u_xpb_out[75][660],u_xpb_out[76][660],u_xpb_out[77][660],u_xpb_out[78][660],u_xpb_out[79][660],u_xpb_out[80][660],u_xpb_out[81][660],u_xpb_out[82][660],u_xpb_out[83][660],u_xpb_out[84][660],u_xpb_out[85][660],u_xpb_out[86][660],u_xpb_out[87][660],u_xpb_out[88][660],u_xpb_out[89][660],u_xpb_out[90][660],u_xpb_out[91][660],u_xpb_out[92][660],u_xpb_out[93][660],u_xpb_out[94][660],u_xpb_out[95][660],u_xpb_out[96][660],u_xpb_out[97][660],u_xpb_out[98][660],u_xpb_out[99][660],u_xpb_out[100][660],u_xpb_out[101][660],u_xpb_out[102][660],u_xpb_out[103][660],u_xpb_out[104][660],u_xpb_out[105][660]};

assign col_out_661 = {u_xpb_out[0][661],u_xpb_out[1][661],u_xpb_out[2][661],u_xpb_out[3][661],u_xpb_out[4][661],u_xpb_out[5][661],u_xpb_out[6][661],u_xpb_out[7][661],u_xpb_out[8][661],u_xpb_out[9][661],u_xpb_out[10][661],u_xpb_out[11][661],u_xpb_out[12][661],u_xpb_out[13][661],u_xpb_out[14][661],u_xpb_out[15][661],u_xpb_out[16][661],u_xpb_out[17][661],u_xpb_out[18][661],u_xpb_out[19][661],u_xpb_out[20][661],u_xpb_out[21][661],u_xpb_out[22][661],u_xpb_out[23][661],u_xpb_out[24][661],u_xpb_out[25][661],u_xpb_out[26][661],u_xpb_out[27][661],u_xpb_out[28][661],u_xpb_out[29][661],u_xpb_out[30][661],u_xpb_out[31][661],u_xpb_out[32][661],u_xpb_out[33][661],u_xpb_out[34][661],u_xpb_out[35][661],u_xpb_out[36][661],u_xpb_out[37][661],u_xpb_out[38][661],u_xpb_out[39][661],u_xpb_out[40][661],u_xpb_out[41][661],u_xpb_out[42][661],u_xpb_out[43][661],u_xpb_out[44][661],u_xpb_out[45][661],u_xpb_out[46][661],u_xpb_out[47][661],u_xpb_out[48][661],u_xpb_out[49][661],u_xpb_out[50][661],u_xpb_out[51][661],u_xpb_out[52][661],u_xpb_out[53][661],u_xpb_out[54][661],u_xpb_out[55][661],u_xpb_out[56][661],u_xpb_out[57][661],u_xpb_out[58][661],u_xpb_out[59][661],u_xpb_out[60][661],u_xpb_out[61][661],u_xpb_out[62][661],u_xpb_out[63][661],u_xpb_out[64][661],u_xpb_out[65][661],u_xpb_out[66][661],u_xpb_out[67][661],u_xpb_out[68][661],u_xpb_out[69][661],u_xpb_out[70][661],u_xpb_out[71][661],u_xpb_out[72][661],u_xpb_out[73][661],u_xpb_out[74][661],u_xpb_out[75][661],u_xpb_out[76][661],u_xpb_out[77][661],u_xpb_out[78][661],u_xpb_out[79][661],u_xpb_out[80][661],u_xpb_out[81][661],u_xpb_out[82][661],u_xpb_out[83][661],u_xpb_out[84][661],u_xpb_out[85][661],u_xpb_out[86][661],u_xpb_out[87][661],u_xpb_out[88][661],u_xpb_out[89][661],u_xpb_out[90][661],u_xpb_out[91][661],u_xpb_out[92][661],u_xpb_out[93][661],u_xpb_out[94][661],u_xpb_out[95][661],u_xpb_out[96][661],u_xpb_out[97][661],u_xpb_out[98][661],u_xpb_out[99][661],u_xpb_out[100][661],u_xpb_out[101][661],u_xpb_out[102][661],u_xpb_out[103][661],u_xpb_out[104][661],u_xpb_out[105][661]};

assign col_out_662 = {u_xpb_out[0][662],u_xpb_out[1][662],u_xpb_out[2][662],u_xpb_out[3][662],u_xpb_out[4][662],u_xpb_out[5][662],u_xpb_out[6][662],u_xpb_out[7][662],u_xpb_out[8][662],u_xpb_out[9][662],u_xpb_out[10][662],u_xpb_out[11][662],u_xpb_out[12][662],u_xpb_out[13][662],u_xpb_out[14][662],u_xpb_out[15][662],u_xpb_out[16][662],u_xpb_out[17][662],u_xpb_out[18][662],u_xpb_out[19][662],u_xpb_out[20][662],u_xpb_out[21][662],u_xpb_out[22][662],u_xpb_out[23][662],u_xpb_out[24][662],u_xpb_out[25][662],u_xpb_out[26][662],u_xpb_out[27][662],u_xpb_out[28][662],u_xpb_out[29][662],u_xpb_out[30][662],u_xpb_out[31][662],u_xpb_out[32][662],u_xpb_out[33][662],u_xpb_out[34][662],u_xpb_out[35][662],u_xpb_out[36][662],u_xpb_out[37][662],u_xpb_out[38][662],u_xpb_out[39][662],u_xpb_out[40][662],u_xpb_out[41][662],u_xpb_out[42][662],u_xpb_out[43][662],u_xpb_out[44][662],u_xpb_out[45][662],u_xpb_out[46][662],u_xpb_out[47][662],u_xpb_out[48][662],u_xpb_out[49][662],u_xpb_out[50][662],u_xpb_out[51][662],u_xpb_out[52][662],u_xpb_out[53][662],u_xpb_out[54][662],u_xpb_out[55][662],u_xpb_out[56][662],u_xpb_out[57][662],u_xpb_out[58][662],u_xpb_out[59][662],u_xpb_out[60][662],u_xpb_out[61][662],u_xpb_out[62][662],u_xpb_out[63][662],u_xpb_out[64][662],u_xpb_out[65][662],u_xpb_out[66][662],u_xpb_out[67][662],u_xpb_out[68][662],u_xpb_out[69][662],u_xpb_out[70][662],u_xpb_out[71][662],u_xpb_out[72][662],u_xpb_out[73][662],u_xpb_out[74][662],u_xpb_out[75][662],u_xpb_out[76][662],u_xpb_out[77][662],u_xpb_out[78][662],u_xpb_out[79][662],u_xpb_out[80][662],u_xpb_out[81][662],u_xpb_out[82][662],u_xpb_out[83][662],u_xpb_out[84][662],u_xpb_out[85][662],u_xpb_out[86][662],u_xpb_out[87][662],u_xpb_out[88][662],u_xpb_out[89][662],u_xpb_out[90][662],u_xpb_out[91][662],u_xpb_out[92][662],u_xpb_out[93][662],u_xpb_out[94][662],u_xpb_out[95][662],u_xpb_out[96][662],u_xpb_out[97][662],u_xpb_out[98][662],u_xpb_out[99][662],u_xpb_out[100][662],u_xpb_out[101][662],u_xpb_out[102][662],u_xpb_out[103][662],u_xpb_out[104][662],u_xpb_out[105][662]};

assign col_out_663 = {u_xpb_out[0][663],u_xpb_out[1][663],u_xpb_out[2][663],u_xpb_out[3][663],u_xpb_out[4][663],u_xpb_out[5][663],u_xpb_out[6][663],u_xpb_out[7][663],u_xpb_out[8][663],u_xpb_out[9][663],u_xpb_out[10][663],u_xpb_out[11][663],u_xpb_out[12][663],u_xpb_out[13][663],u_xpb_out[14][663],u_xpb_out[15][663],u_xpb_out[16][663],u_xpb_out[17][663],u_xpb_out[18][663],u_xpb_out[19][663],u_xpb_out[20][663],u_xpb_out[21][663],u_xpb_out[22][663],u_xpb_out[23][663],u_xpb_out[24][663],u_xpb_out[25][663],u_xpb_out[26][663],u_xpb_out[27][663],u_xpb_out[28][663],u_xpb_out[29][663],u_xpb_out[30][663],u_xpb_out[31][663],u_xpb_out[32][663],u_xpb_out[33][663],u_xpb_out[34][663],u_xpb_out[35][663],u_xpb_out[36][663],u_xpb_out[37][663],u_xpb_out[38][663],u_xpb_out[39][663],u_xpb_out[40][663],u_xpb_out[41][663],u_xpb_out[42][663],u_xpb_out[43][663],u_xpb_out[44][663],u_xpb_out[45][663],u_xpb_out[46][663],u_xpb_out[47][663],u_xpb_out[48][663],u_xpb_out[49][663],u_xpb_out[50][663],u_xpb_out[51][663],u_xpb_out[52][663],u_xpb_out[53][663],u_xpb_out[54][663],u_xpb_out[55][663],u_xpb_out[56][663],u_xpb_out[57][663],u_xpb_out[58][663],u_xpb_out[59][663],u_xpb_out[60][663],u_xpb_out[61][663],u_xpb_out[62][663],u_xpb_out[63][663],u_xpb_out[64][663],u_xpb_out[65][663],u_xpb_out[66][663],u_xpb_out[67][663],u_xpb_out[68][663],u_xpb_out[69][663],u_xpb_out[70][663],u_xpb_out[71][663],u_xpb_out[72][663],u_xpb_out[73][663],u_xpb_out[74][663],u_xpb_out[75][663],u_xpb_out[76][663],u_xpb_out[77][663],u_xpb_out[78][663],u_xpb_out[79][663],u_xpb_out[80][663],u_xpb_out[81][663],u_xpb_out[82][663],u_xpb_out[83][663],u_xpb_out[84][663],u_xpb_out[85][663],u_xpb_out[86][663],u_xpb_out[87][663],u_xpb_out[88][663],u_xpb_out[89][663],u_xpb_out[90][663],u_xpb_out[91][663],u_xpb_out[92][663],u_xpb_out[93][663],u_xpb_out[94][663],u_xpb_out[95][663],u_xpb_out[96][663],u_xpb_out[97][663],u_xpb_out[98][663],u_xpb_out[99][663],u_xpb_out[100][663],u_xpb_out[101][663],u_xpb_out[102][663],u_xpb_out[103][663],u_xpb_out[104][663],u_xpb_out[105][663]};

assign col_out_664 = {u_xpb_out[0][664],u_xpb_out[1][664],u_xpb_out[2][664],u_xpb_out[3][664],u_xpb_out[4][664],u_xpb_out[5][664],u_xpb_out[6][664],u_xpb_out[7][664],u_xpb_out[8][664],u_xpb_out[9][664],u_xpb_out[10][664],u_xpb_out[11][664],u_xpb_out[12][664],u_xpb_out[13][664],u_xpb_out[14][664],u_xpb_out[15][664],u_xpb_out[16][664],u_xpb_out[17][664],u_xpb_out[18][664],u_xpb_out[19][664],u_xpb_out[20][664],u_xpb_out[21][664],u_xpb_out[22][664],u_xpb_out[23][664],u_xpb_out[24][664],u_xpb_out[25][664],u_xpb_out[26][664],u_xpb_out[27][664],u_xpb_out[28][664],u_xpb_out[29][664],u_xpb_out[30][664],u_xpb_out[31][664],u_xpb_out[32][664],u_xpb_out[33][664],u_xpb_out[34][664],u_xpb_out[35][664],u_xpb_out[36][664],u_xpb_out[37][664],u_xpb_out[38][664],u_xpb_out[39][664],u_xpb_out[40][664],u_xpb_out[41][664],u_xpb_out[42][664],u_xpb_out[43][664],u_xpb_out[44][664],u_xpb_out[45][664],u_xpb_out[46][664],u_xpb_out[47][664],u_xpb_out[48][664],u_xpb_out[49][664],u_xpb_out[50][664],u_xpb_out[51][664],u_xpb_out[52][664],u_xpb_out[53][664],u_xpb_out[54][664],u_xpb_out[55][664],u_xpb_out[56][664],u_xpb_out[57][664],u_xpb_out[58][664],u_xpb_out[59][664],u_xpb_out[60][664],u_xpb_out[61][664],u_xpb_out[62][664],u_xpb_out[63][664],u_xpb_out[64][664],u_xpb_out[65][664],u_xpb_out[66][664],u_xpb_out[67][664],u_xpb_out[68][664],u_xpb_out[69][664],u_xpb_out[70][664],u_xpb_out[71][664],u_xpb_out[72][664],u_xpb_out[73][664],u_xpb_out[74][664],u_xpb_out[75][664],u_xpb_out[76][664],u_xpb_out[77][664],u_xpb_out[78][664],u_xpb_out[79][664],u_xpb_out[80][664],u_xpb_out[81][664],u_xpb_out[82][664],u_xpb_out[83][664],u_xpb_out[84][664],u_xpb_out[85][664],u_xpb_out[86][664],u_xpb_out[87][664],u_xpb_out[88][664],u_xpb_out[89][664],u_xpb_out[90][664],u_xpb_out[91][664],u_xpb_out[92][664],u_xpb_out[93][664],u_xpb_out[94][664],u_xpb_out[95][664],u_xpb_out[96][664],u_xpb_out[97][664],u_xpb_out[98][664],u_xpb_out[99][664],u_xpb_out[100][664],u_xpb_out[101][664],u_xpb_out[102][664],u_xpb_out[103][664],u_xpb_out[104][664],u_xpb_out[105][664]};

assign col_out_665 = {u_xpb_out[0][665],u_xpb_out[1][665],u_xpb_out[2][665],u_xpb_out[3][665],u_xpb_out[4][665],u_xpb_out[5][665],u_xpb_out[6][665],u_xpb_out[7][665],u_xpb_out[8][665],u_xpb_out[9][665],u_xpb_out[10][665],u_xpb_out[11][665],u_xpb_out[12][665],u_xpb_out[13][665],u_xpb_out[14][665],u_xpb_out[15][665],u_xpb_out[16][665],u_xpb_out[17][665],u_xpb_out[18][665],u_xpb_out[19][665],u_xpb_out[20][665],u_xpb_out[21][665],u_xpb_out[22][665],u_xpb_out[23][665],u_xpb_out[24][665],u_xpb_out[25][665],u_xpb_out[26][665],u_xpb_out[27][665],u_xpb_out[28][665],u_xpb_out[29][665],u_xpb_out[30][665],u_xpb_out[31][665],u_xpb_out[32][665],u_xpb_out[33][665],u_xpb_out[34][665],u_xpb_out[35][665],u_xpb_out[36][665],u_xpb_out[37][665],u_xpb_out[38][665],u_xpb_out[39][665],u_xpb_out[40][665],u_xpb_out[41][665],u_xpb_out[42][665],u_xpb_out[43][665],u_xpb_out[44][665],u_xpb_out[45][665],u_xpb_out[46][665],u_xpb_out[47][665],u_xpb_out[48][665],u_xpb_out[49][665],u_xpb_out[50][665],u_xpb_out[51][665],u_xpb_out[52][665],u_xpb_out[53][665],u_xpb_out[54][665],u_xpb_out[55][665],u_xpb_out[56][665],u_xpb_out[57][665],u_xpb_out[58][665],u_xpb_out[59][665],u_xpb_out[60][665],u_xpb_out[61][665],u_xpb_out[62][665],u_xpb_out[63][665],u_xpb_out[64][665],u_xpb_out[65][665],u_xpb_out[66][665],u_xpb_out[67][665],u_xpb_out[68][665],u_xpb_out[69][665],u_xpb_out[70][665],u_xpb_out[71][665],u_xpb_out[72][665],u_xpb_out[73][665],u_xpb_out[74][665],u_xpb_out[75][665],u_xpb_out[76][665],u_xpb_out[77][665],u_xpb_out[78][665],u_xpb_out[79][665],u_xpb_out[80][665],u_xpb_out[81][665],u_xpb_out[82][665],u_xpb_out[83][665],u_xpb_out[84][665],u_xpb_out[85][665],u_xpb_out[86][665],u_xpb_out[87][665],u_xpb_out[88][665],u_xpb_out[89][665],u_xpb_out[90][665],u_xpb_out[91][665],u_xpb_out[92][665],u_xpb_out[93][665],u_xpb_out[94][665],u_xpb_out[95][665],u_xpb_out[96][665],u_xpb_out[97][665],u_xpb_out[98][665],u_xpb_out[99][665],u_xpb_out[100][665],u_xpb_out[101][665],u_xpb_out[102][665],u_xpb_out[103][665],u_xpb_out[104][665],u_xpb_out[105][665]};

assign col_out_666 = {u_xpb_out[0][666],u_xpb_out[1][666],u_xpb_out[2][666],u_xpb_out[3][666],u_xpb_out[4][666],u_xpb_out[5][666],u_xpb_out[6][666],u_xpb_out[7][666],u_xpb_out[8][666],u_xpb_out[9][666],u_xpb_out[10][666],u_xpb_out[11][666],u_xpb_out[12][666],u_xpb_out[13][666],u_xpb_out[14][666],u_xpb_out[15][666],u_xpb_out[16][666],u_xpb_out[17][666],u_xpb_out[18][666],u_xpb_out[19][666],u_xpb_out[20][666],u_xpb_out[21][666],u_xpb_out[22][666],u_xpb_out[23][666],u_xpb_out[24][666],u_xpb_out[25][666],u_xpb_out[26][666],u_xpb_out[27][666],u_xpb_out[28][666],u_xpb_out[29][666],u_xpb_out[30][666],u_xpb_out[31][666],u_xpb_out[32][666],u_xpb_out[33][666],u_xpb_out[34][666],u_xpb_out[35][666],u_xpb_out[36][666],u_xpb_out[37][666],u_xpb_out[38][666],u_xpb_out[39][666],u_xpb_out[40][666],u_xpb_out[41][666],u_xpb_out[42][666],u_xpb_out[43][666],u_xpb_out[44][666],u_xpb_out[45][666],u_xpb_out[46][666],u_xpb_out[47][666],u_xpb_out[48][666],u_xpb_out[49][666],u_xpb_out[50][666],u_xpb_out[51][666],u_xpb_out[52][666],u_xpb_out[53][666],u_xpb_out[54][666],u_xpb_out[55][666],u_xpb_out[56][666],u_xpb_out[57][666],u_xpb_out[58][666],u_xpb_out[59][666],u_xpb_out[60][666],u_xpb_out[61][666],u_xpb_out[62][666],u_xpb_out[63][666],u_xpb_out[64][666],u_xpb_out[65][666],u_xpb_out[66][666],u_xpb_out[67][666],u_xpb_out[68][666],u_xpb_out[69][666],u_xpb_out[70][666],u_xpb_out[71][666],u_xpb_out[72][666],u_xpb_out[73][666],u_xpb_out[74][666],u_xpb_out[75][666],u_xpb_out[76][666],u_xpb_out[77][666],u_xpb_out[78][666],u_xpb_out[79][666],u_xpb_out[80][666],u_xpb_out[81][666],u_xpb_out[82][666],u_xpb_out[83][666],u_xpb_out[84][666],u_xpb_out[85][666],u_xpb_out[86][666],u_xpb_out[87][666],u_xpb_out[88][666],u_xpb_out[89][666],u_xpb_out[90][666],u_xpb_out[91][666],u_xpb_out[92][666],u_xpb_out[93][666],u_xpb_out[94][666],u_xpb_out[95][666],u_xpb_out[96][666],u_xpb_out[97][666],u_xpb_out[98][666],u_xpb_out[99][666],u_xpb_out[100][666],u_xpb_out[101][666],u_xpb_out[102][666],u_xpb_out[103][666],u_xpb_out[104][666],u_xpb_out[105][666]};

assign col_out_667 = {u_xpb_out[0][667],u_xpb_out[1][667],u_xpb_out[2][667],u_xpb_out[3][667],u_xpb_out[4][667],u_xpb_out[5][667],u_xpb_out[6][667],u_xpb_out[7][667],u_xpb_out[8][667],u_xpb_out[9][667],u_xpb_out[10][667],u_xpb_out[11][667],u_xpb_out[12][667],u_xpb_out[13][667],u_xpb_out[14][667],u_xpb_out[15][667],u_xpb_out[16][667],u_xpb_out[17][667],u_xpb_out[18][667],u_xpb_out[19][667],u_xpb_out[20][667],u_xpb_out[21][667],u_xpb_out[22][667],u_xpb_out[23][667],u_xpb_out[24][667],u_xpb_out[25][667],u_xpb_out[26][667],u_xpb_out[27][667],u_xpb_out[28][667],u_xpb_out[29][667],u_xpb_out[30][667],u_xpb_out[31][667],u_xpb_out[32][667],u_xpb_out[33][667],u_xpb_out[34][667],u_xpb_out[35][667],u_xpb_out[36][667],u_xpb_out[37][667],u_xpb_out[38][667],u_xpb_out[39][667],u_xpb_out[40][667],u_xpb_out[41][667],u_xpb_out[42][667],u_xpb_out[43][667],u_xpb_out[44][667],u_xpb_out[45][667],u_xpb_out[46][667],u_xpb_out[47][667],u_xpb_out[48][667],u_xpb_out[49][667],u_xpb_out[50][667],u_xpb_out[51][667],u_xpb_out[52][667],u_xpb_out[53][667],u_xpb_out[54][667],u_xpb_out[55][667],u_xpb_out[56][667],u_xpb_out[57][667],u_xpb_out[58][667],u_xpb_out[59][667],u_xpb_out[60][667],u_xpb_out[61][667],u_xpb_out[62][667],u_xpb_out[63][667],u_xpb_out[64][667],u_xpb_out[65][667],u_xpb_out[66][667],u_xpb_out[67][667],u_xpb_out[68][667],u_xpb_out[69][667],u_xpb_out[70][667],u_xpb_out[71][667],u_xpb_out[72][667],u_xpb_out[73][667],u_xpb_out[74][667],u_xpb_out[75][667],u_xpb_out[76][667],u_xpb_out[77][667],u_xpb_out[78][667],u_xpb_out[79][667],u_xpb_out[80][667],u_xpb_out[81][667],u_xpb_out[82][667],u_xpb_out[83][667],u_xpb_out[84][667],u_xpb_out[85][667],u_xpb_out[86][667],u_xpb_out[87][667],u_xpb_out[88][667],u_xpb_out[89][667],u_xpb_out[90][667],u_xpb_out[91][667],u_xpb_out[92][667],u_xpb_out[93][667],u_xpb_out[94][667],u_xpb_out[95][667],u_xpb_out[96][667],u_xpb_out[97][667],u_xpb_out[98][667],u_xpb_out[99][667],u_xpb_out[100][667],u_xpb_out[101][667],u_xpb_out[102][667],u_xpb_out[103][667],u_xpb_out[104][667],u_xpb_out[105][667]};

assign col_out_668 = {u_xpb_out[0][668],u_xpb_out[1][668],u_xpb_out[2][668],u_xpb_out[3][668],u_xpb_out[4][668],u_xpb_out[5][668],u_xpb_out[6][668],u_xpb_out[7][668],u_xpb_out[8][668],u_xpb_out[9][668],u_xpb_out[10][668],u_xpb_out[11][668],u_xpb_out[12][668],u_xpb_out[13][668],u_xpb_out[14][668],u_xpb_out[15][668],u_xpb_out[16][668],u_xpb_out[17][668],u_xpb_out[18][668],u_xpb_out[19][668],u_xpb_out[20][668],u_xpb_out[21][668],u_xpb_out[22][668],u_xpb_out[23][668],u_xpb_out[24][668],u_xpb_out[25][668],u_xpb_out[26][668],u_xpb_out[27][668],u_xpb_out[28][668],u_xpb_out[29][668],u_xpb_out[30][668],u_xpb_out[31][668],u_xpb_out[32][668],u_xpb_out[33][668],u_xpb_out[34][668],u_xpb_out[35][668],u_xpb_out[36][668],u_xpb_out[37][668],u_xpb_out[38][668],u_xpb_out[39][668],u_xpb_out[40][668],u_xpb_out[41][668],u_xpb_out[42][668],u_xpb_out[43][668],u_xpb_out[44][668],u_xpb_out[45][668],u_xpb_out[46][668],u_xpb_out[47][668],u_xpb_out[48][668],u_xpb_out[49][668],u_xpb_out[50][668],u_xpb_out[51][668],u_xpb_out[52][668],u_xpb_out[53][668],u_xpb_out[54][668],u_xpb_out[55][668],u_xpb_out[56][668],u_xpb_out[57][668],u_xpb_out[58][668],u_xpb_out[59][668],u_xpb_out[60][668],u_xpb_out[61][668],u_xpb_out[62][668],u_xpb_out[63][668],u_xpb_out[64][668],u_xpb_out[65][668],u_xpb_out[66][668],u_xpb_out[67][668],u_xpb_out[68][668],u_xpb_out[69][668],u_xpb_out[70][668],u_xpb_out[71][668],u_xpb_out[72][668],u_xpb_out[73][668],u_xpb_out[74][668],u_xpb_out[75][668],u_xpb_out[76][668],u_xpb_out[77][668],u_xpb_out[78][668],u_xpb_out[79][668],u_xpb_out[80][668],u_xpb_out[81][668],u_xpb_out[82][668],u_xpb_out[83][668],u_xpb_out[84][668],u_xpb_out[85][668],u_xpb_out[86][668],u_xpb_out[87][668],u_xpb_out[88][668],u_xpb_out[89][668],u_xpb_out[90][668],u_xpb_out[91][668],u_xpb_out[92][668],u_xpb_out[93][668],u_xpb_out[94][668],u_xpb_out[95][668],u_xpb_out[96][668],u_xpb_out[97][668],u_xpb_out[98][668],u_xpb_out[99][668],u_xpb_out[100][668],u_xpb_out[101][668],u_xpb_out[102][668],u_xpb_out[103][668],u_xpb_out[104][668],u_xpb_out[105][668]};

assign col_out_669 = {u_xpb_out[0][669],u_xpb_out[1][669],u_xpb_out[2][669],u_xpb_out[3][669],u_xpb_out[4][669],u_xpb_out[5][669],u_xpb_out[6][669],u_xpb_out[7][669],u_xpb_out[8][669],u_xpb_out[9][669],u_xpb_out[10][669],u_xpb_out[11][669],u_xpb_out[12][669],u_xpb_out[13][669],u_xpb_out[14][669],u_xpb_out[15][669],u_xpb_out[16][669],u_xpb_out[17][669],u_xpb_out[18][669],u_xpb_out[19][669],u_xpb_out[20][669],u_xpb_out[21][669],u_xpb_out[22][669],u_xpb_out[23][669],u_xpb_out[24][669],u_xpb_out[25][669],u_xpb_out[26][669],u_xpb_out[27][669],u_xpb_out[28][669],u_xpb_out[29][669],u_xpb_out[30][669],u_xpb_out[31][669],u_xpb_out[32][669],u_xpb_out[33][669],u_xpb_out[34][669],u_xpb_out[35][669],u_xpb_out[36][669],u_xpb_out[37][669],u_xpb_out[38][669],u_xpb_out[39][669],u_xpb_out[40][669],u_xpb_out[41][669],u_xpb_out[42][669],u_xpb_out[43][669],u_xpb_out[44][669],u_xpb_out[45][669],u_xpb_out[46][669],u_xpb_out[47][669],u_xpb_out[48][669],u_xpb_out[49][669],u_xpb_out[50][669],u_xpb_out[51][669],u_xpb_out[52][669],u_xpb_out[53][669],u_xpb_out[54][669],u_xpb_out[55][669],u_xpb_out[56][669],u_xpb_out[57][669],u_xpb_out[58][669],u_xpb_out[59][669],u_xpb_out[60][669],u_xpb_out[61][669],u_xpb_out[62][669],u_xpb_out[63][669],u_xpb_out[64][669],u_xpb_out[65][669],u_xpb_out[66][669],u_xpb_out[67][669],u_xpb_out[68][669],u_xpb_out[69][669],u_xpb_out[70][669],u_xpb_out[71][669],u_xpb_out[72][669],u_xpb_out[73][669],u_xpb_out[74][669],u_xpb_out[75][669],u_xpb_out[76][669],u_xpb_out[77][669],u_xpb_out[78][669],u_xpb_out[79][669],u_xpb_out[80][669],u_xpb_out[81][669],u_xpb_out[82][669],u_xpb_out[83][669],u_xpb_out[84][669],u_xpb_out[85][669],u_xpb_out[86][669],u_xpb_out[87][669],u_xpb_out[88][669],u_xpb_out[89][669],u_xpb_out[90][669],u_xpb_out[91][669],u_xpb_out[92][669],u_xpb_out[93][669],u_xpb_out[94][669],u_xpb_out[95][669],u_xpb_out[96][669],u_xpb_out[97][669],u_xpb_out[98][669],u_xpb_out[99][669],u_xpb_out[100][669],u_xpb_out[101][669],u_xpb_out[102][669],u_xpb_out[103][669],u_xpb_out[104][669],u_xpb_out[105][669]};

assign col_out_670 = {u_xpb_out[0][670],u_xpb_out[1][670],u_xpb_out[2][670],u_xpb_out[3][670],u_xpb_out[4][670],u_xpb_out[5][670],u_xpb_out[6][670],u_xpb_out[7][670],u_xpb_out[8][670],u_xpb_out[9][670],u_xpb_out[10][670],u_xpb_out[11][670],u_xpb_out[12][670],u_xpb_out[13][670],u_xpb_out[14][670],u_xpb_out[15][670],u_xpb_out[16][670],u_xpb_out[17][670],u_xpb_out[18][670],u_xpb_out[19][670],u_xpb_out[20][670],u_xpb_out[21][670],u_xpb_out[22][670],u_xpb_out[23][670],u_xpb_out[24][670],u_xpb_out[25][670],u_xpb_out[26][670],u_xpb_out[27][670],u_xpb_out[28][670],u_xpb_out[29][670],u_xpb_out[30][670],u_xpb_out[31][670],u_xpb_out[32][670],u_xpb_out[33][670],u_xpb_out[34][670],u_xpb_out[35][670],u_xpb_out[36][670],u_xpb_out[37][670],u_xpb_out[38][670],u_xpb_out[39][670],u_xpb_out[40][670],u_xpb_out[41][670],u_xpb_out[42][670],u_xpb_out[43][670],u_xpb_out[44][670],u_xpb_out[45][670],u_xpb_out[46][670],u_xpb_out[47][670],u_xpb_out[48][670],u_xpb_out[49][670],u_xpb_out[50][670],u_xpb_out[51][670],u_xpb_out[52][670],u_xpb_out[53][670],u_xpb_out[54][670],u_xpb_out[55][670],u_xpb_out[56][670],u_xpb_out[57][670],u_xpb_out[58][670],u_xpb_out[59][670],u_xpb_out[60][670],u_xpb_out[61][670],u_xpb_out[62][670],u_xpb_out[63][670],u_xpb_out[64][670],u_xpb_out[65][670],u_xpb_out[66][670],u_xpb_out[67][670],u_xpb_out[68][670],u_xpb_out[69][670],u_xpb_out[70][670],u_xpb_out[71][670],u_xpb_out[72][670],u_xpb_out[73][670],u_xpb_out[74][670],u_xpb_out[75][670],u_xpb_out[76][670],u_xpb_out[77][670],u_xpb_out[78][670],u_xpb_out[79][670],u_xpb_out[80][670],u_xpb_out[81][670],u_xpb_out[82][670],u_xpb_out[83][670],u_xpb_out[84][670],u_xpb_out[85][670],u_xpb_out[86][670],u_xpb_out[87][670],u_xpb_out[88][670],u_xpb_out[89][670],u_xpb_out[90][670],u_xpb_out[91][670],u_xpb_out[92][670],u_xpb_out[93][670],u_xpb_out[94][670],u_xpb_out[95][670],u_xpb_out[96][670],u_xpb_out[97][670],u_xpb_out[98][670],u_xpb_out[99][670],u_xpb_out[100][670],u_xpb_out[101][670],u_xpb_out[102][670],u_xpb_out[103][670],u_xpb_out[104][670],u_xpb_out[105][670]};

assign col_out_671 = {u_xpb_out[0][671],u_xpb_out[1][671],u_xpb_out[2][671],u_xpb_out[3][671],u_xpb_out[4][671],u_xpb_out[5][671],u_xpb_out[6][671],u_xpb_out[7][671],u_xpb_out[8][671],u_xpb_out[9][671],u_xpb_out[10][671],u_xpb_out[11][671],u_xpb_out[12][671],u_xpb_out[13][671],u_xpb_out[14][671],u_xpb_out[15][671],u_xpb_out[16][671],u_xpb_out[17][671],u_xpb_out[18][671],u_xpb_out[19][671],u_xpb_out[20][671],u_xpb_out[21][671],u_xpb_out[22][671],u_xpb_out[23][671],u_xpb_out[24][671],u_xpb_out[25][671],u_xpb_out[26][671],u_xpb_out[27][671],u_xpb_out[28][671],u_xpb_out[29][671],u_xpb_out[30][671],u_xpb_out[31][671],u_xpb_out[32][671],u_xpb_out[33][671],u_xpb_out[34][671],u_xpb_out[35][671],u_xpb_out[36][671],u_xpb_out[37][671],u_xpb_out[38][671],u_xpb_out[39][671],u_xpb_out[40][671],u_xpb_out[41][671],u_xpb_out[42][671],u_xpb_out[43][671],u_xpb_out[44][671],u_xpb_out[45][671],u_xpb_out[46][671],u_xpb_out[47][671],u_xpb_out[48][671],u_xpb_out[49][671],u_xpb_out[50][671],u_xpb_out[51][671],u_xpb_out[52][671],u_xpb_out[53][671],u_xpb_out[54][671],u_xpb_out[55][671],u_xpb_out[56][671],u_xpb_out[57][671],u_xpb_out[58][671],u_xpb_out[59][671],u_xpb_out[60][671],u_xpb_out[61][671],u_xpb_out[62][671],u_xpb_out[63][671],u_xpb_out[64][671],u_xpb_out[65][671],u_xpb_out[66][671],u_xpb_out[67][671],u_xpb_out[68][671],u_xpb_out[69][671],u_xpb_out[70][671],u_xpb_out[71][671],u_xpb_out[72][671],u_xpb_out[73][671],u_xpb_out[74][671],u_xpb_out[75][671],u_xpb_out[76][671],u_xpb_out[77][671],u_xpb_out[78][671],u_xpb_out[79][671],u_xpb_out[80][671],u_xpb_out[81][671],u_xpb_out[82][671],u_xpb_out[83][671],u_xpb_out[84][671],u_xpb_out[85][671],u_xpb_out[86][671],u_xpb_out[87][671],u_xpb_out[88][671],u_xpb_out[89][671],u_xpb_out[90][671],u_xpb_out[91][671],u_xpb_out[92][671],u_xpb_out[93][671],u_xpb_out[94][671],u_xpb_out[95][671],u_xpb_out[96][671],u_xpb_out[97][671],u_xpb_out[98][671],u_xpb_out[99][671],u_xpb_out[100][671],u_xpb_out[101][671],u_xpb_out[102][671],u_xpb_out[103][671],u_xpb_out[104][671],u_xpb_out[105][671]};

assign col_out_672 = {u_xpb_out[0][672],u_xpb_out[1][672],u_xpb_out[2][672],u_xpb_out[3][672],u_xpb_out[4][672],u_xpb_out[5][672],u_xpb_out[6][672],u_xpb_out[7][672],u_xpb_out[8][672],u_xpb_out[9][672],u_xpb_out[10][672],u_xpb_out[11][672],u_xpb_out[12][672],u_xpb_out[13][672],u_xpb_out[14][672],u_xpb_out[15][672],u_xpb_out[16][672],u_xpb_out[17][672],u_xpb_out[18][672],u_xpb_out[19][672],u_xpb_out[20][672],u_xpb_out[21][672],u_xpb_out[22][672],u_xpb_out[23][672],u_xpb_out[24][672],u_xpb_out[25][672],u_xpb_out[26][672],u_xpb_out[27][672],u_xpb_out[28][672],u_xpb_out[29][672],u_xpb_out[30][672],u_xpb_out[31][672],u_xpb_out[32][672],u_xpb_out[33][672],u_xpb_out[34][672],u_xpb_out[35][672],u_xpb_out[36][672],u_xpb_out[37][672],u_xpb_out[38][672],u_xpb_out[39][672],u_xpb_out[40][672],u_xpb_out[41][672],u_xpb_out[42][672],u_xpb_out[43][672],u_xpb_out[44][672],u_xpb_out[45][672],u_xpb_out[46][672],u_xpb_out[47][672],u_xpb_out[48][672],u_xpb_out[49][672],u_xpb_out[50][672],u_xpb_out[51][672],u_xpb_out[52][672],u_xpb_out[53][672],u_xpb_out[54][672],u_xpb_out[55][672],u_xpb_out[56][672],u_xpb_out[57][672],u_xpb_out[58][672],u_xpb_out[59][672],u_xpb_out[60][672],u_xpb_out[61][672],u_xpb_out[62][672],u_xpb_out[63][672],u_xpb_out[64][672],u_xpb_out[65][672],u_xpb_out[66][672],u_xpb_out[67][672],u_xpb_out[68][672],u_xpb_out[69][672],u_xpb_out[70][672],u_xpb_out[71][672],u_xpb_out[72][672],u_xpb_out[73][672],u_xpb_out[74][672],u_xpb_out[75][672],u_xpb_out[76][672],u_xpb_out[77][672],u_xpb_out[78][672],u_xpb_out[79][672],u_xpb_out[80][672],u_xpb_out[81][672],u_xpb_out[82][672],u_xpb_out[83][672],u_xpb_out[84][672],u_xpb_out[85][672],u_xpb_out[86][672],u_xpb_out[87][672],u_xpb_out[88][672],u_xpb_out[89][672],u_xpb_out[90][672],u_xpb_out[91][672],u_xpb_out[92][672],u_xpb_out[93][672],u_xpb_out[94][672],u_xpb_out[95][672],u_xpb_out[96][672],u_xpb_out[97][672],u_xpb_out[98][672],u_xpb_out[99][672],u_xpb_out[100][672],u_xpb_out[101][672],u_xpb_out[102][672],u_xpb_out[103][672],u_xpb_out[104][672],u_xpb_out[105][672]};

assign col_out_673 = {u_xpb_out[0][673],u_xpb_out[1][673],u_xpb_out[2][673],u_xpb_out[3][673],u_xpb_out[4][673],u_xpb_out[5][673],u_xpb_out[6][673],u_xpb_out[7][673],u_xpb_out[8][673],u_xpb_out[9][673],u_xpb_out[10][673],u_xpb_out[11][673],u_xpb_out[12][673],u_xpb_out[13][673],u_xpb_out[14][673],u_xpb_out[15][673],u_xpb_out[16][673],u_xpb_out[17][673],u_xpb_out[18][673],u_xpb_out[19][673],u_xpb_out[20][673],u_xpb_out[21][673],u_xpb_out[22][673],u_xpb_out[23][673],u_xpb_out[24][673],u_xpb_out[25][673],u_xpb_out[26][673],u_xpb_out[27][673],u_xpb_out[28][673],u_xpb_out[29][673],u_xpb_out[30][673],u_xpb_out[31][673],u_xpb_out[32][673],u_xpb_out[33][673],u_xpb_out[34][673],u_xpb_out[35][673],u_xpb_out[36][673],u_xpb_out[37][673],u_xpb_out[38][673],u_xpb_out[39][673],u_xpb_out[40][673],u_xpb_out[41][673],u_xpb_out[42][673],u_xpb_out[43][673],u_xpb_out[44][673],u_xpb_out[45][673],u_xpb_out[46][673],u_xpb_out[47][673],u_xpb_out[48][673],u_xpb_out[49][673],u_xpb_out[50][673],u_xpb_out[51][673],u_xpb_out[52][673],u_xpb_out[53][673],u_xpb_out[54][673],u_xpb_out[55][673],u_xpb_out[56][673],u_xpb_out[57][673],u_xpb_out[58][673],u_xpb_out[59][673],u_xpb_out[60][673],u_xpb_out[61][673],u_xpb_out[62][673],u_xpb_out[63][673],u_xpb_out[64][673],u_xpb_out[65][673],u_xpb_out[66][673],u_xpb_out[67][673],u_xpb_out[68][673],u_xpb_out[69][673],u_xpb_out[70][673],u_xpb_out[71][673],u_xpb_out[72][673],u_xpb_out[73][673],u_xpb_out[74][673],u_xpb_out[75][673],u_xpb_out[76][673],u_xpb_out[77][673],u_xpb_out[78][673],u_xpb_out[79][673],u_xpb_out[80][673],u_xpb_out[81][673],u_xpb_out[82][673],u_xpb_out[83][673],u_xpb_out[84][673],u_xpb_out[85][673],u_xpb_out[86][673],u_xpb_out[87][673],u_xpb_out[88][673],u_xpb_out[89][673],u_xpb_out[90][673],u_xpb_out[91][673],u_xpb_out[92][673],u_xpb_out[93][673],u_xpb_out[94][673],u_xpb_out[95][673],u_xpb_out[96][673],u_xpb_out[97][673],u_xpb_out[98][673],u_xpb_out[99][673],u_xpb_out[100][673],u_xpb_out[101][673],u_xpb_out[102][673],u_xpb_out[103][673],u_xpb_out[104][673],u_xpb_out[105][673]};

assign col_out_674 = {u_xpb_out[0][674],u_xpb_out[1][674],u_xpb_out[2][674],u_xpb_out[3][674],u_xpb_out[4][674],u_xpb_out[5][674],u_xpb_out[6][674],u_xpb_out[7][674],u_xpb_out[8][674],u_xpb_out[9][674],u_xpb_out[10][674],u_xpb_out[11][674],u_xpb_out[12][674],u_xpb_out[13][674],u_xpb_out[14][674],u_xpb_out[15][674],u_xpb_out[16][674],u_xpb_out[17][674],u_xpb_out[18][674],u_xpb_out[19][674],u_xpb_out[20][674],u_xpb_out[21][674],u_xpb_out[22][674],u_xpb_out[23][674],u_xpb_out[24][674],u_xpb_out[25][674],u_xpb_out[26][674],u_xpb_out[27][674],u_xpb_out[28][674],u_xpb_out[29][674],u_xpb_out[30][674],u_xpb_out[31][674],u_xpb_out[32][674],u_xpb_out[33][674],u_xpb_out[34][674],u_xpb_out[35][674],u_xpb_out[36][674],u_xpb_out[37][674],u_xpb_out[38][674],u_xpb_out[39][674],u_xpb_out[40][674],u_xpb_out[41][674],u_xpb_out[42][674],u_xpb_out[43][674],u_xpb_out[44][674],u_xpb_out[45][674],u_xpb_out[46][674],u_xpb_out[47][674],u_xpb_out[48][674],u_xpb_out[49][674],u_xpb_out[50][674],u_xpb_out[51][674],u_xpb_out[52][674],u_xpb_out[53][674],u_xpb_out[54][674],u_xpb_out[55][674],u_xpb_out[56][674],u_xpb_out[57][674],u_xpb_out[58][674],u_xpb_out[59][674],u_xpb_out[60][674],u_xpb_out[61][674],u_xpb_out[62][674],u_xpb_out[63][674],u_xpb_out[64][674],u_xpb_out[65][674],u_xpb_out[66][674],u_xpb_out[67][674],u_xpb_out[68][674],u_xpb_out[69][674],u_xpb_out[70][674],u_xpb_out[71][674],u_xpb_out[72][674],u_xpb_out[73][674],u_xpb_out[74][674],u_xpb_out[75][674],u_xpb_out[76][674],u_xpb_out[77][674],u_xpb_out[78][674],u_xpb_out[79][674],u_xpb_out[80][674],u_xpb_out[81][674],u_xpb_out[82][674],u_xpb_out[83][674],u_xpb_out[84][674],u_xpb_out[85][674],u_xpb_out[86][674],u_xpb_out[87][674],u_xpb_out[88][674],u_xpb_out[89][674],u_xpb_out[90][674],u_xpb_out[91][674],u_xpb_out[92][674],u_xpb_out[93][674],u_xpb_out[94][674],u_xpb_out[95][674],u_xpb_out[96][674],u_xpb_out[97][674],u_xpb_out[98][674],u_xpb_out[99][674],u_xpb_out[100][674],u_xpb_out[101][674],u_xpb_out[102][674],u_xpb_out[103][674],u_xpb_out[104][674],u_xpb_out[105][674]};

assign col_out_675 = {u_xpb_out[0][675],u_xpb_out[1][675],u_xpb_out[2][675],u_xpb_out[3][675],u_xpb_out[4][675],u_xpb_out[5][675],u_xpb_out[6][675],u_xpb_out[7][675],u_xpb_out[8][675],u_xpb_out[9][675],u_xpb_out[10][675],u_xpb_out[11][675],u_xpb_out[12][675],u_xpb_out[13][675],u_xpb_out[14][675],u_xpb_out[15][675],u_xpb_out[16][675],u_xpb_out[17][675],u_xpb_out[18][675],u_xpb_out[19][675],u_xpb_out[20][675],u_xpb_out[21][675],u_xpb_out[22][675],u_xpb_out[23][675],u_xpb_out[24][675],u_xpb_out[25][675],u_xpb_out[26][675],u_xpb_out[27][675],u_xpb_out[28][675],u_xpb_out[29][675],u_xpb_out[30][675],u_xpb_out[31][675],u_xpb_out[32][675],u_xpb_out[33][675],u_xpb_out[34][675],u_xpb_out[35][675],u_xpb_out[36][675],u_xpb_out[37][675],u_xpb_out[38][675],u_xpb_out[39][675],u_xpb_out[40][675],u_xpb_out[41][675],u_xpb_out[42][675],u_xpb_out[43][675],u_xpb_out[44][675],u_xpb_out[45][675],u_xpb_out[46][675],u_xpb_out[47][675],u_xpb_out[48][675],u_xpb_out[49][675],u_xpb_out[50][675],u_xpb_out[51][675],u_xpb_out[52][675],u_xpb_out[53][675],u_xpb_out[54][675],u_xpb_out[55][675],u_xpb_out[56][675],u_xpb_out[57][675],u_xpb_out[58][675],u_xpb_out[59][675],u_xpb_out[60][675],u_xpb_out[61][675],u_xpb_out[62][675],u_xpb_out[63][675],u_xpb_out[64][675],u_xpb_out[65][675],u_xpb_out[66][675],u_xpb_out[67][675],u_xpb_out[68][675],u_xpb_out[69][675],u_xpb_out[70][675],u_xpb_out[71][675],u_xpb_out[72][675],u_xpb_out[73][675],u_xpb_out[74][675],u_xpb_out[75][675],u_xpb_out[76][675],u_xpb_out[77][675],u_xpb_out[78][675],u_xpb_out[79][675],u_xpb_out[80][675],u_xpb_out[81][675],u_xpb_out[82][675],u_xpb_out[83][675],u_xpb_out[84][675],u_xpb_out[85][675],u_xpb_out[86][675],u_xpb_out[87][675],u_xpb_out[88][675],u_xpb_out[89][675],u_xpb_out[90][675],u_xpb_out[91][675],u_xpb_out[92][675],u_xpb_out[93][675],u_xpb_out[94][675],u_xpb_out[95][675],u_xpb_out[96][675],u_xpb_out[97][675],u_xpb_out[98][675],u_xpb_out[99][675],u_xpb_out[100][675],u_xpb_out[101][675],u_xpb_out[102][675],u_xpb_out[103][675],u_xpb_out[104][675],u_xpb_out[105][675]};

assign col_out_676 = {u_xpb_out[0][676],u_xpb_out[1][676],u_xpb_out[2][676],u_xpb_out[3][676],u_xpb_out[4][676],u_xpb_out[5][676],u_xpb_out[6][676],u_xpb_out[7][676],u_xpb_out[8][676],u_xpb_out[9][676],u_xpb_out[10][676],u_xpb_out[11][676],u_xpb_out[12][676],u_xpb_out[13][676],u_xpb_out[14][676],u_xpb_out[15][676],u_xpb_out[16][676],u_xpb_out[17][676],u_xpb_out[18][676],u_xpb_out[19][676],u_xpb_out[20][676],u_xpb_out[21][676],u_xpb_out[22][676],u_xpb_out[23][676],u_xpb_out[24][676],u_xpb_out[25][676],u_xpb_out[26][676],u_xpb_out[27][676],u_xpb_out[28][676],u_xpb_out[29][676],u_xpb_out[30][676],u_xpb_out[31][676],u_xpb_out[32][676],u_xpb_out[33][676],u_xpb_out[34][676],u_xpb_out[35][676],u_xpb_out[36][676],u_xpb_out[37][676],u_xpb_out[38][676],u_xpb_out[39][676],u_xpb_out[40][676],u_xpb_out[41][676],u_xpb_out[42][676],u_xpb_out[43][676],u_xpb_out[44][676],u_xpb_out[45][676],u_xpb_out[46][676],u_xpb_out[47][676],u_xpb_out[48][676],u_xpb_out[49][676],u_xpb_out[50][676],u_xpb_out[51][676],u_xpb_out[52][676],u_xpb_out[53][676],u_xpb_out[54][676],u_xpb_out[55][676],u_xpb_out[56][676],u_xpb_out[57][676],u_xpb_out[58][676],u_xpb_out[59][676],u_xpb_out[60][676],u_xpb_out[61][676],u_xpb_out[62][676],u_xpb_out[63][676],u_xpb_out[64][676],u_xpb_out[65][676],u_xpb_out[66][676],u_xpb_out[67][676],u_xpb_out[68][676],u_xpb_out[69][676],u_xpb_out[70][676],u_xpb_out[71][676],u_xpb_out[72][676],u_xpb_out[73][676],u_xpb_out[74][676],u_xpb_out[75][676],u_xpb_out[76][676],u_xpb_out[77][676],u_xpb_out[78][676],u_xpb_out[79][676],u_xpb_out[80][676],u_xpb_out[81][676],u_xpb_out[82][676],u_xpb_out[83][676],u_xpb_out[84][676],u_xpb_out[85][676],u_xpb_out[86][676],u_xpb_out[87][676],u_xpb_out[88][676],u_xpb_out[89][676],u_xpb_out[90][676],u_xpb_out[91][676],u_xpb_out[92][676],u_xpb_out[93][676],u_xpb_out[94][676],u_xpb_out[95][676],u_xpb_out[96][676],u_xpb_out[97][676],u_xpb_out[98][676],u_xpb_out[99][676],u_xpb_out[100][676],u_xpb_out[101][676],u_xpb_out[102][676],u_xpb_out[103][676],u_xpb_out[104][676],u_xpb_out[105][676]};

assign col_out_677 = {u_xpb_out[0][677],u_xpb_out[1][677],u_xpb_out[2][677],u_xpb_out[3][677],u_xpb_out[4][677],u_xpb_out[5][677],u_xpb_out[6][677],u_xpb_out[7][677],u_xpb_out[8][677],u_xpb_out[9][677],u_xpb_out[10][677],u_xpb_out[11][677],u_xpb_out[12][677],u_xpb_out[13][677],u_xpb_out[14][677],u_xpb_out[15][677],u_xpb_out[16][677],u_xpb_out[17][677],u_xpb_out[18][677],u_xpb_out[19][677],u_xpb_out[20][677],u_xpb_out[21][677],u_xpb_out[22][677],u_xpb_out[23][677],u_xpb_out[24][677],u_xpb_out[25][677],u_xpb_out[26][677],u_xpb_out[27][677],u_xpb_out[28][677],u_xpb_out[29][677],u_xpb_out[30][677],u_xpb_out[31][677],u_xpb_out[32][677],u_xpb_out[33][677],u_xpb_out[34][677],u_xpb_out[35][677],u_xpb_out[36][677],u_xpb_out[37][677],u_xpb_out[38][677],u_xpb_out[39][677],u_xpb_out[40][677],u_xpb_out[41][677],u_xpb_out[42][677],u_xpb_out[43][677],u_xpb_out[44][677],u_xpb_out[45][677],u_xpb_out[46][677],u_xpb_out[47][677],u_xpb_out[48][677],u_xpb_out[49][677],u_xpb_out[50][677],u_xpb_out[51][677],u_xpb_out[52][677],u_xpb_out[53][677],u_xpb_out[54][677],u_xpb_out[55][677],u_xpb_out[56][677],u_xpb_out[57][677],u_xpb_out[58][677],u_xpb_out[59][677],u_xpb_out[60][677],u_xpb_out[61][677],u_xpb_out[62][677],u_xpb_out[63][677],u_xpb_out[64][677],u_xpb_out[65][677],u_xpb_out[66][677],u_xpb_out[67][677],u_xpb_out[68][677],u_xpb_out[69][677],u_xpb_out[70][677],u_xpb_out[71][677],u_xpb_out[72][677],u_xpb_out[73][677],u_xpb_out[74][677],u_xpb_out[75][677],u_xpb_out[76][677],u_xpb_out[77][677],u_xpb_out[78][677],u_xpb_out[79][677],u_xpb_out[80][677],u_xpb_out[81][677],u_xpb_out[82][677],u_xpb_out[83][677],u_xpb_out[84][677],u_xpb_out[85][677],u_xpb_out[86][677],u_xpb_out[87][677],u_xpb_out[88][677],u_xpb_out[89][677],u_xpb_out[90][677],u_xpb_out[91][677],u_xpb_out[92][677],u_xpb_out[93][677],u_xpb_out[94][677],u_xpb_out[95][677],u_xpb_out[96][677],u_xpb_out[97][677],u_xpb_out[98][677],u_xpb_out[99][677],u_xpb_out[100][677],u_xpb_out[101][677],u_xpb_out[102][677],u_xpb_out[103][677],u_xpb_out[104][677],u_xpb_out[105][677]};

assign col_out_678 = {u_xpb_out[0][678],u_xpb_out[1][678],u_xpb_out[2][678],u_xpb_out[3][678],u_xpb_out[4][678],u_xpb_out[5][678],u_xpb_out[6][678],u_xpb_out[7][678],u_xpb_out[8][678],u_xpb_out[9][678],u_xpb_out[10][678],u_xpb_out[11][678],u_xpb_out[12][678],u_xpb_out[13][678],u_xpb_out[14][678],u_xpb_out[15][678],u_xpb_out[16][678],u_xpb_out[17][678],u_xpb_out[18][678],u_xpb_out[19][678],u_xpb_out[20][678],u_xpb_out[21][678],u_xpb_out[22][678],u_xpb_out[23][678],u_xpb_out[24][678],u_xpb_out[25][678],u_xpb_out[26][678],u_xpb_out[27][678],u_xpb_out[28][678],u_xpb_out[29][678],u_xpb_out[30][678],u_xpb_out[31][678],u_xpb_out[32][678],u_xpb_out[33][678],u_xpb_out[34][678],u_xpb_out[35][678],u_xpb_out[36][678],u_xpb_out[37][678],u_xpb_out[38][678],u_xpb_out[39][678],u_xpb_out[40][678],u_xpb_out[41][678],u_xpb_out[42][678],u_xpb_out[43][678],u_xpb_out[44][678],u_xpb_out[45][678],u_xpb_out[46][678],u_xpb_out[47][678],u_xpb_out[48][678],u_xpb_out[49][678],u_xpb_out[50][678],u_xpb_out[51][678],u_xpb_out[52][678],u_xpb_out[53][678],u_xpb_out[54][678],u_xpb_out[55][678],u_xpb_out[56][678],u_xpb_out[57][678],u_xpb_out[58][678],u_xpb_out[59][678],u_xpb_out[60][678],u_xpb_out[61][678],u_xpb_out[62][678],u_xpb_out[63][678],u_xpb_out[64][678],u_xpb_out[65][678],u_xpb_out[66][678],u_xpb_out[67][678],u_xpb_out[68][678],u_xpb_out[69][678],u_xpb_out[70][678],u_xpb_out[71][678],u_xpb_out[72][678],u_xpb_out[73][678],u_xpb_out[74][678],u_xpb_out[75][678],u_xpb_out[76][678],u_xpb_out[77][678],u_xpb_out[78][678],u_xpb_out[79][678],u_xpb_out[80][678],u_xpb_out[81][678],u_xpb_out[82][678],u_xpb_out[83][678],u_xpb_out[84][678],u_xpb_out[85][678],u_xpb_out[86][678],u_xpb_out[87][678],u_xpb_out[88][678],u_xpb_out[89][678],u_xpb_out[90][678],u_xpb_out[91][678],u_xpb_out[92][678],u_xpb_out[93][678],u_xpb_out[94][678],u_xpb_out[95][678],u_xpb_out[96][678],u_xpb_out[97][678],u_xpb_out[98][678],u_xpb_out[99][678],u_xpb_out[100][678],u_xpb_out[101][678],u_xpb_out[102][678],u_xpb_out[103][678],u_xpb_out[104][678],u_xpb_out[105][678]};

assign col_out_679 = {u_xpb_out[0][679],u_xpb_out[1][679],u_xpb_out[2][679],u_xpb_out[3][679],u_xpb_out[4][679],u_xpb_out[5][679],u_xpb_out[6][679],u_xpb_out[7][679],u_xpb_out[8][679],u_xpb_out[9][679],u_xpb_out[10][679],u_xpb_out[11][679],u_xpb_out[12][679],u_xpb_out[13][679],u_xpb_out[14][679],u_xpb_out[15][679],u_xpb_out[16][679],u_xpb_out[17][679],u_xpb_out[18][679],u_xpb_out[19][679],u_xpb_out[20][679],u_xpb_out[21][679],u_xpb_out[22][679],u_xpb_out[23][679],u_xpb_out[24][679],u_xpb_out[25][679],u_xpb_out[26][679],u_xpb_out[27][679],u_xpb_out[28][679],u_xpb_out[29][679],u_xpb_out[30][679],u_xpb_out[31][679],u_xpb_out[32][679],u_xpb_out[33][679],u_xpb_out[34][679],u_xpb_out[35][679],u_xpb_out[36][679],u_xpb_out[37][679],u_xpb_out[38][679],u_xpb_out[39][679],u_xpb_out[40][679],u_xpb_out[41][679],u_xpb_out[42][679],u_xpb_out[43][679],u_xpb_out[44][679],u_xpb_out[45][679],u_xpb_out[46][679],u_xpb_out[47][679],u_xpb_out[48][679],u_xpb_out[49][679],u_xpb_out[50][679],u_xpb_out[51][679],u_xpb_out[52][679],u_xpb_out[53][679],u_xpb_out[54][679],u_xpb_out[55][679],u_xpb_out[56][679],u_xpb_out[57][679],u_xpb_out[58][679],u_xpb_out[59][679],u_xpb_out[60][679],u_xpb_out[61][679],u_xpb_out[62][679],u_xpb_out[63][679],u_xpb_out[64][679],u_xpb_out[65][679],u_xpb_out[66][679],u_xpb_out[67][679],u_xpb_out[68][679],u_xpb_out[69][679],u_xpb_out[70][679],u_xpb_out[71][679],u_xpb_out[72][679],u_xpb_out[73][679],u_xpb_out[74][679],u_xpb_out[75][679],u_xpb_out[76][679],u_xpb_out[77][679],u_xpb_out[78][679],u_xpb_out[79][679],u_xpb_out[80][679],u_xpb_out[81][679],u_xpb_out[82][679],u_xpb_out[83][679],u_xpb_out[84][679],u_xpb_out[85][679],u_xpb_out[86][679],u_xpb_out[87][679],u_xpb_out[88][679],u_xpb_out[89][679],u_xpb_out[90][679],u_xpb_out[91][679],u_xpb_out[92][679],u_xpb_out[93][679],u_xpb_out[94][679],u_xpb_out[95][679],u_xpb_out[96][679],u_xpb_out[97][679],u_xpb_out[98][679],u_xpb_out[99][679],u_xpb_out[100][679],u_xpb_out[101][679],u_xpb_out[102][679],u_xpb_out[103][679],u_xpb_out[104][679],u_xpb_out[105][679]};

assign col_out_680 = {u_xpb_out[0][680],u_xpb_out[1][680],u_xpb_out[2][680],u_xpb_out[3][680],u_xpb_out[4][680],u_xpb_out[5][680],u_xpb_out[6][680],u_xpb_out[7][680],u_xpb_out[8][680],u_xpb_out[9][680],u_xpb_out[10][680],u_xpb_out[11][680],u_xpb_out[12][680],u_xpb_out[13][680],u_xpb_out[14][680],u_xpb_out[15][680],u_xpb_out[16][680],u_xpb_out[17][680],u_xpb_out[18][680],u_xpb_out[19][680],u_xpb_out[20][680],u_xpb_out[21][680],u_xpb_out[22][680],u_xpb_out[23][680],u_xpb_out[24][680],u_xpb_out[25][680],u_xpb_out[26][680],u_xpb_out[27][680],u_xpb_out[28][680],u_xpb_out[29][680],u_xpb_out[30][680],u_xpb_out[31][680],u_xpb_out[32][680],u_xpb_out[33][680],u_xpb_out[34][680],u_xpb_out[35][680],u_xpb_out[36][680],u_xpb_out[37][680],u_xpb_out[38][680],u_xpb_out[39][680],u_xpb_out[40][680],u_xpb_out[41][680],u_xpb_out[42][680],u_xpb_out[43][680],u_xpb_out[44][680],u_xpb_out[45][680],u_xpb_out[46][680],u_xpb_out[47][680],u_xpb_out[48][680],u_xpb_out[49][680],u_xpb_out[50][680],u_xpb_out[51][680],u_xpb_out[52][680],u_xpb_out[53][680],u_xpb_out[54][680],u_xpb_out[55][680],u_xpb_out[56][680],u_xpb_out[57][680],u_xpb_out[58][680],u_xpb_out[59][680],u_xpb_out[60][680],u_xpb_out[61][680],u_xpb_out[62][680],u_xpb_out[63][680],u_xpb_out[64][680],u_xpb_out[65][680],u_xpb_out[66][680],u_xpb_out[67][680],u_xpb_out[68][680],u_xpb_out[69][680],u_xpb_out[70][680],u_xpb_out[71][680],u_xpb_out[72][680],u_xpb_out[73][680],u_xpb_out[74][680],u_xpb_out[75][680],u_xpb_out[76][680],u_xpb_out[77][680],u_xpb_out[78][680],u_xpb_out[79][680],u_xpb_out[80][680],u_xpb_out[81][680],u_xpb_out[82][680],u_xpb_out[83][680],u_xpb_out[84][680],u_xpb_out[85][680],u_xpb_out[86][680],u_xpb_out[87][680],u_xpb_out[88][680],u_xpb_out[89][680],u_xpb_out[90][680],u_xpb_out[91][680],u_xpb_out[92][680],u_xpb_out[93][680],u_xpb_out[94][680],u_xpb_out[95][680],u_xpb_out[96][680],u_xpb_out[97][680],u_xpb_out[98][680],u_xpb_out[99][680],u_xpb_out[100][680],u_xpb_out[101][680],u_xpb_out[102][680],u_xpb_out[103][680],u_xpb_out[104][680],u_xpb_out[105][680]};

assign col_out_681 = {u_xpb_out[0][681],u_xpb_out[1][681],u_xpb_out[2][681],u_xpb_out[3][681],u_xpb_out[4][681],u_xpb_out[5][681],u_xpb_out[6][681],u_xpb_out[7][681],u_xpb_out[8][681],u_xpb_out[9][681],u_xpb_out[10][681],u_xpb_out[11][681],u_xpb_out[12][681],u_xpb_out[13][681],u_xpb_out[14][681],u_xpb_out[15][681],u_xpb_out[16][681],u_xpb_out[17][681],u_xpb_out[18][681],u_xpb_out[19][681],u_xpb_out[20][681],u_xpb_out[21][681],u_xpb_out[22][681],u_xpb_out[23][681],u_xpb_out[24][681],u_xpb_out[25][681],u_xpb_out[26][681],u_xpb_out[27][681],u_xpb_out[28][681],u_xpb_out[29][681],u_xpb_out[30][681],u_xpb_out[31][681],u_xpb_out[32][681],u_xpb_out[33][681],u_xpb_out[34][681],u_xpb_out[35][681],u_xpb_out[36][681],u_xpb_out[37][681],u_xpb_out[38][681],u_xpb_out[39][681],u_xpb_out[40][681],u_xpb_out[41][681],u_xpb_out[42][681],u_xpb_out[43][681],u_xpb_out[44][681],u_xpb_out[45][681],u_xpb_out[46][681],u_xpb_out[47][681],u_xpb_out[48][681],u_xpb_out[49][681],u_xpb_out[50][681],u_xpb_out[51][681],u_xpb_out[52][681],u_xpb_out[53][681],u_xpb_out[54][681],u_xpb_out[55][681],u_xpb_out[56][681],u_xpb_out[57][681],u_xpb_out[58][681],u_xpb_out[59][681],u_xpb_out[60][681],u_xpb_out[61][681],u_xpb_out[62][681],u_xpb_out[63][681],u_xpb_out[64][681],u_xpb_out[65][681],u_xpb_out[66][681],u_xpb_out[67][681],u_xpb_out[68][681],u_xpb_out[69][681],u_xpb_out[70][681],u_xpb_out[71][681],u_xpb_out[72][681],u_xpb_out[73][681],u_xpb_out[74][681],u_xpb_out[75][681],u_xpb_out[76][681],u_xpb_out[77][681],u_xpb_out[78][681],u_xpb_out[79][681],u_xpb_out[80][681],u_xpb_out[81][681],u_xpb_out[82][681],u_xpb_out[83][681],u_xpb_out[84][681],u_xpb_out[85][681],u_xpb_out[86][681],u_xpb_out[87][681],u_xpb_out[88][681],u_xpb_out[89][681],u_xpb_out[90][681],u_xpb_out[91][681],u_xpb_out[92][681],u_xpb_out[93][681],u_xpb_out[94][681],u_xpb_out[95][681],u_xpb_out[96][681],u_xpb_out[97][681],u_xpb_out[98][681],u_xpb_out[99][681],u_xpb_out[100][681],u_xpb_out[101][681],u_xpb_out[102][681],u_xpb_out[103][681],u_xpb_out[104][681],u_xpb_out[105][681]};

assign col_out_682 = {u_xpb_out[0][682],u_xpb_out[1][682],u_xpb_out[2][682],u_xpb_out[3][682],u_xpb_out[4][682],u_xpb_out[5][682],u_xpb_out[6][682],u_xpb_out[7][682],u_xpb_out[8][682],u_xpb_out[9][682],u_xpb_out[10][682],u_xpb_out[11][682],u_xpb_out[12][682],u_xpb_out[13][682],u_xpb_out[14][682],u_xpb_out[15][682],u_xpb_out[16][682],u_xpb_out[17][682],u_xpb_out[18][682],u_xpb_out[19][682],u_xpb_out[20][682],u_xpb_out[21][682],u_xpb_out[22][682],u_xpb_out[23][682],u_xpb_out[24][682],u_xpb_out[25][682],u_xpb_out[26][682],u_xpb_out[27][682],u_xpb_out[28][682],u_xpb_out[29][682],u_xpb_out[30][682],u_xpb_out[31][682],u_xpb_out[32][682],u_xpb_out[33][682],u_xpb_out[34][682],u_xpb_out[35][682],u_xpb_out[36][682],u_xpb_out[37][682],u_xpb_out[38][682],u_xpb_out[39][682],u_xpb_out[40][682],u_xpb_out[41][682],u_xpb_out[42][682],u_xpb_out[43][682],u_xpb_out[44][682],u_xpb_out[45][682],u_xpb_out[46][682],u_xpb_out[47][682],u_xpb_out[48][682],u_xpb_out[49][682],u_xpb_out[50][682],u_xpb_out[51][682],u_xpb_out[52][682],u_xpb_out[53][682],u_xpb_out[54][682],u_xpb_out[55][682],u_xpb_out[56][682],u_xpb_out[57][682],u_xpb_out[58][682],u_xpb_out[59][682],u_xpb_out[60][682],u_xpb_out[61][682],u_xpb_out[62][682],u_xpb_out[63][682],u_xpb_out[64][682],u_xpb_out[65][682],u_xpb_out[66][682],u_xpb_out[67][682],u_xpb_out[68][682],u_xpb_out[69][682],u_xpb_out[70][682],u_xpb_out[71][682],u_xpb_out[72][682],u_xpb_out[73][682],u_xpb_out[74][682],u_xpb_out[75][682],u_xpb_out[76][682],u_xpb_out[77][682],u_xpb_out[78][682],u_xpb_out[79][682],u_xpb_out[80][682],u_xpb_out[81][682],u_xpb_out[82][682],u_xpb_out[83][682],u_xpb_out[84][682],u_xpb_out[85][682],u_xpb_out[86][682],u_xpb_out[87][682],u_xpb_out[88][682],u_xpb_out[89][682],u_xpb_out[90][682],u_xpb_out[91][682],u_xpb_out[92][682],u_xpb_out[93][682],u_xpb_out[94][682],u_xpb_out[95][682],u_xpb_out[96][682],u_xpb_out[97][682],u_xpb_out[98][682],u_xpb_out[99][682],u_xpb_out[100][682],u_xpb_out[101][682],u_xpb_out[102][682],u_xpb_out[103][682],u_xpb_out[104][682],u_xpb_out[105][682]};

assign col_out_683 = {u_xpb_out[0][683],u_xpb_out[1][683],u_xpb_out[2][683],u_xpb_out[3][683],u_xpb_out[4][683],u_xpb_out[5][683],u_xpb_out[6][683],u_xpb_out[7][683],u_xpb_out[8][683],u_xpb_out[9][683],u_xpb_out[10][683],u_xpb_out[11][683],u_xpb_out[12][683],u_xpb_out[13][683],u_xpb_out[14][683],u_xpb_out[15][683],u_xpb_out[16][683],u_xpb_out[17][683],u_xpb_out[18][683],u_xpb_out[19][683],u_xpb_out[20][683],u_xpb_out[21][683],u_xpb_out[22][683],u_xpb_out[23][683],u_xpb_out[24][683],u_xpb_out[25][683],u_xpb_out[26][683],u_xpb_out[27][683],u_xpb_out[28][683],u_xpb_out[29][683],u_xpb_out[30][683],u_xpb_out[31][683],u_xpb_out[32][683],u_xpb_out[33][683],u_xpb_out[34][683],u_xpb_out[35][683],u_xpb_out[36][683],u_xpb_out[37][683],u_xpb_out[38][683],u_xpb_out[39][683],u_xpb_out[40][683],u_xpb_out[41][683],u_xpb_out[42][683],u_xpb_out[43][683],u_xpb_out[44][683],u_xpb_out[45][683],u_xpb_out[46][683],u_xpb_out[47][683],u_xpb_out[48][683],u_xpb_out[49][683],u_xpb_out[50][683],u_xpb_out[51][683],u_xpb_out[52][683],u_xpb_out[53][683],u_xpb_out[54][683],u_xpb_out[55][683],u_xpb_out[56][683],u_xpb_out[57][683],u_xpb_out[58][683],u_xpb_out[59][683],u_xpb_out[60][683],u_xpb_out[61][683],u_xpb_out[62][683],u_xpb_out[63][683],u_xpb_out[64][683],u_xpb_out[65][683],u_xpb_out[66][683],u_xpb_out[67][683],u_xpb_out[68][683],u_xpb_out[69][683],u_xpb_out[70][683],u_xpb_out[71][683],u_xpb_out[72][683],u_xpb_out[73][683],u_xpb_out[74][683],u_xpb_out[75][683],u_xpb_out[76][683],u_xpb_out[77][683],u_xpb_out[78][683],u_xpb_out[79][683],u_xpb_out[80][683],u_xpb_out[81][683],u_xpb_out[82][683],u_xpb_out[83][683],u_xpb_out[84][683],u_xpb_out[85][683],u_xpb_out[86][683],u_xpb_out[87][683],u_xpb_out[88][683],u_xpb_out[89][683],u_xpb_out[90][683],u_xpb_out[91][683],u_xpb_out[92][683],u_xpb_out[93][683],u_xpb_out[94][683],u_xpb_out[95][683],u_xpb_out[96][683],u_xpb_out[97][683],u_xpb_out[98][683],u_xpb_out[99][683],u_xpb_out[100][683],u_xpb_out[101][683],u_xpb_out[102][683],u_xpb_out[103][683],u_xpb_out[104][683],u_xpb_out[105][683]};

assign col_out_684 = {u_xpb_out[0][684],u_xpb_out[1][684],u_xpb_out[2][684],u_xpb_out[3][684],u_xpb_out[4][684],u_xpb_out[5][684],u_xpb_out[6][684],u_xpb_out[7][684],u_xpb_out[8][684],u_xpb_out[9][684],u_xpb_out[10][684],u_xpb_out[11][684],u_xpb_out[12][684],u_xpb_out[13][684],u_xpb_out[14][684],u_xpb_out[15][684],u_xpb_out[16][684],u_xpb_out[17][684],u_xpb_out[18][684],u_xpb_out[19][684],u_xpb_out[20][684],u_xpb_out[21][684],u_xpb_out[22][684],u_xpb_out[23][684],u_xpb_out[24][684],u_xpb_out[25][684],u_xpb_out[26][684],u_xpb_out[27][684],u_xpb_out[28][684],u_xpb_out[29][684],u_xpb_out[30][684],u_xpb_out[31][684],u_xpb_out[32][684],u_xpb_out[33][684],u_xpb_out[34][684],u_xpb_out[35][684],u_xpb_out[36][684],u_xpb_out[37][684],u_xpb_out[38][684],u_xpb_out[39][684],u_xpb_out[40][684],u_xpb_out[41][684],u_xpb_out[42][684],u_xpb_out[43][684],u_xpb_out[44][684],u_xpb_out[45][684],u_xpb_out[46][684],u_xpb_out[47][684],u_xpb_out[48][684],u_xpb_out[49][684],u_xpb_out[50][684],u_xpb_out[51][684],u_xpb_out[52][684],u_xpb_out[53][684],u_xpb_out[54][684],u_xpb_out[55][684],u_xpb_out[56][684],u_xpb_out[57][684],u_xpb_out[58][684],u_xpb_out[59][684],u_xpb_out[60][684],u_xpb_out[61][684],u_xpb_out[62][684],u_xpb_out[63][684],u_xpb_out[64][684],u_xpb_out[65][684],u_xpb_out[66][684],u_xpb_out[67][684],u_xpb_out[68][684],u_xpb_out[69][684],u_xpb_out[70][684],u_xpb_out[71][684],u_xpb_out[72][684],u_xpb_out[73][684],u_xpb_out[74][684],u_xpb_out[75][684],u_xpb_out[76][684],u_xpb_out[77][684],u_xpb_out[78][684],u_xpb_out[79][684],u_xpb_out[80][684],u_xpb_out[81][684],u_xpb_out[82][684],u_xpb_out[83][684],u_xpb_out[84][684],u_xpb_out[85][684],u_xpb_out[86][684],u_xpb_out[87][684],u_xpb_out[88][684],u_xpb_out[89][684],u_xpb_out[90][684],u_xpb_out[91][684],u_xpb_out[92][684],u_xpb_out[93][684],u_xpb_out[94][684],u_xpb_out[95][684],u_xpb_out[96][684],u_xpb_out[97][684],u_xpb_out[98][684],u_xpb_out[99][684],u_xpb_out[100][684],u_xpb_out[101][684],u_xpb_out[102][684],u_xpb_out[103][684],u_xpb_out[104][684],u_xpb_out[105][684]};

assign col_out_685 = {u_xpb_out[0][685],u_xpb_out[1][685],u_xpb_out[2][685],u_xpb_out[3][685],u_xpb_out[4][685],u_xpb_out[5][685],u_xpb_out[6][685],u_xpb_out[7][685],u_xpb_out[8][685],u_xpb_out[9][685],u_xpb_out[10][685],u_xpb_out[11][685],u_xpb_out[12][685],u_xpb_out[13][685],u_xpb_out[14][685],u_xpb_out[15][685],u_xpb_out[16][685],u_xpb_out[17][685],u_xpb_out[18][685],u_xpb_out[19][685],u_xpb_out[20][685],u_xpb_out[21][685],u_xpb_out[22][685],u_xpb_out[23][685],u_xpb_out[24][685],u_xpb_out[25][685],u_xpb_out[26][685],u_xpb_out[27][685],u_xpb_out[28][685],u_xpb_out[29][685],u_xpb_out[30][685],u_xpb_out[31][685],u_xpb_out[32][685],u_xpb_out[33][685],u_xpb_out[34][685],u_xpb_out[35][685],u_xpb_out[36][685],u_xpb_out[37][685],u_xpb_out[38][685],u_xpb_out[39][685],u_xpb_out[40][685],u_xpb_out[41][685],u_xpb_out[42][685],u_xpb_out[43][685],u_xpb_out[44][685],u_xpb_out[45][685],u_xpb_out[46][685],u_xpb_out[47][685],u_xpb_out[48][685],u_xpb_out[49][685],u_xpb_out[50][685],u_xpb_out[51][685],u_xpb_out[52][685],u_xpb_out[53][685],u_xpb_out[54][685],u_xpb_out[55][685],u_xpb_out[56][685],u_xpb_out[57][685],u_xpb_out[58][685],u_xpb_out[59][685],u_xpb_out[60][685],u_xpb_out[61][685],u_xpb_out[62][685],u_xpb_out[63][685],u_xpb_out[64][685],u_xpb_out[65][685],u_xpb_out[66][685],u_xpb_out[67][685],u_xpb_out[68][685],u_xpb_out[69][685],u_xpb_out[70][685],u_xpb_out[71][685],u_xpb_out[72][685],u_xpb_out[73][685],u_xpb_out[74][685],u_xpb_out[75][685],u_xpb_out[76][685],u_xpb_out[77][685],u_xpb_out[78][685],u_xpb_out[79][685],u_xpb_out[80][685],u_xpb_out[81][685],u_xpb_out[82][685],u_xpb_out[83][685],u_xpb_out[84][685],u_xpb_out[85][685],u_xpb_out[86][685],u_xpb_out[87][685],u_xpb_out[88][685],u_xpb_out[89][685],u_xpb_out[90][685],u_xpb_out[91][685],u_xpb_out[92][685],u_xpb_out[93][685],u_xpb_out[94][685],u_xpb_out[95][685],u_xpb_out[96][685],u_xpb_out[97][685],u_xpb_out[98][685],u_xpb_out[99][685],u_xpb_out[100][685],u_xpb_out[101][685],u_xpb_out[102][685],u_xpb_out[103][685],u_xpb_out[104][685],u_xpb_out[105][685]};

assign col_out_686 = {u_xpb_out[0][686],u_xpb_out[1][686],u_xpb_out[2][686],u_xpb_out[3][686],u_xpb_out[4][686],u_xpb_out[5][686],u_xpb_out[6][686],u_xpb_out[7][686],u_xpb_out[8][686],u_xpb_out[9][686],u_xpb_out[10][686],u_xpb_out[11][686],u_xpb_out[12][686],u_xpb_out[13][686],u_xpb_out[14][686],u_xpb_out[15][686],u_xpb_out[16][686],u_xpb_out[17][686],u_xpb_out[18][686],u_xpb_out[19][686],u_xpb_out[20][686],u_xpb_out[21][686],u_xpb_out[22][686],u_xpb_out[23][686],u_xpb_out[24][686],u_xpb_out[25][686],u_xpb_out[26][686],u_xpb_out[27][686],u_xpb_out[28][686],u_xpb_out[29][686],u_xpb_out[30][686],u_xpb_out[31][686],u_xpb_out[32][686],u_xpb_out[33][686],u_xpb_out[34][686],u_xpb_out[35][686],u_xpb_out[36][686],u_xpb_out[37][686],u_xpb_out[38][686],u_xpb_out[39][686],u_xpb_out[40][686],u_xpb_out[41][686],u_xpb_out[42][686],u_xpb_out[43][686],u_xpb_out[44][686],u_xpb_out[45][686],u_xpb_out[46][686],u_xpb_out[47][686],u_xpb_out[48][686],u_xpb_out[49][686],u_xpb_out[50][686],u_xpb_out[51][686],u_xpb_out[52][686],u_xpb_out[53][686],u_xpb_out[54][686],u_xpb_out[55][686],u_xpb_out[56][686],u_xpb_out[57][686],u_xpb_out[58][686],u_xpb_out[59][686],u_xpb_out[60][686],u_xpb_out[61][686],u_xpb_out[62][686],u_xpb_out[63][686],u_xpb_out[64][686],u_xpb_out[65][686],u_xpb_out[66][686],u_xpb_out[67][686],u_xpb_out[68][686],u_xpb_out[69][686],u_xpb_out[70][686],u_xpb_out[71][686],u_xpb_out[72][686],u_xpb_out[73][686],u_xpb_out[74][686],u_xpb_out[75][686],u_xpb_out[76][686],u_xpb_out[77][686],u_xpb_out[78][686],u_xpb_out[79][686],u_xpb_out[80][686],u_xpb_out[81][686],u_xpb_out[82][686],u_xpb_out[83][686],u_xpb_out[84][686],u_xpb_out[85][686],u_xpb_out[86][686],u_xpb_out[87][686],u_xpb_out[88][686],u_xpb_out[89][686],u_xpb_out[90][686],u_xpb_out[91][686],u_xpb_out[92][686],u_xpb_out[93][686],u_xpb_out[94][686],u_xpb_out[95][686],u_xpb_out[96][686],u_xpb_out[97][686],u_xpb_out[98][686],u_xpb_out[99][686],u_xpb_out[100][686],u_xpb_out[101][686],u_xpb_out[102][686],u_xpb_out[103][686],u_xpb_out[104][686],u_xpb_out[105][686]};

assign col_out_687 = {u_xpb_out[0][687],u_xpb_out[1][687],u_xpb_out[2][687],u_xpb_out[3][687],u_xpb_out[4][687],u_xpb_out[5][687],u_xpb_out[6][687],u_xpb_out[7][687],u_xpb_out[8][687],u_xpb_out[9][687],u_xpb_out[10][687],u_xpb_out[11][687],u_xpb_out[12][687],u_xpb_out[13][687],u_xpb_out[14][687],u_xpb_out[15][687],u_xpb_out[16][687],u_xpb_out[17][687],u_xpb_out[18][687],u_xpb_out[19][687],u_xpb_out[20][687],u_xpb_out[21][687],u_xpb_out[22][687],u_xpb_out[23][687],u_xpb_out[24][687],u_xpb_out[25][687],u_xpb_out[26][687],u_xpb_out[27][687],u_xpb_out[28][687],u_xpb_out[29][687],u_xpb_out[30][687],u_xpb_out[31][687],u_xpb_out[32][687],u_xpb_out[33][687],u_xpb_out[34][687],u_xpb_out[35][687],u_xpb_out[36][687],u_xpb_out[37][687],u_xpb_out[38][687],u_xpb_out[39][687],u_xpb_out[40][687],u_xpb_out[41][687],u_xpb_out[42][687],u_xpb_out[43][687],u_xpb_out[44][687],u_xpb_out[45][687],u_xpb_out[46][687],u_xpb_out[47][687],u_xpb_out[48][687],u_xpb_out[49][687],u_xpb_out[50][687],u_xpb_out[51][687],u_xpb_out[52][687],u_xpb_out[53][687],u_xpb_out[54][687],u_xpb_out[55][687],u_xpb_out[56][687],u_xpb_out[57][687],u_xpb_out[58][687],u_xpb_out[59][687],u_xpb_out[60][687],u_xpb_out[61][687],u_xpb_out[62][687],u_xpb_out[63][687],u_xpb_out[64][687],u_xpb_out[65][687],u_xpb_out[66][687],u_xpb_out[67][687],u_xpb_out[68][687],u_xpb_out[69][687],u_xpb_out[70][687],u_xpb_out[71][687],u_xpb_out[72][687],u_xpb_out[73][687],u_xpb_out[74][687],u_xpb_out[75][687],u_xpb_out[76][687],u_xpb_out[77][687],u_xpb_out[78][687],u_xpb_out[79][687],u_xpb_out[80][687],u_xpb_out[81][687],u_xpb_out[82][687],u_xpb_out[83][687],u_xpb_out[84][687],u_xpb_out[85][687],u_xpb_out[86][687],u_xpb_out[87][687],u_xpb_out[88][687],u_xpb_out[89][687],u_xpb_out[90][687],u_xpb_out[91][687],u_xpb_out[92][687],u_xpb_out[93][687],u_xpb_out[94][687],u_xpb_out[95][687],u_xpb_out[96][687],u_xpb_out[97][687],u_xpb_out[98][687],u_xpb_out[99][687],u_xpb_out[100][687],u_xpb_out[101][687],u_xpb_out[102][687],u_xpb_out[103][687],u_xpb_out[104][687],u_xpb_out[105][687]};

assign col_out_688 = {u_xpb_out[0][688],u_xpb_out[1][688],u_xpb_out[2][688],u_xpb_out[3][688],u_xpb_out[4][688],u_xpb_out[5][688],u_xpb_out[6][688],u_xpb_out[7][688],u_xpb_out[8][688],u_xpb_out[9][688],u_xpb_out[10][688],u_xpb_out[11][688],u_xpb_out[12][688],u_xpb_out[13][688],u_xpb_out[14][688],u_xpb_out[15][688],u_xpb_out[16][688],u_xpb_out[17][688],u_xpb_out[18][688],u_xpb_out[19][688],u_xpb_out[20][688],u_xpb_out[21][688],u_xpb_out[22][688],u_xpb_out[23][688],u_xpb_out[24][688],u_xpb_out[25][688],u_xpb_out[26][688],u_xpb_out[27][688],u_xpb_out[28][688],u_xpb_out[29][688],u_xpb_out[30][688],u_xpb_out[31][688],u_xpb_out[32][688],u_xpb_out[33][688],u_xpb_out[34][688],u_xpb_out[35][688],u_xpb_out[36][688],u_xpb_out[37][688],u_xpb_out[38][688],u_xpb_out[39][688],u_xpb_out[40][688],u_xpb_out[41][688],u_xpb_out[42][688],u_xpb_out[43][688],u_xpb_out[44][688],u_xpb_out[45][688],u_xpb_out[46][688],u_xpb_out[47][688],u_xpb_out[48][688],u_xpb_out[49][688],u_xpb_out[50][688],u_xpb_out[51][688],u_xpb_out[52][688],u_xpb_out[53][688],u_xpb_out[54][688],u_xpb_out[55][688],u_xpb_out[56][688],u_xpb_out[57][688],u_xpb_out[58][688],u_xpb_out[59][688],u_xpb_out[60][688],u_xpb_out[61][688],u_xpb_out[62][688],u_xpb_out[63][688],u_xpb_out[64][688],u_xpb_out[65][688],u_xpb_out[66][688],u_xpb_out[67][688],u_xpb_out[68][688],u_xpb_out[69][688],u_xpb_out[70][688],u_xpb_out[71][688],u_xpb_out[72][688],u_xpb_out[73][688],u_xpb_out[74][688],u_xpb_out[75][688],u_xpb_out[76][688],u_xpb_out[77][688],u_xpb_out[78][688],u_xpb_out[79][688],u_xpb_out[80][688],u_xpb_out[81][688],u_xpb_out[82][688],u_xpb_out[83][688],u_xpb_out[84][688],u_xpb_out[85][688],u_xpb_out[86][688],u_xpb_out[87][688],u_xpb_out[88][688],u_xpb_out[89][688],u_xpb_out[90][688],u_xpb_out[91][688],u_xpb_out[92][688],u_xpb_out[93][688],u_xpb_out[94][688],u_xpb_out[95][688],u_xpb_out[96][688],u_xpb_out[97][688],u_xpb_out[98][688],u_xpb_out[99][688],u_xpb_out[100][688],u_xpb_out[101][688],u_xpb_out[102][688],u_xpb_out[103][688],u_xpb_out[104][688],u_xpb_out[105][688]};

assign col_out_689 = {u_xpb_out[0][689],u_xpb_out[1][689],u_xpb_out[2][689],u_xpb_out[3][689],u_xpb_out[4][689],u_xpb_out[5][689],u_xpb_out[6][689],u_xpb_out[7][689],u_xpb_out[8][689],u_xpb_out[9][689],u_xpb_out[10][689],u_xpb_out[11][689],u_xpb_out[12][689],u_xpb_out[13][689],u_xpb_out[14][689],u_xpb_out[15][689],u_xpb_out[16][689],u_xpb_out[17][689],u_xpb_out[18][689],u_xpb_out[19][689],u_xpb_out[20][689],u_xpb_out[21][689],u_xpb_out[22][689],u_xpb_out[23][689],u_xpb_out[24][689],u_xpb_out[25][689],u_xpb_out[26][689],u_xpb_out[27][689],u_xpb_out[28][689],u_xpb_out[29][689],u_xpb_out[30][689],u_xpb_out[31][689],u_xpb_out[32][689],u_xpb_out[33][689],u_xpb_out[34][689],u_xpb_out[35][689],u_xpb_out[36][689],u_xpb_out[37][689],u_xpb_out[38][689],u_xpb_out[39][689],u_xpb_out[40][689],u_xpb_out[41][689],u_xpb_out[42][689],u_xpb_out[43][689],u_xpb_out[44][689],u_xpb_out[45][689],u_xpb_out[46][689],u_xpb_out[47][689],u_xpb_out[48][689],u_xpb_out[49][689],u_xpb_out[50][689],u_xpb_out[51][689],u_xpb_out[52][689],u_xpb_out[53][689],u_xpb_out[54][689],u_xpb_out[55][689],u_xpb_out[56][689],u_xpb_out[57][689],u_xpb_out[58][689],u_xpb_out[59][689],u_xpb_out[60][689],u_xpb_out[61][689],u_xpb_out[62][689],u_xpb_out[63][689],u_xpb_out[64][689],u_xpb_out[65][689],u_xpb_out[66][689],u_xpb_out[67][689],u_xpb_out[68][689],u_xpb_out[69][689],u_xpb_out[70][689],u_xpb_out[71][689],u_xpb_out[72][689],u_xpb_out[73][689],u_xpb_out[74][689],u_xpb_out[75][689],u_xpb_out[76][689],u_xpb_out[77][689],u_xpb_out[78][689],u_xpb_out[79][689],u_xpb_out[80][689],u_xpb_out[81][689],u_xpb_out[82][689],u_xpb_out[83][689],u_xpb_out[84][689],u_xpb_out[85][689],u_xpb_out[86][689],u_xpb_out[87][689],u_xpb_out[88][689],u_xpb_out[89][689],u_xpb_out[90][689],u_xpb_out[91][689],u_xpb_out[92][689],u_xpb_out[93][689],u_xpb_out[94][689],u_xpb_out[95][689],u_xpb_out[96][689],u_xpb_out[97][689],u_xpb_out[98][689],u_xpb_out[99][689],u_xpb_out[100][689],u_xpb_out[101][689],u_xpb_out[102][689],u_xpb_out[103][689],u_xpb_out[104][689],u_xpb_out[105][689]};

assign col_out_690 = {u_xpb_out[0][690],u_xpb_out[1][690],u_xpb_out[2][690],u_xpb_out[3][690],u_xpb_out[4][690],u_xpb_out[5][690],u_xpb_out[6][690],u_xpb_out[7][690],u_xpb_out[8][690],u_xpb_out[9][690],u_xpb_out[10][690],u_xpb_out[11][690],u_xpb_out[12][690],u_xpb_out[13][690],u_xpb_out[14][690],u_xpb_out[15][690],u_xpb_out[16][690],u_xpb_out[17][690],u_xpb_out[18][690],u_xpb_out[19][690],u_xpb_out[20][690],u_xpb_out[21][690],u_xpb_out[22][690],u_xpb_out[23][690],u_xpb_out[24][690],u_xpb_out[25][690],u_xpb_out[26][690],u_xpb_out[27][690],u_xpb_out[28][690],u_xpb_out[29][690],u_xpb_out[30][690],u_xpb_out[31][690],u_xpb_out[32][690],u_xpb_out[33][690],u_xpb_out[34][690],u_xpb_out[35][690],u_xpb_out[36][690],u_xpb_out[37][690],u_xpb_out[38][690],u_xpb_out[39][690],u_xpb_out[40][690],u_xpb_out[41][690],u_xpb_out[42][690],u_xpb_out[43][690],u_xpb_out[44][690],u_xpb_out[45][690],u_xpb_out[46][690],u_xpb_out[47][690],u_xpb_out[48][690],u_xpb_out[49][690],u_xpb_out[50][690],u_xpb_out[51][690],u_xpb_out[52][690],u_xpb_out[53][690],u_xpb_out[54][690],u_xpb_out[55][690],u_xpb_out[56][690],u_xpb_out[57][690],u_xpb_out[58][690],u_xpb_out[59][690],u_xpb_out[60][690],u_xpb_out[61][690],u_xpb_out[62][690],u_xpb_out[63][690],u_xpb_out[64][690],u_xpb_out[65][690],u_xpb_out[66][690],u_xpb_out[67][690],u_xpb_out[68][690],u_xpb_out[69][690],u_xpb_out[70][690],u_xpb_out[71][690],u_xpb_out[72][690],u_xpb_out[73][690],u_xpb_out[74][690],u_xpb_out[75][690],u_xpb_out[76][690],u_xpb_out[77][690],u_xpb_out[78][690],u_xpb_out[79][690],u_xpb_out[80][690],u_xpb_out[81][690],u_xpb_out[82][690],u_xpb_out[83][690],u_xpb_out[84][690],u_xpb_out[85][690],u_xpb_out[86][690],u_xpb_out[87][690],u_xpb_out[88][690],u_xpb_out[89][690],u_xpb_out[90][690],u_xpb_out[91][690],u_xpb_out[92][690],u_xpb_out[93][690],u_xpb_out[94][690],u_xpb_out[95][690],u_xpb_out[96][690],u_xpb_out[97][690],u_xpb_out[98][690],u_xpb_out[99][690],u_xpb_out[100][690],u_xpb_out[101][690],u_xpb_out[102][690],u_xpb_out[103][690],u_xpb_out[104][690],u_xpb_out[105][690]};

assign col_out_691 = {u_xpb_out[0][691],u_xpb_out[1][691],u_xpb_out[2][691],u_xpb_out[3][691],u_xpb_out[4][691],u_xpb_out[5][691],u_xpb_out[6][691],u_xpb_out[7][691],u_xpb_out[8][691],u_xpb_out[9][691],u_xpb_out[10][691],u_xpb_out[11][691],u_xpb_out[12][691],u_xpb_out[13][691],u_xpb_out[14][691],u_xpb_out[15][691],u_xpb_out[16][691],u_xpb_out[17][691],u_xpb_out[18][691],u_xpb_out[19][691],u_xpb_out[20][691],u_xpb_out[21][691],u_xpb_out[22][691],u_xpb_out[23][691],u_xpb_out[24][691],u_xpb_out[25][691],u_xpb_out[26][691],u_xpb_out[27][691],u_xpb_out[28][691],u_xpb_out[29][691],u_xpb_out[30][691],u_xpb_out[31][691],u_xpb_out[32][691],u_xpb_out[33][691],u_xpb_out[34][691],u_xpb_out[35][691],u_xpb_out[36][691],u_xpb_out[37][691],u_xpb_out[38][691],u_xpb_out[39][691],u_xpb_out[40][691],u_xpb_out[41][691],u_xpb_out[42][691],u_xpb_out[43][691],u_xpb_out[44][691],u_xpb_out[45][691],u_xpb_out[46][691],u_xpb_out[47][691],u_xpb_out[48][691],u_xpb_out[49][691],u_xpb_out[50][691],u_xpb_out[51][691],u_xpb_out[52][691],u_xpb_out[53][691],u_xpb_out[54][691],u_xpb_out[55][691],u_xpb_out[56][691],u_xpb_out[57][691],u_xpb_out[58][691],u_xpb_out[59][691],u_xpb_out[60][691],u_xpb_out[61][691],u_xpb_out[62][691],u_xpb_out[63][691],u_xpb_out[64][691],u_xpb_out[65][691],u_xpb_out[66][691],u_xpb_out[67][691],u_xpb_out[68][691],u_xpb_out[69][691],u_xpb_out[70][691],u_xpb_out[71][691],u_xpb_out[72][691],u_xpb_out[73][691],u_xpb_out[74][691],u_xpb_out[75][691],u_xpb_out[76][691],u_xpb_out[77][691],u_xpb_out[78][691],u_xpb_out[79][691],u_xpb_out[80][691],u_xpb_out[81][691],u_xpb_out[82][691],u_xpb_out[83][691],u_xpb_out[84][691],u_xpb_out[85][691],u_xpb_out[86][691],u_xpb_out[87][691],u_xpb_out[88][691],u_xpb_out[89][691],u_xpb_out[90][691],u_xpb_out[91][691],u_xpb_out[92][691],u_xpb_out[93][691],u_xpb_out[94][691],u_xpb_out[95][691],u_xpb_out[96][691],u_xpb_out[97][691],u_xpb_out[98][691],u_xpb_out[99][691],u_xpb_out[100][691],u_xpb_out[101][691],u_xpb_out[102][691],u_xpb_out[103][691],u_xpb_out[104][691],u_xpb_out[105][691]};

assign col_out_692 = {u_xpb_out[0][692],u_xpb_out[1][692],u_xpb_out[2][692],u_xpb_out[3][692],u_xpb_out[4][692],u_xpb_out[5][692],u_xpb_out[6][692],u_xpb_out[7][692],u_xpb_out[8][692],u_xpb_out[9][692],u_xpb_out[10][692],u_xpb_out[11][692],u_xpb_out[12][692],u_xpb_out[13][692],u_xpb_out[14][692],u_xpb_out[15][692],u_xpb_out[16][692],u_xpb_out[17][692],u_xpb_out[18][692],u_xpb_out[19][692],u_xpb_out[20][692],u_xpb_out[21][692],u_xpb_out[22][692],u_xpb_out[23][692],u_xpb_out[24][692],u_xpb_out[25][692],u_xpb_out[26][692],u_xpb_out[27][692],u_xpb_out[28][692],u_xpb_out[29][692],u_xpb_out[30][692],u_xpb_out[31][692],u_xpb_out[32][692],u_xpb_out[33][692],u_xpb_out[34][692],u_xpb_out[35][692],u_xpb_out[36][692],u_xpb_out[37][692],u_xpb_out[38][692],u_xpb_out[39][692],u_xpb_out[40][692],u_xpb_out[41][692],u_xpb_out[42][692],u_xpb_out[43][692],u_xpb_out[44][692],u_xpb_out[45][692],u_xpb_out[46][692],u_xpb_out[47][692],u_xpb_out[48][692],u_xpb_out[49][692],u_xpb_out[50][692],u_xpb_out[51][692],u_xpb_out[52][692],u_xpb_out[53][692],u_xpb_out[54][692],u_xpb_out[55][692],u_xpb_out[56][692],u_xpb_out[57][692],u_xpb_out[58][692],u_xpb_out[59][692],u_xpb_out[60][692],u_xpb_out[61][692],u_xpb_out[62][692],u_xpb_out[63][692],u_xpb_out[64][692],u_xpb_out[65][692],u_xpb_out[66][692],u_xpb_out[67][692],u_xpb_out[68][692],u_xpb_out[69][692],u_xpb_out[70][692],u_xpb_out[71][692],u_xpb_out[72][692],u_xpb_out[73][692],u_xpb_out[74][692],u_xpb_out[75][692],u_xpb_out[76][692],u_xpb_out[77][692],u_xpb_out[78][692],u_xpb_out[79][692],u_xpb_out[80][692],u_xpb_out[81][692],u_xpb_out[82][692],u_xpb_out[83][692],u_xpb_out[84][692],u_xpb_out[85][692],u_xpb_out[86][692],u_xpb_out[87][692],u_xpb_out[88][692],u_xpb_out[89][692],u_xpb_out[90][692],u_xpb_out[91][692],u_xpb_out[92][692],u_xpb_out[93][692],u_xpb_out[94][692],u_xpb_out[95][692],u_xpb_out[96][692],u_xpb_out[97][692],u_xpb_out[98][692],u_xpb_out[99][692],u_xpb_out[100][692],u_xpb_out[101][692],u_xpb_out[102][692],u_xpb_out[103][692],u_xpb_out[104][692],u_xpb_out[105][692]};

assign col_out_693 = {u_xpb_out[0][693],u_xpb_out[1][693],u_xpb_out[2][693],u_xpb_out[3][693],u_xpb_out[4][693],u_xpb_out[5][693],u_xpb_out[6][693],u_xpb_out[7][693],u_xpb_out[8][693],u_xpb_out[9][693],u_xpb_out[10][693],u_xpb_out[11][693],u_xpb_out[12][693],u_xpb_out[13][693],u_xpb_out[14][693],u_xpb_out[15][693],u_xpb_out[16][693],u_xpb_out[17][693],u_xpb_out[18][693],u_xpb_out[19][693],u_xpb_out[20][693],u_xpb_out[21][693],u_xpb_out[22][693],u_xpb_out[23][693],u_xpb_out[24][693],u_xpb_out[25][693],u_xpb_out[26][693],u_xpb_out[27][693],u_xpb_out[28][693],u_xpb_out[29][693],u_xpb_out[30][693],u_xpb_out[31][693],u_xpb_out[32][693],u_xpb_out[33][693],u_xpb_out[34][693],u_xpb_out[35][693],u_xpb_out[36][693],u_xpb_out[37][693],u_xpb_out[38][693],u_xpb_out[39][693],u_xpb_out[40][693],u_xpb_out[41][693],u_xpb_out[42][693],u_xpb_out[43][693],u_xpb_out[44][693],u_xpb_out[45][693],u_xpb_out[46][693],u_xpb_out[47][693],u_xpb_out[48][693],u_xpb_out[49][693],u_xpb_out[50][693],u_xpb_out[51][693],u_xpb_out[52][693],u_xpb_out[53][693],u_xpb_out[54][693],u_xpb_out[55][693],u_xpb_out[56][693],u_xpb_out[57][693],u_xpb_out[58][693],u_xpb_out[59][693],u_xpb_out[60][693],u_xpb_out[61][693],u_xpb_out[62][693],u_xpb_out[63][693],u_xpb_out[64][693],u_xpb_out[65][693],u_xpb_out[66][693],u_xpb_out[67][693],u_xpb_out[68][693],u_xpb_out[69][693],u_xpb_out[70][693],u_xpb_out[71][693],u_xpb_out[72][693],u_xpb_out[73][693],u_xpb_out[74][693],u_xpb_out[75][693],u_xpb_out[76][693],u_xpb_out[77][693],u_xpb_out[78][693],u_xpb_out[79][693],u_xpb_out[80][693],u_xpb_out[81][693],u_xpb_out[82][693],u_xpb_out[83][693],u_xpb_out[84][693],u_xpb_out[85][693],u_xpb_out[86][693],u_xpb_out[87][693],u_xpb_out[88][693],u_xpb_out[89][693],u_xpb_out[90][693],u_xpb_out[91][693],u_xpb_out[92][693],u_xpb_out[93][693],u_xpb_out[94][693],u_xpb_out[95][693],u_xpb_out[96][693],u_xpb_out[97][693],u_xpb_out[98][693],u_xpb_out[99][693],u_xpb_out[100][693],u_xpb_out[101][693],u_xpb_out[102][693],u_xpb_out[103][693],u_xpb_out[104][693],u_xpb_out[105][693]};

assign col_out_694 = {u_xpb_out[0][694],u_xpb_out[1][694],u_xpb_out[2][694],u_xpb_out[3][694],u_xpb_out[4][694],u_xpb_out[5][694],u_xpb_out[6][694],u_xpb_out[7][694],u_xpb_out[8][694],u_xpb_out[9][694],u_xpb_out[10][694],u_xpb_out[11][694],u_xpb_out[12][694],u_xpb_out[13][694],u_xpb_out[14][694],u_xpb_out[15][694],u_xpb_out[16][694],u_xpb_out[17][694],u_xpb_out[18][694],u_xpb_out[19][694],u_xpb_out[20][694],u_xpb_out[21][694],u_xpb_out[22][694],u_xpb_out[23][694],u_xpb_out[24][694],u_xpb_out[25][694],u_xpb_out[26][694],u_xpb_out[27][694],u_xpb_out[28][694],u_xpb_out[29][694],u_xpb_out[30][694],u_xpb_out[31][694],u_xpb_out[32][694],u_xpb_out[33][694],u_xpb_out[34][694],u_xpb_out[35][694],u_xpb_out[36][694],u_xpb_out[37][694],u_xpb_out[38][694],u_xpb_out[39][694],u_xpb_out[40][694],u_xpb_out[41][694],u_xpb_out[42][694],u_xpb_out[43][694],u_xpb_out[44][694],u_xpb_out[45][694],u_xpb_out[46][694],u_xpb_out[47][694],u_xpb_out[48][694],u_xpb_out[49][694],u_xpb_out[50][694],u_xpb_out[51][694],u_xpb_out[52][694],u_xpb_out[53][694],u_xpb_out[54][694],u_xpb_out[55][694],u_xpb_out[56][694],u_xpb_out[57][694],u_xpb_out[58][694],u_xpb_out[59][694],u_xpb_out[60][694],u_xpb_out[61][694],u_xpb_out[62][694],u_xpb_out[63][694],u_xpb_out[64][694],u_xpb_out[65][694],u_xpb_out[66][694],u_xpb_out[67][694],u_xpb_out[68][694],u_xpb_out[69][694],u_xpb_out[70][694],u_xpb_out[71][694],u_xpb_out[72][694],u_xpb_out[73][694],u_xpb_out[74][694],u_xpb_out[75][694],u_xpb_out[76][694],u_xpb_out[77][694],u_xpb_out[78][694],u_xpb_out[79][694],u_xpb_out[80][694],u_xpb_out[81][694],u_xpb_out[82][694],u_xpb_out[83][694],u_xpb_out[84][694],u_xpb_out[85][694],u_xpb_out[86][694],u_xpb_out[87][694],u_xpb_out[88][694],u_xpb_out[89][694],u_xpb_out[90][694],u_xpb_out[91][694],u_xpb_out[92][694],u_xpb_out[93][694],u_xpb_out[94][694],u_xpb_out[95][694],u_xpb_out[96][694],u_xpb_out[97][694],u_xpb_out[98][694],u_xpb_out[99][694],u_xpb_out[100][694],u_xpb_out[101][694],u_xpb_out[102][694],u_xpb_out[103][694],u_xpb_out[104][694],u_xpb_out[105][694]};

assign col_out_695 = {u_xpb_out[0][695],u_xpb_out[1][695],u_xpb_out[2][695],u_xpb_out[3][695],u_xpb_out[4][695],u_xpb_out[5][695],u_xpb_out[6][695],u_xpb_out[7][695],u_xpb_out[8][695],u_xpb_out[9][695],u_xpb_out[10][695],u_xpb_out[11][695],u_xpb_out[12][695],u_xpb_out[13][695],u_xpb_out[14][695],u_xpb_out[15][695],u_xpb_out[16][695],u_xpb_out[17][695],u_xpb_out[18][695],u_xpb_out[19][695],u_xpb_out[20][695],u_xpb_out[21][695],u_xpb_out[22][695],u_xpb_out[23][695],u_xpb_out[24][695],u_xpb_out[25][695],u_xpb_out[26][695],u_xpb_out[27][695],u_xpb_out[28][695],u_xpb_out[29][695],u_xpb_out[30][695],u_xpb_out[31][695],u_xpb_out[32][695],u_xpb_out[33][695],u_xpb_out[34][695],u_xpb_out[35][695],u_xpb_out[36][695],u_xpb_out[37][695],u_xpb_out[38][695],u_xpb_out[39][695],u_xpb_out[40][695],u_xpb_out[41][695],u_xpb_out[42][695],u_xpb_out[43][695],u_xpb_out[44][695],u_xpb_out[45][695],u_xpb_out[46][695],u_xpb_out[47][695],u_xpb_out[48][695],u_xpb_out[49][695],u_xpb_out[50][695],u_xpb_out[51][695],u_xpb_out[52][695],u_xpb_out[53][695],u_xpb_out[54][695],u_xpb_out[55][695],u_xpb_out[56][695],u_xpb_out[57][695],u_xpb_out[58][695],u_xpb_out[59][695],u_xpb_out[60][695],u_xpb_out[61][695],u_xpb_out[62][695],u_xpb_out[63][695],u_xpb_out[64][695],u_xpb_out[65][695],u_xpb_out[66][695],u_xpb_out[67][695],u_xpb_out[68][695],u_xpb_out[69][695],u_xpb_out[70][695],u_xpb_out[71][695],u_xpb_out[72][695],u_xpb_out[73][695],u_xpb_out[74][695],u_xpb_out[75][695],u_xpb_out[76][695],u_xpb_out[77][695],u_xpb_out[78][695],u_xpb_out[79][695],u_xpb_out[80][695],u_xpb_out[81][695],u_xpb_out[82][695],u_xpb_out[83][695],u_xpb_out[84][695],u_xpb_out[85][695],u_xpb_out[86][695],u_xpb_out[87][695],u_xpb_out[88][695],u_xpb_out[89][695],u_xpb_out[90][695],u_xpb_out[91][695],u_xpb_out[92][695],u_xpb_out[93][695],u_xpb_out[94][695],u_xpb_out[95][695],u_xpb_out[96][695],u_xpb_out[97][695],u_xpb_out[98][695],u_xpb_out[99][695],u_xpb_out[100][695],u_xpb_out[101][695],u_xpb_out[102][695],u_xpb_out[103][695],u_xpb_out[104][695],u_xpb_out[105][695]};

assign col_out_696 = {u_xpb_out[0][696],u_xpb_out[1][696],u_xpb_out[2][696],u_xpb_out[3][696],u_xpb_out[4][696],u_xpb_out[5][696],u_xpb_out[6][696],u_xpb_out[7][696],u_xpb_out[8][696],u_xpb_out[9][696],u_xpb_out[10][696],u_xpb_out[11][696],u_xpb_out[12][696],u_xpb_out[13][696],u_xpb_out[14][696],u_xpb_out[15][696],u_xpb_out[16][696],u_xpb_out[17][696],u_xpb_out[18][696],u_xpb_out[19][696],u_xpb_out[20][696],u_xpb_out[21][696],u_xpb_out[22][696],u_xpb_out[23][696],u_xpb_out[24][696],u_xpb_out[25][696],u_xpb_out[26][696],u_xpb_out[27][696],u_xpb_out[28][696],u_xpb_out[29][696],u_xpb_out[30][696],u_xpb_out[31][696],u_xpb_out[32][696],u_xpb_out[33][696],u_xpb_out[34][696],u_xpb_out[35][696],u_xpb_out[36][696],u_xpb_out[37][696],u_xpb_out[38][696],u_xpb_out[39][696],u_xpb_out[40][696],u_xpb_out[41][696],u_xpb_out[42][696],u_xpb_out[43][696],u_xpb_out[44][696],u_xpb_out[45][696],u_xpb_out[46][696],u_xpb_out[47][696],u_xpb_out[48][696],u_xpb_out[49][696],u_xpb_out[50][696],u_xpb_out[51][696],u_xpb_out[52][696],u_xpb_out[53][696],u_xpb_out[54][696],u_xpb_out[55][696],u_xpb_out[56][696],u_xpb_out[57][696],u_xpb_out[58][696],u_xpb_out[59][696],u_xpb_out[60][696],u_xpb_out[61][696],u_xpb_out[62][696],u_xpb_out[63][696],u_xpb_out[64][696],u_xpb_out[65][696],u_xpb_out[66][696],u_xpb_out[67][696],u_xpb_out[68][696],u_xpb_out[69][696],u_xpb_out[70][696],u_xpb_out[71][696],u_xpb_out[72][696],u_xpb_out[73][696],u_xpb_out[74][696],u_xpb_out[75][696],u_xpb_out[76][696],u_xpb_out[77][696],u_xpb_out[78][696],u_xpb_out[79][696],u_xpb_out[80][696],u_xpb_out[81][696],u_xpb_out[82][696],u_xpb_out[83][696],u_xpb_out[84][696],u_xpb_out[85][696],u_xpb_out[86][696],u_xpb_out[87][696],u_xpb_out[88][696],u_xpb_out[89][696],u_xpb_out[90][696],u_xpb_out[91][696],u_xpb_out[92][696],u_xpb_out[93][696],u_xpb_out[94][696],u_xpb_out[95][696],u_xpb_out[96][696],u_xpb_out[97][696],u_xpb_out[98][696],u_xpb_out[99][696],u_xpb_out[100][696],u_xpb_out[101][696],u_xpb_out[102][696],u_xpb_out[103][696],u_xpb_out[104][696],u_xpb_out[105][696]};

assign col_out_697 = {u_xpb_out[0][697],u_xpb_out[1][697],u_xpb_out[2][697],u_xpb_out[3][697],u_xpb_out[4][697],u_xpb_out[5][697],u_xpb_out[6][697],u_xpb_out[7][697],u_xpb_out[8][697],u_xpb_out[9][697],u_xpb_out[10][697],u_xpb_out[11][697],u_xpb_out[12][697],u_xpb_out[13][697],u_xpb_out[14][697],u_xpb_out[15][697],u_xpb_out[16][697],u_xpb_out[17][697],u_xpb_out[18][697],u_xpb_out[19][697],u_xpb_out[20][697],u_xpb_out[21][697],u_xpb_out[22][697],u_xpb_out[23][697],u_xpb_out[24][697],u_xpb_out[25][697],u_xpb_out[26][697],u_xpb_out[27][697],u_xpb_out[28][697],u_xpb_out[29][697],u_xpb_out[30][697],u_xpb_out[31][697],u_xpb_out[32][697],u_xpb_out[33][697],u_xpb_out[34][697],u_xpb_out[35][697],u_xpb_out[36][697],u_xpb_out[37][697],u_xpb_out[38][697],u_xpb_out[39][697],u_xpb_out[40][697],u_xpb_out[41][697],u_xpb_out[42][697],u_xpb_out[43][697],u_xpb_out[44][697],u_xpb_out[45][697],u_xpb_out[46][697],u_xpb_out[47][697],u_xpb_out[48][697],u_xpb_out[49][697],u_xpb_out[50][697],u_xpb_out[51][697],u_xpb_out[52][697],u_xpb_out[53][697],u_xpb_out[54][697],u_xpb_out[55][697],u_xpb_out[56][697],u_xpb_out[57][697],u_xpb_out[58][697],u_xpb_out[59][697],u_xpb_out[60][697],u_xpb_out[61][697],u_xpb_out[62][697],u_xpb_out[63][697],u_xpb_out[64][697],u_xpb_out[65][697],u_xpb_out[66][697],u_xpb_out[67][697],u_xpb_out[68][697],u_xpb_out[69][697],u_xpb_out[70][697],u_xpb_out[71][697],u_xpb_out[72][697],u_xpb_out[73][697],u_xpb_out[74][697],u_xpb_out[75][697],u_xpb_out[76][697],u_xpb_out[77][697],u_xpb_out[78][697],u_xpb_out[79][697],u_xpb_out[80][697],u_xpb_out[81][697],u_xpb_out[82][697],u_xpb_out[83][697],u_xpb_out[84][697],u_xpb_out[85][697],u_xpb_out[86][697],u_xpb_out[87][697],u_xpb_out[88][697],u_xpb_out[89][697],u_xpb_out[90][697],u_xpb_out[91][697],u_xpb_out[92][697],u_xpb_out[93][697],u_xpb_out[94][697],u_xpb_out[95][697],u_xpb_out[96][697],u_xpb_out[97][697],u_xpb_out[98][697],u_xpb_out[99][697],u_xpb_out[100][697],u_xpb_out[101][697],u_xpb_out[102][697],u_xpb_out[103][697],u_xpb_out[104][697],u_xpb_out[105][697]};

assign col_out_698 = {u_xpb_out[0][698],u_xpb_out[1][698],u_xpb_out[2][698],u_xpb_out[3][698],u_xpb_out[4][698],u_xpb_out[5][698],u_xpb_out[6][698],u_xpb_out[7][698],u_xpb_out[8][698],u_xpb_out[9][698],u_xpb_out[10][698],u_xpb_out[11][698],u_xpb_out[12][698],u_xpb_out[13][698],u_xpb_out[14][698],u_xpb_out[15][698],u_xpb_out[16][698],u_xpb_out[17][698],u_xpb_out[18][698],u_xpb_out[19][698],u_xpb_out[20][698],u_xpb_out[21][698],u_xpb_out[22][698],u_xpb_out[23][698],u_xpb_out[24][698],u_xpb_out[25][698],u_xpb_out[26][698],u_xpb_out[27][698],u_xpb_out[28][698],u_xpb_out[29][698],u_xpb_out[30][698],u_xpb_out[31][698],u_xpb_out[32][698],u_xpb_out[33][698],u_xpb_out[34][698],u_xpb_out[35][698],u_xpb_out[36][698],u_xpb_out[37][698],u_xpb_out[38][698],u_xpb_out[39][698],u_xpb_out[40][698],u_xpb_out[41][698],u_xpb_out[42][698],u_xpb_out[43][698],u_xpb_out[44][698],u_xpb_out[45][698],u_xpb_out[46][698],u_xpb_out[47][698],u_xpb_out[48][698],u_xpb_out[49][698],u_xpb_out[50][698],u_xpb_out[51][698],u_xpb_out[52][698],u_xpb_out[53][698],u_xpb_out[54][698],u_xpb_out[55][698],u_xpb_out[56][698],u_xpb_out[57][698],u_xpb_out[58][698],u_xpb_out[59][698],u_xpb_out[60][698],u_xpb_out[61][698],u_xpb_out[62][698],u_xpb_out[63][698],u_xpb_out[64][698],u_xpb_out[65][698],u_xpb_out[66][698],u_xpb_out[67][698],u_xpb_out[68][698],u_xpb_out[69][698],u_xpb_out[70][698],u_xpb_out[71][698],u_xpb_out[72][698],u_xpb_out[73][698],u_xpb_out[74][698],u_xpb_out[75][698],u_xpb_out[76][698],u_xpb_out[77][698],u_xpb_out[78][698],u_xpb_out[79][698],u_xpb_out[80][698],u_xpb_out[81][698],u_xpb_out[82][698],u_xpb_out[83][698],u_xpb_out[84][698],u_xpb_out[85][698],u_xpb_out[86][698],u_xpb_out[87][698],u_xpb_out[88][698],u_xpb_out[89][698],u_xpb_out[90][698],u_xpb_out[91][698],u_xpb_out[92][698],u_xpb_out[93][698],u_xpb_out[94][698],u_xpb_out[95][698],u_xpb_out[96][698],u_xpb_out[97][698],u_xpb_out[98][698],u_xpb_out[99][698],u_xpb_out[100][698],u_xpb_out[101][698],u_xpb_out[102][698],u_xpb_out[103][698],u_xpb_out[104][698],u_xpb_out[105][698]};

assign col_out_699 = {u_xpb_out[0][699],u_xpb_out[1][699],u_xpb_out[2][699],u_xpb_out[3][699],u_xpb_out[4][699],u_xpb_out[5][699],u_xpb_out[6][699],u_xpb_out[7][699],u_xpb_out[8][699],u_xpb_out[9][699],u_xpb_out[10][699],u_xpb_out[11][699],u_xpb_out[12][699],u_xpb_out[13][699],u_xpb_out[14][699],u_xpb_out[15][699],u_xpb_out[16][699],u_xpb_out[17][699],u_xpb_out[18][699],u_xpb_out[19][699],u_xpb_out[20][699],u_xpb_out[21][699],u_xpb_out[22][699],u_xpb_out[23][699],u_xpb_out[24][699],u_xpb_out[25][699],u_xpb_out[26][699],u_xpb_out[27][699],u_xpb_out[28][699],u_xpb_out[29][699],u_xpb_out[30][699],u_xpb_out[31][699],u_xpb_out[32][699],u_xpb_out[33][699],u_xpb_out[34][699],u_xpb_out[35][699],u_xpb_out[36][699],u_xpb_out[37][699],u_xpb_out[38][699],u_xpb_out[39][699],u_xpb_out[40][699],u_xpb_out[41][699],u_xpb_out[42][699],u_xpb_out[43][699],u_xpb_out[44][699],u_xpb_out[45][699],u_xpb_out[46][699],u_xpb_out[47][699],u_xpb_out[48][699],u_xpb_out[49][699],u_xpb_out[50][699],u_xpb_out[51][699],u_xpb_out[52][699],u_xpb_out[53][699],u_xpb_out[54][699],u_xpb_out[55][699],u_xpb_out[56][699],u_xpb_out[57][699],u_xpb_out[58][699],u_xpb_out[59][699],u_xpb_out[60][699],u_xpb_out[61][699],u_xpb_out[62][699],u_xpb_out[63][699],u_xpb_out[64][699],u_xpb_out[65][699],u_xpb_out[66][699],u_xpb_out[67][699],u_xpb_out[68][699],u_xpb_out[69][699],u_xpb_out[70][699],u_xpb_out[71][699],u_xpb_out[72][699],u_xpb_out[73][699],u_xpb_out[74][699],u_xpb_out[75][699],u_xpb_out[76][699],u_xpb_out[77][699],u_xpb_out[78][699],u_xpb_out[79][699],u_xpb_out[80][699],u_xpb_out[81][699],u_xpb_out[82][699],u_xpb_out[83][699],u_xpb_out[84][699],u_xpb_out[85][699],u_xpb_out[86][699],u_xpb_out[87][699],u_xpb_out[88][699],u_xpb_out[89][699],u_xpb_out[90][699],u_xpb_out[91][699],u_xpb_out[92][699],u_xpb_out[93][699],u_xpb_out[94][699],u_xpb_out[95][699],u_xpb_out[96][699],u_xpb_out[97][699],u_xpb_out[98][699],u_xpb_out[99][699],u_xpb_out[100][699],u_xpb_out[101][699],u_xpb_out[102][699],u_xpb_out[103][699],u_xpb_out[104][699],u_xpb_out[105][699]};

assign col_out_700 = {u_xpb_out[0][700],u_xpb_out[1][700],u_xpb_out[2][700],u_xpb_out[3][700],u_xpb_out[4][700],u_xpb_out[5][700],u_xpb_out[6][700],u_xpb_out[7][700],u_xpb_out[8][700],u_xpb_out[9][700],u_xpb_out[10][700],u_xpb_out[11][700],u_xpb_out[12][700],u_xpb_out[13][700],u_xpb_out[14][700],u_xpb_out[15][700],u_xpb_out[16][700],u_xpb_out[17][700],u_xpb_out[18][700],u_xpb_out[19][700],u_xpb_out[20][700],u_xpb_out[21][700],u_xpb_out[22][700],u_xpb_out[23][700],u_xpb_out[24][700],u_xpb_out[25][700],u_xpb_out[26][700],u_xpb_out[27][700],u_xpb_out[28][700],u_xpb_out[29][700],u_xpb_out[30][700],u_xpb_out[31][700],u_xpb_out[32][700],u_xpb_out[33][700],u_xpb_out[34][700],u_xpb_out[35][700],u_xpb_out[36][700],u_xpb_out[37][700],u_xpb_out[38][700],u_xpb_out[39][700],u_xpb_out[40][700],u_xpb_out[41][700],u_xpb_out[42][700],u_xpb_out[43][700],u_xpb_out[44][700],u_xpb_out[45][700],u_xpb_out[46][700],u_xpb_out[47][700],u_xpb_out[48][700],u_xpb_out[49][700],u_xpb_out[50][700],u_xpb_out[51][700],u_xpb_out[52][700],u_xpb_out[53][700],u_xpb_out[54][700],u_xpb_out[55][700],u_xpb_out[56][700],u_xpb_out[57][700],u_xpb_out[58][700],u_xpb_out[59][700],u_xpb_out[60][700],u_xpb_out[61][700],u_xpb_out[62][700],u_xpb_out[63][700],u_xpb_out[64][700],u_xpb_out[65][700],u_xpb_out[66][700],u_xpb_out[67][700],u_xpb_out[68][700],u_xpb_out[69][700],u_xpb_out[70][700],u_xpb_out[71][700],u_xpb_out[72][700],u_xpb_out[73][700],u_xpb_out[74][700],u_xpb_out[75][700],u_xpb_out[76][700],u_xpb_out[77][700],u_xpb_out[78][700],u_xpb_out[79][700],u_xpb_out[80][700],u_xpb_out[81][700],u_xpb_out[82][700],u_xpb_out[83][700],u_xpb_out[84][700],u_xpb_out[85][700],u_xpb_out[86][700],u_xpb_out[87][700],u_xpb_out[88][700],u_xpb_out[89][700],u_xpb_out[90][700],u_xpb_out[91][700],u_xpb_out[92][700],u_xpb_out[93][700],u_xpb_out[94][700],u_xpb_out[95][700],u_xpb_out[96][700],u_xpb_out[97][700],u_xpb_out[98][700],u_xpb_out[99][700],u_xpb_out[100][700],u_xpb_out[101][700],u_xpb_out[102][700],u_xpb_out[103][700],u_xpb_out[104][700],u_xpb_out[105][700]};

assign col_out_701 = {u_xpb_out[0][701],u_xpb_out[1][701],u_xpb_out[2][701],u_xpb_out[3][701],u_xpb_out[4][701],u_xpb_out[5][701],u_xpb_out[6][701],u_xpb_out[7][701],u_xpb_out[8][701],u_xpb_out[9][701],u_xpb_out[10][701],u_xpb_out[11][701],u_xpb_out[12][701],u_xpb_out[13][701],u_xpb_out[14][701],u_xpb_out[15][701],u_xpb_out[16][701],u_xpb_out[17][701],u_xpb_out[18][701],u_xpb_out[19][701],u_xpb_out[20][701],u_xpb_out[21][701],u_xpb_out[22][701],u_xpb_out[23][701],u_xpb_out[24][701],u_xpb_out[25][701],u_xpb_out[26][701],u_xpb_out[27][701],u_xpb_out[28][701],u_xpb_out[29][701],u_xpb_out[30][701],u_xpb_out[31][701],u_xpb_out[32][701],u_xpb_out[33][701],u_xpb_out[34][701],u_xpb_out[35][701],u_xpb_out[36][701],u_xpb_out[37][701],u_xpb_out[38][701],u_xpb_out[39][701],u_xpb_out[40][701],u_xpb_out[41][701],u_xpb_out[42][701],u_xpb_out[43][701],u_xpb_out[44][701],u_xpb_out[45][701],u_xpb_out[46][701],u_xpb_out[47][701],u_xpb_out[48][701],u_xpb_out[49][701],u_xpb_out[50][701],u_xpb_out[51][701],u_xpb_out[52][701],u_xpb_out[53][701],u_xpb_out[54][701],u_xpb_out[55][701],u_xpb_out[56][701],u_xpb_out[57][701],u_xpb_out[58][701],u_xpb_out[59][701],u_xpb_out[60][701],u_xpb_out[61][701],u_xpb_out[62][701],u_xpb_out[63][701],u_xpb_out[64][701],u_xpb_out[65][701],u_xpb_out[66][701],u_xpb_out[67][701],u_xpb_out[68][701],u_xpb_out[69][701],u_xpb_out[70][701],u_xpb_out[71][701],u_xpb_out[72][701],u_xpb_out[73][701],u_xpb_out[74][701],u_xpb_out[75][701],u_xpb_out[76][701],u_xpb_out[77][701],u_xpb_out[78][701],u_xpb_out[79][701],u_xpb_out[80][701],u_xpb_out[81][701],u_xpb_out[82][701],u_xpb_out[83][701],u_xpb_out[84][701],u_xpb_out[85][701],u_xpb_out[86][701],u_xpb_out[87][701],u_xpb_out[88][701],u_xpb_out[89][701],u_xpb_out[90][701],u_xpb_out[91][701],u_xpb_out[92][701],u_xpb_out[93][701],u_xpb_out[94][701],u_xpb_out[95][701],u_xpb_out[96][701],u_xpb_out[97][701],u_xpb_out[98][701],u_xpb_out[99][701],u_xpb_out[100][701],u_xpb_out[101][701],u_xpb_out[102][701],u_xpb_out[103][701],u_xpb_out[104][701],u_xpb_out[105][701]};

assign col_out_702 = {u_xpb_out[0][702],u_xpb_out[1][702],u_xpb_out[2][702],u_xpb_out[3][702],u_xpb_out[4][702],u_xpb_out[5][702],u_xpb_out[6][702],u_xpb_out[7][702],u_xpb_out[8][702],u_xpb_out[9][702],u_xpb_out[10][702],u_xpb_out[11][702],u_xpb_out[12][702],u_xpb_out[13][702],u_xpb_out[14][702],u_xpb_out[15][702],u_xpb_out[16][702],u_xpb_out[17][702],u_xpb_out[18][702],u_xpb_out[19][702],u_xpb_out[20][702],u_xpb_out[21][702],u_xpb_out[22][702],u_xpb_out[23][702],u_xpb_out[24][702],u_xpb_out[25][702],u_xpb_out[26][702],u_xpb_out[27][702],u_xpb_out[28][702],u_xpb_out[29][702],u_xpb_out[30][702],u_xpb_out[31][702],u_xpb_out[32][702],u_xpb_out[33][702],u_xpb_out[34][702],u_xpb_out[35][702],u_xpb_out[36][702],u_xpb_out[37][702],u_xpb_out[38][702],u_xpb_out[39][702],u_xpb_out[40][702],u_xpb_out[41][702],u_xpb_out[42][702],u_xpb_out[43][702],u_xpb_out[44][702],u_xpb_out[45][702],u_xpb_out[46][702],u_xpb_out[47][702],u_xpb_out[48][702],u_xpb_out[49][702],u_xpb_out[50][702],u_xpb_out[51][702],u_xpb_out[52][702],u_xpb_out[53][702],u_xpb_out[54][702],u_xpb_out[55][702],u_xpb_out[56][702],u_xpb_out[57][702],u_xpb_out[58][702],u_xpb_out[59][702],u_xpb_out[60][702],u_xpb_out[61][702],u_xpb_out[62][702],u_xpb_out[63][702],u_xpb_out[64][702],u_xpb_out[65][702],u_xpb_out[66][702],u_xpb_out[67][702],u_xpb_out[68][702],u_xpb_out[69][702],u_xpb_out[70][702],u_xpb_out[71][702],u_xpb_out[72][702],u_xpb_out[73][702],u_xpb_out[74][702],u_xpb_out[75][702],u_xpb_out[76][702],u_xpb_out[77][702],u_xpb_out[78][702],u_xpb_out[79][702],u_xpb_out[80][702],u_xpb_out[81][702],u_xpb_out[82][702],u_xpb_out[83][702],u_xpb_out[84][702],u_xpb_out[85][702],u_xpb_out[86][702],u_xpb_out[87][702],u_xpb_out[88][702],u_xpb_out[89][702],u_xpb_out[90][702],u_xpb_out[91][702],u_xpb_out[92][702],u_xpb_out[93][702],u_xpb_out[94][702],u_xpb_out[95][702],u_xpb_out[96][702],u_xpb_out[97][702],u_xpb_out[98][702],u_xpb_out[99][702],u_xpb_out[100][702],u_xpb_out[101][702],u_xpb_out[102][702],u_xpb_out[103][702],u_xpb_out[104][702],u_xpb_out[105][702]};

assign col_out_703 = {u_xpb_out[0][703],u_xpb_out[1][703],u_xpb_out[2][703],u_xpb_out[3][703],u_xpb_out[4][703],u_xpb_out[5][703],u_xpb_out[6][703],u_xpb_out[7][703],u_xpb_out[8][703],u_xpb_out[9][703],u_xpb_out[10][703],u_xpb_out[11][703],u_xpb_out[12][703],u_xpb_out[13][703],u_xpb_out[14][703],u_xpb_out[15][703],u_xpb_out[16][703],u_xpb_out[17][703],u_xpb_out[18][703],u_xpb_out[19][703],u_xpb_out[20][703],u_xpb_out[21][703],u_xpb_out[22][703],u_xpb_out[23][703],u_xpb_out[24][703],u_xpb_out[25][703],u_xpb_out[26][703],u_xpb_out[27][703],u_xpb_out[28][703],u_xpb_out[29][703],u_xpb_out[30][703],u_xpb_out[31][703],u_xpb_out[32][703],u_xpb_out[33][703],u_xpb_out[34][703],u_xpb_out[35][703],u_xpb_out[36][703],u_xpb_out[37][703],u_xpb_out[38][703],u_xpb_out[39][703],u_xpb_out[40][703],u_xpb_out[41][703],u_xpb_out[42][703],u_xpb_out[43][703],u_xpb_out[44][703],u_xpb_out[45][703],u_xpb_out[46][703],u_xpb_out[47][703],u_xpb_out[48][703],u_xpb_out[49][703],u_xpb_out[50][703],u_xpb_out[51][703],u_xpb_out[52][703],u_xpb_out[53][703],u_xpb_out[54][703],u_xpb_out[55][703],u_xpb_out[56][703],u_xpb_out[57][703],u_xpb_out[58][703],u_xpb_out[59][703],u_xpb_out[60][703],u_xpb_out[61][703],u_xpb_out[62][703],u_xpb_out[63][703],u_xpb_out[64][703],u_xpb_out[65][703],u_xpb_out[66][703],u_xpb_out[67][703],u_xpb_out[68][703],u_xpb_out[69][703],u_xpb_out[70][703],u_xpb_out[71][703],u_xpb_out[72][703],u_xpb_out[73][703],u_xpb_out[74][703],u_xpb_out[75][703],u_xpb_out[76][703],u_xpb_out[77][703],u_xpb_out[78][703],u_xpb_out[79][703],u_xpb_out[80][703],u_xpb_out[81][703],u_xpb_out[82][703],u_xpb_out[83][703],u_xpb_out[84][703],u_xpb_out[85][703],u_xpb_out[86][703],u_xpb_out[87][703],u_xpb_out[88][703],u_xpb_out[89][703],u_xpb_out[90][703],u_xpb_out[91][703],u_xpb_out[92][703],u_xpb_out[93][703],u_xpb_out[94][703],u_xpb_out[95][703],u_xpb_out[96][703],u_xpb_out[97][703],u_xpb_out[98][703],u_xpb_out[99][703],u_xpb_out[100][703],u_xpb_out[101][703],u_xpb_out[102][703],u_xpb_out[103][703],u_xpb_out[104][703],u_xpb_out[105][703]};

assign col_out_704 = {u_xpb_out[0][704],u_xpb_out[1][704],u_xpb_out[2][704],u_xpb_out[3][704],u_xpb_out[4][704],u_xpb_out[5][704],u_xpb_out[6][704],u_xpb_out[7][704],u_xpb_out[8][704],u_xpb_out[9][704],u_xpb_out[10][704],u_xpb_out[11][704],u_xpb_out[12][704],u_xpb_out[13][704],u_xpb_out[14][704],u_xpb_out[15][704],u_xpb_out[16][704],u_xpb_out[17][704],u_xpb_out[18][704],u_xpb_out[19][704],u_xpb_out[20][704],u_xpb_out[21][704],u_xpb_out[22][704],u_xpb_out[23][704],u_xpb_out[24][704],u_xpb_out[25][704],u_xpb_out[26][704],u_xpb_out[27][704],u_xpb_out[28][704],u_xpb_out[29][704],u_xpb_out[30][704],u_xpb_out[31][704],u_xpb_out[32][704],u_xpb_out[33][704],u_xpb_out[34][704],u_xpb_out[35][704],u_xpb_out[36][704],u_xpb_out[37][704],u_xpb_out[38][704],u_xpb_out[39][704],u_xpb_out[40][704],u_xpb_out[41][704],u_xpb_out[42][704],u_xpb_out[43][704],u_xpb_out[44][704],u_xpb_out[45][704],u_xpb_out[46][704],u_xpb_out[47][704],u_xpb_out[48][704],u_xpb_out[49][704],u_xpb_out[50][704],u_xpb_out[51][704],u_xpb_out[52][704],u_xpb_out[53][704],u_xpb_out[54][704],u_xpb_out[55][704],u_xpb_out[56][704],u_xpb_out[57][704],u_xpb_out[58][704],u_xpb_out[59][704],u_xpb_out[60][704],u_xpb_out[61][704],u_xpb_out[62][704],u_xpb_out[63][704],u_xpb_out[64][704],u_xpb_out[65][704],u_xpb_out[66][704],u_xpb_out[67][704],u_xpb_out[68][704],u_xpb_out[69][704],u_xpb_out[70][704],u_xpb_out[71][704],u_xpb_out[72][704],u_xpb_out[73][704],u_xpb_out[74][704],u_xpb_out[75][704],u_xpb_out[76][704],u_xpb_out[77][704],u_xpb_out[78][704],u_xpb_out[79][704],u_xpb_out[80][704],u_xpb_out[81][704],u_xpb_out[82][704],u_xpb_out[83][704],u_xpb_out[84][704],u_xpb_out[85][704],u_xpb_out[86][704],u_xpb_out[87][704],u_xpb_out[88][704],u_xpb_out[89][704],u_xpb_out[90][704],u_xpb_out[91][704],u_xpb_out[92][704],u_xpb_out[93][704],u_xpb_out[94][704],u_xpb_out[95][704],u_xpb_out[96][704],u_xpb_out[97][704],u_xpb_out[98][704],u_xpb_out[99][704],u_xpb_out[100][704],u_xpb_out[101][704],u_xpb_out[102][704],u_xpb_out[103][704],u_xpb_out[104][704],u_xpb_out[105][704]};

assign col_out_705 = {u_xpb_out[0][705],u_xpb_out[1][705],u_xpb_out[2][705],u_xpb_out[3][705],u_xpb_out[4][705],u_xpb_out[5][705],u_xpb_out[6][705],u_xpb_out[7][705],u_xpb_out[8][705],u_xpb_out[9][705],u_xpb_out[10][705],u_xpb_out[11][705],u_xpb_out[12][705],u_xpb_out[13][705],u_xpb_out[14][705],u_xpb_out[15][705],u_xpb_out[16][705],u_xpb_out[17][705],u_xpb_out[18][705],u_xpb_out[19][705],u_xpb_out[20][705],u_xpb_out[21][705],u_xpb_out[22][705],u_xpb_out[23][705],u_xpb_out[24][705],u_xpb_out[25][705],u_xpb_out[26][705],u_xpb_out[27][705],u_xpb_out[28][705],u_xpb_out[29][705],u_xpb_out[30][705],u_xpb_out[31][705],u_xpb_out[32][705],u_xpb_out[33][705],u_xpb_out[34][705],u_xpb_out[35][705],u_xpb_out[36][705],u_xpb_out[37][705],u_xpb_out[38][705],u_xpb_out[39][705],u_xpb_out[40][705],u_xpb_out[41][705],u_xpb_out[42][705],u_xpb_out[43][705],u_xpb_out[44][705],u_xpb_out[45][705],u_xpb_out[46][705],u_xpb_out[47][705],u_xpb_out[48][705],u_xpb_out[49][705],u_xpb_out[50][705],u_xpb_out[51][705],u_xpb_out[52][705],u_xpb_out[53][705],u_xpb_out[54][705],u_xpb_out[55][705],u_xpb_out[56][705],u_xpb_out[57][705],u_xpb_out[58][705],u_xpb_out[59][705],u_xpb_out[60][705],u_xpb_out[61][705],u_xpb_out[62][705],u_xpb_out[63][705],u_xpb_out[64][705],u_xpb_out[65][705],u_xpb_out[66][705],u_xpb_out[67][705],u_xpb_out[68][705],u_xpb_out[69][705],u_xpb_out[70][705],u_xpb_out[71][705],u_xpb_out[72][705],u_xpb_out[73][705],u_xpb_out[74][705],u_xpb_out[75][705],u_xpb_out[76][705],u_xpb_out[77][705],u_xpb_out[78][705],u_xpb_out[79][705],u_xpb_out[80][705],u_xpb_out[81][705],u_xpb_out[82][705],u_xpb_out[83][705],u_xpb_out[84][705],u_xpb_out[85][705],u_xpb_out[86][705],u_xpb_out[87][705],u_xpb_out[88][705],u_xpb_out[89][705],u_xpb_out[90][705],u_xpb_out[91][705],u_xpb_out[92][705],u_xpb_out[93][705],u_xpb_out[94][705],u_xpb_out[95][705],u_xpb_out[96][705],u_xpb_out[97][705],u_xpb_out[98][705],u_xpb_out[99][705],u_xpb_out[100][705],u_xpb_out[101][705],u_xpb_out[102][705],u_xpb_out[103][705],u_xpb_out[104][705],u_xpb_out[105][705]};

assign col_out_706 = {u_xpb_out[0][706],u_xpb_out[1][706],u_xpb_out[2][706],u_xpb_out[3][706],u_xpb_out[4][706],u_xpb_out[5][706],u_xpb_out[6][706],u_xpb_out[7][706],u_xpb_out[8][706],u_xpb_out[9][706],u_xpb_out[10][706],u_xpb_out[11][706],u_xpb_out[12][706],u_xpb_out[13][706],u_xpb_out[14][706],u_xpb_out[15][706],u_xpb_out[16][706],u_xpb_out[17][706],u_xpb_out[18][706],u_xpb_out[19][706],u_xpb_out[20][706],u_xpb_out[21][706],u_xpb_out[22][706],u_xpb_out[23][706],u_xpb_out[24][706],u_xpb_out[25][706],u_xpb_out[26][706],u_xpb_out[27][706],u_xpb_out[28][706],u_xpb_out[29][706],u_xpb_out[30][706],u_xpb_out[31][706],u_xpb_out[32][706],u_xpb_out[33][706],u_xpb_out[34][706],u_xpb_out[35][706],u_xpb_out[36][706],u_xpb_out[37][706],u_xpb_out[38][706],u_xpb_out[39][706],u_xpb_out[40][706],u_xpb_out[41][706],u_xpb_out[42][706],u_xpb_out[43][706],u_xpb_out[44][706],u_xpb_out[45][706],u_xpb_out[46][706],u_xpb_out[47][706],u_xpb_out[48][706],u_xpb_out[49][706],u_xpb_out[50][706],u_xpb_out[51][706],u_xpb_out[52][706],u_xpb_out[53][706],u_xpb_out[54][706],u_xpb_out[55][706],u_xpb_out[56][706],u_xpb_out[57][706],u_xpb_out[58][706],u_xpb_out[59][706],u_xpb_out[60][706],u_xpb_out[61][706],u_xpb_out[62][706],u_xpb_out[63][706],u_xpb_out[64][706],u_xpb_out[65][706],u_xpb_out[66][706],u_xpb_out[67][706],u_xpb_out[68][706],u_xpb_out[69][706],u_xpb_out[70][706],u_xpb_out[71][706],u_xpb_out[72][706],u_xpb_out[73][706],u_xpb_out[74][706],u_xpb_out[75][706],u_xpb_out[76][706],u_xpb_out[77][706],u_xpb_out[78][706],u_xpb_out[79][706],u_xpb_out[80][706],u_xpb_out[81][706],u_xpb_out[82][706],u_xpb_out[83][706],u_xpb_out[84][706],u_xpb_out[85][706],u_xpb_out[86][706],u_xpb_out[87][706],u_xpb_out[88][706],u_xpb_out[89][706],u_xpb_out[90][706],u_xpb_out[91][706],u_xpb_out[92][706],u_xpb_out[93][706],u_xpb_out[94][706],u_xpb_out[95][706],u_xpb_out[96][706],u_xpb_out[97][706],u_xpb_out[98][706],u_xpb_out[99][706],u_xpb_out[100][706],u_xpb_out[101][706],u_xpb_out[102][706],u_xpb_out[103][706],u_xpb_out[104][706],u_xpb_out[105][706]};

assign col_out_707 = {u_xpb_out[0][707],u_xpb_out[1][707],u_xpb_out[2][707],u_xpb_out[3][707],u_xpb_out[4][707],u_xpb_out[5][707],u_xpb_out[6][707],u_xpb_out[7][707],u_xpb_out[8][707],u_xpb_out[9][707],u_xpb_out[10][707],u_xpb_out[11][707],u_xpb_out[12][707],u_xpb_out[13][707],u_xpb_out[14][707],u_xpb_out[15][707],u_xpb_out[16][707],u_xpb_out[17][707],u_xpb_out[18][707],u_xpb_out[19][707],u_xpb_out[20][707],u_xpb_out[21][707],u_xpb_out[22][707],u_xpb_out[23][707],u_xpb_out[24][707],u_xpb_out[25][707],u_xpb_out[26][707],u_xpb_out[27][707],u_xpb_out[28][707],u_xpb_out[29][707],u_xpb_out[30][707],u_xpb_out[31][707],u_xpb_out[32][707],u_xpb_out[33][707],u_xpb_out[34][707],u_xpb_out[35][707],u_xpb_out[36][707],u_xpb_out[37][707],u_xpb_out[38][707],u_xpb_out[39][707],u_xpb_out[40][707],u_xpb_out[41][707],u_xpb_out[42][707],u_xpb_out[43][707],u_xpb_out[44][707],u_xpb_out[45][707],u_xpb_out[46][707],u_xpb_out[47][707],u_xpb_out[48][707],u_xpb_out[49][707],u_xpb_out[50][707],u_xpb_out[51][707],u_xpb_out[52][707],u_xpb_out[53][707],u_xpb_out[54][707],u_xpb_out[55][707],u_xpb_out[56][707],u_xpb_out[57][707],u_xpb_out[58][707],u_xpb_out[59][707],u_xpb_out[60][707],u_xpb_out[61][707],u_xpb_out[62][707],u_xpb_out[63][707],u_xpb_out[64][707],u_xpb_out[65][707],u_xpb_out[66][707],u_xpb_out[67][707],u_xpb_out[68][707],u_xpb_out[69][707],u_xpb_out[70][707],u_xpb_out[71][707],u_xpb_out[72][707],u_xpb_out[73][707],u_xpb_out[74][707],u_xpb_out[75][707],u_xpb_out[76][707],u_xpb_out[77][707],u_xpb_out[78][707],u_xpb_out[79][707],u_xpb_out[80][707],u_xpb_out[81][707],u_xpb_out[82][707],u_xpb_out[83][707],u_xpb_out[84][707],u_xpb_out[85][707],u_xpb_out[86][707],u_xpb_out[87][707],u_xpb_out[88][707],u_xpb_out[89][707],u_xpb_out[90][707],u_xpb_out[91][707],u_xpb_out[92][707],u_xpb_out[93][707],u_xpb_out[94][707],u_xpb_out[95][707],u_xpb_out[96][707],u_xpb_out[97][707],u_xpb_out[98][707],u_xpb_out[99][707],u_xpb_out[100][707],u_xpb_out[101][707],u_xpb_out[102][707],u_xpb_out[103][707],u_xpb_out[104][707],u_xpb_out[105][707]};

assign col_out_708 = {u_xpb_out[0][708],u_xpb_out[1][708],u_xpb_out[2][708],u_xpb_out[3][708],u_xpb_out[4][708],u_xpb_out[5][708],u_xpb_out[6][708],u_xpb_out[7][708],u_xpb_out[8][708],u_xpb_out[9][708],u_xpb_out[10][708],u_xpb_out[11][708],u_xpb_out[12][708],u_xpb_out[13][708],u_xpb_out[14][708],u_xpb_out[15][708],u_xpb_out[16][708],u_xpb_out[17][708],u_xpb_out[18][708],u_xpb_out[19][708],u_xpb_out[20][708],u_xpb_out[21][708],u_xpb_out[22][708],u_xpb_out[23][708],u_xpb_out[24][708],u_xpb_out[25][708],u_xpb_out[26][708],u_xpb_out[27][708],u_xpb_out[28][708],u_xpb_out[29][708],u_xpb_out[30][708],u_xpb_out[31][708],u_xpb_out[32][708],u_xpb_out[33][708],u_xpb_out[34][708],u_xpb_out[35][708],u_xpb_out[36][708],u_xpb_out[37][708],u_xpb_out[38][708],u_xpb_out[39][708],u_xpb_out[40][708],u_xpb_out[41][708],u_xpb_out[42][708],u_xpb_out[43][708],u_xpb_out[44][708],u_xpb_out[45][708],u_xpb_out[46][708],u_xpb_out[47][708],u_xpb_out[48][708],u_xpb_out[49][708],u_xpb_out[50][708],u_xpb_out[51][708],u_xpb_out[52][708],u_xpb_out[53][708],u_xpb_out[54][708],u_xpb_out[55][708],u_xpb_out[56][708],u_xpb_out[57][708],u_xpb_out[58][708],u_xpb_out[59][708],u_xpb_out[60][708],u_xpb_out[61][708],u_xpb_out[62][708],u_xpb_out[63][708],u_xpb_out[64][708],u_xpb_out[65][708],u_xpb_out[66][708],u_xpb_out[67][708],u_xpb_out[68][708],u_xpb_out[69][708],u_xpb_out[70][708],u_xpb_out[71][708],u_xpb_out[72][708],u_xpb_out[73][708],u_xpb_out[74][708],u_xpb_out[75][708],u_xpb_out[76][708],u_xpb_out[77][708],u_xpb_out[78][708],u_xpb_out[79][708],u_xpb_out[80][708],u_xpb_out[81][708],u_xpb_out[82][708],u_xpb_out[83][708],u_xpb_out[84][708],u_xpb_out[85][708],u_xpb_out[86][708],u_xpb_out[87][708],u_xpb_out[88][708],u_xpb_out[89][708],u_xpb_out[90][708],u_xpb_out[91][708],u_xpb_out[92][708],u_xpb_out[93][708],u_xpb_out[94][708],u_xpb_out[95][708],u_xpb_out[96][708],u_xpb_out[97][708],u_xpb_out[98][708],u_xpb_out[99][708],u_xpb_out[100][708],u_xpb_out[101][708],u_xpb_out[102][708],u_xpb_out[103][708],u_xpb_out[104][708],u_xpb_out[105][708]};

assign col_out_709 = {u_xpb_out[0][709],u_xpb_out[1][709],u_xpb_out[2][709],u_xpb_out[3][709],u_xpb_out[4][709],u_xpb_out[5][709],u_xpb_out[6][709],u_xpb_out[7][709],u_xpb_out[8][709],u_xpb_out[9][709],u_xpb_out[10][709],u_xpb_out[11][709],u_xpb_out[12][709],u_xpb_out[13][709],u_xpb_out[14][709],u_xpb_out[15][709],u_xpb_out[16][709],u_xpb_out[17][709],u_xpb_out[18][709],u_xpb_out[19][709],u_xpb_out[20][709],u_xpb_out[21][709],u_xpb_out[22][709],u_xpb_out[23][709],u_xpb_out[24][709],u_xpb_out[25][709],u_xpb_out[26][709],u_xpb_out[27][709],u_xpb_out[28][709],u_xpb_out[29][709],u_xpb_out[30][709],u_xpb_out[31][709],u_xpb_out[32][709],u_xpb_out[33][709],u_xpb_out[34][709],u_xpb_out[35][709],u_xpb_out[36][709],u_xpb_out[37][709],u_xpb_out[38][709],u_xpb_out[39][709],u_xpb_out[40][709],u_xpb_out[41][709],u_xpb_out[42][709],u_xpb_out[43][709],u_xpb_out[44][709],u_xpb_out[45][709],u_xpb_out[46][709],u_xpb_out[47][709],u_xpb_out[48][709],u_xpb_out[49][709],u_xpb_out[50][709],u_xpb_out[51][709],u_xpb_out[52][709],u_xpb_out[53][709],u_xpb_out[54][709],u_xpb_out[55][709],u_xpb_out[56][709],u_xpb_out[57][709],u_xpb_out[58][709],u_xpb_out[59][709],u_xpb_out[60][709],u_xpb_out[61][709],u_xpb_out[62][709],u_xpb_out[63][709],u_xpb_out[64][709],u_xpb_out[65][709],u_xpb_out[66][709],u_xpb_out[67][709],u_xpb_out[68][709],u_xpb_out[69][709],u_xpb_out[70][709],u_xpb_out[71][709],u_xpb_out[72][709],u_xpb_out[73][709],u_xpb_out[74][709],u_xpb_out[75][709],u_xpb_out[76][709],u_xpb_out[77][709],u_xpb_out[78][709],u_xpb_out[79][709],u_xpb_out[80][709],u_xpb_out[81][709],u_xpb_out[82][709],u_xpb_out[83][709],u_xpb_out[84][709],u_xpb_out[85][709],u_xpb_out[86][709],u_xpb_out[87][709],u_xpb_out[88][709],u_xpb_out[89][709],u_xpb_out[90][709],u_xpb_out[91][709],u_xpb_out[92][709],u_xpb_out[93][709],u_xpb_out[94][709],u_xpb_out[95][709],u_xpb_out[96][709],u_xpb_out[97][709],u_xpb_out[98][709],u_xpb_out[99][709],u_xpb_out[100][709],u_xpb_out[101][709],u_xpb_out[102][709],u_xpb_out[103][709],u_xpb_out[104][709],u_xpb_out[105][709]};

assign col_out_710 = {u_xpb_out[0][710],u_xpb_out[1][710],u_xpb_out[2][710],u_xpb_out[3][710],u_xpb_out[4][710],u_xpb_out[5][710],u_xpb_out[6][710],u_xpb_out[7][710],u_xpb_out[8][710],u_xpb_out[9][710],u_xpb_out[10][710],u_xpb_out[11][710],u_xpb_out[12][710],u_xpb_out[13][710],u_xpb_out[14][710],u_xpb_out[15][710],u_xpb_out[16][710],u_xpb_out[17][710],u_xpb_out[18][710],u_xpb_out[19][710],u_xpb_out[20][710],u_xpb_out[21][710],u_xpb_out[22][710],u_xpb_out[23][710],u_xpb_out[24][710],u_xpb_out[25][710],u_xpb_out[26][710],u_xpb_out[27][710],u_xpb_out[28][710],u_xpb_out[29][710],u_xpb_out[30][710],u_xpb_out[31][710],u_xpb_out[32][710],u_xpb_out[33][710],u_xpb_out[34][710],u_xpb_out[35][710],u_xpb_out[36][710],u_xpb_out[37][710],u_xpb_out[38][710],u_xpb_out[39][710],u_xpb_out[40][710],u_xpb_out[41][710],u_xpb_out[42][710],u_xpb_out[43][710],u_xpb_out[44][710],u_xpb_out[45][710],u_xpb_out[46][710],u_xpb_out[47][710],u_xpb_out[48][710],u_xpb_out[49][710],u_xpb_out[50][710],u_xpb_out[51][710],u_xpb_out[52][710],u_xpb_out[53][710],u_xpb_out[54][710],u_xpb_out[55][710],u_xpb_out[56][710],u_xpb_out[57][710],u_xpb_out[58][710],u_xpb_out[59][710],u_xpb_out[60][710],u_xpb_out[61][710],u_xpb_out[62][710],u_xpb_out[63][710],u_xpb_out[64][710],u_xpb_out[65][710],u_xpb_out[66][710],u_xpb_out[67][710],u_xpb_out[68][710],u_xpb_out[69][710],u_xpb_out[70][710],u_xpb_out[71][710],u_xpb_out[72][710],u_xpb_out[73][710],u_xpb_out[74][710],u_xpb_out[75][710],u_xpb_out[76][710],u_xpb_out[77][710],u_xpb_out[78][710],u_xpb_out[79][710],u_xpb_out[80][710],u_xpb_out[81][710],u_xpb_out[82][710],u_xpb_out[83][710],u_xpb_out[84][710],u_xpb_out[85][710],u_xpb_out[86][710],u_xpb_out[87][710],u_xpb_out[88][710],u_xpb_out[89][710],u_xpb_out[90][710],u_xpb_out[91][710],u_xpb_out[92][710],u_xpb_out[93][710],u_xpb_out[94][710],u_xpb_out[95][710],u_xpb_out[96][710],u_xpb_out[97][710],u_xpb_out[98][710],u_xpb_out[99][710],u_xpb_out[100][710],u_xpb_out[101][710],u_xpb_out[102][710],u_xpb_out[103][710],u_xpb_out[104][710],u_xpb_out[105][710]};

assign col_out_711 = {u_xpb_out[0][711],u_xpb_out[1][711],u_xpb_out[2][711],u_xpb_out[3][711],u_xpb_out[4][711],u_xpb_out[5][711],u_xpb_out[6][711],u_xpb_out[7][711],u_xpb_out[8][711],u_xpb_out[9][711],u_xpb_out[10][711],u_xpb_out[11][711],u_xpb_out[12][711],u_xpb_out[13][711],u_xpb_out[14][711],u_xpb_out[15][711],u_xpb_out[16][711],u_xpb_out[17][711],u_xpb_out[18][711],u_xpb_out[19][711],u_xpb_out[20][711],u_xpb_out[21][711],u_xpb_out[22][711],u_xpb_out[23][711],u_xpb_out[24][711],u_xpb_out[25][711],u_xpb_out[26][711],u_xpb_out[27][711],u_xpb_out[28][711],u_xpb_out[29][711],u_xpb_out[30][711],u_xpb_out[31][711],u_xpb_out[32][711],u_xpb_out[33][711],u_xpb_out[34][711],u_xpb_out[35][711],u_xpb_out[36][711],u_xpb_out[37][711],u_xpb_out[38][711],u_xpb_out[39][711],u_xpb_out[40][711],u_xpb_out[41][711],u_xpb_out[42][711],u_xpb_out[43][711],u_xpb_out[44][711],u_xpb_out[45][711],u_xpb_out[46][711],u_xpb_out[47][711],u_xpb_out[48][711],u_xpb_out[49][711],u_xpb_out[50][711],u_xpb_out[51][711],u_xpb_out[52][711],u_xpb_out[53][711],u_xpb_out[54][711],u_xpb_out[55][711],u_xpb_out[56][711],u_xpb_out[57][711],u_xpb_out[58][711],u_xpb_out[59][711],u_xpb_out[60][711],u_xpb_out[61][711],u_xpb_out[62][711],u_xpb_out[63][711],u_xpb_out[64][711],u_xpb_out[65][711],u_xpb_out[66][711],u_xpb_out[67][711],u_xpb_out[68][711],u_xpb_out[69][711],u_xpb_out[70][711],u_xpb_out[71][711],u_xpb_out[72][711],u_xpb_out[73][711],u_xpb_out[74][711],u_xpb_out[75][711],u_xpb_out[76][711],u_xpb_out[77][711],u_xpb_out[78][711],u_xpb_out[79][711],u_xpb_out[80][711],u_xpb_out[81][711],u_xpb_out[82][711],u_xpb_out[83][711],u_xpb_out[84][711],u_xpb_out[85][711],u_xpb_out[86][711],u_xpb_out[87][711],u_xpb_out[88][711],u_xpb_out[89][711],u_xpb_out[90][711],u_xpb_out[91][711],u_xpb_out[92][711],u_xpb_out[93][711],u_xpb_out[94][711],u_xpb_out[95][711],u_xpb_out[96][711],u_xpb_out[97][711],u_xpb_out[98][711],u_xpb_out[99][711],u_xpb_out[100][711],u_xpb_out[101][711],u_xpb_out[102][711],u_xpb_out[103][711],u_xpb_out[104][711],u_xpb_out[105][711]};

assign col_out_712 = {u_xpb_out[0][712],u_xpb_out[1][712],u_xpb_out[2][712],u_xpb_out[3][712],u_xpb_out[4][712],u_xpb_out[5][712],u_xpb_out[6][712],u_xpb_out[7][712],u_xpb_out[8][712],u_xpb_out[9][712],u_xpb_out[10][712],u_xpb_out[11][712],u_xpb_out[12][712],u_xpb_out[13][712],u_xpb_out[14][712],u_xpb_out[15][712],u_xpb_out[16][712],u_xpb_out[17][712],u_xpb_out[18][712],u_xpb_out[19][712],u_xpb_out[20][712],u_xpb_out[21][712],u_xpb_out[22][712],u_xpb_out[23][712],u_xpb_out[24][712],u_xpb_out[25][712],u_xpb_out[26][712],u_xpb_out[27][712],u_xpb_out[28][712],u_xpb_out[29][712],u_xpb_out[30][712],u_xpb_out[31][712],u_xpb_out[32][712],u_xpb_out[33][712],u_xpb_out[34][712],u_xpb_out[35][712],u_xpb_out[36][712],u_xpb_out[37][712],u_xpb_out[38][712],u_xpb_out[39][712],u_xpb_out[40][712],u_xpb_out[41][712],u_xpb_out[42][712],u_xpb_out[43][712],u_xpb_out[44][712],u_xpb_out[45][712],u_xpb_out[46][712],u_xpb_out[47][712],u_xpb_out[48][712],u_xpb_out[49][712],u_xpb_out[50][712],u_xpb_out[51][712],u_xpb_out[52][712],u_xpb_out[53][712],u_xpb_out[54][712],u_xpb_out[55][712],u_xpb_out[56][712],u_xpb_out[57][712],u_xpb_out[58][712],u_xpb_out[59][712],u_xpb_out[60][712],u_xpb_out[61][712],u_xpb_out[62][712],u_xpb_out[63][712],u_xpb_out[64][712],u_xpb_out[65][712],u_xpb_out[66][712],u_xpb_out[67][712],u_xpb_out[68][712],u_xpb_out[69][712],u_xpb_out[70][712],u_xpb_out[71][712],u_xpb_out[72][712],u_xpb_out[73][712],u_xpb_out[74][712],u_xpb_out[75][712],u_xpb_out[76][712],u_xpb_out[77][712],u_xpb_out[78][712],u_xpb_out[79][712],u_xpb_out[80][712],u_xpb_out[81][712],u_xpb_out[82][712],u_xpb_out[83][712],u_xpb_out[84][712],u_xpb_out[85][712],u_xpb_out[86][712],u_xpb_out[87][712],u_xpb_out[88][712],u_xpb_out[89][712],u_xpb_out[90][712],u_xpb_out[91][712],u_xpb_out[92][712],u_xpb_out[93][712],u_xpb_out[94][712],u_xpb_out[95][712],u_xpb_out[96][712],u_xpb_out[97][712],u_xpb_out[98][712],u_xpb_out[99][712],u_xpb_out[100][712],u_xpb_out[101][712],u_xpb_out[102][712],u_xpb_out[103][712],u_xpb_out[104][712],u_xpb_out[105][712]};

assign col_out_713 = {u_xpb_out[0][713],u_xpb_out[1][713],u_xpb_out[2][713],u_xpb_out[3][713],u_xpb_out[4][713],u_xpb_out[5][713],u_xpb_out[6][713],u_xpb_out[7][713],u_xpb_out[8][713],u_xpb_out[9][713],u_xpb_out[10][713],u_xpb_out[11][713],u_xpb_out[12][713],u_xpb_out[13][713],u_xpb_out[14][713],u_xpb_out[15][713],u_xpb_out[16][713],u_xpb_out[17][713],u_xpb_out[18][713],u_xpb_out[19][713],u_xpb_out[20][713],u_xpb_out[21][713],u_xpb_out[22][713],u_xpb_out[23][713],u_xpb_out[24][713],u_xpb_out[25][713],u_xpb_out[26][713],u_xpb_out[27][713],u_xpb_out[28][713],u_xpb_out[29][713],u_xpb_out[30][713],u_xpb_out[31][713],u_xpb_out[32][713],u_xpb_out[33][713],u_xpb_out[34][713],u_xpb_out[35][713],u_xpb_out[36][713],u_xpb_out[37][713],u_xpb_out[38][713],u_xpb_out[39][713],u_xpb_out[40][713],u_xpb_out[41][713],u_xpb_out[42][713],u_xpb_out[43][713],u_xpb_out[44][713],u_xpb_out[45][713],u_xpb_out[46][713],u_xpb_out[47][713],u_xpb_out[48][713],u_xpb_out[49][713],u_xpb_out[50][713],u_xpb_out[51][713],u_xpb_out[52][713],u_xpb_out[53][713],u_xpb_out[54][713],u_xpb_out[55][713],u_xpb_out[56][713],u_xpb_out[57][713],u_xpb_out[58][713],u_xpb_out[59][713],u_xpb_out[60][713],u_xpb_out[61][713],u_xpb_out[62][713],u_xpb_out[63][713],u_xpb_out[64][713],u_xpb_out[65][713],u_xpb_out[66][713],u_xpb_out[67][713],u_xpb_out[68][713],u_xpb_out[69][713],u_xpb_out[70][713],u_xpb_out[71][713],u_xpb_out[72][713],u_xpb_out[73][713],u_xpb_out[74][713],u_xpb_out[75][713],u_xpb_out[76][713],u_xpb_out[77][713],u_xpb_out[78][713],u_xpb_out[79][713],u_xpb_out[80][713],u_xpb_out[81][713],u_xpb_out[82][713],u_xpb_out[83][713],u_xpb_out[84][713],u_xpb_out[85][713],u_xpb_out[86][713],u_xpb_out[87][713],u_xpb_out[88][713],u_xpb_out[89][713],u_xpb_out[90][713],u_xpb_out[91][713],u_xpb_out[92][713],u_xpb_out[93][713],u_xpb_out[94][713],u_xpb_out[95][713],u_xpb_out[96][713],u_xpb_out[97][713],u_xpb_out[98][713],u_xpb_out[99][713],u_xpb_out[100][713],u_xpb_out[101][713],u_xpb_out[102][713],u_xpb_out[103][713],u_xpb_out[104][713],u_xpb_out[105][713]};

assign col_out_714 = {u_xpb_out[0][714],u_xpb_out[1][714],u_xpb_out[2][714],u_xpb_out[3][714],u_xpb_out[4][714],u_xpb_out[5][714],u_xpb_out[6][714],u_xpb_out[7][714],u_xpb_out[8][714],u_xpb_out[9][714],u_xpb_out[10][714],u_xpb_out[11][714],u_xpb_out[12][714],u_xpb_out[13][714],u_xpb_out[14][714],u_xpb_out[15][714],u_xpb_out[16][714],u_xpb_out[17][714],u_xpb_out[18][714],u_xpb_out[19][714],u_xpb_out[20][714],u_xpb_out[21][714],u_xpb_out[22][714],u_xpb_out[23][714],u_xpb_out[24][714],u_xpb_out[25][714],u_xpb_out[26][714],u_xpb_out[27][714],u_xpb_out[28][714],u_xpb_out[29][714],u_xpb_out[30][714],u_xpb_out[31][714],u_xpb_out[32][714],u_xpb_out[33][714],u_xpb_out[34][714],u_xpb_out[35][714],u_xpb_out[36][714],u_xpb_out[37][714],u_xpb_out[38][714],u_xpb_out[39][714],u_xpb_out[40][714],u_xpb_out[41][714],u_xpb_out[42][714],u_xpb_out[43][714],u_xpb_out[44][714],u_xpb_out[45][714],u_xpb_out[46][714],u_xpb_out[47][714],u_xpb_out[48][714],u_xpb_out[49][714],u_xpb_out[50][714],u_xpb_out[51][714],u_xpb_out[52][714],u_xpb_out[53][714],u_xpb_out[54][714],u_xpb_out[55][714],u_xpb_out[56][714],u_xpb_out[57][714],u_xpb_out[58][714],u_xpb_out[59][714],u_xpb_out[60][714],u_xpb_out[61][714],u_xpb_out[62][714],u_xpb_out[63][714],u_xpb_out[64][714],u_xpb_out[65][714],u_xpb_out[66][714],u_xpb_out[67][714],u_xpb_out[68][714],u_xpb_out[69][714],u_xpb_out[70][714],u_xpb_out[71][714],u_xpb_out[72][714],u_xpb_out[73][714],u_xpb_out[74][714],u_xpb_out[75][714],u_xpb_out[76][714],u_xpb_out[77][714],u_xpb_out[78][714],u_xpb_out[79][714],u_xpb_out[80][714],u_xpb_out[81][714],u_xpb_out[82][714],u_xpb_out[83][714],u_xpb_out[84][714],u_xpb_out[85][714],u_xpb_out[86][714],u_xpb_out[87][714],u_xpb_out[88][714],u_xpb_out[89][714],u_xpb_out[90][714],u_xpb_out[91][714],u_xpb_out[92][714],u_xpb_out[93][714],u_xpb_out[94][714],u_xpb_out[95][714],u_xpb_out[96][714],u_xpb_out[97][714],u_xpb_out[98][714],u_xpb_out[99][714],u_xpb_out[100][714],u_xpb_out[101][714],u_xpb_out[102][714],u_xpb_out[103][714],u_xpb_out[104][714],u_xpb_out[105][714]};

assign col_out_715 = {u_xpb_out[0][715],u_xpb_out[1][715],u_xpb_out[2][715],u_xpb_out[3][715],u_xpb_out[4][715],u_xpb_out[5][715],u_xpb_out[6][715],u_xpb_out[7][715],u_xpb_out[8][715],u_xpb_out[9][715],u_xpb_out[10][715],u_xpb_out[11][715],u_xpb_out[12][715],u_xpb_out[13][715],u_xpb_out[14][715],u_xpb_out[15][715],u_xpb_out[16][715],u_xpb_out[17][715],u_xpb_out[18][715],u_xpb_out[19][715],u_xpb_out[20][715],u_xpb_out[21][715],u_xpb_out[22][715],u_xpb_out[23][715],u_xpb_out[24][715],u_xpb_out[25][715],u_xpb_out[26][715],u_xpb_out[27][715],u_xpb_out[28][715],u_xpb_out[29][715],u_xpb_out[30][715],u_xpb_out[31][715],u_xpb_out[32][715],u_xpb_out[33][715],u_xpb_out[34][715],u_xpb_out[35][715],u_xpb_out[36][715],u_xpb_out[37][715],u_xpb_out[38][715],u_xpb_out[39][715],u_xpb_out[40][715],u_xpb_out[41][715],u_xpb_out[42][715],u_xpb_out[43][715],u_xpb_out[44][715],u_xpb_out[45][715],u_xpb_out[46][715],u_xpb_out[47][715],u_xpb_out[48][715],u_xpb_out[49][715],u_xpb_out[50][715],u_xpb_out[51][715],u_xpb_out[52][715],u_xpb_out[53][715],u_xpb_out[54][715],u_xpb_out[55][715],u_xpb_out[56][715],u_xpb_out[57][715],u_xpb_out[58][715],u_xpb_out[59][715],u_xpb_out[60][715],u_xpb_out[61][715],u_xpb_out[62][715],u_xpb_out[63][715],u_xpb_out[64][715],u_xpb_out[65][715],u_xpb_out[66][715],u_xpb_out[67][715],u_xpb_out[68][715],u_xpb_out[69][715],u_xpb_out[70][715],u_xpb_out[71][715],u_xpb_out[72][715],u_xpb_out[73][715],u_xpb_out[74][715],u_xpb_out[75][715],u_xpb_out[76][715],u_xpb_out[77][715],u_xpb_out[78][715],u_xpb_out[79][715],u_xpb_out[80][715],u_xpb_out[81][715],u_xpb_out[82][715],u_xpb_out[83][715],u_xpb_out[84][715],u_xpb_out[85][715],u_xpb_out[86][715],u_xpb_out[87][715],u_xpb_out[88][715],u_xpb_out[89][715],u_xpb_out[90][715],u_xpb_out[91][715],u_xpb_out[92][715],u_xpb_out[93][715],u_xpb_out[94][715],u_xpb_out[95][715],u_xpb_out[96][715],u_xpb_out[97][715],u_xpb_out[98][715],u_xpb_out[99][715],u_xpb_out[100][715],u_xpb_out[101][715],u_xpb_out[102][715],u_xpb_out[103][715],u_xpb_out[104][715],u_xpb_out[105][715]};

assign col_out_716 = {u_xpb_out[0][716],u_xpb_out[1][716],u_xpb_out[2][716],u_xpb_out[3][716],u_xpb_out[4][716],u_xpb_out[5][716],u_xpb_out[6][716],u_xpb_out[7][716],u_xpb_out[8][716],u_xpb_out[9][716],u_xpb_out[10][716],u_xpb_out[11][716],u_xpb_out[12][716],u_xpb_out[13][716],u_xpb_out[14][716],u_xpb_out[15][716],u_xpb_out[16][716],u_xpb_out[17][716],u_xpb_out[18][716],u_xpb_out[19][716],u_xpb_out[20][716],u_xpb_out[21][716],u_xpb_out[22][716],u_xpb_out[23][716],u_xpb_out[24][716],u_xpb_out[25][716],u_xpb_out[26][716],u_xpb_out[27][716],u_xpb_out[28][716],u_xpb_out[29][716],u_xpb_out[30][716],u_xpb_out[31][716],u_xpb_out[32][716],u_xpb_out[33][716],u_xpb_out[34][716],u_xpb_out[35][716],u_xpb_out[36][716],u_xpb_out[37][716],u_xpb_out[38][716],u_xpb_out[39][716],u_xpb_out[40][716],u_xpb_out[41][716],u_xpb_out[42][716],u_xpb_out[43][716],u_xpb_out[44][716],u_xpb_out[45][716],u_xpb_out[46][716],u_xpb_out[47][716],u_xpb_out[48][716],u_xpb_out[49][716],u_xpb_out[50][716],u_xpb_out[51][716],u_xpb_out[52][716],u_xpb_out[53][716],u_xpb_out[54][716],u_xpb_out[55][716],u_xpb_out[56][716],u_xpb_out[57][716],u_xpb_out[58][716],u_xpb_out[59][716],u_xpb_out[60][716],u_xpb_out[61][716],u_xpb_out[62][716],u_xpb_out[63][716],u_xpb_out[64][716],u_xpb_out[65][716],u_xpb_out[66][716],u_xpb_out[67][716],u_xpb_out[68][716],u_xpb_out[69][716],u_xpb_out[70][716],u_xpb_out[71][716],u_xpb_out[72][716],u_xpb_out[73][716],u_xpb_out[74][716],u_xpb_out[75][716],u_xpb_out[76][716],u_xpb_out[77][716],u_xpb_out[78][716],u_xpb_out[79][716],u_xpb_out[80][716],u_xpb_out[81][716],u_xpb_out[82][716],u_xpb_out[83][716],u_xpb_out[84][716],u_xpb_out[85][716],u_xpb_out[86][716],u_xpb_out[87][716],u_xpb_out[88][716],u_xpb_out[89][716],u_xpb_out[90][716],u_xpb_out[91][716],u_xpb_out[92][716],u_xpb_out[93][716],u_xpb_out[94][716],u_xpb_out[95][716],u_xpb_out[96][716],u_xpb_out[97][716],u_xpb_out[98][716],u_xpb_out[99][716],u_xpb_out[100][716],u_xpb_out[101][716],u_xpb_out[102][716],u_xpb_out[103][716],u_xpb_out[104][716],u_xpb_out[105][716]};

assign col_out_717 = {u_xpb_out[0][717],u_xpb_out[1][717],u_xpb_out[2][717],u_xpb_out[3][717],u_xpb_out[4][717],u_xpb_out[5][717],u_xpb_out[6][717],u_xpb_out[7][717],u_xpb_out[8][717],u_xpb_out[9][717],u_xpb_out[10][717],u_xpb_out[11][717],u_xpb_out[12][717],u_xpb_out[13][717],u_xpb_out[14][717],u_xpb_out[15][717],u_xpb_out[16][717],u_xpb_out[17][717],u_xpb_out[18][717],u_xpb_out[19][717],u_xpb_out[20][717],u_xpb_out[21][717],u_xpb_out[22][717],u_xpb_out[23][717],u_xpb_out[24][717],u_xpb_out[25][717],u_xpb_out[26][717],u_xpb_out[27][717],u_xpb_out[28][717],u_xpb_out[29][717],u_xpb_out[30][717],u_xpb_out[31][717],u_xpb_out[32][717],u_xpb_out[33][717],u_xpb_out[34][717],u_xpb_out[35][717],u_xpb_out[36][717],u_xpb_out[37][717],u_xpb_out[38][717],u_xpb_out[39][717],u_xpb_out[40][717],u_xpb_out[41][717],u_xpb_out[42][717],u_xpb_out[43][717],u_xpb_out[44][717],u_xpb_out[45][717],u_xpb_out[46][717],u_xpb_out[47][717],u_xpb_out[48][717],u_xpb_out[49][717],u_xpb_out[50][717],u_xpb_out[51][717],u_xpb_out[52][717],u_xpb_out[53][717],u_xpb_out[54][717],u_xpb_out[55][717],u_xpb_out[56][717],u_xpb_out[57][717],u_xpb_out[58][717],u_xpb_out[59][717],u_xpb_out[60][717],u_xpb_out[61][717],u_xpb_out[62][717],u_xpb_out[63][717],u_xpb_out[64][717],u_xpb_out[65][717],u_xpb_out[66][717],u_xpb_out[67][717],u_xpb_out[68][717],u_xpb_out[69][717],u_xpb_out[70][717],u_xpb_out[71][717],u_xpb_out[72][717],u_xpb_out[73][717],u_xpb_out[74][717],u_xpb_out[75][717],u_xpb_out[76][717],u_xpb_out[77][717],u_xpb_out[78][717],u_xpb_out[79][717],u_xpb_out[80][717],u_xpb_out[81][717],u_xpb_out[82][717],u_xpb_out[83][717],u_xpb_out[84][717],u_xpb_out[85][717],u_xpb_out[86][717],u_xpb_out[87][717],u_xpb_out[88][717],u_xpb_out[89][717],u_xpb_out[90][717],u_xpb_out[91][717],u_xpb_out[92][717],u_xpb_out[93][717],u_xpb_out[94][717],u_xpb_out[95][717],u_xpb_out[96][717],u_xpb_out[97][717],u_xpb_out[98][717],u_xpb_out[99][717],u_xpb_out[100][717],u_xpb_out[101][717],u_xpb_out[102][717],u_xpb_out[103][717],u_xpb_out[104][717],u_xpb_out[105][717]};

assign col_out_718 = {u_xpb_out[0][718],u_xpb_out[1][718],u_xpb_out[2][718],u_xpb_out[3][718],u_xpb_out[4][718],u_xpb_out[5][718],u_xpb_out[6][718],u_xpb_out[7][718],u_xpb_out[8][718],u_xpb_out[9][718],u_xpb_out[10][718],u_xpb_out[11][718],u_xpb_out[12][718],u_xpb_out[13][718],u_xpb_out[14][718],u_xpb_out[15][718],u_xpb_out[16][718],u_xpb_out[17][718],u_xpb_out[18][718],u_xpb_out[19][718],u_xpb_out[20][718],u_xpb_out[21][718],u_xpb_out[22][718],u_xpb_out[23][718],u_xpb_out[24][718],u_xpb_out[25][718],u_xpb_out[26][718],u_xpb_out[27][718],u_xpb_out[28][718],u_xpb_out[29][718],u_xpb_out[30][718],u_xpb_out[31][718],u_xpb_out[32][718],u_xpb_out[33][718],u_xpb_out[34][718],u_xpb_out[35][718],u_xpb_out[36][718],u_xpb_out[37][718],u_xpb_out[38][718],u_xpb_out[39][718],u_xpb_out[40][718],u_xpb_out[41][718],u_xpb_out[42][718],u_xpb_out[43][718],u_xpb_out[44][718],u_xpb_out[45][718],u_xpb_out[46][718],u_xpb_out[47][718],u_xpb_out[48][718],u_xpb_out[49][718],u_xpb_out[50][718],u_xpb_out[51][718],u_xpb_out[52][718],u_xpb_out[53][718],u_xpb_out[54][718],u_xpb_out[55][718],u_xpb_out[56][718],u_xpb_out[57][718],u_xpb_out[58][718],u_xpb_out[59][718],u_xpb_out[60][718],u_xpb_out[61][718],u_xpb_out[62][718],u_xpb_out[63][718],u_xpb_out[64][718],u_xpb_out[65][718],u_xpb_out[66][718],u_xpb_out[67][718],u_xpb_out[68][718],u_xpb_out[69][718],u_xpb_out[70][718],u_xpb_out[71][718],u_xpb_out[72][718],u_xpb_out[73][718],u_xpb_out[74][718],u_xpb_out[75][718],u_xpb_out[76][718],u_xpb_out[77][718],u_xpb_out[78][718],u_xpb_out[79][718],u_xpb_out[80][718],u_xpb_out[81][718],u_xpb_out[82][718],u_xpb_out[83][718],u_xpb_out[84][718],u_xpb_out[85][718],u_xpb_out[86][718],u_xpb_out[87][718],u_xpb_out[88][718],u_xpb_out[89][718],u_xpb_out[90][718],u_xpb_out[91][718],u_xpb_out[92][718],u_xpb_out[93][718],u_xpb_out[94][718],u_xpb_out[95][718],u_xpb_out[96][718],u_xpb_out[97][718],u_xpb_out[98][718],u_xpb_out[99][718],u_xpb_out[100][718],u_xpb_out[101][718],u_xpb_out[102][718],u_xpb_out[103][718],u_xpb_out[104][718],u_xpb_out[105][718]};

assign col_out_719 = {u_xpb_out[0][719],u_xpb_out[1][719],u_xpb_out[2][719],u_xpb_out[3][719],u_xpb_out[4][719],u_xpb_out[5][719],u_xpb_out[6][719],u_xpb_out[7][719],u_xpb_out[8][719],u_xpb_out[9][719],u_xpb_out[10][719],u_xpb_out[11][719],u_xpb_out[12][719],u_xpb_out[13][719],u_xpb_out[14][719],u_xpb_out[15][719],u_xpb_out[16][719],u_xpb_out[17][719],u_xpb_out[18][719],u_xpb_out[19][719],u_xpb_out[20][719],u_xpb_out[21][719],u_xpb_out[22][719],u_xpb_out[23][719],u_xpb_out[24][719],u_xpb_out[25][719],u_xpb_out[26][719],u_xpb_out[27][719],u_xpb_out[28][719],u_xpb_out[29][719],u_xpb_out[30][719],u_xpb_out[31][719],u_xpb_out[32][719],u_xpb_out[33][719],u_xpb_out[34][719],u_xpb_out[35][719],u_xpb_out[36][719],u_xpb_out[37][719],u_xpb_out[38][719],u_xpb_out[39][719],u_xpb_out[40][719],u_xpb_out[41][719],u_xpb_out[42][719],u_xpb_out[43][719],u_xpb_out[44][719],u_xpb_out[45][719],u_xpb_out[46][719],u_xpb_out[47][719],u_xpb_out[48][719],u_xpb_out[49][719],u_xpb_out[50][719],u_xpb_out[51][719],u_xpb_out[52][719],u_xpb_out[53][719],u_xpb_out[54][719],u_xpb_out[55][719],u_xpb_out[56][719],u_xpb_out[57][719],u_xpb_out[58][719],u_xpb_out[59][719],u_xpb_out[60][719],u_xpb_out[61][719],u_xpb_out[62][719],u_xpb_out[63][719],u_xpb_out[64][719],u_xpb_out[65][719],u_xpb_out[66][719],u_xpb_out[67][719],u_xpb_out[68][719],u_xpb_out[69][719],u_xpb_out[70][719],u_xpb_out[71][719],u_xpb_out[72][719],u_xpb_out[73][719],u_xpb_out[74][719],u_xpb_out[75][719],u_xpb_out[76][719],u_xpb_out[77][719],u_xpb_out[78][719],u_xpb_out[79][719],u_xpb_out[80][719],u_xpb_out[81][719],u_xpb_out[82][719],u_xpb_out[83][719],u_xpb_out[84][719],u_xpb_out[85][719],u_xpb_out[86][719],u_xpb_out[87][719],u_xpb_out[88][719],u_xpb_out[89][719],u_xpb_out[90][719],u_xpb_out[91][719],u_xpb_out[92][719],u_xpb_out[93][719],u_xpb_out[94][719],u_xpb_out[95][719],u_xpb_out[96][719],u_xpb_out[97][719],u_xpb_out[98][719],u_xpb_out[99][719],u_xpb_out[100][719],u_xpb_out[101][719],u_xpb_out[102][719],u_xpb_out[103][719],u_xpb_out[104][719],u_xpb_out[105][719]};

assign col_out_720 = {u_xpb_out[0][720],u_xpb_out[1][720],u_xpb_out[2][720],u_xpb_out[3][720],u_xpb_out[4][720],u_xpb_out[5][720],u_xpb_out[6][720],u_xpb_out[7][720],u_xpb_out[8][720],u_xpb_out[9][720],u_xpb_out[10][720],u_xpb_out[11][720],u_xpb_out[12][720],u_xpb_out[13][720],u_xpb_out[14][720],u_xpb_out[15][720],u_xpb_out[16][720],u_xpb_out[17][720],u_xpb_out[18][720],u_xpb_out[19][720],u_xpb_out[20][720],u_xpb_out[21][720],u_xpb_out[22][720],u_xpb_out[23][720],u_xpb_out[24][720],u_xpb_out[25][720],u_xpb_out[26][720],u_xpb_out[27][720],u_xpb_out[28][720],u_xpb_out[29][720],u_xpb_out[30][720],u_xpb_out[31][720],u_xpb_out[32][720],u_xpb_out[33][720],u_xpb_out[34][720],u_xpb_out[35][720],u_xpb_out[36][720],u_xpb_out[37][720],u_xpb_out[38][720],u_xpb_out[39][720],u_xpb_out[40][720],u_xpb_out[41][720],u_xpb_out[42][720],u_xpb_out[43][720],u_xpb_out[44][720],u_xpb_out[45][720],u_xpb_out[46][720],u_xpb_out[47][720],u_xpb_out[48][720],u_xpb_out[49][720],u_xpb_out[50][720],u_xpb_out[51][720],u_xpb_out[52][720],u_xpb_out[53][720],u_xpb_out[54][720],u_xpb_out[55][720],u_xpb_out[56][720],u_xpb_out[57][720],u_xpb_out[58][720],u_xpb_out[59][720],u_xpb_out[60][720],u_xpb_out[61][720],u_xpb_out[62][720],u_xpb_out[63][720],u_xpb_out[64][720],u_xpb_out[65][720],u_xpb_out[66][720],u_xpb_out[67][720],u_xpb_out[68][720],u_xpb_out[69][720],u_xpb_out[70][720],u_xpb_out[71][720],u_xpb_out[72][720],u_xpb_out[73][720],u_xpb_out[74][720],u_xpb_out[75][720],u_xpb_out[76][720],u_xpb_out[77][720],u_xpb_out[78][720],u_xpb_out[79][720],u_xpb_out[80][720],u_xpb_out[81][720],u_xpb_out[82][720],u_xpb_out[83][720],u_xpb_out[84][720],u_xpb_out[85][720],u_xpb_out[86][720],u_xpb_out[87][720],u_xpb_out[88][720],u_xpb_out[89][720],u_xpb_out[90][720],u_xpb_out[91][720],u_xpb_out[92][720],u_xpb_out[93][720],u_xpb_out[94][720],u_xpb_out[95][720],u_xpb_out[96][720],u_xpb_out[97][720],u_xpb_out[98][720],u_xpb_out[99][720],u_xpb_out[100][720],u_xpb_out[101][720],u_xpb_out[102][720],u_xpb_out[103][720],u_xpb_out[104][720],u_xpb_out[105][720]};

assign col_out_721 = {u_xpb_out[0][721],u_xpb_out[1][721],u_xpb_out[2][721],u_xpb_out[3][721],u_xpb_out[4][721],u_xpb_out[5][721],u_xpb_out[6][721],u_xpb_out[7][721],u_xpb_out[8][721],u_xpb_out[9][721],u_xpb_out[10][721],u_xpb_out[11][721],u_xpb_out[12][721],u_xpb_out[13][721],u_xpb_out[14][721],u_xpb_out[15][721],u_xpb_out[16][721],u_xpb_out[17][721],u_xpb_out[18][721],u_xpb_out[19][721],u_xpb_out[20][721],u_xpb_out[21][721],u_xpb_out[22][721],u_xpb_out[23][721],u_xpb_out[24][721],u_xpb_out[25][721],u_xpb_out[26][721],u_xpb_out[27][721],u_xpb_out[28][721],u_xpb_out[29][721],u_xpb_out[30][721],u_xpb_out[31][721],u_xpb_out[32][721],u_xpb_out[33][721],u_xpb_out[34][721],u_xpb_out[35][721],u_xpb_out[36][721],u_xpb_out[37][721],u_xpb_out[38][721],u_xpb_out[39][721],u_xpb_out[40][721],u_xpb_out[41][721],u_xpb_out[42][721],u_xpb_out[43][721],u_xpb_out[44][721],u_xpb_out[45][721],u_xpb_out[46][721],u_xpb_out[47][721],u_xpb_out[48][721],u_xpb_out[49][721],u_xpb_out[50][721],u_xpb_out[51][721],u_xpb_out[52][721],u_xpb_out[53][721],u_xpb_out[54][721],u_xpb_out[55][721],u_xpb_out[56][721],u_xpb_out[57][721],u_xpb_out[58][721],u_xpb_out[59][721],u_xpb_out[60][721],u_xpb_out[61][721],u_xpb_out[62][721],u_xpb_out[63][721],u_xpb_out[64][721],u_xpb_out[65][721],u_xpb_out[66][721],u_xpb_out[67][721],u_xpb_out[68][721],u_xpb_out[69][721],u_xpb_out[70][721],u_xpb_out[71][721],u_xpb_out[72][721],u_xpb_out[73][721],u_xpb_out[74][721],u_xpb_out[75][721],u_xpb_out[76][721],u_xpb_out[77][721],u_xpb_out[78][721],u_xpb_out[79][721],u_xpb_out[80][721],u_xpb_out[81][721],u_xpb_out[82][721],u_xpb_out[83][721],u_xpb_out[84][721],u_xpb_out[85][721],u_xpb_out[86][721],u_xpb_out[87][721],u_xpb_out[88][721],u_xpb_out[89][721],u_xpb_out[90][721],u_xpb_out[91][721],u_xpb_out[92][721],u_xpb_out[93][721],u_xpb_out[94][721],u_xpb_out[95][721],u_xpb_out[96][721],u_xpb_out[97][721],u_xpb_out[98][721],u_xpb_out[99][721],u_xpb_out[100][721],u_xpb_out[101][721],u_xpb_out[102][721],u_xpb_out[103][721],u_xpb_out[104][721],u_xpb_out[105][721]};

assign col_out_722 = {u_xpb_out[0][722],u_xpb_out[1][722],u_xpb_out[2][722],u_xpb_out[3][722],u_xpb_out[4][722],u_xpb_out[5][722],u_xpb_out[6][722],u_xpb_out[7][722],u_xpb_out[8][722],u_xpb_out[9][722],u_xpb_out[10][722],u_xpb_out[11][722],u_xpb_out[12][722],u_xpb_out[13][722],u_xpb_out[14][722],u_xpb_out[15][722],u_xpb_out[16][722],u_xpb_out[17][722],u_xpb_out[18][722],u_xpb_out[19][722],u_xpb_out[20][722],u_xpb_out[21][722],u_xpb_out[22][722],u_xpb_out[23][722],u_xpb_out[24][722],u_xpb_out[25][722],u_xpb_out[26][722],u_xpb_out[27][722],u_xpb_out[28][722],u_xpb_out[29][722],u_xpb_out[30][722],u_xpb_out[31][722],u_xpb_out[32][722],u_xpb_out[33][722],u_xpb_out[34][722],u_xpb_out[35][722],u_xpb_out[36][722],u_xpb_out[37][722],u_xpb_out[38][722],u_xpb_out[39][722],u_xpb_out[40][722],u_xpb_out[41][722],u_xpb_out[42][722],u_xpb_out[43][722],u_xpb_out[44][722],u_xpb_out[45][722],u_xpb_out[46][722],u_xpb_out[47][722],u_xpb_out[48][722],u_xpb_out[49][722],u_xpb_out[50][722],u_xpb_out[51][722],u_xpb_out[52][722],u_xpb_out[53][722],u_xpb_out[54][722],u_xpb_out[55][722],u_xpb_out[56][722],u_xpb_out[57][722],u_xpb_out[58][722],u_xpb_out[59][722],u_xpb_out[60][722],u_xpb_out[61][722],u_xpb_out[62][722],u_xpb_out[63][722],u_xpb_out[64][722],u_xpb_out[65][722],u_xpb_out[66][722],u_xpb_out[67][722],u_xpb_out[68][722],u_xpb_out[69][722],u_xpb_out[70][722],u_xpb_out[71][722],u_xpb_out[72][722],u_xpb_out[73][722],u_xpb_out[74][722],u_xpb_out[75][722],u_xpb_out[76][722],u_xpb_out[77][722],u_xpb_out[78][722],u_xpb_out[79][722],u_xpb_out[80][722],u_xpb_out[81][722],u_xpb_out[82][722],u_xpb_out[83][722],u_xpb_out[84][722],u_xpb_out[85][722],u_xpb_out[86][722],u_xpb_out[87][722],u_xpb_out[88][722],u_xpb_out[89][722],u_xpb_out[90][722],u_xpb_out[91][722],u_xpb_out[92][722],u_xpb_out[93][722],u_xpb_out[94][722],u_xpb_out[95][722],u_xpb_out[96][722],u_xpb_out[97][722],u_xpb_out[98][722],u_xpb_out[99][722],u_xpb_out[100][722],u_xpb_out[101][722],u_xpb_out[102][722],u_xpb_out[103][722],u_xpb_out[104][722],u_xpb_out[105][722]};

assign col_out_723 = {u_xpb_out[0][723],u_xpb_out[1][723],u_xpb_out[2][723],u_xpb_out[3][723],u_xpb_out[4][723],u_xpb_out[5][723],u_xpb_out[6][723],u_xpb_out[7][723],u_xpb_out[8][723],u_xpb_out[9][723],u_xpb_out[10][723],u_xpb_out[11][723],u_xpb_out[12][723],u_xpb_out[13][723],u_xpb_out[14][723],u_xpb_out[15][723],u_xpb_out[16][723],u_xpb_out[17][723],u_xpb_out[18][723],u_xpb_out[19][723],u_xpb_out[20][723],u_xpb_out[21][723],u_xpb_out[22][723],u_xpb_out[23][723],u_xpb_out[24][723],u_xpb_out[25][723],u_xpb_out[26][723],u_xpb_out[27][723],u_xpb_out[28][723],u_xpb_out[29][723],u_xpb_out[30][723],u_xpb_out[31][723],u_xpb_out[32][723],u_xpb_out[33][723],u_xpb_out[34][723],u_xpb_out[35][723],u_xpb_out[36][723],u_xpb_out[37][723],u_xpb_out[38][723],u_xpb_out[39][723],u_xpb_out[40][723],u_xpb_out[41][723],u_xpb_out[42][723],u_xpb_out[43][723],u_xpb_out[44][723],u_xpb_out[45][723],u_xpb_out[46][723],u_xpb_out[47][723],u_xpb_out[48][723],u_xpb_out[49][723],u_xpb_out[50][723],u_xpb_out[51][723],u_xpb_out[52][723],u_xpb_out[53][723],u_xpb_out[54][723],u_xpb_out[55][723],u_xpb_out[56][723],u_xpb_out[57][723],u_xpb_out[58][723],u_xpb_out[59][723],u_xpb_out[60][723],u_xpb_out[61][723],u_xpb_out[62][723],u_xpb_out[63][723],u_xpb_out[64][723],u_xpb_out[65][723],u_xpb_out[66][723],u_xpb_out[67][723],u_xpb_out[68][723],u_xpb_out[69][723],u_xpb_out[70][723],u_xpb_out[71][723],u_xpb_out[72][723],u_xpb_out[73][723],u_xpb_out[74][723],u_xpb_out[75][723],u_xpb_out[76][723],u_xpb_out[77][723],u_xpb_out[78][723],u_xpb_out[79][723],u_xpb_out[80][723],u_xpb_out[81][723],u_xpb_out[82][723],u_xpb_out[83][723],u_xpb_out[84][723],u_xpb_out[85][723],u_xpb_out[86][723],u_xpb_out[87][723],u_xpb_out[88][723],u_xpb_out[89][723],u_xpb_out[90][723],u_xpb_out[91][723],u_xpb_out[92][723],u_xpb_out[93][723],u_xpb_out[94][723],u_xpb_out[95][723],u_xpb_out[96][723],u_xpb_out[97][723],u_xpb_out[98][723],u_xpb_out[99][723],u_xpb_out[100][723],u_xpb_out[101][723],u_xpb_out[102][723],u_xpb_out[103][723],u_xpb_out[104][723],u_xpb_out[105][723]};

assign col_out_724 = {u_xpb_out[0][724],u_xpb_out[1][724],u_xpb_out[2][724],u_xpb_out[3][724],u_xpb_out[4][724],u_xpb_out[5][724],u_xpb_out[6][724],u_xpb_out[7][724],u_xpb_out[8][724],u_xpb_out[9][724],u_xpb_out[10][724],u_xpb_out[11][724],u_xpb_out[12][724],u_xpb_out[13][724],u_xpb_out[14][724],u_xpb_out[15][724],u_xpb_out[16][724],u_xpb_out[17][724],u_xpb_out[18][724],u_xpb_out[19][724],u_xpb_out[20][724],u_xpb_out[21][724],u_xpb_out[22][724],u_xpb_out[23][724],u_xpb_out[24][724],u_xpb_out[25][724],u_xpb_out[26][724],u_xpb_out[27][724],u_xpb_out[28][724],u_xpb_out[29][724],u_xpb_out[30][724],u_xpb_out[31][724],u_xpb_out[32][724],u_xpb_out[33][724],u_xpb_out[34][724],u_xpb_out[35][724],u_xpb_out[36][724],u_xpb_out[37][724],u_xpb_out[38][724],u_xpb_out[39][724],u_xpb_out[40][724],u_xpb_out[41][724],u_xpb_out[42][724],u_xpb_out[43][724],u_xpb_out[44][724],u_xpb_out[45][724],u_xpb_out[46][724],u_xpb_out[47][724],u_xpb_out[48][724],u_xpb_out[49][724],u_xpb_out[50][724],u_xpb_out[51][724],u_xpb_out[52][724],u_xpb_out[53][724],u_xpb_out[54][724],u_xpb_out[55][724],u_xpb_out[56][724],u_xpb_out[57][724],u_xpb_out[58][724],u_xpb_out[59][724],u_xpb_out[60][724],u_xpb_out[61][724],u_xpb_out[62][724],u_xpb_out[63][724],u_xpb_out[64][724],u_xpb_out[65][724],u_xpb_out[66][724],u_xpb_out[67][724],u_xpb_out[68][724],u_xpb_out[69][724],u_xpb_out[70][724],u_xpb_out[71][724],u_xpb_out[72][724],u_xpb_out[73][724],u_xpb_out[74][724],u_xpb_out[75][724],u_xpb_out[76][724],u_xpb_out[77][724],u_xpb_out[78][724],u_xpb_out[79][724],u_xpb_out[80][724],u_xpb_out[81][724],u_xpb_out[82][724],u_xpb_out[83][724],u_xpb_out[84][724],u_xpb_out[85][724],u_xpb_out[86][724],u_xpb_out[87][724],u_xpb_out[88][724],u_xpb_out[89][724],u_xpb_out[90][724],u_xpb_out[91][724],u_xpb_out[92][724],u_xpb_out[93][724],u_xpb_out[94][724],u_xpb_out[95][724],u_xpb_out[96][724],u_xpb_out[97][724],u_xpb_out[98][724],u_xpb_out[99][724],u_xpb_out[100][724],u_xpb_out[101][724],u_xpb_out[102][724],u_xpb_out[103][724],u_xpb_out[104][724],u_xpb_out[105][724]};

assign col_out_725 = {u_xpb_out[0][725],u_xpb_out[1][725],u_xpb_out[2][725],u_xpb_out[3][725],u_xpb_out[4][725],u_xpb_out[5][725],u_xpb_out[6][725],u_xpb_out[7][725],u_xpb_out[8][725],u_xpb_out[9][725],u_xpb_out[10][725],u_xpb_out[11][725],u_xpb_out[12][725],u_xpb_out[13][725],u_xpb_out[14][725],u_xpb_out[15][725],u_xpb_out[16][725],u_xpb_out[17][725],u_xpb_out[18][725],u_xpb_out[19][725],u_xpb_out[20][725],u_xpb_out[21][725],u_xpb_out[22][725],u_xpb_out[23][725],u_xpb_out[24][725],u_xpb_out[25][725],u_xpb_out[26][725],u_xpb_out[27][725],u_xpb_out[28][725],u_xpb_out[29][725],u_xpb_out[30][725],u_xpb_out[31][725],u_xpb_out[32][725],u_xpb_out[33][725],u_xpb_out[34][725],u_xpb_out[35][725],u_xpb_out[36][725],u_xpb_out[37][725],u_xpb_out[38][725],u_xpb_out[39][725],u_xpb_out[40][725],u_xpb_out[41][725],u_xpb_out[42][725],u_xpb_out[43][725],u_xpb_out[44][725],u_xpb_out[45][725],u_xpb_out[46][725],u_xpb_out[47][725],u_xpb_out[48][725],u_xpb_out[49][725],u_xpb_out[50][725],u_xpb_out[51][725],u_xpb_out[52][725],u_xpb_out[53][725],u_xpb_out[54][725],u_xpb_out[55][725],u_xpb_out[56][725],u_xpb_out[57][725],u_xpb_out[58][725],u_xpb_out[59][725],u_xpb_out[60][725],u_xpb_out[61][725],u_xpb_out[62][725],u_xpb_out[63][725],u_xpb_out[64][725],u_xpb_out[65][725],u_xpb_out[66][725],u_xpb_out[67][725],u_xpb_out[68][725],u_xpb_out[69][725],u_xpb_out[70][725],u_xpb_out[71][725],u_xpb_out[72][725],u_xpb_out[73][725],u_xpb_out[74][725],u_xpb_out[75][725],u_xpb_out[76][725],u_xpb_out[77][725],u_xpb_out[78][725],u_xpb_out[79][725],u_xpb_out[80][725],u_xpb_out[81][725],u_xpb_out[82][725],u_xpb_out[83][725],u_xpb_out[84][725],u_xpb_out[85][725],u_xpb_out[86][725],u_xpb_out[87][725],u_xpb_out[88][725],u_xpb_out[89][725],u_xpb_out[90][725],u_xpb_out[91][725],u_xpb_out[92][725],u_xpb_out[93][725],u_xpb_out[94][725],u_xpb_out[95][725],u_xpb_out[96][725],u_xpb_out[97][725],u_xpb_out[98][725],u_xpb_out[99][725],u_xpb_out[100][725],u_xpb_out[101][725],u_xpb_out[102][725],u_xpb_out[103][725],u_xpb_out[104][725],u_xpb_out[105][725]};

assign col_out_726 = {u_xpb_out[0][726],u_xpb_out[1][726],u_xpb_out[2][726],u_xpb_out[3][726],u_xpb_out[4][726],u_xpb_out[5][726],u_xpb_out[6][726],u_xpb_out[7][726],u_xpb_out[8][726],u_xpb_out[9][726],u_xpb_out[10][726],u_xpb_out[11][726],u_xpb_out[12][726],u_xpb_out[13][726],u_xpb_out[14][726],u_xpb_out[15][726],u_xpb_out[16][726],u_xpb_out[17][726],u_xpb_out[18][726],u_xpb_out[19][726],u_xpb_out[20][726],u_xpb_out[21][726],u_xpb_out[22][726],u_xpb_out[23][726],u_xpb_out[24][726],u_xpb_out[25][726],u_xpb_out[26][726],u_xpb_out[27][726],u_xpb_out[28][726],u_xpb_out[29][726],u_xpb_out[30][726],u_xpb_out[31][726],u_xpb_out[32][726],u_xpb_out[33][726],u_xpb_out[34][726],u_xpb_out[35][726],u_xpb_out[36][726],u_xpb_out[37][726],u_xpb_out[38][726],u_xpb_out[39][726],u_xpb_out[40][726],u_xpb_out[41][726],u_xpb_out[42][726],u_xpb_out[43][726],u_xpb_out[44][726],u_xpb_out[45][726],u_xpb_out[46][726],u_xpb_out[47][726],u_xpb_out[48][726],u_xpb_out[49][726],u_xpb_out[50][726],u_xpb_out[51][726],u_xpb_out[52][726],u_xpb_out[53][726],u_xpb_out[54][726],u_xpb_out[55][726],u_xpb_out[56][726],u_xpb_out[57][726],u_xpb_out[58][726],u_xpb_out[59][726],u_xpb_out[60][726],u_xpb_out[61][726],u_xpb_out[62][726],u_xpb_out[63][726],u_xpb_out[64][726],u_xpb_out[65][726],u_xpb_out[66][726],u_xpb_out[67][726],u_xpb_out[68][726],u_xpb_out[69][726],u_xpb_out[70][726],u_xpb_out[71][726],u_xpb_out[72][726],u_xpb_out[73][726],u_xpb_out[74][726],u_xpb_out[75][726],u_xpb_out[76][726],u_xpb_out[77][726],u_xpb_out[78][726],u_xpb_out[79][726],u_xpb_out[80][726],u_xpb_out[81][726],u_xpb_out[82][726],u_xpb_out[83][726],u_xpb_out[84][726],u_xpb_out[85][726],u_xpb_out[86][726],u_xpb_out[87][726],u_xpb_out[88][726],u_xpb_out[89][726],u_xpb_out[90][726],u_xpb_out[91][726],u_xpb_out[92][726],u_xpb_out[93][726],u_xpb_out[94][726],u_xpb_out[95][726],u_xpb_out[96][726],u_xpb_out[97][726],u_xpb_out[98][726],u_xpb_out[99][726],u_xpb_out[100][726],u_xpb_out[101][726],u_xpb_out[102][726],u_xpb_out[103][726],u_xpb_out[104][726],u_xpb_out[105][726]};

assign col_out_727 = {u_xpb_out[0][727],u_xpb_out[1][727],u_xpb_out[2][727],u_xpb_out[3][727],u_xpb_out[4][727],u_xpb_out[5][727],u_xpb_out[6][727],u_xpb_out[7][727],u_xpb_out[8][727],u_xpb_out[9][727],u_xpb_out[10][727],u_xpb_out[11][727],u_xpb_out[12][727],u_xpb_out[13][727],u_xpb_out[14][727],u_xpb_out[15][727],u_xpb_out[16][727],u_xpb_out[17][727],u_xpb_out[18][727],u_xpb_out[19][727],u_xpb_out[20][727],u_xpb_out[21][727],u_xpb_out[22][727],u_xpb_out[23][727],u_xpb_out[24][727],u_xpb_out[25][727],u_xpb_out[26][727],u_xpb_out[27][727],u_xpb_out[28][727],u_xpb_out[29][727],u_xpb_out[30][727],u_xpb_out[31][727],u_xpb_out[32][727],u_xpb_out[33][727],u_xpb_out[34][727],u_xpb_out[35][727],u_xpb_out[36][727],u_xpb_out[37][727],u_xpb_out[38][727],u_xpb_out[39][727],u_xpb_out[40][727],u_xpb_out[41][727],u_xpb_out[42][727],u_xpb_out[43][727],u_xpb_out[44][727],u_xpb_out[45][727],u_xpb_out[46][727],u_xpb_out[47][727],u_xpb_out[48][727],u_xpb_out[49][727],u_xpb_out[50][727],u_xpb_out[51][727],u_xpb_out[52][727],u_xpb_out[53][727],u_xpb_out[54][727],u_xpb_out[55][727],u_xpb_out[56][727],u_xpb_out[57][727],u_xpb_out[58][727],u_xpb_out[59][727],u_xpb_out[60][727],u_xpb_out[61][727],u_xpb_out[62][727],u_xpb_out[63][727],u_xpb_out[64][727],u_xpb_out[65][727],u_xpb_out[66][727],u_xpb_out[67][727],u_xpb_out[68][727],u_xpb_out[69][727],u_xpb_out[70][727],u_xpb_out[71][727],u_xpb_out[72][727],u_xpb_out[73][727],u_xpb_out[74][727],u_xpb_out[75][727],u_xpb_out[76][727],u_xpb_out[77][727],u_xpb_out[78][727],u_xpb_out[79][727],u_xpb_out[80][727],u_xpb_out[81][727],u_xpb_out[82][727],u_xpb_out[83][727],u_xpb_out[84][727],u_xpb_out[85][727],u_xpb_out[86][727],u_xpb_out[87][727],u_xpb_out[88][727],u_xpb_out[89][727],u_xpb_out[90][727],u_xpb_out[91][727],u_xpb_out[92][727],u_xpb_out[93][727],u_xpb_out[94][727],u_xpb_out[95][727],u_xpb_out[96][727],u_xpb_out[97][727],u_xpb_out[98][727],u_xpb_out[99][727],u_xpb_out[100][727],u_xpb_out[101][727],u_xpb_out[102][727],u_xpb_out[103][727],u_xpb_out[104][727],u_xpb_out[105][727]};

assign col_out_728 = {u_xpb_out[0][728],u_xpb_out[1][728],u_xpb_out[2][728],u_xpb_out[3][728],u_xpb_out[4][728],u_xpb_out[5][728],u_xpb_out[6][728],u_xpb_out[7][728],u_xpb_out[8][728],u_xpb_out[9][728],u_xpb_out[10][728],u_xpb_out[11][728],u_xpb_out[12][728],u_xpb_out[13][728],u_xpb_out[14][728],u_xpb_out[15][728],u_xpb_out[16][728],u_xpb_out[17][728],u_xpb_out[18][728],u_xpb_out[19][728],u_xpb_out[20][728],u_xpb_out[21][728],u_xpb_out[22][728],u_xpb_out[23][728],u_xpb_out[24][728],u_xpb_out[25][728],u_xpb_out[26][728],u_xpb_out[27][728],u_xpb_out[28][728],u_xpb_out[29][728],u_xpb_out[30][728],u_xpb_out[31][728],u_xpb_out[32][728],u_xpb_out[33][728],u_xpb_out[34][728],u_xpb_out[35][728],u_xpb_out[36][728],u_xpb_out[37][728],u_xpb_out[38][728],u_xpb_out[39][728],u_xpb_out[40][728],u_xpb_out[41][728],u_xpb_out[42][728],u_xpb_out[43][728],u_xpb_out[44][728],u_xpb_out[45][728],u_xpb_out[46][728],u_xpb_out[47][728],u_xpb_out[48][728],u_xpb_out[49][728],u_xpb_out[50][728],u_xpb_out[51][728],u_xpb_out[52][728],u_xpb_out[53][728],u_xpb_out[54][728],u_xpb_out[55][728],u_xpb_out[56][728],u_xpb_out[57][728],u_xpb_out[58][728],u_xpb_out[59][728],u_xpb_out[60][728],u_xpb_out[61][728],u_xpb_out[62][728],u_xpb_out[63][728],u_xpb_out[64][728],u_xpb_out[65][728],u_xpb_out[66][728],u_xpb_out[67][728],u_xpb_out[68][728],u_xpb_out[69][728],u_xpb_out[70][728],u_xpb_out[71][728],u_xpb_out[72][728],u_xpb_out[73][728],u_xpb_out[74][728],u_xpb_out[75][728],u_xpb_out[76][728],u_xpb_out[77][728],u_xpb_out[78][728],u_xpb_out[79][728],u_xpb_out[80][728],u_xpb_out[81][728],u_xpb_out[82][728],u_xpb_out[83][728],u_xpb_out[84][728],u_xpb_out[85][728],u_xpb_out[86][728],u_xpb_out[87][728],u_xpb_out[88][728],u_xpb_out[89][728],u_xpb_out[90][728],u_xpb_out[91][728],u_xpb_out[92][728],u_xpb_out[93][728],u_xpb_out[94][728],u_xpb_out[95][728],u_xpb_out[96][728],u_xpb_out[97][728],u_xpb_out[98][728],u_xpb_out[99][728],u_xpb_out[100][728],u_xpb_out[101][728],u_xpb_out[102][728],u_xpb_out[103][728],u_xpb_out[104][728],u_xpb_out[105][728]};

assign col_out_729 = {u_xpb_out[0][729],u_xpb_out[1][729],u_xpb_out[2][729],u_xpb_out[3][729],u_xpb_out[4][729],u_xpb_out[5][729],u_xpb_out[6][729],u_xpb_out[7][729],u_xpb_out[8][729],u_xpb_out[9][729],u_xpb_out[10][729],u_xpb_out[11][729],u_xpb_out[12][729],u_xpb_out[13][729],u_xpb_out[14][729],u_xpb_out[15][729],u_xpb_out[16][729],u_xpb_out[17][729],u_xpb_out[18][729],u_xpb_out[19][729],u_xpb_out[20][729],u_xpb_out[21][729],u_xpb_out[22][729],u_xpb_out[23][729],u_xpb_out[24][729],u_xpb_out[25][729],u_xpb_out[26][729],u_xpb_out[27][729],u_xpb_out[28][729],u_xpb_out[29][729],u_xpb_out[30][729],u_xpb_out[31][729],u_xpb_out[32][729],u_xpb_out[33][729],u_xpb_out[34][729],u_xpb_out[35][729],u_xpb_out[36][729],u_xpb_out[37][729],u_xpb_out[38][729],u_xpb_out[39][729],u_xpb_out[40][729],u_xpb_out[41][729],u_xpb_out[42][729],u_xpb_out[43][729],u_xpb_out[44][729],u_xpb_out[45][729],u_xpb_out[46][729],u_xpb_out[47][729],u_xpb_out[48][729],u_xpb_out[49][729],u_xpb_out[50][729],u_xpb_out[51][729],u_xpb_out[52][729],u_xpb_out[53][729],u_xpb_out[54][729],u_xpb_out[55][729],u_xpb_out[56][729],u_xpb_out[57][729],u_xpb_out[58][729],u_xpb_out[59][729],u_xpb_out[60][729],u_xpb_out[61][729],u_xpb_out[62][729],u_xpb_out[63][729],u_xpb_out[64][729],u_xpb_out[65][729],u_xpb_out[66][729],u_xpb_out[67][729],u_xpb_out[68][729],u_xpb_out[69][729],u_xpb_out[70][729],u_xpb_out[71][729],u_xpb_out[72][729],u_xpb_out[73][729],u_xpb_out[74][729],u_xpb_out[75][729],u_xpb_out[76][729],u_xpb_out[77][729],u_xpb_out[78][729],u_xpb_out[79][729],u_xpb_out[80][729],u_xpb_out[81][729],u_xpb_out[82][729],u_xpb_out[83][729],u_xpb_out[84][729],u_xpb_out[85][729],u_xpb_out[86][729],u_xpb_out[87][729],u_xpb_out[88][729],u_xpb_out[89][729],u_xpb_out[90][729],u_xpb_out[91][729],u_xpb_out[92][729],u_xpb_out[93][729],u_xpb_out[94][729],u_xpb_out[95][729],u_xpb_out[96][729],u_xpb_out[97][729],u_xpb_out[98][729],u_xpb_out[99][729],u_xpb_out[100][729],u_xpb_out[101][729],u_xpb_out[102][729],u_xpb_out[103][729],u_xpb_out[104][729],u_xpb_out[105][729]};

assign col_out_730 = {u_xpb_out[0][730],u_xpb_out[1][730],u_xpb_out[2][730],u_xpb_out[3][730],u_xpb_out[4][730],u_xpb_out[5][730],u_xpb_out[6][730],u_xpb_out[7][730],u_xpb_out[8][730],u_xpb_out[9][730],u_xpb_out[10][730],u_xpb_out[11][730],u_xpb_out[12][730],u_xpb_out[13][730],u_xpb_out[14][730],u_xpb_out[15][730],u_xpb_out[16][730],u_xpb_out[17][730],u_xpb_out[18][730],u_xpb_out[19][730],u_xpb_out[20][730],u_xpb_out[21][730],u_xpb_out[22][730],u_xpb_out[23][730],u_xpb_out[24][730],u_xpb_out[25][730],u_xpb_out[26][730],u_xpb_out[27][730],u_xpb_out[28][730],u_xpb_out[29][730],u_xpb_out[30][730],u_xpb_out[31][730],u_xpb_out[32][730],u_xpb_out[33][730],u_xpb_out[34][730],u_xpb_out[35][730],u_xpb_out[36][730],u_xpb_out[37][730],u_xpb_out[38][730],u_xpb_out[39][730],u_xpb_out[40][730],u_xpb_out[41][730],u_xpb_out[42][730],u_xpb_out[43][730],u_xpb_out[44][730],u_xpb_out[45][730],u_xpb_out[46][730],u_xpb_out[47][730],u_xpb_out[48][730],u_xpb_out[49][730],u_xpb_out[50][730],u_xpb_out[51][730],u_xpb_out[52][730],u_xpb_out[53][730],u_xpb_out[54][730],u_xpb_out[55][730],u_xpb_out[56][730],u_xpb_out[57][730],u_xpb_out[58][730],u_xpb_out[59][730],u_xpb_out[60][730],u_xpb_out[61][730],u_xpb_out[62][730],u_xpb_out[63][730],u_xpb_out[64][730],u_xpb_out[65][730],u_xpb_out[66][730],u_xpb_out[67][730],u_xpb_out[68][730],u_xpb_out[69][730],u_xpb_out[70][730],u_xpb_out[71][730],u_xpb_out[72][730],u_xpb_out[73][730],u_xpb_out[74][730],u_xpb_out[75][730],u_xpb_out[76][730],u_xpb_out[77][730],u_xpb_out[78][730],u_xpb_out[79][730],u_xpb_out[80][730],u_xpb_out[81][730],u_xpb_out[82][730],u_xpb_out[83][730],u_xpb_out[84][730],u_xpb_out[85][730],u_xpb_out[86][730],u_xpb_out[87][730],u_xpb_out[88][730],u_xpb_out[89][730],u_xpb_out[90][730],u_xpb_out[91][730],u_xpb_out[92][730],u_xpb_out[93][730],u_xpb_out[94][730],u_xpb_out[95][730],u_xpb_out[96][730],u_xpb_out[97][730],u_xpb_out[98][730],u_xpb_out[99][730],u_xpb_out[100][730],u_xpb_out[101][730],u_xpb_out[102][730],u_xpb_out[103][730],u_xpb_out[104][730],u_xpb_out[105][730]};

assign col_out_731 = {u_xpb_out[0][731],u_xpb_out[1][731],u_xpb_out[2][731],u_xpb_out[3][731],u_xpb_out[4][731],u_xpb_out[5][731],u_xpb_out[6][731],u_xpb_out[7][731],u_xpb_out[8][731],u_xpb_out[9][731],u_xpb_out[10][731],u_xpb_out[11][731],u_xpb_out[12][731],u_xpb_out[13][731],u_xpb_out[14][731],u_xpb_out[15][731],u_xpb_out[16][731],u_xpb_out[17][731],u_xpb_out[18][731],u_xpb_out[19][731],u_xpb_out[20][731],u_xpb_out[21][731],u_xpb_out[22][731],u_xpb_out[23][731],u_xpb_out[24][731],u_xpb_out[25][731],u_xpb_out[26][731],u_xpb_out[27][731],u_xpb_out[28][731],u_xpb_out[29][731],u_xpb_out[30][731],u_xpb_out[31][731],u_xpb_out[32][731],u_xpb_out[33][731],u_xpb_out[34][731],u_xpb_out[35][731],u_xpb_out[36][731],u_xpb_out[37][731],u_xpb_out[38][731],u_xpb_out[39][731],u_xpb_out[40][731],u_xpb_out[41][731],u_xpb_out[42][731],u_xpb_out[43][731],u_xpb_out[44][731],u_xpb_out[45][731],u_xpb_out[46][731],u_xpb_out[47][731],u_xpb_out[48][731],u_xpb_out[49][731],u_xpb_out[50][731],u_xpb_out[51][731],u_xpb_out[52][731],u_xpb_out[53][731],u_xpb_out[54][731],u_xpb_out[55][731],u_xpb_out[56][731],u_xpb_out[57][731],u_xpb_out[58][731],u_xpb_out[59][731],u_xpb_out[60][731],u_xpb_out[61][731],u_xpb_out[62][731],u_xpb_out[63][731],u_xpb_out[64][731],u_xpb_out[65][731],u_xpb_out[66][731],u_xpb_out[67][731],u_xpb_out[68][731],u_xpb_out[69][731],u_xpb_out[70][731],u_xpb_out[71][731],u_xpb_out[72][731],u_xpb_out[73][731],u_xpb_out[74][731],u_xpb_out[75][731],u_xpb_out[76][731],u_xpb_out[77][731],u_xpb_out[78][731],u_xpb_out[79][731],u_xpb_out[80][731],u_xpb_out[81][731],u_xpb_out[82][731],u_xpb_out[83][731],u_xpb_out[84][731],u_xpb_out[85][731],u_xpb_out[86][731],u_xpb_out[87][731],u_xpb_out[88][731],u_xpb_out[89][731],u_xpb_out[90][731],u_xpb_out[91][731],u_xpb_out[92][731],u_xpb_out[93][731],u_xpb_out[94][731],u_xpb_out[95][731],u_xpb_out[96][731],u_xpb_out[97][731],u_xpb_out[98][731],u_xpb_out[99][731],u_xpb_out[100][731],u_xpb_out[101][731],u_xpb_out[102][731],u_xpb_out[103][731],u_xpb_out[104][731],u_xpb_out[105][731]};

assign col_out_732 = {u_xpb_out[0][732],u_xpb_out[1][732],u_xpb_out[2][732],u_xpb_out[3][732],u_xpb_out[4][732],u_xpb_out[5][732],u_xpb_out[6][732],u_xpb_out[7][732],u_xpb_out[8][732],u_xpb_out[9][732],u_xpb_out[10][732],u_xpb_out[11][732],u_xpb_out[12][732],u_xpb_out[13][732],u_xpb_out[14][732],u_xpb_out[15][732],u_xpb_out[16][732],u_xpb_out[17][732],u_xpb_out[18][732],u_xpb_out[19][732],u_xpb_out[20][732],u_xpb_out[21][732],u_xpb_out[22][732],u_xpb_out[23][732],u_xpb_out[24][732],u_xpb_out[25][732],u_xpb_out[26][732],u_xpb_out[27][732],u_xpb_out[28][732],u_xpb_out[29][732],u_xpb_out[30][732],u_xpb_out[31][732],u_xpb_out[32][732],u_xpb_out[33][732],u_xpb_out[34][732],u_xpb_out[35][732],u_xpb_out[36][732],u_xpb_out[37][732],u_xpb_out[38][732],u_xpb_out[39][732],u_xpb_out[40][732],u_xpb_out[41][732],u_xpb_out[42][732],u_xpb_out[43][732],u_xpb_out[44][732],u_xpb_out[45][732],u_xpb_out[46][732],u_xpb_out[47][732],u_xpb_out[48][732],u_xpb_out[49][732],u_xpb_out[50][732],u_xpb_out[51][732],u_xpb_out[52][732],u_xpb_out[53][732],u_xpb_out[54][732],u_xpb_out[55][732],u_xpb_out[56][732],u_xpb_out[57][732],u_xpb_out[58][732],u_xpb_out[59][732],u_xpb_out[60][732],u_xpb_out[61][732],u_xpb_out[62][732],u_xpb_out[63][732],u_xpb_out[64][732],u_xpb_out[65][732],u_xpb_out[66][732],u_xpb_out[67][732],u_xpb_out[68][732],u_xpb_out[69][732],u_xpb_out[70][732],u_xpb_out[71][732],u_xpb_out[72][732],u_xpb_out[73][732],u_xpb_out[74][732],u_xpb_out[75][732],u_xpb_out[76][732],u_xpb_out[77][732],u_xpb_out[78][732],u_xpb_out[79][732],u_xpb_out[80][732],u_xpb_out[81][732],u_xpb_out[82][732],u_xpb_out[83][732],u_xpb_out[84][732],u_xpb_out[85][732],u_xpb_out[86][732],u_xpb_out[87][732],u_xpb_out[88][732],u_xpb_out[89][732],u_xpb_out[90][732],u_xpb_out[91][732],u_xpb_out[92][732],u_xpb_out[93][732],u_xpb_out[94][732],u_xpb_out[95][732],u_xpb_out[96][732],u_xpb_out[97][732],u_xpb_out[98][732],u_xpb_out[99][732],u_xpb_out[100][732],u_xpb_out[101][732],u_xpb_out[102][732],u_xpb_out[103][732],u_xpb_out[104][732],u_xpb_out[105][732]};

assign col_out_733 = {u_xpb_out[0][733],u_xpb_out[1][733],u_xpb_out[2][733],u_xpb_out[3][733],u_xpb_out[4][733],u_xpb_out[5][733],u_xpb_out[6][733],u_xpb_out[7][733],u_xpb_out[8][733],u_xpb_out[9][733],u_xpb_out[10][733],u_xpb_out[11][733],u_xpb_out[12][733],u_xpb_out[13][733],u_xpb_out[14][733],u_xpb_out[15][733],u_xpb_out[16][733],u_xpb_out[17][733],u_xpb_out[18][733],u_xpb_out[19][733],u_xpb_out[20][733],u_xpb_out[21][733],u_xpb_out[22][733],u_xpb_out[23][733],u_xpb_out[24][733],u_xpb_out[25][733],u_xpb_out[26][733],u_xpb_out[27][733],u_xpb_out[28][733],u_xpb_out[29][733],u_xpb_out[30][733],u_xpb_out[31][733],u_xpb_out[32][733],u_xpb_out[33][733],u_xpb_out[34][733],u_xpb_out[35][733],u_xpb_out[36][733],u_xpb_out[37][733],u_xpb_out[38][733],u_xpb_out[39][733],u_xpb_out[40][733],u_xpb_out[41][733],u_xpb_out[42][733],u_xpb_out[43][733],u_xpb_out[44][733],u_xpb_out[45][733],u_xpb_out[46][733],u_xpb_out[47][733],u_xpb_out[48][733],u_xpb_out[49][733],u_xpb_out[50][733],u_xpb_out[51][733],u_xpb_out[52][733],u_xpb_out[53][733],u_xpb_out[54][733],u_xpb_out[55][733],u_xpb_out[56][733],u_xpb_out[57][733],u_xpb_out[58][733],u_xpb_out[59][733],u_xpb_out[60][733],u_xpb_out[61][733],u_xpb_out[62][733],u_xpb_out[63][733],u_xpb_out[64][733],u_xpb_out[65][733],u_xpb_out[66][733],u_xpb_out[67][733],u_xpb_out[68][733],u_xpb_out[69][733],u_xpb_out[70][733],u_xpb_out[71][733],u_xpb_out[72][733],u_xpb_out[73][733],u_xpb_out[74][733],u_xpb_out[75][733],u_xpb_out[76][733],u_xpb_out[77][733],u_xpb_out[78][733],u_xpb_out[79][733],u_xpb_out[80][733],u_xpb_out[81][733],u_xpb_out[82][733],u_xpb_out[83][733],u_xpb_out[84][733],u_xpb_out[85][733],u_xpb_out[86][733],u_xpb_out[87][733],u_xpb_out[88][733],u_xpb_out[89][733],u_xpb_out[90][733],u_xpb_out[91][733],u_xpb_out[92][733],u_xpb_out[93][733],u_xpb_out[94][733],u_xpb_out[95][733],u_xpb_out[96][733],u_xpb_out[97][733],u_xpb_out[98][733],u_xpb_out[99][733],u_xpb_out[100][733],u_xpb_out[101][733],u_xpb_out[102][733],u_xpb_out[103][733],u_xpb_out[104][733],u_xpb_out[105][733]};

assign col_out_734 = {u_xpb_out[0][734],u_xpb_out[1][734],u_xpb_out[2][734],u_xpb_out[3][734],u_xpb_out[4][734],u_xpb_out[5][734],u_xpb_out[6][734],u_xpb_out[7][734],u_xpb_out[8][734],u_xpb_out[9][734],u_xpb_out[10][734],u_xpb_out[11][734],u_xpb_out[12][734],u_xpb_out[13][734],u_xpb_out[14][734],u_xpb_out[15][734],u_xpb_out[16][734],u_xpb_out[17][734],u_xpb_out[18][734],u_xpb_out[19][734],u_xpb_out[20][734],u_xpb_out[21][734],u_xpb_out[22][734],u_xpb_out[23][734],u_xpb_out[24][734],u_xpb_out[25][734],u_xpb_out[26][734],u_xpb_out[27][734],u_xpb_out[28][734],u_xpb_out[29][734],u_xpb_out[30][734],u_xpb_out[31][734],u_xpb_out[32][734],u_xpb_out[33][734],u_xpb_out[34][734],u_xpb_out[35][734],u_xpb_out[36][734],u_xpb_out[37][734],u_xpb_out[38][734],u_xpb_out[39][734],u_xpb_out[40][734],u_xpb_out[41][734],u_xpb_out[42][734],u_xpb_out[43][734],u_xpb_out[44][734],u_xpb_out[45][734],u_xpb_out[46][734],u_xpb_out[47][734],u_xpb_out[48][734],u_xpb_out[49][734],u_xpb_out[50][734],u_xpb_out[51][734],u_xpb_out[52][734],u_xpb_out[53][734],u_xpb_out[54][734],u_xpb_out[55][734],u_xpb_out[56][734],u_xpb_out[57][734],u_xpb_out[58][734],u_xpb_out[59][734],u_xpb_out[60][734],u_xpb_out[61][734],u_xpb_out[62][734],u_xpb_out[63][734],u_xpb_out[64][734],u_xpb_out[65][734],u_xpb_out[66][734],u_xpb_out[67][734],u_xpb_out[68][734],u_xpb_out[69][734],u_xpb_out[70][734],u_xpb_out[71][734],u_xpb_out[72][734],u_xpb_out[73][734],u_xpb_out[74][734],u_xpb_out[75][734],u_xpb_out[76][734],u_xpb_out[77][734],u_xpb_out[78][734],u_xpb_out[79][734],u_xpb_out[80][734],u_xpb_out[81][734],u_xpb_out[82][734],u_xpb_out[83][734],u_xpb_out[84][734],u_xpb_out[85][734],u_xpb_out[86][734],u_xpb_out[87][734],u_xpb_out[88][734],u_xpb_out[89][734],u_xpb_out[90][734],u_xpb_out[91][734],u_xpb_out[92][734],u_xpb_out[93][734],u_xpb_out[94][734],u_xpb_out[95][734],u_xpb_out[96][734],u_xpb_out[97][734],u_xpb_out[98][734],u_xpb_out[99][734],u_xpb_out[100][734],u_xpb_out[101][734],u_xpb_out[102][734],u_xpb_out[103][734],u_xpb_out[104][734],u_xpb_out[105][734]};

assign col_out_735 = {u_xpb_out[0][735],u_xpb_out[1][735],u_xpb_out[2][735],u_xpb_out[3][735],u_xpb_out[4][735],u_xpb_out[5][735],u_xpb_out[6][735],u_xpb_out[7][735],u_xpb_out[8][735],u_xpb_out[9][735],u_xpb_out[10][735],u_xpb_out[11][735],u_xpb_out[12][735],u_xpb_out[13][735],u_xpb_out[14][735],u_xpb_out[15][735],u_xpb_out[16][735],u_xpb_out[17][735],u_xpb_out[18][735],u_xpb_out[19][735],u_xpb_out[20][735],u_xpb_out[21][735],u_xpb_out[22][735],u_xpb_out[23][735],u_xpb_out[24][735],u_xpb_out[25][735],u_xpb_out[26][735],u_xpb_out[27][735],u_xpb_out[28][735],u_xpb_out[29][735],u_xpb_out[30][735],u_xpb_out[31][735],u_xpb_out[32][735],u_xpb_out[33][735],u_xpb_out[34][735],u_xpb_out[35][735],u_xpb_out[36][735],u_xpb_out[37][735],u_xpb_out[38][735],u_xpb_out[39][735],u_xpb_out[40][735],u_xpb_out[41][735],u_xpb_out[42][735],u_xpb_out[43][735],u_xpb_out[44][735],u_xpb_out[45][735],u_xpb_out[46][735],u_xpb_out[47][735],u_xpb_out[48][735],u_xpb_out[49][735],u_xpb_out[50][735],u_xpb_out[51][735],u_xpb_out[52][735],u_xpb_out[53][735],u_xpb_out[54][735],u_xpb_out[55][735],u_xpb_out[56][735],u_xpb_out[57][735],u_xpb_out[58][735],u_xpb_out[59][735],u_xpb_out[60][735],u_xpb_out[61][735],u_xpb_out[62][735],u_xpb_out[63][735],u_xpb_out[64][735],u_xpb_out[65][735],u_xpb_out[66][735],u_xpb_out[67][735],u_xpb_out[68][735],u_xpb_out[69][735],u_xpb_out[70][735],u_xpb_out[71][735],u_xpb_out[72][735],u_xpb_out[73][735],u_xpb_out[74][735],u_xpb_out[75][735],u_xpb_out[76][735],u_xpb_out[77][735],u_xpb_out[78][735],u_xpb_out[79][735],u_xpb_out[80][735],u_xpb_out[81][735],u_xpb_out[82][735],u_xpb_out[83][735],u_xpb_out[84][735],u_xpb_out[85][735],u_xpb_out[86][735],u_xpb_out[87][735],u_xpb_out[88][735],u_xpb_out[89][735],u_xpb_out[90][735],u_xpb_out[91][735],u_xpb_out[92][735],u_xpb_out[93][735],u_xpb_out[94][735],u_xpb_out[95][735],u_xpb_out[96][735],u_xpb_out[97][735],u_xpb_out[98][735],u_xpb_out[99][735],u_xpb_out[100][735],u_xpb_out[101][735],u_xpb_out[102][735],u_xpb_out[103][735],u_xpb_out[104][735],u_xpb_out[105][735]};

assign col_out_736 = {u_xpb_out[0][736],u_xpb_out[1][736],u_xpb_out[2][736],u_xpb_out[3][736],u_xpb_out[4][736],u_xpb_out[5][736],u_xpb_out[6][736],u_xpb_out[7][736],u_xpb_out[8][736],u_xpb_out[9][736],u_xpb_out[10][736],u_xpb_out[11][736],u_xpb_out[12][736],u_xpb_out[13][736],u_xpb_out[14][736],u_xpb_out[15][736],u_xpb_out[16][736],u_xpb_out[17][736],u_xpb_out[18][736],u_xpb_out[19][736],u_xpb_out[20][736],u_xpb_out[21][736],u_xpb_out[22][736],u_xpb_out[23][736],u_xpb_out[24][736],u_xpb_out[25][736],u_xpb_out[26][736],u_xpb_out[27][736],u_xpb_out[28][736],u_xpb_out[29][736],u_xpb_out[30][736],u_xpb_out[31][736],u_xpb_out[32][736],u_xpb_out[33][736],u_xpb_out[34][736],u_xpb_out[35][736],u_xpb_out[36][736],u_xpb_out[37][736],u_xpb_out[38][736],u_xpb_out[39][736],u_xpb_out[40][736],u_xpb_out[41][736],u_xpb_out[42][736],u_xpb_out[43][736],u_xpb_out[44][736],u_xpb_out[45][736],u_xpb_out[46][736],u_xpb_out[47][736],u_xpb_out[48][736],u_xpb_out[49][736],u_xpb_out[50][736],u_xpb_out[51][736],u_xpb_out[52][736],u_xpb_out[53][736],u_xpb_out[54][736],u_xpb_out[55][736],u_xpb_out[56][736],u_xpb_out[57][736],u_xpb_out[58][736],u_xpb_out[59][736],u_xpb_out[60][736],u_xpb_out[61][736],u_xpb_out[62][736],u_xpb_out[63][736],u_xpb_out[64][736],u_xpb_out[65][736],u_xpb_out[66][736],u_xpb_out[67][736],u_xpb_out[68][736],u_xpb_out[69][736],u_xpb_out[70][736],u_xpb_out[71][736],u_xpb_out[72][736],u_xpb_out[73][736],u_xpb_out[74][736],u_xpb_out[75][736],u_xpb_out[76][736],u_xpb_out[77][736],u_xpb_out[78][736],u_xpb_out[79][736],u_xpb_out[80][736],u_xpb_out[81][736],u_xpb_out[82][736],u_xpb_out[83][736],u_xpb_out[84][736],u_xpb_out[85][736],u_xpb_out[86][736],u_xpb_out[87][736],u_xpb_out[88][736],u_xpb_out[89][736],u_xpb_out[90][736],u_xpb_out[91][736],u_xpb_out[92][736],u_xpb_out[93][736],u_xpb_out[94][736],u_xpb_out[95][736],u_xpb_out[96][736],u_xpb_out[97][736],u_xpb_out[98][736],u_xpb_out[99][736],u_xpb_out[100][736],u_xpb_out[101][736],u_xpb_out[102][736],u_xpb_out[103][736],u_xpb_out[104][736],u_xpb_out[105][736]};

assign col_out_737 = {u_xpb_out[0][737],u_xpb_out[1][737],u_xpb_out[2][737],u_xpb_out[3][737],u_xpb_out[4][737],u_xpb_out[5][737],u_xpb_out[6][737],u_xpb_out[7][737],u_xpb_out[8][737],u_xpb_out[9][737],u_xpb_out[10][737],u_xpb_out[11][737],u_xpb_out[12][737],u_xpb_out[13][737],u_xpb_out[14][737],u_xpb_out[15][737],u_xpb_out[16][737],u_xpb_out[17][737],u_xpb_out[18][737],u_xpb_out[19][737],u_xpb_out[20][737],u_xpb_out[21][737],u_xpb_out[22][737],u_xpb_out[23][737],u_xpb_out[24][737],u_xpb_out[25][737],u_xpb_out[26][737],u_xpb_out[27][737],u_xpb_out[28][737],u_xpb_out[29][737],u_xpb_out[30][737],u_xpb_out[31][737],u_xpb_out[32][737],u_xpb_out[33][737],u_xpb_out[34][737],u_xpb_out[35][737],u_xpb_out[36][737],u_xpb_out[37][737],u_xpb_out[38][737],u_xpb_out[39][737],u_xpb_out[40][737],u_xpb_out[41][737],u_xpb_out[42][737],u_xpb_out[43][737],u_xpb_out[44][737],u_xpb_out[45][737],u_xpb_out[46][737],u_xpb_out[47][737],u_xpb_out[48][737],u_xpb_out[49][737],u_xpb_out[50][737],u_xpb_out[51][737],u_xpb_out[52][737],u_xpb_out[53][737],u_xpb_out[54][737],u_xpb_out[55][737],u_xpb_out[56][737],u_xpb_out[57][737],u_xpb_out[58][737],u_xpb_out[59][737],u_xpb_out[60][737],u_xpb_out[61][737],u_xpb_out[62][737],u_xpb_out[63][737],u_xpb_out[64][737],u_xpb_out[65][737],u_xpb_out[66][737],u_xpb_out[67][737],u_xpb_out[68][737],u_xpb_out[69][737],u_xpb_out[70][737],u_xpb_out[71][737],u_xpb_out[72][737],u_xpb_out[73][737],u_xpb_out[74][737],u_xpb_out[75][737],u_xpb_out[76][737],u_xpb_out[77][737],u_xpb_out[78][737],u_xpb_out[79][737],u_xpb_out[80][737],u_xpb_out[81][737],u_xpb_out[82][737],u_xpb_out[83][737],u_xpb_out[84][737],u_xpb_out[85][737],u_xpb_out[86][737],u_xpb_out[87][737],u_xpb_out[88][737],u_xpb_out[89][737],u_xpb_out[90][737],u_xpb_out[91][737],u_xpb_out[92][737],u_xpb_out[93][737],u_xpb_out[94][737],u_xpb_out[95][737],u_xpb_out[96][737],u_xpb_out[97][737],u_xpb_out[98][737],u_xpb_out[99][737],u_xpb_out[100][737],u_xpb_out[101][737],u_xpb_out[102][737],u_xpb_out[103][737],u_xpb_out[104][737],u_xpb_out[105][737]};

assign col_out_738 = {u_xpb_out[0][738],u_xpb_out[1][738],u_xpb_out[2][738],u_xpb_out[3][738],u_xpb_out[4][738],u_xpb_out[5][738],u_xpb_out[6][738],u_xpb_out[7][738],u_xpb_out[8][738],u_xpb_out[9][738],u_xpb_out[10][738],u_xpb_out[11][738],u_xpb_out[12][738],u_xpb_out[13][738],u_xpb_out[14][738],u_xpb_out[15][738],u_xpb_out[16][738],u_xpb_out[17][738],u_xpb_out[18][738],u_xpb_out[19][738],u_xpb_out[20][738],u_xpb_out[21][738],u_xpb_out[22][738],u_xpb_out[23][738],u_xpb_out[24][738],u_xpb_out[25][738],u_xpb_out[26][738],u_xpb_out[27][738],u_xpb_out[28][738],u_xpb_out[29][738],u_xpb_out[30][738],u_xpb_out[31][738],u_xpb_out[32][738],u_xpb_out[33][738],u_xpb_out[34][738],u_xpb_out[35][738],u_xpb_out[36][738],u_xpb_out[37][738],u_xpb_out[38][738],u_xpb_out[39][738],u_xpb_out[40][738],u_xpb_out[41][738],u_xpb_out[42][738],u_xpb_out[43][738],u_xpb_out[44][738],u_xpb_out[45][738],u_xpb_out[46][738],u_xpb_out[47][738],u_xpb_out[48][738],u_xpb_out[49][738],u_xpb_out[50][738],u_xpb_out[51][738],u_xpb_out[52][738],u_xpb_out[53][738],u_xpb_out[54][738],u_xpb_out[55][738],u_xpb_out[56][738],u_xpb_out[57][738],u_xpb_out[58][738],u_xpb_out[59][738],u_xpb_out[60][738],u_xpb_out[61][738],u_xpb_out[62][738],u_xpb_out[63][738],u_xpb_out[64][738],u_xpb_out[65][738],u_xpb_out[66][738],u_xpb_out[67][738],u_xpb_out[68][738],u_xpb_out[69][738],u_xpb_out[70][738],u_xpb_out[71][738],u_xpb_out[72][738],u_xpb_out[73][738],u_xpb_out[74][738],u_xpb_out[75][738],u_xpb_out[76][738],u_xpb_out[77][738],u_xpb_out[78][738],u_xpb_out[79][738],u_xpb_out[80][738],u_xpb_out[81][738],u_xpb_out[82][738],u_xpb_out[83][738],u_xpb_out[84][738],u_xpb_out[85][738],u_xpb_out[86][738],u_xpb_out[87][738],u_xpb_out[88][738],u_xpb_out[89][738],u_xpb_out[90][738],u_xpb_out[91][738],u_xpb_out[92][738],u_xpb_out[93][738],u_xpb_out[94][738],u_xpb_out[95][738],u_xpb_out[96][738],u_xpb_out[97][738],u_xpb_out[98][738],u_xpb_out[99][738],u_xpb_out[100][738],u_xpb_out[101][738],u_xpb_out[102][738],u_xpb_out[103][738],u_xpb_out[104][738],u_xpb_out[105][738]};

assign col_out_739 = {u_xpb_out[0][739],u_xpb_out[1][739],u_xpb_out[2][739],u_xpb_out[3][739],u_xpb_out[4][739],u_xpb_out[5][739],u_xpb_out[6][739],u_xpb_out[7][739],u_xpb_out[8][739],u_xpb_out[9][739],u_xpb_out[10][739],u_xpb_out[11][739],u_xpb_out[12][739],u_xpb_out[13][739],u_xpb_out[14][739],u_xpb_out[15][739],u_xpb_out[16][739],u_xpb_out[17][739],u_xpb_out[18][739],u_xpb_out[19][739],u_xpb_out[20][739],u_xpb_out[21][739],u_xpb_out[22][739],u_xpb_out[23][739],u_xpb_out[24][739],u_xpb_out[25][739],u_xpb_out[26][739],u_xpb_out[27][739],u_xpb_out[28][739],u_xpb_out[29][739],u_xpb_out[30][739],u_xpb_out[31][739],u_xpb_out[32][739],u_xpb_out[33][739],u_xpb_out[34][739],u_xpb_out[35][739],u_xpb_out[36][739],u_xpb_out[37][739],u_xpb_out[38][739],u_xpb_out[39][739],u_xpb_out[40][739],u_xpb_out[41][739],u_xpb_out[42][739],u_xpb_out[43][739],u_xpb_out[44][739],u_xpb_out[45][739],u_xpb_out[46][739],u_xpb_out[47][739],u_xpb_out[48][739],u_xpb_out[49][739],u_xpb_out[50][739],u_xpb_out[51][739],u_xpb_out[52][739],u_xpb_out[53][739],u_xpb_out[54][739],u_xpb_out[55][739],u_xpb_out[56][739],u_xpb_out[57][739],u_xpb_out[58][739],u_xpb_out[59][739],u_xpb_out[60][739],u_xpb_out[61][739],u_xpb_out[62][739],u_xpb_out[63][739],u_xpb_out[64][739],u_xpb_out[65][739],u_xpb_out[66][739],u_xpb_out[67][739],u_xpb_out[68][739],u_xpb_out[69][739],u_xpb_out[70][739],u_xpb_out[71][739],u_xpb_out[72][739],u_xpb_out[73][739],u_xpb_out[74][739],u_xpb_out[75][739],u_xpb_out[76][739],u_xpb_out[77][739],u_xpb_out[78][739],u_xpb_out[79][739],u_xpb_out[80][739],u_xpb_out[81][739],u_xpb_out[82][739],u_xpb_out[83][739],u_xpb_out[84][739],u_xpb_out[85][739],u_xpb_out[86][739],u_xpb_out[87][739],u_xpb_out[88][739],u_xpb_out[89][739],u_xpb_out[90][739],u_xpb_out[91][739],u_xpb_out[92][739],u_xpb_out[93][739],u_xpb_out[94][739],u_xpb_out[95][739],u_xpb_out[96][739],u_xpb_out[97][739],u_xpb_out[98][739],u_xpb_out[99][739],u_xpb_out[100][739],u_xpb_out[101][739],u_xpb_out[102][739],u_xpb_out[103][739],u_xpb_out[104][739],u_xpb_out[105][739]};

assign col_out_740 = {u_xpb_out[0][740],u_xpb_out[1][740],u_xpb_out[2][740],u_xpb_out[3][740],u_xpb_out[4][740],u_xpb_out[5][740],u_xpb_out[6][740],u_xpb_out[7][740],u_xpb_out[8][740],u_xpb_out[9][740],u_xpb_out[10][740],u_xpb_out[11][740],u_xpb_out[12][740],u_xpb_out[13][740],u_xpb_out[14][740],u_xpb_out[15][740],u_xpb_out[16][740],u_xpb_out[17][740],u_xpb_out[18][740],u_xpb_out[19][740],u_xpb_out[20][740],u_xpb_out[21][740],u_xpb_out[22][740],u_xpb_out[23][740],u_xpb_out[24][740],u_xpb_out[25][740],u_xpb_out[26][740],u_xpb_out[27][740],u_xpb_out[28][740],u_xpb_out[29][740],u_xpb_out[30][740],u_xpb_out[31][740],u_xpb_out[32][740],u_xpb_out[33][740],u_xpb_out[34][740],u_xpb_out[35][740],u_xpb_out[36][740],u_xpb_out[37][740],u_xpb_out[38][740],u_xpb_out[39][740],u_xpb_out[40][740],u_xpb_out[41][740],u_xpb_out[42][740],u_xpb_out[43][740],u_xpb_out[44][740],u_xpb_out[45][740],u_xpb_out[46][740],u_xpb_out[47][740],u_xpb_out[48][740],u_xpb_out[49][740],u_xpb_out[50][740],u_xpb_out[51][740],u_xpb_out[52][740],u_xpb_out[53][740],u_xpb_out[54][740],u_xpb_out[55][740],u_xpb_out[56][740],u_xpb_out[57][740],u_xpb_out[58][740],u_xpb_out[59][740],u_xpb_out[60][740],u_xpb_out[61][740],u_xpb_out[62][740],u_xpb_out[63][740],u_xpb_out[64][740],u_xpb_out[65][740],u_xpb_out[66][740],u_xpb_out[67][740],u_xpb_out[68][740],u_xpb_out[69][740],u_xpb_out[70][740],u_xpb_out[71][740],u_xpb_out[72][740],u_xpb_out[73][740],u_xpb_out[74][740],u_xpb_out[75][740],u_xpb_out[76][740],u_xpb_out[77][740],u_xpb_out[78][740],u_xpb_out[79][740],u_xpb_out[80][740],u_xpb_out[81][740],u_xpb_out[82][740],u_xpb_out[83][740],u_xpb_out[84][740],u_xpb_out[85][740],u_xpb_out[86][740],u_xpb_out[87][740],u_xpb_out[88][740],u_xpb_out[89][740],u_xpb_out[90][740],u_xpb_out[91][740],u_xpb_out[92][740],u_xpb_out[93][740],u_xpb_out[94][740],u_xpb_out[95][740],u_xpb_out[96][740],u_xpb_out[97][740],u_xpb_out[98][740],u_xpb_out[99][740],u_xpb_out[100][740],u_xpb_out[101][740],u_xpb_out[102][740],u_xpb_out[103][740],u_xpb_out[104][740],u_xpb_out[105][740]};

assign col_out_741 = {u_xpb_out[0][741],u_xpb_out[1][741],u_xpb_out[2][741],u_xpb_out[3][741],u_xpb_out[4][741],u_xpb_out[5][741],u_xpb_out[6][741],u_xpb_out[7][741],u_xpb_out[8][741],u_xpb_out[9][741],u_xpb_out[10][741],u_xpb_out[11][741],u_xpb_out[12][741],u_xpb_out[13][741],u_xpb_out[14][741],u_xpb_out[15][741],u_xpb_out[16][741],u_xpb_out[17][741],u_xpb_out[18][741],u_xpb_out[19][741],u_xpb_out[20][741],u_xpb_out[21][741],u_xpb_out[22][741],u_xpb_out[23][741],u_xpb_out[24][741],u_xpb_out[25][741],u_xpb_out[26][741],u_xpb_out[27][741],u_xpb_out[28][741],u_xpb_out[29][741],u_xpb_out[30][741],u_xpb_out[31][741],u_xpb_out[32][741],u_xpb_out[33][741],u_xpb_out[34][741],u_xpb_out[35][741],u_xpb_out[36][741],u_xpb_out[37][741],u_xpb_out[38][741],u_xpb_out[39][741],u_xpb_out[40][741],u_xpb_out[41][741],u_xpb_out[42][741],u_xpb_out[43][741],u_xpb_out[44][741],u_xpb_out[45][741],u_xpb_out[46][741],u_xpb_out[47][741],u_xpb_out[48][741],u_xpb_out[49][741],u_xpb_out[50][741],u_xpb_out[51][741],u_xpb_out[52][741],u_xpb_out[53][741],u_xpb_out[54][741],u_xpb_out[55][741],u_xpb_out[56][741],u_xpb_out[57][741],u_xpb_out[58][741],u_xpb_out[59][741],u_xpb_out[60][741],u_xpb_out[61][741],u_xpb_out[62][741],u_xpb_out[63][741],u_xpb_out[64][741],u_xpb_out[65][741],u_xpb_out[66][741],u_xpb_out[67][741],u_xpb_out[68][741],u_xpb_out[69][741],u_xpb_out[70][741],u_xpb_out[71][741],u_xpb_out[72][741],u_xpb_out[73][741],u_xpb_out[74][741],u_xpb_out[75][741],u_xpb_out[76][741],u_xpb_out[77][741],u_xpb_out[78][741],u_xpb_out[79][741],u_xpb_out[80][741],u_xpb_out[81][741],u_xpb_out[82][741],u_xpb_out[83][741],u_xpb_out[84][741],u_xpb_out[85][741],u_xpb_out[86][741],u_xpb_out[87][741],u_xpb_out[88][741],u_xpb_out[89][741],u_xpb_out[90][741],u_xpb_out[91][741],u_xpb_out[92][741],u_xpb_out[93][741],u_xpb_out[94][741],u_xpb_out[95][741],u_xpb_out[96][741],u_xpb_out[97][741],u_xpb_out[98][741],u_xpb_out[99][741],u_xpb_out[100][741],u_xpb_out[101][741],u_xpb_out[102][741],u_xpb_out[103][741],u_xpb_out[104][741],u_xpb_out[105][741]};

assign col_out_742 = {u_xpb_out[0][742],u_xpb_out[1][742],u_xpb_out[2][742],u_xpb_out[3][742],u_xpb_out[4][742],u_xpb_out[5][742],u_xpb_out[6][742],u_xpb_out[7][742],u_xpb_out[8][742],u_xpb_out[9][742],u_xpb_out[10][742],u_xpb_out[11][742],u_xpb_out[12][742],u_xpb_out[13][742],u_xpb_out[14][742],u_xpb_out[15][742],u_xpb_out[16][742],u_xpb_out[17][742],u_xpb_out[18][742],u_xpb_out[19][742],u_xpb_out[20][742],u_xpb_out[21][742],u_xpb_out[22][742],u_xpb_out[23][742],u_xpb_out[24][742],u_xpb_out[25][742],u_xpb_out[26][742],u_xpb_out[27][742],u_xpb_out[28][742],u_xpb_out[29][742],u_xpb_out[30][742],u_xpb_out[31][742],u_xpb_out[32][742],u_xpb_out[33][742],u_xpb_out[34][742],u_xpb_out[35][742],u_xpb_out[36][742],u_xpb_out[37][742],u_xpb_out[38][742],u_xpb_out[39][742],u_xpb_out[40][742],u_xpb_out[41][742],u_xpb_out[42][742],u_xpb_out[43][742],u_xpb_out[44][742],u_xpb_out[45][742],u_xpb_out[46][742],u_xpb_out[47][742],u_xpb_out[48][742],u_xpb_out[49][742],u_xpb_out[50][742],u_xpb_out[51][742],u_xpb_out[52][742],u_xpb_out[53][742],u_xpb_out[54][742],u_xpb_out[55][742],u_xpb_out[56][742],u_xpb_out[57][742],u_xpb_out[58][742],u_xpb_out[59][742],u_xpb_out[60][742],u_xpb_out[61][742],u_xpb_out[62][742],u_xpb_out[63][742],u_xpb_out[64][742],u_xpb_out[65][742],u_xpb_out[66][742],u_xpb_out[67][742],u_xpb_out[68][742],u_xpb_out[69][742],u_xpb_out[70][742],u_xpb_out[71][742],u_xpb_out[72][742],u_xpb_out[73][742],u_xpb_out[74][742],u_xpb_out[75][742],u_xpb_out[76][742],u_xpb_out[77][742],u_xpb_out[78][742],u_xpb_out[79][742],u_xpb_out[80][742],u_xpb_out[81][742],u_xpb_out[82][742],u_xpb_out[83][742],u_xpb_out[84][742],u_xpb_out[85][742],u_xpb_out[86][742],u_xpb_out[87][742],u_xpb_out[88][742],u_xpb_out[89][742],u_xpb_out[90][742],u_xpb_out[91][742],u_xpb_out[92][742],u_xpb_out[93][742],u_xpb_out[94][742],u_xpb_out[95][742],u_xpb_out[96][742],u_xpb_out[97][742],u_xpb_out[98][742],u_xpb_out[99][742],u_xpb_out[100][742],u_xpb_out[101][742],u_xpb_out[102][742],u_xpb_out[103][742],u_xpb_out[104][742],u_xpb_out[105][742]};

assign col_out_743 = {u_xpb_out[0][743],u_xpb_out[1][743],u_xpb_out[2][743],u_xpb_out[3][743],u_xpb_out[4][743],u_xpb_out[5][743],u_xpb_out[6][743],u_xpb_out[7][743],u_xpb_out[8][743],u_xpb_out[9][743],u_xpb_out[10][743],u_xpb_out[11][743],u_xpb_out[12][743],u_xpb_out[13][743],u_xpb_out[14][743],u_xpb_out[15][743],u_xpb_out[16][743],u_xpb_out[17][743],u_xpb_out[18][743],u_xpb_out[19][743],u_xpb_out[20][743],u_xpb_out[21][743],u_xpb_out[22][743],u_xpb_out[23][743],u_xpb_out[24][743],u_xpb_out[25][743],u_xpb_out[26][743],u_xpb_out[27][743],u_xpb_out[28][743],u_xpb_out[29][743],u_xpb_out[30][743],u_xpb_out[31][743],u_xpb_out[32][743],u_xpb_out[33][743],u_xpb_out[34][743],u_xpb_out[35][743],u_xpb_out[36][743],u_xpb_out[37][743],u_xpb_out[38][743],u_xpb_out[39][743],u_xpb_out[40][743],u_xpb_out[41][743],u_xpb_out[42][743],u_xpb_out[43][743],u_xpb_out[44][743],u_xpb_out[45][743],u_xpb_out[46][743],u_xpb_out[47][743],u_xpb_out[48][743],u_xpb_out[49][743],u_xpb_out[50][743],u_xpb_out[51][743],u_xpb_out[52][743],u_xpb_out[53][743],u_xpb_out[54][743],u_xpb_out[55][743],u_xpb_out[56][743],u_xpb_out[57][743],u_xpb_out[58][743],u_xpb_out[59][743],u_xpb_out[60][743],u_xpb_out[61][743],u_xpb_out[62][743],u_xpb_out[63][743],u_xpb_out[64][743],u_xpb_out[65][743],u_xpb_out[66][743],u_xpb_out[67][743],u_xpb_out[68][743],u_xpb_out[69][743],u_xpb_out[70][743],u_xpb_out[71][743],u_xpb_out[72][743],u_xpb_out[73][743],u_xpb_out[74][743],u_xpb_out[75][743],u_xpb_out[76][743],u_xpb_out[77][743],u_xpb_out[78][743],u_xpb_out[79][743],u_xpb_out[80][743],u_xpb_out[81][743],u_xpb_out[82][743],u_xpb_out[83][743],u_xpb_out[84][743],u_xpb_out[85][743],u_xpb_out[86][743],u_xpb_out[87][743],u_xpb_out[88][743],u_xpb_out[89][743],u_xpb_out[90][743],u_xpb_out[91][743],u_xpb_out[92][743],u_xpb_out[93][743],u_xpb_out[94][743],u_xpb_out[95][743],u_xpb_out[96][743],u_xpb_out[97][743],u_xpb_out[98][743],u_xpb_out[99][743],u_xpb_out[100][743],u_xpb_out[101][743],u_xpb_out[102][743],u_xpb_out[103][743],u_xpb_out[104][743],u_xpb_out[105][743]};

assign col_out_744 = {u_xpb_out[0][744],u_xpb_out[1][744],u_xpb_out[2][744],u_xpb_out[3][744],u_xpb_out[4][744],u_xpb_out[5][744],u_xpb_out[6][744],u_xpb_out[7][744],u_xpb_out[8][744],u_xpb_out[9][744],u_xpb_out[10][744],u_xpb_out[11][744],u_xpb_out[12][744],u_xpb_out[13][744],u_xpb_out[14][744],u_xpb_out[15][744],u_xpb_out[16][744],u_xpb_out[17][744],u_xpb_out[18][744],u_xpb_out[19][744],u_xpb_out[20][744],u_xpb_out[21][744],u_xpb_out[22][744],u_xpb_out[23][744],u_xpb_out[24][744],u_xpb_out[25][744],u_xpb_out[26][744],u_xpb_out[27][744],u_xpb_out[28][744],u_xpb_out[29][744],u_xpb_out[30][744],u_xpb_out[31][744],u_xpb_out[32][744],u_xpb_out[33][744],u_xpb_out[34][744],u_xpb_out[35][744],u_xpb_out[36][744],u_xpb_out[37][744],u_xpb_out[38][744],u_xpb_out[39][744],u_xpb_out[40][744],u_xpb_out[41][744],u_xpb_out[42][744],u_xpb_out[43][744],u_xpb_out[44][744],u_xpb_out[45][744],u_xpb_out[46][744],u_xpb_out[47][744],u_xpb_out[48][744],u_xpb_out[49][744],u_xpb_out[50][744],u_xpb_out[51][744],u_xpb_out[52][744],u_xpb_out[53][744],u_xpb_out[54][744],u_xpb_out[55][744],u_xpb_out[56][744],u_xpb_out[57][744],u_xpb_out[58][744],u_xpb_out[59][744],u_xpb_out[60][744],u_xpb_out[61][744],u_xpb_out[62][744],u_xpb_out[63][744],u_xpb_out[64][744],u_xpb_out[65][744],u_xpb_out[66][744],u_xpb_out[67][744],u_xpb_out[68][744],u_xpb_out[69][744],u_xpb_out[70][744],u_xpb_out[71][744],u_xpb_out[72][744],u_xpb_out[73][744],u_xpb_out[74][744],u_xpb_out[75][744],u_xpb_out[76][744],u_xpb_out[77][744],u_xpb_out[78][744],u_xpb_out[79][744],u_xpb_out[80][744],u_xpb_out[81][744],u_xpb_out[82][744],u_xpb_out[83][744],u_xpb_out[84][744],u_xpb_out[85][744],u_xpb_out[86][744],u_xpb_out[87][744],u_xpb_out[88][744],u_xpb_out[89][744],u_xpb_out[90][744],u_xpb_out[91][744],u_xpb_out[92][744],u_xpb_out[93][744],u_xpb_out[94][744],u_xpb_out[95][744],u_xpb_out[96][744],u_xpb_out[97][744],u_xpb_out[98][744],u_xpb_out[99][744],u_xpb_out[100][744],u_xpb_out[101][744],u_xpb_out[102][744],u_xpb_out[103][744],u_xpb_out[104][744],u_xpb_out[105][744]};

assign col_out_745 = {u_xpb_out[0][745],u_xpb_out[1][745],u_xpb_out[2][745],u_xpb_out[3][745],u_xpb_out[4][745],u_xpb_out[5][745],u_xpb_out[6][745],u_xpb_out[7][745],u_xpb_out[8][745],u_xpb_out[9][745],u_xpb_out[10][745],u_xpb_out[11][745],u_xpb_out[12][745],u_xpb_out[13][745],u_xpb_out[14][745],u_xpb_out[15][745],u_xpb_out[16][745],u_xpb_out[17][745],u_xpb_out[18][745],u_xpb_out[19][745],u_xpb_out[20][745],u_xpb_out[21][745],u_xpb_out[22][745],u_xpb_out[23][745],u_xpb_out[24][745],u_xpb_out[25][745],u_xpb_out[26][745],u_xpb_out[27][745],u_xpb_out[28][745],u_xpb_out[29][745],u_xpb_out[30][745],u_xpb_out[31][745],u_xpb_out[32][745],u_xpb_out[33][745],u_xpb_out[34][745],u_xpb_out[35][745],u_xpb_out[36][745],u_xpb_out[37][745],u_xpb_out[38][745],u_xpb_out[39][745],u_xpb_out[40][745],u_xpb_out[41][745],u_xpb_out[42][745],u_xpb_out[43][745],u_xpb_out[44][745],u_xpb_out[45][745],u_xpb_out[46][745],u_xpb_out[47][745],u_xpb_out[48][745],u_xpb_out[49][745],u_xpb_out[50][745],u_xpb_out[51][745],u_xpb_out[52][745],u_xpb_out[53][745],u_xpb_out[54][745],u_xpb_out[55][745],u_xpb_out[56][745],u_xpb_out[57][745],u_xpb_out[58][745],u_xpb_out[59][745],u_xpb_out[60][745],u_xpb_out[61][745],u_xpb_out[62][745],u_xpb_out[63][745],u_xpb_out[64][745],u_xpb_out[65][745],u_xpb_out[66][745],u_xpb_out[67][745],u_xpb_out[68][745],u_xpb_out[69][745],u_xpb_out[70][745],u_xpb_out[71][745],u_xpb_out[72][745],u_xpb_out[73][745],u_xpb_out[74][745],u_xpb_out[75][745],u_xpb_out[76][745],u_xpb_out[77][745],u_xpb_out[78][745],u_xpb_out[79][745],u_xpb_out[80][745],u_xpb_out[81][745],u_xpb_out[82][745],u_xpb_out[83][745],u_xpb_out[84][745],u_xpb_out[85][745],u_xpb_out[86][745],u_xpb_out[87][745],u_xpb_out[88][745],u_xpb_out[89][745],u_xpb_out[90][745],u_xpb_out[91][745],u_xpb_out[92][745],u_xpb_out[93][745],u_xpb_out[94][745],u_xpb_out[95][745],u_xpb_out[96][745],u_xpb_out[97][745],u_xpb_out[98][745],u_xpb_out[99][745],u_xpb_out[100][745],u_xpb_out[101][745],u_xpb_out[102][745],u_xpb_out[103][745],u_xpb_out[104][745],u_xpb_out[105][745]};

assign col_out_746 = {u_xpb_out[0][746],u_xpb_out[1][746],u_xpb_out[2][746],u_xpb_out[3][746],u_xpb_out[4][746],u_xpb_out[5][746],u_xpb_out[6][746],u_xpb_out[7][746],u_xpb_out[8][746],u_xpb_out[9][746],u_xpb_out[10][746],u_xpb_out[11][746],u_xpb_out[12][746],u_xpb_out[13][746],u_xpb_out[14][746],u_xpb_out[15][746],u_xpb_out[16][746],u_xpb_out[17][746],u_xpb_out[18][746],u_xpb_out[19][746],u_xpb_out[20][746],u_xpb_out[21][746],u_xpb_out[22][746],u_xpb_out[23][746],u_xpb_out[24][746],u_xpb_out[25][746],u_xpb_out[26][746],u_xpb_out[27][746],u_xpb_out[28][746],u_xpb_out[29][746],u_xpb_out[30][746],u_xpb_out[31][746],u_xpb_out[32][746],u_xpb_out[33][746],u_xpb_out[34][746],u_xpb_out[35][746],u_xpb_out[36][746],u_xpb_out[37][746],u_xpb_out[38][746],u_xpb_out[39][746],u_xpb_out[40][746],u_xpb_out[41][746],u_xpb_out[42][746],u_xpb_out[43][746],u_xpb_out[44][746],u_xpb_out[45][746],u_xpb_out[46][746],u_xpb_out[47][746],u_xpb_out[48][746],u_xpb_out[49][746],u_xpb_out[50][746],u_xpb_out[51][746],u_xpb_out[52][746],u_xpb_out[53][746],u_xpb_out[54][746],u_xpb_out[55][746],u_xpb_out[56][746],u_xpb_out[57][746],u_xpb_out[58][746],u_xpb_out[59][746],u_xpb_out[60][746],u_xpb_out[61][746],u_xpb_out[62][746],u_xpb_out[63][746],u_xpb_out[64][746],u_xpb_out[65][746],u_xpb_out[66][746],u_xpb_out[67][746],u_xpb_out[68][746],u_xpb_out[69][746],u_xpb_out[70][746],u_xpb_out[71][746],u_xpb_out[72][746],u_xpb_out[73][746],u_xpb_out[74][746],u_xpb_out[75][746],u_xpb_out[76][746],u_xpb_out[77][746],u_xpb_out[78][746],u_xpb_out[79][746],u_xpb_out[80][746],u_xpb_out[81][746],u_xpb_out[82][746],u_xpb_out[83][746],u_xpb_out[84][746],u_xpb_out[85][746],u_xpb_out[86][746],u_xpb_out[87][746],u_xpb_out[88][746],u_xpb_out[89][746],u_xpb_out[90][746],u_xpb_out[91][746],u_xpb_out[92][746],u_xpb_out[93][746],u_xpb_out[94][746],u_xpb_out[95][746],u_xpb_out[96][746],u_xpb_out[97][746],u_xpb_out[98][746],u_xpb_out[99][746],u_xpb_out[100][746],u_xpb_out[101][746],u_xpb_out[102][746],u_xpb_out[103][746],u_xpb_out[104][746],u_xpb_out[105][746]};

assign col_out_747 = {u_xpb_out[0][747],u_xpb_out[1][747],u_xpb_out[2][747],u_xpb_out[3][747],u_xpb_out[4][747],u_xpb_out[5][747],u_xpb_out[6][747],u_xpb_out[7][747],u_xpb_out[8][747],u_xpb_out[9][747],u_xpb_out[10][747],u_xpb_out[11][747],u_xpb_out[12][747],u_xpb_out[13][747],u_xpb_out[14][747],u_xpb_out[15][747],u_xpb_out[16][747],u_xpb_out[17][747],u_xpb_out[18][747],u_xpb_out[19][747],u_xpb_out[20][747],u_xpb_out[21][747],u_xpb_out[22][747],u_xpb_out[23][747],u_xpb_out[24][747],u_xpb_out[25][747],u_xpb_out[26][747],u_xpb_out[27][747],u_xpb_out[28][747],u_xpb_out[29][747],u_xpb_out[30][747],u_xpb_out[31][747],u_xpb_out[32][747],u_xpb_out[33][747],u_xpb_out[34][747],u_xpb_out[35][747],u_xpb_out[36][747],u_xpb_out[37][747],u_xpb_out[38][747],u_xpb_out[39][747],u_xpb_out[40][747],u_xpb_out[41][747],u_xpb_out[42][747],u_xpb_out[43][747],u_xpb_out[44][747],u_xpb_out[45][747],u_xpb_out[46][747],u_xpb_out[47][747],u_xpb_out[48][747],u_xpb_out[49][747],u_xpb_out[50][747],u_xpb_out[51][747],u_xpb_out[52][747],u_xpb_out[53][747],u_xpb_out[54][747],u_xpb_out[55][747],u_xpb_out[56][747],u_xpb_out[57][747],u_xpb_out[58][747],u_xpb_out[59][747],u_xpb_out[60][747],u_xpb_out[61][747],u_xpb_out[62][747],u_xpb_out[63][747],u_xpb_out[64][747],u_xpb_out[65][747],u_xpb_out[66][747],u_xpb_out[67][747],u_xpb_out[68][747],u_xpb_out[69][747],u_xpb_out[70][747],u_xpb_out[71][747],u_xpb_out[72][747],u_xpb_out[73][747],u_xpb_out[74][747],u_xpb_out[75][747],u_xpb_out[76][747],u_xpb_out[77][747],u_xpb_out[78][747],u_xpb_out[79][747],u_xpb_out[80][747],u_xpb_out[81][747],u_xpb_out[82][747],u_xpb_out[83][747],u_xpb_out[84][747],u_xpb_out[85][747],u_xpb_out[86][747],u_xpb_out[87][747],u_xpb_out[88][747],u_xpb_out[89][747],u_xpb_out[90][747],u_xpb_out[91][747],u_xpb_out[92][747],u_xpb_out[93][747],u_xpb_out[94][747],u_xpb_out[95][747],u_xpb_out[96][747],u_xpb_out[97][747],u_xpb_out[98][747],u_xpb_out[99][747],u_xpb_out[100][747],u_xpb_out[101][747],u_xpb_out[102][747],u_xpb_out[103][747],u_xpb_out[104][747],u_xpb_out[105][747]};

assign col_out_748 = {u_xpb_out[0][748],u_xpb_out[1][748],u_xpb_out[2][748],u_xpb_out[3][748],u_xpb_out[4][748],u_xpb_out[5][748],u_xpb_out[6][748],u_xpb_out[7][748],u_xpb_out[8][748],u_xpb_out[9][748],u_xpb_out[10][748],u_xpb_out[11][748],u_xpb_out[12][748],u_xpb_out[13][748],u_xpb_out[14][748],u_xpb_out[15][748],u_xpb_out[16][748],u_xpb_out[17][748],u_xpb_out[18][748],u_xpb_out[19][748],u_xpb_out[20][748],u_xpb_out[21][748],u_xpb_out[22][748],u_xpb_out[23][748],u_xpb_out[24][748],u_xpb_out[25][748],u_xpb_out[26][748],u_xpb_out[27][748],u_xpb_out[28][748],u_xpb_out[29][748],u_xpb_out[30][748],u_xpb_out[31][748],u_xpb_out[32][748],u_xpb_out[33][748],u_xpb_out[34][748],u_xpb_out[35][748],u_xpb_out[36][748],u_xpb_out[37][748],u_xpb_out[38][748],u_xpb_out[39][748],u_xpb_out[40][748],u_xpb_out[41][748],u_xpb_out[42][748],u_xpb_out[43][748],u_xpb_out[44][748],u_xpb_out[45][748],u_xpb_out[46][748],u_xpb_out[47][748],u_xpb_out[48][748],u_xpb_out[49][748],u_xpb_out[50][748],u_xpb_out[51][748],u_xpb_out[52][748],u_xpb_out[53][748],u_xpb_out[54][748],u_xpb_out[55][748],u_xpb_out[56][748],u_xpb_out[57][748],u_xpb_out[58][748],u_xpb_out[59][748],u_xpb_out[60][748],u_xpb_out[61][748],u_xpb_out[62][748],u_xpb_out[63][748],u_xpb_out[64][748],u_xpb_out[65][748],u_xpb_out[66][748],u_xpb_out[67][748],u_xpb_out[68][748],u_xpb_out[69][748],u_xpb_out[70][748],u_xpb_out[71][748],u_xpb_out[72][748],u_xpb_out[73][748],u_xpb_out[74][748],u_xpb_out[75][748],u_xpb_out[76][748],u_xpb_out[77][748],u_xpb_out[78][748],u_xpb_out[79][748],u_xpb_out[80][748],u_xpb_out[81][748],u_xpb_out[82][748],u_xpb_out[83][748],u_xpb_out[84][748],u_xpb_out[85][748],u_xpb_out[86][748],u_xpb_out[87][748],u_xpb_out[88][748],u_xpb_out[89][748],u_xpb_out[90][748],u_xpb_out[91][748],u_xpb_out[92][748],u_xpb_out[93][748],u_xpb_out[94][748],u_xpb_out[95][748],u_xpb_out[96][748],u_xpb_out[97][748],u_xpb_out[98][748],u_xpb_out[99][748],u_xpb_out[100][748],u_xpb_out[101][748],u_xpb_out[102][748],u_xpb_out[103][748],u_xpb_out[104][748],u_xpb_out[105][748]};

assign col_out_749 = {u_xpb_out[0][749],u_xpb_out[1][749],u_xpb_out[2][749],u_xpb_out[3][749],u_xpb_out[4][749],u_xpb_out[5][749],u_xpb_out[6][749],u_xpb_out[7][749],u_xpb_out[8][749],u_xpb_out[9][749],u_xpb_out[10][749],u_xpb_out[11][749],u_xpb_out[12][749],u_xpb_out[13][749],u_xpb_out[14][749],u_xpb_out[15][749],u_xpb_out[16][749],u_xpb_out[17][749],u_xpb_out[18][749],u_xpb_out[19][749],u_xpb_out[20][749],u_xpb_out[21][749],u_xpb_out[22][749],u_xpb_out[23][749],u_xpb_out[24][749],u_xpb_out[25][749],u_xpb_out[26][749],u_xpb_out[27][749],u_xpb_out[28][749],u_xpb_out[29][749],u_xpb_out[30][749],u_xpb_out[31][749],u_xpb_out[32][749],u_xpb_out[33][749],u_xpb_out[34][749],u_xpb_out[35][749],u_xpb_out[36][749],u_xpb_out[37][749],u_xpb_out[38][749],u_xpb_out[39][749],u_xpb_out[40][749],u_xpb_out[41][749],u_xpb_out[42][749],u_xpb_out[43][749],u_xpb_out[44][749],u_xpb_out[45][749],u_xpb_out[46][749],u_xpb_out[47][749],u_xpb_out[48][749],u_xpb_out[49][749],u_xpb_out[50][749],u_xpb_out[51][749],u_xpb_out[52][749],u_xpb_out[53][749],u_xpb_out[54][749],u_xpb_out[55][749],u_xpb_out[56][749],u_xpb_out[57][749],u_xpb_out[58][749],u_xpb_out[59][749],u_xpb_out[60][749],u_xpb_out[61][749],u_xpb_out[62][749],u_xpb_out[63][749],u_xpb_out[64][749],u_xpb_out[65][749],u_xpb_out[66][749],u_xpb_out[67][749],u_xpb_out[68][749],u_xpb_out[69][749],u_xpb_out[70][749],u_xpb_out[71][749],u_xpb_out[72][749],u_xpb_out[73][749],u_xpb_out[74][749],u_xpb_out[75][749],u_xpb_out[76][749],u_xpb_out[77][749],u_xpb_out[78][749],u_xpb_out[79][749],u_xpb_out[80][749],u_xpb_out[81][749],u_xpb_out[82][749],u_xpb_out[83][749],u_xpb_out[84][749],u_xpb_out[85][749],u_xpb_out[86][749],u_xpb_out[87][749],u_xpb_out[88][749],u_xpb_out[89][749],u_xpb_out[90][749],u_xpb_out[91][749],u_xpb_out[92][749],u_xpb_out[93][749],u_xpb_out[94][749],u_xpb_out[95][749],u_xpb_out[96][749],u_xpb_out[97][749],u_xpb_out[98][749],u_xpb_out[99][749],u_xpb_out[100][749],u_xpb_out[101][749],u_xpb_out[102][749],u_xpb_out[103][749],u_xpb_out[104][749],u_xpb_out[105][749]};

assign col_out_750 = {u_xpb_out[0][750],u_xpb_out[1][750],u_xpb_out[2][750],u_xpb_out[3][750],u_xpb_out[4][750],u_xpb_out[5][750],u_xpb_out[6][750],u_xpb_out[7][750],u_xpb_out[8][750],u_xpb_out[9][750],u_xpb_out[10][750],u_xpb_out[11][750],u_xpb_out[12][750],u_xpb_out[13][750],u_xpb_out[14][750],u_xpb_out[15][750],u_xpb_out[16][750],u_xpb_out[17][750],u_xpb_out[18][750],u_xpb_out[19][750],u_xpb_out[20][750],u_xpb_out[21][750],u_xpb_out[22][750],u_xpb_out[23][750],u_xpb_out[24][750],u_xpb_out[25][750],u_xpb_out[26][750],u_xpb_out[27][750],u_xpb_out[28][750],u_xpb_out[29][750],u_xpb_out[30][750],u_xpb_out[31][750],u_xpb_out[32][750],u_xpb_out[33][750],u_xpb_out[34][750],u_xpb_out[35][750],u_xpb_out[36][750],u_xpb_out[37][750],u_xpb_out[38][750],u_xpb_out[39][750],u_xpb_out[40][750],u_xpb_out[41][750],u_xpb_out[42][750],u_xpb_out[43][750],u_xpb_out[44][750],u_xpb_out[45][750],u_xpb_out[46][750],u_xpb_out[47][750],u_xpb_out[48][750],u_xpb_out[49][750],u_xpb_out[50][750],u_xpb_out[51][750],u_xpb_out[52][750],u_xpb_out[53][750],u_xpb_out[54][750],u_xpb_out[55][750],u_xpb_out[56][750],u_xpb_out[57][750],u_xpb_out[58][750],u_xpb_out[59][750],u_xpb_out[60][750],u_xpb_out[61][750],u_xpb_out[62][750],u_xpb_out[63][750],u_xpb_out[64][750],u_xpb_out[65][750],u_xpb_out[66][750],u_xpb_out[67][750],u_xpb_out[68][750],u_xpb_out[69][750],u_xpb_out[70][750],u_xpb_out[71][750],u_xpb_out[72][750],u_xpb_out[73][750],u_xpb_out[74][750],u_xpb_out[75][750],u_xpb_out[76][750],u_xpb_out[77][750],u_xpb_out[78][750],u_xpb_out[79][750],u_xpb_out[80][750],u_xpb_out[81][750],u_xpb_out[82][750],u_xpb_out[83][750],u_xpb_out[84][750],u_xpb_out[85][750],u_xpb_out[86][750],u_xpb_out[87][750],u_xpb_out[88][750],u_xpb_out[89][750],u_xpb_out[90][750],u_xpb_out[91][750],u_xpb_out[92][750],u_xpb_out[93][750],u_xpb_out[94][750],u_xpb_out[95][750],u_xpb_out[96][750],u_xpb_out[97][750],u_xpb_out[98][750],u_xpb_out[99][750],u_xpb_out[100][750],u_xpb_out[101][750],u_xpb_out[102][750],u_xpb_out[103][750],u_xpb_out[104][750],u_xpb_out[105][750]};

assign col_out_751 = {u_xpb_out[0][751],u_xpb_out[1][751],u_xpb_out[2][751],u_xpb_out[3][751],u_xpb_out[4][751],u_xpb_out[5][751],u_xpb_out[6][751],u_xpb_out[7][751],u_xpb_out[8][751],u_xpb_out[9][751],u_xpb_out[10][751],u_xpb_out[11][751],u_xpb_out[12][751],u_xpb_out[13][751],u_xpb_out[14][751],u_xpb_out[15][751],u_xpb_out[16][751],u_xpb_out[17][751],u_xpb_out[18][751],u_xpb_out[19][751],u_xpb_out[20][751],u_xpb_out[21][751],u_xpb_out[22][751],u_xpb_out[23][751],u_xpb_out[24][751],u_xpb_out[25][751],u_xpb_out[26][751],u_xpb_out[27][751],u_xpb_out[28][751],u_xpb_out[29][751],u_xpb_out[30][751],u_xpb_out[31][751],u_xpb_out[32][751],u_xpb_out[33][751],u_xpb_out[34][751],u_xpb_out[35][751],u_xpb_out[36][751],u_xpb_out[37][751],u_xpb_out[38][751],u_xpb_out[39][751],u_xpb_out[40][751],u_xpb_out[41][751],u_xpb_out[42][751],u_xpb_out[43][751],u_xpb_out[44][751],u_xpb_out[45][751],u_xpb_out[46][751],u_xpb_out[47][751],u_xpb_out[48][751],u_xpb_out[49][751],u_xpb_out[50][751],u_xpb_out[51][751],u_xpb_out[52][751],u_xpb_out[53][751],u_xpb_out[54][751],u_xpb_out[55][751],u_xpb_out[56][751],u_xpb_out[57][751],u_xpb_out[58][751],u_xpb_out[59][751],u_xpb_out[60][751],u_xpb_out[61][751],u_xpb_out[62][751],u_xpb_out[63][751],u_xpb_out[64][751],u_xpb_out[65][751],u_xpb_out[66][751],u_xpb_out[67][751],u_xpb_out[68][751],u_xpb_out[69][751],u_xpb_out[70][751],u_xpb_out[71][751],u_xpb_out[72][751],u_xpb_out[73][751],u_xpb_out[74][751],u_xpb_out[75][751],u_xpb_out[76][751],u_xpb_out[77][751],u_xpb_out[78][751],u_xpb_out[79][751],u_xpb_out[80][751],u_xpb_out[81][751],u_xpb_out[82][751],u_xpb_out[83][751],u_xpb_out[84][751],u_xpb_out[85][751],u_xpb_out[86][751],u_xpb_out[87][751],u_xpb_out[88][751],u_xpb_out[89][751],u_xpb_out[90][751],u_xpb_out[91][751],u_xpb_out[92][751],u_xpb_out[93][751],u_xpb_out[94][751],u_xpb_out[95][751],u_xpb_out[96][751],u_xpb_out[97][751],u_xpb_out[98][751],u_xpb_out[99][751],u_xpb_out[100][751],u_xpb_out[101][751],u_xpb_out[102][751],u_xpb_out[103][751],u_xpb_out[104][751],u_xpb_out[105][751]};

assign col_out_752 = {u_xpb_out[0][752],u_xpb_out[1][752],u_xpb_out[2][752],u_xpb_out[3][752],u_xpb_out[4][752],u_xpb_out[5][752],u_xpb_out[6][752],u_xpb_out[7][752],u_xpb_out[8][752],u_xpb_out[9][752],u_xpb_out[10][752],u_xpb_out[11][752],u_xpb_out[12][752],u_xpb_out[13][752],u_xpb_out[14][752],u_xpb_out[15][752],u_xpb_out[16][752],u_xpb_out[17][752],u_xpb_out[18][752],u_xpb_out[19][752],u_xpb_out[20][752],u_xpb_out[21][752],u_xpb_out[22][752],u_xpb_out[23][752],u_xpb_out[24][752],u_xpb_out[25][752],u_xpb_out[26][752],u_xpb_out[27][752],u_xpb_out[28][752],u_xpb_out[29][752],u_xpb_out[30][752],u_xpb_out[31][752],u_xpb_out[32][752],u_xpb_out[33][752],u_xpb_out[34][752],u_xpb_out[35][752],u_xpb_out[36][752],u_xpb_out[37][752],u_xpb_out[38][752],u_xpb_out[39][752],u_xpb_out[40][752],u_xpb_out[41][752],u_xpb_out[42][752],u_xpb_out[43][752],u_xpb_out[44][752],u_xpb_out[45][752],u_xpb_out[46][752],u_xpb_out[47][752],u_xpb_out[48][752],u_xpb_out[49][752],u_xpb_out[50][752],u_xpb_out[51][752],u_xpb_out[52][752],u_xpb_out[53][752],u_xpb_out[54][752],u_xpb_out[55][752],u_xpb_out[56][752],u_xpb_out[57][752],u_xpb_out[58][752],u_xpb_out[59][752],u_xpb_out[60][752],u_xpb_out[61][752],u_xpb_out[62][752],u_xpb_out[63][752],u_xpb_out[64][752],u_xpb_out[65][752],u_xpb_out[66][752],u_xpb_out[67][752],u_xpb_out[68][752],u_xpb_out[69][752],u_xpb_out[70][752],u_xpb_out[71][752],u_xpb_out[72][752],u_xpb_out[73][752],u_xpb_out[74][752],u_xpb_out[75][752],u_xpb_out[76][752],u_xpb_out[77][752],u_xpb_out[78][752],u_xpb_out[79][752],u_xpb_out[80][752],u_xpb_out[81][752],u_xpb_out[82][752],u_xpb_out[83][752],u_xpb_out[84][752],u_xpb_out[85][752],u_xpb_out[86][752],u_xpb_out[87][752],u_xpb_out[88][752],u_xpb_out[89][752],u_xpb_out[90][752],u_xpb_out[91][752],u_xpb_out[92][752],u_xpb_out[93][752],u_xpb_out[94][752],u_xpb_out[95][752],u_xpb_out[96][752],u_xpb_out[97][752],u_xpb_out[98][752],u_xpb_out[99][752],u_xpb_out[100][752],u_xpb_out[101][752],u_xpb_out[102][752],u_xpb_out[103][752],u_xpb_out[104][752],u_xpb_out[105][752]};

assign col_out_753 = {u_xpb_out[0][753],u_xpb_out[1][753],u_xpb_out[2][753],u_xpb_out[3][753],u_xpb_out[4][753],u_xpb_out[5][753],u_xpb_out[6][753],u_xpb_out[7][753],u_xpb_out[8][753],u_xpb_out[9][753],u_xpb_out[10][753],u_xpb_out[11][753],u_xpb_out[12][753],u_xpb_out[13][753],u_xpb_out[14][753],u_xpb_out[15][753],u_xpb_out[16][753],u_xpb_out[17][753],u_xpb_out[18][753],u_xpb_out[19][753],u_xpb_out[20][753],u_xpb_out[21][753],u_xpb_out[22][753],u_xpb_out[23][753],u_xpb_out[24][753],u_xpb_out[25][753],u_xpb_out[26][753],u_xpb_out[27][753],u_xpb_out[28][753],u_xpb_out[29][753],u_xpb_out[30][753],u_xpb_out[31][753],u_xpb_out[32][753],u_xpb_out[33][753],u_xpb_out[34][753],u_xpb_out[35][753],u_xpb_out[36][753],u_xpb_out[37][753],u_xpb_out[38][753],u_xpb_out[39][753],u_xpb_out[40][753],u_xpb_out[41][753],u_xpb_out[42][753],u_xpb_out[43][753],u_xpb_out[44][753],u_xpb_out[45][753],u_xpb_out[46][753],u_xpb_out[47][753],u_xpb_out[48][753],u_xpb_out[49][753],u_xpb_out[50][753],u_xpb_out[51][753],u_xpb_out[52][753],u_xpb_out[53][753],u_xpb_out[54][753],u_xpb_out[55][753],u_xpb_out[56][753],u_xpb_out[57][753],u_xpb_out[58][753],u_xpb_out[59][753],u_xpb_out[60][753],u_xpb_out[61][753],u_xpb_out[62][753],u_xpb_out[63][753],u_xpb_out[64][753],u_xpb_out[65][753],u_xpb_out[66][753],u_xpb_out[67][753],u_xpb_out[68][753],u_xpb_out[69][753],u_xpb_out[70][753],u_xpb_out[71][753],u_xpb_out[72][753],u_xpb_out[73][753],u_xpb_out[74][753],u_xpb_out[75][753],u_xpb_out[76][753],u_xpb_out[77][753],u_xpb_out[78][753],u_xpb_out[79][753],u_xpb_out[80][753],u_xpb_out[81][753],u_xpb_out[82][753],u_xpb_out[83][753],u_xpb_out[84][753],u_xpb_out[85][753],u_xpb_out[86][753],u_xpb_out[87][753],u_xpb_out[88][753],u_xpb_out[89][753],u_xpb_out[90][753],u_xpb_out[91][753],u_xpb_out[92][753],u_xpb_out[93][753],u_xpb_out[94][753],u_xpb_out[95][753],u_xpb_out[96][753],u_xpb_out[97][753],u_xpb_out[98][753],u_xpb_out[99][753],u_xpb_out[100][753],u_xpb_out[101][753],u_xpb_out[102][753],u_xpb_out[103][753],u_xpb_out[104][753],u_xpb_out[105][753]};

assign col_out_754 = {u_xpb_out[0][754],u_xpb_out[1][754],u_xpb_out[2][754],u_xpb_out[3][754],u_xpb_out[4][754],u_xpb_out[5][754],u_xpb_out[6][754],u_xpb_out[7][754],u_xpb_out[8][754],u_xpb_out[9][754],u_xpb_out[10][754],u_xpb_out[11][754],u_xpb_out[12][754],u_xpb_out[13][754],u_xpb_out[14][754],u_xpb_out[15][754],u_xpb_out[16][754],u_xpb_out[17][754],u_xpb_out[18][754],u_xpb_out[19][754],u_xpb_out[20][754],u_xpb_out[21][754],u_xpb_out[22][754],u_xpb_out[23][754],u_xpb_out[24][754],u_xpb_out[25][754],u_xpb_out[26][754],u_xpb_out[27][754],u_xpb_out[28][754],u_xpb_out[29][754],u_xpb_out[30][754],u_xpb_out[31][754],u_xpb_out[32][754],u_xpb_out[33][754],u_xpb_out[34][754],u_xpb_out[35][754],u_xpb_out[36][754],u_xpb_out[37][754],u_xpb_out[38][754],u_xpb_out[39][754],u_xpb_out[40][754],u_xpb_out[41][754],u_xpb_out[42][754],u_xpb_out[43][754],u_xpb_out[44][754],u_xpb_out[45][754],u_xpb_out[46][754],u_xpb_out[47][754],u_xpb_out[48][754],u_xpb_out[49][754],u_xpb_out[50][754],u_xpb_out[51][754],u_xpb_out[52][754],u_xpb_out[53][754],u_xpb_out[54][754],u_xpb_out[55][754],u_xpb_out[56][754],u_xpb_out[57][754],u_xpb_out[58][754],u_xpb_out[59][754],u_xpb_out[60][754],u_xpb_out[61][754],u_xpb_out[62][754],u_xpb_out[63][754],u_xpb_out[64][754],u_xpb_out[65][754],u_xpb_out[66][754],u_xpb_out[67][754],u_xpb_out[68][754],u_xpb_out[69][754],u_xpb_out[70][754],u_xpb_out[71][754],u_xpb_out[72][754],u_xpb_out[73][754],u_xpb_out[74][754],u_xpb_out[75][754],u_xpb_out[76][754],u_xpb_out[77][754],u_xpb_out[78][754],u_xpb_out[79][754],u_xpb_out[80][754],u_xpb_out[81][754],u_xpb_out[82][754],u_xpb_out[83][754],u_xpb_out[84][754],u_xpb_out[85][754],u_xpb_out[86][754],u_xpb_out[87][754],u_xpb_out[88][754],u_xpb_out[89][754],u_xpb_out[90][754],u_xpb_out[91][754],u_xpb_out[92][754],u_xpb_out[93][754],u_xpb_out[94][754],u_xpb_out[95][754],u_xpb_out[96][754],u_xpb_out[97][754],u_xpb_out[98][754],u_xpb_out[99][754],u_xpb_out[100][754],u_xpb_out[101][754],u_xpb_out[102][754],u_xpb_out[103][754],u_xpb_out[104][754],u_xpb_out[105][754]};

assign col_out_755 = {u_xpb_out[0][755],u_xpb_out[1][755],u_xpb_out[2][755],u_xpb_out[3][755],u_xpb_out[4][755],u_xpb_out[5][755],u_xpb_out[6][755],u_xpb_out[7][755],u_xpb_out[8][755],u_xpb_out[9][755],u_xpb_out[10][755],u_xpb_out[11][755],u_xpb_out[12][755],u_xpb_out[13][755],u_xpb_out[14][755],u_xpb_out[15][755],u_xpb_out[16][755],u_xpb_out[17][755],u_xpb_out[18][755],u_xpb_out[19][755],u_xpb_out[20][755],u_xpb_out[21][755],u_xpb_out[22][755],u_xpb_out[23][755],u_xpb_out[24][755],u_xpb_out[25][755],u_xpb_out[26][755],u_xpb_out[27][755],u_xpb_out[28][755],u_xpb_out[29][755],u_xpb_out[30][755],u_xpb_out[31][755],u_xpb_out[32][755],u_xpb_out[33][755],u_xpb_out[34][755],u_xpb_out[35][755],u_xpb_out[36][755],u_xpb_out[37][755],u_xpb_out[38][755],u_xpb_out[39][755],u_xpb_out[40][755],u_xpb_out[41][755],u_xpb_out[42][755],u_xpb_out[43][755],u_xpb_out[44][755],u_xpb_out[45][755],u_xpb_out[46][755],u_xpb_out[47][755],u_xpb_out[48][755],u_xpb_out[49][755],u_xpb_out[50][755],u_xpb_out[51][755],u_xpb_out[52][755],u_xpb_out[53][755],u_xpb_out[54][755],u_xpb_out[55][755],u_xpb_out[56][755],u_xpb_out[57][755],u_xpb_out[58][755],u_xpb_out[59][755],u_xpb_out[60][755],u_xpb_out[61][755],u_xpb_out[62][755],u_xpb_out[63][755],u_xpb_out[64][755],u_xpb_out[65][755],u_xpb_out[66][755],u_xpb_out[67][755],u_xpb_out[68][755],u_xpb_out[69][755],u_xpb_out[70][755],u_xpb_out[71][755],u_xpb_out[72][755],u_xpb_out[73][755],u_xpb_out[74][755],u_xpb_out[75][755],u_xpb_out[76][755],u_xpb_out[77][755],u_xpb_out[78][755],u_xpb_out[79][755],u_xpb_out[80][755],u_xpb_out[81][755],u_xpb_out[82][755],u_xpb_out[83][755],u_xpb_out[84][755],u_xpb_out[85][755],u_xpb_out[86][755],u_xpb_out[87][755],u_xpb_out[88][755],u_xpb_out[89][755],u_xpb_out[90][755],u_xpb_out[91][755],u_xpb_out[92][755],u_xpb_out[93][755],u_xpb_out[94][755],u_xpb_out[95][755],u_xpb_out[96][755],u_xpb_out[97][755],u_xpb_out[98][755],u_xpb_out[99][755],u_xpb_out[100][755],u_xpb_out[101][755],u_xpb_out[102][755],u_xpb_out[103][755],u_xpb_out[104][755],u_xpb_out[105][755]};

assign col_out_756 = {u_xpb_out[0][756],u_xpb_out[1][756],u_xpb_out[2][756],u_xpb_out[3][756],u_xpb_out[4][756],u_xpb_out[5][756],u_xpb_out[6][756],u_xpb_out[7][756],u_xpb_out[8][756],u_xpb_out[9][756],u_xpb_out[10][756],u_xpb_out[11][756],u_xpb_out[12][756],u_xpb_out[13][756],u_xpb_out[14][756],u_xpb_out[15][756],u_xpb_out[16][756],u_xpb_out[17][756],u_xpb_out[18][756],u_xpb_out[19][756],u_xpb_out[20][756],u_xpb_out[21][756],u_xpb_out[22][756],u_xpb_out[23][756],u_xpb_out[24][756],u_xpb_out[25][756],u_xpb_out[26][756],u_xpb_out[27][756],u_xpb_out[28][756],u_xpb_out[29][756],u_xpb_out[30][756],u_xpb_out[31][756],u_xpb_out[32][756],u_xpb_out[33][756],u_xpb_out[34][756],u_xpb_out[35][756],u_xpb_out[36][756],u_xpb_out[37][756],u_xpb_out[38][756],u_xpb_out[39][756],u_xpb_out[40][756],u_xpb_out[41][756],u_xpb_out[42][756],u_xpb_out[43][756],u_xpb_out[44][756],u_xpb_out[45][756],u_xpb_out[46][756],u_xpb_out[47][756],u_xpb_out[48][756],u_xpb_out[49][756],u_xpb_out[50][756],u_xpb_out[51][756],u_xpb_out[52][756],u_xpb_out[53][756],u_xpb_out[54][756],u_xpb_out[55][756],u_xpb_out[56][756],u_xpb_out[57][756],u_xpb_out[58][756],u_xpb_out[59][756],u_xpb_out[60][756],u_xpb_out[61][756],u_xpb_out[62][756],u_xpb_out[63][756],u_xpb_out[64][756],u_xpb_out[65][756],u_xpb_out[66][756],u_xpb_out[67][756],u_xpb_out[68][756],u_xpb_out[69][756],u_xpb_out[70][756],u_xpb_out[71][756],u_xpb_out[72][756],u_xpb_out[73][756],u_xpb_out[74][756],u_xpb_out[75][756],u_xpb_out[76][756],u_xpb_out[77][756],u_xpb_out[78][756],u_xpb_out[79][756],u_xpb_out[80][756],u_xpb_out[81][756],u_xpb_out[82][756],u_xpb_out[83][756],u_xpb_out[84][756],u_xpb_out[85][756],u_xpb_out[86][756],u_xpb_out[87][756],u_xpb_out[88][756],u_xpb_out[89][756],u_xpb_out[90][756],u_xpb_out[91][756],u_xpb_out[92][756],u_xpb_out[93][756],u_xpb_out[94][756],u_xpb_out[95][756],u_xpb_out[96][756],u_xpb_out[97][756],u_xpb_out[98][756],u_xpb_out[99][756],u_xpb_out[100][756],u_xpb_out[101][756],u_xpb_out[102][756],u_xpb_out[103][756],u_xpb_out[104][756],u_xpb_out[105][756]};

assign col_out_757 = {u_xpb_out[0][757],u_xpb_out[1][757],u_xpb_out[2][757],u_xpb_out[3][757],u_xpb_out[4][757],u_xpb_out[5][757],u_xpb_out[6][757],u_xpb_out[7][757],u_xpb_out[8][757],u_xpb_out[9][757],u_xpb_out[10][757],u_xpb_out[11][757],u_xpb_out[12][757],u_xpb_out[13][757],u_xpb_out[14][757],u_xpb_out[15][757],u_xpb_out[16][757],u_xpb_out[17][757],u_xpb_out[18][757],u_xpb_out[19][757],u_xpb_out[20][757],u_xpb_out[21][757],u_xpb_out[22][757],u_xpb_out[23][757],u_xpb_out[24][757],u_xpb_out[25][757],u_xpb_out[26][757],u_xpb_out[27][757],u_xpb_out[28][757],u_xpb_out[29][757],u_xpb_out[30][757],u_xpb_out[31][757],u_xpb_out[32][757],u_xpb_out[33][757],u_xpb_out[34][757],u_xpb_out[35][757],u_xpb_out[36][757],u_xpb_out[37][757],u_xpb_out[38][757],u_xpb_out[39][757],u_xpb_out[40][757],u_xpb_out[41][757],u_xpb_out[42][757],u_xpb_out[43][757],u_xpb_out[44][757],u_xpb_out[45][757],u_xpb_out[46][757],u_xpb_out[47][757],u_xpb_out[48][757],u_xpb_out[49][757],u_xpb_out[50][757],u_xpb_out[51][757],u_xpb_out[52][757],u_xpb_out[53][757],u_xpb_out[54][757],u_xpb_out[55][757],u_xpb_out[56][757],u_xpb_out[57][757],u_xpb_out[58][757],u_xpb_out[59][757],u_xpb_out[60][757],u_xpb_out[61][757],u_xpb_out[62][757],u_xpb_out[63][757],u_xpb_out[64][757],u_xpb_out[65][757],u_xpb_out[66][757],u_xpb_out[67][757],u_xpb_out[68][757],u_xpb_out[69][757],u_xpb_out[70][757],u_xpb_out[71][757],u_xpb_out[72][757],u_xpb_out[73][757],u_xpb_out[74][757],u_xpb_out[75][757],u_xpb_out[76][757],u_xpb_out[77][757],u_xpb_out[78][757],u_xpb_out[79][757],u_xpb_out[80][757],u_xpb_out[81][757],u_xpb_out[82][757],u_xpb_out[83][757],u_xpb_out[84][757],u_xpb_out[85][757],u_xpb_out[86][757],u_xpb_out[87][757],u_xpb_out[88][757],u_xpb_out[89][757],u_xpb_out[90][757],u_xpb_out[91][757],u_xpb_out[92][757],u_xpb_out[93][757],u_xpb_out[94][757],u_xpb_out[95][757],u_xpb_out[96][757],u_xpb_out[97][757],u_xpb_out[98][757],u_xpb_out[99][757],u_xpb_out[100][757],u_xpb_out[101][757],u_xpb_out[102][757],u_xpb_out[103][757],u_xpb_out[104][757],u_xpb_out[105][757]};

assign col_out_758 = {u_xpb_out[0][758],u_xpb_out[1][758],u_xpb_out[2][758],u_xpb_out[3][758],u_xpb_out[4][758],u_xpb_out[5][758],u_xpb_out[6][758],u_xpb_out[7][758],u_xpb_out[8][758],u_xpb_out[9][758],u_xpb_out[10][758],u_xpb_out[11][758],u_xpb_out[12][758],u_xpb_out[13][758],u_xpb_out[14][758],u_xpb_out[15][758],u_xpb_out[16][758],u_xpb_out[17][758],u_xpb_out[18][758],u_xpb_out[19][758],u_xpb_out[20][758],u_xpb_out[21][758],u_xpb_out[22][758],u_xpb_out[23][758],u_xpb_out[24][758],u_xpb_out[25][758],u_xpb_out[26][758],u_xpb_out[27][758],u_xpb_out[28][758],u_xpb_out[29][758],u_xpb_out[30][758],u_xpb_out[31][758],u_xpb_out[32][758],u_xpb_out[33][758],u_xpb_out[34][758],u_xpb_out[35][758],u_xpb_out[36][758],u_xpb_out[37][758],u_xpb_out[38][758],u_xpb_out[39][758],u_xpb_out[40][758],u_xpb_out[41][758],u_xpb_out[42][758],u_xpb_out[43][758],u_xpb_out[44][758],u_xpb_out[45][758],u_xpb_out[46][758],u_xpb_out[47][758],u_xpb_out[48][758],u_xpb_out[49][758],u_xpb_out[50][758],u_xpb_out[51][758],u_xpb_out[52][758],u_xpb_out[53][758],u_xpb_out[54][758],u_xpb_out[55][758],u_xpb_out[56][758],u_xpb_out[57][758],u_xpb_out[58][758],u_xpb_out[59][758],u_xpb_out[60][758],u_xpb_out[61][758],u_xpb_out[62][758],u_xpb_out[63][758],u_xpb_out[64][758],u_xpb_out[65][758],u_xpb_out[66][758],u_xpb_out[67][758],u_xpb_out[68][758],u_xpb_out[69][758],u_xpb_out[70][758],u_xpb_out[71][758],u_xpb_out[72][758],u_xpb_out[73][758],u_xpb_out[74][758],u_xpb_out[75][758],u_xpb_out[76][758],u_xpb_out[77][758],u_xpb_out[78][758],u_xpb_out[79][758],u_xpb_out[80][758],u_xpb_out[81][758],u_xpb_out[82][758],u_xpb_out[83][758],u_xpb_out[84][758],u_xpb_out[85][758],u_xpb_out[86][758],u_xpb_out[87][758],u_xpb_out[88][758],u_xpb_out[89][758],u_xpb_out[90][758],u_xpb_out[91][758],u_xpb_out[92][758],u_xpb_out[93][758],u_xpb_out[94][758],u_xpb_out[95][758],u_xpb_out[96][758],u_xpb_out[97][758],u_xpb_out[98][758],u_xpb_out[99][758],u_xpb_out[100][758],u_xpb_out[101][758],u_xpb_out[102][758],u_xpb_out[103][758],u_xpb_out[104][758],u_xpb_out[105][758]};

assign col_out_759 = {u_xpb_out[0][759],u_xpb_out[1][759],u_xpb_out[2][759],u_xpb_out[3][759],u_xpb_out[4][759],u_xpb_out[5][759],u_xpb_out[6][759],u_xpb_out[7][759],u_xpb_out[8][759],u_xpb_out[9][759],u_xpb_out[10][759],u_xpb_out[11][759],u_xpb_out[12][759],u_xpb_out[13][759],u_xpb_out[14][759],u_xpb_out[15][759],u_xpb_out[16][759],u_xpb_out[17][759],u_xpb_out[18][759],u_xpb_out[19][759],u_xpb_out[20][759],u_xpb_out[21][759],u_xpb_out[22][759],u_xpb_out[23][759],u_xpb_out[24][759],u_xpb_out[25][759],u_xpb_out[26][759],u_xpb_out[27][759],u_xpb_out[28][759],u_xpb_out[29][759],u_xpb_out[30][759],u_xpb_out[31][759],u_xpb_out[32][759],u_xpb_out[33][759],u_xpb_out[34][759],u_xpb_out[35][759],u_xpb_out[36][759],u_xpb_out[37][759],u_xpb_out[38][759],u_xpb_out[39][759],u_xpb_out[40][759],u_xpb_out[41][759],u_xpb_out[42][759],u_xpb_out[43][759],u_xpb_out[44][759],u_xpb_out[45][759],u_xpb_out[46][759],u_xpb_out[47][759],u_xpb_out[48][759],u_xpb_out[49][759],u_xpb_out[50][759],u_xpb_out[51][759],u_xpb_out[52][759],u_xpb_out[53][759],u_xpb_out[54][759],u_xpb_out[55][759],u_xpb_out[56][759],u_xpb_out[57][759],u_xpb_out[58][759],u_xpb_out[59][759],u_xpb_out[60][759],u_xpb_out[61][759],u_xpb_out[62][759],u_xpb_out[63][759],u_xpb_out[64][759],u_xpb_out[65][759],u_xpb_out[66][759],u_xpb_out[67][759],u_xpb_out[68][759],u_xpb_out[69][759],u_xpb_out[70][759],u_xpb_out[71][759],u_xpb_out[72][759],u_xpb_out[73][759],u_xpb_out[74][759],u_xpb_out[75][759],u_xpb_out[76][759],u_xpb_out[77][759],u_xpb_out[78][759],u_xpb_out[79][759],u_xpb_out[80][759],u_xpb_out[81][759],u_xpb_out[82][759],u_xpb_out[83][759],u_xpb_out[84][759],u_xpb_out[85][759],u_xpb_out[86][759],u_xpb_out[87][759],u_xpb_out[88][759],u_xpb_out[89][759],u_xpb_out[90][759],u_xpb_out[91][759],u_xpb_out[92][759],u_xpb_out[93][759],u_xpb_out[94][759],u_xpb_out[95][759],u_xpb_out[96][759],u_xpb_out[97][759],u_xpb_out[98][759],u_xpb_out[99][759],u_xpb_out[100][759],u_xpb_out[101][759],u_xpb_out[102][759],u_xpb_out[103][759],u_xpb_out[104][759],u_xpb_out[105][759]};

assign col_out_760 = {u_xpb_out[0][760],u_xpb_out[1][760],u_xpb_out[2][760],u_xpb_out[3][760],u_xpb_out[4][760],u_xpb_out[5][760],u_xpb_out[6][760],u_xpb_out[7][760],u_xpb_out[8][760],u_xpb_out[9][760],u_xpb_out[10][760],u_xpb_out[11][760],u_xpb_out[12][760],u_xpb_out[13][760],u_xpb_out[14][760],u_xpb_out[15][760],u_xpb_out[16][760],u_xpb_out[17][760],u_xpb_out[18][760],u_xpb_out[19][760],u_xpb_out[20][760],u_xpb_out[21][760],u_xpb_out[22][760],u_xpb_out[23][760],u_xpb_out[24][760],u_xpb_out[25][760],u_xpb_out[26][760],u_xpb_out[27][760],u_xpb_out[28][760],u_xpb_out[29][760],u_xpb_out[30][760],u_xpb_out[31][760],u_xpb_out[32][760],u_xpb_out[33][760],u_xpb_out[34][760],u_xpb_out[35][760],u_xpb_out[36][760],u_xpb_out[37][760],u_xpb_out[38][760],u_xpb_out[39][760],u_xpb_out[40][760],u_xpb_out[41][760],u_xpb_out[42][760],u_xpb_out[43][760],u_xpb_out[44][760],u_xpb_out[45][760],u_xpb_out[46][760],u_xpb_out[47][760],u_xpb_out[48][760],u_xpb_out[49][760],u_xpb_out[50][760],u_xpb_out[51][760],u_xpb_out[52][760],u_xpb_out[53][760],u_xpb_out[54][760],u_xpb_out[55][760],u_xpb_out[56][760],u_xpb_out[57][760],u_xpb_out[58][760],u_xpb_out[59][760],u_xpb_out[60][760],u_xpb_out[61][760],u_xpb_out[62][760],u_xpb_out[63][760],u_xpb_out[64][760],u_xpb_out[65][760],u_xpb_out[66][760],u_xpb_out[67][760],u_xpb_out[68][760],u_xpb_out[69][760],u_xpb_out[70][760],u_xpb_out[71][760],u_xpb_out[72][760],u_xpb_out[73][760],u_xpb_out[74][760],u_xpb_out[75][760],u_xpb_out[76][760],u_xpb_out[77][760],u_xpb_out[78][760],u_xpb_out[79][760],u_xpb_out[80][760],u_xpb_out[81][760],u_xpb_out[82][760],u_xpb_out[83][760],u_xpb_out[84][760],u_xpb_out[85][760],u_xpb_out[86][760],u_xpb_out[87][760],u_xpb_out[88][760],u_xpb_out[89][760],u_xpb_out[90][760],u_xpb_out[91][760],u_xpb_out[92][760],u_xpb_out[93][760],u_xpb_out[94][760],u_xpb_out[95][760],u_xpb_out[96][760],u_xpb_out[97][760],u_xpb_out[98][760],u_xpb_out[99][760],u_xpb_out[100][760],u_xpb_out[101][760],u_xpb_out[102][760],u_xpb_out[103][760],u_xpb_out[104][760],u_xpb_out[105][760]};

assign col_out_761 = {u_xpb_out[0][761],u_xpb_out[1][761],u_xpb_out[2][761],u_xpb_out[3][761],u_xpb_out[4][761],u_xpb_out[5][761],u_xpb_out[6][761],u_xpb_out[7][761],u_xpb_out[8][761],u_xpb_out[9][761],u_xpb_out[10][761],u_xpb_out[11][761],u_xpb_out[12][761],u_xpb_out[13][761],u_xpb_out[14][761],u_xpb_out[15][761],u_xpb_out[16][761],u_xpb_out[17][761],u_xpb_out[18][761],u_xpb_out[19][761],u_xpb_out[20][761],u_xpb_out[21][761],u_xpb_out[22][761],u_xpb_out[23][761],u_xpb_out[24][761],u_xpb_out[25][761],u_xpb_out[26][761],u_xpb_out[27][761],u_xpb_out[28][761],u_xpb_out[29][761],u_xpb_out[30][761],u_xpb_out[31][761],u_xpb_out[32][761],u_xpb_out[33][761],u_xpb_out[34][761],u_xpb_out[35][761],u_xpb_out[36][761],u_xpb_out[37][761],u_xpb_out[38][761],u_xpb_out[39][761],u_xpb_out[40][761],u_xpb_out[41][761],u_xpb_out[42][761],u_xpb_out[43][761],u_xpb_out[44][761],u_xpb_out[45][761],u_xpb_out[46][761],u_xpb_out[47][761],u_xpb_out[48][761],u_xpb_out[49][761],u_xpb_out[50][761],u_xpb_out[51][761],u_xpb_out[52][761],u_xpb_out[53][761],u_xpb_out[54][761],u_xpb_out[55][761],u_xpb_out[56][761],u_xpb_out[57][761],u_xpb_out[58][761],u_xpb_out[59][761],u_xpb_out[60][761],u_xpb_out[61][761],u_xpb_out[62][761],u_xpb_out[63][761],u_xpb_out[64][761],u_xpb_out[65][761],u_xpb_out[66][761],u_xpb_out[67][761],u_xpb_out[68][761],u_xpb_out[69][761],u_xpb_out[70][761],u_xpb_out[71][761],u_xpb_out[72][761],u_xpb_out[73][761],u_xpb_out[74][761],u_xpb_out[75][761],u_xpb_out[76][761],u_xpb_out[77][761],u_xpb_out[78][761],u_xpb_out[79][761],u_xpb_out[80][761],u_xpb_out[81][761],u_xpb_out[82][761],u_xpb_out[83][761],u_xpb_out[84][761],u_xpb_out[85][761],u_xpb_out[86][761],u_xpb_out[87][761],u_xpb_out[88][761],u_xpb_out[89][761],u_xpb_out[90][761],u_xpb_out[91][761],u_xpb_out[92][761],u_xpb_out[93][761],u_xpb_out[94][761],u_xpb_out[95][761],u_xpb_out[96][761],u_xpb_out[97][761],u_xpb_out[98][761],u_xpb_out[99][761],u_xpb_out[100][761],u_xpb_out[101][761],u_xpb_out[102][761],u_xpb_out[103][761],u_xpb_out[104][761],u_xpb_out[105][761]};

assign col_out_762 = {u_xpb_out[0][762],u_xpb_out[1][762],u_xpb_out[2][762],u_xpb_out[3][762],u_xpb_out[4][762],u_xpb_out[5][762],u_xpb_out[6][762],u_xpb_out[7][762],u_xpb_out[8][762],u_xpb_out[9][762],u_xpb_out[10][762],u_xpb_out[11][762],u_xpb_out[12][762],u_xpb_out[13][762],u_xpb_out[14][762],u_xpb_out[15][762],u_xpb_out[16][762],u_xpb_out[17][762],u_xpb_out[18][762],u_xpb_out[19][762],u_xpb_out[20][762],u_xpb_out[21][762],u_xpb_out[22][762],u_xpb_out[23][762],u_xpb_out[24][762],u_xpb_out[25][762],u_xpb_out[26][762],u_xpb_out[27][762],u_xpb_out[28][762],u_xpb_out[29][762],u_xpb_out[30][762],u_xpb_out[31][762],u_xpb_out[32][762],u_xpb_out[33][762],u_xpb_out[34][762],u_xpb_out[35][762],u_xpb_out[36][762],u_xpb_out[37][762],u_xpb_out[38][762],u_xpb_out[39][762],u_xpb_out[40][762],u_xpb_out[41][762],u_xpb_out[42][762],u_xpb_out[43][762],u_xpb_out[44][762],u_xpb_out[45][762],u_xpb_out[46][762],u_xpb_out[47][762],u_xpb_out[48][762],u_xpb_out[49][762],u_xpb_out[50][762],u_xpb_out[51][762],u_xpb_out[52][762],u_xpb_out[53][762],u_xpb_out[54][762],u_xpb_out[55][762],u_xpb_out[56][762],u_xpb_out[57][762],u_xpb_out[58][762],u_xpb_out[59][762],u_xpb_out[60][762],u_xpb_out[61][762],u_xpb_out[62][762],u_xpb_out[63][762],u_xpb_out[64][762],u_xpb_out[65][762],u_xpb_out[66][762],u_xpb_out[67][762],u_xpb_out[68][762],u_xpb_out[69][762],u_xpb_out[70][762],u_xpb_out[71][762],u_xpb_out[72][762],u_xpb_out[73][762],u_xpb_out[74][762],u_xpb_out[75][762],u_xpb_out[76][762],u_xpb_out[77][762],u_xpb_out[78][762],u_xpb_out[79][762],u_xpb_out[80][762],u_xpb_out[81][762],u_xpb_out[82][762],u_xpb_out[83][762],u_xpb_out[84][762],u_xpb_out[85][762],u_xpb_out[86][762],u_xpb_out[87][762],u_xpb_out[88][762],u_xpb_out[89][762],u_xpb_out[90][762],u_xpb_out[91][762],u_xpb_out[92][762],u_xpb_out[93][762],u_xpb_out[94][762],u_xpb_out[95][762],u_xpb_out[96][762],u_xpb_out[97][762],u_xpb_out[98][762],u_xpb_out[99][762],u_xpb_out[100][762],u_xpb_out[101][762],u_xpb_out[102][762],u_xpb_out[103][762],u_xpb_out[104][762],u_xpb_out[105][762]};

assign col_out_763 = {u_xpb_out[0][763],u_xpb_out[1][763],u_xpb_out[2][763],u_xpb_out[3][763],u_xpb_out[4][763],u_xpb_out[5][763],u_xpb_out[6][763],u_xpb_out[7][763],u_xpb_out[8][763],u_xpb_out[9][763],u_xpb_out[10][763],u_xpb_out[11][763],u_xpb_out[12][763],u_xpb_out[13][763],u_xpb_out[14][763],u_xpb_out[15][763],u_xpb_out[16][763],u_xpb_out[17][763],u_xpb_out[18][763],u_xpb_out[19][763],u_xpb_out[20][763],u_xpb_out[21][763],u_xpb_out[22][763],u_xpb_out[23][763],u_xpb_out[24][763],u_xpb_out[25][763],u_xpb_out[26][763],u_xpb_out[27][763],u_xpb_out[28][763],u_xpb_out[29][763],u_xpb_out[30][763],u_xpb_out[31][763],u_xpb_out[32][763],u_xpb_out[33][763],u_xpb_out[34][763],u_xpb_out[35][763],u_xpb_out[36][763],u_xpb_out[37][763],u_xpb_out[38][763],u_xpb_out[39][763],u_xpb_out[40][763],u_xpb_out[41][763],u_xpb_out[42][763],u_xpb_out[43][763],u_xpb_out[44][763],u_xpb_out[45][763],u_xpb_out[46][763],u_xpb_out[47][763],u_xpb_out[48][763],u_xpb_out[49][763],u_xpb_out[50][763],u_xpb_out[51][763],u_xpb_out[52][763],u_xpb_out[53][763],u_xpb_out[54][763],u_xpb_out[55][763],u_xpb_out[56][763],u_xpb_out[57][763],u_xpb_out[58][763],u_xpb_out[59][763],u_xpb_out[60][763],u_xpb_out[61][763],u_xpb_out[62][763],u_xpb_out[63][763],u_xpb_out[64][763],u_xpb_out[65][763],u_xpb_out[66][763],u_xpb_out[67][763],u_xpb_out[68][763],u_xpb_out[69][763],u_xpb_out[70][763],u_xpb_out[71][763],u_xpb_out[72][763],u_xpb_out[73][763],u_xpb_out[74][763],u_xpb_out[75][763],u_xpb_out[76][763],u_xpb_out[77][763],u_xpb_out[78][763],u_xpb_out[79][763],u_xpb_out[80][763],u_xpb_out[81][763],u_xpb_out[82][763],u_xpb_out[83][763],u_xpb_out[84][763],u_xpb_out[85][763],u_xpb_out[86][763],u_xpb_out[87][763],u_xpb_out[88][763],u_xpb_out[89][763],u_xpb_out[90][763],u_xpb_out[91][763],u_xpb_out[92][763],u_xpb_out[93][763],u_xpb_out[94][763],u_xpb_out[95][763],u_xpb_out[96][763],u_xpb_out[97][763],u_xpb_out[98][763],u_xpb_out[99][763],u_xpb_out[100][763],u_xpb_out[101][763],u_xpb_out[102][763],u_xpb_out[103][763],u_xpb_out[104][763],u_xpb_out[105][763]};

assign col_out_764 = {u_xpb_out[0][764],u_xpb_out[1][764],u_xpb_out[2][764],u_xpb_out[3][764],u_xpb_out[4][764],u_xpb_out[5][764],u_xpb_out[6][764],u_xpb_out[7][764],u_xpb_out[8][764],u_xpb_out[9][764],u_xpb_out[10][764],u_xpb_out[11][764],u_xpb_out[12][764],u_xpb_out[13][764],u_xpb_out[14][764],u_xpb_out[15][764],u_xpb_out[16][764],u_xpb_out[17][764],u_xpb_out[18][764],u_xpb_out[19][764],u_xpb_out[20][764],u_xpb_out[21][764],u_xpb_out[22][764],u_xpb_out[23][764],u_xpb_out[24][764],u_xpb_out[25][764],u_xpb_out[26][764],u_xpb_out[27][764],u_xpb_out[28][764],u_xpb_out[29][764],u_xpb_out[30][764],u_xpb_out[31][764],u_xpb_out[32][764],u_xpb_out[33][764],u_xpb_out[34][764],u_xpb_out[35][764],u_xpb_out[36][764],u_xpb_out[37][764],u_xpb_out[38][764],u_xpb_out[39][764],u_xpb_out[40][764],u_xpb_out[41][764],u_xpb_out[42][764],u_xpb_out[43][764],u_xpb_out[44][764],u_xpb_out[45][764],u_xpb_out[46][764],u_xpb_out[47][764],u_xpb_out[48][764],u_xpb_out[49][764],u_xpb_out[50][764],u_xpb_out[51][764],u_xpb_out[52][764],u_xpb_out[53][764],u_xpb_out[54][764],u_xpb_out[55][764],u_xpb_out[56][764],u_xpb_out[57][764],u_xpb_out[58][764],u_xpb_out[59][764],u_xpb_out[60][764],u_xpb_out[61][764],u_xpb_out[62][764],u_xpb_out[63][764],u_xpb_out[64][764],u_xpb_out[65][764],u_xpb_out[66][764],u_xpb_out[67][764],u_xpb_out[68][764],u_xpb_out[69][764],u_xpb_out[70][764],u_xpb_out[71][764],u_xpb_out[72][764],u_xpb_out[73][764],u_xpb_out[74][764],u_xpb_out[75][764],u_xpb_out[76][764],u_xpb_out[77][764],u_xpb_out[78][764],u_xpb_out[79][764],u_xpb_out[80][764],u_xpb_out[81][764],u_xpb_out[82][764],u_xpb_out[83][764],u_xpb_out[84][764],u_xpb_out[85][764],u_xpb_out[86][764],u_xpb_out[87][764],u_xpb_out[88][764],u_xpb_out[89][764],u_xpb_out[90][764],u_xpb_out[91][764],u_xpb_out[92][764],u_xpb_out[93][764],u_xpb_out[94][764],u_xpb_out[95][764],u_xpb_out[96][764],u_xpb_out[97][764],u_xpb_out[98][764],u_xpb_out[99][764],u_xpb_out[100][764],u_xpb_out[101][764],u_xpb_out[102][764],u_xpb_out[103][764],u_xpb_out[104][764],u_xpb_out[105][764]};

assign col_out_765 = {u_xpb_out[0][765],u_xpb_out[1][765],u_xpb_out[2][765],u_xpb_out[3][765],u_xpb_out[4][765],u_xpb_out[5][765],u_xpb_out[6][765],u_xpb_out[7][765],u_xpb_out[8][765],u_xpb_out[9][765],u_xpb_out[10][765],u_xpb_out[11][765],u_xpb_out[12][765],u_xpb_out[13][765],u_xpb_out[14][765],u_xpb_out[15][765],u_xpb_out[16][765],u_xpb_out[17][765],u_xpb_out[18][765],u_xpb_out[19][765],u_xpb_out[20][765],u_xpb_out[21][765],u_xpb_out[22][765],u_xpb_out[23][765],u_xpb_out[24][765],u_xpb_out[25][765],u_xpb_out[26][765],u_xpb_out[27][765],u_xpb_out[28][765],u_xpb_out[29][765],u_xpb_out[30][765],u_xpb_out[31][765],u_xpb_out[32][765],u_xpb_out[33][765],u_xpb_out[34][765],u_xpb_out[35][765],u_xpb_out[36][765],u_xpb_out[37][765],u_xpb_out[38][765],u_xpb_out[39][765],u_xpb_out[40][765],u_xpb_out[41][765],u_xpb_out[42][765],u_xpb_out[43][765],u_xpb_out[44][765],u_xpb_out[45][765],u_xpb_out[46][765],u_xpb_out[47][765],u_xpb_out[48][765],u_xpb_out[49][765],u_xpb_out[50][765],u_xpb_out[51][765],u_xpb_out[52][765],u_xpb_out[53][765],u_xpb_out[54][765],u_xpb_out[55][765],u_xpb_out[56][765],u_xpb_out[57][765],u_xpb_out[58][765],u_xpb_out[59][765],u_xpb_out[60][765],u_xpb_out[61][765],u_xpb_out[62][765],u_xpb_out[63][765],u_xpb_out[64][765],u_xpb_out[65][765],u_xpb_out[66][765],u_xpb_out[67][765],u_xpb_out[68][765],u_xpb_out[69][765],u_xpb_out[70][765],u_xpb_out[71][765],u_xpb_out[72][765],u_xpb_out[73][765],u_xpb_out[74][765],u_xpb_out[75][765],u_xpb_out[76][765],u_xpb_out[77][765],u_xpb_out[78][765],u_xpb_out[79][765],u_xpb_out[80][765],u_xpb_out[81][765],u_xpb_out[82][765],u_xpb_out[83][765],u_xpb_out[84][765],u_xpb_out[85][765],u_xpb_out[86][765],u_xpb_out[87][765],u_xpb_out[88][765],u_xpb_out[89][765],u_xpb_out[90][765],u_xpb_out[91][765],u_xpb_out[92][765],u_xpb_out[93][765],u_xpb_out[94][765],u_xpb_out[95][765],u_xpb_out[96][765],u_xpb_out[97][765],u_xpb_out[98][765],u_xpb_out[99][765],u_xpb_out[100][765],u_xpb_out[101][765],u_xpb_out[102][765],u_xpb_out[103][765],u_xpb_out[104][765],u_xpb_out[105][765]};

assign col_out_766 = {u_xpb_out[0][766],u_xpb_out[1][766],u_xpb_out[2][766],u_xpb_out[3][766],u_xpb_out[4][766],u_xpb_out[5][766],u_xpb_out[6][766],u_xpb_out[7][766],u_xpb_out[8][766],u_xpb_out[9][766],u_xpb_out[10][766],u_xpb_out[11][766],u_xpb_out[12][766],u_xpb_out[13][766],u_xpb_out[14][766],u_xpb_out[15][766],u_xpb_out[16][766],u_xpb_out[17][766],u_xpb_out[18][766],u_xpb_out[19][766],u_xpb_out[20][766],u_xpb_out[21][766],u_xpb_out[22][766],u_xpb_out[23][766],u_xpb_out[24][766],u_xpb_out[25][766],u_xpb_out[26][766],u_xpb_out[27][766],u_xpb_out[28][766],u_xpb_out[29][766],u_xpb_out[30][766],u_xpb_out[31][766],u_xpb_out[32][766],u_xpb_out[33][766],u_xpb_out[34][766],u_xpb_out[35][766],u_xpb_out[36][766],u_xpb_out[37][766],u_xpb_out[38][766],u_xpb_out[39][766],u_xpb_out[40][766],u_xpb_out[41][766],u_xpb_out[42][766],u_xpb_out[43][766],u_xpb_out[44][766],u_xpb_out[45][766],u_xpb_out[46][766],u_xpb_out[47][766],u_xpb_out[48][766],u_xpb_out[49][766],u_xpb_out[50][766],u_xpb_out[51][766],u_xpb_out[52][766],u_xpb_out[53][766],u_xpb_out[54][766],u_xpb_out[55][766],u_xpb_out[56][766],u_xpb_out[57][766],u_xpb_out[58][766],u_xpb_out[59][766],u_xpb_out[60][766],u_xpb_out[61][766],u_xpb_out[62][766],u_xpb_out[63][766],u_xpb_out[64][766],u_xpb_out[65][766],u_xpb_out[66][766],u_xpb_out[67][766],u_xpb_out[68][766],u_xpb_out[69][766],u_xpb_out[70][766],u_xpb_out[71][766],u_xpb_out[72][766],u_xpb_out[73][766],u_xpb_out[74][766],u_xpb_out[75][766],u_xpb_out[76][766],u_xpb_out[77][766],u_xpb_out[78][766],u_xpb_out[79][766],u_xpb_out[80][766],u_xpb_out[81][766],u_xpb_out[82][766],u_xpb_out[83][766],u_xpb_out[84][766],u_xpb_out[85][766],u_xpb_out[86][766],u_xpb_out[87][766],u_xpb_out[88][766],u_xpb_out[89][766],u_xpb_out[90][766],u_xpb_out[91][766],u_xpb_out[92][766],u_xpb_out[93][766],u_xpb_out[94][766],u_xpb_out[95][766],u_xpb_out[96][766],u_xpb_out[97][766],u_xpb_out[98][766],u_xpb_out[99][766],u_xpb_out[100][766],u_xpb_out[101][766],u_xpb_out[102][766],u_xpb_out[103][766],u_xpb_out[104][766],u_xpb_out[105][766]};

assign col_out_767 = {u_xpb_out[0][767],u_xpb_out[1][767],u_xpb_out[2][767],u_xpb_out[3][767],u_xpb_out[4][767],u_xpb_out[5][767],u_xpb_out[6][767],u_xpb_out[7][767],u_xpb_out[8][767],u_xpb_out[9][767],u_xpb_out[10][767],u_xpb_out[11][767],u_xpb_out[12][767],u_xpb_out[13][767],u_xpb_out[14][767],u_xpb_out[15][767],u_xpb_out[16][767],u_xpb_out[17][767],u_xpb_out[18][767],u_xpb_out[19][767],u_xpb_out[20][767],u_xpb_out[21][767],u_xpb_out[22][767],u_xpb_out[23][767],u_xpb_out[24][767],u_xpb_out[25][767],u_xpb_out[26][767],u_xpb_out[27][767],u_xpb_out[28][767],u_xpb_out[29][767],u_xpb_out[30][767],u_xpb_out[31][767],u_xpb_out[32][767],u_xpb_out[33][767],u_xpb_out[34][767],u_xpb_out[35][767],u_xpb_out[36][767],u_xpb_out[37][767],u_xpb_out[38][767],u_xpb_out[39][767],u_xpb_out[40][767],u_xpb_out[41][767],u_xpb_out[42][767],u_xpb_out[43][767],u_xpb_out[44][767],u_xpb_out[45][767],u_xpb_out[46][767],u_xpb_out[47][767],u_xpb_out[48][767],u_xpb_out[49][767],u_xpb_out[50][767],u_xpb_out[51][767],u_xpb_out[52][767],u_xpb_out[53][767],u_xpb_out[54][767],u_xpb_out[55][767],u_xpb_out[56][767],u_xpb_out[57][767],u_xpb_out[58][767],u_xpb_out[59][767],u_xpb_out[60][767],u_xpb_out[61][767],u_xpb_out[62][767],u_xpb_out[63][767],u_xpb_out[64][767],u_xpb_out[65][767],u_xpb_out[66][767],u_xpb_out[67][767],u_xpb_out[68][767],u_xpb_out[69][767],u_xpb_out[70][767],u_xpb_out[71][767],u_xpb_out[72][767],u_xpb_out[73][767],u_xpb_out[74][767],u_xpb_out[75][767],u_xpb_out[76][767],u_xpb_out[77][767],u_xpb_out[78][767],u_xpb_out[79][767],u_xpb_out[80][767],u_xpb_out[81][767],u_xpb_out[82][767],u_xpb_out[83][767],u_xpb_out[84][767],u_xpb_out[85][767],u_xpb_out[86][767],u_xpb_out[87][767],u_xpb_out[88][767],u_xpb_out[89][767],u_xpb_out[90][767],u_xpb_out[91][767],u_xpb_out[92][767],u_xpb_out[93][767],u_xpb_out[94][767],u_xpb_out[95][767],u_xpb_out[96][767],u_xpb_out[97][767],u_xpb_out[98][767],u_xpb_out[99][767],u_xpb_out[100][767],u_xpb_out[101][767],u_xpb_out[102][767],u_xpb_out[103][767],u_xpb_out[104][767],u_xpb_out[105][767]};

assign col_out_768 = {u_xpb_out[0][768],u_xpb_out[1][768],u_xpb_out[2][768],u_xpb_out[3][768],u_xpb_out[4][768],u_xpb_out[5][768],u_xpb_out[6][768],u_xpb_out[7][768],u_xpb_out[8][768],u_xpb_out[9][768],u_xpb_out[10][768],u_xpb_out[11][768],u_xpb_out[12][768],u_xpb_out[13][768],u_xpb_out[14][768],u_xpb_out[15][768],u_xpb_out[16][768],u_xpb_out[17][768],u_xpb_out[18][768],u_xpb_out[19][768],u_xpb_out[20][768],u_xpb_out[21][768],u_xpb_out[22][768],u_xpb_out[23][768],u_xpb_out[24][768],u_xpb_out[25][768],u_xpb_out[26][768],u_xpb_out[27][768],u_xpb_out[28][768],u_xpb_out[29][768],u_xpb_out[30][768],u_xpb_out[31][768],u_xpb_out[32][768],u_xpb_out[33][768],u_xpb_out[34][768],u_xpb_out[35][768],u_xpb_out[36][768],u_xpb_out[37][768],u_xpb_out[38][768],u_xpb_out[39][768],u_xpb_out[40][768],u_xpb_out[41][768],u_xpb_out[42][768],u_xpb_out[43][768],u_xpb_out[44][768],u_xpb_out[45][768],u_xpb_out[46][768],u_xpb_out[47][768],u_xpb_out[48][768],u_xpb_out[49][768],u_xpb_out[50][768],u_xpb_out[51][768],u_xpb_out[52][768],u_xpb_out[53][768],u_xpb_out[54][768],u_xpb_out[55][768],u_xpb_out[56][768],u_xpb_out[57][768],u_xpb_out[58][768],u_xpb_out[59][768],u_xpb_out[60][768],u_xpb_out[61][768],u_xpb_out[62][768],u_xpb_out[63][768],u_xpb_out[64][768],u_xpb_out[65][768],u_xpb_out[66][768],u_xpb_out[67][768],u_xpb_out[68][768],u_xpb_out[69][768],u_xpb_out[70][768],u_xpb_out[71][768],u_xpb_out[72][768],u_xpb_out[73][768],u_xpb_out[74][768],u_xpb_out[75][768],u_xpb_out[76][768],u_xpb_out[77][768],u_xpb_out[78][768],u_xpb_out[79][768],u_xpb_out[80][768],u_xpb_out[81][768],u_xpb_out[82][768],u_xpb_out[83][768],u_xpb_out[84][768],u_xpb_out[85][768],u_xpb_out[86][768],u_xpb_out[87][768],u_xpb_out[88][768],u_xpb_out[89][768],u_xpb_out[90][768],u_xpb_out[91][768],u_xpb_out[92][768],u_xpb_out[93][768],u_xpb_out[94][768],u_xpb_out[95][768],u_xpb_out[96][768],u_xpb_out[97][768],u_xpb_out[98][768],u_xpb_out[99][768],u_xpb_out[100][768],u_xpb_out[101][768],u_xpb_out[102][768],u_xpb_out[103][768],u_xpb_out[104][768],u_xpb_out[105][768]};

assign col_out_769 = {u_xpb_out[0][769],u_xpb_out[1][769],u_xpb_out[2][769],u_xpb_out[3][769],u_xpb_out[4][769],u_xpb_out[5][769],u_xpb_out[6][769],u_xpb_out[7][769],u_xpb_out[8][769],u_xpb_out[9][769],u_xpb_out[10][769],u_xpb_out[11][769],u_xpb_out[12][769],u_xpb_out[13][769],u_xpb_out[14][769],u_xpb_out[15][769],u_xpb_out[16][769],u_xpb_out[17][769],u_xpb_out[18][769],u_xpb_out[19][769],u_xpb_out[20][769],u_xpb_out[21][769],u_xpb_out[22][769],u_xpb_out[23][769],u_xpb_out[24][769],u_xpb_out[25][769],u_xpb_out[26][769],u_xpb_out[27][769],u_xpb_out[28][769],u_xpb_out[29][769],u_xpb_out[30][769],u_xpb_out[31][769],u_xpb_out[32][769],u_xpb_out[33][769],u_xpb_out[34][769],u_xpb_out[35][769],u_xpb_out[36][769],u_xpb_out[37][769],u_xpb_out[38][769],u_xpb_out[39][769],u_xpb_out[40][769],u_xpb_out[41][769],u_xpb_out[42][769],u_xpb_out[43][769],u_xpb_out[44][769],u_xpb_out[45][769],u_xpb_out[46][769],u_xpb_out[47][769],u_xpb_out[48][769],u_xpb_out[49][769],u_xpb_out[50][769],u_xpb_out[51][769],u_xpb_out[52][769],u_xpb_out[53][769],u_xpb_out[54][769],u_xpb_out[55][769],u_xpb_out[56][769],u_xpb_out[57][769],u_xpb_out[58][769],u_xpb_out[59][769],u_xpb_out[60][769],u_xpb_out[61][769],u_xpb_out[62][769],u_xpb_out[63][769],u_xpb_out[64][769],u_xpb_out[65][769],u_xpb_out[66][769],u_xpb_out[67][769],u_xpb_out[68][769],u_xpb_out[69][769],u_xpb_out[70][769],u_xpb_out[71][769],u_xpb_out[72][769],u_xpb_out[73][769],u_xpb_out[74][769],u_xpb_out[75][769],u_xpb_out[76][769],u_xpb_out[77][769],u_xpb_out[78][769],u_xpb_out[79][769],u_xpb_out[80][769],u_xpb_out[81][769],u_xpb_out[82][769],u_xpb_out[83][769],u_xpb_out[84][769],u_xpb_out[85][769],u_xpb_out[86][769],u_xpb_out[87][769],u_xpb_out[88][769],u_xpb_out[89][769],u_xpb_out[90][769],u_xpb_out[91][769],u_xpb_out[92][769],u_xpb_out[93][769],u_xpb_out[94][769],u_xpb_out[95][769],u_xpb_out[96][769],u_xpb_out[97][769],u_xpb_out[98][769],u_xpb_out[99][769],u_xpb_out[100][769],u_xpb_out[101][769],u_xpb_out[102][769],u_xpb_out[103][769],u_xpb_out[104][769],u_xpb_out[105][769]};

assign col_out_770 = {u_xpb_out[0][770],u_xpb_out[1][770],u_xpb_out[2][770],u_xpb_out[3][770],u_xpb_out[4][770],u_xpb_out[5][770],u_xpb_out[6][770],u_xpb_out[7][770],u_xpb_out[8][770],u_xpb_out[9][770],u_xpb_out[10][770],u_xpb_out[11][770],u_xpb_out[12][770],u_xpb_out[13][770],u_xpb_out[14][770],u_xpb_out[15][770],u_xpb_out[16][770],u_xpb_out[17][770],u_xpb_out[18][770],u_xpb_out[19][770],u_xpb_out[20][770],u_xpb_out[21][770],u_xpb_out[22][770],u_xpb_out[23][770],u_xpb_out[24][770],u_xpb_out[25][770],u_xpb_out[26][770],u_xpb_out[27][770],u_xpb_out[28][770],u_xpb_out[29][770],u_xpb_out[30][770],u_xpb_out[31][770],u_xpb_out[32][770],u_xpb_out[33][770],u_xpb_out[34][770],u_xpb_out[35][770],u_xpb_out[36][770],u_xpb_out[37][770],u_xpb_out[38][770],u_xpb_out[39][770],u_xpb_out[40][770],u_xpb_out[41][770],u_xpb_out[42][770],u_xpb_out[43][770],u_xpb_out[44][770],u_xpb_out[45][770],u_xpb_out[46][770],u_xpb_out[47][770],u_xpb_out[48][770],u_xpb_out[49][770],u_xpb_out[50][770],u_xpb_out[51][770],u_xpb_out[52][770],u_xpb_out[53][770],u_xpb_out[54][770],u_xpb_out[55][770],u_xpb_out[56][770],u_xpb_out[57][770],u_xpb_out[58][770],u_xpb_out[59][770],u_xpb_out[60][770],u_xpb_out[61][770],u_xpb_out[62][770],u_xpb_out[63][770],u_xpb_out[64][770],u_xpb_out[65][770],u_xpb_out[66][770],u_xpb_out[67][770],u_xpb_out[68][770],u_xpb_out[69][770],u_xpb_out[70][770],u_xpb_out[71][770],u_xpb_out[72][770],u_xpb_out[73][770],u_xpb_out[74][770],u_xpb_out[75][770],u_xpb_out[76][770],u_xpb_out[77][770],u_xpb_out[78][770],u_xpb_out[79][770],u_xpb_out[80][770],u_xpb_out[81][770],u_xpb_out[82][770],u_xpb_out[83][770],u_xpb_out[84][770],u_xpb_out[85][770],u_xpb_out[86][770],u_xpb_out[87][770],u_xpb_out[88][770],u_xpb_out[89][770],u_xpb_out[90][770],u_xpb_out[91][770],u_xpb_out[92][770],u_xpb_out[93][770],u_xpb_out[94][770],u_xpb_out[95][770],u_xpb_out[96][770],u_xpb_out[97][770],u_xpb_out[98][770],u_xpb_out[99][770],u_xpb_out[100][770],u_xpb_out[101][770],u_xpb_out[102][770],u_xpb_out[103][770],u_xpb_out[104][770],u_xpb_out[105][770]};

assign col_out_771 = {u_xpb_out[0][771],u_xpb_out[1][771],u_xpb_out[2][771],u_xpb_out[3][771],u_xpb_out[4][771],u_xpb_out[5][771],u_xpb_out[6][771],u_xpb_out[7][771],u_xpb_out[8][771],u_xpb_out[9][771],u_xpb_out[10][771],u_xpb_out[11][771],u_xpb_out[12][771],u_xpb_out[13][771],u_xpb_out[14][771],u_xpb_out[15][771],u_xpb_out[16][771],u_xpb_out[17][771],u_xpb_out[18][771],u_xpb_out[19][771],u_xpb_out[20][771],u_xpb_out[21][771],u_xpb_out[22][771],u_xpb_out[23][771],u_xpb_out[24][771],u_xpb_out[25][771],u_xpb_out[26][771],u_xpb_out[27][771],u_xpb_out[28][771],u_xpb_out[29][771],u_xpb_out[30][771],u_xpb_out[31][771],u_xpb_out[32][771],u_xpb_out[33][771],u_xpb_out[34][771],u_xpb_out[35][771],u_xpb_out[36][771],u_xpb_out[37][771],u_xpb_out[38][771],u_xpb_out[39][771],u_xpb_out[40][771],u_xpb_out[41][771],u_xpb_out[42][771],u_xpb_out[43][771],u_xpb_out[44][771],u_xpb_out[45][771],u_xpb_out[46][771],u_xpb_out[47][771],u_xpb_out[48][771],u_xpb_out[49][771],u_xpb_out[50][771],u_xpb_out[51][771],u_xpb_out[52][771],u_xpb_out[53][771],u_xpb_out[54][771],u_xpb_out[55][771],u_xpb_out[56][771],u_xpb_out[57][771],u_xpb_out[58][771],u_xpb_out[59][771],u_xpb_out[60][771],u_xpb_out[61][771],u_xpb_out[62][771],u_xpb_out[63][771],u_xpb_out[64][771],u_xpb_out[65][771],u_xpb_out[66][771],u_xpb_out[67][771],u_xpb_out[68][771],u_xpb_out[69][771],u_xpb_out[70][771],u_xpb_out[71][771],u_xpb_out[72][771],u_xpb_out[73][771],u_xpb_out[74][771],u_xpb_out[75][771],u_xpb_out[76][771],u_xpb_out[77][771],u_xpb_out[78][771],u_xpb_out[79][771],u_xpb_out[80][771],u_xpb_out[81][771],u_xpb_out[82][771],u_xpb_out[83][771],u_xpb_out[84][771],u_xpb_out[85][771],u_xpb_out[86][771],u_xpb_out[87][771],u_xpb_out[88][771],u_xpb_out[89][771],u_xpb_out[90][771],u_xpb_out[91][771],u_xpb_out[92][771],u_xpb_out[93][771],u_xpb_out[94][771],u_xpb_out[95][771],u_xpb_out[96][771],u_xpb_out[97][771],u_xpb_out[98][771],u_xpb_out[99][771],u_xpb_out[100][771],u_xpb_out[101][771],u_xpb_out[102][771],u_xpb_out[103][771],u_xpb_out[104][771],u_xpb_out[105][771]};

assign col_out_772 = {u_xpb_out[0][772],u_xpb_out[1][772],u_xpb_out[2][772],u_xpb_out[3][772],u_xpb_out[4][772],u_xpb_out[5][772],u_xpb_out[6][772],u_xpb_out[7][772],u_xpb_out[8][772],u_xpb_out[9][772],u_xpb_out[10][772],u_xpb_out[11][772],u_xpb_out[12][772],u_xpb_out[13][772],u_xpb_out[14][772],u_xpb_out[15][772],u_xpb_out[16][772],u_xpb_out[17][772],u_xpb_out[18][772],u_xpb_out[19][772],u_xpb_out[20][772],u_xpb_out[21][772],u_xpb_out[22][772],u_xpb_out[23][772],u_xpb_out[24][772],u_xpb_out[25][772],u_xpb_out[26][772],u_xpb_out[27][772],u_xpb_out[28][772],u_xpb_out[29][772],u_xpb_out[30][772],u_xpb_out[31][772],u_xpb_out[32][772],u_xpb_out[33][772],u_xpb_out[34][772],u_xpb_out[35][772],u_xpb_out[36][772],u_xpb_out[37][772],u_xpb_out[38][772],u_xpb_out[39][772],u_xpb_out[40][772],u_xpb_out[41][772],u_xpb_out[42][772],u_xpb_out[43][772],u_xpb_out[44][772],u_xpb_out[45][772],u_xpb_out[46][772],u_xpb_out[47][772],u_xpb_out[48][772],u_xpb_out[49][772],u_xpb_out[50][772],u_xpb_out[51][772],u_xpb_out[52][772],u_xpb_out[53][772],u_xpb_out[54][772],u_xpb_out[55][772],u_xpb_out[56][772],u_xpb_out[57][772],u_xpb_out[58][772],u_xpb_out[59][772],u_xpb_out[60][772],u_xpb_out[61][772],u_xpb_out[62][772],u_xpb_out[63][772],u_xpb_out[64][772],u_xpb_out[65][772],u_xpb_out[66][772],u_xpb_out[67][772],u_xpb_out[68][772],u_xpb_out[69][772],u_xpb_out[70][772],u_xpb_out[71][772],u_xpb_out[72][772],u_xpb_out[73][772],u_xpb_out[74][772],u_xpb_out[75][772],u_xpb_out[76][772],u_xpb_out[77][772],u_xpb_out[78][772],u_xpb_out[79][772],u_xpb_out[80][772],u_xpb_out[81][772],u_xpb_out[82][772],u_xpb_out[83][772],u_xpb_out[84][772],u_xpb_out[85][772],u_xpb_out[86][772],u_xpb_out[87][772],u_xpb_out[88][772],u_xpb_out[89][772],u_xpb_out[90][772],u_xpb_out[91][772],u_xpb_out[92][772],u_xpb_out[93][772],u_xpb_out[94][772],u_xpb_out[95][772],u_xpb_out[96][772],u_xpb_out[97][772],u_xpb_out[98][772],u_xpb_out[99][772],u_xpb_out[100][772],u_xpb_out[101][772],u_xpb_out[102][772],u_xpb_out[103][772],u_xpb_out[104][772],u_xpb_out[105][772]};

assign col_out_773 = {u_xpb_out[0][773],u_xpb_out[1][773],u_xpb_out[2][773],u_xpb_out[3][773],u_xpb_out[4][773],u_xpb_out[5][773],u_xpb_out[6][773],u_xpb_out[7][773],u_xpb_out[8][773],u_xpb_out[9][773],u_xpb_out[10][773],u_xpb_out[11][773],u_xpb_out[12][773],u_xpb_out[13][773],u_xpb_out[14][773],u_xpb_out[15][773],u_xpb_out[16][773],u_xpb_out[17][773],u_xpb_out[18][773],u_xpb_out[19][773],u_xpb_out[20][773],u_xpb_out[21][773],u_xpb_out[22][773],u_xpb_out[23][773],u_xpb_out[24][773],u_xpb_out[25][773],u_xpb_out[26][773],u_xpb_out[27][773],u_xpb_out[28][773],u_xpb_out[29][773],u_xpb_out[30][773],u_xpb_out[31][773],u_xpb_out[32][773],u_xpb_out[33][773],u_xpb_out[34][773],u_xpb_out[35][773],u_xpb_out[36][773],u_xpb_out[37][773],u_xpb_out[38][773],u_xpb_out[39][773],u_xpb_out[40][773],u_xpb_out[41][773],u_xpb_out[42][773],u_xpb_out[43][773],u_xpb_out[44][773],u_xpb_out[45][773],u_xpb_out[46][773],u_xpb_out[47][773],u_xpb_out[48][773],u_xpb_out[49][773],u_xpb_out[50][773],u_xpb_out[51][773],u_xpb_out[52][773],u_xpb_out[53][773],u_xpb_out[54][773],u_xpb_out[55][773],u_xpb_out[56][773],u_xpb_out[57][773],u_xpb_out[58][773],u_xpb_out[59][773],u_xpb_out[60][773],u_xpb_out[61][773],u_xpb_out[62][773],u_xpb_out[63][773],u_xpb_out[64][773],u_xpb_out[65][773],u_xpb_out[66][773],u_xpb_out[67][773],u_xpb_out[68][773],u_xpb_out[69][773],u_xpb_out[70][773],u_xpb_out[71][773],u_xpb_out[72][773],u_xpb_out[73][773],u_xpb_out[74][773],u_xpb_out[75][773],u_xpb_out[76][773],u_xpb_out[77][773],u_xpb_out[78][773],u_xpb_out[79][773],u_xpb_out[80][773],u_xpb_out[81][773],u_xpb_out[82][773],u_xpb_out[83][773],u_xpb_out[84][773],u_xpb_out[85][773],u_xpb_out[86][773],u_xpb_out[87][773],u_xpb_out[88][773],u_xpb_out[89][773],u_xpb_out[90][773],u_xpb_out[91][773],u_xpb_out[92][773],u_xpb_out[93][773],u_xpb_out[94][773],u_xpb_out[95][773],u_xpb_out[96][773],u_xpb_out[97][773],u_xpb_out[98][773],u_xpb_out[99][773],u_xpb_out[100][773],u_xpb_out[101][773],u_xpb_out[102][773],u_xpb_out[103][773],u_xpb_out[104][773],u_xpb_out[105][773]};

assign col_out_774 = {u_xpb_out[0][774],u_xpb_out[1][774],u_xpb_out[2][774],u_xpb_out[3][774],u_xpb_out[4][774],u_xpb_out[5][774],u_xpb_out[6][774],u_xpb_out[7][774],u_xpb_out[8][774],u_xpb_out[9][774],u_xpb_out[10][774],u_xpb_out[11][774],u_xpb_out[12][774],u_xpb_out[13][774],u_xpb_out[14][774],u_xpb_out[15][774],u_xpb_out[16][774],u_xpb_out[17][774],u_xpb_out[18][774],u_xpb_out[19][774],u_xpb_out[20][774],u_xpb_out[21][774],u_xpb_out[22][774],u_xpb_out[23][774],u_xpb_out[24][774],u_xpb_out[25][774],u_xpb_out[26][774],u_xpb_out[27][774],u_xpb_out[28][774],u_xpb_out[29][774],u_xpb_out[30][774],u_xpb_out[31][774],u_xpb_out[32][774],u_xpb_out[33][774],u_xpb_out[34][774],u_xpb_out[35][774],u_xpb_out[36][774],u_xpb_out[37][774],u_xpb_out[38][774],u_xpb_out[39][774],u_xpb_out[40][774],u_xpb_out[41][774],u_xpb_out[42][774],u_xpb_out[43][774],u_xpb_out[44][774],u_xpb_out[45][774],u_xpb_out[46][774],u_xpb_out[47][774],u_xpb_out[48][774],u_xpb_out[49][774],u_xpb_out[50][774],u_xpb_out[51][774],u_xpb_out[52][774],u_xpb_out[53][774],u_xpb_out[54][774],u_xpb_out[55][774],u_xpb_out[56][774],u_xpb_out[57][774],u_xpb_out[58][774],u_xpb_out[59][774],u_xpb_out[60][774],u_xpb_out[61][774],u_xpb_out[62][774],u_xpb_out[63][774],u_xpb_out[64][774],u_xpb_out[65][774],u_xpb_out[66][774],u_xpb_out[67][774],u_xpb_out[68][774],u_xpb_out[69][774],u_xpb_out[70][774],u_xpb_out[71][774],u_xpb_out[72][774],u_xpb_out[73][774],u_xpb_out[74][774],u_xpb_out[75][774],u_xpb_out[76][774],u_xpb_out[77][774],u_xpb_out[78][774],u_xpb_out[79][774],u_xpb_out[80][774],u_xpb_out[81][774],u_xpb_out[82][774],u_xpb_out[83][774],u_xpb_out[84][774],u_xpb_out[85][774],u_xpb_out[86][774],u_xpb_out[87][774],u_xpb_out[88][774],u_xpb_out[89][774],u_xpb_out[90][774],u_xpb_out[91][774],u_xpb_out[92][774],u_xpb_out[93][774],u_xpb_out[94][774],u_xpb_out[95][774],u_xpb_out[96][774],u_xpb_out[97][774],u_xpb_out[98][774],u_xpb_out[99][774],u_xpb_out[100][774],u_xpb_out[101][774],u_xpb_out[102][774],u_xpb_out[103][774],u_xpb_out[104][774],u_xpb_out[105][774]};

assign col_out_775 = {u_xpb_out[0][775],u_xpb_out[1][775],u_xpb_out[2][775],u_xpb_out[3][775],u_xpb_out[4][775],u_xpb_out[5][775],u_xpb_out[6][775],u_xpb_out[7][775],u_xpb_out[8][775],u_xpb_out[9][775],u_xpb_out[10][775],u_xpb_out[11][775],u_xpb_out[12][775],u_xpb_out[13][775],u_xpb_out[14][775],u_xpb_out[15][775],u_xpb_out[16][775],u_xpb_out[17][775],u_xpb_out[18][775],u_xpb_out[19][775],u_xpb_out[20][775],u_xpb_out[21][775],u_xpb_out[22][775],u_xpb_out[23][775],u_xpb_out[24][775],u_xpb_out[25][775],u_xpb_out[26][775],u_xpb_out[27][775],u_xpb_out[28][775],u_xpb_out[29][775],u_xpb_out[30][775],u_xpb_out[31][775],u_xpb_out[32][775],u_xpb_out[33][775],u_xpb_out[34][775],u_xpb_out[35][775],u_xpb_out[36][775],u_xpb_out[37][775],u_xpb_out[38][775],u_xpb_out[39][775],u_xpb_out[40][775],u_xpb_out[41][775],u_xpb_out[42][775],u_xpb_out[43][775],u_xpb_out[44][775],u_xpb_out[45][775],u_xpb_out[46][775],u_xpb_out[47][775],u_xpb_out[48][775],u_xpb_out[49][775],u_xpb_out[50][775],u_xpb_out[51][775],u_xpb_out[52][775],u_xpb_out[53][775],u_xpb_out[54][775],u_xpb_out[55][775],u_xpb_out[56][775],u_xpb_out[57][775],u_xpb_out[58][775],u_xpb_out[59][775],u_xpb_out[60][775],u_xpb_out[61][775],u_xpb_out[62][775],u_xpb_out[63][775],u_xpb_out[64][775],u_xpb_out[65][775],u_xpb_out[66][775],u_xpb_out[67][775],u_xpb_out[68][775],u_xpb_out[69][775],u_xpb_out[70][775],u_xpb_out[71][775],u_xpb_out[72][775],u_xpb_out[73][775],u_xpb_out[74][775],u_xpb_out[75][775],u_xpb_out[76][775],u_xpb_out[77][775],u_xpb_out[78][775],u_xpb_out[79][775],u_xpb_out[80][775],u_xpb_out[81][775],u_xpb_out[82][775],u_xpb_out[83][775],u_xpb_out[84][775],u_xpb_out[85][775],u_xpb_out[86][775],u_xpb_out[87][775],u_xpb_out[88][775],u_xpb_out[89][775],u_xpb_out[90][775],u_xpb_out[91][775],u_xpb_out[92][775],u_xpb_out[93][775],u_xpb_out[94][775],u_xpb_out[95][775],u_xpb_out[96][775],u_xpb_out[97][775],u_xpb_out[98][775],u_xpb_out[99][775],u_xpb_out[100][775],u_xpb_out[101][775],u_xpb_out[102][775],u_xpb_out[103][775],u_xpb_out[104][775],u_xpb_out[105][775]};

assign col_out_776 = {u_xpb_out[0][776],u_xpb_out[1][776],u_xpb_out[2][776],u_xpb_out[3][776],u_xpb_out[4][776],u_xpb_out[5][776],u_xpb_out[6][776],u_xpb_out[7][776],u_xpb_out[8][776],u_xpb_out[9][776],u_xpb_out[10][776],u_xpb_out[11][776],u_xpb_out[12][776],u_xpb_out[13][776],u_xpb_out[14][776],u_xpb_out[15][776],u_xpb_out[16][776],u_xpb_out[17][776],u_xpb_out[18][776],u_xpb_out[19][776],u_xpb_out[20][776],u_xpb_out[21][776],u_xpb_out[22][776],u_xpb_out[23][776],u_xpb_out[24][776],u_xpb_out[25][776],u_xpb_out[26][776],u_xpb_out[27][776],u_xpb_out[28][776],u_xpb_out[29][776],u_xpb_out[30][776],u_xpb_out[31][776],u_xpb_out[32][776],u_xpb_out[33][776],u_xpb_out[34][776],u_xpb_out[35][776],u_xpb_out[36][776],u_xpb_out[37][776],u_xpb_out[38][776],u_xpb_out[39][776],u_xpb_out[40][776],u_xpb_out[41][776],u_xpb_out[42][776],u_xpb_out[43][776],u_xpb_out[44][776],u_xpb_out[45][776],u_xpb_out[46][776],u_xpb_out[47][776],u_xpb_out[48][776],u_xpb_out[49][776],u_xpb_out[50][776],u_xpb_out[51][776],u_xpb_out[52][776],u_xpb_out[53][776],u_xpb_out[54][776],u_xpb_out[55][776],u_xpb_out[56][776],u_xpb_out[57][776],u_xpb_out[58][776],u_xpb_out[59][776],u_xpb_out[60][776],u_xpb_out[61][776],u_xpb_out[62][776],u_xpb_out[63][776],u_xpb_out[64][776],u_xpb_out[65][776],u_xpb_out[66][776],u_xpb_out[67][776],u_xpb_out[68][776],u_xpb_out[69][776],u_xpb_out[70][776],u_xpb_out[71][776],u_xpb_out[72][776],u_xpb_out[73][776],u_xpb_out[74][776],u_xpb_out[75][776],u_xpb_out[76][776],u_xpb_out[77][776],u_xpb_out[78][776],u_xpb_out[79][776],u_xpb_out[80][776],u_xpb_out[81][776],u_xpb_out[82][776],u_xpb_out[83][776],u_xpb_out[84][776],u_xpb_out[85][776],u_xpb_out[86][776],u_xpb_out[87][776],u_xpb_out[88][776],u_xpb_out[89][776],u_xpb_out[90][776],u_xpb_out[91][776],u_xpb_out[92][776],u_xpb_out[93][776],u_xpb_out[94][776],u_xpb_out[95][776],u_xpb_out[96][776],u_xpb_out[97][776],u_xpb_out[98][776],u_xpb_out[99][776],u_xpb_out[100][776],u_xpb_out[101][776],u_xpb_out[102][776],u_xpb_out[103][776],u_xpb_out[104][776],u_xpb_out[105][776]};

assign col_out_777 = {u_xpb_out[0][777],u_xpb_out[1][777],u_xpb_out[2][777],u_xpb_out[3][777],u_xpb_out[4][777],u_xpb_out[5][777],u_xpb_out[6][777],u_xpb_out[7][777],u_xpb_out[8][777],u_xpb_out[9][777],u_xpb_out[10][777],u_xpb_out[11][777],u_xpb_out[12][777],u_xpb_out[13][777],u_xpb_out[14][777],u_xpb_out[15][777],u_xpb_out[16][777],u_xpb_out[17][777],u_xpb_out[18][777],u_xpb_out[19][777],u_xpb_out[20][777],u_xpb_out[21][777],u_xpb_out[22][777],u_xpb_out[23][777],u_xpb_out[24][777],u_xpb_out[25][777],u_xpb_out[26][777],u_xpb_out[27][777],u_xpb_out[28][777],u_xpb_out[29][777],u_xpb_out[30][777],u_xpb_out[31][777],u_xpb_out[32][777],u_xpb_out[33][777],u_xpb_out[34][777],u_xpb_out[35][777],u_xpb_out[36][777],u_xpb_out[37][777],u_xpb_out[38][777],u_xpb_out[39][777],u_xpb_out[40][777],u_xpb_out[41][777],u_xpb_out[42][777],u_xpb_out[43][777],u_xpb_out[44][777],u_xpb_out[45][777],u_xpb_out[46][777],u_xpb_out[47][777],u_xpb_out[48][777],u_xpb_out[49][777],u_xpb_out[50][777],u_xpb_out[51][777],u_xpb_out[52][777],u_xpb_out[53][777],u_xpb_out[54][777],u_xpb_out[55][777],u_xpb_out[56][777],u_xpb_out[57][777],u_xpb_out[58][777],u_xpb_out[59][777],u_xpb_out[60][777],u_xpb_out[61][777],u_xpb_out[62][777],u_xpb_out[63][777],u_xpb_out[64][777],u_xpb_out[65][777],u_xpb_out[66][777],u_xpb_out[67][777],u_xpb_out[68][777],u_xpb_out[69][777],u_xpb_out[70][777],u_xpb_out[71][777],u_xpb_out[72][777],u_xpb_out[73][777],u_xpb_out[74][777],u_xpb_out[75][777],u_xpb_out[76][777],u_xpb_out[77][777],u_xpb_out[78][777],u_xpb_out[79][777],u_xpb_out[80][777],u_xpb_out[81][777],u_xpb_out[82][777],u_xpb_out[83][777],u_xpb_out[84][777],u_xpb_out[85][777],u_xpb_out[86][777],u_xpb_out[87][777],u_xpb_out[88][777],u_xpb_out[89][777],u_xpb_out[90][777],u_xpb_out[91][777],u_xpb_out[92][777],u_xpb_out[93][777],u_xpb_out[94][777],u_xpb_out[95][777],u_xpb_out[96][777],u_xpb_out[97][777],u_xpb_out[98][777],u_xpb_out[99][777],u_xpb_out[100][777],u_xpb_out[101][777],u_xpb_out[102][777],u_xpb_out[103][777],u_xpb_out[104][777],u_xpb_out[105][777]};

assign col_out_778 = {u_xpb_out[0][778],u_xpb_out[1][778],u_xpb_out[2][778],u_xpb_out[3][778],u_xpb_out[4][778],u_xpb_out[5][778],u_xpb_out[6][778],u_xpb_out[7][778],u_xpb_out[8][778],u_xpb_out[9][778],u_xpb_out[10][778],u_xpb_out[11][778],u_xpb_out[12][778],u_xpb_out[13][778],u_xpb_out[14][778],u_xpb_out[15][778],u_xpb_out[16][778],u_xpb_out[17][778],u_xpb_out[18][778],u_xpb_out[19][778],u_xpb_out[20][778],u_xpb_out[21][778],u_xpb_out[22][778],u_xpb_out[23][778],u_xpb_out[24][778],u_xpb_out[25][778],u_xpb_out[26][778],u_xpb_out[27][778],u_xpb_out[28][778],u_xpb_out[29][778],u_xpb_out[30][778],u_xpb_out[31][778],u_xpb_out[32][778],u_xpb_out[33][778],u_xpb_out[34][778],u_xpb_out[35][778],u_xpb_out[36][778],u_xpb_out[37][778],u_xpb_out[38][778],u_xpb_out[39][778],u_xpb_out[40][778],u_xpb_out[41][778],u_xpb_out[42][778],u_xpb_out[43][778],u_xpb_out[44][778],u_xpb_out[45][778],u_xpb_out[46][778],u_xpb_out[47][778],u_xpb_out[48][778],u_xpb_out[49][778],u_xpb_out[50][778],u_xpb_out[51][778],u_xpb_out[52][778],u_xpb_out[53][778],u_xpb_out[54][778],u_xpb_out[55][778],u_xpb_out[56][778],u_xpb_out[57][778],u_xpb_out[58][778],u_xpb_out[59][778],u_xpb_out[60][778],u_xpb_out[61][778],u_xpb_out[62][778],u_xpb_out[63][778],u_xpb_out[64][778],u_xpb_out[65][778],u_xpb_out[66][778],u_xpb_out[67][778],u_xpb_out[68][778],u_xpb_out[69][778],u_xpb_out[70][778],u_xpb_out[71][778],u_xpb_out[72][778],u_xpb_out[73][778],u_xpb_out[74][778],u_xpb_out[75][778],u_xpb_out[76][778],u_xpb_out[77][778],u_xpb_out[78][778],u_xpb_out[79][778],u_xpb_out[80][778],u_xpb_out[81][778],u_xpb_out[82][778],u_xpb_out[83][778],u_xpb_out[84][778],u_xpb_out[85][778],u_xpb_out[86][778],u_xpb_out[87][778],u_xpb_out[88][778],u_xpb_out[89][778],u_xpb_out[90][778],u_xpb_out[91][778],u_xpb_out[92][778],u_xpb_out[93][778],u_xpb_out[94][778],u_xpb_out[95][778],u_xpb_out[96][778],u_xpb_out[97][778],u_xpb_out[98][778],u_xpb_out[99][778],u_xpb_out[100][778],u_xpb_out[101][778],u_xpb_out[102][778],u_xpb_out[103][778],u_xpb_out[104][778],u_xpb_out[105][778]};

assign col_out_779 = {u_xpb_out[0][779],u_xpb_out[1][779],u_xpb_out[2][779],u_xpb_out[3][779],u_xpb_out[4][779],u_xpb_out[5][779],u_xpb_out[6][779],u_xpb_out[7][779],u_xpb_out[8][779],u_xpb_out[9][779],u_xpb_out[10][779],u_xpb_out[11][779],u_xpb_out[12][779],u_xpb_out[13][779],u_xpb_out[14][779],u_xpb_out[15][779],u_xpb_out[16][779],u_xpb_out[17][779],u_xpb_out[18][779],u_xpb_out[19][779],u_xpb_out[20][779],u_xpb_out[21][779],u_xpb_out[22][779],u_xpb_out[23][779],u_xpb_out[24][779],u_xpb_out[25][779],u_xpb_out[26][779],u_xpb_out[27][779],u_xpb_out[28][779],u_xpb_out[29][779],u_xpb_out[30][779],u_xpb_out[31][779],u_xpb_out[32][779],u_xpb_out[33][779],u_xpb_out[34][779],u_xpb_out[35][779],u_xpb_out[36][779],u_xpb_out[37][779],u_xpb_out[38][779],u_xpb_out[39][779],u_xpb_out[40][779],u_xpb_out[41][779],u_xpb_out[42][779],u_xpb_out[43][779],u_xpb_out[44][779],u_xpb_out[45][779],u_xpb_out[46][779],u_xpb_out[47][779],u_xpb_out[48][779],u_xpb_out[49][779],u_xpb_out[50][779],u_xpb_out[51][779],u_xpb_out[52][779],u_xpb_out[53][779],u_xpb_out[54][779],u_xpb_out[55][779],u_xpb_out[56][779],u_xpb_out[57][779],u_xpb_out[58][779],u_xpb_out[59][779],u_xpb_out[60][779],u_xpb_out[61][779],u_xpb_out[62][779],u_xpb_out[63][779],u_xpb_out[64][779],u_xpb_out[65][779],u_xpb_out[66][779],u_xpb_out[67][779],u_xpb_out[68][779],u_xpb_out[69][779],u_xpb_out[70][779],u_xpb_out[71][779],u_xpb_out[72][779],u_xpb_out[73][779],u_xpb_out[74][779],u_xpb_out[75][779],u_xpb_out[76][779],u_xpb_out[77][779],u_xpb_out[78][779],u_xpb_out[79][779],u_xpb_out[80][779],u_xpb_out[81][779],u_xpb_out[82][779],u_xpb_out[83][779],u_xpb_out[84][779],u_xpb_out[85][779],u_xpb_out[86][779],u_xpb_out[87][779],u_xpb_out[88][779],u_xpb_out[89][779],u_xpb_out[90][779],u_xpb_out[91][779],u_xpb_out[92][779],u_xpb_out[93][779],u_xpb_out[94][779],u_xpb_out[95][779],u_xpb_out[96][779],u_xpb_out[97][779],u_xpb_out[98][779],u_xpb_out[99][779],u_xpb_out[100][779],u_xpb_out[101][779],u_xpb_out[102][779],u_xpb_out[103][779],u_xpb_out[104][779],u_xpb_out[105][779]};

assign col_out_780 = {u_xpb_out[0][780],u_xpb_out[1][780],u_xpb_out[2][780],u_xpb_out[3][780],u_xpb_out[4][780],u_xpb_out[5][780],u_xpb_out[6][780],u_xpb_out[7][780],u_xpb_out[8][780],u_xpb_out[9][780],u_xpb_out[10][780],u_xpb_out[11][780],u_xpb_out[12][780],u_xpb_out[13][780],u_xpb_out[14][780],u_xpb_out[15][780],u_xpb_out[16][780],u_xpb_out[17][780],u_xpb_out[18][780],u_xpb_out[19][780],u_xpb_out[20][780],u_xpb_out[21][780],u_xpb_out[22][780],u_xpb_out[23][780],u_xpb_out[24][780],u_xpb_out[25][780],u_xpb_out[26][780],u_xpb_out[27][780],u_xpb_out[28][780],u_xpb_out[29][780],u_xpb_out[30][780],u_xpb_out[31][780],u_xpb_out[32][780],u_xpb_out[33][780],u_xpb_out[34][780],u_xpb_out[35][780],u_xpb_out[36][780],u_xpb_out[37][780],u_xpb_out[38][780],u_xpb_out[39][780],u_xpb_out[40][780],u_xpb_out[41][780],u_xpb_out[42][780],u_xpb_out[43][780],u_xpb_out[44][780],u_xpb_out[45][780],u_xpb_out[46][780],u_xpb_out[47][780],u_xpb_out[48][780],u_xpb_out[49][780],u_xpb_out[50][780],u_xpb_out[51][780],u_xpb_out[52][780],u_xpb_out[53][780],u_xpb_out[54][780],u_xpb_out[55][780],u_xpb_out[56][780],u_xpb_out[57][780],u_xpb_out[58][780],u_xpb_out[59][780],u_xpb_out[60][780],u_xpb_out[61][780],u_xpb_out[62][780],u_xpb_out[63][780],u_xpb_out[64][780],u_xpb_out[65][780],u_xpb_out[66][780],u_xpb_out[67][780],u_xpb_out[68][780],u_xpb_out[69][780],u_xpb_out[70][780],u_xpb_out[71][780],u_xpb_out[72][780],u_xpb_out[73][780],u_xpb_out[74][780],u_xpb_out[75][780],u_xpb_out[76][780],u_xpb_out[77][780],u_xpb_out[78][780],u_xpb_out[79][780],u_xpb_out[80][780],u_xpb_out[81][780],u_xpb_out[82][780],u_xpb_out[83][780],u_xpb_out[84][780],u_xpb_out[85][780],u_xpb_out[86][780],u_xpb_out[87][780],u_xpb_out[88][780],u_xpb_out[89][780],u_xpb_out[90][780],u_xpb_out[91][780],u_xpb_out[92][780],u_xpb_out[93][780],u_xpb_out[94][780],u_xpb_out[95][780],u_xpb_out[96][780],u_xpb_out[97][780],u_xpb_out[98][780],u_xpb_out[99][780],u_xpb_out[100][780],u_xpb_out[101][780],u_xpb_out[102][780],u_xpb_out[103][780],u_xpb_out[104][780],u_xpb_out[105][780]};

assign col_out_781 = {u_xpb_out[0][781],u_xpb_out[1][781],u_xpb_out[2][781],u_xpb_out[3][781],u_xpb_out[4][781],u_xpb_out[5][781],u_xpb_out[6][781],u_xpb_out[7][781],u_xpb_out[8][781],u_xpb_out[9][781],u_xpb_out[10][781],u_xpb_out[11][781],u_xpb_out[12][781],u_xpb_out[13][781],u_xpb_out[14][781],u_xpb_out[15][781],u_xpb_out[16][781],u_xpb_out[17][781],u_xpb_out[18][781],u_xpb_out[19][781],u_xpb_out[20][781],u_xpb_out[21][781],u_xpb_out[22][781],u_xpb_out[23][781],u_xpb_out[24][781],u_xpb_out[25][781],u_xpb_out[26][781],u_xpb_out[27][781],u_xpb_out[28][781],u_xpb_out[29][781],u_xpb_out[30][781],u_xpb_out[31][781],u_xpb_out[32][781],u_xpb_out[33][781],u_xpb_out[34][781],u_xpb_out[35][781],u_xpb_out[36][781],u_xpb_out[37][781],u_xpb_out[38][781],u_xpb_out[39][781],u_xpb_out[40][781],u_xpb_out[41][781],u_xpb_out[42][781],u_xpb_out[43][781],u_xpb_out[44][781],u_xpb_out[45][781],u_xpb_out[46][781],u_xpb_out[47][781],u_xpb_out[48][781],u_xpb_out[49][781],u_xpb_out[50][781],u_xpb_out[51][781],u_xpb_out[52][781],u_xpb_out[53][781],u_xpb_out[54][781],u_xpb_out[55][781],u_xpb_out[56][781],u_xpb_out[57][781],u_xpb_out[58][781],u_xpb_out[59][781],u_xpb_out[60][781],u_xpb_out[61][781],u_xpb_out[62][781],u_xpb_out[63][781],u_xpb_out[64][781],u_xpb_out[65][781],u_xpb_out[66][781],u_xpb_out[67][781],u_xpb_out[68][781],u_xpb_out[69][781],u_xpb_out[70][781],u_xpb_out[71][781],u_xpb_out[72][781],u_xpb_out[73][781],u_xpb_out[74][781],u_xpb_out[75][781],u_xpb_out[76][781],u_xpb_out[77][781],u_xpb_out[78][781],u_xpb_out[79][781],u_xpb_out[80][781],u_xpb_out[81][781],u_xpb_out[82][781],u_xpb_out[83][781],u_xpb_out[84][781],u_xpb_out[85][781],u_xpb_out[86][781],u_xpb_out[87][781],u_xpb_out[88][781],u_xpb_out[89][781],u_xpb_out[90][781],u_xpb_out[91][781],u_xpb_out[92][781],u_xpb_out[93][781],u_xpb_out[94][781],u_xpb_out[95][781],u_xpb_out[96][781],u_xpb_out[97][781],u_xpb_out[98][781],u_xpb_out[99][781],u_xpb_out[100][781],u_xpb_out[101][781],u_xpb_out[102][781],u_xpb_out[103][781],u_xpb_out[104][781],u_xpb_out[105][781]};

assign col_out_782 = {u_xpb_out[0][782],u_xpb_out[1][782],u_xpb_out[2][782],u_xpb_out[3][782],u_xpb_out[4][782],u_xpb_out[5][782],u_xpb_out[6][782],u_xpb_out[7][782],u_xpb_out[8][782],u_xpb_out[9][782],u_xpb_out[10][782],u_xpb_out[11][782],u_xpb_out[12][782],u_xpb_out[13][782],u_xpb_out[14][782],u_xpb_out[15][782],u_xpb_out[16][782],u_xpb_out[17][782],u_xpb_out[18][782],u_xpb_out[19][782],u_xpb_out[20][782],u_xpb_out[21][782],u_xpb_out[22][782],u_xpb_out[23][782],u_xpb_out[24][782],u_xpb_out[25][782],u_xpb_out[26][782],u_xpb_out[27][782],u_xpb_out[28][782],u_xpb_out[29][782],u_xpb_out[30][782],u_xpb_out[31][782],u_xpb_out[32][782],u_xpb_out[33][782],u_xpb_out[34][782],u_xpb_out[35][782],u_xpb_out[36][782],u_xpb_out[37][782],u_xpb_out[38][782],u_xpb_out[39][782],u_xpb_out[40][782],u_xpb_out[41][782],u_xpb_out[42][782],u_xpb_out[43][782],u_xpb_out[44][782],u_xpb_out[45][782],u_xpb_out[46][782],u_xpb_out[47][782],u_xpb_out[48][782],u_xpb_out[49][782],u_xpb_out[50][782],u_xpb_out[51][782],u_xpb_out[52][782],u_xpb_out[53][782],u_xpb_out[54][782],u_xpb_out[55][782],u_xpb_out[56][782],u_xpb_out[57][782],u_xpb_out[58][782],u_xpb_out[59][782],u_xpb_out[60][782],u_xpb_out[61][782],u_xpb_out[62][782],u_xpb_out[63][782],u_xpb_out[64][782],u_xpb_out[65][782],u_xpb_out[66][782],u_xpb_out[67][782],u_xpb_out[68][782],u_xpb_out[69][782],u_xpb_out[70][782],u_xpb_out[71][782],u_xpb_out[72][782],u_xpb_out[73][782],u_xpb_out[74][782],u_xpb_out[75][782],u_xpb_out[76][782],u_xpb_out[77][782],u_xpb_out[78][782],u_xpb_out[79][782],u_xpb_out[80][782],u_xpb_out[81][782],u_xpb_out[82][782],u_xpb_out[83][782],u_xpb_out[84][782],u_xpb_out[85][782],u_xpb_out[86][782],u_xpb_out[87][782],u_xpb_out[88][782],u_xpb_out[89][782],u_xpb_out[90][782],u_xpb_out[91][782],u_xpb_out[92][782],u_xpb_out[93][782],u_xpb_out[94][782],u_xpb_out[95][782],u_xpb_out[96][782],u_xpb_out[97][782],u_xpb_out[98][782],u_xpb_out[99][782],u_xpb_out[100][782],u_xpb_out[101][782],u_xpb_out[102][782],u_xpb_out[103][782],u_xpb_out[104][782],u_xpb_out[105][782]};

assign col_out_783 = {u_xpb_out[0][783],u_xpb_out[1][783],u_xpb_out[2][783],u_xpb_out[3][783],u_xpb_out[4][783],u_xpb_out[5][783],u_xpb_out[6][783],u_xpb_out[7][783],u_xpb_out[8][783],u_xpb_out[9][783],u_xpb_out[10][783],u_xpb_out[11][783],u_xpb_out[12][783],u_xpb_out[13][783],u_xpb_out[14][783],u_xpb_out[15][783],u_xpb_out[16][783],u_xpb_out[17][783],u_xpb_out[18][783],u_xpb_out[19][783],u_xpb_out[20][783],u_xpb_out[21][783],u_xpb_out[22][783],u_xpb_out[23][783],u_xpb_out[24][783],u_xpb_out[25][783],u_xpb_out[26][783],u_xpb_out[27][783],u_xpb_out[28][783],u_xpb_out[29][783],u_xpb_out[30][783],u_xpb_out[31][783],u_xpb_out[32][783],u_xpb_out[33][783],u_xpb_out[34][783],u_xpb_out[35][783],u_xpb_out[36][783],u_xpb_out[37][783],u_xpb_out[38][783],u_xpb_out[39][783],u_xpb_out[40][783],u_xpb_out[41][783],u_xpb_out[42][783],u_xpb_out[43][783],u_xpb_out[44][783],u_xpb_out[45][783],u_xpb_out[46][783],u_xpb_out[47][783],u_xpb_out[48][783],u_xpb_out[49][783],u_xpb_out[50][783],u_xpb_out[51][783],u_xpb_out[52][783],u_xpb_out[53][783],u_xpb_out[54][783],u_xpb_out[55][783],u_xpb_out[56][783],u_xpb_out[57][783],u_xpb_out[58][783],u_xpb_out[59][783],u_xpb_out[60][783],u_xpb_out[61][783],u_xpb_out[62][783],u_xpb_out[63][783],u_xpb_out[64][783],u_xpb_out[65][783],u_xpb_out[66][783],u_xpb_out[67][783],u_xpb_out[68][783],u_xpb_out[69][783],u_xpb_out[70][783],u_xpb_out[71][783],u_xpb_out[72][783],u_xpb_out[73][783],u_xpb_out[74][783],u_xpb_out[75][783],u_xpb_out[76][783],u_xpb_out[77][783],u_xpb_out[78][783],u_xpb_out[79][783],u_xpb_out[80][783],u_xpb_out[81][783],u_xpb_out[82][783],u_xpb_out[83][783],u_xpb_out[84][783],u_xpb_out[85][783],u_xpb_out[86][783],u_xpb_out[87][783],u_xpb_out[88][783],u_xpb_out[89][783],u_xpb_out[90][783],u_xpb_out[91][783],u_xpb_out[92][783],u_xpb_out[93][783],u_xpb_out[94][783],u_xpb_out[95][783],u_xpb_out[96][783],u_xpb_out[97][783],u_xpb_out[98][783],u_xpb_out[99][783],u_xpb_out[100][783],u_xpb_out[101][783],u_xpb_out[102][783],u_xpb_out[103][783],u_xpb_out[104][783],u_xpb_out[105][783]};

assign col_out_784 = {u_xpb_out[0][784],u_xpb_out[1][784],u_xpb_out[2][784],u_xpb_out[3][784],u_xpb_out[4][784],u_xpb_out[5][784],u_xpb_out[6][784],u_xpb_out[7][784],u_xpb_out[8][784],u_xpb_out[9][784],u_xpb_out[10][784],u_xpb_out[11][784],u_xpb_out[12][784],u_xpb_out[13][784],u_xpb_out[14][784],u_xpb_out[15][784],u_xpb_out[16][784],u_xpb_out[17][784],u_xpb_out[18][784],u_xpb_out[19][784],u_xpb_out[20][784],u_xpb_out[21][784],u_xpb_out[22][784],u_xpb_out[23][784],u_xpb_out[24][784],u_xpb_out[25][784],u_xpb_out[26][784],u_xpb_out[27][784],u_xpb_out[28][784],u_xpb_out[29][784],u_xpb_out[30][784],u_xpb_out[31][784],u_xpb_out[32][784],u_xpb_out[33][784],u_xpb_out[34][784],u_xpb_out[35][784],u_xpb_out[36][784],u_xpb_out[37][784],u_xpb_out[38][784],u_xpb_out[39][784],u_xpb_out[40][784],u_xpb_out[41][784],u_xpb_out[42][784],u_xpb_out[43][784],u_xpb_out[44][784],u_xpb_out[45][784],u_xpb_out[46][784],u_xpb_out[47][784],u_xpb_out[48][784],u_xpb_out[49][784],u_xpb_out[50][784],u_xpb_out[51][784],u_xpb_out[52][784],u_xpb_out[53][784],u_xpb_out[54][784],u_xpb_out[55][784],u_xpb_out[56][784],u_xpb_out[57][784],u_xpb_out[58][784],u_xpb_out[59][784],u_xpb_out[60][784],u_xpb_out[61][784],u_xpb_out[62][784],u_xpb_out[63][784],u_xpb_out[64][784],u_xpb_out[65][784],u_xpb_out[66][784],u_xpb_out[67][784],u_xpb_out[68][784],u_xpb_out[69][784],u_xpb_out[70][784],u_xpb_out[71][784],u_xpb_out[72][784],u_xpb_out[73][784],u_xpb_out[74][784],u_xpb_out[75][784],u_xpb_out[76][784],u_xpb_out[77][784],u_xpb_out[78][784],u_xpb_out[79][784],u_xpb_out[80][784],u_xpb_out[81][784],u_xpb_out[82][784],u_xpb_out[83][784],u_xpb_out[84][784],u_xpb_out[85][784],u_xpb_out[86][784],u_xpb_out[87][784],u_xpb_out[88][784],u_xpb_out[89][784],u_xpb_out[90][784],u_xpb_out[91][784],u_xpb_out[92][784],u_xpb_out[93][784],u_xpb_out[94][784],u_xpb_out[95][784],u_xpb_out[96][784],u_xpb_out[97][784],u_xpb_out[98][784],u_xpb_out[99][784],u_xpb_out[100][784],u_xpb_out[101][784],u_xpb_out[102][784],u_xpb_out[103][784],u_xpb_out[104][784],u_xpb_out[105][784]};

assign col_out_785 = {u_xpb_out[0][785],u_xpb_out[1][785],u_xpb_out[2][785],u_xpb_out[3][785],u_xpb_out[4][785],u_xpb_out[5][785],u_xpb_out[6][785],u_xpb_out[7][785],u_xpb_out[8][785],u_xpb_out[9][785],u_xpb_out[10][785],u_xpb_out[11][785],u_xpb_out[12][785],u_xpb_out[13][785],u_xpb_out[14][785],u_xpb_out[15][785],u_xpb_out[16][785],u_xpb_out[17][785],u_xpb_out[18][785],u_xpb_out[19][785],u_xpb_out[20][785],u_xpb_out[21][785],u_xpb_out[22][785],u_xpb_out[23][785],u_xpb_out[24][785],u_xpb_out[25][785],u_xpb_out[26][785],u_xpb_out[27][785],u_xpb_out[28][785],u_xpb_out[29][785],u_xpb_out[30][785],u_xpb_out[31][785],u_xpb_out[32][785],u_xpb_out[33][785],u_xpb_out[34][785],u_xpb_out[35][785],u_xpb_out[36][785],u_xpb_out[37][785],u_xpb_out[38][785],u_xpb_out[39][785],u_xpb_out[40][785],u_xpb_out[41][785],u_xpb_out[42][785],u_xpb_out[43][785],u_xpb_out[44][785],u_xpb_out[45][785],u_xpb_out[46][785],u_xpb_out[47][785],u_xpb_out[48][785],u_xpb_out[49][785],u_xpb_out[50][785],u_xpb_out[51][785],u_xpb_out[52][785],u_xpb_out[53][785],u_xpb_out[54][785],u_xpb_out[55][785],u_xpb_out[56][785],u_xpb_out[57][785],u_xpb_out[58][785],u_xpb_out[59][785],u_xpb_out[60][785],u_xpb_out[61][785],u_xpb_out[62][785],u_xpb_out[63][785],u_xpb_out[64][785],u_xpb_out[65][785],u_xpb_out[66][785],u_xpb_out[67][785],u_xpb_out[68][785],u_xpb_out[69][785],u_xpb_out[70][785],u_xpb_out[71][785],u_xpb_out[72][785],u_xpb_out[73][785],u_xpb_out[74][785],u_xpb_out[75][785],u_xpb_out[76][785],u_xpb_out[77][785],u_xpb_out[78][785],u_xpb_out[79][785],u_xpb_out[80][785],u_xpb_out[81][785],u_xpb_out[82][785],u_xpb_out[83][785],u_xpb_out[84][785],u_xpb_out[85][785],u_xpb_out[86][785],u_xpb_out[87][785],u_xpb_out[88][785],u_xpb_out[89][785],u_xpb_out[90][785],u_xpb_out[91][785],u_xpb_out[92][785],u_xpb_out[93][785],u_xpb_out[94][785],u_xpb_out[95][785],u_xpb_out[96][785],u_xpb_out[97][785],u_xpb_out[98][785],u_xpb_out[99][785],u_xpb_out[100][785],u_xpb_out[101][785],u_xpb_out[102][785],u_xpb_out[103][785],u_xpb_out[104][785],u_xpb_out[105][785]};

assign col_out_786 = {u_xpb_out[0][786],u_xpb_out[1][786],u_xpb_out[2][786],u_xpb_out[3][786],u_xpb_out[4][786],u_xpb_out[5][786],u_xpb_out[6][786],u_xpb_out[7][786],u_xpb_out[8][786],u_xpb_out[9][786],u_xpb_out[10][786],u_xpb_out[11][786],u_xpb_out[12][786],u_xpb_out[13][786],u_xpb_out[14][786],u_xpb_out[15][786],u_xpb_out[16][786],u_xpb_out[17][786],u_xpb_out[18][786],u_xpb_out[19][786],u_xpb_out[20][786],u_xpb_out[21][786],u_xpb_out[22][786],u_xpb_out[23][786],u_xpb_out[24][786],u_xpb_out[25][786],u_xpb_out[26][786],u_xpb_out[27][786],u_xpb_out[28][786],u_xpb_out[29][786],u_xpb_out[30][786],u_xpb_out[31][786],u_xpb_out[32][786],u_xpb_out[33][786],u_xpb_out[34][786],u_xpb_out[35][786],u_xpb_out[36][786],u_xpb_out[37][786],u_xpb_out[38][786],u_xpb_out[39][786],u_xpb_out[40][786],u_xpb_out[41][786],u_xpb_out[42][786],u_xpb_out[43][786],u_xpb_out[44][786],u_xpb_out[45][786],u_xpb_out[46][786],u_xpb_out[47][786],u_xpb_out[48][786],u_xpb_out[49][786],u_xpb_out[50][786],u_xpb_out[51][786],u_xpb_out[52][786],u_xpb_out[53][786],u_xpb_out[54][786],u_xpb_out[55][786],u_xpb_out[56][786],u_xpb_out[57][786],u_xpb_out[58][786],u_xpb_out[59][786],u_xpb_out[60][786],u_xpb_out[61][786],u_xpb_out[62][786],u_xpb_out[63][786],u_xpb_out[64][786],u_xpb_out[65][786],u_xpb_out[66][786],u_xpb_out[67][786],u_xpb_out[68][786],u_xpb_out[69][786],u_xpb_out[70][786],u_xpb_out[71][786],u_xpb_out[72][786],u_xpb_out[73][786],u_xpb_out[74][786],u_xpb_out[75][786],u_xpb_out[76][786],u_xpb_out[77][786],u_xpb_out[78][786],u_xpb_out[79][786],u_xpb_out[80][786],u_xpb_out[81][786],u_xpb_out[82][786],u_xpb_out[83][786],u_xpb_out[84][786],u_xpb_out[85][786],u_xpb_out[86][786],u_xpb_out[87][786],u_xpb_out[88][786],u_xpb_out[89][786],u_xpb_out[90][786],u_xpb_out[91][786],u_xpb_out[92][786],u_xpb_out[93][786],u_xpb_out[94][786],u_xpb_out[95][786],u_xpb_out[96][786],u_xpb_out[97][786],u_xpb_out[98][786],u_xpb_out[99][786],u_xpb_out[100][786],u_xpb_out[101][786],u_xpb_out[102][786],u_xpb_out[103][786],u_xpb_out[104][786],u_xpb_out[105][786]};

assign col_out_787 = {u_xpb_out[0][787],u_xpb_out[1][787],u_xpb_out[2][787],u_xpb_out[3][787],u_xpb_out[4][787],u_xpb_out[5][787],u_xpb_out[6][787],u_xpb_out[7][787],u_xpb_out[8][787],u_xpb_out[9][787],u_xpb_out[10][787],u_xpb_out[11][787],u_xpb_out[12][787],u_xpb_out[13][787],u_xpb_out[14][787],u_xpb_out[15][787],u_xpb_out[16][787],u_xpb_out[17][787],u_xpb_out[18][787],u_xpb_out[19][787],u_xpb_out[20][787],u_xpb_out[21][787],u_xpb_out[22][787],u_xpb_out[23][787],u_xpb_out[24][787],u_xpb_out[25][787],u_xpb_out[26][787],u_xpb_out[27][787],u_xpb_out[28][787],u_xpb_out[29][787],u_xpb_out[30][787],u_xpb_out[31][787],u_xpb_out[32][787],u_xpb_out[33][787],u_xpb_out[34][787],u_xpb_out[35][787],u_xpb_out[36][787],u_xpb_out[37][787],u_xpb_out[38][787],u_xpb_out[39][787],u_xpb_out[40][787],u_xpb_out[41][787],u_xpb_out[42][787],u_xpb_out[43][787],u_xpb_out[44][787],u_xpb_out[45][787],u_xpb_out[46][787],u_xpb_out[47][787],u_xpb_out[48][787],u_xpb_out[49][787],u_xpb_out[50][787],u_xpb_out[51][787],u_xpb_out[52][787],u_xpb_out[53][787],u_xpb_out[54][787],u_xpb_out[55][787],u_xpb_out[56][787],u_xpb_out[57][787],u_xpb_out[58][787],u_xpb_out[59][787],u_xpb_out[60][787],u_xpb_out[61][787],u_xpb_out[62][787],u_xpb_out[63][787],u_xpb_out[64][787],u_xpb_out[65][787],u_xpb_out[66][787],u_xpb_out[67][787],u_xpb_out[68][787],u_xpb_out[69][787],u_xpb_out[70][787],u_xpb_out[71][787],u_xpb_out[72][787],u_xpb_out[73][787],u_xpb_out[74][787],u_xpb_out[75][787],u_xpb_out[76][787],u_xpb_out[77][787],u_xpb_out[78][787],u_xpb_out[79][787],u_xpb_out[80][787],u_xpb_out[81][787],u_xpb_out[82][787],u_xpb_out[83][787],u_xpb_out[84][787],u_xpb_out[85][787],u_xpb_out[86][787],u_xpb_out[87][787],u_xpb_out[88][787],u_xpb_out[89][787],u_xpb_out[90][787],u_xpb_out[91][787],u_xpb_out[92][787],u_xpb_out[93][787],u_xpb_out[94][787],u_xpb_out[95][787],u_xpb_out[96][787],u_xpb_out[97][787],u_xpb_out[98][787],u_xpb_out[99][787],u_xpb_out[100][787],u_xpb_out[101][787],u_xpb_out[102][787],u_xpb_out[103][787],u_xpb_out[104][787],u_xpb_out[105][787]};

assign col_out_788 = {u_xpb_out[0][788],u_xpb_out[1][788],u_xpb_out[2][788],u_xpb_out[3][788],u_xpb_out[4][788],u_xpb_out[5][788],u_xpb_out[6][788],u_xpb_out[7][788],u_xpb_out[8][788],u_xpb_out[9][788],u_xpb_out[10][788],u_xpb_out[11][788],u_xpb_out[12][788],u_xpb_out[13][788],u_xpb_out[14][788],u_xpb_out[15][788],u_xpb_out[16][788],u_xpb_out[17][788],u_xpb_out[18][788],u_xpb_out[19][788],u_xpb_out[20][788],u_xpb_out[21][788],u_xpb_out[22][788],u_xpb_out[23][788],u_xpb_out[24][788],u_xpb_out[25][788],u_xpb_out[26][788],u_xpb_out[27][788],u_xpb_out[28][788],u_xpb_out[29][788],u_xpb_out[30][788],u_xpb_out[31][788],u_xpb_out[32][788],u_xpb_out[33][788],u_xpb_out[34][788],u_xpb_out[35][788],u_xpb_out[36][788],u_xpb_out[37][788],u_xpb_out[38][788],u_xpb_out[39][788],u_xpb_out[40][788],u_xpb_out[41][788],u_xpb_out[42][788],u_xpb_out[43][788],u_xpb_out[44][788],u_xpb_out[45][788],u_xpb_out[46][788],u_xpb_out[47][788],u_xpb_out[48][788],u_xpb_out[49][788],u_xpb_out[50][788],u_xpb_out[51][788],u_xpb_out[52][788],u_xpb_out[53][788],u_xpb_out[54][788],u_xpb_out[55][788],u_xpb_out[56][788],u_xpb_out[57][788],u_xpb_out[58][788],u_xpb_out[59][788],u_xpb_out[60][788],u_xpb_out[61][788],u_xpb_out[62][788],u_xpb_out[63][788],u_xpb_out[64][788],u_xpb_out[65][788],u_xpb_out[66][788],u_xpb_out[67][788],u_xpb_out[68][788],u_xpb_out[69][788],u_xpb_out[70][788],u_xpb_out[71][788],u_xpb_out[72][788],u_xpb_out[73][788],u_xpb_out[74][788],u_xpb_out[75][788],u_xpb_out[76][788],u_xpb_out[77][788],u_xpb_out[78][788],u_xpb_out[79][788],u_xpb_out[80][788],u_xpb_out[81][788],u_xpb_out[82][788],u_xpb_out[83][788],u_xpb_out[84][788],u_xpb_out[85][788],u_xpb_out[86][788],u_xpb_out[87][788],u_xpb_out[88][788],u_xpb_out[89][788],u_xpb_out[90][788],u_xpb_out[91][788],u_xpb_out[92][788],u_xpb_out[93][788],u_xpb_out[94][788],u_xpb_out[95][788],u_xpb_out[96][788],u_xpb_out[97][788],u_xpb_out[98][788],u_xpb_out[99][788],u_xpb_out[100][788],u_xpb_out[101][788],u_xpb_out[102][788],u_xpb_out[103][788],u_xpb_out[104][788],u_xpb_out[105][788]};

assign col_out_789 = {u_xpb_out[0][789],u_xpb_out[1][789],u_xpb_out[2][789],u_xpb_out[3][789],u_xpb_out[4][789],u_xpb_out[5][789],u_xpb_out[6][789],u_xpb_out[7][789],u_xpb_out[8][789],u_xpb_out[9][789],u_xpb_out[10][789],u_xpb_out[11][789],u_xpb_out[12][789],u_xpb_out[13][789],u_xpb_out[14][789],u_xpb_out[15][789],u_xpb_out[16][789],u_xpb_out[17][789],u_xpb_out[18][789],u_xpb_out[19][789],u_xpb_out[20][789],u_xpb_out[21][789],u_xpb_out[22][789],u_xpb_out[23][789],u_xpb_out[24][789],u_xpb_out[25][789],u_xpb_out[26][789],u_xpb_out[27][789],u_xpb_out[28][789],u_xpb_out[29][789],u_xpb_out[30][789],u_xpb_out[31][789],u_xpb_out[32][789],u_xpb_out[33][789],u_xpb_out[34][789],u_xpb_out[35][789],u_xpb_out[36][789],u_xpb_out[37][789],u_xpb_out[38][789],u_xpb_out[39][789],u_xpb_out[40][789],u_xpb_out[41][789],u_xpb_out[42][789],u_xpb_out[43][789],u_xpb_out[44][789],u_xpb_out[45][789],u_xpb_out[46][789],u_xpb_out[47][789],u_xpb_out[48][789],u_xpb_out[49][789],u_xpb_out[50][789],u_xpb_out[51][789],u_xpb_out[52][789],u_xpb_out[53][789],u_xpb_out[54][789],u_xpb_out[55][789],u_xpb_out[56][789],u_xpb_out[57][789],u_xpb_out[58][789],u_xpb_out[59][789],u_xpb_out[60][789],u_xpb_out[61][789],u_xpb_out[62][789],u_xpb_out[63][789],u_xpb_out[64][789],u_xpb_out[65][789],u_xpb_out[66][789],u_xpb_out[67][789],u_xpb_out[68][789],u_xpb_out[69][789],u_xpb_out[70][789],u_xpb_out[71][789],u_xpb_out[72][789],u_xpb_out[73][789],u_xpb_out[74][789],u_xpb_out[75][789],u_xpb_out[76][789],u_xpb_out[77][789],u_xpb_out[78][789],u_xpb_out[79][789],u_xpb_out[80][789],u_xpb_out[81][789],u_xpb_out[82][789],u_xpb_out[83][789],u_xpb_out[84][789],u_xpb_out[85][789],u_xpb_out[86][789],u_xpb_out[87][789],u_xpb_out[88][789],u_xpb_out[89][789],u_xpb_out[90][789],u_xpb_out[91][789],u_xpb_out[92][789],u_xpb_out[93][789],u_xpb_out[94][789],u_xpb_out[95][789],u_xpb_out[96][789],u_xpb_out[97][789],u_xpb_out[98][789],u_xpb_out[99][789],u_xpb_out[100][789],u_xpb_out[101][789],u_xpb_out[102][789],u_xpb_out[103][789],u_xpb_out[104][789],u_xpb_out[105][789]};

assign col_out_790 = {u_xpb_out[0][790],u_xpb_out[1][790],u_xpb_out[2][790],u_xpb_out[3][790],u_xpb_out[4][790],u_xpb_out[5][790],u_xpb_out[6][790],u_xpb_out[7][790],u_xpb_out[8][790],u_xpb_out[9][790],u_xpb_out[10][790],u_xpb_out[11][790],u_xpb_out[12][790],u_xpb_out[13][790],u_xpb_out[14][790],u_xpb_out[15][790],u_xpb_out[16][790],u_xpb_out[17][790],u_xpb_out[18][790],u_xpb_out[19][790],u_xpb_out[20][790],u_xpb_out[21][790],u_xpb_out[22][790],u_xpb_out[23][790],u_xpb_out[24][790],u_xpb_out[25][790],u_xpb_out[26][790],u_xpb_out[27][790],u_xpb_out[28][790],u_xpb_out[29][790],u_xpb_out[30][790],u_xpb_out[31][790],u_xpb_out[32][790],u_xpb_out[33][790],u_xpb_out[34][790],u_xpb_out[35][790],u_xpb_out[36][790],u_xpb_out[37][790],u_xpb_out[38][790],u_xpb_out[39][790],u_xpb_out[40][790],u_xpb_out[41][790],u_xpb_out[42][790],u_xpb_out[43][790],u_xpb_out[44][790],u_xpb_out[45][790],u_xpb_out[46][790],u_xpb_out[47][790],u_xpb_out[48][790],u_xpb_out[49][790],u_xpb_out[50][790],u_xpb_out[51][790],u_xpb_out[52][790],u_xpb_out[53][790],u_xpb_out[54][790],u_xpb_out[55][790],u_xpb_out[56][790],u_xpb_out[57][790],u_xpb_out[58][790],u_xpb_out[59][790],u_xpb_out[60][790],u_xpb_out[61][790],u_xpb_out[62][790],u_xpb_out[63][790],u_xpb_out[64][790],u_xpb_out[65][790],u_xpb_out[66][790],u_xpb_out[67][790],u_xpb_out[68][790],u_xpb_out[69][790],u_xpb_out[70][790],u_xpb_out[71][790],u_xpb_out[72][790],u_xpb_out[73][790],u_xpb_out[74][790],u_xpb_out[75][790],u_xpb_out[76][790],u_xpb_out[77][790],u_xpb_out[78][790],u_xpb_out[79][790],u_xpb_out[80][790],u_xpb_out[81][790],u_xpb_out[82][790],u_xpb_out[83][790],u_xpb_out[84][790],u_xpb_out[85][790],u_xpb_out[86][790],u_xpb_out[87][790],u_xpb_out[88][790],u_xpb_out[89][790],u_xpb_out[90][790],u_xpb_out[91][790],u_xpb_out[92][790],u_xpb_out[93][790],u_xpb_out[94][790],u_xpb_out[95][790],u_xpb_out[96][790],u_xpb_out[97][790],u_xpb_out[98][790],u_xpb_out[99][790],u_xpb_out[100][790],u_xpb_out[101][790],u_xpb_out[102][790],u_xpb_out[103][790],u_xpb_out[104][790],u_xpb_out[105][790]};

assign col_out_791 = {u_xpb_out[0][791],u_xpb_out[1][791],u_xpb_out[2][791],u_xpb_out[3][791],u_xpb_out[4][791],u_xpb_out[5][791],u_xpb_out[6][791],u_xpb_out[7][791],u_xpb_out[8][791],u_xpb_out[9][791],u_xpb_out[10][791],u_xpb_out[11][791],u_xpb_out[12][791],u_xpb_out[13][791],u_xpb_out[14][791],u_xpb_out[15][791],u_xpb_out[16][791],u_xpb_out[17][791],u_xpb_out[18][791],u_xpb_out[19][791],u_xpb_out[20][791],u_xpb_out[21][791],u_xpb_out[22][791],u_xpb_out[23][791],u_xpb_out[24][791],u_xpb_out[25][791],u_xpb_out[26][791],u_xpb_out[27][791],u_xpb_out[28][791],u_xpb_out[29][791],u_xpb_out[30][791],u_xpb_out[31][791],u_xpb_out[32][791],u_xpb_out[33][791],u_xpb_out[34][791],u_xpb_out[35][791],u_xpb_out[36][791],u_xpb_out[37][791],u_xpb_out[38][791],u_xpb_out[39][791],u_xpb_out[40][791],u_xpb_out[41][791],u_xpb_out[42][791],u_xpb_out[43][791],u_xpb_out[44][791],u_xpb_out[45][791],u_xpb_out[46][791],u_xpb_out[47][791],u_xpb_out[48][791],u_xpb_out[49][791],u_xpb_out[50][791],u_xpb_out[51][791],u_xpb_out[52][791],u_xpb_out[53][791],u_xpb_out[54][791],u_xpb_out[55][791],u_xpb_out[56][791],u_xpb_out[57][791],u_xpb_out[58][791],u_xpb_out[59][791],u_xpb_out[60][791],u_xpb_out[61][791],u_xpb_out[62][791],u_xpb_out[63][791],u_xpb_out[64][791],u_xpb_out[65][791],u_xpb_out[66][791],u_xpb_out[67][791],u_xpb_out[68][791],u_xpb_out[69][791],u_xpb_out[70][791],u_xpb_out[71][791],u_xpb_out[72][791],u_xpb_out[73][791],u_xpb_out[74][791],u_xpb_out[75][791],u_xpb_out[76][791],u_xpb_out[77][791],u_xpb_out[78][791],u_xpb_out[79][791],u_xpb_out[80][791],u_xpb_out[81][791],u_xpb_out[82][791],u_xpb_out[83][791],u_xpb_out[84][791],u_xpb_out[85][791],u_xpb_out[86][791],u_xpb_out[87][791],u_xpb_out[88][791],u_xpb_out[89][791],u_xpb_out[90][791],u_xpb_out[91][791],u_xpb_out[92][791],u_xpb_out[93][791],u_xpb_out[94][791],u_xpb_out[95][791],u_xpb_out[96][791],u_xpb_out[97][791],u_xpb_out[98][791],u_xpb_out[99][791],u_xpb_out[100][791],u_xpb_out[101][791],u_xpb_out[102][791],u_xpb_out[103][791],u_xpb_out[104][791],u_xpb_out[105][791]};

assign col_out_792 = {u_xpb_out[0][792],u_xpb_out[1][792],u_xpb_out[2][792],u_xpb_out[3][792],u_xpb_out[4][792],u_xpb_out[5][792],u_xpb_out[6][792],u_xpb_out[7][792],u_xpb_out[8][792],u_xpb_out[9][792],u_xpb_out[10][792],u_xpb_out[11][792],u_xpb_out[12][792],u_xpb_out[13][792],u_xpb_out[14][792],u_xpb_out[15][792],u_xpb_out[16][792],u_xpb_out[17][792],u_xpb_out[18][792],u_xpb_out[19][792],u_xpb_out[20][792],u_xpb_out[21][792],u_xpb_out[22][792],u_xpb_out[23][792],u_xpb_out[24][792],u_xpb_out[25][792],u_xpb_out[26][792],u_xpb_out[27][792],u_xpb_out[28][792],u_xpb_out[29][792],u_xpb_out[30][792],u_xpb_out[31][792],u_xpb_out[32][792],u_xpb_out[33][792],u_xpb_out[34][792],u_xpb_out[35][792],u_xpb_out[36][792],u_xpb_out[37][792],u_xpb_out[38][792],u_xpb_out[39][792],u_xpb_out[40][792],u_xpb_out[41][792],u_xpb_out[42][792],u_xpb_out[43][792],u_xpb_out[44][792],u_xpb_out[45][792],u_xpb_out[46][792],u_xpb_out[47][792],u_xpb_out[48][792],u_xpb_out[49][792],u_xpb_out[50][792],u_xpb_out[51][792],u_xpb_out[52][792],u_xpb_out[53][792],u_xpb_out[54][792],u_xpb_out[55][792],u_xpb_out[56][792],u_xpb_out[57][792],u_xpb_out[58][792],u_xpb_out[59][792],u_xpb_out[60][792],u_xpb_out[61][792],u_xpb_out[62][792],u_xpb_out[63][792],u_xpb_out[64][792],u_xpb_out[65][792],u_xpb_out[66][792],u_xpb_out[67][792],u_xpb_out[68][792],u_xpb_out[69][792],u_xpb_out[70][792],u_xpb_out[71][792],u_xpb_out[72][792],u_xpb_out[73][792],u_xpb_out[74][792],u_xpb_out[75][792],u_xpb_out[76][792],u_xpb_out[77][792],u_xpb_out[78][792],u_xpb_out[79][792],u_xpb_out[80][792],u_xpb_out[81][792],u_xpb_out[82][792],u_xpb_out[83][792],u_xpb_out[84][792],u_xpb_out[85][792],u_xpb_out[86][792],u_xpb_out[87][792],u_xpb_out[88][792],u_xpb_out[89][792],u_xpb_out[90][792],u_xpb_out[91][792],u_xpb_out[92][792],u_xpb_out[93][792],u_xpb_out[94][792],u_xpb_out[95][792],u_xpb_out[96][792],u_xpb_out[97][792],u_xpb_out[98][792],u_xpb_out[99][792],u_xpb_out[100][792],u_xpb_out[101][792],u_xpb_out[102][792],u_xpb_out[103][792],u_xpb_out[104][792],u_xpb_out[105][792]};

assign col_out_793 = {u_xpb_out[0][793],u_xpb_out[1][793],u_xpb_out[2][793],u_xpb_out[3][793],u_xpb_out[4][793],u_xpb_out[5][793],u_xpb_out[6][793],u_xpb_out[7][793],u_xpb_out[8][793],u_xpb_out[9][793],u_xpb_out[10][793],u_xpb_out[11][793],u_xpb_out[12][793],u_xpb_out[13][793],u_xpb_out[14][793],u_xpb_out[15][793],u_xpb_out[16][793],u_xpb_out[17][793],u_xpb_out[18][793],u_xpb_out[19][793],u_xpb_out[20][793],u_xpb_out[21][793],u_xpb_out[22][793],u_xpb_out[23][793],u_xpb_out[24][793],u_xpb_out[25][793],u_xpb_out[26][793],u_xpb_out[27][793],u_xpb_out[28][793],u_xpb_out[29][793],u_xpb_out[30][793],u_xpb_out[31][793],u_xpb_out[32][793],u_xpb_out[33][793],u_xpb_out[34][793],u_xpb_out[35][793],u_xpb_out[36][793],u_xpb_out[37][793],u_xpb_out[38][793],u_xpb_out[39][793],u_xpb_out[40][793],u_xpb_out[41][793],u_xpb_out[42][793],u_xpb_out[43][793],u_xpb_out[44][793],u_xpb_out[45][793],u_xpb_out[46][793],u_xpb_out[47][793],u_xpb_out[48][793],u_xpb_out[49][793],u_xpb_out[50][793],u_xpb_out[51][793],u_xpb_out[52][793],u_xpb_out[53][793],u_xpb_out[54][793],u_xpb_out[55][793],u_xpb_out[56][793],u_xpb_out[57][793],u_xpb_out[58][793],u_xpb_out[59][793],u_xpb_out[60][793],u_xpb_out[61][793],u_xpb_out[62][793],u_xpb_out[63][793],u_xpb_out[64][793],u_xpb_out[65][793],u_xpb_out[66][793],u_xpb_out[67][793],u_xpb_out[68][793],u_xpb_out[69][793],u_xpb_out[70][793],u_xpb_out[71][793],u_xpb_out[72][793],u_xpb_out[73][793],u_xpb_out[74][793],u_xpb_out[75][793],u_xpb_out[76][793],u_xpb_out[77][793],u_xpb_out[78][793],u_xpb_out[79][793],u_xpb_out[80][793],u_xpb_out[81][793],u_xpb_out[82][793],u_xpb_out[83][793],u_xpb_out[84][793],u_xpb_out[85][793],u_xpb_out[86][793],u_xpb_out[87][793],u_xpb_out[88][793],u_xpb_out[89][793],u_xpb_out[90][793],u_xpb_out[91][793],u_xpb_out[92][793],u_xpb_out[93][793],u_xpb_out[94][793],u_xpb_out[95][793],u_xpb_out[96][793],u_xpb_out[97][793],u_xpb_out[98][793],u_xpb_out[99][793],u_xpb_out[100][793],u_xpb_out[101][793],u_xpb_out[102][793],u_xpb_out[103][793],u_xpb_out[104][793],u_xpb_out[105][793]};

assign col_out_794 = {u_xpb_out[0][794],u_xpb_out[1][794],u_xpb_out[2][794],u_xpb_out[3][794],u_xpb_out[4][794],u_xpb_out[5][794],u_xpb_out[6][794],u_xpb_out[7][794],u_xpb_out[8][794],u_xpb_out[9][794],u_xpb_out[10][794],u_xpb_out[11][794],u_xpb_out[12][794],u_xpb_out[13][794],u_xpb_out[14][794],u_xpb_out[15][794],u_xpb_out[16][794],u_xpb_out[17][794],u_xpb_out[18][794],u_xpb_out[19][794],u_xpb_out[20][794],u_xpb_out[21][794],u_xpb_out[22][794],u_xpb_out[23][794],u_xpb_out[24][794],u_xpb_out[25][794],u_xpb_out[26][794],u_xpb_out[27][794],u_xpb_out[28][794],u_xpb_out[29][794],u_xpb_out[30][794],u_xpb_out[31][794],u_xpb_out[32][794],u_xpb_out[33][794],u_xpb_out[34][794],u_xpb_out[35][794],u_xpb_out[36][794],u_xpb_out[37][794],u_xpb_out[38][794],u_xpb_out[39][794],u_xpb_out[40][794],u_xpb_out[41][794],u_xpb_out[42][794],u_xpb_out[43][794],u_xpb_out[44][794],u_xpb_out[45][794],u_xpb_out[46][794],u_xpb_out[47][794],u_xpb_out[48][794],u_xpb_out[49][794],u_xpb_out[50][794],u_xpb_out[51][794],u_xpb_out[52][794],u_xpb_out[53][794],u_xpb_out[54][794],u_xpb_out[55][794],u_xpb_out[56][794],u_xpb_out[57][794],u_xpb_out[58][794],u_xpb_out[59][794],u_xpb_out[60][794],u_xpb_out[61][794],u_xpb_out[62][794],u_xpb_out[63][794],u_xpb_out[64][794],u_xpb_out[65][794],u_xpb_out[66][794],u_xpb_out[67][794],u_xpb_out[68][794],u_xpb_out[69][794],u_xpb_out[70][794],u_xpb_out[71][794],u_xpb_out[72][794],u_xpb_out[73][794],u_xpb_out[74][794],u_xpb_out[75][794],u_xpb_out[76][794],u_xpb_out[77][794],u_xpb_out[78][794],u_xpb_out[79][794],u_xpb_out[80][794],u_xpb_out[81][794],u_xpb_out[82][794],u_xpb_out[83][794],u_xpb_out[84][794],u_xpb_out[85][794],u_xpb_out[86][794],u_xpb_out[87][794],u_xpb_out[88][794],u_xpb_out[89][794],u_xpb_out[90][794],u_xpb_out[91][794],u_xpb_out[92][794],u_xpb_out[93][794],u_xpb_out[94][794],u_xpb_out[95][794],u_xpb_out[96][794],u_xpb_out[97][794],u_xpb_out[98][794],u_xpb_out[99][794],u_xpb_out[100][794],u_xpb_out[101][794],u_xpb_out[102][794],u_xpb_out[103][794],u_xpb_out[104][794],u_xpb_out[105][794]};

assign col_out_795 = {u_xpb_out[0][795],u_xpb_out[1][795],u_xpb_out[2][795],u_xpb_out[3][795],u_xpb_out[4][795],u_xpb_out[5][795],u_xpb_out[6][795],u_xpb_out[7][795],u_xpb_out[8][795],u_xpb_out[9][795],u_xpb_out[10][795],u_xpb_out[11][795],u_xpb_out[12][795],u_xpb_out[13][795],u_xpb_out[14][795],u_xpb_out[15][795],u_xpb_out[16][795],u_xpb_out[17][795],u_xpb_out[18][795],u_xpb_out[19][795],u_xpb_out[20][795],u_xpb_out[21][795],u_xpb_out[22][795],u_xpb_out[23][795],u_xpb_out[24][795],u_xpb_out[25][795],u_xpb_out[26][795],u_xpb_out[27][795],u_xpb_out[28][795],u_xpb_out[29][795],u_xpb_out[30][795],u_xpb_out[31][795],u_xpb_out[32][795],u_xpb_out[33][795],u_xpb_out[34][795],u_xpb_out[35][795],u_xpb_out[36][795],u_xpb_out[37][795],u_xpb_out[38][795],u_xpb_out[39][795],u_xpb_out[40][795],u_xpb_out[41][795],u_xpb_out[42][795],u_xpb_out[43][795],u_xpb_out[44][795],u_xpb_out[45][795],u_xpb_out[46][795],u_xpb_out[47][795],u_xpb_out[48][795],u_xpb_out[49][795],u_xpb_out[50][795],u_xpb_out[51][795],u_xpb_out[52][795],u_xpb_out[53][795],u_xpb_out[54][795],u_xpb_out[55][795],u_xpb_out[56][795],u_xpb_out[57][795],u_xpb_out[58][795],u_xpb_out[59][795],u_xpb_out[60][795],u_xpb_out[61][795],u_xpb_out[62][795],u_xpb_out[63][795],u_xpb_out[64][795],u_xpb_out[65][795],u_xpb_out[66][795],u_xpb_out[67][795],u_xpb_out[68][795],u_xpb_out[69][795],u_xpb_out[70][795],u_xpb_out[71][795],u_xpb_out[72][795],u_xpb_out[73][795],u_xpb_out[74][795],u_xpb_out[75][795],u_xpb_out[76][795],u_xpb_out[77][795],u_xpb_out[78][795],u_xpb_out[79][795],u_xpb_out[80][795],u_xpb_out[81][795],u_xpb_out[82][795],u_xpb_out[83][795],u_xpb_out[84][795],u_xpb_out[85][795],u_xpb_out[86][795],u_xpb_out[87][795],u_xpb_out[88][795],u_xpb_out[89][795],u_xpb_out[90][795],u_xpb_out[91][795],u_xpb_out[92][795],u_xpb_out[93][795],u_xpb_out[94][795],u_xpb_out[95][795],u_xpb_out[96][795],u_xpb_out[97][795],u_xpb_out[98][795],u_xpb_out[99][795],u_xpb_out[100][795],u_xpb_out[101][795],u_xpb_out[102][795],u_xpb_out[103][795],u_xpb_out[104][795],u_xpb_out[105][795]};

assign col_out_796 = {u_xpb_out[0][796],u_xpb_out[1][796],u_xpb_out[2][796],u_xpb_out[3][796],u_xpb_out[4][796],u_xpb_out[5][796],u_xpb_out[6][796],u_xpb_out[7][796],u_xpb_out[8][796],u_xpb_out[9][796],u_xpb_out[10][796],u_xpb_out[11][796],u_xpb_out[12][796],u_xpb_out[13][796],u_xpb_out[14][796],u_xpb_out[15][796],u_xpb_out[16][796],u_xpb_out[17][796],u_xpb_out[18][796],u_xpb_out[19][796],u_xpb_out[20][796],u_xpb_out[21][796],u_xpb_out[22][796],u_xpb_out[23][796],u_xpb_out[24][796],u_xpb_out[25][796],u_xpb_out[26][796],u_xpb_out[27][796],u_xpb_out[28][796],u_xpb_out[29][796],u_xpb_out[30][796],u_xpb_out[31][796],u_xpb_out[32][796],u_xpb_out[33][796],u_xpb_out[34][796],u_xpb_out[35][796],u_xpb_out[36][796],u_xpb_out[37][796],u_xpb_out[38][796],u_xpb_out[39][796],u_xpb_out[40][796],u_xpb_out[41][796],u_xpb_out[42][796],u_xpb_out[43][796],u_xpb_out[44][796],u_xpb_out[45][796],u_xpb_out[46][796],u_xpb_out[47][796],u_xpb_out[48][796],u_xpb_out[49][796],u_xpb_out[50][796],u_xpb_out[51][796],u_xpb_out[52][796],u_xpb_out[53][796],u_xpb_out[54][796],u_xpb_out[55][796],u_xpb_out[56][796],u_xpb_out[57][796],u_xpb_out[58][796],u_xpb_out[59][796],u_xpb_out[60][796],u_xpb_out[61][796],u_xpb_out[62][796],u_xpb_out[63][796],u_xpb_out[64][796],u_xpb_out[65][796],u_xpb_out[66][796],u_xpb_out[67][796],u_xpb_out[68][796],u_xpb_out[69][796],u_xpb_out[70][796],u_xpb_out[71][796],u_xpb_out[72][796],u_xpb_out[73][796],u_xpb_out[74][796],u_xpb_out[75][796],u_xpb_out[76][796],u_xpb_out[77][796],u_xpb_out[78][796],u_xpb_out[79][796],u_xpb_out[80][796],u_xpb_out[81][796],u_xpb_out[82][796],u_xpb_out[83][796],u_xpb_out[84][796],u_xpb_out[85][796],u_xpb_out[86][796],u_xpb_out[87][796],u_xpb_out[88][796],u_xpb_out[89][796],u_xpb_out[90][796],u_xpb_out[91][796],u_xpb_out[92][796],u_xpb_out[93][796],u_xpb_out[94][796],u_xpb_out[95][796],u_xpb_out[96][796],u_xpb_out[97][796],u_xpb_out[98][796],u_xpb_out[99][796],u_xpb_out[100][796],u_xpb_out[101][796],u_xpb_out[102][796],u_xpb_out[103][796],u_xpb_out[104][796],u_xpb_out[105][796]};

assign col_out_797 = {u_xpb_out[0][797],u_xpb_out[1][797],u_xpb_out[2][797],u_xpb_out[3][797],u_xpb_out[4][797],u_xpb_out[5][797],u_xpb_out[6][797],u_xpb_out[7][797],u_xpb_out[8][797],u_xpb_out[9][797],u_xpb_out[10][797],u_xpb_out[11][797],u_xpb_out[12][797],u_xpb_out[13][797],u_xpb_out[14][797],u_xpb_out[15][797],u_xpb_out[16][797],u_xpb_out[17][797],u_xpb_out[18][797],u_xpb_out[19][797],u_xpb_out[20][797],u_xpb_out[21][797],u_xpb_out[22][797],u_xpb_out[23][797],u_xpb_out[24][797],u_xpb_out[25][797],u_xpb_out[26][797],u_xpb_out[27][797],u_xpb_out[28][797],u_xpb_out[29][797],u_xpb_out[30][797],u_xpb_out[31][797],u_xpb_out[32][797],u_xpb_out[33][797],u_xpb_out[34][797],u_xpb_out[35][797],u_xpb_out[36][797],u_xpb_out[37][797],u_xpb_out[38][797],u_xpb_out[39][797],u_xpb_out[40][797],u_xpb_out[41][797],u_xpb_out[42][797],u_xpb_out[43][797],u_xpb_out[44][797],u_xpb_out[45][797],u_xpb_out[46][797],u_xpb_out[47][797],u_xpb_out[48][797],u_xpb_out[49][797],u_xpb_out[50][797],u_xpb_out[51][797],u_xpb_out[52][797],u_xpb_out[53][797],u_xpb_out[54][797],u_xpb_out[55][797],u_xpb_out[56][797],u_xpb_out[57][797],u_xpb_out[58][797],u_xpb_out[59][797],u_xpb_out[60][797],u_xpb_out[61][797],u_xpb_out[62][797],u_xpb_out[63][797],u_xpb_out[64][797],u_xpb_out[65][797],u_xpb_out[66][797],u_xpb_out[67][797],u_xpb_out[68][797],u_xpb_out[69][797],u_xpb_out[70][797],u_xpb_out[71][797],u_xpb_out[72][797],u_xpb_out[73][797],u_xpb_out[74][797],u_xpb_out[75][797],u_xpb_out[76][797],u_xpb_out[77][797],u_xpb_out[78][797],u_xpb_out[79][797],u_xpb_out[80][797],u_xpb_out[81][797],u_xpb_out[82][797],u_xpb_out[83][797],u_xpb_out[84][797],u_xpb_out[85][797],u_xpb_out[86][797],u_xpb_out[87][797],u_xpb_out[88][797],u_xpb_out[89][797],u_xpb_out[90][797],u_xpb_out[91][797],u_xpb_out[92][797],u_xpb_out[93][797],u_xpb_out[94][797],u_xpb_out[95][797],u_xpb_out[96][797],u_xpb_out[97][797],u_xpb_out[98][797],u_xpb_out[99][797],u_xpb_out[100][797],u_xpb_out[101][797],u_xpb_out[102][797],u_xpb_out[103][797],u_xpb_out[104][797],u_xpb_out[105][797]};

assign col_out_798 = {u_xpb_out[0][798],u_xpb_out[1][798],u_xpb_out[2][798],u_xpb_out[3][798],u_xpb_out[4][798],u_xpb_out[5][798],u_xpb_out[6][798],u_xpb_out[7][798],u_xpb_out[8][798],u_xpb_out[9][798],u_xpb_out[10][798],u_xpb_out[11][798],u_xpb_out[12][798],u_xpb_out[13][798],u_xpb_out[14][798],u_xpb_out[15][798],u_xpb_out[16][798],u_xpb_out[17][798],u_xpb_out[18][798],u_xpb_out[19][798],u_xpb_out[20][798],u_xpb_out[21][798],u_xpb_out[22][798],u_xpb_out[23][798],u_xpb_out[24][798],u_xpb_out[25][798],u_xpb_out[26][798],u_xpb_out[27][798],u_xpb_out[28][798],u_xpb_out[29][798],u_xpb_out[30][798],u_xpb_out[31][798],u_xpb_out[32][798],u_xpb_out[33][798],u_xpb_out[34][798],u_xpb_out[35][798],u_xpb_out[36][798],u_xpb_out[37][798],u_xpb_out[38][798],u_xpb_out[39][798],u_xpb_out[40][798],u_xpb_out[41][798],u_xpb_out[42][798],u_xpb_out[43][798],u_xpb_out[44][798],u_xpb_out[45][798],u_xpb_out[46][798],u_xpb_out[47][798],u_xpb_out[48][798],u_xpb_out[49][798],u_xpb_out[50][798],u_xpb_out[51][798],u_xpb_out[52][798],u_xpb_out[53][798],u_xpb_out[54][798],u_xpb_out[55][798],u_xpb_out[56][798],u_xpb_out[57][798],u_xpb_out[58][798],u_xpb_out[59][798],u_xpb_out[60][798],u_xpb_out[61][798],u_xpb_out[62][798],u_xpb_out[63][798],u_xpb_out[64][798],u_xpb_out[65][798],u_xpb_out[66][798],u_xpb_out[67][798],u_xpb_out[68][798],u_xpb_out[69][798],u_xpb_out[70][798],u_xpb_out[71][798],u_xpb_out[72][798],u_xpb_out[73][798],u_xpb_out[74][798],u_xpb_out[75][798],u_xpb_out[76][798],u_xpb_out[77][798],u_xpb_out[78][798],u_xpb_out[79][798],u_xpb_out[80][798],u_xpb_out[81][798],u_xpb_out[82][798],u_xpb_out[83][798],u_xpb_out[84][798],u_xpb_out[85][798],u_xpb_out[86][798],u_xpb_out[87][798],u_xpb_out[88][798],u_xpb_out[89][798],u_xpb_out[90][798],u_xpb_out[91][798],u_xpb_out[92][798],u_xpb_out[93][798],u_xpb_out[94][798],u_xpb_out[95][798],u_xpb_out[96][798],u_xpb_out[97][798],u_xpb_out[98][798],u_xpb_out[99][798],u_xpb_out[100][798],u_xpb_out[101][798],u_xpb_out[102][798],u_xpb_out[103][798],u_xpb_out[104][798],u_xpb_out[105][798]};

assign col_out_799 = {u_xpb_out[0][799],u_xpb_out[1][799],u_xpb_out[2][799],u_xpb_out[3][799],u_xpb_out[4][799],u_xpb_out[5][799],u_xpb_out[6][799],u_xpb_out[7][799],u_xpb_out[8][799],u_xpb_out[9][799],u_xpb_out[10][799],u_xpb_out[11][799],u_xpb_out[12][799],u_xpb_out[13][799],u_xpb_out[14][799],u_xpb_out[15][799],u_xpb_out[16][799],u_xpb_out[17][799],u_xpb_out[18][799],u_xpb_out[19][799],u_xpb_out[20][799],u_xpb_out[21][799],u_xpb_out[22][799],u_xpb_out[23][799],u_xpb_out[24][799],u_xpb_out[25][799],u_xpb_out[26][799],u_xpb_out[27][799],u_xpb_out[28][799],u_xpb_out[29][799],u_xpb_out[30][799],u_xpb_out[31][799],u_xpb_out[32][799],u_xpb_out[33][799],u_xpb_out[34][799],u_xpb_out[35][799],u_xpb_out[36][799],u_xpb_out[37][799],u_xpb_out[38][799],u_xpb_out[39][799],u_xpb_out[40][799],u_xpb_out[41][799],u_xpb_out[42][799],u_xpb_out[43][799],u_xpb_out[44][799],u_xpb_out[45][799],u_xpb_out[46][799],u_xpb_out[47][799],u_xpb_out[48][799],u_xpb_out[49][799],u_xpb_out[50][799],u_xpb_out[51][799],u_xpb_out[52][799],u_xpb_out[53][799],u_xpb_out[54][799],u_xpb_out[55][799],u_xpb_out[56][799],u_xpb_out[57][799],u_xpb_out[58][799],u_xpb_out[59][799],u_xpb_out[60][799],u_xpb_out[61][799],u_xpb_out[62][799],u_xpb_out[63][799],u_xpb_out[64][799],u_xpb_out[65][799],u_xpb_out[66][799],u_xpb_out[67][799],u_xpb_out[68][799],u_xpb_out[69][799],u_xpb_out[70][799],u_xpb_out[71][799],u_xpb_out[72][799],u_xpb_out[73][799],u_xpb_out[74][799],u_xpb_out[75][799],u_xpb_out[76][799],u_xpb_out[77][799],u_xpb_out[78][799],u_xpb_out[79][799],u_xpb_out[80][799],u_xpb_out[81][799],u_xpb_out[82][799],u_xpb_out[83][799],u_xpb_out[84][799],u_xpb_out[85][799],u_xpb_out[86][799],u_xpb_out[87][799],u_xpb_out[88][799],u_xpb_out[89][799],u_xpb_out[90][799],u_xpb_out[91][799],u_xpb_out[92][799],u_xpb_out[93][799],u_xpb_out[94][799],u_xpb_out[95][799],u_xpb_out[96][799],u_xpb_out[97][799],u_xpb_out[98][799],u_xpb_out[99][799],u_xpb_out[100][799],u_xpb_out[101][799],u_xpb_out[102][799],u_xpb_out[103][799],u_xpb_out[104][799],u_xpb_out[105][799]};

assign col_out_800 = {u_xpb_out[0][800],u_xpb_out[1][800],u_xpb_out[2][800],u_xpb_out[3][800],u_xpb_out[4][800],u_xpb_out[5][800],u_xpb_out[6][800],u_xpb_out[7][800],u_xpb_out[8][800],u_xpb_out[9][800],u_xpb_out[10][800],u_xpb_out[11][800],u_xpb_out[12][800],u_xpb_out[13][800],u_xpb_out[14][800],u_xpb_out[15][800],u_xpb_out[16][800],u_xpb_out[17][800],u_xpb_out[18][800],u_xpb_out[19][800],u_xpb_out[20][800],u_xpb_out[21][800],u_xpb_out[22][800],u_xpb_out[23][800],u_xpb_out[24][800],u_xpb_out[25][800],u_xpb_out[26][800],u_xpb_out[27][800],u_xpb_out[28][800],u_xpb_out[29][800],u_xpb_out[30][800],u_xpb_out[31][800],u_xpb_out[32][800],u_xpb_out[33][800],u_xpb_out[34][800],u_xpb_out[35][800],u_xpb_out[36][800],u_xpb_out[37][800],u_xpb_out[38][800],u_xpb_out[39][800],u_xpb_out[40][800],u_xpb_out[41][800],u_xpb_out[42][800],u_xpb_out[43][800],u_xpb_out[44][800],u_xpb_out[45][800],u_xpb_out[46][800],u_xpb_out[47][800],u_xpb_out[48][800],u_xpb_out[49][800],u_xpb_out[50][800],u_xpb_out[51][800],u_xpb_out[52][800],u_xpb_out[53][800],u_xpb_out[54][800],u_xpb_out[55][800],u_xpb_out[56][800],u_xpb_out[57][800],u_xpb_out[58][800],u_xpb_out[59][800],u_xpb_out[60][800],u_xpb_out[61][800],u_xpb_out[62][800],u_xpb_out[63][800],u_xpb_out[64][800],u_xpb_out[65][800],u_xpb_out[66][800],u_xpb_out[67][800],u_xpb_out[68][800],u_xpb_out[69][800],u_xpb_out[70][800],u_xpb_out[71][800],u_xpb_out[72][800],u_xpb_out[73][800],u_xpb_out[74][800],u_xpb_out[75][800],u_xpb_out[76][800],u_xpb_out[77][800],u_xpb_out[78][800],u_xpb_out[79][800],u_xpb_out[80][800],u_xpb_out[81][800],u_xpb_out[82][800],u_xpb_out[83][800],u_xpb_out[84][800],u_xpb_out[85][800],u_xpb_out[86][800],u_xpb_out[87][800],u_xpb_out[88][800],u_xpb_out[89][800],u_xpb_out[90][800],u_xpb_out[91][800],u_xpb_out[92][800],u_xpb_out[93][800],u_xpb_out[94][800],u_xpb_out[95][800],u_xpb_out[96][800],u_xpb_out[97][800],u_xpb_out[98][800],u_xpb_out[99][800],u_xpb_out[100][800],u_xpb_out[101][800],u_xpb_out[102][800],u_xpb_out[103][800],u_xpb_out[104][800],u_xpb_out[105][800]};

assign col_out_801 = {u_xpb_out[0][801],u_xpb_out[1][801],u_xpb_out[2][801],u_xpb_out[3][801],u_xpb_out[4][801],u_xpb_out[5][801],u_xpb_out[6][801],u_xpb_out[7][801],u_xpb_out[8][801],u_xpb_out[9][801],u_xpb_out[10][801],u_xpb_out[11][801],u_xpb_out[12][801],u_xpb_out[13][801],u_xpb_out[14][801],u_xpb_out[15][801],u_xpb_out[16][801],u_xpb_out[17][801],u_xpb_out[18][801],u_xpb_out[19][801],u_xpb_out[20][801],u_xpb_out[21][801],u_xpb_out[22][801],u_xpb_out[23][801],u_xpb_out[24][801],u_xpb_out[25][801],u_xpb_out[26][801],u_xpb_out[27][801],u_xpb_out[28][801],u_xpb_out[29][801],u_xpb_out[30][801],u_xpb_out[31][801],u_xpb_out[32][801],u_xpb_out[33][801],u_xpb_out[34][801],u_xpb_out[35][801],u_xpb_out[36][801],u_xpb_out[37][801],u_xpb_out[38][801],u_xpb_out[39][801],u_xpb_out[40][801],u_xpb_out[41][801],u_xpb_out[42][801],u_xpb_out[43][801],u_xpb_out[44][801],u_xpb_out[45][801],u_xpb_out[46][801],u_xpb_out[47][801],u_xpb_out[48][801],u_xpb_out[49][801],u_xpb_out[50][801],u_xpb_out[51][801],u_xpb_out[52][801],u_xpb_out[53][801],u_xpb_out[54][801],u_xpb_out[55][801],u_xpb_out[56][801],u_xpb_out[57][801],u_xpb_out[58][801],u_xpb_out[59][801],u_xpb_out[60][801],u_xpb_out[61][801],u_xpb_out[62][801],u_xpb_out[63][801],u_xpb_out[64][801],u_xpb_out[65][801],u_xpb_out[66][801],u_xpb_out[67][801],u_xpb_out[68][801],u_xpb_out[69][801],u_xpb_out[70][801],u_xpb_out[71][801],u_xpb_out[72][801],u_xpb_out[73][801],u_xpb_out[74][801],u_xpb_out[75][801],u_xpb_out[76][801],u_xpb_out[77][801],u_xpb_out[78][801],u_xpb_out[79][801],u_xpb_out[80][801],u_xpb_out[81][801],u_xpb_out[82][801],u_xpb_out[83][801],u_xpb_out[84][801],u_xpb_out[85][801],u_xpb_out[86][801],u_xpb_out[87][801],u_xpb_out[88][801],u_xpb_out[89][801],u_xpb_out[90][801],u_xpb_out[91][801],u_xpb_out[92][801],u_xpb_out[93][801],u_xpb_out[94][801],u_xpb_out[95][801],u_xpb_out[96][801],u_xpb_out[97][801],u_xpb_out[98][801],u_xpb_out[99][801],u_xpb_out[100][801],u_xpb_out[101][801],u_xpb_out[102][801],u_xpb_out[103][801],u_xpb_out[104][801],u_xpb_out[105][801]};

assign col_out_802 = {u_xpb_out[0][802],u_xpb_out[1][802],u_xpb_out[2][802],u_xpb_out[3][802],u_xpb_out[4][802],u_xpb_out[5][802],u_xpb_out[6][802],u_xpb_out[7][802],u_xpb_out[8][802],u_xpb_out[9][802],u_xpb_out[10][802],u_xpb_out[11][802],u_xpb_out[12][802],u_xpb_out[13][802],u_xpb_out[14][802],u_xpb_out[15][802],u_xpb_out[16][802],u_xpb_out[17][802],u_xpb_out[18][802],u_xpb_out[19][802],u_xpb_out[20][802],u_xpb_out[21][802],u_xpb_out[22][802],u_xpb_out[23][802],u_xpb_out[24][802],u_xpb_out[25][802],u_xpb_out[26][802],u_xpb_out[27][802],u_xpb_out[28][802],u_xpb_out[29][802],u_xpb_out[30][802],u_xpb_out[31][802],u_xpb_out[32][802],u_xpb_out[33][802],u_xpb_out[34][802],u_xpb_out[35][802],u_xpb_out[36][802],u_xpb_out[37][802],u_xpb_out[38][802],u_xpb_out[39][802],u_xpb_out[40][802],u_xpb_out[41][802],u_xpb_out[42][802],u_xpb_out[43][802],u_xpb_out[44][802],u_xpb_out[45][802],u_xpb_out[46][802],u_xpb_out[47][802],u_xpb_out[48][802],u_xpb_out[49][802],u_xpb_out[50][802],u_xpb_out[51][802],u_xpb_out[52][802],u_xpb_out[53][802],u_xpb_out[54][802],u_xpb_out[55][802],u_xpb_out[56][802],u_xpb_out[57][802],u_xpb_out[58][802],u_xpb_out[59][802],u_xpb_out[60][802],u_xpb_out[61][802],u_xpb_out[62][802],u_xpb_out[63][802],u_xpb_out[64][802],u_xpb_out[65][802],u_xpb_out[66][802],u_xpb_out[67][802],u_xpb_out[68][802],u_xpb_out[69][802],u_xpb_out[70][802],u_xpb_out[71][802],u_xpb_out[72][802],u_xpb_out[73][802],u_xpb_out[74][802],u_xpb_out[75][802],u_xpb_out[76][802],u_xpb_out[77][802],u_xpb_out[78][802],u_xpb_out[79][802],u_xpb_out[80][802],u_xpb_out[81][802],u_xpb_out[82][802],u_xpb_out[83][802],u_xpb_out[84][802],u_xpb_out[85][802],u_xpb_out[86][802],u_xpb_out[87][802],u_xpb_out[88][802],u_xpb_out[89][802],u_xpb_out[90][802],u_xpb_out[91][802],u_xpb_out[92][802],u_xpb_out[93][802],u_xpb_out[94][802],u_xpb_out[95][802],u_xpb_out[96][802],u_xpb_out[97][802],u_xpb_out[98][802],u_xpb_out[99][802],u_xpb_out[100][802],u_xpb_out[101][802],u_xpb_out[102][802],u_xpb_out[103][802],u_xpb_out[104][802],u_xpb_out[105][802]};

assign col_out_803 = {u_xpb_out[0][803],u_xpb_out[1][803],u_xpb_out[2][803],u_xpb_out[3][803],u_xpb_out[4][803],u_xpb_out[5][803],u_xpb_out[6][803],u_xpb_out[7][803],u_xpb_out[8][803],u_xpb_out[9][803],u_xpb_out[10][803],u_xpb_out[11][803],u_xpb_out[12][803],u_xpb_out[13][803],u_xpb_out[14][803],u_xpb_out[15][803],u_xpb_out[16][803],u_xpb_out[17][803],u_xpb_out[18][803],u_xpb_out[19][803],u_xpb_out[20][803],u_xpb_out[21][803],u_xpb_out[22][803],u_xpb_out[23][803],u_xpb_out[24][803],u_xpb_out[25][803],u_xpb_out[26][803],u_xpb_out[27][803],u_xpb_out[28][803],u_xpb_out[29][803],u_xpb_out[30][803],u_xpb_out[31][803],u_xpb_out[32][803],u_xpb_out[33][803],u_xpb_out[34][803],u_xpb_out[35][803],u_xpb_out[36][803],u_xpb_out[37][803],u_xpb_out[38][803],u_xpb_out[39][803],u_xpb_out[40][803],u_xpb_out[41][803],u_xpb_out[42][803],u_xpb_out[43][803],u_xpb_out[44][803],u_xpb_out[45][803],u_xpb_out[46][803],u_xpb_out[47][803],u_xpb_out[48][803],u_xpb_out[49][803],u_xpb_out[50][803],u_xpb_out[51][803],u_xpb_out[52][803],u_xpb_out[53][803],u_xpb_out[54][803],u_xpb_out[55][803],u_xpb_out[56][803],u_xpb_out[57][803],u_xpb_out[58][803],u_xpb_out[59][803],u_xpb_out[60][803],u_xpb_out[61][803],u_xpb_out[62][803],u_xpb_out[63][803],u_xpb_out[64][803],u_xpb_out[65][803],u_xpb_out[66][803],u_xpb_out[67][803],u_xpb_out[68][803],u_xpb_out[69][803],u_xpb_out[70][803],u_xpb_out[71][803],u_xpb_out[72][803],u_xpb_out[73][803],u_xpb_out[74][803],u_xpb_out[75][803],u_xpb_out[76][803],u_xpb_out[77][803],u_xpb_out[78][803],u_xpb_out[79][803],u_xpb_out[80][803],u_xpb_out[81][803],u_xpb_out[82][803],u_xpb_out[83][803],u_xpb_out[84][803],u_xpb_out[85][803],u_xpb_out[86][803],u_xpb_out[87][803],u_xpb_out[88][803],u_xpb_out[89][803],u_xpb_out[90][803],u_xpb_out[91][803],u_xpb_out[92][803],u_xpb_out[93][803],u_xpb_out[94][803],u_xpb_out[95][803],u_xpb_out[96][803],u_xpb_out[97][803],u_xpb_out[98][803],u_xpb_out[99][803],u_xpb_out[100][803],u_xpb_out[101][803],u_xpb_out[102][803],u_xpb_out[103][803],u_xpb_out[104][803],u_xpb_out[105][803]};

assign col_out_804 = {u_xpb_out[0][804],u_xpb_out[1][804],u_xpb_out[2][804],u_xpb_out[3][804],u_xpb_out[4][804],u_xpb_out[5][804],u_xpb_out[6][804],u_xpb_out[7][804],u_xpb_out[8][804],u_xpb_out[9][804],u_xpb_out[10][804],u_xpb_out[11][804],u_xpb_out[12][804],u_xpb_out[13][804],u_xpb_out[14][804],u_xpb_out[15][804],u_xpb_out[16][804],u_xpb_out[17][804],u_xpb_out[18][804],u_xpb_out[19][804],u_xpb_out[20][804],u_xpb_out[21][804],u_xpb_out[22][804],u_xpb_out[23][804],u_xpb_out[24][804],u_xpb_out[25][804],u_xpb_out[26][804],u_xpb_out[27][804],u_xpb_out[28][804],u_xpb_out[29][804],u_xpb_out[30][804],u_xpb_out[31][804],u_xpb_out[32][804],u_xpb_out[33][804],u_xpb_out[34][804],u_xpb_out[35][804],u_xpb_out[36][804],u_xpb_out[37][804],u_xpb_out[38][804],u_xpb_out[39][804],u_xpb_out[40][804],u_xpb_out[41][804],u_xpb_out[42][804],u_xpb_out[43][804],u_xpb_out[44][804],u_xpb_out[45][804],u_xpb_out[46][804],u_xpb_out[47][804],u_xpb_out[48][804],u_xpb_out[49][804],u_xpb_out[50][804],u_xpb_out[51][804],u_xpb_out[52][804],u_xpb_out[53][804],u_xpb_out[54][804],u_xpb_out[55][804],u_xpb_out[56][804],u_xpb_out[57][804],u_xpb_out[58][804],u_xpb_out[59][804],u_xpb_out[60][804],u_xpb_out[61][804],u_xpb_out[62][804],u_xpb_out[63][804],u_xpb_out[64][804],u_xpb_out[65][804],u_xpb_out[66][804],u_xpb_out[67][804],u_xpb_out[68][804],u_xpb_out[69][804],u_xpb_out[70][804],u_xpb_out[71][804],u_xpb_out[72][804],u_xpb_out[73][804],u_xpb_out[74][804],u_xpb_out[75][804],u_xpb_out[76][804],u_xpb_out[77][804],u_xpb_out[78][804],u_xpb_out[79][804],u_xpb_out[80][804],u_xpb_out[81][804],u_xpb_out[82][804],u_xpb_out[83][804],u_xpb_out[84][804],u_xpb_out[85][804],u_xpb_out[86][804],u_xpb_out[87][804],u_xpb_out[88][804],u_xpb_out[89][804],u_xpb_out[90][804],u_xpb_out[91][804],u_xpb_out[92][804],u_xpb_out[93][804],u_xpb_out[94][804],u_xpb_out[95][804],u_xpb_out[96][804],u_xpb_out[97][804],u_xpb_out[98][804],u_xpb_out[99][804],u_xpb_out[100][804],u_xpb_out[101][804],u_xpb_out[102][804],u_xpb_out[103][804],u_xpb_out[104][804],u_xpb_out[105][804]};

assign col_out_805 = {u_xpb_out[0][805],u_xpb_out[1][805],u_xpb_out[2][805],u_xpb_out[3][805],u_xpb_out[4][805],u_xpb_out[5][805],u_xpb_out[6][805],u_xpb_out[7][805],u_xpb_out[8][805],u_xpb_out[9][805],u_xpb_out[10][805],u_xpb_out[11][805],u_xpb_out[12][805],u_xpb_out[13][805],u_xpb_out[14][805],u_xpb_out[15][805],u_xpb_out[16][805],u_xpb_out[17][805],u_xpb_out[18][805],u_xpb_out[19][805],u_xpb_out[20][805],u_xpb_out[21][805],u_xpb_out[22][805],u_xpb_out[23][805],u_xpb_out[24][805],u_xpb_out[25][805],u_xpb_out[26][805],u_xpb_out[27][805],u_xpb_out[28][805],u_xpb_out[29][805],u_xpb_out[30][805],u_xpb_out[31][805],u_xpb_out[32][805],u_xpb_out[33][805],u_xpb_out[34][805],u_xpb_out[35][805],u_xpb_out[36][805],u_xpb_out[37][805],u_xpb_out[38][805],u_xpb_out[39][805],u_xpb_out[40][805],u_xpb_out[41][805],u_xpb_out[42][805],u_xpb_out[43][805],u_xpb_out[44][805],u_xpb_out[45][805],u_xpb_out[46][805],u_xpb_out[47][805],u_xpb_out[48][805],u_xpb_out[49][805],u_xpb_out[50][805],u_xpb_out[51][805],u_xpb_out[52][805],u_xpb_out[53][805],u_xpb_out[54][805],u_xpb_out[55][805],u_xpb_out[56][805],u_xpb_out[57][805],u_xpb_out[58][805],u_xpb_out[59][805],u_xpb_out[60][805],u_xpb_out[61][805],u_xpb_out[62][805],u_xpb_out[63][805],u_xpb_out[64][805],u_xpb_out[65][805],u_xpb_out[66][805],u_xpb_out[67][805],u_xpb_out[68][805],u_xpb_out[69][805],u_xpb_out[70][805],u_xpb_out[71][805],u_xpb_out[72][805],u_xpb_out[73][805],u_xpb_out[74][805],u_xpb_out[75][805],u_xpb_out[76][805],u_xpb_out[77][805],u_xpb_out[78][805],u_xpb_out[79][805],u_xpb_out[80][805],u_xpb_out[81][805],u_xpb_out[82][805],u_xpb_out[83][805],u_xpb_out[84][805],u_xpb_out[85][805],u_xpb_out[86][805],u_xpb_out[87][805],u_xpb_out[88][805],u_xpb_out[89][805],u_xpb_out[90][805],u_xpb_out[91][805],u_xpb_out[92][805],u_xpb_out[93][805],u_xpb_out[94][805],u_xpb_out[95][805],u_xpb_out[96][805],u_xpb_out[97][805],u_xpb_out[98][805],u_xpb_out[99][805],u_xpb_out[100][805],u_xpb_out[101][805],u_xpb_out[102][805],u_xpb_out[103][805],u_xpb_out[104][805],u_xpb_out[105][805]};

assign col_out_806 = {u_xpb_out[0][806],u_xpb_out[1][806],u_xpb_out[2][806],u_xpb_out[3][806],u_xpb_out[4][806],u_xpb_out[5][806],u_xpb_out[6][806],u_xpb_out[7][806],u_xpb_out[8][806],u_xpb_out[9][806],u_xpb_out[10][806],u_xpb_out[11][806],u_xpb_out[12][806],u_xpb_out[13][806],u_xpb_out[14][806],u_xpb_out[15][806],u_xpb_out[16][806],u_xpb_out[17][806],u_xpb_out[18][806],u_xpb_out[19][806],u_xpb_out[20][806],u_xpb_out[21][806],u_xpb_out[22][806],u_xpb_out[23][806],u_xpb_out[24][806],u_xpb_out[25][806],u_xpb_out[26][806],u_xpb_out[27][806],u_xpb_out[28][806],u_xpb_out[29][806],u_xpb_out[30][806],u_xpb_out[31][806],u_xpb_out[32][806],u_xpb_out[33][806],u_xpb_out[34][806],u_xpb_out[35][806],u_xpb_out[36][806],u_xpb_out[37][806],u_xpb_out[38][806],u_xpb_out[39][806],u_xpb_out[40][806],u_xpb_out[41][806],u_xpb_out[42][806],u_xpb_out[43][806],u_xpb_out[44][806],u_xpb_out[45][806],u_xpb_out[46][806],u_xpb_out[47][806],u_xpb_out[48][806],u_xpb_out[49][806],u_xpb_out[50][806],u_xpb_out[51][806],u_xpb_out[52][806],u_xpb_out[53][806],u_xpb_out[54][806],u_xpb_out[55][806],u_xpb_out[56][806],u_xpb_out[57][806],u_xpb_out[58][806],u_xpb_out[59][806],u_xpb_out[60][806],u_xpb_out[61][806],u_xpb_out[62][806],u_xpb_out[63][806],u_xpb_out[64][806],u_xpb_out[65][806],u_xpb_out[66][806],u_xpb_out[67][806],u_xpb_out[68][806],u_xpb_out[69][806],u_xpb_out[70][806],u_xpb_out[71][806],u_xpb_out[72][806],u_xpb_out[73][806],u_xpb_out[74][806],u_xpb_out[75][806],u_xpb_out[76][806],u_xpb_out[77][806],u_xpb_out[78][806],u_xpb_out[79][806],u_xpb_out[80][806],u_xpb_out[81][806],u_xpb_out[82][806],u_xpb_out[83][806],u_xpb_out[84][806],u_xpb_out[85][806],u_xpb_out[86][806],u_xpb_out[87][806],u_xpb_out[88][806],u_xpb_out[89][806],u_xpb_out[90][806],u_xpb_out[91][806],u_xpb_out[92][806],u_xpb_out[93][806],u_xpb_out[94][806],u_xpb_out[95][806],u_xpb_out[96][806],u_xpb_out[97][806],u_xpb_out[98][806],u_xpb_out[99][806],u_xpb_out[100][806],u_xpb_out[101][806],u_xpb_out[102][806],u_xpb_out[103][806],u_xpb_out[104][806],u_xpb_out[105][806]};

assign col_out_807 = {u_xpb_out[0][807],u_xpb_out[1][807],u_xpb_out[2][807],u_xpb_out[3][807],u_xpb_out[4][807],u_xpb_out[5][807],u_xpb_out[6][807],u_xpb_out[7][807],u_xpb_out[8][807],u_xpb_out[9][807],u_xpb_out[10][807],u_xpb_out[11][807],u_xpb_out[12][807],u_xpb_out[13][807],u_xpb_out[14][807],u_xpb_out[15][807],u_xpb_out[16][807],u_xpb_out[17][807],u_xpb_out[18][807],u_xpb_out[19][807],u_xpb_out[20][807],u_xpb_out[21][807],u_xpb_out[22][807],u_xpb_out[23][807],u_xpb_out[24][807],u_xpb_out[25][807],u_xpb_out[26][807],u_xpb_out[27][807],u_xpb_out[28][807],u_xpb_out[29][807],u_xpb_out[30][807],u_xpb_out[31][807],u_xpb_out[32][807],u_xpb_out[33][807],u_xpb_out[34][807],u_xpb_out[35][807],u_xpb_out[36][807],u_xpb_out[37][807],u_xpb_out[38][807],u_xpb_out[39][807],u_xpb_out[40][807],u_xpb_out[41][807],u_xpb_out[42][807],u_xpb_out[43][807],u_xpb_out[44][807],u_xpb_out[45][807],u_xpb_out[46][807],u_xpb_out[47][807],u_xpb_out[48][807],u_xpb_out[49][807],u_xpb_out[50][807],u_xpb_out[51][807],u_xpb_out[52][807],u_xpb_out[53][807],u_xpb_out[54][807],u_xpb_out[55][807],u_xpb_out[56][807],u_xpb_out[57][807],u_xpb_out[58][807],u_xpb_out[59][807],u_xpb_out[60][807],u_xpb_out[61][807],u_xpb_out[62][807],u_xpb_out[63][807],u_xpb_out[64][807],u_xpb_out[65][807],u_xpb_out[66][807],u_xpb_out[67][807],u_xpb_out[68][807],u_xpb_out[69][807],u_xpb_out[70][807],u_xpb_out[71][807],u_xpb_out[72][807],u_xpb_out[73][807],u_xpb_out[74][807],u_xpb_out[75][807],u_xpb_out[76][807],u_xpb_out[77][807],u_xpb_out[78][807],u_xpb_out[79][807],u_xpb_out[80][807],u_xpb_out[81][807],u_xpb_out[82][807],u_xpb_out[83][807],u_xpb_out[84][807],u_xpb_out[85][807],u_xpb_out[86][807],u_xpb_out[87][807],u_xpb_out[88][807],u_xpb_out[89][807],u_xpb_out[90][807],u_xpb_out[91][807],u_xpb_out[92][807],u_xpb_out[93][807],u_xpb_out[94][807],u_xpb_out[95][807],u_xpb_out[96][807],u_xpb_out[97][807],u_xpb_out[98][807],u_xpb_out[99][807],u_xpb_out[100][807],u_xpb_out[101][807],u_xpb_out[102][807],u_xpb_out[103][807],u_xpb_out[104][807],u_xpb_out[105][807]};

assign col_out_808 = {u_xpb_out[0][808],u_xpb_out[1][808],u_xpb_out[2][808],u_xpb_out[3][808],u_xpb_out[4][808],u_xpb_out[5][808],u_xpb_out[6][808],u_xpb_out[7][808],u_xpb_out[8][808],u_xpb_out[9][808],u_xpb_out[10][808],u_xpb_out[11][808],u_xpb_out[12][808],u_xpb_out[13][808],u_xpb_out[14][808],u_xpb_out[15][808],u_xpb_out[16][808],u_xpb_out[17][808],u_xpb_out[18][808],u_xpb_out[19][808],u_xpb_out[20][808],u_xpb_out[21][808],u_xpb_out[22][808],u_xpb_out[23][808],u_xpb_out[24][808],u_xpb_out[25][808],u_xpb_out[26][808],u_xpb_out[27][808],u_xpb_out[28][808],u_xpb_out[29][808],u_xpb_out[30][808],u_xpb_out[31][808],u_xpb_out[32][808],u_xpb_out[33][808],u_xpb_out[34][808],u_xpb_out[35][808],u_xpb_out[36][808],u_xpb_out[37][808],u_xpb_out[38][808],u_xpb_out[39][808],u_xpb_out[40][808],u_xpb_out[41][808],u_xpb_out[42][808],u_xpb_out[43][808],u_xpb_out[44][808],u_xpb_out[45][808],u_xpb_out[46][808],u_xpb_out[47][808],u_xpb_out[48][808],u_xpb_out[49][808],u_xpb_out[50][808],u_xpb_out[51][808],u_xpb_out[52][808],u_xpb_out[53][808],u_xpb_out[54][808],u_xpb_out[55][808],u_xpb_out[56][808],u_xpb_out[57][808],u_xpb_out[58][808],u_xpb_out[59][808],u_xpb_out[60][808],u_xpb_out[61][808],u_xpb_out[62][808],u_xpb_out[63][808],u_xpb_out[64][808],u_xpb_out[65][808],u_xpb_out[66][808],u_xpb_out[67][808],u_xpb_out[68][808],u_xpb_out[69][808],u_xpb_out[70][808],u_xpb_out[71][808],u_xpb_out[72][808],u_xpb_out[73][808],u_xpb_out[74][808],u_xpb_out[75][808],u_xpb_out[76][808],u_xpb_out[77][808],u_xpb_out[78][808],u_xpb_out[79][808],u_xpb_out[80][808],u_xpb_out[81][808],u_xpb_out[82][808],u_xpb_out[83][808],u_xpb_out[84][808],u_xpb_out[85][808],u_xpb_out[86][808],u_xpb_out[87][808],u_xpb_out[88][808],u_xpb_out[89][808],u_xpb_out[90][808],u_xpb_out[91][808],u_xpb_out[92][808],u_xpb_out[93][808],u_xpb_out[94][808],u_xpb_out[95][808],u_xpb_out[96][808],u_xpb_out[97][808],u_xpb_out[98][808],u_xpb_out[99][808],u_xpb_out[100][808],u_xpb_out[101][808],u_xpb_out[102][808],u_xpb_out[103][808],u_xpb_out[104][808],u_xpb_out[105][808]};

assign col_out_809 = {u_xpb_out[0][809],u_xpb_out[1][809],u_xpb_out[2][809],u_xpb_out[3][809],u_xpb_out[4][809],u_xpb_out[5][809],u_xpb_out[6][809],u_xpb_out[7][809],u_xpb_out[8][809],u_xpb_out[9][809],u_xpb_out[10][809],u_xpb_out[11][809],u_xpb_out[12][809],u_xpb_out[13][809],u_xpb_out[14][809],u_xpb_out[15][809],u_xpb_out[16][809],u_xpb_out[17][809],u_xpb_out[18][809],u_xpb_out[19][809],u_xpb_out[20][809],u_xpb_out[21][809],u_xpb_out[22][809],u_xpb_out[23][809],u_xpb_out[24][809],u_xpb_out[25][809],u_xpb_out[26][809],u_xpb_out[27][809],u_xpb_out[28][809],u_xpb_out[29][809],u_xpb_out[30][809],u_xpb_out[31][809],u_xpb_out[32][809],u_xpb_out[33][809],u_xpb_out[34][809],u_xpb_out[35][809],u_xpb_out[36][809],u_xpb_out[37][809],u_xpb_out[38][809],u_xpb_out[39][809],u_xpb_out[40][809],u_xpb_out[41][809],u_xpb_out[42][809],u_xpb_out[43][809],u_xpb_out[44][809],u_xpb_out[45][809],u_xpb_out[46][809],u_xpb_out[47][809],u_xpb_out[48][809],u_xpb_out[49][809],u_xpb_out[50][809],u_xpb_out[51][809],u_xpb_out[52][809],u_xpb_out[53][809],u_xpb_out[54][809],u_xpb_out[55][809],u_xpb_out[56][809],u_xpb_out[57][809],u_xpb_out[58][809],u_xpb_out[59][809],u_xpb_out[60][809],u_xpb_out[61][809],u_xpb_out[62][809],u_xpb_out[63][809],u_xpb_out[64][809],u_xpb_out[65][809],u_xpb_out[66][809],u_xpb_out[67][809],u_xpb_out[68][809],u_xpb_out[69][809],u_xpb_out[70][809],u_xpb_out[71][809],u_xpb_out[72][809],u_xpb_out[73][809],u_xpb_out[74][809],u_xpb_out[75][809],u_xpb_out[76][809],u_xpb_out[77][809],u_xpb_out[78][809],u_xpb_out[79][809],u_xpb_out[80][809],u_xpb_out[81][809],u_xpb_out[82][809],u_xpb_out[83][809],u_xpb_out[84][809],u_xpb_out[85][809],u_xpb_out[86][809],u_xpb_out[87][809],u_xpb_out[88][809],u_xpb_out[89][809],u_xpb_out[90][809],u_xpb_out[91][809],u_xpb_out[92][809],u_xpb_out[93][809],u_xpb_out[94][809],u_xpb_out[95][809],u_xpb_out[96][809],u_xpb_out[97][809],u_xpb_out[98][809],u_xpb_out[99][809],u_xpb_out[100][809],u_xpb_out[101][809],u_xpb_out[102][809],u_xpb_out[103][809],u_xpb_out[104][809],u_xpb_out[105][809]};

assign col_out_810 = {u_xpb_out[0][810],u_xpb_out[1][810],u_xpb_out[2][810],u_xpb_out[3][810],u_xpb_out[4][810],u_xpb_out[5][810],u_xpb_out[6][810],u_xpb_out[7][810],u_xpb_out[8][810],u_xpb_out[9][810],u_xpb_out[10][810],u_xpb_out[11][810],u_xpb_out[12][810],u_xpb_out[13][810],u_xpb_out[14][810],u_xpb_out[15][810],u_xpb_out[16][810],u_xpb_out[17][810],u_xpb_out[18][810],u_xpb_out[19][810],u_xpb_out[20][810],u_xpb_out[21][810],u_xpb_out[22][810],u_xpb_out[23][810],u_xpb_out[24][810],u_xpb_out[25][810],u_xpb_out[26][810],u_xpb_out[27][810],u_xpb_out[28][810],u_xpb_out[29][810],u_xpb_out[30][810],u_xpb_out[31][810],u_xpb_out[32][810],u_xpb_out[33][810],u_xpb_out[34][810],u_xpb_out[35][810],u_xpb_out[36][810],u_xpb_out[37][810],u_xpb_out[38][810],u_xpb_out[39][810],u_xpb_out[40][810],u_xpb_out[41][810],u_xpb_out[42][810],u_xpb_out[43][810],u_xpb_out[44][810],u_xpb_out[45][810],u_xpb_out[46][810],u_xpb_out[47][810],u_xpb_out[48][810],u_xpb_out[49][810],u_xpb_out[50][810],u_xpb_out[51][810],u_xpb_out[52][810],u_xpb_out[53][810],u_xpb_out[54][810],u_xpb_out[55][810],u_xpb_out[56][810],u_xpb_out[57][810],u_xpb_out[58][810],u_xpb_out[59][810],u_xpb_out[60][810],u_xpb_out[61][810],u_xpb_out[62][810],u_xpb_out[63][810],u_xpb_out[64][810],u_xpb_out[65][810],u_xpb_out[66][810],u_xpb_out[67][810],u_xpb_out[68][810],u_xpb_out[69][810],u_xpb_out[70][810],u_xpb_out[71][810],u_xpb_out[72][810],u_xpb_out[73][810],u_xpb_out[74][810],u_xpb_out[75][810],u_xpb_out[76][810],u_xpb_out[77][810],u_xpb_out[78][810],u_xpb_out[79][810],u_xpb_out[80][810],u_xpb_out[81][810],u_xpb_out[82][810],u_xpb_out[83][810],u_xpb_out[84][810],u_xpb_out[85][810],u_xpb_out[86][810],u_xpb_out[87][810],u_xpb_out[88][810],u_xpb_out[89][810],u_xpb_out[90][810],u_xpb_out[91][810],u_xpb_out[92][810],u_xpb_out[93][810],u_xpb_out[94][810],u_xpb_out[95][810],u_xpb_out[96][810],u_xpb_out[97][810],u_xpb_out[98][810],u_xpb_out[99][810],u_xpb_out[100][810],u_xpb_out[101][810],u_xpb_out[102][810],u_xpb_out[103][810],u_xpb_out[104][810],u_xpb_out[105][810]};

assign col_out_811 = {u_xpb_out[0][811],u_xpb_out[1][811],u_xpb_out[2][811],u_xpb_out[3][811],u_xpb_out[4][811],u_xpb_out[5][811],u_xpb_out[6][811],u_xpb_out[7][811],u_xpb_out[8][811],u_xpb_out[9][811],u_xpb_out[10][811],u_xpb_out[11][811],u_xpb_out[12][811],u_xpb_out[13][811],u_xpb_out[14][811],u_xpb_out[15][811],u_xpb_out[16][811],u_xpb_out[17][811],u_xpb_out[18][811],u_xpb_out[19][811],u_xpb_out[20][811],u_xpb_out[21][811],u_xpb_out[22][811],u_xpb_out[23][811],u_xpb_out[24][811],u_xpb_out[25][811],u_xpb_out[26][811],u_xpb_out[27][811],u_xpb_out[28][811],u_xpb_out[29][811],u_xpb_out[30][811],u_xpb_out[31][811],u_xpb_out[32][811],u_xpb_out[33][811],u_xpb_out[34][811],u_xpb_out[35][811],u_xpb_out[36][811],u_xpb_out[37][811],u_xpb_out[38][811],u_xpb_out[39][811],u_xpb_out[40][811],u_xpb_out[41][811],u_xpb_out[42][811],u_xpb_out[43][811],u_xpb_out[44][811],u_xpb_out[45][811],u_xpb_out[46][811],u_xpb_out[47][811],u_xpb_out[48][811],u_xpb_out[49][811],u_xpb_out[50][811],u_xpb_out[51][811],u_xpb_out[52][811],u_xpb_out[53][811],u_xpb_out[54][811],u_xpb_out[55][811],u_xpb_out[56][811],u_xpb_out[57][811],u_xpb_out[58][811],u_xpb_out[59][811],u_xpb_out[60][811],u_xpb_out[61][811],u_xpb_out[62][811],u_xpb_out[63][811],u_xpb_out[64][811],u_xpb_out[65][811],u_xpb_out[66][811],u_xpb_out[67][811],u_xpb_out[68][811],u_xpb_out[69][811],u_xpb_out[70][811],u_xpb_out[71][811],u_xpb_out[72][811],u_xpb_out[73][811],u_xpb_out[74][811],u_xpb_out[75][811],u_xpb_out[76][811],u_xpb_out[77][811],u_xpb_out[78][811],u_xpb_out[79][811],u_xpb_out[80][811],u_xpb_out[81][811],u_xpb_out[82][811],u_xpb_out[83][811],u_xpb_out[84][811],u_xpb_out[85][811],u_xpb_out[86][811],u_xpb_out[87][811],u_xpb_out[88][811],u_xpb_out[89][811],u_xpb_out[90][811],u_xpb_out[91][811],u_xpb_out[92][811],u_xpb_out[93][811],u_xpb_out[94][811],u_xpb_out[95][811],u_xpb_out[96][811],u_xpb_out[97][811],u_xpb_out[98][811],u_xpb_out[99][811],u_xpb_out[100][811],u_xpb_out[101][811],u_xpb_out[102][811],u_xpb_out[103][811],u_xpb_out[104][811],u_xpb_out[105][811]};

assign col_out_812 = {u_xpb_out[0][812],u_xpb_out[1][812],u_xpb_out[2][812],u_xpb_out[3][812],u_xpb_out[4][812],u_xpb_out[5][812],u_xpb_out[6][812],u_xpb_out[7][812],u_xpb_out[8][812],u_xpb_out[9][812],u_xpb_out[10][812],u_xpb_out[11][812],u_xpb_out[12][812],u_xpb_out[13][812],u_xpb_out[14][812],u_xpb_out[15][812],u_xpb_out[16][812],u_xpb_out[17][812],u_xpb_out[18][812],u_xpb_out[19][812],u_xpb_out[20][812],u_xpb_out[21][812],u_xpb_out[22][812],u_xpb_out[23][812],u_xpb_out[24][812],u_xpb_out[25][812],u_xpb_out[26][812],u_xpb_out[27][812],u_xpb_out[28][812],u_xpb_out[29][812],u_xpb_out[30][812],u_xpb_out[31][812],u_xpb_out[32][812],u_xpb_out[33][812],u_xpb_out[34][812],u_xpb_out[35][812],u_xpb_out[36][812],u_xpb_out[37][812],u_xpb_out[38][812],u_xpb_out[39][812],u_xpb_out[40][812],u_xpb_out[41][812],u_xpb_out[42][812],u_xpb_out[43][812],u_xpb_out[44][812],u_xpb_out[45][812],u_xpb_out[46][812],u_xpb_out[47][812],u_xpb_out[48][812],u_xpb_out[49][812],u_xpb_out[50][812],u_xpb_out[51][812],u_xpb_out[52][812],u_xpb_out[53][812],u_xpb_out[54][812],u_xpb_out[55][812],u_xpb_out[56][812],u_xpb_out[57][812],u_xpb_out[58][812],u_xpb_out[59][812],u_xpb_out[60][812],u_xpb_out[61][812],u_xpb_out[62][812],u_xpb_out[63][812],u_xpb_out[64][812],u_xpb_out[65][812],u_xpb_out[66][812],u_xpb_out[67][812],u_xpb_out[68][812],u_xpb_out[69][812],u_xpb_out[70][812],u_xpb_out[71][812],u_xpb_out[72][812],u_xpb_out[73][812],u_xpb_out[74][812],u_xpb_out[75][812],u_xpb_out[76][812],u_xpb_out[77][812],u_xpb_out[78][812],u_xpb_out[79][812],u_xpb_out[80][812],u_xpb_out[81][812],u_xpb_out[82][812],u_xpb_out[83][812],u_xpb_out[84][812],u_xpb_out[85][812],u_xpb_out[86][812],u_xpb_out[87][812],u_xpb_out[88][812],u_xpb_out[89][812],u_xpb_out[90][812],u_xpb_out[91][812],u_xpb_out[92][812],u_xpb_out[93][812],u_xpb_out[94][812],u_xpb_out[95][812],u_xpb_out[96][812],u_xpb_out[97][812],u_xpb_out[98][812],u_xpb_out[99][812],u_xpb_out[100][812],u_xpb_out[101][812],u_xpb_out[102][812],u_xpb_out[103][812],u_xpb_out[104][812],u_xpb_out[105][812]};

assign col_out_813 = {u_xpb_out[0][813],u_xpb_out[1][813],u_xpb_out[2][813],u_xpb_out[3][813],u_xpb_out[4][813],u_xpb_out[5][813],u_xpb_out[6][813],u_xpb_out[7][813],u_xpb_out[8][813],u_xpb_out[9][813],u_xpb_out[10][813],u_xpb_out[11][813],u_xpb_out[12][813],u_xpb_out[13][813],u_xpb_out[14][813],u_xpb_out[15][813],u_xpb_out[16][813],u_xpb_out[17][813],u_xpb_out[18][813],u_xpb_out[19][813],u_xpb_out[20][813],u_xpb_out[21][813],u_xpb_out[22][813],u_xpb_out[23][813],u_xpb_out[24][813],u_xpb_out[25][813],u_xpb_out[26][813],u_xpb_out[27][813],u_xpb_out[28][813],u_xpb_out[29][813],u_xpb_out[30][813],u_xpb_out[31][813],u_xpb_out[32][813],u_xpb_out[33][813],u_xpb_out[34][813],u_xpb_out[35][813],u_xpb_out[36][813],u_xpb_out[37][813],u_xpb_out[38][813],u_xpb_out[39][813],u_xpb_out[40][813],u_xpb_out[41][813],u_xpb_out[42][813],u_xpb_out[43][813],u_xpb_out[44][813],u_xpb_out[45][813],u_xpb_out[46][813],u_xpb_out[47][813],u_xpb_out[48][813],u_xpb_out[49][813],u_xpb_out[50][813],u_xpb_out[51][813],u_xpb_out[52][813],u_xpb_out[53][813],u_xpb_out[54][813],u_xpb_out[55][813],u_xpb_out[56][813],u_xpb_out[57][813],u_xpb_out[58][813],u_xpb_out[59][813],u_xpb_out[60][813],u_xpb_out[61][813],u_xpb_out[62][813],u_xpb_out[63][813],u_xpb_out[64][813],u_xpb_out[65][813],u_xpb_out[66][813],u_xpb_out[67][813],u_xpb_out[68][813],u_xpb_out[69][813],u_xpb_out[70][813],u_xpb_out[71][813],u_xpb_out[72][813],u_xpb_out[73][813],u_xpb_out[74][813],u_xpb_out[75][813],u_xpb_out[76][813],u_xpb_out[77][813],u_xpb_out[78][813],u_xpb_out[79][813],u_xpb_out[80][813],u_xpb_out[81][813],u_xpb_out[82][813],u_xpb_out[83][813],u_xpb_out[84][813],u_xpb_out[85][813],u_xpb_out[86][813],u_xpb_out[87][813],u_xpb_out[88][813],u_xpb_out[89][813],u_xpb_out[90][813],u_xpb_out[91][813],u_xpb_out[92][813],u_xpb_out[93][813],u_xpb_out[94][813],u_xpb_out[95][813],u_xpb_out[96][813],u_xpb_out[97][813],u_xpb_out[98][813],u_xpb_out[99][813],u_xpb_out[100][813],u_xpb_out[101][813],u_xpb_out[102][813],u_xpb_out[103][813],u_xpb_out[104][813],u_xpb_out[105][813]};

assign col_out_814 = {u_xpb_out[0][814],u_xpb_out[1][814],u_xpb_out[2][814],u_xpb_out[3][814],u_xpb_out[4][814],u_xpb_out[5][814],u_xpb_out[6][814],u_xpb_out[7][814],u_xpb_out[8][814],u_xpb_out[9][814],u_xpb_out[10][814],u_xpb_out[11][814],u_xpb_out[12][814],u_xpb_out[13][814],u_xpb_out[14][814],u_xpb_out[15][814],u_xpb_out[16][814],u_xpb_out[17][814],u_xpb_out[18][814],u_xpb_out[19][814],u_xpb_out[20][814],u_xpb_out[21][814],u_xpb_out[22][814],u_xpb_out[23][814],u_xpb_out[24][814],u_xpb_out[25][814],u_xpb_out[26][814],u_xpb_out[27][814],u_xpb_out[28][814],u_xpb_out[29][814],u_xpb_out[30][814],u_xpb_out[31][814],u_xpb_out[32][814],u_xpb_out[33][814],u_xpb_out[34][814],u_xpb_out[35][814],u_xpb_out[36][814],u_xpb_out[37][814],u_xpb_out[38][814],u_xpb_out[39][814],u_xpb_out[40][814],u_xpb_out[41][814],u_xpb_out[42][814],u_xpb_out[43][814],u_xpb_out[44][814],u_xpb_out[45][814],u_xpb_out[46][814],u_xpb_out[47][814],u_xpb_out[48][814],u_xpb_out[49][814],u_xpb_out[50][814],u_xpb_out[51][814],u_xpb_out[52][814],u_xpb_out[53][814],u_xpb_out[54][814],u_xpb_out[55][814],u_xpb_out[56][814],u_xpb_out[57][814],u_xpb_out[58][814],u_xpb_out[59][814],u_xpb_out[60][814],u_xpb_out[61][814],u_xpb_out[62][814],u_xpb_out[63][814],u_xpb_out[64][814],u_xpb_out[65][814],u_xpb_out[66][814],u_xpb_out[67][814],u_xpb_out[68][814],u_xpb_out[69][814],u_xpb_out[70][814],u_xpb_out[71][814],u_xpb_out[72][814],u_xpb_out[73][814],u_xpb_out[74][814],u_xpb_out[75][814],u_xpb_out[76][814],u_xpb_out[77][814],u_xpb_out[78][814],u_xpb_out[79][814],u_xpb_out[80][814],u_xpb_out[81][814],u_xpb_out[82][814],u_xpb_out[83][814],u_xpb_out[84][814],u_xpb_out[85][814],u_xpb_out[86][814],u_xpb_out[87][814],u_xpb_out[88][814],u_xpb_out[89][814],u_xpb_out[90][814],u_xpb_out[91][814],u_xpb_out[92][814],u_xpb_out[93][814],u_xpb_out[94][814],u_xpb_out[95][814],u_xpb_out[96][814],u_xpb_out[97][814],u_xpb_out[98][814],u_xpb_out[99][814],u_xpb_out[100][814],u_xpb_out[101][814],u_xpb_out[102][814],u_xpb_out[103][814],u_xpb_out[104][814],u_xpb_out[105][814]};

assign col_out_815 = {u_xpb_out[0][815],u_xpb_out[1][815],u_xpb_out[2][815],u_xpb_out[3][815],u_xpb_out[4][815],u_xpb_out[5][815],u_xpb_out[6][815],u_xpb_out[7][815],u_xpb_out[8][815],u_xpb_out[9][815],u_xpb_out[10][815],u_xpb_out[11][815],u_xpb_out[12][815],u_xpb_out[13][815],u_xpb_out[14][815],u_xpb_out[15][815],u_xpb_out[16][815],u_xpb_out[17][815],u_xpb_out[18][815],u_xpb_out[19][815],u_xpb_out[20][815],u_xpb_out[21][815],u_xpb_out[22][815],u_xpb_out[23][815],u_xpb_out[24][815],u_xpb_out[25][815],u_xpb_out[26][815],u_xpb_out[27][815],u_xpb_out[28][815],u_xpb_out[29][815],u_xpb_out[30][815],u_xpb_out[31][815],u_xpb_out[32][815],u_xpb_out[33][815],u_xpb_out[34][815],u_xpb_out[35][815],u_xpb_out[36][815],u_xpb_out[37][815],u_xpb_out[38][815],u_xpb_out[39][815],u_xpb_out[40][815],u_xpb_out[41][815],u_xpb_out[42][815],u_xpb_out[43][815],u_xpb_out[44][815],u_xpb_out[45][815],u_xpb_out[46][815],u_xpb_out[47][815],u_xpb_out[48][815],u_xpb_out[49][815],u_xpb_out[50][815],u_xpb_out[51][815],u_xpb_out[52][815],u_xpb_out[53][815],u_xpb_out[54][815],u_xpb_out[55][815],u_xpb_out[56][815],u_xpb_out[57][815],u_xpb_out[58][815],u_xpb_out[59][815],u_xpb_out[60][815],u_xpb_out[61][815],u_xpb_out[62][815],u_xpb_out[63][815],u_xpb_out[64][815],u_xpb_out[65][815],u_xpb_out[66][815],u_xpb_out[67][815],u_xpb_out[68][815],u_xpb_out[69][815],u_xpb_out[70][815],u_xpb_out[71][815],u_xpb_out[72][815],u_xpb_out[73][815],u_xpb_out[74][815],u_xpb_out[75][815],u_xpb_out[76][815],u_xpb_out[77][815],u_xpb_out[78][815],u_xpb_out[79][815],u_xpb_out[80][815],u_xpb_out[81][815],u_xpb_out[82][815],u_xpb_out[83][815],u_xpb_out[84][815],u_xpb_out[85][815],u_xpb_out[86][815],u_xpb_out[87][815],u_xpb_out[88][815],u_xpb_out[89][815],u_xpb_out[90][815],u_xpb_out[91][815],u_xpb_out[92][815],u_xpb_out[93][815],u_xpb_out[94][815],u_xpb_out[95][815],u_xpb_out[96][815],u_xpb_out[97][815],u_xpb_out[98][815],u_xpb_out[99][815],u_xpb_out[100][815],u_xpb_out[101][815],u_xpb_out[102][815],u_xpb_out[103][815],u_xpb_out[104][815],u_xpb_out[105][815]};

assign col_out_816 = {u_xpb_out[0][816],u_xpb_out[1][816],u_xpb_out[2][816],u_xpb_out[3][816],u_xpb_out[4][816],u_xpb_out[5][816],u_xpb_out[6][816],u_xpb_out[7][816],u_xpb_out[8][816],u_xpb_out[9][816],u_xpb_out[10][816],u_xpb_out[11][816],u_xpb_out[12][816],u_xpb_out[13][816],u_xpb_out[14][816],u_xpb_out[15][816],u_xpb_out[16][816],u_xpb_out[17][816],u_xpb_out[18][816],u_xpb_out[19][816],u_xpb_out[20][816],u_xpb_out[21][816],u_xpb_out[22][816],u_xpb_out[23][816],u_xpb_out[24][816],u_xpb_out[25][816],u_xpb_out[26][816],u_xpb_out[27][816],u_xpb_out[28][816],u_xpb_out[29][816],u_xpb_out[30][816],u_xpb_out[31][816],u_xpb_out[32][816],u_xpb_out[33][816],u_xpb_out[34][816],u_xpb_out[35][816],u_xpb_out[36][816],u_xpb_out[37][816],u_xpb_out[38][816],u_xpb_out[39][816],u_xpb_out[40][816],u_xpb_out[41][816],u_xpb_out[42][816],u_xpb_out[43][816],u_xpb_out[44][816],u_xpb_out[45][816],u_xpb_out[46][816],u_xpb_out[47][816],u_xpb_out[48][816],u_xpb_out[49][816],u_xpb_out[50][816],u_xpb_out[51][816],u_xpb_out[52][816],u_xpb_out[53][816],u_xpb_out[54][816],u_xpb_out[55][816],u_xpb_out[56][816],u_xpb_out[57][816],u_xpb_out[58][816],u_xpb_out[59][816],u_xpb_out[60][816],u_xpb_out[61][816],u_xpb_out[62][816],u_xpb_out[63][816],u_xpb_out[64][816],u_xpb_out[65][816],u_xpb_out[66][816],u_xpb_out[67][816],u_xpb_out[68][816],u_xpb_out[69][816],u_xpb_out[70][816],u_xpb_out[71][816],u_xpb_out[72][816],u_xpb_out[73][816],u_xpb_out[74][816],u_xpb_out[75][816],u_xpb_out[76][816],u_xpb_out[77][816],u_xpb_out[78][816],u_xpb_out[79][816],u_xpb_out[80][816],u_xpb_out[81][816],u_xpb_out[82][816],u_xpb_out[83][816],u_xpb_out[84][816],u_xpb_out[85][816],u_xpb_out[86][816],u_xpb_out[87][816],u_xpb_out[88][816],u_xpb_out[89][816],u_xpb_out[90][816],u_xpb_out[91][816],u_xpb_out[92][816],u_xpb_out[93][816],u_xpb_out[94][816],u_xpb_out[95][816],u_xpb_out[96][816],u_xpb_out[97][816],u_xpb_out[98][816],u_xpb_out[99][816],u_xpb_out[100][816],u_xpb_out[101][816],u_xpb_out[102][816],u_xpb_out[103][816],u_xpb_out[104][816],u_xpb_out[105][816]};

assign col_out_817 = {u_xpb_out[0][817],u_xpb_out[1][817],u_xpb_out[2][817],u_xpb_out[3][817],u_xpb_out[4][817],u_xpb_out[5][817],u_xpb_out[6][817],u_xpb_out[7][817],u_xpb_out[8][817],u_xpb_out[9][817],u_xpb_out[10][817],u_xpb_out[11][817],u_xpb_out[12][817],u_xpb_out[13][817],u_xpb_out[14][817],u_xpb_out[15][817],u_xpb_out[16][817],u_xpb_out[17][817],u_xpb_out[18][817],u_xpb_out[19][817],u_xpb_out[20][817],u_xpb_out[21][817],u_xpb_out[22][817],u_xpb_out[23][817],u_xpb_out[24][817],u_xpb_out[25][817],u_xpb_out[26][817],u_xpb_out[27][817],u_xpb_out[28][817],u_xpb_out[29][817],u_xpb_out[30][817],u_xpb_out[31][817],u_xpb_out[32][817],u_xpb_out[33][817],u_xpb_out[34][817],u_xpb_out[35][817],u_xpb_out[36][817],u_xpb_out[37][817],u_xpb_out[38][817],u_xpb_out[39][817],u_xpb_out[40][817],u_xpb_out[41][817],u_xpb_out[42][817],u_xpb_out[43][817],u_xpb_out[44][817],u_xpb_out[45][817],u_xpb_out[46][817],u_xpb_out[47][817],u_xpb_out[48][817],u_xpb_out[49][817],u_xpb_out[50][817],u_xpb_out[51][817],u_xpb_out[52][817],u_xpb_out[53][817],u_xpb_out[54][817],u_xpb_out[55][817],u_xpb_out[56][817],u_xpb_out[57][817],u_xpb_out[58][817],u_xpb_out[59][817],u_xpb_out[60][817],u_xpb_out[61][817],u_xpb_out[62][817],u_xpb_out[63][817],u_xpb_out[64][817],u_xpb_out[65][817],u_xpb_out[66][817],u_xpb_out[67][817],u_xpb_out[68][817],u_xpb_out[69][817],u_xpb_out[70][817],u_xpb_out[71][817],u_xpb_out[72][817],u_xpb_out[73][817],u_xpb_out[74][817],u_xpb_out[75][817],u_xpb_out[76][817],u_xpb_out[77][817],u_xpb_out[78][817],u_xpb_out[79][817],u_xpb_out[80][817],u_xpb_out[81][817],u_xpb_out[82][817],u_xpb_out[83][817],u_xpb_out[84][817],u_xpb_out[85][817],u_xpb_out[86][817],u_xpb_out[87][817],u_xpb_out[88][817],u_xpb_out[89][817],u_xpb_out[90][817],u_xpb_out[91][817],u_xpb_out[92][817],u_xpb_out[93][817],u_xpb_out[94][817],u_xpb_out[95][817],u_xpb_out[96][817],u_xpb_out[97][817],u_xpb_out[98][817],u_xpb_out[99][817],u_xpb_out[100][817],u_xpb_out[101][817],u_xpb_out[102][817],u_xpb_out[103][817],u_xpb_out[104][817],u_xpb_out[105][817]};

assign col_out_818 = {u_xpb_out[0][818],u_xpb_out[1][818],u_xpb_out[2][818],u_xpb_out[3][818],u_xpb_out[4][818],u_xpb_out[5][818],u_xpb_out[6][818],u_xpb_out[7][818],u_xpb_out[8][818],u_xpb_out[9][818],u_xpb_out[10][818],u_xpb_out[11][818],u_xpb_out[12][818],u_xpb_out[13][818],u_xpb_out[14][818],u_xpb_out[15][818],u_xpb_out[16][818],u_xpb_out[17][818],u_xpb_out[18][818],u_xpb_out[19][818],u_xpb_out[20][818],u_xpb_out[21][818],u_xpb_out[22][818],u_xpb_out[23][818],u_xpb_out[24][818],u_xpb_out[25][818],u_xpb_out[26][818],u_xpb_out[27][818],u_xpb_out[28][818],u_xpb_out[29][818],u_xpb_out[30][818],u_xpb_out[31][818],u_xpb_out[32][818],u_xpb_out[33][818],u_xpb_out[34][818],u_xpb_out[35][818],u_xpb_out[36][818],u_xpb_out[37][818],u_xpb_out[38][818],u_xpb_out[39][818],u_xpb_out[40][818],u_xpb_out[41][818],u_xpb_out[42][818],u_xpb_out[43][818],u_xpb_out[44][818],u_xpb_out[45][818],u_xpb_out[46][818],u_xpb_out[47][818],u_xpb_out[48][818],u_xpb_out[49][818],u_xpb_out[50][818],u_xpb_out[51][818],u_xpb_out[52][818],u_xpb_out[53][818],u_xpb_out[54][818],u_xpb_out[55][818],u_xpb_out[56][818],u_xpb_out[57][818],u_xpb_out[58][818],u_xpb_out[59][818],u_xpb_out[60][818],u_xpb_out[61][818],u_xpb_out[62][818],u_xpb_out[63][818],u_xpb_out[64][818],u_xpb_out[65][818],u_xpb_out[66][818],u_xpb_out[67][818],u_xpb_out[68][818],u_xpb_out[69][818],u_xpb_out[70][818],u_xpb_out[71][818],u_xpb_out[72][818],u_xpb_out[73][818],u_xpb_out[74][818],u_xpb_out[75][818],u_xpb_out[76][818],u_xpb_out[77][818],u_xpb_out[78][818],u_xpb_out[79][818],u_xpb_out[80][818],u_xpb_out[81][818],u_xpb_out[82][818],u_xpb_out[83][818],u_xpb_out[84][818],u_xpb_out[85][818],u_xpb_out[86][818],u_xpb_out[87][818],u_xpb_out[88][818],u_xpb_out[89][818],u_xpb_out[90][818],u_xpb_out[91][818],u_xpb_out[92][818],u_xpb_out[93][818],u_xpb_out[94][818],u_xpb_out[95][818],u_xpb_out[96][818],u_xpb_out[97][818],u_xpb_out[98][818],u_xpb_out[99][818],u_xpb_out[100][818],u_xpb_out[101][818],u_xpb_out[102][818],u_xpb_out[103][818],u_xpb_out[104][818],u_xpb_out[105][818]};

assign col_out_819 = {u_xpb_out[0][819],u_xpb_out[1][819],u_xpb_out[2][819],u_xpb_out[3][819],u_xpb_out[4][819],u_xpb_out[5][819],u_xpb_out[6][819],u_xpb_out[7][819],u_xpb_out[8][819],u_xpb_out[9][819],u_xpb_out[10][819],u_xpb_out[11][819],u_xpb_out[12][819],u_xpb_out[13][819],u_xpb_out[14][819],u_xpb_out[15][819],u_xpb_out[16][819],u_xpb_out[17][819],u_xpb_out[18][819],u_xpb_out[19][819],u_xpb_out[20][819],u_xpb_out[21][819],u_xpb_out[22][819],u_xpb_out[23][819],u_xpb_out[24][819],u_xpb_out[25][819],u_xpb_out[26][819],u_xpb_out[27][819],u_xpb_out[28][819],u_xpb_out[29][819],u_xpb_out[30][819],u_xpb_out[31][819],u_xpb_out[32][819],u_xpb_out[33][819],u_xpb_out[34][819],u_xpb_out[35][819],u_xpb_out[36][819],u_xpb_out[37][819],u_xpb_out[38][819],u_xpb_out[39][819],u_xpb_out[40][819],u_xpb_out[41][819],u_xpb_out[42][819],u_xpb_out[43][819],u_xpb_out[44][819],u_xpb_out[45][819],u_xpb_out[46][819],u_xpb_out[47][819],u_xpb_out[48][819],u_xpb_out[49][819],u_xpb_out[50][819],u_xpb_out[51][819],u_xpb_out[52][819],u_xpb_out[53][819],u_xpb_out[54][819],u_xpb_out[55][819],u_xpb_out[56][819],u_xpb_out[57][819],u_xpb_out[58][819],u_xpb_out[59][819],u_xpb_out[60][819],u_xpb_out[61][819],u_xpb_out[62][819],u_xpb_out[63][819],u_xpb_out[64][819],u_xpb_out[65][819],u_xpb_out[66][819],u_xpb_out[67][819],u_xpb_out[68][819],u_xpb_out[69][819],u_xpb_out[70][819],u_xpb_out[71][819],u_xpb_out[72][819],u_xpb_out[73][819],u_xpb_out[74][819],u_xpb_out[75][819],u_xpb_out[76][819],u_xpb_out[77][819],u_xpb_out[78][819],u_xpb_out[79][819],u_xpb_out[80][819],u_xpb_out[81][819],u_xpb_out[82][819],u_xpb_out[83][819],u_xpb_out[84][819],u_xpb_out[85][819],u_xpb_out[86][819],u_xpb_out[87][819],u_xpb_out[88][819],u_xpb_out[89][819],u_xpb_out[90][819],u_xpb_out[91][819],u_xpb_out[92][819],u_xpb_out[93][819],u_xpb_out[94][819],u_xpb_out[95][819],u_xpb_out[96][819],u_xpb_out[97][819],u_xpb_out[98][819],u_xpb_out[99][819],u_xpb_out[100][819],u_xpb_out[101][819],u_xpb_out[102][819],u_xpb_out[103][819],u_xpb_out[104][819],u_xpb_out[105][819]};

assign col_out_820 = {u_xpb_out[0][820],u_xpb_out[1][820],u_xpb_out[2][820],u_xpb_out[3][820],u_xpb_out[4][820],u_xpb_out[5][820],u_xpb_out[6][820],u_xpb_out[7][820],u_xpb_out[8][820],u_xpb_out[9][820],u_xpb_out[10][820],u_xpb_out[11][820],u_xpb_out[12][820],u_xpb_out[13][820],u_xpb_out[14][820],u_xpb_out[15][820],u_xpb_out[16][820],u_xpb_out[17][820],u_xpb_out[18][820],u_xpb_out[19][820],u_xpb_out[20][820],u_xpb_out[21][820],u_xpb_out[22][820],u_xpb_out[23][820],u_xpb_out[24][820],u_xpb_out[25][820],u_xpb_out[26][820],u_xpb_out[27][820],u_xpb_out[28][820],u_xpb_out[29][820],u_xpb_out[30][820],u_xpb_out[31][820],u_xpb_out[32][820],u_xpb_out[33][820],u_xpb_out[34][820],u_xpb_out[35][820],u_xpb_out[36][820],u_xpb_out[37][820],u_xpb_out[38][820],u_xpb_out[39][820],u_xpb_out[40][820],u_xpb_out[41][820],u_xpb_out[42][820],u_xpb_out[43][820],u_xpb_out[44][820],u_xpb_out[45][820],u_xpb_out[46][820],u_xpb_out[47][820],u_xpb_out[48][820],u_xpb_out[49][820],u_xpb_out[50][820],u_xpb_out[51][820],u_xpb_out[52][820],u_xpb_out[53][820],u_xpb_out[54][820],u_xpb_out[55][820],u_xpb_out[56][820],u_xpb_out[57][820],u_xpb_out[58][820],u_xpb_out[59][820],u_xpb_out[60][820],u_xpb_out[61][820],u_xpb_out[62][820],u_xpb_out[63][820],u_xpb_out[64][820],u_xpb_out[65][820],u_xpb_out[66][820],u_xpb_out[67][820],u_xpb_out[68][820],u_xpb_out[69][820],u_xpb_out[70][820],u_xpb_out[71][820],u_xpb_out[72][820],u_xpb_out[73][820],u_xpb_out[74][820],u_xpb_out[75][820],u_xpb_out[76][820],u_xpb_out[77][820],u_xpb_out[78][820],u_xpb_out[79][820],u_xpb_out[80][820],u_xpb_out[81][820],u_xpb_out[82][820],u_xpb_out[83][820],u_xpb_out[84][820],u_xpb_out[85][820],u_xpb_out[86][820],u_xpb_out[87][820],u_xpb_out[88][820],u_xpb_out[89][820],u_xpb_out[90][820],u_xpb_out[91][820],u_xpb_out[92][820],u_xpb_out[93][820],u_xpb_out[94][820],u_xpb_out[95][820],u_xpb_out[96][820],u_xpb_out[97][820],u_xpb_out[98][820],u_xpb_out[99][820],u_xpb_out[100][820],u_xpb_out[101][820],u_xpb_out[102][820],u_xpb_out[103][820],u_xpb_out[104][820],u_xpb_out[105][820]};

assign col_out_821 = {u_xpb_out[0][821],u_xpb_out[1][821],u_xpb_out[2][821],u_xpb_out[3][821],u_xpb_out[4][821],u_xpb_out[5][821],u_xpb_out[6][821],u_xpb_out[7][821],u_xpb_out[8][821],u_xpb_out[9][821],u_xpb_out[10][821],u_xpb_out[11][821],u_xpb_out[12][821],u_xpb_out[13][821],u_xpb_out[14][821],u_xpb_out[15][821],u_xpb_out[16][821],u_xpb_out[17][821],u_xpb_out[18][821],u_xpb_out[19][821],u_xpb_out[20][821],u_xpb_out[21][821],u_xpb_out[22][821],u_xpb_out[23][821],u_xpb_out[24][821],u_xpb_out[25][821],u_xpb_out[26][821],u_xpb_out[27][821],u_xpb_out[28][821],u_xpb_out[29][821],u_xpb_out[30][821],u_xpb_out[31][821],u_xpb_out[32][821],u_xpb_out[33][821],u_xpb_out[34][821],u_xpb_out[35][821],u_xpb_out[36][821],u_xpb_out[37][821],u_xpb_out[38][821],u_xpb_out[39][821],u_xpb_out[40][821],u_xpb_out[41][821],u_xpb_out[42][821],u_xpb_out[43][821],u_xpb_out[44][821],u_xpb_out[45][821],u_xpb_out[46][821],u_xpb_out[47][821],u_xpb_out[48][821],u_xpb_out[49][821],u_xpb_out[50][821],u_xpb_out[51][821],u_xpb_out[52][821],u_xpb_out[53][821],u_xpb_out[54][821],u_xpb_out[55][821],u_xpb_out[56][821],u_xpb_out[57][821],u_xpb_out[58][821],u_xpb_out[59][821],u_xpb_out[60][821],u_xpb_out[61][821],u_xpb_out[62][821],u_xpb_out[63][821],u_xpb_out[64][821],u_xpb_out[65][821],u_xpb_out[66][821],u_xpb_out[67][821],u_xpb_out[68][821],u_xpb_out[69][821],u_xpb_out[70][821],u_xpb_out[71][821],u_xpb_out[72][821],u_xpb_out[73][821],u_xpb_out[74][821],u_xpb_out[75][821],u_xpb_out[76][821],u_xpb_out[77][821],u_xpb_out[78][821],u_xpb_out[79][821],u_xpb_out[80][821],u_xpb_out[81][821],u_xpb_out[82][821],u_xpb_out[83][821],u_xpb_out[84][821],u_xpb_out[85][821],u_xpb_out[86][821],u_xpb_out[87][821],u_xpb_out[88][821],u_xpb_out[89][821],u_xpb_out[90][821],u_xpb_out[91][821],u_xpb_out[92][821],u_xpb_out[93][821],u_xpb_out[94][821],u_xpb_out[95][821],u_xpb_out[96][821],u_xpb_out[97][821],u_xpb_out[98][821],u_xpb_out[99][821],u_xpb_out[100][821],u_xpb_out[101][821],u_xpb_out[102][821],u_xpb_out[103][821],u_xpb_out[104][821],u_xpb_out[105][821]};

assign col_out_822 = {u_xpb_out[0][822],u_xpb_out[1][822],u_xpb_out[2][822],u_xpb_out[3][822],u_xpb_out[4][822],u_xpb_out[5][822],u_xpb_out[6][822],u_xpb_out[7][822],u_xpb_out[8][822],u_xpb_out[9][822],u_xpb_out[10][822],u_xpb_out[11][822],u_xpb_out[12][822],u_xpb_out[13][822],u_xpb_out[14][822],u_xpb_out[15][822],u_xpb_out[16][822],u_xpb_out[17][822],u_xpb_out[18][822],u_xpb_out[19][822],u_xpb_out[20][822],u_xpb_out[21][822],u_xpb_out[22][822],u_xpb_out[23][822],u_xpb_out[24][822],u_xpb_out[25][822],u_xpb_out[26][822],u_xpb_out[27][822],u_xpb_out[28][822],u_xpb_out[29][822],u_xpb_out[30][822],u_xpb_out[31][822],u_xpb_out[32][822],u_xpb_out[33][822],u_xpb_out[34][822],u_xpb_out[35][822],u_xpb_out[36][822],u_xpb_out[37][822],u_xpb_out[38][822],u_xpb_out[39][822],u_xpb_out[40][822],u_xpb_out[41][822],u_xpb_out[42][822],u_xpb_out[43][822],u_xpb_out[44][822],u_xpb_out[45][822],u_xpb_out[46][822],u_xpb_out[47][822],u_xpb_out[48][822],u_xpb_out[49][822],u_xpb_out[50][822],u_xpb_out[51][822],u_xpb_out[52][822],u_xpb_out[53][822],u_xpb_out[54][822],u_xpb_out[55][822],u_xpb_out[56][822],u_xpb_out[57][822],u_xpb_out[58][822],u_xpb_out[59][822],u_xpb_out[60][822],u_xpb_out[61][822],u_xpb_out[62][822],u_xpb_out[63][822],u_xpb_out[64][822],u_xpb_out[65][822],u_xpb_out[66][822],u_xpb_out[67][822],u_xpb_out[68][822],u_xpb_out[69][822],u_xpb_out[70][822],u_xpb_out[71][822],u_xpb_out[72][822],u_xpb_out[73][822],u_xpb_out[74][822],u_xpb_out[75][822],u_xpb_out[76][822],u_xpb_out[77][822],u_xpb_out[78][822],u_xpb_out[79][822],u_xpb_out[80][822],u_xpb_out[81][822],u_xpb_out[82][822],u_xpb_out[83][822],u_xpb_out[84][822],u_xpb_out[85][822],u_xpb_out[86][822],u_xpb_out[87][822],u_xpb_out[88][822],u_xpb_out[89][822],u_xpb_out[90][822],u_xpb_out[91][822],u_xpb_out[92][822],u_xpb_out[93][822],u_xpb_out[94][822],u_xpb_out[95][822],u_xpb_out[96][822],u_xpb_out[97][822],u_xpb_out[98][822],u_xpb_out[99][822],u_xpb_out[100][822],u_xpb_out[101][822],u_xpb_out[102][822],u_xpb_out[103][822],u_xpb_out[104][822],u_xpb_out[105][822]};

assign col_out_823 = {u_xpb_out[0][823],u_xpb_out[1][823],u_xpb_out[2][823],u_xpb_out[3][823],u_xpb_out[4][823],u_xpb_out[5][823],u_xpb_out[6][823],u_xpb_out[7][823],u_xpb_out[8][823],u_xpb_out[9][823],u_xpb_out[10][823],u_xpb_out[11][823],u_xpb_out[12][823],u_xpb_out[13][823],u_xpb_out[14][823],u_xpb_out[15][823],u_xpb_out[16][823],u_xpb_out[17][823],u_xpb_out[18][823],u_xpb_out[19][823],u_xpb_out[20][823],u_xpb_out[21][823],u_xpb_out[22][823],u_xpb_out[23][823],u_xpb_out[24][823],u_xpb_out[25][823],u_xpb_out[26][823],u_xpb_out[27][823],u_xpb_out[28][823],u_xpb_out[29][823],u_xpb_out[30][823],u_xpb_out[31][823],u_xpb_out[32][823],u_xpb_out[33][823],u_xpb_out[34][823],u_xpb_out[35][823],u_xpb_out[36][823],u_xpb_out[37][823],u_xpb_out[38][823],u_xpb_out[39][823],u_xpb_out[40][823],u_xpb_out[41][823],u_xpb_out[42][823],u_xpb_out[43][823],u_xpb_out[44][823],u_xpb_out[45][823],u_xpb_out[46][823],u_xpb_out[47][823],u_xpb_out[48][823],u_xpb_out[49][823],u_xpb_out[50][823],u_xpb_out[51][823],u_xpb_out[52][823],u_xpb_out[53][823],u_xpb_out[54][823],u_xpb_out[55][823],u_xpb_out[56][823],u_xpb_out[57][823],u_xpb_out[58][823],u_xpb_out[59][823],u_xpb_out[60][823],u_xpb_out[61][823],u_xpb_out[62][823],u_xpb_out[63][823],u_xpb_out[64][823],u_xpb_out[65][823],u_xpb_out[66][823],u_xpb_out[67][823],u_xpb_out[68][823],u_xpb_out[69][823],u_xpb_out[70][823],u_xpb_out[71][823],u_xpb_out[72][823],u_xpb_out[73][823],u_xpb_out[74][823],u_xpb_out[75][823],u_xpb_out[76][823],u_xpb_out[77][823],u_xpb_out[78][823],u_xpb_out[79][823],u_xpb_out[80][823],u_xpb_out[81][823],u_xpb_out[82][823],u_xpb_out[83][823],u_xpb_out[84][823],u_xpb_out[85][823],u_xpb_out[86][823],u_xpb_out[87][823],u_xpb_out[88][823],u_xpb_out[89][823],u_xpb_out[90][823],u_xpb_out[91][823],u_xpb_out[92][823],u_xpb_out[93][823],u_xpb_out[94][823],u_xpb_out[95][823],u_xpb_out[96][823],u_xpb_out[97][823],u_xpb_out[98][823],u_xpb_out[99][823],u_xpb_out[100][823],u_xpb_out[101][823],u_xpb_out[102][823],u_xpb_out[103][823],u_xpb_out[104][823],u_xpb_out[105][823]};

assign col_out_824 = {u_xpb_out[0][824],u_xpb_out[1][824],u_xpb_out[2][824],u_xpb_out[3][824],u_xpb_out[4][824],u_xpb_out[5][824],u_xpb_out[6][824],u_xpb_out[7][824],u_xpb_out[8][824],u_xpb_out[9][824],u_xpb_out[10][824],u_xpb_out[11][824],u_xpb_out[12][824],u_xpb_out[13][824],u_xpb_out[14][824],u_xpb_out[15][824],u_xpb_out[16][824],u_xpb_out[17][824],u_xpb_out[18][824],u_xpb_out[19][824],u_xpb_out[20][824],u_xpb_out[21][824],u_xpb_out[22][824],u_xpb_out[23][824],u_xpb_out[24][824],u_xpb_out[25][824],u_xpb_out[26][824],u_xpb_out[27][824],u_xpb_out[28][824],u_xpb_out[29][824],u_xpb_out[30][824],u_xpb_out[31][824],u_xpb_out[32][824],u_xpb_out[33][824],u_xpb_out[34][824],u_xpb_out[35][824],u_xpb_out[36][824],u_xpb_out[37][824],u_xpb_out[38][824],u_xpb_out[39][824],u_xpb_out[40][824],u_xpb_out[41][824],u_xpb_out[42][824],u_xpb_out[43][824],u_xpb_out[44][824],u_xpb_out[45][824],u_xpb_out[46][824],u_xpb_out[47][824],u_xpb_out[48][824],u_xpb_out[49][824],u_xpb_out[50][824],u_xpb_out[51][824],u_xpb_out[52][824],u_xpb_out[53][824],u_xpb_out[54][824],u_xpb_out[55][824],u_xpb_out[56][824],u_xpb_out[57][824],u_xpb_out[58][824],u_xpb_out[59][824],u_xpb_out[60][824],u_xpb_out[61][824],u_xpb_out[62][824],u_xpb_out[63][824],u_xpb_out[64][824],u_xpb_out[65][824],u_xpb_out[66][824],u_xpb_out[67][824],u_xpb_out[68][824],u_xpb_out[69][824],u_xpb_out[70][824],u_xpb_out[71][824],u_xpb_out[72][824],u_xpb_out[73][824],u_xpb_out[74][824],u_xpb_out[75][824],u_xpb_out[76][824],u_xpb_out[77][824],u_xpb_out[78][824],u_xpb_out[79][824],u_xpb_out[80][824],u_xpb_out[81][824],u_xpb_out[82][824],u_xpb_out[83][824],u_xpb_out[84][824],u_xpb_out[85][824],u_xpb_out[86][824],u_xpb_out[87][824],u_xpb_out[88][824],u_xpb_out[89][824],u_xpb_out[90][824],u_xpb_out[91][824],u_xpb_out[92][824],u_xpb_out[93][824],u_xpb_out[94][824],u_xpb_out[95][824],u_xpb_out[96][824],u_xpb_out[97][824],u_xpb_out[98][824],u_xpb_out[99][824],u_xpb_out[100][824],u_xpb_out[101][824],u_xpb_out[102][824],u_xpb_out[103][824],u_xpb_out[104][824],u_xpb_out[105][824]};

assign col_out_825 = {u_xpb_out[0][825],u_xpb_out[1][825],u_xpb_out[2][825],u_xpb_out[3][825],u_xpb_out[4][825],u_xpb_out[5][825],u_xpb_out[6][825],u_xpb_out[7][825],u_xpb_out[8][825],u_xpb_out[9][825],u_xpb_out[10][825],u_xpb_out[11][825],u_xpb_out[12][825],u_xpb_out[13][825],u_xpb_out[14][825],u_xpb_out[15][825],u_xpb_out[16][825],u_xpb_out[17][825],u_xpb_out[18][825],u_xpb_out[19][825],u_xpb_out[20][825],u_xpb_out[21][825],u_xpb_out[22][825],u_xpb_out[23][825],u_xpb_out[24][825],u_xpb_out[25][825],u_xpb_out[26][825],u_xpb_out[27][825],u_xpb_out[28][825],u_xpb_out[29][825],u_xpb_out[30][825],u_xpb_out[31][825],u_xpb_out[32][825],u_xpb_out[33][825],u_xpb_out[34][825],u_xpb_out[35][825],u_xpb_out[36][825],u_xpb_out[37][825],u_xpb_out[38][825],u_xpb_out[39][825],u_xpb_out[40][825],u_xpb_out[41][825],u_xpb_out[42][825],u_xpb_out[43][825],u_xpb_out[44][825],u_xpb_out[45][825],u_xpb_out[46][825],u_xpb_out[47][825],u_xpb_out[48][825],u_xpb_out[49][825],u_xpb_out[50][825],u_xpb_out[51][825],u_xpb_out[52][825],u_xpb_out[53][825],u_xpb_out[54][825],u_xpb_out[55][825],u_xpb_out[56][825],u_xpb_out[57][825],u_xpb_out[58][825],u_xpb_out[59][825],u_xpb_out[60][825],u_xpb_out[61][825],u_xpb_out[62][825],u_xpb_out[63][825],u_xpb_out[64][825],u_xpb_out[65][825],u_xpb_out[66][825],u_xpb_out[67][825],u_xpb_out[68][825],u_xpb_out[69][825],u_xpb_out[70][825],u_xpb_out[71][825],u_xpb_out[72][825],u_xpb_out[73][825],u_xpb_out[74][825],u_xpb_out[75][825],u_xpb_out[76][825],u_xpb_out[77][825],u_xpb_out[78][825],u_xpb_out[79][825],u_xpb_out[80][825],u_xpb_out[81][825],u_xpb_out[82][825],u_xpb_out[83][825],u_xpb_out[84][825],u_xpb_out[85][825],u_xpb_out[86][825],u_xpb_out[87][825],u_xpb_out[88][825],u_xpb_out[89][825],u_xpb_out[90][825],u_xpb_out[91][825],u_xpb_out[92][825],u_xpb_out[93][825],u_xpb_out[94][825],u_xpb_out[95][825],u_xpb_out[96][825],u_xpb_out[97][825],u_xpb_out[98][825],u_xpb_out[99][825],u_xpb_out[100][825],u_xpb_out[101][825],u_xpb_out[102][825],u_xpb_out[103][825],u_xpb_out[104][825],u_xpb_out[105][825]};

assign col_out_826 = {u_xpb_out[0][826],u_xpb_out[1][826],u_xpb_out[2][826],u_xpb_out[3][826],u_xpb_out[4][826],u_xpb_out[5][826],u_xpb_out[6][826],u_xpb_out[7][826],u_xpb_out[8][826],u_xpb_out[9][826],u_xpb_out[10][826],u_xpb_out[11][826],u_xpb_out[12][826],u_xpb_out[13][826],u_xpb_out[14][826],u_xpb_out[15][826],u_xpb_out[16][826],u_xpb_out[17][826],u_xpb_out[18][826],u_xpb_out[19][826],u_xpb_out[20][826],u_xpb_out[21][826],u_xpb_out[22][826],u_xpb_out[23][826],u_xpb_out[24][826],u_xpb_out[25][826],u_xpb_out[26][826],u_xpb_out[27][826],u_xpb_out[28][826],u_xpb_out[29][826],u_xpb_out[30][826],u_xpb_out[31][826],u_xpb_out[32][826],u_xpb_out[33][826],u_xpb_out[34][826],u_xpb_out[35][826],u_xpb_out[36][826],u_xpb_out[37][826],u_xpb_out[38][826],u_xpb_out[39][826],u_xpb_out[40][826],u_xpb_out[41][826],u_xpb_out[42][826],u_xpb_out[43][826],u_xpb_out[44][826],u_xpb_out[45][826],u_xpb_out[46][826],u_xpb_out[47][826],u_xpb_out[48][826],u_xpb_out[49][826],u_xpb_out[50][826],u_xpb_out[51][826],u_xpb_out[52][826],u_xpb_out[53][826],u_xpb_out[54][826],u_xpb_out[55][826],u_xpb_out[56][826],u_xpb_out[57][826],u_xpb_out[58][826],u_xpb_out[59][826],u_xpb_out[60][826],u_xpb_out[61][826],u_xpb_out[62][826],u_xpb_out[63][826],u_xpb_out[64][826],u_xpb_out[65][826],u_xpb_out[66][826],u_xpb_out[67][826],u_xpb_out[68][826],u_xpb_out[69][826],u_xpb_out[70][826],u_xpb_out[71][826],u_xpb_out[72][826],u_xpb_out[73][826],u_xpb_out[74][826],u_xpb_out[75][826],u_xpb_out[76][826],u_xpb_out[77][826],u_xpb_out[78][826],u_xpb_out[79][826],u_xpb_out[80][826],u_xpb_out[81][826],u_xpb_out[82][826],u_xpb_out[83][826],u_xpb_out[84][826],u_xpb_out[85][826],u_xpb_out[86][826],u_xpb_out[87][826],u_xpb_out[88][826],u_xpb_out[89][826],u_xpb_out[90][826],u_xpb_out[91][826],u_xpb_out[92][826],u_xpb_out[93][826],u_xpb_out[94][826],u_xpb_out[95][826],u_xpb_out[96][826],u_xpb_out[97][826],u_xpb_out[98][826],u_xpb_out[99][826],u_xpb_out[100][826],u_xpb_out[101][826],u_xpb_out[102][826],u_xpb_out[103][826],u_xpb_out[104][826],u_xpb_out[105][826]};

assign col_out_827 = {u_xpb_out[0][827],u_xpb_out[1][827],u_xpb_out[2][827],u_xpb_out[3][827],u_xpb_out[4][827],u_xpb_out[5][827],u_xpb_out[6][827],u_xpb_out[7][827],u_xpb_out[8][827],u_xpb_out[9][827],u_xpb_out[10][827],u_xpb_out[11][827],u_xpb_out[12][827],u_xpb_out[13][827],u_xpb_out[14][827],u_xpb_out[15][827],u_xpb_out[16][827],u_xpb_out[17][827],u_xpb_out[18][827],u_xpb_out[19][827],u_xpb_out[20][827],u_xpb_out[21][827],u_xpb_out[22][827],u_xpb_out[23][827],u_xpb_out[24][827],u_xpb_out[25][827],u_xpb_out[26][827],u_xpb_out[27][827],u_xpb_out[28][827],u_xpb_out[29][827],u_xpb_out[30][827],u_xpb_out[31][827],u_xpb_out[32][827],u_xpb_out[33][827],u_xpb_out[34][827],u_xpb_out[35][827],u_xpb_out[36][827],u_xpb_out[37][827],u_xpb_out[38][827],u_xpb_out[39][827],u_xpb_out[40][827],u_xpb_out[41][827],u_xpb_out[42][827],u_xpb_out[43][827],u_xpb_out[44][827],u_xpb_out[45][827],u_xpb_out[46][827],u_xpb_out[47][827],u_xpb_out[48][827],u_xpb_out[49][827],u_xpb_out[50][827],u_xpb_out[51][827],u_xpb_out[52][827],u_xpb_out[53][827],u_xpb_out[54][827],u_xpb_out[55][827],u_xpb_out[56][827],u_xpb_out[57][827],u_xpb_out[58][827],u_xpb_out[59][827],u_xpb_out[60][827],u_xpb_out[61][827],u_xpb_out[62][827],u_xpb_out[63][827],u_xpb_out[64][827],u_xpb_out[65][827],u_xpb_out[66][827],u_xpb_out[67][827],u_xpb_out[68][827],u_xpb_out[69][827],u_xpb_out[70][827],u_xpb_out[71][827],u_xpb_out[72][827],u_xpb_out[73][827],u_xpb_out[74][827],u_xpb_out[75][827],u_xpb_out[76][827],u_xpb_out[77][827],u_xpb_out[78][827],u_xpb_out[79][827],u_xpb_out[80][827],u_xpb_out[81][827],u_xpb_out[82][827],u_xpb_out[83][827],u_xpb_out[84][827],u_xpb_out[85][827],u_xpb_out[86][827],u_xpb_out[87][827],u_xpb_out[88][827],u_xpb_out[89][827],u_xpb_out[90][827],u_xpb_out[91][827],u_xpb_out[92][827],u_xpb_out[93][827],u_xpb_out[94][827],u_xpb_out[95][827],u_xpb_out[96][827],u_xpb_out[97][827],u_xpb_out[98][827],u_xpb_out[99][827],u_xpb_out[100][827],u_xpb_out[101][827],u_xpb_out[102][827],u_xpb_out[103][827],u_xpb_out[104][827],u_xpb_out[105][827]};

assign col_out_828 = {u_xpb_out[0][828],u_xpb_out[1][828],u_xpb_out[2][828],u_xpb_out[3][828],u_xpb_out[4][828],u_xpb_out[5][828],u_xpb_out[6][828],u_xpb_out[7][828],u_xpb_out[8][828],u_xpb_out[9][828],u_xpb_out[10][828],u_xpb_out[11][828],u_xpb_out[12][828],u_xpb_out[13][828],u_xpb_out[14][828],u_xpb_out[15][828],u_xpb_out[16][828],u_xpb_out[17][828],u_xpb_out[18][828],u_xpb_out[19][828],u_xpb_out[20][828],u_xpb_out[21][828],u_xpb_out[22][828],u_xpb_out[23][828],u_xpb_out[24][828],u_xpb_out[25][828],u_xpb_out[26][828],u_xpb_out[27][828],u_xpb_out[28][828],u_xpb_out[29][828],u_xpb_out[30][828],u_xpb_out[31][828],u_xpb_out[32][828],u_xpb_out[33][828],u_xpb_out[34][828],u_xpb_out[35][828],u_xpb_out[36][828],u_xpb_out[37][828],u_xpb_out[38][828],u_xpb_out[39][828],u_xpb_out[40][828],u_xpb_out[41][828],u_xpb_out[42][828],u_xpb_out[43][828],u_xpb_out[44][828],u_xpb_out[45][828],u_xpb_out[46][828],u_xpb_out[47][828],u_xpb_out[48][828],u_xpb_out[49][828],u_xpb_out[50][828],u_xpb_out[51][828],u_xpb_out[52][828],u_xpb_out[53][828],u_xpb_out[54][828],u_xpb_out[55][828],u_xpb_out[56][828],u_xpb_out[57][828],u_xpb_out[58][828],u_xpb_out[59][828],u_xpb_out[60][828],u_xpb_out[61][828],u_xpb_out[62][828],u_xpb_out[63][828],u_xpb_out[64][828],u_xpb_out[65][828],u_xpb_out[66][828],u_xpb_out[67][828],u_xpb_out[68][828],u_xpb_out[69][828],u_xpb_out[70][828],u_xpb_out[71][828],u_xpb_out[72][828],u_xpb_out[73][828],u_xpb_out[74][828],u_xpb_out[75][828],u_xpb_out[76][828],u_xpb_out[77][828],u_xpb_out[78][828],u_xpb_out[79][828],u_xpb_out[80][828],u_xpb_out[81][828],u_xpb_out[82][828],u_xpb_out[83][828],u_xpb_out[84][828],u_xpb_out[85][828],u_xpb_out[86][828],u_xpb_out[87][828],u_xpb_out[88][828],u_xpb_out[89][828],u_xpb_out[90][828],u_xpb_out[91][828],u_xpb_out[92][828],u_xpb_out[93][828],u_xpb_out[94][828],u_xpb_out[95][828],u_xpb_out[96][828],u_xpb_out[97][828],u_xpb_out[98][828],u_xpb_out[99][828],u_xpb_out[100][828],u_xpb_out[101][828],u_xpb_out[102][828],u_xpb_out[103][828],u_xpb_out[104][828],u_xpb_out[105][828]};

assign col_out_829 = {u_xpb_out[0][829],u_xpb_out[1][829],u_xpb_out[2][829],u_xpb_out[3][829],u_xpb_out[4][829],u_xpb_out[5][829],u_xpb_out[6][829],u_xpb_out[7][829],u_xpb_out[8][829],u_xpb_out[9][829],u_xpb_out[10][829],u_xpb_out[11][829],u_xpb_out[12][829],u_xpb_out[13][829],u_xpb_out[14][829],u_xpb_out[15][829],u_xpb_out[16][829],u_xpb_out[17][829],u_xpb_out[18][829],u_xpb_out[19][829],u_xpb_out[20][829],u_xpb_out[21][829],u_xpb_out[22][829],u_xpb_out[23][829],u_xpb_out[24][829],u_xpb_out[25][829],u_xpb_out[26][829],u_xpb_out[27][829],u_xpb_out[28][829],u_xpb_out[29][829],u_xpb_out[30][829],u_xpb_out[31][829],u_xpb_out[32][829],u_xpb_out[33][829],u_xpb_out[34][829],u_xpb_out[35][829],u_xpb_out[36][829],u_xpb_out[37][829],u_xpb_out[38][829],u_xpb_out[39][829],u_xpb_out[40][829],u_xpb_out[41][829],u_xpb_out[42][829],u_xpb_out[43][829],u_xpb_out[44][829],u_xpb_out[45][829],u_xpb_out[46][829],u_xpb_out[47][829],u_xpb_out[48][829],u_xpb_out[49][829],u_xpb_out[50][829],u_xpb_out[51][829],u_xpb_out[52][829],u_xpb_out[53][829],u_xpb_out[54][829],u_xpb_out[55][829],u_xpb_out[56][829],u_xpb_out[57][829],u_xpb_out[58][829],u_xpb_out[59][829],u_xpb_out[60][829],u_xpb_out[61][829],u_xpb_out[62][829],u_xpb_out[63][829],u_xpb_out[64][829],u_xpb_out[65][829],u_xpb_out[66][829],u_xpb_out[67][829],u_xpb_out[68][829],u_xpb_out[69][829],u_xpb_out[70][829],u_xpb_out[71][829],u_xpb_out[72][829],u_xpb_out[73][829],u_xpb_out[74][829],u_xpb_out[75][829],u_xpb_out[76][829],u_xpb_out[77][829],u_xpb_out[78][829],u_xpb_out[79][829],u_xpb_out[80][829],u_xpb_out[81][829],u_xpb_out[82][829],u_xpb_out[83][829],u_xpb_out[84][829],u_xpb_out[85][829],u_xpb_out[86][829],u_xpb_out[87][829],u_xpb_out[88][829],u_xpb_out[89][829],u_xpb_out[90][829],u_xpb_out[91][829],u_xpb_out[92][829],u_xpb_out[93][829],u_xpb_out[94][829],u_xpb_out[95][829],u_xpb_out[96][829],u_xpb_out[97][829],u_xpb_out[98][829],u_xpb_out[99][829],u_xpb_out[100][829],u_xpb_out[101][829],u_xpb_out[102][829],u_xpb_out[103][829],u_xpb_out[104][829],u_xpb_out[105][829]};

assign col_out_830 = {u_xpb_out[0][830],u_xpb_out[1][830],u_xpb_out[2][830],u_xpb_out[3][830],u_xpb_out[4][830],u_xpb_out[5][830],u_xpb_out[6][830],u_xpb_out[7][830],u_xpb_out[8][830],u_xpb_out[9][830],u_xpb_out[10][830],u_xpb_out[11][830],u_xpb_out[12][830],u_xpb_out[13][830],u_xpb_out[14][830],u_xpb_out[15][830],u_xpb_out[16][830],u_xpb_out[17][830],u_xpb_out[18][830],u_xpb_out[19][830],u_xpb_out[20][830],u_xpb_out[21][830],u_xpb_out[22][830],u_xpb_out[23][830],u_xpb_out[24][830],u_xpb_out[25][830],u_xpb_out[26][830],u_xpb_out[27][830],u_xpb_out[28][830],u_xpb_out[29][830],u_xpb_out[30][830],u_xpb_out[31][830],u_xpb_out[32][830],u_xpb_out[33][830],u_xpb_out[34][830],u_xpb_out[35][830],u_xpb_out[36][830],u_xpb_out[37][830],u_xpb_out[38][830],u_xpb_out[39][830],u_xpb_out[40][830],u_xpb_out[41][830],u_xpb_out[42][830],u_xpb_out[43][830],u_xpb_out[44][830],u_xpb_out[45][830],u_xpb_out[46][830],u_xpb_out[47][830],u_xpb_out[48][830],u_xpb_out[49][830],u_xpb_out[50][830],u_xpb_out[51][830],u_xpb_out[52][830],u_xpb_out[53][830],u_xpb_out[54][830],u_xpb_out[55][830],u_xpb_out[56][830],u_xpb_out[57][830],u_xpb_out[58][830],u_xpb_out[59][830],u_xpb_out[60][830],u_xpb_out[61][830],u_xpb_out[62][830],u_xpb_out[63][830],u_xpb_out[64][830],u_xpb_out[65][830],u_xpb_out[66][830],u_xpb_out[67][830],u_xpb_out[68][830],u_xpb_out[69][830],u_xpb_out[70][830],u_xpb_out[71][830],u_xpb_out[72][830],u_xpb_out[73][830],u_xpb_out[74][830],u_xpb_out[75][830],u_xpb_out[76][830],u_xpb_out[77][830],u_xpb_out[78][830],u_xpb_out[79][830],u_xpb_out[80][830],u_xpb_out[81][830],u_xpb_out[82][830],u_xpb_out[83][830],u_xpb_out[84][830],u_xpb_out[85][830],u_xpb_out[86][830],u_xpb_out[87][830],u_xpb_out[88][830],u_xpb_out[89][830],u_xpb_out[90][830],u_xpb_out[91][830],u_xpb_out[92][830],u_xpb_out[93][830],u_xpb_out[94][830],u_xpb_out[95][830],u_xpb_out[96][830],u_xpb_out[97][830],u_xpb_out[98][830],u_xpb_out[99][830],u_xpb_out[100][830],u_xpb_out[101][830],u_xpb_out[102][830],u_xpb_out[103][830],u_xpb_out[104][830],u_xpb_out[105][830]};

assign col_out_831 = {u_xpb_out[0][831],u_xpb_out[1][831],u_xpb_out[2][831],u_xpb_out[3][831],u_xpb_out[4][831],u_xpb_out[5][831],u_xpb_out[6][831],u_xpb_out[7][831],u_xpb_out[8][831],u_xpb_out[9][831],u_xpb_out[10][831],u_xpb_out[11][831],u_xpb_out[12][831],u_xpb_out[13][831],u_xpb_out[14][831],u_xpb_out[15][831],u_xpb_out[16][831],u_xpb_out[17][831],u_xpb_out[18][831],u_xpb_out[19][831],u_xpb_out[20][831],u_xpb_out[21][831],u_xpb_out[22][831],u_xpb_out[23][831],u_xpb_out[24][831],u_xpb_out[25][831],u_xpb_out[26][831],u_xpb_out[27][831],u_xpb_out[28][831],u_xpb_out[29][831],u_xpb_out[30][831],u_xpb_out[31][831],u_xpb_out[32][831],u_xpb_out[33][831],u_xpb_out[34][831],u_xpb_out[35][831],u_xpb_out[36][831],u_xpb_out[37][831],u_xpb_out[38][831],u_xpb_out[39][831],u_xpb_out[40][831],u_xpb_out[41][831],u_xpb_out[42][831],u_xpb_out[43][831],u_xpb_out[44][831],u_xpb_out[45][831],u_xpb_out[46][831],u_xpb_out[47][831],u_xpb_out[48][831],u_xpb_out[49][831],u_xpb_out[50][831],u_xpb_out[51][831],u_xpb_out[52][831],u_xpb_out[53][831],u_xpb_out[54][831],u_xpb_out[55][831],u_xpb_out[56][831],u_xpb_out[57][831],u_xpb_out[58][831],u_xpb_out[59][831],u_xpb_out[60][831],u_xpb_out[61][831],u_xpb_out[62][831],u_xpb_out[63][831],u_xpb_out[64][831],u_xpb_out[65][831],u_xpb_out[66][831],u_xpb_out[67][831],u_xpb_out[68][831],u_xpb_out[69][831],u_xpb_out[70][831],u_xpb_out[71][831],u_xpb_out[72][831],u_xpb_out[73][831],u_xpb_out[74][831],u_xpb_out[75][831],u_xpb_out[76][831],u_xpb_out[77][831],u_xpb_out[78][831],u_xpb_out[79][831],u_xpb_out[80][831],u_xpb_out[81][831],u_xpb_out[82][831],u_xpb_out[83][831],u_xpb_out[84][831],u_xpb_out[85][831],u_xpb_out[86][831],u_xpb_out[87][831],u_xpb_out[88][831],u_xpb_out[89][831],u_xpb_out[90][831],u_xpb_out[91][831],u_xpb_out[92][831],u_xpb_out[93][831],u_xpb_out[94][831],u_xpb_out[95][831],u_xpb_out[96][831],u_xpb_out[97][831],u_xpb_out[98][831],u_xpb_out[99][831],u_xpb_out[100][831],u_xpb_out[101][831],u_xpb_out[102][831],u_xpb_out[103][831],u_xpb_out[104][831],u_xpb_out[105][831]};

assign col_out_832 = {u_xpb_out[0][832],u_xpb_out[1][832],u_xpb_out[2][832],u_xpb_out[3][832],u_xpb_out[4][832],u_xpb_out[5][832],u_xpb_out[6][832],u_xpb_out[7][832],u_xpb_out[8][832],u_xpb_out[9][832],u_xpb_out[10][832],u_xpb_out[11][832],u_xpb_out[12][832],u_xpb_out[13][832],u_xpb_out[14][832],u_xpb_out[15][832],u_xpb_out[16][832],u_xpb_out[17][832],u_xpb_out[18][832],u_xpb_out[19][832],u_xpb_out[20][832],u_xpb_out[21][832],u_xpb_out[22][832],u_xpb_out[23][832],u_xpb_out[24][832],u_xpb_out[25][832],u_xpb_out[26][832],u_xpb_out[27][832],u_xpb_out[28][832],u_xpb_out[29][832],u_xpb_out[30][832],u_xpb_out[31][832],u_xpb_out[32][832],u_xpb_out[33][832],u_xpb_out[34][832],u_xpb_out[35][832],u_xpb_out[36][832],u_xpb_out[37][832],u_xpb_out[38][832],u_xpb_out[39][832],u_xpb_out[40][832],u_xpb_out[41][832],u_xpb_out[42][832],u_xpb_out[43][832],u_xpb_out[44][832],u_xpb_out[45][832],u_xpb_out[46][832],u_xpb_out[47][832],u_xpb_out[48][832],u_xpb_out[49][832],u_xpb_out[50][832],u_xpb_out[51][832],u_xpb_out[52][832],u_xpb_out[53][832],u_xpb_out[54][832],u_xpb_out[55][832],u_xpb_out[56][832],u_xpb_out[57][832],u_xpb_out[58][832],u_xpb_out[59][832],u_xpb_out[60][832],u_xpb_out[61][832],u_xpb_out[62][832],u_xpb_out[63][832],u_xpb_out[64][832],u_xpb_out[65][832],u_xpb_out[66][832],u_xpb_out[67][832],u_xpb_out[68][832],u_xpb_out[69][832],u_xpb_out[70][832],u_xpb_out[71][832],u_xpb_out[72][832],u_xpb_out[73][832],u_xpb_out[74][832],u_xpb_out[75][832],u_xpb_out[76][832],u_xpb_out[77][832],u_xpb_out[78][832],u_xpb_out[79][832],u_xpb_out[80][832],u_xpb_out[81][832],u_xpb_out[82][832],u_xpb_out[83][832],u_xpb_out[84][832],u_xpb_out[85][832],u_xpb_out[86][832],u_xpb_out[87][832],u_xpb_out[88][832],u_xpb_out[89][832],u_xpb_out[90][832],u_xpb_out[91][832],u_xpb_out[92][832],u_xpb_out[93][832],u_xpb_out[94][832],u_xpb_out[95][832],u_xpb_out[96][832],u_xpb_out[97][832],u_xpb_out[98][832],u_xpb_out[99][832],u_xpb_out[100][832],u_xpb_out[101][832],u_xpb_out[102][832],u_xpb_out[103][832],u_xpb_out[104][832],u_xpb_out[105][832]};

assign col_out_833 = {u_xpb_out[0][833],u_xpb_out[1][833],u_xpb_out[2][833],u_xpb_out[3][833],u_xpb_out[4][833],u_xpb_out[5][833],u_xpb_out[6][833],u_xpb_out[7][833],u_xpb_out[8][833],u_xpb_out[9][833],u_xpb_out[10][833],u_xpb_out[11][833],u_xpb_out[12][833],u_xpb_out[13][833],u_xpb_out[14][833],u_xpb_out[15][833],u_xpb_out[16][833],u_xpb_out[17][833],u_xpb_out[18][833],u_xpb_out[19][833],u_xpb_out[20][833],u_xpb_out[21][833],u_xpb_out[22][833],u_xpb_out[23][833],u_xpb_out[24][833],u_xpb_out[25][833],u_xpb_out[26][833],u_xpb_out[27][833],u_xpb_out[28][833],u_xpb_out[29][833],u_xpb_out[30][833],u_xpb_out[31][833],u_xpb_out[32][833],u_xpb_out[33][833],u_xpb_out[34][833],u_xpb_out[35][833],u_xpb_out[36][833],u_xpb_out[37][833],u_xpb_out[38][833],u_xpb_out[39][833],u_xpb_out[40][833],u_xpb_out[41][833],u_xpb_out[42][833],u_xpb_out[43][833],u_xpb_out[44][833],u_xpb_out[45][833],u_xpb_out[46][833],u_xpb_out[47][833],u_xpb_out[48][833],u_xpb_out[49][833],u_xpb_out[50][833],u_xpb_out[51][833],u_xpb_out[52][833],u_xpb_out[53][833],u_xpb_out[54][833],u_xpb_out[55][833],u_xpb_out[56][833],u_xpb_out[57][833],u_xpb_out[58][833],u_xpb_out[59][833],u_xpb_out[60][833],u_xpb_out[61][833],u_xpb_out[62][833],u_xpb_out[63][833],u_xpb_out[64][833],u_xpb_out[65][833],u_xpb_out[66][833],u_xpb_out[67][833],u_xpb_out[68][833],u_xpb_out[69][833],u_xpb_out[70][833],u_xpb_out[71][833],u_xpb_out[72][833],u_xpb_out[73][833],u_xpb_out[74][833],u_xpb_out[75][833],u_xpb_out[76][833],u_xpb_out[77][833],u_xpb_out[78][833],u_xpb_out[79][833],u_xpb_out[80][833],u_xpb_out[81][833],u_xpb_out[82][833],u_xpb_out[83][833],u_xpb_out[84][833],u_xpb_out[85][833],u_xpb_out[86][833],u_xpb_out[87][833],u_xpb_out[88][833],u_xpb_out[89][833],u_xpb_out[90][833],u_xpb_out[91][833],u_xpb_out[92][833],u_xpb_out[93][833],u_xpb_out[94][833],u_xpb_out[95][833],u_xpb_out[96][833],u_xpb_out[97][833],u_xpb_out[98][833],u_xpb_out[99][833],u_xpb_out[100][833],u_xpb_out[101][833],u_xpb_out[102][833],u_xpb_out[103][833],u_xpb_out[104][833],u_xpb_out[105][833]};

assign col_out_834 = {u_xpb_out[0][834],u_xpb_out[1][834],u_xpb_out[2][834],u_xpb_out[3][834],u_xpb_out[4][834],u_xpb_out[5][834],u_xpb_out[6][834],u_xpb_out[7][834],u_xpb_out[8][834],u_xpb_out[9][834],u_xpb_out[10][834],u_xpb_out[11][834],u_xpb_out[12][834],u_xpb_out[13][834],u_xpb_out[14][834],u_xpb_out[15][834],u_xpb_out[16][834],u_xpb_out[17][834],u_xpb_out[18][834],u_xpb_out[19][834],u_xpb_out[20][834],u_xpb_out[21][834],u_xpb_out[22][834],u_xpb_out[23][834],u_xpb_out[24][834],u_xpb_out[25][834],u_xpb_out[26][834],u_xpb_out[27][834],u_xpb_out[28][834],u_xpb_out[29][834],u_xpb_out[30][834],u_xpb_out[31][834],u_xpb_out[32][834],u_xpb_out[33][834],u_xpb_out[34][834],u_xpb_out[35][834],u_xpb_out[36][834],u_xpb_out[37][834],u_xpb_out[38][834],u_xpb_out[39][834],u_xpb_out[40][834],u_xpb_out[41][834],u_xpb_out[42][834],u_xpb_out[43][834],u_xpb_out[44][834],u_xpb_out[45][834],u_xpb_out[46][834],u_xpb_out[47][834],u_xpb_out[48][834],u_xpb_out[49][834],u_xpb_out[50][834],u_xpb_out[51][834],u_xpb_out[52][834],u_xpb_out[53][834],u_xpb_out[54][834],u_xpb_out[55][834],u_xpb_out[56][834],u_xpb_out[57][834],u_xpb_out[58][834],u_xpb_out[59][834],u_xpb_out[60][834],u_xpb_out[61][834],u_xpb_out[62][834],u_xpb_out[63][834],u_xpb_out[64][834],u_xpb_out[65][834],u_xpb_out[66][834],u_xpb_out[67][834],u_xpb_out[68][834],u_xpb_out[69][834],u_xpb_out[70][834],u_xpb_out[71][834],u_xpb_out[72][834],u_xpb_out[73][834],u_xpb_out[74][834],u_xpb_out[75][834],u_xpb_out[76][834],u_xpb_out[77][834],u_xpb_out[78][834],u_xpb_out[79][834],u_xpb_out[80][834],u_xpb_out[81][834],u_xpb_out[82][834],u_xpb_out[83][834],u_xpb_out[84][834],u_xpb_out[85][834],u_xpb_out[86][834],u_xpb_out[87][834],u_xpb_out[88][834],u_xpb_out[89][834],u_xpb_out[90][834],u_xpb_out[91][834],u_xpb_out[92][834],u_xpb_out[93][834],u_xpb_out[94][834],u_xpb_out[95][834],u_xpb_out[96][834],u_xpb_out[97][834],u_xpb_out[98][834],u_xpb_out[99][834],u_xpb_out[100][834],u_xpb_out[101][834],u_xpb_out[102][834],u_xpb_out[103][834],u_xpb_out[104][834],u_xpb_out[105][834]};

assign col_out_835 = {u_xpb_out[0][835],u_xpb_out[1][835],u_xpb_out[2][835],u_xpb_out[3][835],u_xpb_out[4][835],u_xpb_out[5][835],u_xpb_out[6][835],u_xpb_out[7][835],u_xpb_out[8][835],u_xpb_out[9][835],u_xpb_out[10][835],u_xpb_out[11][835],u_xpb_out[12][835],u_xpb_out[13][835],u_xpb_out[14][835],u_xpb_out[15][835],u_xpb_out[16][835],u_xpb_out[17][835],u_xpb_out[18][835],u_xpb_out[19][835],u_xpb_out[20][835],u_xpb_out[21][835],u_xpb_out[22][835],u_xpb_out[23][835],u_xpb_out[24][835],u_xpb_out[25][835],u_xpb_out[26][835],u_xpb_out[27][835],u_xpb_out[28][835],u_xpb_out[29][835],u_xpb_out[30][835],u_xpb_out[31][835],u_xpb_out[32][835],u_xpb_out[33][835],u_xpb_out[34][835],u_xpb_out[35][835],u_xpb_out[36][835],u_xpb_out[37][835],u_xpb_out[38][835],u_xpb_out[39][835],u_xpb_out[40][835],u_xpb_out[41][835],u_xpb_out[42][835],u_xpb_out[43][835],u_xpb_out[44][835],u_xpb_out[45][835],u_xpb_out[46][835],u_xpb_out[47][835],u_xpb_out[48][835],u_xpb_out[49][835],u_xpb_out[50][835],u_xpb_out[51][835],u_xpb_out[52][835],u_xpb_out[53][835],u_xpb_out[54][835],u_xpb_out[55][835],u_xpb_out[56][835],u_xpb_out[57][835],u_xpb_out[58][835],u_xpb_out[59][835],u_xpb_out[60][835],u_xpb_out[61][835],u_xpb_out[62][835],u_xpb_out[63][835],u_xpb_out[64][835],u_xpb_out[65][835],u_xpb_out[66][835],u_xpb_out[67][835],u_xpb_out[68][835],u_xpb_out[69][835],u_xpb_out[70][835],u_xpb_out[71][835],u_xpb_out[72][835],u_xpb_out[73][835],u_xpb_out[74][835],u_xpb_out[75][835],u_xpb_out[76][835],u_xpb_out[77][835],u_xpb_out[78][835],u_xpb_out[79][835],u_xpb_out[80][835],u_xpb_out[81][835],u_xpb_out[82][835],u_xpb_out[83][835],u_xpb_out[84][835],u_xpb_out[85][835],u_xpb_out[86][835],u_xpb_out[87][835],u_xpb_out[88][835],u_xpb_out[89][835],u_xpb_out[90][835],u_xpb_out[91][835],u_xpb_out[92][835],u_xpb_out[93][835],u_xpb_out[94][835],u_xpb_out[95][835],u_xpb_out[96][835],u_xpb_out[97][835],u_xpb_out[98][835],u_xpb_out[99][835],u_xpb_out[100][835],u_xpb_out[101][835],u_xpb_out[102][835],u_xpb_out[103][835],u_xpb_out[104][835],u_xpb_out[105][835]};

assign col_out_836 = {u_xpb_out[0][836],u_xpb_out[1][836],u_xpb_out[2][836],u_xpb_out[3][836],u_xpb_out[4][836],u_xpb_out[5][836],u_xpb_out[6][836],u_xpb_out[7][836],u_xpb_out[8][836],u_xpb_out[9][836],u_xpb_out[10][836],u_xpb_out[11][836],u_xpb_out[12][836],u_xpb_out[13][836],u_xpb_out[14][836],u_xpb_out[15][836],u_xpb_out[16][836],u_xpb_out[17][836],u_xpb_out[18][836],u_xpb_out[19][836],u_xpb_out[20][836],u_xpb_out[21][836],u_xpb_out[22][836],u_xpb_out[23][836],u_xpb_out[24][836],u_xpb_out[25][836],u_xpb_out[26][836],u_xpb_out[27][836],u_xpb_out[28][836],u_xpb_out[29][836],u_xpb_out[30][836],u_xpb_out[31][836],u_xpb_out[32][836],u_xpb_out[33][836],u_xpb_out[34][836],u_xpb_out[35][836],u_xpb_out[36][836],u_xpb_out[37][836],u_xpb_out[38][836],u_xpb_out[39][836],u_xpb_out[40][836],u_xpb_out[41][836],u_xpb_out[42][836],u_xpb_out[43][836],u_xpb_out[44][836],u_xpb_out[45][836],u_xpb_out[46][836],u_xpb_out[47][836],u_xpb_out[48][836],u_xpb_out[49][836],u_xpb_out[50][836],u_xpb_out[51][836],u_xpb_out[52][836],u_xpb_out[53][836],u_xpb_out[54][836],u_xpb_out[55][836],u_xpb_out[56][836],u_xpb_out[57][836],u_xpb_out[58][836],u_xpb_out[59][836],u_xpb_out[60][836],u_xpb_out[61][836],u_xpb_out[62][836],u_xpb_out[63][836],u_xpb_out[64][836],u_xpb_out[65][836],u_xpb_out[66][836],u_xpb_out[67][836],u_xpb_out[68][836],u_xpb_out[69][836],u_xpb_out[70][836],u_xpb_out[71][836],u_xpb_out[72][836],u_xpb_out[73][836],u_xpb_out[74][836],u_xpb_out[75][836],u_xpb_out[76][836],u_xpb_out[77][836],u_xpb_out[78][836],u_xpb_out[79][836],u_xpb_out[80][836],u_xpb_out[81][836],u_xpb_out[82][836],u_xpb_out[83][836],u_xpb_out[84][836],u_xpb_out[85][836],u_xpb_out[86][836],u_xpb_out[87][836],u_xpb_out[88][836],u_xpb_out[89][836],u_xpb_out[90][836],u_xpb_out[91][836],u_xpb_out[92][836],u_xpb_out[93][836],u_xpb_out[94][836],u_xpb_out[95][836],u_xpb_out[96][836],u_xpb_out[97][836],u_xpb_out[98][836],u_xpb_out[99][836],u_xpb_out[100][836],u_xpb_out[101][836],u_xpb_out[102][836],u_xpb_out[103][836],u_xpb_out[104][836],u_xpb_out[105][836]};

assign col_out_837 = {u_xpb_out[0][837],u_xpb_out[1][837],u_xpb_out[2][837],u_xpb_out[3][837],u_xpb_out[4][837],u_xpb_out[5][837],u_xpb_out[6][837],u_xpb_out[7][837],u_xpb_out[8][837],u_xpb_out[9][837],u_xpb_out[10][837],u_xpb_out[11][837],u_xpb_out[12][837],u_xpb_out[13][837],u_xpb_out[14][837],u_xpb_out[15][837],u_xpb_out[16][837],u_xpb_out[17][837],u_xpb_out[18][837],u_xpb_out[19][837],u_xpb_out[20][837],u_xpb_out[21][837],u_xpb_out[22][837],u_xpb_out[23][837],u_xpb_out[24][837],u_xpb_out[25][837],u_xpb_out[26][837],u_xpb_out[27][837],u_xpb_out[28][837],u_xpb_out[29][837],u_xpb_out[30][837],u_xpb_out[31][837],u_xpb_out[32][837],u_xpb_out[33][837],u_xpb_out[34][837],u_xpb_out[35][837],u_xpb_out[36][837],u_xpb_out[37][837],u_xpb_out[38][837],u_xpb_out[39][837],u_xpb_out[40][837],u_xpb_out[41][837],u_xpb_out[42][837],u_xpb_out[43][837],u_xpb_out[44][837],u_xpb_out[45][837],u_xpb_out[46][837],u_xpb_out[47][837],u_xpb_out[48][837],u_xpb_out[49][837],u_xpb_out[50][837],u_xpb_out[51][837],u_xpb_out[52][837],u_xpb_out[53][837],u_xpb_out[54][837],u_xpb_out[55][837],u_xpb_out[56][837],u_xpb_out[57][837],u_xpb_out[58][837],u_xpb_out[59][837],u_xpb_out[60][837],u_xpb_out[61][837],u_xpb_out[62][837],u_xpb_out[63][837],u_xpb_out[64][837],u_xpb_out[65][837],u_xpb_out[66][837],u_xpb_out[67][837],u_xpb_out[68][837],u_xpb_out[69][837],u_xpb_out[70][837],u_xpb_out[71][837],u_xpb_out[72][837],u_xpb_out[73][837],u_xpb_out[74][837],u_xpb_out[75][837],u_xpb_out[76][837],u_xpb_out[77][837],u_xpb_out[78][837],u_xpb_out[79][837],u_xpb_out[80][837],u_xpb_out[81][837],u_xpb_out[82][837],u_xpb_out[83][837],u_xpb_out[84][837],u_xpb_out[85][837],u_xpb_out[86][837],u_xpb_out[87][837],u_xpb_out[88][837],u_xpb_out[89][837],u_xpb_out[90][837],u_xpb_out[91][837],u_xpb_out[92][837],u_xpb_out[93][837],u_xpb_out[94][837],u_xpb_out[95][837],u_xpb_out[96][837],u_xpb_out[97][837],u_xpb_out[98][837],u_xpb_out[99][837],u_xpb_out[100][837],u_xpb_out[101][837],u_xpb_out[102][837],u_xpb_out[103][837],u_xpb_out[104][837],u_xpb_out[105][837]};

assign col_out_838 = {u_xpb_out[0][838],u_xpb_out[1][838],u_xpb_out[2][838],u_xpb_out[3][838],u_xpb_out[4][838],u_xpb_out[5][838],u_xpb_out[6][838],u_xpb_out[7][838],u_xpb_out[8][838],u_xpb_out[9][838],u_xpb_out[10][838],u_xpb_out[11][838],u_xpb_out[12][838],u_xpb_out[13][838],u_xpb_out[14][838],u_xpb_out[15][838],u_xpb_out[16][838],u_xpb_out[17][838],u_xpb_out[18][838],u_xpb_out[19][838],u_xpb_out[20][838],u_xpb_out[21][838],u_xpb_out[22][838],u_xpb_out[23][838],u_xpb_out[24][838],u_xpb_out[25][838],u_xpb_out[26][838],u_xpb_out[27][838],u_xpb_out[28][838],u_xpb_out[29][838],u_xpb_out[30][838],u_xpb_out[31][838],u_xpb_out[32][838],u_xpb_out[33][838],u_xpb_out[34][838],u_xpb_out[35][838],u_xpb_out[36][838],u_xpb_out[37][838],u_xpb_out[38][838],u_xpb_out[39][838],u_xpb_out[40][838],u_xpb_out[41][838],u_xpb_out[42][838],u_xpb_out[43][838],u_xpb_out[44][838],u_xpb_out[45][838],u_xpb_out[46][838],u_xpb_out[47][838],u_xpb_out[48][838],u_xpb_out[49][838],u_xpb_out[50][838],u_xpb_out[51][838],u_xpb_out[52][838],u_xpb_out[53][838],u_xpb_out[54][838],u_xpb_out[55][838],u_xpb_out[56][838],u_xpb_out[57][838],u_xpb_out[58][838],u_xpb_out[59][838],u_xpb_out[60][838],u_xpb_out[61][838],u_xpb_out[62][838],u_xpb_out[63][838],u_xpb_out[64][838],u_xpb_out[65][838],u_xpb_out[66][838],u_xpb_out[67][838],u_xpb_out[68][838],u_xpb_out[69][838],u_xpb_out[70][838],u_xpb_out[71][838],u_xpb_out[72][838],u_xpb_out[73][838],u_xpb_out[74][838],u_xpb_out[75][838],u_xpb_out[76][838],u_xpb_out[77][838],u_xpb_out[78][838],u_xpb_out[79][838],u_xpb_out[80][838],u_xpb_out[81][838],u_xpb_out[82][838],u_xpb_out[83][838],u_xpb_out[84][838],u_xpb_out[85][838],u_xpb_out[86][838],u_xpb_out[87][838],u_xpb_out[88][838],u_xpb_out[89][838],u_xpb_out[90][838],u_xpb_out[91][838],u_xpb_out[92][838],u_xpb_out[93][838],u_xpb_out[94][838],u_xpb_out[95][838],u_xpb_out[96][838],u_xpb_out[97][838],u_xpb_out[98][838],u_xpb_out[99][838],u_xpb_out[100][838],u_xpb_out[101][838],u_xpb_out[102][838],u_xpb_out[103][838],u_xpb_out[104][838],u_xpb_out[105][838]};

assign col_out_839 = {u_xpb_out[0][839],u_xpb_out[1][839],u_xpb_out[2][839],u_xpb_out[3][839],u_xpb_out[4][839],u_xpb_out[5][839],u_xpb_out[6][839],u_xpb_out[7][839],u_xpb_out[8][839],u_xpb_out[9][839],u_xpb_out[10][839],u_xpb_out[11][839],u_xpb_out[12][839],u_xpb_out[13][839],u_xpb_out[14][839],u_xpb_out[15][839],u_xpb_out[16][839],u_xpb_out[17][839],u_xpb_out[18][839],u_xpb_out[19][839],u_xpb_out[20][839],u_xpb_out[21][839],u_xpb_out[22][839],u_xpb_out[23][839],u_xpb_out[24][839],u_xpb_out[25][839],u_xpb_out[26][839],u_xpb_out[27][839],u_xpb_out[28][839],u_xpb_out[29][839],u_xpb_out[30][839],u_xpb_out[31][839],u_xpb_out[32][839],u_xpb_out[33][839],u_xpb_out[34][839],u_xpb_out[35][839],u_xpb_out[36][839],u_xpb_out[37][839],u_xpb_out[38][839],u_xpb_out[39][839],u_xpb_out[40][839],u_xpb_out[41][839],u_xpb_out[42][839],u_xpb_out[43][839],u_xpb_out[44][839],u_xpb_out[45][839],u_xpb_out[46][839],u_xpb_out[47][839],u_xpb_out[48][839],u_xpb_out[49][839],u_xpb_out[50][839],u_xpb_out[51][839],u_xpb_out[52][839],u_xpb_out[53][839],u_xpb_out[54][839],u_xpb_out[55][839],u_xpb_out[56][839],u_xpb_out[57][839],u_xpb_out[58][839],u_xpb_out[59][839],u_xpb_out[60][839],u_xpb_out[61][839],u_xpb_out[62][839],u_xpb_out[63][839],u_xpb_out[64][839],u_xpb_out[65][839],u_xpb_out[66][839],u_xpb_out[67][839],u_xpb_out[68][839],u_xpb_out[69][839],u_xpb_out[70][839],u_xpb_out[71][839],u_xpb_out[72][839],u_xpb_out[73][839],u_xpb_out[74][839],u_xpb_out[75][839],u_xpb_out[76][839],u_xpb_out[77][839],u_xpb_out[78][839],u_xpb_out[79][839],u_xpb_out[80][839],u_xpb_out[81][839],u_xpb_out[82][839],u_xpb_out[83][839],u_xpb_out[84][839],u_xpb_out[85][839],u_xpb_out[86][839],u_xpb_out[87][839],u_xpb_out[88][839],u_xpb_out[89][839],u_xpb_out[90][839],u_xpb_out[91][839],u_xpb_out[92][839],u_xpb_out[93][839],u_xpb_out[94][839],u_xpb_out[95][839],u_xpb_out[96][839],u_xpb_out[97][839],u_xpb_out[98][839],u_xpb_out[99][839],u_xpb_out[100][839],u_xpb_out[101][839],u_xpb_out[102][839],u_xpb_out[103][839],u_xpb_out[104][839],u_xpb_out[105][839]};

assign col_out_840 = {u_xpb_out[0][840],u_xpb_out[1][840],u_xpb_out[2][840],u_xpb_out[3][840],u_xpb_out[4][840],u_xpb_out[5][840],u_xpb_out[6][840],u_xpb_out[7][840],u_xpb_out[8][840],u_xpb_out[9][840],u_xpb_out[10][840],u_xpb_out[11][840],u_xpb_out[12][840],u_xpb_out[13][840],u_xpb_out[14][840],u_xpb_out[15][840],u_xpb_out[16][840],u_xpb_out[17][840],u_xpb_out[18][840],u_xpb_out[19][840],u_xpb_out[20][840],u_xpb_out[21][840],u_xpb_out[22][840],u_xpb_out[23][840],u_xpb_out[24][840],u_xpb_out[25][840],u_xpb_out[26][840],u_xpb_out[27][840],u_xpb_out[28][840],u_xpb_out[29][840],u_xpb_out[30][840],u_xpb_out[31][840],u_xpb_out[32][840],u_xpb_out[33][840],u_xpb_out[34][840],u_xpb_out[35][840],u_xpb_out[36][840],u_xpb_out[37][840],u_xpb_out[38][840],u_xpb_out[39][840],u_xpb_out[40][840],u_xpb_out[41][840],u_xpb_out[42][840],u_xpb_out[43][840],u_xpb_out[44][840],u_xpb_out[45][840],u_xpb_out[46][840],u_xpb_out[47][840],u_xpb_out[48][840],u_xpb_out[49][840],u_xpb_out[50][840],u_xpb_out[51][840],u_xpb_out[52][840],u_xpb_out[53][840],u_xpb_out[54][840],u_xpb_out[55][840],u_xpb_out[56][840],u_xpb_out[57][840],u_xpb_out[58][840],u_xpb_out[59][840],u_xpb_out[60][840],u_xpb_out[61][840],u_xpb_out[62][840],u_xpb_out[63][840],u_xpb_out[64][840],u_xpb_out[65][840],u_xpb_out[66][840],u_xpb_out[67][840],u_xpb_out[68][840],u_xpb_out[69][840],u_xpb_out[70][840],u_xpb_out[71][840],u_xpb_out[72][840],u_xpb_out[73][840],u_xpb_out[74][840],u_xpb_out[75][840],u_xpb_out[76][840],u_xpb_out[77][840],u_xpb_out[78][840],u_xpb_out[79][840],u_xpb_out[80][840],u_xpb_out[81][840],u_xpb_out[82][840],u_xpb_out[83][840],u_xpb_out[84][840],u_xpb_out[85][840],u_xpb_out[86][840],u_xpb_out[87][840],u_xpb_out[88][840],u_xpb_out[89][840],u_xpb_out[90][840],u_xpb_out[91][840],u_xpb_out[92][840],u_xpb_out[93][840],u_xpb_out[94][840],u_xpb_out[95][840],u_xpb_out[96][840],u_xpb_out[97][840],u_xpb_out[98][840],u_xpb_out[99][840],u_xpb_out[100][840],u_xpb_out[101][840],u_xpb_out[102][840],u_xpb_out[103][840],u_xpb_out[104][840],u_xpb_out[105][840]};

assign col_out_841 = {u_xpb_out[0][841],u_xpb_out[1][841],u_xpb_out[2][841],u_xpb_out[3][841],u_xpb_out[4][841],u_xpb_out[5][841],u_xpb_out[6][841],u_xpb_out[7][841],u_xpb_out[8][841],u_xpb_out[9][841],u_xpb_out[10][841],u_xpb_out[11][841],u_xpb_out[12][841],u_xpb_out[13][841],u_xpb_out[14][841],u_xpb_out[15][841],u_xpb_out[16][841],u_xpb_out[17][841],u_xpb_out[18][841],u_xpb_out[19][841],u_xpb_out[20][841],u_xpb_out[21][841],u_xpb_out[22][841],u_xpb_out[23][841],u_xpb_out[24][841],u_xpb_out[25][841],u_xpb_out[26][841],u_xpb_out[27][841],u_xpb_out[28][841],u_xpb_out[29][841],u_xpb_out[30][841],u_xpb_out[31][841],u_xpb_out[32][841],u_xpb_out[33][841],u_xpb_out[34][841],u_xpb_out[35][841],u_xpb_out[36][841],u_xpb_out[37][841],u_xpb_out[38][841],u_xpb_out[39][841],u_xpb_out[40][841],u_xpb_out[41][841],u_xpb_out[42][841],u_xpb_out[43][841],u_xpb_out[44][841],u_xpb_out[45][841],u_xpb_out[46][841],u_xpb_out[47][841],u_xpb_out[48][841],u_xpb_out[49][841],u_xpb_out[50][841],u_xpb_out[51][841],u_xpb_out[52][841],u_xpb_out[53][841],u_xpb_out[54][841],u_xpb_out[55][841],u_xpb_out[56][841],u_xpb_out[57][841],u_xpb_out[58][841],u_xpb_out[59][841],u_xpb_out[60][841],u_xpb_out[61][841],u_xpb_out[62][841],u_xpb_out[63][841],u_xpb_out[64][841],u_xpb_out[65][841],u_xpb_out[66][841],u_xpb_out[67][841],u_xpb_out[68][841],u_xpb_out[69][841],u_xpb_out[70][841],u_xpb_out[71][841],u_xpb_out[72][841],u_xpb_out[73][841],u_xpb_out[74][841],u_xpb_out[75][841],u_xpb_out[76][841],u_xpb_out[77][841],u_xpb_out[78][841],u_xpb_out[79][841],u_xpb_out[80][841],u_xpb_out[81][841],u_xpb_out[82][841],u_xpb_out[83][841],u_xpb_out[84][841],u_xpb_out[85][841],u_xpb_out[86][841],u_xpb_out[87][841],u_xpb_out[88][841],u_xpb_out[89][841],u_xpb_out[90][841],u_xpb_out[91][841],u_xpb_out[92][841],u_xpb_out[93][841],u_xpb_out[94][841],u_xpb_out[95][841],u_xpb_out[96][841],u_xpb_out[97][841],u_xpb_out[98][841],u_xpb_out[99][841],u_xpb_out[100][841],u_xpb_out[101][841],u_xpb_out[102][841],u_xpb_out[103][841],u_xpb_out[104][841],u_xpb_out[105][841]};

assign col_out_842 = {u_xpb_out[0][842],u_xpb_out[1][842],u_xpb_out[2][842],u_xpb_out[3][842],u_xpb_out[4][842],u_xpb_out[5][842],u_xpb_out[6][842],u_xpb_out[7][842],u_xpb_out[8][842],u_xpb_out[9][842],u_xpb_out[10][842],u_xpb_out[11][842],u_xpb_out[12][842],u_xpb_out[13][842],u_xpb_out[14][842],u_xpb_out[15][842],u_xpb_out[16][842],u_xpb_out[17][842],u_xpb_out[18][842],u_xpb_out[19][842],u_xpb_out[20][842],u_xpb_out[21][842],u_xpb_out[22][842],u_xpb_out[23][842],u_xpb_out[24][842],u_xpb_out[25][842],u_xpb_out[26][842],u_xpb_out[27][842],u_xpb_out[28][842],u_xpb_out[29][842],u_xpb_out[30][842],u_xpb_out[31][842],u_xpb_out[32][842],u_xpb_out[33][842],u_xpb_out[34][842],u_xpb_out[35][842],u_xpb_out[36][842],u_xpb_out[37][842],u_xpb_out[38][842],u_xpb_out[39][842],u_xpb_out[40][842],u_xpb_out[41][842],u_xpb_out[42][842],u_xpb_out[43][842],u_xpb_out[44][842],u_xpb_out[45][842],u_xpb_out[46][842],u_xpb_out[47][842],u_xpb_out[48][842],u_xpb_out[49][842],u_xpb_out[50][842],u_xpb_out[51][842],u_xpb_out[52][842],u_xpb_out[53][842],u_xpb_out[54][842],u_xpb_out[55][842],u_xpb_out[56][842],u_xpb_out[57][842],u_xpb_out[58][842],u_xpb_out[59][842],u_xpb_out[60][842],u_xpb_out[61][842],u_xpb_out[62][842],u_xpb_out[63][842],u_xpb_out[64][842],u_xpb_out[65][842],u_xpb_out[66][842],u_xpb_out[67][842],u_xpb_out[68][842],u_xpb_out[69][842],u_xpb_out[70][842],u_xpb_out[71][842],u_xpb_out[72][842],u_xpb_out[73][842],u_xpb_out[74][842],u_xpb_out[75][842],u_xpb_out[76][842],u_xpb_out[77][842],u_xpb_out[78][842],u_xpb_out[79][842],u_xpb_out[80][842],u_xpb_out[81][842],u_xpb_out[82][842],u_xpb_out[83][842],u_xpb_out[84][842],u_xpb_out[85][842],u_xpb_out[86][842],u_xpb_out[87][842],u_xpb_out[88][842],u_xpb_out[89][842],u_xpb_out[90][842],u_xpb_out[91][842],u_xpb_out[92][842],u_xpb_out[93][842],u_xpb_out[94][842],u_xpb_out[95][842],u_xpb_out[96][842],u_xpb_out[97][842],u_xpb_out[98][842],u_xpb_out[99][842],u_xpb_out[100][842],u_xpb_out[101][842],u_xpb_out[102][842],u_xpb_out[103][842],u_xpb_out[104][842],u_xpb_out[105][842]};

assign col_out_843 = {u_xpb_out[0][843],u_xpb_out[1][843],u_xpb_out[2][843],u_xpb_out[3][843],u_xpb_out[4][843],u_xpb_out[5][843],u_xpb_out[6][843],u_xpb_out[7][843],u_xpb_out[8][843],u_xpb_out[9][843],u_xpb_out[10][843],u_xpb_out[11][843],u_xpb_out[12][843],u_xpb_out[13][843],u_xpb_out[14][843],u_xpb_out[15][843],u_xpb_out[16][843],u_xpb_out[17][843],u_xpb_out[18][843],u_xpb_out[19][843],u_xpb_out[20][843],u_xpb_out[21][843],u_xpb_out[22][843],u_xpb_out[23][843],u_xpb_out[24][843],u_xpb_out[25][843],u_xpb_out[26][843],u_xpb_out[27][843],u_xpb_out[28][843],u_xpb_out[29][843],u_xpb_out[30][843],u_xpb_out[31][843],u_xpb_out[32][843],u_xpb_out[33][843],u_xpb_out[34][843],u_xpb_out[35][843],u_xpb_out[36][843],u_xpb_out[37][843],u_xpb_out[38][843],u_xpb_out[39][843],u_xpb_out[40][843],u_xpb_out[41][843],u_xpb_out[42][843],u_xpb_out[43][843],u_xpb_out[44][843],u_xpb_out[45][843],u_xpb_out[46][843],u_xpb_out[47][843],u_xpb_out[48][843],u_xpb_out[49][843],u_xpb_out[50][843],u_xpb_out[51][843],u_xpb_out[52][843],u_xpb_out[53][843],u_xpb_out[54][843],u_xpb_out[55][843],u_xpb_out[56][843],u_xpb_out[57][843],u_xpb_out[58][843],u_xpb_out[59][843],u_xpb_out[60][843],u_xpb_out[61][843],u_xpb_out[62][843],u_xpb_out[63][843],u_xpb_out[64][843],u_xpb_out[65][843],u_xpb_out[66][843],u_xpb_out[67][843],u_xpb_out[68][843],u_xpb_out[69][843],u_xpb_out[70][843],u_xpb_out[71][843],u_xpb_out[72][843],u_xpb_out[73][843],u_xpb_out[74][843],u_xpb_out[75][843],u_xpb_out[76][843],u_xpb_out[77][843],u_xpb_out[78][843],u_xpb_out[79][843],u_xpb_out[80][843],u_xpb_out[81][843],u_xpb_out[82][843],u_xpb_out[83][843],u_xpb_out[84][843],u_xpb_out[85][843],u_xpb_out[86][843],u_xpb_out[87][843],u_xpb_out[88][843],u_xpb_out[89][843],u_xpb_out[90][843],u_xpb_out[91][843],u_xpb_out[92][843],u_xpb_out[93][843],u_xpb_out[94][843],u_xpb_out[95][843],u_xpb_out[96][843],u_xpb_out[97][843],u_xpb_out[98][843],u_xpb_out[99][843],u_xpb_out[100][843],u_xpb_out[101][843],u_xpb_out[102][843],u_xpb_out[103][843],u_xpb_out[104][843],u_xpb_out[105][843]};

assign col_out_844 = {u_xpb_out[0][844],u_xpb_out[1][844],u_xpb_out[2][844],u_xpb_out[3][844],u_xpb_out[4][844],u_xpb_out[5][844],u_xpb_out[6][844],u_xpb_out[7][844],u_xpb_out[8][844],u_xpb_out[9][844],u_xpb_out[10][844],u_xpb_out[11][844],u_xpb_out[12][844],u_xpb_out[13][844],u_xpb_out[14][844],u_xpb_out[15][844],u_xpb_out[16][844],u_xpb_out[17][844],u_xpb_out[18][844],u_xpb_out[19][844],u_xpb_out[20][844],u_xpb_out[21][844],u_xpb_out[22][844],u_xpb_out[23][844],u_xpb_out[24][844],u_xpb_out[25][844],u_xpb_out[26][844],u_xpb_out[27][844],u_xpb_out[28][844],u_xpb_out[29][844],u_xpb_out[30][844],u_xpb_out[31][844],u_xpb_out[32][844],u_xpb_out[33][844],u_xpb_out[34][844],u_xpb_out[35][844],u_xpb_out[36][844],u_xpb_out[37][844],u_xpb_out[38][844],u_xpb_out[39][844],u_xpb_out[40][844],u_xpb_out[41][844],u_xpb_out[42][844],u_xpb_out[43][844],u_xpb_out[44][844],u_xpb_out[45][844],u_xpb_out[46][844],u_xpb_out[47][844],u_xpb_out[48][844],u_xpb_out[49][844],u_xpb_out[50][844],u_xpb_out[51][844],u_xpb_out[52][844],u_xpb_out[53][844],u_xpb_out[54][844],u_xpb_out[55][844],u_xpb_out[56][844],u_xpb_out[57][844],u_xpb_out[58][844],u_xpb_out[59][844],u_xpb_out[60][844],u_xpb_out[61][844],u_xpb_out[62][844],u_xpb_out[63][844],u_xpb_out[64][844],u_xpb_out[65][844],u_xpb_out[66][844],u_xpb_out[67][844],u_xpb_out[68][844],u_xpb_out[69][844],u_xpb_out[70][844],u_xpb_out[71][844],u_xpb_out[72][844],u_xpb_out[73][844],u_xpb_out[74][844],u_xpb_out[75][844],u_xpb_out[76][844],u_xpb_out[77][844],u_xpb_out[78][844],u_xpb_out[79][844],u_xpb_out[80][844],u_xpb_out[81][844],u_xpb_out[82][844],u_xpb_out[83][844],u_xpb_out[84][844],u_xpb_out[85][844],u_xpb_out[86][844],u_xpb_out[87][844],u_xpb_out[88][844],u_xpb_out[89][844],u_xpb_out[90][844],u_xpb_out[91][844],u_xpb_out[92][844],u_xpb_out[93][844],u_xpb_out[94][844],u_xpb_out[95][844],u_xpb_out[96][844],u_xpb_out[97][844],u_xpb_out[98][844],u_xpb_out[99][844],u_xpb_out[100][844],u_xpb_out[101][844],u_xpb_out[102][844],u_xpb_out[103][844],u_xpb_out[104][844],u_xpb_out[105][844]};

assign col_out_845 = {u_xpb_out[0][845],u_xpb_out[1][845],u_xpb_out[2][845],u_xpb_out[3][845],u_xpb_out[4][845],u_xpb_out[5][845],u_xpb_out[6][845],u_xpb_out[7][845],u_xpb_out[8][845],u_xpb_out[9][845],u_xpb_out[10][845],u_xpb_out[11][845],u_xpb_out[12][845],u_xpb_out[13][845],u_xpb_out[14][845],u_xpb_out[15][845],u_xpb_out[16][845],u_xpb_out[17][845],u_xpb_out[18][845],u_xpb_out[19][845],u_xpb_out[20][845],u_xpb_out[21][845],u_xpb_out[22][845],u_xpb_out[23][845],u_xpb_out[24][845],u_xpb_out[25][845],u_xpb_out[26][845],u_xpb_out[27][845],u_xpb_out[28][845],u_xpb_out[29][845],u_xpb_out[30][845],u_xpb_out[31][845],u_xpb_out[32][845],u_xpb_out[33][845],u_xpb_out[34][845],u_xpb_out[35][845],u_xpb_out[36][845],u_xpb_out[37][845],u_xpb_out[38][845],u_xpb_out[39][845],u_xpb_out[40][845],u_xpb_out[41][845],u_xpb_out[42][845],u_xpb_out[43][845],u_xpb_out[44][845],u_xpb_out[45][845],u_xpb_out[46][845],u_xpb_out[47][845],u_xpb_out[48][845],u_xpb_out[49][845],u_xpb_out[50][845],u_xpb_out[51][845],u_xpb_out[52][845],u_xpb_out[53][845],u_xpb_out[54][845],u_xpb_out[55][845],u_xpb_out[56][845],u_xpb_out[57][845],u_xpb_out[58][845],u_xpb_out[59][845],u_xpb_out[60][845],u_xpb_out[61][845],u_xpb_out[62][845],u_xpb_out[63][845],u_xpb_out[64][845],u_xpb_out[65][845],u_xpb_out[66][845],u_xpb_out[67][845],u_xpb_out[68][845],u_xpb_out[69][845],u_xpb_out[70][845],u_xpb_out[71][845],u_xpb_out[72][845],u_xpb_out[73][845],u_xpb_out[74][845],u_xpb_out[75][845],u_xpb_out[76][845],u_xpb_out[77][845],u_xpb_out[78][845],u_xpb_out[79][845],u_xpb_out[80][845],u_xpb_out[81][845],u_xpb_out[82][845],u_xpb_out[83][845],u_xpb_out[84][845],u_xpb_out[85][845],u_xpb_out[86][845],u_xpb_out[87][845],u_xpb_out[88][845],u_xpb_out[89][845],u_xpb_out[90][845],u_xpb_out[91][845],u_xpb_out[92][845],u_xpb_out[93][845],u_xpb_out[94][845],u_xpb_out[95][845],u_xpb_out[96][845],u_xpb_out[97][845],u_xpb_out[98][845],u_xpb_out[99][845],u_xpb_out[100][845],u_xpb_out[101][845],u_xpb_out[102][845],u_xpb_out[103][845],u_xpb_out[104][845],u_xpb_out[105][845]};

assign col_out_846 = {u_xpb_out[0][846],u_xpb_out[1][846],u_xpb_out[2][846],u_xpb_out[3][846],u_xpb_out[4][846],u_xpb_out[5][846],u_xpb_out[6][846],u_xpb_out[7][846],u_xpb_out[8][846],u_xpb_out[9][846],u_xpb_out[10][846],u_xpb_out[11][846],u_xpb_out[12][846],u_xpb_out[13][846],u_xpb_out[14][846],u_xpb_out[15][846],u_xpb_out[16][846],u_xpb_out[17][846],u_xpb_out[18][846],u_xpb_out[19][846],u_xpb_out[20][846],u_xpb_out[21][846],u_xpb_out[22][846],u_xpb_out[23][846],u_xpb_out[24][846],u_xpb_out[25][846],u_xpb_out[26][846],u_xpb_out[27][846],u_xpb_out[28][846],u_xpb_out[29][846],u_xpb_out[30][846],u_xpb_out[31][846],u_xpb_out[32][846],u_xpb_out[33][846],u_xpb_out[34][846],u_xpb_out[35][846],u_xpb_out[36][846],u_xpb_out[37][846],u_xpb_out[38][846],u_xpb_out[39][846],u_xpb_out[40][846],u_xpb_out[41][846],u_xpb_out[42][846],u_xpb_out[43][846],u_xpb_out[44][846],u_xpb_out[45][846],u_xpb_out[46][846],u_xpb_out[47][846],u_xpb_out[48][846],u_xpb_out[49][846],u_xpb_out[50][846],u_xpb_out[51][846],u_xpb_out[52][846],u_xpb_out[53][846],u_xpb_out[54][846],u_xpb_out[55][846],u_xpb_out[56][846],u_xpb_out[57][846],u_xpb_out[58][846],u_xpb_out[59][846],u_xpb_out[60][846],u_xpb_out[61][846],u_xpb_out[62][846],u_xpb_out[63][846],u_xpb_out[64][846],u_xpb_out[65][846],u_xpb_out[66][846],u_xpb_out[67][846],u_xpb_out[68][846],u_xpb_out[69][846],u_xpb_out[70][846],u_xpb_out[71][846],u_xpb_out[72][846],u_xpb_out[73][846],u_xpb_out[74][846],u_xpb_out[75][846],u_xpb_out[76][846],u_xpb_out[77][846],u_xpb_out[78][846],u_xpb_out[79][846],u_xpb_out[80][846],u_xpb_out[81][846],u_xpb_out[82][846],u_xpb_out[83][846],u_xpb_out[84][846],u_xpb_out[85][846],u_xpb_out[86][846],u_xpb_out[87][846],u_xpb_out[88][846],u_xpb_out[89][846],u_xpb_out[90][846],u_xpb_out[91][846],u_xpb_out[92][846],u_xpb_out[93][846],u_xpb_out[94][846],u_xpb_out[95][846],u_xpb_out[96][846],u_xpb_out[97][846],u_xpb_out[98][846],u_xpb_out[99][846],u_xpb_out[100][846],u_xpb_out[101][846],u_xpb_out[102][846],u_xpb_out[103][846],u_xpb_out[104][846],u_xpb_out[105][846]};

assign col_out_847 = {u_xpb_out[0][847],u_xpb_out[1][847],u_xpb_out[2][847],u_xpb_out[3][847],u_xpb_out[4][847],u_xpb_out[5][847],u_xpb_out[6][847],u_xpb_out[7][847],u_xpb_out[8][847],u_xpb_out[9][847],u_xpb_out[10][847],u_xpb_out[11][847],u_xpb_out[12][847],u_xpb_out[13][847],u_xpb_out[14][847],u_xpb_out[15][847],u_xpb_out[16][847],u_xpb_out[17][847],u_xpb_out[18][847],u_xpb_out[19][847],u_xpb_out[20][847],u_xpb_out[21][847],u_xpb_out[22][847],u_xpb_out[23][847],u_xpb_out[24][847],u_xpb_out[25][847],u_xpb_out[26][847],u_xpb_out[27][847],u_xpb_out[28][847],u_xpb_out[29][847],u_xpb_out[30][847],u_xpb_out[31][847],u_xpb_out[32][847],u_xpb_out[33][847],u_xpb_out[34][847],u_xpb_out[35][847],u_xpb_out[36][847],u_xpb_out[37][847],u_xpb_out[38][847],u_xpb_out[39][847],u_xpb_out[40][847],u_xpb_out[41][847],u_xpb_out[42][847],u_xpb_out[43][847],u_xpb_out[44][847],u_xpb_out[45][847],u_xpb_out[46][847],u_xpb_out[47][847],u_xpb_out[48][847],u_xpb_out[49][847],u_xpb_out[50][847],u_xpb_out[51][847],u_xpb_out[52][847],u_xpb_out[53][847],u_xpb_out[54][847],u_xpb_out[55][847],u_xpb_out[56][847],u_xpb_out[57][847],u_xpb_out[58][847],u_xpb_out[59][847],u_xpb_out[60][847],u_xpb_out[61][847],u_xpb_out[62][847],u_xpb_out[63][847],u_xpb_out[64][847],u_xpb_out[65][847],u_xpb_out[66][847],u_xpb_out[67][847],u_xpb_out[68][847],u_xpb_out[69][847],u_xpb_out[70][847],u_xpb_out[71][847],u_xpb_out[72][847],u_xpb_out[73][847],u_xpb_out[74][847],u_xpb_out[75][847],u_xpb_out[76][847],u_xpb_out[77][847],u_xpb_out[78][847],u_xpb_out[79][847],u_xpb_out[80][847],u_xpb_out[81][847],u_xpb_out[82][847],u_xpb_out[83][847],u_xpb_out[84][847],u_xpb_out[85][847],u_xpb_out[86][847],u_xpb_out[87][847],u_xpb_out[88][847],u_xpb_out[89][847],u_xpb_out[90][847],u_xpb_out[91][847],u_xpb_out[92][847],u_xpb_out[93][847],u_xpb_out[94][847],u_xpb_out[95][847],u_xpb_out[96][847],u_xpb_out[97][847],u_xpb_out[98][847],u_xpb_out[99][847],u_xpb_out[100][847],u_xpb_out[101][847],u_xpb_out[102][847],u_xpb_out[103][847],u_xpb_out[104][847],u_xpb_out[105][847]};

assign col_out_848 = {u_xpb_out[0][848],u_xpb_out[1][848],u_xpb_out[2][848],u_xpb_out[3][848],u_xpb_out[4][848],u_xpb_out[5][848],u_xpb_out[6][848],u_xpb_out[7][848],u_xpb_out[8][848],u_xpb_out[9][848],u_xpb_out[10][848],u_xpb_out[11][848],u_xpb_out[12][848],u_xpb_out[13][848],u_xpb_out[14][848],u_xpb_out[15][848],u_xpb_out[16][848],u_xpb_out[17][848],u_xpb_out[18][848],u_xpb_out[19][848],u_xpb_out[20][848],u_xpb_out[21][848],u_xpb_out[22][848],u_xpb_out[23][848],u_xpb_out[24][848],u_xpb_out[25][848],u_xpb_out[26][848],u_xpb_out[27][848],u_xpb_out[28][848],u_xpb_out[29][848],u_xpb_out[30][848],u_xpb_out[31][848],u_xpb_out[32][848],u_xpb_out[33][848],u_xpb_out[34][848],u_xpb_out[35][848],u_xpb_out[36][848],u_xpb_out[37][848],u_xpb_out[38][848],u_xpb_out[39][848],u_xpb_out[40][848],u_xpb_out[41][848],u_xpb_out[42][848],u_xpb_out[43][848],u_xpb_out[44][848],u_xpb_out[45][848],u_xpb_out[46][848],u_xpb_out[47][848],u_xpb_out[48][848],u_xpb_out[49][848],u_xpb_out[50][848],u_xpb_out[51][848],u_xpb_out[52][848],u_xpb_out[53][848],u_xpb_out[54][848],u_xpb_out[55][848],u_xpb_out[56][848],u_xpb_out[57][848],u_xpb_out[58][848],u_xpb_out[59][848],u_xpb_out[60][848],u_xpb_out[61][848],u_xpb_out[62][848],u_xpb_out[63][848],u_xpb_out[64][848],u_xpb_out[65][848],u_xpb_out[66][848],u_xpb_out[67][848],u_xpb_out[68][848],u_xpb_out[69][848],u_xpb_out[70][848],u_xpb_out[71][848],u_xpb_out[72][848],u_xpb_out[73][848],u_xpb_out[74][848],u_xpb_out[75][848],u_xpb_out[76][848],u_xpb_out[77][848],u_xpb_out[78][848],u_xpb_out[79][848],u_xpb_out[80][848],u_xpb_out[81][848],u_xpb_out[82][848],u_xpb_out[83][848],u_xpb_out[84][848],u_xpb_out[85][848],u_xpb_out[86][848],u_xpb_out[87][848],u_xpb_out[88][848],u_xpb_out[89][848],u_xpb_out[90][848],u_xpb_out[91][848],u_xpb_out[92][848],u_xpb_out[93][848],u_xpb_out[94][848],u_xpb_out[95][848],u_xpb_out[96][848],u_xpb_out[97][848],u_xpb_out[98][848],u_xpb_out[99][848],u_xpb_out[100][848],u_xpb_out[101][848],u_xpb_out[102][848],u_xpb_out[103][848],u_xpb_out[104][848],u_xpb_out[105][848]};

assign col_out_849 = {u_xpb_out[0][849],u_xpb_out[1][849],u_xpb_out[2][849],u_xpb_out[3][849],u_xpb_out[4][849],u_xpb_out[5][849],u_xpb_out[6][849],u_xpb_out[7][849],u_xpb_out[8][849],u_xpb_out[9][849],u_xpb_out[10][849],u_xpb_out[11][849],u_xpb_out[12][849],u_xpb_out[13][849],u_xpb_out[14][849],u_xpb_out[15][849],u_xpb_out[16][849],u_xpb_out[17][849],u_xpb_out[18][849],u_xpb_out[19][849],u_xpb_out[20][849],u_xpb_out[21][849],u_xpb_out[22][849],u_xpb_out[23][849],u_xpb_out[24][849],u_xpb_out[25][849],u_xpb_out[26][849],u_xpb_out[27][849],u_xpb_out[28][849],u_xpb_out[29][849],u_xpb_out[30][849],u_xpb_out[31][849],u_xpb_out[32][849],u_xpb_out[33][849],u_xpb_out[34][849],u_xpb_out[35][849],u_xpb_out[36][849],u_xpb_out[37][849],u_xpb_out[38][849],u_xpb_out[39][849],u_xpb_out[40][849],u_xpb_out[41][849],u_xpb_out[42][849],u_xpb_out[43][849],u_xpb_out[44][849],u_xpb_out[45][849],u_xpb_out[46][849],u_xpb_out[47][849],u_xpb_out[48][849],u_xpb_out[49][849],u_xpb_out[50][849],u_xpb_out[51][849],u_xpb_out[52][849],u_xpb_out[53][849],u_xpb_out[54][849],u_xpb_out[55][849],u_xpb_out[56][849],u_xpb_out[57][849],u_xpb_out[58][849],u_xpb_out[59][849],u_xpb_out[60][849],u_xpb_out[61][849],u_xpb_out[62][849],u_xpb_out[63][849],u_xpb_out[64][849],u_xpb_out[65][849],u_xpb_out[66][849],u_xpb_out[67][849],u_xpb_out[68][849],u_xpb_out[69][849],u_xpb_out[70][849],u_xpb_out[71][849],u_xpb_out[72][849],u_xpb_out[73][849],u_xpb_out[74][849],u_xpb_out[75][849],u_xpb_out[76][849],u_xpb_out[77][849],u_xpb_out[78][849],u_xpb_out[79][849],u_xpb_out[80][849],u_xpb_out[81][849],u_xpb_out[82][849],u_xpb_out[83][849],u_xpb_out[84][849],u_xpb_out[85][849],u_xpb_out[86][849],u_xpb_out[87][849],u_xpb_out[88][849],u_xpb_out[89][849],u_xpb_out[90][849],u_xpb_out[91][849],u_xpb_out[92][849],u_xpb_out[93][849],u_xpb_out[94][849],u_xpb_out[95][849],u_xpb_out[96][849],u_xpb_out[97][849],u_xpb_out[98][849],u_xpb_out[99][849],u_xpb_out[100][849],u_xpb_out[101][849],u_xpb_out[102][849],u_xpb_out[103][849],u_xpb_out[104][849],u_xpb_out[105][849]};

assign col_out_850 = {u_xpb_out[0][850],u_xpb_out[1][850],u_xpb_out[2][850],u_xpb_out[3][850],u_xpb_out[4][850],u_xpb_out[5][850],u_xpb_out[6][850],u_xpb_out[7][850],u_xpb_out[8][850],u_xpb_out[9][850],u_xpb_out[10][850],u_xpb_out[11][850],u_xpb_out[12][850],u_xpb_out[13][850],u_xpb_out[14][850],u_xpb_out[15][850],u_xpb_out[16][850],u_xpb_out[17][850],u_xpb_out[18][850],u_xpb_out[19][850],u_xpb_out[20][850],u_xpb_out[21][850],u_xpb_out[22][850],u_xpb_out[23][850],u_xpb_out[24][850],u_xpb_out[25][850],u_xpb_out[26][850],u_xpb_out[27][850],u_xpb_out[28][850],u_xpb_out[29][850],u_xpb_out[30][850],u_xpb_out[31][850],u_xpb_out[32][850],u_xpb_out[33][850],u_xpb_out[34][850],u_xpb_out[35][850],u_xpb_out[36][850],u_xpb_out[37][850],u_xpb_out[38][850],u_xpb_out[39][850],u_xpb_out[40][850],u_xpb_out[41][850],u_xpb_out[42][850],u_xpb_out[43][850],u_xpb_out[44][850],u_xpb_out[45][850],u_xpb_out[46][850],u_xpb_out[47][850],u_xpb_out[48][850],u_xpb_out[49][850],u_xpb_out[50][850],u_xpb_out[51][850],u_xpb_out[52][850],u_xpb_out[53][850],u_xpb_out[54][850],u_xpb_out[55][850],u_xpb_out[56][850],u_xpb_out[57][850],u_xpb_out[58][850],u_xpb_out[59][850],u_xpb_out[60][850],u_xpb_out[61][850],u_xpb_out[62][850],u_xpb_out[63][850],u_xpb_out[64][850],u_xpb_out[65][850],u_xpb_out[66][850],u_xpb_out[67][850],u_xpb_out[68][850],u_xpb_out[69][850],u_xpb_out[70][850],u_xpb_out[71][850],u_xpb_out[72][850],u_xpb_out[73][850],u_xpb_out[74][850],u_xpb_out[75][850],u_xpb_out[76][850],u_xpb_out[77][850],u_xpb_out[78][850],u_xpb_out[79][850],u_xpb_out[80][850],u_xpb_out[81][850],u_xpb_out[82][850],u_xpb_out[83][850],u_xpb_out[84][850],u_xpb_out[85][850],u_xpb_out[86][850],u_xpb_out[87][850],u_xpb_out[88][850],u_xpb_out[89][850],u_xpb_out[90][850],u_xpb_out[91][850],u_xpb_out[92][850],u_xpb_out[93][850],u_xpb_out[94][850],u_xpb_out[95][850],u_xpb_out[96][850],u_xpb_out[97][850],u_xpb_out[98][850],u_xpb_out[99][850],u_xpb_out[100][850],u_xpb_out[101][850],u_xpb_out[102][850],u_xpb_out[103][850],u_xpb_out[104][850],u_xpb_out[105][850]};

assign col_out_851 = {u_xpb_out[0][851],u_xpb_out[1][851],u_xpb_out[2][851],u_xpb_out[3][851],u_xpb_out[4][851],u_xpb_out[5][851],u_xpb_out[6][851],u_xpb_out[7][851],u_xpb_out[8][851],u_xpb_out[9][851],u_xpb_out[10][851],u_xpb_out[11][851],u_xpb_out[12][851],u_xpb_out[13][851],u_xpb_out[14][851],u_xpb_out[15][851],u_xpb_out[16][851],u_xpb_out[17][851],u_xpb_out[18][851],u_xpb_out[19][851],u_xpb_out[20][851],u_xpb_out[21][851],u_xpb_out[22][851],u_xpb_out[23][851],u_xpb_out[24][851],u_xpb_out[25][851],u_xpb_out[26][851],u_xpb_out[27][851],u_xpb_out[28][851],u_xpb_out[29][851],u_xpb_out[30][851],u_xpb_out[31][851],u_xpb_out[32][851],u_xpb_out[33][851],u_xpb_out[34][851],u_xpb_out[35][851],u_xpb_out[36][851],u_xpb_out[37][851],u_xpb_out[38][851],u_xpb_out[39][851],u_xpb_out[40][851],u_xpb_out[41][851],u_xpb_out[42][851],u_xpb_out[43][851],u_xpb_out[44][851],u_xpb_out[45][851],u_xpb_out[46][851],u_xpb_out[47][851],u_xpb_out[48][851],u_xpb_out[49][851],u_xpb_out[50][851],u_xpb_out[51][851],u_xpb_out[52][851],u_xpb_out[53][851],u_xpb_out[54][851],u_xpb_out[55][851],u_xpb_out[56][851],u_xpb_out[57][851],u_xpb_out[58][851],u_xpb_out[59][851],u_xpb_out[60][851],u_xpb_out[61][851],u_xpb_out[62][851],u_xpb_out[63][851],u_xpb_out[64][851],u_xpb_out[65][851],u_xpb_out[66][851],u_xpb_out[67][851],u_xpb_out[68][851],u_xpb_out[69][851],u_xpb_out[70][851],u_xpb_out[71][851],u_xpb_out[72][851],u_xpb_out[73][851],u_xpb_out[74][851],u_xpb_out[75][851],u_xpb_out[76][851],u_xpb_out[77][851],u_xpb_out[78][851],u_xpb_out[79][851],u_xpb_out[80][851],u_xpb_out[81][851],u_xpb_out[82][851],u_xpb_out[83][851],u_xpb_out[84][851],u_xpb_out[85][851],u_xpb_out[86][851],u_xpb_out[87][851],u_xpb_out[88][851],u_xpb_out[89][851],u_xpb_out[90][851],u_xpb_out[91][851],u_xpb_out[92][851],u_xpb_out[93][851],u_xpb_out[94][851],u_xpb_out[95][851],u_xpb_out[96][851],u_xpb_out[97][851],u_xpb_out[98][851],u_xpb_out[99][851],u_xpb_out[100][851],u_xpb_out[101][851],u_xpb_out[102][851],u_xpb_out[103][851],u_xpb_out[104][851],u_xpb_out[105][851]};

assign col_out_852 = {u_xpb_out[0][852],u_xpb_out[1][852],u_xpb_out[2][852],u_xpb_out[3][852],u_xpb_out[4][852],u_xpb_out[5][852],u_xpb_out[6][852],u_xpb_out[7][852],u_xpb_out[8][852],u_xpb_out[9][852],u_xpb_out[10][852],u_xpb_out[11][852],u_xpb_out[12][852],u_xpb_out[13][852],u_xpb_out[14][852],u_xpb_out[15][852],u_xpb_out[16][852],u_xpb_out[17][852],u_xpb_out[18][852],u_xpb_out[19][852],u_xpb_out[20][852],u_xpb_out[21][852],u_xpb_out[22][852],u_xpb_out[23][852],u_xpb_out[24][852],u_xpb_out[25][852],u_xpb_out[26][852],u_xpb_out[27][852],u_xpb_out[28][852],u_xpb_out[29][852],u_xpb_out[30][852],u_xpb_out[31][852],u_xpb_out[32][852],u_xpb_out[33][852],u_xpb_out[34][852],u_xpb_out[35][852],u_xpb_out[36][852],u_xpb_out[37][852],u_xpb_out[38][852],u_xpb_out[39][852],u_xpb_out[40][852],u_xpb_out[41][852],u_xpb_out[42][852],u_xpb_out[43][852],u_xpb_out[44][852],u_xpb_out[45][852],u_xpb_out[46][852],u_xpb_out[47][852],u_xpb_out[48][852],u_xpb_out[49][852],u_xpb_out[50][852],u_xpb_out[51][852],u_xpb_out[52][852],u_xpb_out[53][852],u_xpb_out[54][852],u_xpb_out[55][852],u_xpb_out[56][852],u_xpb_out[57][852],u_xpb_out[58][852],u_xpb_out[59][852],u_xpb_out[60][852],u_xpb_out[61][852],u_xpb_out[62][852],u_xpb_out[63][852],u_xpb_out[64][852],u_xpb_out[65][852],u_xpb_out[66][852],u_xpb_out[67][852],u_xpb_out[68][852],u_xpb_out[69][852],u_xpb_out[70][852],u_xpb_out[71][852],u_xpb_out[72][852],u_xpb_out[73][852],u_xpb_out[74][852],u_xpb_out[75][852],u_xpb_out[76][852],u_xpb_out[77][852],u_xpb_out[78][852],u_xpb_out[79][852],u_xpb_out[80][852],u_xpb_out[81][852],u_xpb_out[82][852],u_xpb_out[83][852],u_xpb_out[84][852],u_xpb_out[85][852],u_xpb_out[86][852],u_xpb_out[87][852],u_xpb_out[88][852],u_xpb_out[89][852],u_xpb_out[90][852],u_xpb_out[91][852],u_xpb_out[92][852],u_xpb_out[93][852],u_xpb_out[94][852],u_xpb_out[95][852],u_xpb_out[96][852],u_xpb_out[97][852],u_xpb_out[98][852],u_xpb_out[99][852],u_xpb_out[100][852],u_xpb_out[101][852],u_xpb_out[102][852],u_xpb_out[103][852],u_xpb_out[104][852],u_xpb_out[105][852]};

assign col_out_853 = {u_xpb_out[0][853],u_xpb_out[1][853],u_xpb_out[2][853],u_xpb_out[3][853],u_xpb_out[4][853],u_xpb_out[5][853],u_xpb_out[6][853],u_xpb_out[7][853],u_xpb_out[8][853],u_xpb_out[9][853],u_xpb_out[10][853],u_xpb_out[11][853],u_xpb_out[12][853],u_xpb_out[13][853],u_xpb_out[14][853],u_xpb_out[15][853],u_xpb_out[16][853],u_xpb_out[17][853],u_xpb_out[18][853],u_xpb_out[19][853],u_xpb_out[20][853],u_xpb_out[21][853],u_xpb_out[22][853],u_xpb_out[23][853],u_xpb_out[24][853],u_xpb_out[25][853],u_xpb_out[26][853],u_xpb_out[27][853],u_xpb_out[28][853],u_xpb_out[29][853],u_xpb_out[30][853],u_xpb_out[31][853],u_xpb_out[32][853],u_xpb_out[33][853],u_xpb_out[34][853],u_xpb_out[35][853],u_xpb_out[36][853],u_xpb_out[37][853],u_xpb_out[38][853],u_xpb_out[39][853],u_xpb_out[40][853],u_xpb_out[41][853],u_xpb_out[42][853],u_xpb_out[43][853],u_xpb_out[44][853],u_xpb_out[45][853],u_xpb_out[46][853],u_xpb_out[47][853],u_xpb_out[48][853],u_xpb_out[49][853],u_xpb_out[50][853],u_xpb_out[51][853],u_xpb_out[52][853],u_xpb_out[53][853],u_xpb_out[54][853],u_xpb_out[55][853],u_xpb_out[56][853],u_xpb_out[57][853],u_xpb_out[58][853],u_xpb_out[59][853],u_xpb_out[60][853],u_xpb_out[61][853],u_xpb_out[62][853],u_xpb_out[63][853],u_xpb_out[64][853],u_xpb_out[65][853],u_xpb_out[66][853],u_xpb_out[67][853],u_xpb_out[68][853],u_xpb_out[69][853],u_xpb_out[70][853],u_xpb_out[71][853],u_xpb_out[72][853],u_xpb_out[73][853],u_xpb_out[74][853],u_xpb_out[75][853],u_xpb_out[76][853],u_xpb_out[77][853],u_xpb_out[78][853],u_xpb_out[79][853],u_xpb_out[80][853],u_xpb_out[81][853],u_xpb_out[82][853],u_xpb_out[83][853],u_xpb_out[84][853],u_xpb_out[85][853],u_xpb_out[86][853],u_xpb_out[87][853],u_xpb_out[88][853],u_xpb_out[89][853],u_xpb_out[90][853],u_xpb_out[91][853],u_xpb_out[92][853],u_xpb_out[93][853],u_xpb_out[94][853],u_xpb_out[95][853],u_xpb_out[96][853],u_xpb_out[97][853],u_xpb_out[98][853],u_xpb_out[99][853],u_xpb_out[100][853],u_xpb_out[101][853],u_xpb_out[102][853],u_xpb_out[103][853],u_xpb_out[104][853],u_xpb_out[105][853]};

assign col_out_854 = {u_xpb_out[0][854],u_xpb_out[1][854],u_xpb_out[2][854],u_xpb_out[3][854],u_xpb_out[4][854],u_xpb_out[5][854],u_xpb_out[6][854],u_xpb_out[7][854],u_xpb_out[8][854],u_xpb_out[9][854],u_xpb_out[10][854],u_xpb_out[11][854],u_xpb_out[12][854],u_xpb_out[13][854],u_xpb_out[14][854],u_xpb_out[15][854],u_xpb_out[16][854],u_xpb_out[17][854],u_xpb_out[18][854],u_xpb_out[19][854],u_xpb_out[20][854],u_xpb_out[21][854],u_xpb_out[22][854],u_xpb_out[23][854],u_xpb_out[24][854],u_xpb_out[25][854],u_xpb_out[26][854],u_xpb_out[27][854],u_xpb_out[28][854],u_xpb_out[29][854],u_xpb_out[30][854],u_xpb_out[31][854],u_xpb_out[32][854],u_xpb_out[33][854],u_xpb_out[34][854],u_xpb_out[35][854],u_xpb_out[36][854],u_xpb_out[37][854],u_xpb_out[38][854],u_xpb_out[39][854],u_xpb_out[40][854],u_xpb_out[41][854],u_xpb_out[42][854],u_xpb_out[43][854],u_xpb_out[44][854],u_xpb_out[45][854],u_xpb_out[46][854],u_xpb_out[47][854],u_xpb_out[48][854],u_xpb_out[49][854],u_xpb_out[50][854],u_xpb_out[51][854],u_xpb_out[52][854],u_xpb_out[53][854],u_xpb_out[54][854],u_xpb_out[55][854],u_xpb_out[56][854],u_xpb_out[57][854],u_xpb_out[58][854],u_xpb_out[59][854],u_xpb_out[60][854],u_xpb_out[61][854],u_xpb_out[62][854],u_xpb_out[63][854],u_xpb_out[64][854],u_xpb_out[65][854],u_xpb_out[66][854],u_xpb_out[67][854],u_xpb_out[68][854],u_xpb_out[69][854],u_xpb_out[70][854],u_xpb_out[71][854],u_xpb_out[72][854],u_xpb_out[73][854],u_xpb_out[74][854],u_xpb_out[75][854],u_xpb_out[76][854],u_xpb_out[77][854],u_xpb_out[78][854],u_xpb_out[79][854],u_xpb_out[80][854],u_xpb_out[81][854],u_xpb_out[82][854],u_xpb_out[83][854],u_xpb_out[84][854],u_xpb_out[85][854],u_xpb_out[86][854],u_xpb_out[87][854],u_xpb_out[88][854],u_xpb_out[89][854],u_xpb_out[90][854],u_xpb_out[91][854],u_xpb_out[92][854],u_xpb_out[93][854],u_xpb_out[94][854],u_xpb_out[95][854],u_xpb_out[96][854],u_xpb_out[97][854],u_xpb_out[98][854],u_xpb_out[99][854],u_xpb_out[100][854],u_xpb_out[101][854],u_xpb_out[102][854],u_xpb_out[103][854],u_xpb_out[104][854],u_xpb_out[105][854]};

assign col_out_855 = {u_xpb_out[0][855],u_xpb_out[1][855],u_xpb_out[2][855],u_xpb_out[3][855],u_xpb_out[4][855],u_xpb_out[5][855],u_xpb_out[6][855],u_xpb_out[7][855],u_xpb_out[8][855],u_xpb_out[9][855],u_xpb_out[10][855],u_xpb_out[11][855],u_xpb_out[12][855],u_xpb_out[13][855],u_xpb_out[14][855],u_xpb_out[15][855],u_xpb_out[16][855],u_xpb_out[17][855],u_xpb_out[18][855],u_xpb_out[19][855],u_xpb_out[20][855],u_xpb_out[21][855],u_xpb_out[22][855],u_xpb_out[23][855],u_xpb_out[24][855],u_xpb_out[25][855],u_xpb_out[26][855],u_xpb_out[27][855],u_xpb_out[28][855],u_xpb_out[29][855],u_xpb_out[30][855],u_xpb_out[31][855],u_xpb_out[32][855],u_xpb_out[33][855],u_xpb_out[34][855],u_xpb_out[35][855],u_xpb_out[36][855],u_xpb_out[37][855],u_xpb_out[38][855],u_xpb_out[39][855],u_xpb_out[40][855],u_xpb_out[41][855],u_xpb_out[42][855],u_xpb_out[43][855],u_xpb_out[44][855],u_xpb_out[45][855],u_xpb_out[46][855],u_xpb_out[47][855],u_xpb_out[48][855],u_xpb_out[49][855],u_xpb_out[50][855],u_xpb_out[51][855],u_xpb_out[52][855],u_xpb_out[53][855],u_xpb_out[54][855],u_xpb_out[55][855],u_xpb_out[56][855],u_xpb_out[57][855],u_xpb_out[58][855],u_xpb_out[59][855],u_xpb_out[60][855],u_xpb_out[61][855],u_xpb_out[62][855],u_xpb_out[63][855],u_xpb_out[64][855],u_xpb_out[65][855],u_xpb_out[66][855],u_xpb_out[67][855],u_xpb_out[68][855],u_xpb_out[69][855],u_xpb_out[70][855],u_xpb_out[71][855],u_xpb_out[72][855],u_xpb_out[73][855],u_xpb_out[74][855],u_xpb_out[75][855],u_xpb_out[76][855],u_xpb_out[77][855],u_xpb_out[78][855],u_xpb_out[79][855],u_xpb_out[80][855],u_xpb_out[81][855],u_xpb_out[82][855],u_xpb_out[83][855],u_xpb_out[84][855],u_xpb_out[85][855],u_xpb_out[86][855],u_xpb_out[87][855],u_xpb_out[88][855],u_xpb_out[89][855],u_xpb_out[90][855],u_xpb_out[91][855],u_xpb_out[92][855],u_xpb_out[93][855],u_xpb_out[94][855],u_xpb_out[95][855],u_xpb_out[96][855],u_xpb_out[97][855],u_xpb_out[98][855],u_xpb_out[99][855],u_xpb_out[100][855],u_xpb_out[101][855],u_xpb_out[102][855],u_xpb_out[103][855],u_xpb_out[104][855],u_xpb_out[105][855]};

assign col_out_856 = {u_xpb_out[0][856],u_xpb_out[1][856],u_xpb_out[2][856],u_xpb_out[3][856],u_xpb_out[4][856],u_xpb_out[5][856],u_xpb_out[6][856],u_xpb_out[7][856],u_xpb_out[8][856],u_xpb_out[9][856],u_xpb_out[10][856],u_xpb_out[11][856],u_xpb_out[12][856],u_xpb_out[13][856],u_xpb_out[14][856],u_xpb_out[15][856],u_xpb_out[16][856],u_xpb_out[17][856],u_xpb_out[18][856],u_xpb_out[19][856],u_xpb_out[20][856],u_xpb_out[21][856],u_xpb_out[22][856],u_xpb_out[23][856],u_xpb_out[24][856],u_xpb_out[25][856],u_xpb_out[26][856],u_xpb_out[27][856],u_xpb_out[28][856],u_xpb_out[29][856],u_xpb_out[30][856],u_xpb_out[31][856],u_xpb_out[32][856],u_xpb_out[33][856],u_xpb_out[34][856],u_xpb_out[35][856],u_xpb_out[36][856],u_xpb_out[37][856],u_xpb_out[38][856],u_xpb_out[39][856],u_xpb_out[40][856],u_xpb_out[41][856],u_xpb_out[42][856],u_xpb_out[43][856],u_xpb_out[44][856],u_xpb_out[45][856],u_xpb_out[46][856],u_xpb_out[47][856],u_xpb_out[48][856],u_xpb_out[49][856],u_xpb_out[50][856],u_xpb_out[51][856],u_xpb_out[52][856],u_xpb_out[53][856],u_xpb_out[54][856],u_xpb_out[55][856],u_xpb_out[56][856],u_xpb_out[57][856],u_xpb_out[58][856],u_xpb_out[59][856],u_xpb_out[60][856],u_xpb_out[61][856],u_xpb_out[62][856],u_xpb_out[63][856],u_xpb_out[64][856],u_xpb_out[65][856],u_xpb_out[66][856],u_xpb_out[67][856],u_xpb_out[68][856],u_xpb_out[69][856],u_xpb_out[70][856],u_xpb_out[71][856],u_xpb_out[72][856],u_xpb_out[73][856],u_xpb_out[74][856],u_xpb_out[75][856],u_xpb_out[76][856],u_xpb_out[77][856],u_xpb_out[78][856],u_xpb_out[79][856],u_xpb_out[80][856],u_xpb_out[81][856],u_xpb_out[82][856],u_xpb_out[83][856],u_xpb_out[84][856],u_xpb_out[85][856],u_xpb_out[86][856],u_xpb_out[87][856],u_xpb_out[88][856],u_xpb_out[89][856],u_xpb_out[90][856],u_xpb_out[91][856],u_xpb_out[92][856],u_xpb_out[93][856],u_xpb_out[94][856],u_xpb_out[95][856],u_xpb_out[96][856],u_xpb_out[97][856],u_xpb_out[98][856],u_xpb_out[99][856],u_xpb_out[100][856],u_xpb_out[101][856],u_xpb_out[102][856],u_xpb_out[103][856],u_xpb_out[104][856],u_xpb_out[105][856]};

assign col_out_857 = {u_xpb_out[0][857],u_xpb_out[1][857],u_xpb_out[2][857],u_xpb_out[3][857],u_xpb_out[4][857],u_xpb_out[5][857],u_xpb_out[6][857],u_xpb_out[7][857],u_xpb_out[8][857],u_xpb_out[9][857],u_xpb_out[10][857],u_xpb_out[11][857],u_xpb_out[12][857],u_xpb_out[13][857],u_xpb_out[14][857],u_xpb_out[15][857],u_xpb_out[16][857],u_xpb_out[17][857],u_xpb_out[18][857],u_xpb_out[19][857],u_xpb_out[20][857],u_xpb_out[21][857],u_xpb_out[22][857],u_xpb_out[23][857],u_xpb_out[24][857],u_xpb_out[25][857],u_xpb_out[26][857],u_xpb_out[27][857],u_xpb_out[28][857],u_xpb_out[29][857],u_xpb_out[30][857],u_xpb_out[31][857],u_xpb_out[32][857],u_xpb_out[33][857],u_xpb_out[34][857],u_xpb_out[35][857],u_xpb_out[36][857],u_xpb_out[37][857],u_xpb_out[38][857],u_xpb_out[39][857],u_xpb_out[40][857],u_xpb_out[41][857],u_xpb_out[42][857],u_xpb_out[43][857],u_xpb_out[44][857],u_xpb_out[45][857],u_xpb_out[46][857],u_xpb_out[47][857],u_xpb_out[48][857],u_xpb_out[49][857],u_xpb_out[50][857],u_xpb_out[51][857],u_xpb_out[52][857],u_xpb_out[53][857],u_xpb_out[54][857],u_xpb_out[55][857],u_xpb_out[56][857],u_xpb_out[57][857],u_xpb_out[58][857],u_xpb_out[59][857],u_xpb_out[60][857],u_xpb_out[61][857],u_xpb_out[62][857],u_xpb_out[63][857],u_xpb_out[64][857],u_xpb_out[65][857],u_xpb_out[66][857],u_xpb_out[67][857],u_xpb_out[68][857],u_xpb_out[69][857],u_xpb_out[70][857],u_xpb_out[71][857],u_xpb_out[72][857],u_xpb_out[73][857],u_xpb_out[74][857],u_xpb_out[75][857],u_xpb_out[76][857],u_xpb_out[77][857],u_xpb_out[78][857],u_xpb_out[79][857],u_xpb_out[80][857],u_xpb_out[81][857],u_xpb_out[82][857],u_xpb_out[83][857],u_xpb_out[84][857],u_xpb_out[85][857],u_xpb_out[86][857],u_xpb_out[87][857],u_xpb_out[88][857],u_xpb_out[89][857],u_xpb_out[90][857],u_xpb_out[91][857],u_xpb_out[92][857],u_xpb_out[93][857],u_xpb_out[94][857],u_xpb_out[95][857],u_xpb_out[96][857],u_xpb_out[97][857],u_xpb_out[98][857],u_xpb_out[99][857],u_xpb_out[100][857],u_xpb_out[101][857],u_xpb_out[102][857],u_xpb_out[103][857],u_xpb_out[104][857],u_xpb_out[105][857]};

assign col_out_858 = {u_xpb_out[0][858],u_xpb_out[1][858],u_xpb_out[2][858],u_xpb_out[3][858],u_xpb_out[4][858],u_xpb_out[5][858],u_xpb_out[6][858],u_xpb_out[7][858],u_xpb_out[8][858],u_xpb_out[9][858],u_xpb_out[10][858],u_xpb_out[11][858],u_xpb_out[12][858],u_xpb_out[13][858],u_xpb_out[14][858],u_xpb_out[15][858],u_xpb_out[16][858],u_xpb_out[17][858],u_xpb_out[18][858],u_xpb_out[19][858],u_xpb_out[20][858],u_xpb_out[21][858],u_xpb_out[22][858],u_xpb_out[23][858],u_xpb_out[24][858],u_xpb_out[25][858],u_xpb_out[26][858],u_xpb_out[27][858],u_xpb_out[28][858],u_xpb_out[29][858],u_xpb_out[30][858],u_xpb_out[31][858],u_xpb_out[32][858],u_xpb_out[33][858],u_xpb_out[34][858],u_xpb_out[35][858],u_xpb_out[36][858],u_xpb_out[37][858],u_xpb_out[38][858],u_xpb_out[39][858],u_xpb_out[40][858],u_xpb_out[41][858],u_xpb_out[42][858],u_xpb_out[43][858],u_xpb_out[44][858],u_xpb_out[45][858],u_xpb_out[46][858],u_xpb_out[47][858],u_xpb_out[48][858],u_xpb_out[49][858],u_xpb_out[50][858],u_xpb_out[51][858],u_xpb_out[52][858],u_xpb_out[53][858],u_xpb_out[54][858],u_xpb_out[55][858],u_xpb_out[56][858],u_xpb_out[57][858],u_xpb_out[58][858],u_xpb_out[59][858],u_xpb_out[60][858],u_xpb_out[61][858],u_xpb_out[62][858],u_xpb_out[63][858],u_xpb_out[64][858],u_xpb_out[65][858],u_xpb_out[66][858],u_xpb_out[67][858],u_xpb_out[68][858],u_xpb_out[69][858],u_xpb_out[70][858],u_xpb_out[71][858],u_xpb_out[72][858],u_xpb_out[73][858],u_xpb_out[74][858],u_xpb_out[75][858],u_xpb_out[76][858],u_xpb_out[77][858],u_xpb_out[78][858],u_xpb_out[79][858],u_xpb_out[80][858],u_xpb_out[81][858],u_xpb_out[82][858],u_xpb_out[83][858],u_xpb_out[84][858],u_xpb_out[85][858],u_xpb_out[86][858],u_xpb_out[87][858],u_xpb_out[88][858],u_xpb_out[89][858],u_xpb_out[90][858],u_xpb_out[91][858],u_xpb_out[92][858],u_xpb_out[93][858],u_xpb_out[94][858],u_xpb_out[95][858],u_xpb_out[96][858],u_xpb_out[97][858],u_xpb_out[98][858],u_xpb_out[99][858],u_xpb_out[100][858],u_xpb_out[101][858],u_xpb_out[102][858],u_xpb_out[103][858],u_xpb_out[104][858],u_xpb_out[105][858]};

assign col_out_859 = {u_xpb_out[0][859],u_xpb_out[1][859],u_xpb_out[2][859],u_xpb_out[3][859],u_xpb_out[4][859],u_xpb_out[5][859],u_xpb_out[6][859],u_xpb_out[7][859],u_xpb_out[8][859],u_xpb_out[9][859],u_xpb_out[10][859],u_xpb_out[11][859],u_xpb_out[12][859],u_xpb_out[13][859],u_xpb_out[14][859],u_xpb_out[15][859],u_xpb_out[16][859],u_xpb_out[17][859],u_xpb_out[18][859],u_xpb_out[19][859],u_xpb_out[20][859],u_xpb_out[21][859],u_xpb_out[22][859],u_xpb_out[23][859],u_xpb_out[24][859],u_xpb_out[25][859],u_xpb_out[26][859],u_xpb_out[27][859],u_xpb_out[28][859],u_xpb_out[29][859],u_xpb_out[30][859],u_xpb_out[31][859],u_xpb_out[32][859],u_xpb_out[33][859],u_xpb_out[34][859],u_xpb_out[35][859],u_xpb_out[36][859],u_xpb_out[37][859],u_xpb_out[38][859],u_xpb_out[39][859],u_xpb_out[40][859],u_xpb_out[41][859],u_xpb_out[42][859],u_xpb_out[43][859],u_xpb_out[44][859],u_xpb_out[45][859],u_xpb_out[46][859],u_xpb_out[47][859],u_xpb_out[48][859],u_xpb_out[49][859],u_xpb_out[50][859],u_xpb_out[51][859],u_xpb_out[52][859],u_xpb_out[53][859],u_xpb_out[54][859],u_xpb_out[55][859],u_xpb_out[56][859],u_xpb_out[57][859],u_xpb_out[58][859],u_xpb_out[59][859],u_xpb_out[60][859],u_xpb_out[61][859],u_xpb_out[62][859],u_xpb_out[63][859],u_xpb_out[64][859],u_xpb_out[65][859],u_xpb_out[66][859],u_xpb_out[67][859],u_xpb_out[68][859],u_xpb_out[69][859],u_xpb_out[70][859],u_xpb_out[71][859],u_xpb_out[72][859],u_xpb_out[73][859],u_xpb_out[74][859],u_xpb_out[75][859],u_xpb_out[76][859],u_xpb_out[77][859],u_xpb_out[78][859],u_xpb_out[79][859],u_xpb_out[80][859],u_xpb_out[81][859],u_xpb_out[82][859],u_xpb_out[83][859],u_xpb_out[84][859],u_xpb_out[85][859],u_xpb_out[86][859],u_xpb_out[87][859],u_xpb_out[88][859],u_xpb_out[89][859],u_xpb_out[90][859],u_xpb_out[91][859],u_xpb_out[92][859],u_xpb_out[93][859],u_xpb_out[94][859],u_xpb_out[95][859],u_xpb_out[96][859],u_xpb_out[97][859],u_xpb_out[98][859],u_xpb_out[99][859],u_xpb_out[100][859],u_xpb_out[101][859],u_xpb_out[102][859],u_xpb_out[103][859],u_xpb_out[104][859],u_xpb_out[105][859]};

assign col_out_860 = {u_xpb_out[0][860],u_xpb_out[1][860],u_xpb_out[2][860],u_xpb_out[3][860],u_xpb_out[4][860],u_xpb_out[5][860],u_xpb_out[6][860],u_xpb_out[7][860],u_xpb_out[8][860],u_xpb_out[9][860],u_xpb_out[10][860],u_xpb_out[11][860],u_xpb_out[12][860],u_xpb_out[13][860],u_xpb_out[14][860],u_xpb_out[15][860],u_xpb_out[16][860],u_xpb_out[17][860],u_xpb_out[18][860],u_xpb_out[19][860],u_xpb_out[20][860],u_xpb_out[21][860],u_xpb_out[22][860],u_xpb_out[23][860],u_xpb_out[24][860],u_xpb_out[25][860],u_xpb_out[26][860],u_xpb_out[27][860],u_xpb_out[28][860],u_xpb_out[29][860],u_xpb_out[30][860],u_xpb_out[31][860],u_xpb_out[32][860],u_xpb_out[33][860],u_xpb_out[34][860],u_xpb_out[35][860],u_xpb_out[36][860],u_xpb_out[37][860],u_xpb_out[38][860],u_xpb_out[39][860],u_xpb_out[40][860],u_xpb_out[41][860],u_xpb_out[42][860],u_xpb_out[43][860],u_xpb_out[44][860],u_xpb_out[45][860],u_xpb_out[46][860],u_xpb_out[47][860],u_xpb_out[48][860],u_xpb_out[49][860],u_xpb_out[50][860],u_xpb_out[51][860],u_xpb_out[52][860],u_xpb_out[53][860],u_xpb_out[54][860],u_xpb_out[55][860],u_xpb_out[56][860],u_xpb_out[57][860],u_xpb_out[58][860],u_xpb_out[59][860],u_xpb_out[60][860],u_xpb_out[61][860],u_xpb_out[62][860],u_xpb_out[63][860],u_xpb_out[64][860],u_xpb_out[65][860],u_xpb_out[66][860],u_xpb_out[67][860],u_xpb_out[68][860],u_xpb_out[69][860],u_xpb_out[70][860],u_xpb_out[71][860],u_xpb_out[72][860],u_xpb_out[73][860],u_xpb_out[74][860],u_xpb_out[75][860],u_xpb_out[76][860],u_xpb_out[77][860],u_xpb_out[78][860],u_xpb_out[79][860],u_xpb_out[80][860],u_xpb_out[81][860],u_xpb_out[82][860],u_xpb_out[83][860],u_xpb_out[84][860],u_xpb_out[85][860],u_xpb_out[86][860],u_xpb_out[87][860],u_xpb_out[88][860],u_xpb_out[89][860],u_xpb_out[90][860],u_xpb_out[91][860],u_xpb_out[92][860],u_xpb_out[93][860],u_xpb_out[94][860],u_xpb_out[95][860],u_xpb_out[96][860],u_xpb_out[97][860],u_xpb_out[98][860],u_xpb_out[99][860],u_xpb_out[100][860],u_xpb_out[101][860],u_xpb_out[102][860],u_xpb_out[103][860],u_xpb_out[104][860],u_xpb_out[105][860]};

assign col_out_861 = {u_xpb_out[0][861],u_xpb_out[1][861],u_xpb_out[2][861],u_xpb_out[3][861],u_xpb_out[4][861],u_xpb_out[5][861],u_xpb_out[6][861],u_xpb_out[7][861],u_xpb_out[8][861],u_xpb_out[9][861],u_xpb_out[10][861],u_xpb_out[11][861],u_xpb_out[12][861],u_xpb_out[13][861],u_xpb_out[14][861],u_xpb_out[15][861],u_xpb_out[16][861],u_xpb_out[17][861],u_xpb_out[18][861],u_xpb_out[19][861],u_xpb_out[20][861],u_xpb_out[21][861],u_xpb_out[22][861],u_xpb_out[23][861],u_xpb_out[24][861],u_xpb_out[25][861],u_xpb_out[26][861],u_xpb_out[27][861],u_xpb_out[28][861],u_xpb_out[29][861],u_xpb_out[30][861],u_xpb_out[31][861],u_xpb_out[32][861],u_xpb_out[33][861],u_xpb_out[34][861],u_xpb_out[35][861],u_xpb_out[36][861],u_xpb_out[37][861],u_xpb_out[38][861],u_xpb_out[39][861],u_xpb_out[40][861],u_xpb_out[41][861],u_xpb_out[42][861],u_xpb_out[43][861],u_xpb_out[44][861],u_xpb_out[45][861],u_xpb_out[46][861],u_xpb_out[47][861],u_xpb_out[48][861],u_xpb_out[49][861],u_xpb_out[50][861],u_xpb_out[51][861],u_xpb_out[52][861],u_xpb_out[53][861],u_xpb_out[54][861],u_xpb_out[55][861],u_xpb_out[56][861],u_xpb_out[57][861],u_xpb_out[58][861],u_xpb_out[59][861],u_xpb_out[60][861],u_xpb_out[61][861],u_xpb_out[62][861],u_xpb_out[63][861],u_xpb_out[64][861],u_xpb_out[65][861],u_xpb_out[66][861],u_xpb_out[67][861],u_xpb_out[68][861],u_xpb_out[69][861],u_xpb_out[70][861],u_xpb_out[71][861],u_xpb_out[72][861],u_xpb_out[73][861],u_xpb_out[74][861],u_xpb_out[75][861],u_xpb_out[76][861],u_xpb_out[77][861],u_xpb_out[78][861],u_xpb_out[79][861],u_xpb_out[80][861],u_xpb_out[81][861],u_xpb_out[82][861],u_xpb_out[83][861],u_xpb_out[84][861],u_xpb_out[85][861],u_xpb_out[86][861],u_xpb_out[87][861],u_xpb_out[88][861],u_xpb_out[89][861],u_xpb_out[90][861],u_xpb_out[91][861],u_xpb_out[92][861],u_xpb_out[93][861],u_xpb_out[94][861],u_xpb_out[95][861],u_xpb_out[96][861],u_xpb_out[97][861],u_xpb_out[98][861],u_xpb_out[99][861],u_xpb_out[100][861],u_xpb_out[101][861],u_xpb_out[102][861],u_xpb_out[103][861],u_xpb_out[104][861],u_xpb_out[105][861]};

assign col_out_862 = {u_xpb_out[0][862],u_xpb_out[1][862],u_xpb_out[2][862],u_xpb_out[3][862],u_xpb_out[4][862],u_xpb_out[5][862],u_xpb_out[6][862],u_xpb_out[7][862],u_xpb_out[8][862],u_xpb_out[9][862],u_xpb_out[10][862],u_xpb_out[11][862],u_xpb_out[12][862],u_xpb_out[13][862],u_xpb_out[14][862],u_xpb_out[15][862],u_xpb_out[16][862],u_xpb_out[17][862],u_xpb_out[18][862],u_xpb_out[19][862],u_xpb_out[20][862],u_xpb_out[21][862],u_xpb_out[22][862],u_xpb_out[23][862],u_xpb_out[24][862],u_xpb_out[25][862],u_xpb_out[26][862],u_xpb_out[27][862],u_xpb_out[28][862],u_xpb_out[29][862],u_xpb_out[30][862],u_xpb_out[31][862],u_xpb_out[32][862],u_xpb_out[33][862],u_xpb_out[34][862],u_xpb_out[35][862],u_xpb_out[36][862],u_xpb_out[37][862],u_xpb_out[38][862],u_xpb_out[39][862],u_xpb_out[40][862],u_xpb_out[41][862],u_xpb_out[42][862],u_xpb_out[43][862],u_xpb_out[44][862],u_xpb_out[45][862],u_xpb_out[46][862],u_xpb_out[47][862],u_xpb_out[48][862],u_xpb_out[49][862],u_xpb_out[50][862],u_xpb_out[51][862],u_xpb_out[52][862],u_xpb_out[53][862],u_xpb_out[54][862],u_xpb_out[55][862],u_xpb_out[56][862],u_xpb_out[57][862],u_xpb_out[58][862],u_xpb_out[59][862],u_xpb_out[60][862],u_xpb_out[61][862],u_xpb_out[62][862],u_xpb_out[63][862],u_xpb_out[64][862],u_xpb_out[65][862],u_xpb_out[66][862],u_xpb_out[67][862],u_xpb_out[68][862],u_xpb_out[69][862],u_xpb_out[70][862],u_xpb_out[71][862],u_xpb_out[72][862],u_xpb_out[73][862],u_xpb_out[74][862],u_xpb_out[75][862],u_xpb_out[76][862],u_xpb_out[77][862],u_xpb_out[78][862],u_xpb_out[79][862],u_xpb_out[80][862],u_xpb_out[81][862],u_xpb_out[82][862],u_xpb_out[83][862],u_xpb_out[84][862],u_xpb_out[85][862],u_xpb_out[86][862],u_xpb_out[87][862],u_xpb_out[88][862],u_xpb_out[89][862],u_xpb_out[90][862],u_xpb_out[91][862],u_xpb_out[92][862],u_xpb_out[93][862],u_xpb_out[94][862],u_xpb_out[95][862],u_xpb_out[96][862],u_xpb_out[97][862],u_xpb_out[98][862],u_xpb_out[99][862],u_xpb_out[100][862],u_xpb_out[101][862],u_xpb_out[102][862],u_xpb_out[103][862],u_xpb_out[104][862],u_xpb_out[105][862]};

assign col_out_863 = {u_xpb_out[0][863],u_xpb_out[1][863],u_xpb_out[2][863],u_xpb_out[3][863],u_xpb_out[4][863],u_xpb_out[5][863],u_xpb_out[6][863],u_xpb_out[7][863],u_xpb_out[8][863],u_xpb_out[9][863],u_xpb_out[10][863],u_xpb_out[11][863],u_xpb_out[12][863],u_xpb_out[13][863],u_xpb_out[14][863],u_xpb_out[15][863],u_xpb_out[16][863],u_xpb_out[17][863],u_xpb_out[18][863],u_xpb_out[19][863],u_xpb_out[20][863],u_xpb_out[21][863],u_xpb_out[22][863],u_xpb_out[23][863],u_xpb_out[24][863],u_xpb_out[25][863],u_xpb_out[26][863],u_xpb_out[27][863],u_xpb_out[28][863],u_xpb_out[29][863],u_xpb_out[30][863],u_xpb_out[31][863],u_xpb_out[32][863],u_xpb_out[33][863],u_xpb_out[34][863],u_xpb_out[35][863],u_xpb_out[36][863],u_xpb_out[37][863],u_xpb_out[38][863],u_xpb_out[39][863],u_xpb_out[40][863],u_xpb_out[41][863],u_xpb_out[42][863],u_xpb_out[43][863],u_xpb_out[44][863],u_xpb_out[45][863],u_xpb_out[46][863],u_xpb_out[47][863],u_xpb_out[48][863],u_xpb_out[49][863],u_xpb_out[50][863],u_xpb_out[51][863],u_xpb_out[52][863],u_xpb_out[53][863],u_xpb_out[54][863],u_xpb_out[55][863],u_xpb_out[56][863],u_xpb_out[57][863],u_xpb_out[58][863],u_xpb_out[59][863],u_xpb_out[60][863],u_xpb_out[61][863],u_xpb_out[62][863],u_xpb_out[63][863],u_xpb_out[64][863],u_xpb_out[65][863],u_xpb_out[66][863],u_xpb_out[67][863],u_xpb_out[68][863],u_xpb_out[69][863],u_xpb_out[70][863],u_xpb_out[71][863],u_xpb_out[72][863],u_xpb_out[73][863],u_xpb_out[74][863],u_xpb_out[75][863],u_xpb_out[76][863],u_xpb_out[77][863],u_xpb_out[78][863],u_xpb_out[79][863],u_xpb_out[80][863],u_xpb_out[81][863],u_xpb_out[82][863],u_xpb_out[83][863],u_xpb_out[84][863],u_xpb_out[85][863],u_xpb_out[86][863],u_xpb_out[87][863],u_xpb_out[88][863],u_xpb_out[89][863],u_xpb_out[90][863],u_xpb_out[91][863],u_xpb_out[92][863],u_xpb_out[93][863],u_xpb_out[94][863],u_xpb_out[95][863],u_xpb_out[96][863],u_xpb_out[97][863],u_xpb_out[98][863],u_xpb_out[99][863],u_xpb_out[100][863],u_xpb_out[101][863],u_xpb_out[102][863],u_xpb_out[103][863],u_xpb_out[104][863],u_xpb_out[105][863]};

assign col_out_864 = {u_xpb_out[0][864],u_xpb_out[1][864],u_xpb_out[2][864],u_xpb_out[3][864],u_xpb_out[4][864],u_xpb_out[5][864],u_xpb_out[6][864],u_xpb_out[7][864],u_xpb_out[8][864],u_xpb_out[9][864],u_xpb_out[10][864],u_xpb_out[11][864],u_xpb_out[12][864],u_xpb_out[13][864],u_xpb_out[14][864],u_xpb_out[15][864],u_xpb_out[16][864],u_xpb_out[17][864],u_xpb_out[18][864],u_xpb_out[19][864],u_xpb_out[20][864],u_xpb_out[21][864],u_xpb_out[22][864],u_xpb_out[23][864],u_xpb_out[24][864],u_xpb_out[25][864],u_xpb_out[26][864],u_xpb_out[27][864],u_xpb_out[28][864],u_xpb_out[29][864],u_xpb_out[30][864],u_xpb_out[31][864],u_xpb_out[32][864],u_xpb_out[33][864],u_xpb_out[34][864],u_xpb_out[35][864],u_xpb_out[36][864],u_xpb_out[37][864],u_xpb_out[38][864],u_xpb_out[39][864],u_xpb_out[40][864],u_xpb_out[41][864],u_xpb_out[42][864],u_xpb_out[43][864],u_xpb_out[44][864],u_xpb_out[45][864],u_xpb_out[46][864],u_xpb_out[47][864],u_xpb_out[48][864],u_xpb_out[49][864],u_xpb_out[50][864],u_xpb_out[51][864],u_xpb_out[52][864],u_xpb_out[53][864],u_xpb_out[54][864],u_xpb_out[55][864],u_xpb_out[56][864],u_xpb_out[57][864],u_xpb_out[58][864],u_xpb_out[59][864],u_xpb_out[60][864],u_xpb_out[61][864],u_xpb_out[62][864],u_xpb_out[63][864],u_xpb_out[64][864],u_xpb_out[65][864],u_xpb_out[66][864],u_xpb_out[67][864],u_xpb_out[68][864],u_xpb_out[69][864],u_xpb_out[70][864],u_xpb_out[71][864],u_xpb_out[72][864],u_xpb_out[73][864],u_xpb_out[74][864],u_xpb_out[75][864],u_xpb_out[76][864],u_xpb_out[77][864],u_xpb_out[78][864],u_xpb_out[79][864],u_xpb_out[80][864],u_xpb_out[81][864],u_xpb_out[82][864],u_xpb_out[83][864],u_xpb_out[84][864],u_xpb_out[85][864],u_xpb_out[86][864],u_xpb_out[87][864],u_xpb_out[88][864],u_xpb_out[89][864],u_xpb_out[90][864],u_xpb_out[91][864],u_xpb_out[92][864],u_xpb_out[93][864],u_xpb_out[94][864],u_xpb_out[95][864],u_xpb_out[96][864],u_xpb_out[97][864],u_xpb_out[98][864],u_xpb_out[99][864],u_xpb_out[100][864],u_xpb_out[101][864],u_xpb_out[102][864],u_xpb_out[103][864],u_xpb_out[104][864],u_xpb_out[105][864]};

assign col_out_865 = {u_xpb_out[0][865],u_xpb_out[1][865],u_xpb_out[2][865],u_xpb_out[3][865],u_xpb_out[4][865],u_xpb_out[5][865],u_xpb_out[6][865],u_xpb_out[7][865],u_xpb_out[8][865],u_xpb_out[9][865],u_xpb_out[10][865],u_xpb_out[11][865],u_xpb_out[12][865],u_xpb_out[13][865],u_xpb_out[14][865],u_xpb_out[15][865],u_xpb_out[16][865],u_xpb_out[17][865],u_xpb_out[18][865],u_xpb_out[19][865],u_xpb_out[20][865],u_xpb_out[21][865],u_xpb_out[22][865],u_xpb_out[23][865],u_xpb_out[24][865],u_xpb_out[25][865],u_xpb_out[26][865],u_xpb_out[27][865],u_xpb_out[28][865],u_xpb_out[29][865],u_xpb_out[30][865],u_xpb_out[31][865],u_xpb_out[32][865],u_xpb_out[33][865],u_xpb_out[34][865],u_xpb_out[35][865],u_xpb_out[36][865],u_xpb_out[37][865],u_xpb_out[38][865],u_xpb_out[39][865],u_xpb_out[40][865],u_xpb_out[41][865],u_xpb_out[42][865],u_xpb_out[43][865],u_xpb_out[44][865],u_xpb_out[45][865],u_xpb_out[46][865],u_xpb_out[47][865],u_xpb_out[48][865],u_xpb_out[49][865],u_xpb_out[50][865],u_xpb_out[51][865],u_xpb_out[52][865],u_xpb_out[53][865],u_xpb_out[54][865],u_xpb_out[55][865],u_xpb_out[56][865],u_xpb_out[57][865],u_xpb_out[58][865],u_xpb_out[59][865],u_xpb_out[60][865],u_xpb_out[61][865],u_xpb_out[62][865],u_xpb_out[63][865],u_xpb_out[64][865],u_xpb_out[65][865],u_xpb_out[66][865],u_xpb_out[67][865],u_xpb_out[68][865],u_xpb_out[69][865],u_xpb_out[70][865],u_xpb_out[71][865],u_xpb_out[72][865],u_xpb_out[73][865],u_xpb_out[74][865],u_xpb_out[75][865],u_xpb_out[76][865],u_xpb_out[77][865],u_xpb_out[78][865],u_xpb_out[79][865],u_xpb_out[80][865],u_xpb_out[81][865],u_xpb_out[82][865],u_xpb_out[83][865],u_xpb_out[84][865],u_xpb_out[85][865],u_xpb_out[86][865],u_xpb_out[87][865],u_xpb_out[88][865],u_xpb_out[89][865],u_xpb_out[90][865],u_xpb_out[91][865],u_xpb_out[92][865],u_xpb_out[93][865],u_xpb_out[94][865],u_xpb_out[95][865],u_xpb_out[96][865],u_xpb_out[97][865],u_xpb_out[98][865],u_xpb_out[99][865],u_xpb_out[100][865],u_xpb_out[101][865],u_xpb_out[102][865],u_xpb_out[103][865],u_xpb_out[104][865],u_xpb_out[105][865]};

assign col_out_866 = {u_xpb_out[0][866],u_xpb_out[1][866],u_xpb_out[2][866],u_xpb_out[3][866],u_xpb_out[4][866],u_xpb_out[5][866],u_xpb_out[6][866],u_xpb_out[7][866],u_xpb_out[8][866],u_xpb_out[9][866],u_xpb_out[10][866],u_xpb_out[11][866],u_xpb_out[12][866],u_xpb_out[13][866],u_xpb_out[14][866],u_xpb_out[15][866],u_xpb_out[16][866],u_xpb_out[17][866],u_xpb_out[18][866],u_xpb_out[19][866],u_xpb_out[20][866],u_xpb_out[21][866],u_xpb_out[22][866],u_xpb_out[23][866],u_xpb_out[24][866],u_xpb_out[25][866],u_xpb_out[26][866],u_xpb_out[27][866],u_xpb_out[28][866],u_xpb_out[29][866],u_xpb_out[30][866],u_xpb_out[31][866],u_xpb_out[32][866],u_xpb_out[33][866],u_xpb_out[34][866],u_xpb_out[35][866],u_xpb_out[36][866],u_xpb_out[37][866],u_xpb_out[38][866],u_xpb_out[39][866],u_xpb_out[40][866],u_xpb_out[41][866],u_xpb_out[42][866],u_xpb_out[43][866],u_xpb_out[44][866],u_xpb_out[45][866],u_xpb_out[46][866],u_xpb_out[47][866],u_xpb_out[48][866],u_xpb_out[49][866],u_xpb_out[50][866],u_xpb_out[51][866],u_xpb_out[52][866],u_xpb_out[53][866],u_xpb_out[54][866],u_xpb_out[55][866],u_xpb_out[56][866],u_xpb_out[57][866],u_xpb_out[58][866],u_xpb_out[59][866],u_xpb_out[60][866],u_xpb_out[61][866],u_xpb_out[62][866],u_xpb_out[63][866],u_xpb_out[64][866],u_xpb_out[65][866],u_xpb_out[66][866],u_xpb_out[67][866],u_xpb_out[68][866],u_xpb_out[69][866],u_xpb_out[70][866],u_xpb_out[71][866],u_xpb_out[72][866],u_xpb_out[73][866],u_xpb_out[74][866],u_xpb_out[75][866],u_xpb_out[76][866],u_xpb_out[77][866],u_xpb_out[78][866],u_xpb_out[79][866],u_xpb_out[80][866],u_xpb_out[81][866],u_xpb_out[82][866],u_xpb_out[83][866],u_xpb_out[84][866],u_xpb_out[85][866],u_xpb_out[86][866],u_xpb_out[87][866],u_xpb_out[88][866],u_xpb_out[89][866],u_xpb_out[90][866],u_xpb_out[91][866],u_xpb_out[92][866],u_xpb_out[93][866],u_xpb_out[94][866],u_xpb_out[95][866],u_xpb_out[96][866],u_xpb_out[97][866],u_xpb_out[98][866],u_xpb_out[99][866],u_xpb_out[100][866],u_xpb_out[101][866],u_xpb_out[102][866],u_xpb_out[103][866],u_xpb_out[104][866],u_xpb_out[105][866]};

assign col_out_867 = {u_xpb_out[0][867],u_xpb_out[1][867],u_xpb_out[2][867],u_xpb_out[3][867],u_xpb_out[4][867],u_xpb_out[5][867],u_xpb_out[6][867],u_xpb_out[7][867],u_xpb_out[8][867],u_xpb_out[9][867],u_xpb_out[10][867],u_xpb_out[11][867],u_xpb_out[12][867],u_xpb_out[13][867],u_xpb_out[14][867],u_xpb_out[15][867],u_xpb_out[16][867],u_xpb_out[17][867],u_xpb_out[18][867],u_xpb_out[19][867],u_xpb_out[20][867],u_xpb_out[21][867],u_xpb_out[22][867],u_xpb_out[23][867],u_xpb_out[24][867],u_xpb_out[25][867],u_xpb_out[26][867],u_xpb_out[27][867],u_xpb_out[28][867],u_xpb_out[29][867],u_xpb_out[30][867],u_xpb_out[31][867],u_xpb_out[32][867],u_xpb_out[33][867],u_xpb_out[34][867],u_xpb_out[35][867],u_xpb_out[36][867],u_xpb_out[37][867],u_xpb_out[38][867],u_xpb_out[39][867],u_xpb_out[40][867],u_xpb_out[41][867],u_xpb_out[42][867],u_xpb_out[43][867],u_xpb_out[44][867],u_xpb_out[45][867],u_xpb_out[46][867],u_xpb_out[47][867],u_xpb_out[48][867],u_xpb_out[49][867],u_xpb_out[50][867],u_xpb_out[51][867],u_xpb_out[52][867],u_xpb_out[53][867],u_xpb_out[54][867],u_xpb_out[55][867],u_xpb_out[56][867],u_xpb_out[57][867],u_xpb_out[58][867],u_xpb_out[59][867],u_xpb_out[60][867],u_xpb_out[61][867],u_xpb_out[62][867],u_xpb_out[63][867],u_xpb_out[64][867],u_xpb_out[65][867],u_xpb_out[66][867],u_xpb_out[67][867],u_xpb_out[68][867],u_xpb_out[69][867],u_xpb_out[70][867],u_xpb_out[71][867],u_xpb_out[72][867],u_xpb_out[73][867],u_xpb_out[74][867],u_xpb_out[75][867],u_xpb_out[76][867],u_xpb_out[77][867],u_xpb_out[78][867],u_xpb_out[79][867],u_xpb_out[80][867],u_xpb_out[81][867],u_xpb_out[82][867],u_xpb_out[83][867],u_xpb_out[84][867],u_xpb_out[85][867],u_xpb_out[86][867],u_xpb_out[87][867],u_xpb_out[88][867],u_xpb_out[89][867],u_xpb_out[90][867],u_xpb_out[91][867],u_xpb_out[92][867],u_xpb_out[93][867],u_xpb_out[94][867],u_xpb_out[95][867],u_xpb_out[96][867],u_xpb_out[97][867],u_xpb_out[98][867],u_xpb_out[99][867],u_xpb_out[100][867],u_xpb_out[101][867],u_xpb_out[102][867],u_xpb_out[103][867],u_xpb_out[104][867],u_xpb_out[105][867]};

assign col_out_868 = {u_xpb_out[0][868],u_xpb_out[1][868],u_xpb_out[2][868],u_xpb_out[3][868],u_xpb_out[4][868],u_xpb_out[5][868],u_xpb_out[6][868],u_xpb_out[7][868],u_xpb_out[8][868],u_xpb_out[9][868],u_xpb_out[10][868],u_xpb_out[11][868],u_xpb_out[12][868],u_xpb_out[13][868],u_xpb_out[14][868],u_xpb_out[15][868],u_xpb_out[16][868],u_xpb_out[17][868],u_xpb_out[18][868],u_xpb_out[19][868],u_xpb_out[20][868],u_xpb_out[21][868],u_xpb_out[22][868],u_xpb_out[23][868],u_xpb_out[24][868],u_xpb_out[25][868],u_xpb_out[26][868],u_xpb_out[27][868],u_xpb_out[28][868],u_xpb_out[29][868],u_xpb_out[30][868],u_xpb_out[31][868],u_xpb_out[32][868],u_xpb_out[33][868],u_xpb_out[34][868],u_xpb_out[35][868],u_xpb_out[36][868],u_xpb_out[37][868],u_xpb_out[38][868],u_xpb_out[39][868],u_xpb_out[40][868],u_xpb_out[41][868],u_xpb_out[42][868],u_xpb_out[43][868],u_xpb_out[44][868],u_xpb_out[45][868],u_xpb_out[46][868],u_xpb_out[47][868],u_xpb_out[48][868],u_xpb_out[49][868],u_xpb_out[50][868],u_xpb_out[51][868],u_xpb_out[52][868],u_xpb_out[53][868],u_xpb_out[54][868],u_xpb_out[55][868],u_xpb_out[56][868],u_xpb_out[57][868],u_xpb_out[58][868],u_xpb_out[59][868],u_xpb_out[60][868],u_xpb_out[61][868],u_xpb_out[62][868],u_xpb_out[63][868],u_xpb_out[64][868],u_xpb_out[65][868],u_xpb_out[66][868],u_xpb_out[67][868],u_xpb_out[68][868],u_xpb_out[69][868],u_xpb_out[70][868],u_xpb_out[71][868],u_xpb_out[72][868],u_xpb_out[73][868],u_xpb_out[74][868],u_xpb_out[75][868],u_xpb_out[76][868],u_xpb_out[77][868],u_xpb_out[78][868],u_xpb_out[79][868],u_xpb_out[80][868],u_xpb_out[81][868],u_xpb_out[82][868],u_xpb_out[83][868],u_xpb_out[84][868],u_xpb_out[85][868],u_xpb_out[86][868],u_xpb_out[87][868],u_xpb_out[88][868],u_xpb_out[89][868],u_xpb_out[90][868],u_xpb_out[91][868],u_xpb_out[92][868],u_xpb_out[93][868],u_xpb_out[94][868],u_xpb_out[95][868],u_xpb_out[96][868],u_xpb_out[97][868],u_xpb_out[98][868],u_xpb_out[99][868],u_xpb_out[100][868],u_xpb_out[101][868],u_xpb_out[102][868],u_xpb_out[103][868],u_xpb_out[104][868],u_xpb_out[105][868]};

assign col_out_869 = {u_xpb_out[0][869],u_xpb_out[1][869],u_xpb_out[2][869],u_xpb_out[3][869],u_xpb_out[4][869],u_xpb_out[5][869],u_xpb_out[6][869],u_xpb_out[7][869],u_xpb_out[8][869],u_xpb_out[9][869],u_xpb_out[10][869],u_xpb_out[11][869],u_xpb_out[12][869],u_xpb_out[13][869],u_xpb_out[14][869],u_xpb_out[15][869],u_xpb_out[16][869],u_xpb_out[17][869],u_xpb_out[18][869],u_xpb_out[19][869],u_xpb_out[20][869],u_xpb_out[21][869],u_xpb_out[22][869],u_xpb_out[23][869],u_xpb_out[24][869],u_xpb_out[25][869],u_xpb_out[26][869],u_xpb_out[27][869],u_xpb_out[28][869],u_xpb_out[29][869],u_xpb_out[30][869],u_xpb_out[31][869],u_xpb_out[32][869],u_xpb_out[33][869],u_xpb_out[34][869],u_xpb_out[35][869],u_xpb_out[36][869],u_xpb_out[37][869],u_xpb_out[38][869],u_xpb_out[39][869],u_xpb_out[40][869],u_xpb_out[41][869],u_xpb_out[42][869],u_xpb_out[43][869],u_xpb_out[44][869],u_xpb_out[45][869],u_xpb_out[46][869],u_xpb_out[47][869],u_xpb_out[48][869],u_xpb_out[49][869],u_xpb_out[50][869],u_xpb_out[51][869],u_xpb_out[52][869],u_xpb_out[53][869],u_xpb_out[54][869],u_xpb_out[55][869],u_xpb_out[56][869],u_xpb_out[57][869],u_xpb_out[58][869],u_xpb_out[59][869],u_xpb_out[60][869],u_xpb_out[61][869],u_xpb_out[62][869],u_xpb_out[63][869],u_xpb_out[64][869],u_xpb_out[65][869],u_xpb_out[66][869],u_xpb_out[67][869],u_xpb_out[68][869],u_xpb_out[69][869],u_xpb_out[70][869],u_xpb_out[71][869],u_xpb_out[72][869],u_xpb_out[73][869],u_xpb_out[74][869],u_xpb_out[75][869],u_xpb_out[76][869],u_xpb_out[77][869],u_xpb_out[78][869],u_xpb_out[79][869],u_xpb_out[80][869],u_xpb_out[81][869],u_xpb_out[82][869],u_xpb_out[83][869],u_xpb_out[84][869],u_xpb_out[85][869],u_xpb_out[86][869],u_xpb_out[87][869],u_xpb_out[88][869],u_xpb_out[89][869],u_xpb_out[90][869],u_xpb_out[91][869],u_xpb_out[92][869],u_xpb_out[93][869],u_xpb_out[94][869],u_xpb_out[95][869],u_xpb_out[96][869],u_xpb_out[97][869],u_xpb_out[98][869],u_xpb_out[99][869],u_xpb_out[100][869],u_xpb_out[101][869],u_xpb_out[102][869],u_xpb_out[103][869],u_xpb_out[104][869],u_xpb_out[105][869]};

assign col_out_870 = {u_xpb_out[0][870],u_xpb_out[1][870],u_xpb_out[2][870],u_xpb_out[3][870],u_xpb_out[4][870],u_xpb_out[5][870],u_xpb_out[6][870],u_xpb_out[7][870],u_xpb_out[8][870],u_xpb_out[9][870],u_xpb_out[10][870],u_xpb_out[11][870],u_xpb_out[12][870],u_xpb_out[13][870],u_xpb_out[14][870],u_xpb_out[15][870],u_xpb_out[16][870],u_xpb_out[17][870],u_xpb_out[18][870],u_xpb_out[19][870],u_xpb_out[20][870],u_xpb_out[21][870],u_xpb_out[22][870],u_xpb_out[23][870],u_xpb_out[24][870],u_xpb_out[25][870],u_xpb_out[26][870],u_xpb_out[27][870],u_xpb_out[28][870],u_xpb_out[29][870],u_xpb_out[30][870],u_xpb_out[31][870],u_xpb_out[32][870],u_xpb_out[33][870],u_xpb_out[34][870],u_xpb_out[35][870],u_xpb_out[36][870],u_xpb_out[37][870],u_xpb_out[38][870],u_xpb_out[39][870],u_xpb_out[40][870],u_xpb_out[41][870],u_xpb_out[42][870],u_xpb_out[43][870],u_xpb_out[44][870],u_xpb_out[45][870],u_xpb_out[46][870],u_xpb_out[47][870],u_xpb_out[48][870],u_xpb_out[49][870],u_xpb_out[50][870],u_xpb_out[51][870],u_xpb_out[52][870],u_xpb_out[53][870],u_xpb_out[54][870],u_xpb_out[55][870],u_xpb_out[56][870],u_xpb_out[57][870],u_xpb_out[58][870],u_xpb_out[59][870],u_xpb_out[60][870],u_xpb_out[61][870],u_xpb_out[62][870],u_xpb_out[63][870],u_xpb_out[64][870],u_xpb_out[65][870],u_xpb_out[66][870],u_xpb_out[67][870],u_xpb_out[68][870],u_xpb_out[69][870],u_xpb_out[70][870],u_xpb_out[71][870],u_xpb_out[72][870],u_xpb_out[73][870],u_xpb_out[74][870],u_xpb_out[75][870],u_xpb_out[76][870],u_xpb_out[77][870],u_xpb_out[78][870],u_xpb_out[79][870],u_xpb_out[80][870],u_xpb_out[81][870],u_xpb_out[82][870],u_xpb_out[83][870],u_xpb_out[84][870],u_xpb_out[85][870],u_xpb_out[86][870],u_xpb_out[87][870],u_xpb_out[88][870],u_xpb_out[89][870],u_xpb_out[90][870],u_xpb_out[91][870],u_xpb_out[92][870],u_xpb_out[93][870],u_xpb_out[94][870],u_xpb_out[95][870],u_xpb_out[96][870],u_xpb_out[97][870],u_xpb_out[98][870],u_xpb_out[99][870],u_xpb_out[100][870],u_xpb_out[101][870],u_xpb_out[102][870],u_xpb_out[103][870],u_xpb_out[104][870],u_xpb_out[105][870]};

assign col_out_871 = {u_xpb_out[0][871],u_xpb_out[1][871],u_xpb_out[2][871],u_xpb_out[3][871],u_xpb_out[4][871],u_xpb_out[5][871],u_xpb_out[6][871],u_xpb_out[7][871],u_xpb_out[8][871],u_xpb_out[9][871],u_xpb_out[10][871],u_xpb_out[11][871],u_xpb_out[12][871],u_xpb_out[13][871],u_xpb_out[14][871],u_xpb_out[15][871],u_xpb_out[16][871],u_xpb_out[17][871],u_xpb_out[18][871],u_xpb_out[19][871],u_xpb_out[20][871],u_xpb_out[21][871],u_xpb_out[22][871],u_xpb_out[23][871],u_xpb_out[24][871],u_xpb_out[25][871],u_xpb_out[26][871],u_xpb_out[27][871],u_xpb_out[28][871],u_xpb_out[29][871],u_xpb_out[30][871],u_xpb_out[31][871],u_xpb_out[32][871],u_xpb_out[33][871],u_xpb_out[34][871],u_xpb_out[35][871],u_xpb_out[36][871],u_xpb_out[37][871],u_xpb_out[38][871],u_xpb_out[39][871],u_xpb_out[40][871],u_xpb_out[41][871],u_xpb_out[42][871],u_xpb_out[43][871],u_xpb_out[44][871],u_xpb_out[45][871],u_xpb_out[46][871],u_xpb_out[47][871],u_xpb_out[48][871],u_xpb_out[49][871],u_xpb_out[50][871],u_xpb_out[51][871],u_xpb_out[52][871],u_xpb_out[53][871],u_xpb_out[54][871],u_xpb_out[55][871],u_xpb_out[56][871],u_xpb_out[57][871],u_xpb_out[58][871],u_xpb_out[59][871],u_xpb_out[60][871],u_xpb_out[61][871],u_xpb_out[62][871],u_xpb_out[63][871],u_xpb_out[64][871],u_xpb_out[65][871],u_xpb_out[66][871],u_xpb_out[67][871],u_xpb_out[68][871],u_xpb_out[69][871],u_xpb_out[70][871],u_xpb_out[71][871],u_xpb_out[72][871],u_xpb_out[73][871],u_xpb_out[74][871],u_xpb_out[75][871],u_xpb_out[76][871],u_xpb_out[77][871],u_xpb_out[78][871],u_xpb_out[79][871],u_xpb_out[80][871],u_xpb_out[81][871],u_xpb_out[82][871],u_xpb_out[83][871],u_xpb_out[84][871],u_xpb_out[85][871],u_xpb_out[86][871],u_xpb_out[87][871],u_xpb_out[88][871],u_xpb_out[89][871],u_xpb_out[90][871],u_xpb_out[91][871],u_xpb_out[92][871],u_xpb_out[93][871],u_xpb_out[94][871],u_xpb_out[95][871],u_xpb_out[96][871],u_xpb_out[97][871],u_xpb_out[98][871],u_xpb_out[99][871],u_xpb_out[100][871],u_xpb_out[101][871],u_xpb_out[102][871],u_xpb_out[103][871],u_xpb_out[104][871],u_xpb_out[105][871]};

assign col_out_872 = {u_xpb_out[0][872],u_xpb_out[1][872],u_xpb_out[2][872],u_xpb_out[3][872],u_xpb_out[4][872],u_xpb_out[5][872],u_xpb_out[6][872],u_xpb_out[7][872],u_xpb_out[8][872],u_xpb_out[9][872],u_xpb_out[10][872],u_xpb_out[11][872],u_xpb_out[12][872],u_xpb_out[13][872],u_xpb_out[14][872],u_xpb_out[15][872],u_xpb_out[16][872],u_xpb_out[17][872],u_xpb_out[18][872],u_xpb_out[19][872],u_xpb_out[20][872],u_xpb_out[21][872],u_xpb_out[22][872],u_xpb_out[23][872],u_xpb_out[24][872],u_xpb_out[25][872],u_xpb_out[26][872],u_xpb_out[27][872],u_xpb_out[28][872],u_xpb_out[29][872],u_xpb_out[30][872],u_xpb_out[31][872],u_xpb_out[32][872],u_xpb_out[33][872],u_xpb_out[34][872],u_xpb_out[35][872],u_xpb_out[36][872],u_xpb_out[37][872],u_xpb_out[38][872],u_xpb_out[39][872],u_xpb_out[40][872],u_xpb_out[41][872],u_xpb_out[42][872],u_xpb_out[43][872],u_xpb_out[44][872],u_xpb_out[45][872],u_xpb_out[46][872],u_xpb_out[47][872],u_xpb_out[48][872],u_xpb_out[49][872],u_xpb_out[50][872],u_xpb_out[51][872],u_xpb_out[52][872],u_xpb_out[53][872],u_xpb_out[54][872],u_xpb_out[55][872],u_xpb_out[56][872],u_xpb_out[57][872],u_xpb_out[58][872],u_xpb_out[59][872],u_xpb_out[60][872],u_xpb_out[61][872],u_xpb_out[62][872],u_xpb_out[63][872],u_xpb_out[64][872],u_xpb_out[65][872],u_xpb_out[66][872],u_xpb_out[67][872],u_xpb_out[68][872],u_xpb_out[69][872],u_xpb_out[70][872],u_xpb_out[71][872],u_xpb_out[72][872],u_xpb_out[73][872],u_xpb_out[74][872],u_xpb_out[75][872],u_xpb_out[76][872],u_xpb_out[77][872],u_xpb_out[78][872],u_xpb_out[79][872],u_xpb_out[80][872],u_xpb_out[81][872],u_xpb_out[82][872],u_xpb_out[83][872],u_xpb_out[84][872],u_xpb_out[85][872],u_xpb_out[86][872],u_xpb_out[87][872],u_xpb_out[88][872],u_xpb_out[89][872],u_xpb_out[90][872],u_xpb_out[91][872],u_xpb_out[92][872],u_xpb_out[93][872],u_xpb_out[94][872],u_xpb_out[95][872],u_xpb_out[96][872],u_xpb_out[97][872],u_xpb_out[98][872],u_xpb_out[99][872],u_xpb_out[100][872],u_xpb_out[101][872],u_xpb_out[102][872],u_xpb_out[103][872],u_xpb_out[104][872],u_xpb_out[105][872]};

assign col_out_873 = {u_xpb_out[0][873],u_xpb_out[1][873],u_xpb_out[2][873],u_xpb_out[3][873],u_xpb_out[4][873],u_xpb_out[5][873],u_xpb_out[6][873],u_xpb_out[7][873],u_xpb_out[8][873],u_xpb_out[9][873],u_xpb_out[10][873],u_xpb_out[11][873],u_xpb_out[12][873],u_xpb_out[13][873],u_xpb_out[14][873],u_xpb_out[15][873],u_xpb_out[16][873],u_xpb_out[17][873],u_xpb_out[18][873],u_xpb_out[19][873],u_xpb_out[20][873],u_xpb_out[21][873],u_xpb_out[22][873],u_xpb_out[23][873],u_xpb_out[24][873],u_xpb_out[25][873],u_xpb_out[26][873],u_xpb_out[27][873],u_xpb_out[28][873],u_xpb_out[29][873],u_xpb_out[30][873],u_xpb_out[31][873],u_xpb_out[32][873],u_xpb_out[33][873],u_xpb_out[34][873],u_xpb_out[35][873],u_xpb_out[36][873],u_xpb_out[37][873],u_xpb_out[38][873],u_xpb_out[39][873],u_xpb_out[40][873],u_xpb_out[41][873],u_xpb_out[42][873],u_xpb_out[43][873],u_xpb_out[44][873],u_xpb_out[45][873],u_xpb_out[46][873],u_xpb_out[47][873],u_xpb_out[48][873],u_xpb_out[49][873],u_xpb_out[50][873],u_xpb_out[51][873],u_xpb_out[52][873],u_xpb_out[53][873],u_xpb_out[54][873],u_xpb_out[55][873],u_xpb_out[56][873],u_xpb_out[57][873],u_xpb_out[58][873],u_xpb_out[59][873],u_xpb_out[60][873],u_xpb_out[61][873],u_xpb_out[62][873],u_xpb_out[63][873],u_xpb_out[64][873],u_xpb_out[65][873],u_xpb_out[66][873],u_xpb_out[67][873],u_xpb_out[68][873],u_xpb_out[69][873],u_xpb_out[70][873],u_xpb_out[71][873],u_xpb_out[72][873],u_xpb_out[73][873],u_xpb_out[74][873],u_xpb_out[75][873],u_xpb_out[76][873],u_xpb_out[77][873],u_xpb_out[78][873],u_xpb_out[79][873],u_xpb_out[80][873],u_xpb_out[81][873],u_xpb_out[82][873],u_xpb_out[83][873],u_xpb_out[84][873],u_xpb_out[85][873],u_xpb_out[86][873],u_xpb_out[87][873],u_xpb_out[88][873],u_xpb_out[89][873],u_xpb_out[90][873],u_xpb_out[91][873],u_xpb_out[92][873],u_xpb_out[93][873],u_xpb_out[94][873],u_xpb_out[95][873],u_xpb_out[96][873],u_xpb_out[97][873],u_xpb_out[98][873],u_xpb_out[99][873],u_xpb_out[100][873],u_xpb_out[101][873],u_xpb_out[102][873],u_xpb_out[103][873],u_xpb_out[104][873],u_xpb_out[105][873]};

assign col_out_874 = {u_xpb_out[0][874],u_xpb_out[1][874],u_xpb_out[2][874],u_xpb_out[3][874],u_xpb_out[4][874],u_xpb_out[5][874],u_xpb_out[6][874],u_xpb_out[7][874],u_xpb_out[8][874],u_xpb_out[9][874],u_xpb_out[10][874],u_xpb_out[11][874],u_xpb_out[12][874],u_xpb_out[13][874],u_xpb_out[14][874],u_xpb_out[15][874],u_xpb_out[16][874],u_xpb_out[17][874],u_xpb_out[18][874],u_xpb_out[19][874],u_xpb_out[20][874],u_xpb_out[21][874],u_xpb_out[22][874],u_xpb_out[23][874],u_xpb_out[24][874],u_xpb_out[25][874],u_xpb_out[26][874],u_xpb_out[27][874],u_xpb_out[28][874],u_xpb_out[29][874],u_xpb_out[30][874],u_xpb_out[31][874],u_xpb_out[32][874],u_xpb_out[33][874],u_xpb_out[34][874],u_xpb_out[35][874],u_xpb_out[36][874],u_xpb_out[37][874],u_xpb_out[38][874],u_xpb_out[39][874],u_xpb_out[40][874],u_xpb_out[41][874],u_xpb_out[42][874],u_xpb_out[43][874],u_xpb_out[44][874],u_xpb_out[45][874],u_xpb_out[46][874],u_xpb_out[47][874],u_xpb_out[48][874],u_xpb_out[49][874],u_xpb_out[50][874],u_xpb_out[51][874],u_xpb_out[52][874],u_xpb_out[53][874],u_xpb_out[54][874],u_xpb_out[55][874],u_xpb_out[56][874],u_xpb_out[57][874],u_xpb_out[58][874],u_xpb_out[59][874],u_xpb_out[60][874],u_xpb_out[61][874],u_xpb_out[62][874],u_xpb_out[63][874],u_xpb_out[64][874],u_xpb_out[65][874],u_xpb_out[66][874],u_xpb_out[67][874],u_xpb_out[68][874],u_xpb_out[69][874],u_xpb_out[70][874],u_xpb_out[71][874],u_xpb_out[72][874],u_xpb_out[73][874],u_xpb_out[74][874],u_xpb_out[75][874],u_xpb_out[76][874],u_xpb_out[77][874],u_xpb_out[78][874],u_xpb_out[79][874],u_xpb_out[80][874],u_xpb_out[81][874],u_xpb_out[82][874],u_xpb_out[83][874],u_xpb_out[84][874],u_xpb_out[85][874],u_xpb_out[86][874],u_xpb_out[87][874],u_xpb_out[88][874],u_xpb_out[89][874],u_xpb_out[90][874],u_xpb_out[91][874],u_xpb_out[92][874],u_xpb_out[93][874],u_xpb_out[94][874],u_xpb_out[95][874],u_xpb_out[96][874],u_xpb_out[97][874],u_xpb_out[98][874],u_xpb_out[99][874],u_xpb_out[100][874],u_xpb_out[101][874],u_xpb_out[102][874],u_xpb_out[103][874],u_xpb_out[104][874],u_xpb_out[105][874]};

assign col_out_875 = {u_xpb_out[0][875],u_xpb_out[1][875],u_xpb_out[2][875],u_xpb_out[3][875],u_xpb_out[4][875],u_xpb_out[5][875],u_xpb_out[6][875],u_xpb_out[7][875],u_xpb_out[8][875],u_xpb_out[9][875],u_xpb_out[10][875],u_xpb_out[11][875],u_xpb_out[12][875],u_xpb_out[13][875],u_xpb_out[14][875],u_xpb_out[15][875],u_xpb_out[16][875],u_xpb_out[17][875],u_xpb_out[18][875],u_xpb_out[19][875],u_xpb_out[20][875],u_xpb_out[21][875],u_xpb_out[22][875],u_xpb_out[23][875],u_xpb_out[24][875],u_xpb_out[25][875],u_xpb_out[26][875],u_xpb_out[27][875],u_xpb_out[28][875],u_xpb_out[29][875],u_xpb_out[30][875],u_xpb_out[31][875],u_xpb_out[32][875],u_xpb_out[33][875],u_xpb_out[34][875],u_xpb_out[35][875],u_xpb_out[36][875],u_xpb_out[37][875],u_xpb_out[38][875],u_xpb_out[39][875],u_xpb_out[40][875],u_xpb_out[41][875],u_xpb_out[42][875],u_xpb_out[43][875],u_xpb_out[44][875],u_xpb_out[45][875],u_xpb_out[46][875],u_xpb_out[47][875],u_xpb_out[48][875],u_xpb_out[49][875],u_xpb_out[50][875],u_xpb_out[51][875],u_xpb_out[52][875],u_xpb_out[53][875],u_xpb_out[54][875],u_xpb_out[55][875],u_xpb_out[56][875],u_xpb_out[57][875],u_xpb_out[58][875],u_xpb_out[59][875],u_xpb_out[60][875],u_xpb_out[61][875],u_xpb_out[62][875],u_xpb_out[63][875],u_xpb_out[64][875],u_xpb_out[65][875],u_xpb_out[66][875],u_xpb_out[67][875],u_xpb_out[68][875],u_xpb_out[69][875],u_xpb_out[70][875],u_xpb_out[71][875],u_xpb_out[72][875],u_xpb_out[73][875],u_xpb_out[74][875],u_xpb_out[75][875],u_xpb_out[76][875],u_xpb_out[77][875],u_xpb_out[78][875],u_xpb_out[79][875],u_xpb_out[80][875],u_xpb_out[81][875],u_xpb_out[82][875],u_xpb_out[83][875],u_xpb_out[84][875],u_xpb_out[85][875],u_xpb_out[86][875],u_xpb_out[87][875],u_xpb_out[88][875],u_xpb_out[89][875],u_xpb_out[90][875],u_xpb_out[91][875],u_xpb_out[92][875],u_xpb_out[93][875],u_xpb_out[94][875],u_xpb_out[95][875],u_xpb_out[96][875],u_xpb_out[97][875],u_xpb_out[98][875],u_xpb_out[99][875],u_xpb_out[100][875],u_xpb_out[101][875],u_xpb_out[102][875],u_xpb_out[103][875],u_xpb_out[104][875],u_xpb_out[105][875]};

assign col_out_876 = {u_xpb_out[0][876],u_xpb_out[1][876],u_xpb_out[2][876],u_xpb_out[3][876],u_xpb_out[4][876],u_xpb_out[5][876],u_xpb_out[6][876],u_xpb_out[7][876],u_xpb_out[8][876],u_xpb_out[9][876],u_xpb_out[10][876],u_xpb_out[11][876],u_xpb_out[12][876],u_xpb_out[13][876],u_xpb_out[14][876],u_xpb_out[15][876],u_xpb_out[16][876],u_xpb_out[17][876],u_xpb_out[18][876],u_xpb_out[19][876],u_xpb_out[20][876],u_xpb_out[21][876],u_xpb_out[22][876],u_xpb_out[23][876],u_xpb_out[24][876],u_xpb_out[25][876],u_xpb_out[26][876],u_xpb_out[27][876],u_xpb_out[28][876],u_xpb_out[29][876],u_xpb_out[30][876],u_xpb_out[31][876],u_xpb_out[32][876],u_xpb_out[33][876],u_xpb_out[34][876],u_xpb_out[35][876],u_xpb_out[36][876],u_xpb_out[37][876],u_xpb_out[38][876],u_xpb_out[39][876],u_xpb_out[40][876],u_xpb_out[41][876],u_xpb_out[42][876],u_xpb_out[43][876],u_xpb_out[44][876],u_xpb_out[45][876],u_xpb_out[46][876],u_xpb_out[47][876],u_xpb_out[48][876],u_xpb_out[49][876],u_xpb_out[50][876],u_xpb_out[51][876],u_xpb_out[52][876],u_xpb_out[53][876],u_xpb_out[54][876],u_xpb_out[55][876],u_xpb_out[56][876],u_xpb_out[57][876],u_xpb_out[58][876],u_xpb_out[59][876],u_xpb_out[60][876],u_xpb_out[61][876],u_xpb_out[62][876],u_xpb_out[63][876],u_xpb_out[64][876],u_xpb_out[65][876],u_xpb_out[66][876],u_xpb_out[67][876],u_xpb_out[68][876],u_xpb_out[69][876],u_xpb_out[70][876],u_xpb_out[71][876],u_xpb_out[72][876],u_xpb_out[73][876],u_xpb_out[74][876],u_xpb_out[75][876],u_xpb_out[76][876],u_xpb_out[77][876],u_xpb_out[78][876],u_xpb_out[79][876],u_xpb_out[80][876],u_xpb_out[81][876],u_xpb_out[82][876],u_xpb_out[83][876],u_xpb_out[84][876],u_xpb_out[85][876],u_xpb_out[86][876],u_xpb_out[87][876],u_xpb_out[88][876],u_xpb_out[89][876],u_xpb_out[90][876],u_xpb_out[91][876],u_xpb_out[92][876],u_xpb_out[93][876],u_xpb_out[94][876],u_xpb_out[95][876],u_xpb_out[96][876],u_xpb_out[97][876],u_xpb_out[98][876],u_xpb_out[99][876],u_xpb_out[100][876],u_xpb_out[101][876],u_xpb_out[102][876],u_xpb_out[103][876],u_xpb_out[104][876],u_xpb_out[105][876]};

assign col_out_877 = {u_xpb_out[0][877],u_xpb_out[1][877],u_xpb_out[2][877],u_xpb_out[3][877],u_xpb_out[4][877],u_xpb_out[5][877],u_xpb_out[6][877],u_xpb_out[7][877],u_xpb_out[8][877],u_xpb_out[9][877],u_xpb_out[10][877],u_xpb_out[11][877],u_xpb_out[12][877],u_xpb_out[13][877],u_xpb_out[14][877],u_xpb_out[15][877],u_xpb_out[16][877],u_xpb_out[17][877],u_xpb_out[18][877],u_xpb_out[19][877],u_xpb_out[20][877],u_xpb_out[21][877],u_xpb_out[22][877],u_xpb_out[23][877],u_xpb_out[24][877],u_xpb_out[25][877],u_xpb_out[26][877],u_xpb_out[27][877],u_xpb_out[28][877],u_xpb_out[29][877],u_xpb_out[30][877],u_xpb_out[31][877],u_xpb_out[32][877],u_xpb_out[33][877],u_xpb_out[34][877],u_xpb_out[35][877],u_xpb_out[36][877],u_xpb_out[37][877],u_xpb_out[38][877],u_xpb_out[39][877],u_xpb_out[40][877],u_xpb_out[41][877],u_xpb_out[42][877],u_xpb_out[43][877],u_xpb_out[44][877],u_xpb_out[45][877],u_xpb_out[46][877],u_xpb_out[47][877],u_xpb_out[48][877],u_xpb_out[49][877],u_xpb_out[50][877],u_xpb_out[51][877],u_xpb_out[52][877],u_xpb_out[53][877],u_xpb_out[54][877],u_xpb_out[55][877],u_xpb_out[56][877],u_xpb_out[57][877],u_xpb_out[58][877],u_xpb_out[59][877],u_xpb_out[60][877],u_xpb_out[61][877],u_xpb_out[62][877],u_xpb_out[63][877],u_xpb_out[64][877],u_xpb_out[65][877],u_xpb_out[66][877],u_xpb_out[67][877],u_xpb_out[68][877],u_xpb_out[69][877],u_xpb_out[70][877],u_xpb_out[71][877],u_xpb_out[72][877],u_xpb_out[73][877],u_xpb_out[74][877],u_xpb_out[75][877],u_xpb_out[76][877],u_xpb_out[77][877],u_xpb_out[78][877],u_xpb_out[79][877],u_xpb_out[80][877],u_xpb_out[81][877],u_xpb_out[82][877],u_xpb_out[83][877],u_xpb_out[84][877],u_xpb_out[85][877],u_xpb_out[86][877],u_xpb_out[87][877],u_xpb_out[88][877],u_xpb_out[89][877],u_xpb_out[90][877],u_xpb_out[91][877],u_xpb_out[92][877],u_xpb_out[93][877],u_xpb_out[94][877],u_xpb_out[95][877],u_xpb_out[96][877],u_xpb_out[97][877],u_xpb_out[98][877],u_xpb_out[99][877],u_xpb_out[100][877],u_xpb_out[101][877],u_xpb_out[102][877],u_xpb_out[103][877],u_xpb_out[104][877],u_xpb_out[105][877]};

assign col_out_878 = {u_xpb_out[0][878],u_xpb_out[1][878],u_xpb_out[2][878],u_xpb_out[3][878],u_xpb_out[4][878],u_xpb_out[5][878],u_xpb_out[6][878],u_xpb_out[7][878],u_xpb_out[8][878],u_xpb_out[9][878],u_xpb_out[10][878],u_xpb_out[11][878],u_xpb_out[12][878],u_xpb_out[13][878],u_xpb_out[14][878],u_xpb_out[15][878],u_xpb_out[16][878],u_xpb_out[17][878],u_xpb_out[18][878],u_xpb_out[19][878],u_xpb_out[20][878],u_xpb_out[21][878],u_xpb_out[22][878],u_xpb_out[23][878],u_xpb_out[24][878],u_xpb_out[25][878],u_xpb_out[26][878],u_xpb_out[27][878],u_xpb_out[28][878],u_xpb_out[29][878],u_xpb_out[30][878],u_xpb_out[31][878],u_xpb_out[32][878],u_xpb_out[33][878],u_xpb_out[34][878],u_xpb_out[35][878],u_xpb_out[36][878],u_xpb_out[37][878],u_xpb_out[38][878],u_xpb_out[39][878],u_xpb_out[40][878],u_xpb_out[41][878],u_xpb_out[42][878],u_xpb_out[43][878],u_xpb_out[44][878],u_xpb_out[45][878],u_xpb_out[46][878],u_xpb_out[47][878],u_xpb_out[48][878],u_xpb_out[49][878],u_xpb_out[50][878],u_xpb_out[51][878],u_xpb_out[52][878],u_xpb_out[53][878],u_xpb_out[54][878],u_xpb_out[55][878],u_xpb_out[56][878],u_xpb_out[57][878],u_xpb_out[58][878],u_xpb_out[59][878],u_xpb_out[60][878],u_xpb_out[61][878],u_xpb_out[62][878],u_xpb_out[63][878],u_xpb_out[64][878],u_xpb_out[65][878],u_xpb_out[66][878],u_xpb_out[67][878],u_xpb_out[68][878],u_xpb_out[69][878],u_xpb_out[70][878],u_xpb_out[71][878],u_xpb_out[72][878],u_xpb_out[73][878],u_xpb_out[74][878],u_xpb_out[75][878],u_xpb_out[76][878],u_xpb_out[77][878],u_xpb_out[78][878],u_xpb_out[79][878],u_xpb_out[80][878],u_xpb_out[81][878],u_xpb_out[82][878],u_xpb_out[83][878],u_xpb_out[84][878],u_xpb_out[85][878],u_xpb_out[86][878],u_xpb_out[87][878],u_xpb_out[88][878],u_xpb_out[89][878],u_xpb_out[90][878],u_xpb_out[91][878],u_xpb_out[92][878],u_xpb_out[93][878],u_xpb_out[94][878],u_xpb_out[95][878],u_xpb_out[96][878],u_xpb_out[97][878],u_xpb_out[98][878],u_xpb_out[99][878],u_xpb_out[100][878],u_xpb_out[101][878],u_xpb_out[102][878],u_xpb_out[103][878],u_xpb_out[104][878],u_xpb_out[105][878]};

assign col_out_879 = {u_xpb_out[0][879],u_xpb_out[1][879],u_xpb_out[2][879],u_xpb_out[3][879],u_xpb_out[4][879],u_xpb_out[5][879],u_xpb_out[6][879],u_xpb_out[7][879],u_xpb_out[8][879],u_xpb_out[9][879],u_xpb_out[10][879],u_xpb_out[11][879],u_xpb_out[12][879],u_xpb_out[13][879],u_xpb_out[14][879],u_xpb_out[15][879],u_xpb_out[16][879],u_xpb_out[17][879],u_xpb_out[18][879],u_xpb_out[19][879],u_xpb_out[20][879],u_xpb_out[21][879],u_xpb_out[22][879],u_xpb_out[23][879],u_xpb_out[24][879],u_xpb_out[25][879],u_xpb_out[26][879],u_xpb_out[27][879],u_xpb_out[28][879],u_xpb_out[29][879],u_xpb_out[30][879],u_xpb_out[31][879],u_xpb_out[32][879],u_xpb_out[33][879],u_xpb_out[34][879],u_xpb_out[35][879],u_xpb_out[36][879],u_xpb_out[37][879],u_xpb_out[38][879],u_xpb_out[39][879],u_xpb_out[40][879],u_xpb_out[41][879],u_xpb_out[42][879],u_xpb_out[43][879],u_xpb_out[44][879],u_xpb_out[45][879],u_xpb_out[46][879],u_xpb_out[47][879],u_xpb_out[48][879],u_xpb_out[49][879],u_xpb_out[50][879],u_xpb_out[51][879],u_xpb_out[52][879],u_xpb_out[53][879],u_xpb_out[54][879],u_xpb_out[55][879],u_xpb_out[56][879],u_xpb_out[57][879],u_xpb_out[58][879],u_xpb_out[59][879],u_xpb_out[60][879],u_xpb_out[61][879],u_xpb_out[62][879],u_xpb_out[63][879],u_xpb_out[64][879],u_xpb_out[65][879],u_xpb_out[66][879],u_xpb_out[67][879],u_xpb_out[68][879],u_xpb_out[69][879],u_xpb_out[70][879],u_xpb_out[71][879],u_xpb_out[72][879],u_xpb_out[73][879],u_xpb_out[74][879],u_xpb_out[75][879],u_xpb_out[76][879],u_xpb_out[77][879],u_xpb_out[78][879],u_xpb_out[79][879],u_xpb_out[80][879],u_xpb_out[81][879],u_xpb_out[82][879],u_xpb_out[83][879],u_xpb_out[84][879],u_xpb_out[85][879],u_xpb_out[86][879],u_xpb_out[87][879],u_xpb_out[88][879],u_xpb_out[89][879],u_xpb_out[90][879],u_xpb_out[91][879],u_xpb_out[92][879],u_xpb_out[93][879],u_xpb_out[94][879],u_xpb_out[95][879],u_xpb_out[96][879],u_xpb_out[97][879],u_xpb_out[98][879],u_xpb_out[99][879],u_xpb_out[100][879],u_xpb_out[101][879],u_xpb_out[102][879],u_xpb_out[103][879],u_xpb_out[104][879],u_xpb_out[105][879]};

assign col_out_880 = {u_xpb_out[0][880],u_xpb_out[1][880],u_xpb_out[2][880],u_xpb_out[3][880],u_xpb_out[4][880],u_xpb_out[5][880],u_xpb_out[6][880],u_xpb_out[7][880],u_xpb_out[8][880],u_xpb_out[9][880],u_xpb_out[10][880],u_xpb_out[11][880],u_xpb_out[12][880],u_xpb_out[13][880],u_xpb_out[14][880],u_xpb_out[15][880],u_xpb_out[16][880],u_xpb_out[17][880],u_xpb_out[18][880],u_xpb_out[19][880],u_xpb_out[20][880],u_xpb_out[21][880],u_xpb_out[22][880],u_xpb_out[23][880],u_xpb_out[24][880],u_xpb_out[25][880],u_xpb_out[26][880],u_xpb_out[27][880],u_xpb_out[28][880],u_xpb_out[29][880],u_xpb_out[30][880],u_xpb_out[31][880],u_xpb_out[32][880],u_xpb_out[33][880],u_xpb_out[34][880],u_xpb_out[35][880],u_xpb_out[36][880],u_xpb_out[37][880],u_xpb_out[38][880],u_xpb_out[39][880],u_xpb_out[40][880],u_xpb_out[41][880],u_xpb_out[42][880],u_xpb_out[43][880],u_xpb_out[44][880],u_xpb_out[45][880],u_xpb_out[46][880],u_xpb_out[47][880],u_xpb_out[48][880],u_xpb_out[49][880],u_xpb_out[50][880],u_xpb_out[51][880],u_xpb_out[52][880],u_xpb_out[53][880],u_xpb_out[54][880],u_xpb_out[55][880],u_xpb_out[56][880],u_xpb_out[57][880],u_xpb_out[58][880],u_xpb_out[59][880],u_xpb_out[60][880],u_xpb_out[61][880],u_xpb_out[62][880],u_xpb_out[63][880],u_xpb_out[64][880],u_xpb_out[65][880],u_xpb_out[66][880],u_xpb_out[67][880],u_xpb_out[68][880],u_xpb_out[69][880],u_xpb_out[70][880],u_xpb_out[71][880],u_xpb_out[72][880],u_xpb_out[73][880],u_xpb_out[74][880],u_xpb_out[75][880],u_xpb_out[76][880],u_xpb_out[77][880],u_xpb_out[78][880],u_xpb_out[79][880],u_xpb_out[80][880],u_xpb_out[81][880],u_xpb_out[82][880],u_xpb_out[83][880],u_xpb_out[84][880],u_xpb_out[85][880],u_xpb_out[86][880],u_xpb_out[87][880],u_xpb_out[88][880],u_xpb_out[89][880],u_xpb_out[90][880],u_xpb_out[91][880],u_xpb_out[92][880],u_xpb_out[93][880],u_xpb_out[94][880],u_xpb_out[95][880],u_xpb_out[96][880],u_xpb_out[97][880],u_xpb_out[98][880],u_xpb_out[99][880],u_xpb_out[100][880],u_xpb_out[101][880],u_xpb_out[102][880],u_xpb_out[103][880],u_xpb_out[104][880],u_xpb_out[105][880]};

assign col_out_881 = {u_xpb_out[0][881],u_xpb_out[1][881],u_xpb_out[2][881],u_xpb_out[3][881],u_xpb_out[4][881],u_xpb_out[5][881],u_xpb_out[6][881],u_xpb_out[7][881],u_xpb_out[8][881],u_xpb_out[9][881],u_xpb_out[10][881],u_xpb_out[11][881],u_xpb_out[12][881],u_xpb_out[13][881],u_xpb_out[14][881],u_xpb_out[15][881],u_xpb_out[16][881],u_xpb_out[17][881],u_xpb_out[18][881],u_xpb_out[19][881],u_xpb_out[20][881],u_xpb_out[21][881],u_xpb_out[22][881],u_xpb_out[23][881],u_xpb_out[24][881],u_xpb_out[25][881],u_xpb_out[26][881],u_xpb_out[27][881],u_xpb_out[28][881],u_xpb_out[29][881],u_xpb_out[30][881],u_xpb_out[31][881],u_xpb_out[32][881],u_xpb_out[33][881],u_xpb_out[34][881],u_xpb_out[35][881],u_xpb_out[36][881],u_xpb_out[37][881],u_xpb_out[38][881],u_xpb_out[39][881],u_xpb_out[40][881],u_xpb_out[41][881],u_xpb_out[42][881],u_xpb_out[43][881],u_xpb_out[44][881],u_xpb_out[45][881],u_xpb_out[46][881],u_xpb_out[47][881],u_xpb_out[48][881],u_xpb_out[49][881],u_xpb_out[50][881],u_xpb_out[51][881],u_xpb_out[52][881],u_xpb_out[53][881],u_xpb_out[54][881],u_xpb_out[55][881],u_xpb_out[56][881],u_xpb_out[57][881],u_xpb_out[58][881],u_xpb_out[59][881],u_xpb_out[60][881],u_xpb_out[61][881],u_xpb_out[62][881],u_xpb_out[63][881],u_xpb_out[64][881],u_xpb_out[65][881],u_xpb_out[66][881],u_xpb_out[67][881],u_xpb_out[68][881],u_xpb_out[69][881],u_xpb_out[70][881],u_xpb_out[71][881],u_xpb_out[72][881],u_xpb_out[73][881],u_xpb_out[74][881],u_xpb_out[75][881],u_xpb_out[76][881],u_xpb_out[77][881],u_xpb_out[78][881],u_xpb_out[79][881],u_xpb_out[80][881],u_xpb_out[81][881],u_xpb_out[82][881],u_xpb_out[83][881],u_xpb_out[84][881],u_xpb_out[85][881],u_xpb_out[86][881],u_xpb_out[87][881],u_xpb_out[88][881],u_xpb_out[89][881],u_xpb_out[90][881],u_xpb_out[91][881],u_xpb_out[92][881],u_xpb_out[93][881],u_xpb_out[94][881],u_xpb_out[95][881],u_xpb_out[96][881],u_xpb_out[97][881],u_xpb_out[98][881],u_xpb_out[99][881],u_xpb_out[100][881],u_xpb_out[101][881],u_xpb_out[102][881],u_xpb_out[103][881],u_xpb_out[104][881],u_xpb_out[105][881]};

assign col_out_882 = {u_xpb_out[0][882],u_xpb_out[1][882],u_xpb_out[2][882],u_xpb_out[3][882],u_xpb_out[4][882],u_xpb_out[5][882],u_xpb_out[6][882],u_xpb_out[7][882],u_xpb_out[8][882],u_xpb_out[9][882],u_xpb_out[10][882],u_xpb_out[11][882],u_xpb_out[12][882],u_xpb_out[13][882],u_xpb_out[14][882],u_xpb_out[15][882],u_xpb_out[16][882],u_xpb_out[17][882],u_xpb_out[18][882],u_xpb_out[19][882],u_xpb_out[20][882],u_xpb_out[21][882],u_xpb_out[22][882],u_xpb_out[23][882],u_xpb_out[24][882],u_xpb_out[25][882],u_xpb_out[26][882],u_xpb_out[27][882],u_xpb_out[28][882],u_xpb_out[29][882],u_xpb_out[30][882],u_xpb_out[31][882],u_xpb_out[32][882],u_xpb_out[33][882],u_xpb_out[34][882],u_xpb_out[35][882],u_xpb_out[36][882],u_xpb_out[37][882],u_xpb_out[38][882],u_xpb_out[39][882],u_xpb_out[40][882],u_xpb_out[41][882],u_xpb_out[42][882],u_xpb_out[43][882],u_xpb_out[44][882],u_xpb_out[45][882],u_xpb_out[46][882],u_xpb_out[47][882],u_xpb_out[48][882],u_xpb_out[49][882],u_xpb_out[50][882],u_xpb_out[51][882],u_xpb_out[52][882],u_xpb_out[53][882],u_xpb_out[54][882],u_xpb_out[55][882],u_xpb_out[56][882],u_xpb_out[57][882],u_xpb_out[58][882],u_xpb_out[59][882],u_xpb_out[60][882],u_xpb_out[61][882],u_xpb_out[62][882],u_xpb_out[63][882],u_xpb_out[64][882],u_xpb_out[65][882],u_xpb_out[66][882],u_xpb_out[67][882],u_xpb_out[68][882],u_xpb_out[69][882],u_xpb_out[70][882],u_xpb_out[71][882],u_xpb_out[72][882],u_xpb_out[73][882],u_xpb_out[74][882],u_xpb_out[75][882],u_xpb_out[76][882],u_xpb_out[77][882],u_xpb_out[78][882],u_xpb_out[79][882],u_xpb_out[80][882],u_xpb_out[81][882],u_xpb_out[82][882],u_xpb_out[83][882],u_xpb_out[84][882],u_xpb_out[85][882],u_xpb_out[86][882],u_xpb_out[87][882],u_xpb_out[88][882],u_xpb_out[89][882],u_xpb_out[90][882],u_xpb_out[91][882],u_xpb_out[92][882],u_xpb_out[93][882],u_xpb_out[94][882],u_xpb_out[95][882],u_xpb_out[96][882],u_xpb_out[97][882],u_xpb_out[98][882],u_xpb_out[99][882],u_xpb_out[100][882],u_xpb_out[101][882],u_xpb_out[102][882],u_xpb_out[103][882],u_xpb_out[104][882],u_xpb_out[105][882]};

assign col_out_883 = {u_xpb_out[0][883],u_xpb_out[1][883],u_xpb_out[2][883],u_xpb_out[3][883],u_xpb_out[4][883],u_xpb_out[5][883],u_xpb_out[6][883],u_xpb_out[7][883],u_xpb_out[8][883],u_xpb_out[9][883],u_xpb_out[10][883],u_xpb_out[11][883],u_xpb_out[12][883],u_xpb_out[13][883],u_xpb_out[14][883],u_xpb_out[15][883],u_xpb_out[16][883],u_xpb_out[17][883],u_xpb_out[18][883],u_xpb_out[19][883],u_xpb_out[20][883],u_xpb_out[21][883],u_xpb_out[22][883],u_xpb_out[23][883],u_xpb_out[24][883],u_xpb_out[25][883],u_xpb_out[26][883],u_xpb_out[27][883],u_xpb_out[28][883],u_xpb_out[29][883],u_xpb_out[30][883],u_xpb_out[31][883],u_xpb_out[32][883],u_xpb_out[33][883],u_xpb_out[34][883],u_xpb_out[35][883],u_xpb_out[36][883],u_xpb_out[37][883],u_xpb_out[38][883],u_xpb_out[39][883],u_xpb_out[40][883],u_xpb_out[41][883],u_xpb_out[42][883],u_xpb_out[43][883],u_xpb_out[44][883],u_xpb_out[45][883],u_xpb_out[46][883],u_xpb_out[47][883],u_xpb_out[48][883],u_xpb_out[49][883],u_xpb_out[50][883],u_xpb_out[51][883],u_xpb_out[52][883],u_xpb_out[53][883],u_xpb_out[54][883],u_xpb_out[55][883],u_xpb_out[56][883],u_xpb_out[57][883],u_xpb_out[58][883],u_xpb_out[59][883],u_xpb_out[60][883],u_xpb_out[61][883],u_xpb_out[62][883],u_xpb_out[63][883],u_xpb_out[64][883],u_xpb_out[65][883],u_xpb_out[66][883],u_xpb_out[67][883],u_xpb_out[68][883],u_xpb_out[69][883],u_xpb_out[70][883],u_xpb_out[71][883],u_xpb_out[72][883],u_xpb_out[73][883],u_xpb_out[74][883],u_xpb_out[75][883],u_xpb_out[76][883],u_xpb_out[77][883],u_xpb_out[78][883],u_xpb_out[79][883],u_xpb_out[80][883],u_xpb_out[81][883],u_xpb_out[82][883],u_xpb_out[83][883],u_xpb_out[84][883],u_xpb_out[85][883],u_xpb_out[86][883],u_xpb_out[87][883],u_xpb_out[88][883],u_xpb_out[89][883],u_xpb_out[90][883],u_xpb_out[91][883],u_xpb_out[92][883],u_xpb_out[93][883],u_xpb_out[94][883],u_xpb_out[95][883],u_xpb_out[96][883],u_xpb_out[97][883],u_xpb_out[98][883],u_xpb_out[99][883],u_xpb_out[100][883],u_xpb_out[101][883],u_xpb_out[102][883],u_xpb_out[103][883],u_xpb_out[104][883],u_xpb_out[105][883]};

assign col_out_884 = {u_xpb_out[0][884],u_xpb_out[1][884],u_xpb_out[2][884],u_xpb_out[3][884],u_xpb_out[4][884],u_xpb_out[5][884],u_xpb_out[6][884],u_xpb_out[7][884],u_xpb_out[8][884],u_xpb_out[9][884],u_xpb_out[10][884],u_xpb_out[11][884],u_xpb_out[12][884],u_xpb_out[13][884],u_xpb_out[14][884],u_xpb_out[15][884],u_xpb_out[16][884],u_xpb_out[17][884],u_xpb_out[18][884],u_xpb_out[19][884],u_xpb_out[20][884],u_xpb_out[21][884],u_xpb_out[22][884],u_xpb_out[23][884],u_xpb_out[24][884],u_xpb_out[25][884],u_xpb_out[26][884],u_xpb_out[27][884],u_xpb_out[28][884],u_xpb_out[29][884],u_xpb_out[30][884],u_xpb_out[31][884],u_xpb_out[32][884],u_xpb_out[33][884],u_xpb_out[34][884],u_xpb_out[35][884],u_xpb_out[36][884],u_xpb_out[37][884],u_xpb_out[38][884],u_xpb_out[39][884],u_xpb_out[40][884],u_xpb_out[41][884],u_xpb_out[42][884],u_xpb_out[43][884],u_xpb_out[44][884],u_xpb_out[45][884],u_xpb_out[46][884],u_xpb_out[47][884],u_xpb_out[48][884],u_xpb_out[49][884],u_xpb_out[50][884],u_xpb_out[51][884],u_xpb_out[52][884],u_xpb_out[53][884],u_xpb_out[54][884],u_xpb_out[55][884],u_xpb_out[56][884],u_xpb_out[57][884],u_xpb_out[58][884],u_xpb_out[59][884],u_xpb_out[60][884],u_xpb_out[61][884],u_xpb_out[62][884],u_xpb_out[63][884],u_xpb_out[64][884],u_xpb_out[65][884],u_xpb_out[66][884],u_xpb_out[67][884],u_xpb_out[68][884],u_xpb_out[69][884],u_xpb_out[70][884],u_xpb_out[71][884],u_xpb_out[72][884],u_xpb_out[73][884],u_xpb_out[74][884],u_xpb_out[75][884],u_xpb_out[76][884],u_xpb_out[77][884],u_xpb_out[78][884],u_xpb_out[79][884],u_xpb_out[80][884],u_xpb_out[81][884],u_xpb_out[82][884],u_xpb_out[83][884],u_xpb_out[84][884],u_xpb_out[85][884],u_xpb_out[86][884],u_xpb_out[87][884],u_xpb_out[88][884],u_xpb_out[89][884],u_xpb_out[90][884],u_xpb_out[91][884],u_xpb_out[92][884],u_xpb_out[93][884],u_xpb_out[94][884],u_xpb_out[95][884],u_xpb_out[96][884],u_xpb_out[97][884],u_xpb_out[98][884],u_xpb_out[99][884],u_xpb_out[100][884],u_xpb_out[101][884],u_xpb_out[102][884],u_xpb_out[103][884],u_xpb_out[104][884],u_xpb_out[105][884]};

assign col_out_885 = {u_xpb_out[0][885],u_xpb_out[1][885],u_xpb_out[2][885],u_xpb_out[3][885],u_xpb_out[4][885],u_xpb_out[5][885],u_xpb_out[6][885],u_xpb_out[7][885],u_xpb_out[8][885],u_xpb_out[9][885],u_xpb_out[10][885],u_xpb_out[11][885],u_xpb_out[12][885],u_xpb_out[13][885],u_xpb_out[14][885],u_xpb_out[15][885],u_xpb_out[16][885],u_xpb_out[17][885],u_xpb_out[18][885],u_xpb_out[19][885],u_xpb_out[20][885],u_xpb_out[21][885],u_xpb_out[22][885],u_xpb_out[23][885],u_xpb_out[24][885],u_xpb_out[25][885],u_xpb_out[26][885],u_xpb_out[27][885],u_xpb_out[28][885],u_xpb_out[29][885],u_xpb_out[30][885],u_xpb_out[31][885],u_xpb_out[32][885],u_xpb_out[33][885],u_xpb_out[34][885],u_xpb_out[35][885],u_xpb_out[36][885],u_xpb_out[37][885],u_xpb_out[38][885],u_xpb_out[39][885],u_xpb_out[40][885],u_xpb_out[41][885],u_xpb_out[42][885],u_xpb_out[43][885],u_xpb_out[44][885],u_xpb_out[45][885],u_xpb_out[46][885],u_xpb_out[47][885],u_xpb_out[48][885],u_xpb_out[49][885],u_xpb_out[50][885],u_xpb_out[51][885],u_xpb_out[52][885],u_xpb_out[53][885],u_xpb_out[54][885],u_xpb_out[55][885],u_xpb_out[56][885],u_xpb_out[57][885],u_xpb_out[58][885],u_xpb_out[59][885],u_xpb_out[60][885],u_xpb_out[61][885],u_xpb_out[62][885],u_xpb_out[63][885],u_xpb_out[64][885],u_xpb_out[65][885],u_xpb_out[66][885],u_xpb_out[67][885],u_xpb_out[68][885],u_xpb_out[69][885],u_xpb_out[70][885],u_xpb_out[71][885],u_xpb_out[72][885],u_xpb_out[73][885],u_xpb_out[74][885],u_xpb_out[75][885],u_xpb_out[76][885],u_xpb_out[77][885],u_xpb_out[78][885],u_xpb_out[79][885],u_xpb_out[80][885],u_xpb_out[81][885],u_xpb_out[82][885],u_xpb_out[83][885],u_xpb_out[84][885],u_xpb_out[85][885],u_xpb_out[86][885],u_xpb_out[87][885],u_xpb_out[88][885],u_xpb_out[89][885],u_xpb_out[90][885],u_xpb_out[91][885],u_xpb_out[92][885],u_xpb_out[93][885],u_xpb_out[94][885],u_xpb_out[95][885],u_xpb_out[96][885],u_xpb_out[97][885],u_xpb_out[98][885],u_xpb_out[99][885],u_xpb_out[100][885],u_xpb_out[101][885],u_xpb_out[102][885],u_xpb_out[103][885],u_xpb_out[104][885],u_xpb_out[105][885]};

assign col_out_886 = {u_xpb_out[0][886],u_xpb_out[1][886],u_xpb_out[2][886],u_xpb_out[3][886],u_xpb_out[4][886],u_xpb_out[5][886],u_xpb_out[6][886],u_xpb_out[7][886],u_xpb_out[8][886],u_xpb_out[9][886],u_xpb_out[10][886],u_xpb_out[11][886],u_xpb_out[12][886],u_xpb_out[13][886],u_xpb_out[14][886],u_xpb_out[15][886],u_xpb_out[16][886],u_xpb_out[17][886],u_xpb_out[18][886],u_xpb_out[19][886],u_xpb_out[20][886],u_xpb_out[21][886],u_xpb_out[22][886],u_xpb_out[23][886],u_xpb_out[24][886],u_xpb_out[25][886],u_xpb_out[26][886],u_xpb_out[27][886],u_xpb_out[28][886],u_xpb_out[29][886],u_xpb_out[30][886],u_xpb_out[31][886],u_xpb_out[32][886],u_xpb_out[33][886],u_xpb_out[34][886],u_xpb_out[35][886],u_xpb_out[36][886],u_xpb_out[37][886],u_xpb_out[38][886],u_xpb_out[39][886],u_xpb_out[40][886],u_xpb_out[41][886],u_xpb_out[42][886],u_xpb_out[43][886],u_xpb_out[44][886],u_xpb_out[45][886],u_xpb_out[46][886],u_xpb_out[47][886],u_xpb_out[48][886],u_xpb_out[49][886],u_xpb_out[50][886],u_xpb_out[51][886],u_xpb_out[52][886],u_xpb_out[53][886],u_xpb_out[54][886],u_xpb_out[55][886],u_xpb_out[56][886],u_xpb_out[57][886],u_xpb_out[58][886],u_xpb_out[59][886],u_xpb_out[60][886],u_xpb_out[61][886],u_xpb_out[62][886],u_xpb_out[63][886],u_xpb_out[64][886],u_xpb_out[65][886],u_xpb_out[66][886],u_xpb_out[67][886],u_xpb_out[68][886],u_xpb_out[69][886],u_xpb_out[70][886],u_xpb_out[71][886],u_xpb_out[72][886],u_xpb_out[73][886],u_xpb_out[74][886],u_xpb_out[75][886],u_xpb_out[76][886],u_xpb_out[77][886],u_xpb_out[78][886],u_xpb_out[79][886],u_xpb_out[80][886],u_xpb_out[81][886],u_xpb_out[82][886],u_xpb_out[83][886],u_xpb_out[84][886],u_xpb_out[85][886],u_xpb_out[86][886],u_xpb_out[87][886],u_xpb_out[88][886],u_xpb_out[89][886],u_xpb_out[90][886],u_xpb_out[91][886],u_xpb_out[92][886],u_xpb_out[93][886],u_xpb_out[94][886],u_xpb_out[95][886],u_xpb_out[96][886],u_xpb_out[97][886],u_xpb_out[98][886],u_xpb_out[99][886],u_xpb_out[100][886],u_xpb_out[101][886],u_xpb_out[102][886],u_xpb_out[103][886],u_xpb_out[104][886],u_xpb_out[105][886]};

assign col_out_887 = {u_xpb_out[0][887],u_xpb_out[1][887],u_xpb_out[2][887],u_xpb_out[3][887],u_xpb_out[4][887],u_xpb_out[5][887],u_xpb_out[6][887],u_xpb_out[7][887],u_xpb_out[8][887],u_xpb_out[9][887],u_xpb_out[10][887],u_xpb_out[11][887],u_xpb_out[12][887],u_xpb_out[13][887],u_xpb_out[14][887],u_xpb_out[15][887],u_xpb_out[16][887],u_xpb_out[17][887],u_xpb_out[18][887],u_xpb_out[19][887],u_xpb_out[20][887],u_xpb_out[21][887],u_xpb_out[22][887],u_xpb_out[23][887],u_xpb_out[24][887],u_xpb_out[25][887],u_xpb_out[26][887],u_xpb_out[27][887],u_xpb_out[28][887],u_xpb_out[29][887],u_xpb_out[30][887],u_xpb_out[31][887],u_xpb_out[32][887],u_xpb_out[33][887],u_xpb_out[34][887],u_xpb_out[35][887],u_xpb_out[36][887],u_xpb_out[37][887],u_xpb_out[38][887],u_xpb_out[39][887],u_xpb_out[40][887],u_xpb_out[41][887],u_xpb_out[42][887],u_xpb_out[43][887],u_xpb_out[44][887],u_xpb_out[45][887],u_xpb_out[46][887],u_xpb_out[47][887],u_xpb_out[48][887],u_xpb_out[49][887],u_xpb_out[50][887],u_xpb_out[51][887],u_xpb_out[52][887],u_xpb_out[53][887],u_xpb_out[54][887],u_xpb_out[55][887],u_xpb_out[56][887],u_xpb_out[57][887],u_xpb_out[58][887],u_xpb_out[59][887],u_xpb_out[60][887],u_xpb_out[61][887],u_xpb_out[62][887],u_xpb_out[63][887],u_xpb_out[64][887],u_xpb_out[65][887],u_xpb_out[66][887],u_xpb_out[67][887],u_xpb_out[68][887],u_xpb_out[69][887],u_xpb_out[70][887],u_xpb_out[71][887],u_xpb_out[72][887],u_xpb_out[73][887],u_xpb_out[74][887],u_xpb_out[75][887],u_xpb_out[76][887],u_xpb_out[77][887],u_xpb_out[78][887],u_xpb_out[79][887],u_xpb_out[80][887],u_xpb_out[81][887],u_xpb_out[82][887],u_xpb_out[83][887],u_xpb_out[84][887],u_xpb_out[85][887],u_xpb_out[86][887],u_xpb_out[87][887],u_xpb_out[88][887],u_xpb_out[89][887],u_xpb_out[90][887],u_xpb_out[91][887],u_xpb_out[92][887],u_xpb_out[93][887],u_xpb_out[94][887],u_xpb_out[95][887],u_xpb_out[96][887],u_xpb_out[97][887],u_xpb_out[98][887],u_xpb_out[99][887],u_xpb_out[100][887],u_xpb_out[101][887],u_xpb_out[102][887],u_xpb_out[103][887],u_xpb_out[104][887],u_xpb_out[105][887]};

assign col_out_888 = {u_xpb_out[0][888],u_xpb_out[1][888],u_xpb_out[2][888],u_xpb_out[3][888],u_xpb_out[4][888],u_xpb_out[5][888],u_xpb_out[6][888],u_xpb_out[7][888],u_xpb_out[8][888],u_xpb_out[9][888],u_xpb_out[10][888],u_xpb_out[11][888],u_xpb_out[12][888],u_xpb_out[13][888],u_xpb_out[14][888],u_xpb_out[15][888],u_xpb_out[16][888],u_xpb_out[17][888],u_xpb_out[18][888],u_xpb_out[19][888],u_xpb_out[20][888],u_xpb_out[21][888],u_xpb_out[22][888],u_xpb_out[23][888],u_xpb_out[24][888],u_xpb_out[25][888],u_xpb_out[26][888],u_xpb_out[27][888],u_xpb_out[28][888],u_xpb_out[29][888],u_xpb_out[30][888],u_xpb_out[31][888],u_xpb_out[32][888],u_xpb_out[33][888],u_xpb_out[34][888],u_xpb_out[35][888],u_xpb_out[36][888],u_xpb_out[37][888],u_xpb_out[38][888],u_xpb_out[39][888],u_xpb_out[40][888],u_xpb_out[41][888],u_xpb_out[42][888],u_xpb_out[43][888],u_xpb_out[44][888],u_xpb_out[45][888],u_xpb_out[46][888],u_xpb_out[47][888],u_xpb_out[48][888],u_xpb_out[49][888],u_xpb_out[50][888],u_xpb_out[51][888],u_xpb_out[52][888],u_xpb_out[53][888],u_xpb_out[54][888],u_xpb_out[55][888],u_xpb_out[56][888],u_xpb_out[57][888],u_xpb_out[58][888],u_xpb_out[59][888],u_xpb_out[60][888],u_xpb_out[61][888],u_xpb_out[62][888],u_xpb_out[63][888],u_xpb_out[64][888],u_xpb_out[65][888],u_xpb_out[66][888],u_xpb_out[67][888],u_xpb_out[68][888],u_xpb_out[69][888],u_xpb_out[70][888],u_xpb_out[71][888],u_xpb_out[72][888],u_xpb_out[73][888],u_xpb_out[74][888],u_xpb_out[75][888],u_xpb_out[76][888],u_xpb_out[77][888],u_xpb_out[78][888],u_xpb_out[79][888],u_xpb_out[80][888],u_xpb_out[81][888],u_xpb_out[82][888],u_xpb_out[83][888],u_xpb_out[84][888],u_xpb_out[85][888],u_xpb_out[86][888],u_xpb_out[87][888],u_xpb_out[88][888],u_xpb_out[89][888],u_xpb_out[90][888],u_xpb_out[91][888],u_xpb_out[92][888],u_xpb_out[93][888],u_xpb_out[94][888],u_xpb_out[95][888],u_xpb_out[96][888],u_xpb_out[97][888],u_xpb_out[98][888],u_xpb_out[99][888],u_xpb_out[100][888],u_xpb_out[101][888],u_xpb_out[102][888],u_xpb_out[103][888],u_xpb_out[104][888],u_xpb_out[105][888]};

assign col_out_889 = {u_xpb_out[0][889],u_xpb_out[1][889],u_xpb_out[2][889],u_xpb_out[3][889],u_xpb_out[4][889],u_xpb_out[5][889],u_xpb_out[6][889],u_xpb_out[7][889],u_xpb_out[8][889],u_xpb_out[9][889],u_xpb_out[10][889],u_xpb_out[11][889],u_xpb_out[12][889],u_xpb_out[13][889],u_xpb_out[14][889],u_xpb_out[15][889],u_xpb_out[16][889],u_xpb_out[17][889],u_xpb_out[18][889],u_xpb_out[19][889],u_xpb_out[20][889],u_xpb_out[21][889],u_xpb_out[22][889],u_xpb_out[23][889],u_xpb_out[24][889],u_xpb_out[25][889],u_xpb_out[26][889],u_xpb_out[27][889],u_xpb_out[28][889],u_xpb_out[29][889],u_xpb_out[30][889],u_xpb_out[31][889],u_xpb_out[32][889],u_xpb_out[33][889],u_xpb_out[34][889],u_xpb_out[35][889],u_xpb_out[36][889],u_xpb_out[37][889],u_xpb_out[38][889],u_xpb_out[39][889],u_xpb_out[40][889],u_xpb_out[41][889],u_xpb_out[42][889],u_xpb_out[43][889],u_xpb_out[44][889],u_xpb_out[45][889],u_xpb_out[46][889],u_xpb_out[47][889],u_xpb_out[48][889],u_xpb_out[49][889],u_xpb_out[50][889],u_xpb_out[51][889],u_xpb_out[52][889],u_xpb_out[53][889],u_xpb_out[54][889],u_xpb_out[55][889],u_xpb_out[56][889],u_xpb_out[57][889],u_xpb_out[58][889],u_xpb_out[59][889],u_xpb_out[60][889],u_xpb_out[61][889],u_xpb_out[62][889],u_xpb_out[63][889],u_xpb_out[64][889],u_xpb_out[65][889],u_xpb_out[66][889],u_xpb_out[67][889],u_xpb_out[68][889],u_xpb_out[69][889],u_xpb_out[70][889],u_xpb_out[71][889],u_xpb_out[72][889],u_xpb_out[73][889],u_xpb_out[74][889],u_xpb_out[75][889],u_xpb_out[76][889],u_xpb_out[77][889],u_xpb_out[78][889],u_xpb_out[79][889],u_xpb_out[80][889],u_xpb_out[81][889],u_xpb_out[82][889],u_xpb_out[83][889],u_xpb_out[84][889],u_xpb_out[85][889],u_xpb_out[86][889],u_xpb_out[87][889],u_xpb_out[88][889],u_xpb_out[89][889],u_xpb_out[90][889],u_xpb_out[91][889],u_xpb_out[92][889],u_xpb_out[93][889],u_xpb_out[94][889],u_xpb_out[95][889],u_xpb_out[96][889],u_xpb_out[97][889],u_xpb_out[98][889],u_xpb_out[99][889],u_xpb_out[100][889],u_xpb_out[101][889],u_xpb_out[102][889],u_xpb_out[103][889],u_xpb_out[104][889],u_xpb_out[105][889]};

assign col_out_890 = {u_xpb_out[0][890],u_xpb_out[1][890],u_xpb_out[2][890],u_xpb_out[3][890],u_xpb_out[4][890],u_xpb_out[5][890],u_xpb_out[6][890],u_xpb_out[7][890],u_xpb_out[8][890],u_xpb_out[9][890],u_xpb_out[10][890],u_xpb_out[11][890],u_xpb_out[12][890],u_xpb_out[13][890],u_xpb_out[14][890],u_xpb_out[15][890],u_xpb_out[16][890],u_xpb_out[17][890],u_xpb_out[18][890],u_xpb_out[19][890],u_xpb_out[20][890],u_xpb_out[21][890],u_xpb_out[22][890],u_xpb_out[23][890],u_xpb_out[24][890],u_xpb_out[25][890],u_xpb_out[26][890],u_xpb_out[27][890],u_xpb_out[28][890],u_xpb_out[29][890],u_xpb_out[30][890],u_xpb_out[31][890],u_xpb_out[32][890],u_xpb_out[33][890],u_xpb_out[34][890],u_xpb_out[35][890],u_xpb_out[36][890],u_xpb_out[37][890],u_xpb_out[38][890],u_xpb_out[39][890],u_xpb_out[40][890],u_xpb_out[41][890],u_xpb_out[42][890],u_xpb_out[43][890],u_xpb_out[44][890],u_xpb_out[45][890],u_xpb_out[46][890],u_xpb_out[47][890],u_xpb_out[48][890],u_xpb_out[49][890],u_xpb_out[50][890],u_xpb_out[51][890],u_xpb_out[52][890],u_xpb_out[53][890],u_xpb_out[54][890],u_xpb_out[55][890],u_xpb_out[56][890],u_xpb_out[57][890],u_xpb_out[58][890],u_xpb_out[59][890],u_xpb_out[60][890],u_xpb_out[61][890],u_xpb_out[62][890],u_xpb_out[63][890],u_xpb_out[64][890],u_xpb_out[65][890],u_xpb_out[66][890],u_xpb_out[67][890],u_xpb_out[68][890],u_xpb_out[69][890],u_xpb_out[70][890],u_xpb_out[71][890],u_xpb_out[72][890],u_xpb_out[73][890],u_xpb_out[74][890],u_xpb_out[75][890],u_xpb_out[76][890],u_xpb_out[77][890],u_xpb_out[78][890],u_xpb_out[79][890],u_xpb_out[80][890],u_xpb_out[81][890],u_xpb_out[82][890],u_xpb_out[83][890],u_xpb_out[84][890],u_xpb_out[85][890],u_xpb_out[86][890],u_xpb_out[87][890],u_xpb_out[88][890],u_xpb_out[89][890],u_xpb_out[90][890],u_xpb_out[91][890],u_xpb_out[92][890],u_xpb_out[93][890],u_xpb_out[94][890],u_xpb_out[95][890],u_xpb_out[96][890],u_xpb_out[97][890],u_xpb_out[98][890],u_xpb_out[99][890],u_xpb_out[100][890],u_xpb_out[101][890],u_xpb_out[102][890],u_xpb_out[103][890],u_xpb_out[104][890],u_xpb_out[105][890]};

assign col_out_891 = {u_xpb_out[0][891],u_xpb_out[1][891],u_xpb_out[2][891],u_xpb_out[3][891],u_xpb_out[4][891],u_xpb_out[5][891],u_xpb_out[6][891],u_xpb_out[7][891],u_xpb_out[8][891],u_xpb_out[9][891],u_xpb_out[10][891],u_xpb_out[11][891],u_xpb_out[12][891],u_xpb_out[13][891],u_xpb_out[14][891],u_xpb_out[15][891],u_xpb_out[16][891],u_xpb_out[17][891],u_xpb_out[18][891],u_xpb_out[19][891],u_xpb_out[20][891],u_xpb_out[21][891],u_xpb_out[22][891],u_xpb_out[23][891],u_xpb_out[24][891],u_xpb_out[25][891],u_xpb_out[26][891],u_xpb_out[27][891],u_xpb_out[28][891],u_xpb_out[29][891],u_xpb_out[30][891],u_xpb_out[31][891],u_xpb_out[32][891],u_xpb_out[33][891],u_xpb_out[34][891],u_xpb_out[35][891],u_xpb_out[36][891],u_xpb_out[37][891],u_xpb_out[38][891],u_xpb_out[39][891],u_xpb_out[40][891],u_xpb_out[41][891],u_xpb_out[42][891],u_xpb_out[43][891],u_xpb_out[44][891],u_xpb_out[45][891],u_xpb_out[46][891],u_xpb_out[47][891],u_xpb_out[48][891],u_xpb_out[49][891],u_xpb_out[50][891],u_xpb_out[51][891],u_xpb_out[52][891],u_xpb_out[53][891],u_xpb_out[54][891],u_xpb_out[55][891],u_xpb_out[56][891],u_xpb_out[57][891],u_xpb_out[58][891],u_xpb_out[59][891],u_xpb_out[60][891],u_xpb_out[61][891],u_xpb_out[62][891],u_xpb_out[63][891],u_xpb_out[64][891],u_xpb_out[65][891],u_xpb_out[66][891],u_xpb_out[67][891],u_xpb_out[68][891],u_xpb_out[69][891],u_xpb_out[70][891],u_xpb_out[71][891],u_xpb_out[72][891],u_xpb_out[73][891],u_xpb_out[74][891],u_xpb_out[75][891],u_xpb_out[76][891],u_xpb_out[77][891],u_xpb_out[78][891],u_xpb_out[79][891],u_xpb_out[80][891],u_xpb_out[81][891],u_xpb_out[82][891],u_xpb_out[83][891],u_xpb_out[84][891],u_xpb_out[85][891],u_xpb_out[86][891],u_xpb_out[87][891],u_xpb_out[88][891],u_xpb_out[89][891],u_xpb_out[90][891],u_xpb_out[91][891],u_xpb_out[92][891],u_xpb_out[93][891],u_xpb_out[94][891],u_xpb_out[95][891],u_xpb_out[96][891],u_xpb_out[97][891],u_xpb_out[98][891],u_xpb_out[99][891],u_xpb_out[100][891],u_xpb_out[101][891],u_xpb_out[102][891],u_xpb_out[103][891],u_xpb_out[104][891],u_xpb_out[105][891]};

assign col_out_892 = {u_xpb_out[0][892],u_xpb_out[1][892],u_xpb_out[2][892],u_xpb_out[3][892],u_xpb_out[4][892],u_xpb_out[5][892],u_xpb_out[6][892],u_xpb_out[7][892],u_xpb_out[8][892],u_xpb_out[9][892],u_xpb_out[10][892],u_xpb_out[11][892],u_xpb_out[12][892],u_xpb_out[13][892],u_xpb_out[14][892],u_xpb_out[15][892],u_xpb_out[16][892],u_xpb_out[17][892],u_xpb_out[18][892],u_xpb_out[19][892],u_xpb_out[20][892],u_xpb_out[21][892],u_xpb_out[22][892],u_xpb_out[23][892],u_xpb_out[24][892],u_xpb_out[25][892],u_xpb_out[26][892],u_xpb_out[27][892],u_xpb_out[28][892],u_xpb_out[29][892],u_xpb_out[30][892],u_xpb_out[31][892],u_xpb_out[32][892],u_xpb_out[33][892],u_xpb_out[34][892],u_xpb_out[35][892],u_xpb_out[36][892],u_xpb_out[37][892],u_xpb_out[38][892],u_xpb_out[39][892],u_xpb_out[40][892],u_xpb_out[41][892],u_xpb_out[42][892],u_xpb_out[43][892],u_xpb_out[44][892],u_xpb_out[45][892],u_xpb_out[46][892],u_xpb_out[47][892],u_xpb_out[48][892],u_xpb_out[49][892],u_xpb_out[50][892],u_xpb_out[51][892],u_xpb_out[52][892],u_xpb_out[53][892],u_xpb_out[54][892],u_xpb_out[55][892],u_xpb_out[56][892],u_xpb_out[57][892],u_xpb_out[58][892],u_xpb_out[59][892],u_xpb_out[60][892],u_xpb_out[61][892],u_xpb_out[62][892],u_xpb_out[63][892],u_xpb_out[64][892],u_xpb_out[65][892],u_xpb_out[66][892],u_xpb_out[67][892],u_xpb_out[68][892],u_xpb_out[69][892],u_xpb_out[70][892],u_xpb_out[71][892],u_xpb_out[72][892],u_xpb_out[73][892],u_xpb_out[74][892],u_xpb_out[75][892],u_xpb_out[76][892],u_xpb_out[77][892],u_xpb_out[78][892],u_xpb_out[79][892],u_xpb_out[80][892],u_xpb_out[81][892],u_xpb_out[82][892],u_xpb_out[83][892],u_xpb_out[84][892],u_xpb_out[85][892],u_xpb_out[86][892],u_xpb_out[87][892],u_xpb_out[88][892],u_xpb_out[89][892],u_xpb_out[90][892],u_xpb_out[91][892],u_xpb_out[92][892],u_xpb_out[93][892],u_xpb_out[94][892],u_xpb_out[95][892],u_xpb_out[96][892],u_xpb_out[97][892],u_xpb_out[98][892],u_xpb_out[99][892],u_xpb_out[100][892],u_xpb_out[101][892],u_xpb_out[102][892],u_xpb_out[103][892],u_xpb_out[104][892],u_xpb_out[105][892]};

assign col_out_893 = {u_xpb_out[0][893],u_xpb_out[1][893],u_xpb_out[2][893],u_xpb_out[3][893],u_xpb_out[4][893],u_xpb_out[5][893],u_xpb_out[6][893],u_xpb_out[7][893],u_xpb_out[8][893],u_xpb_out[9][893],u_xpb_out[10][893],u_xpb_out[11][893],u_xpb_out[12][893],u_xpb_out[13][893],u_xpb_out[14][893],u_xpb_out[15][893],u_xpb_out[16][893],u_xpb_out[17][893],u_xpb_out[18][893],u_xpb_out[19][893],u_xpb_out[20][893],u_xpb_out[21][893],u_xpb_out[22][893],u_xpb_out[23][893],u_xpb_out[24][893],u_xpb_out[25][893],u_xpb_out[26][893],u_xpb_out[27][893],u_xpb_out[28][893],u_xpb_out[29][893],u_xpb_out[30][893],u_xpb_out[31][893],u_xpb_out[32][893],u_xpb_out[33][893],u_xpb_out[34][893],u_xpb_out[35][893],u_xpb_out[36][893],u_xpb_out[37][893],u_xpb_out[38][893],u_xpb_out[39][893],u_xpb_out[40][893],u_xpb_out[41][893],u_xpb_out[42][893],u_xpb_out[43][893],u_xpb_out[44][893],u_xpb_out[45][893],u_xpb_out[46][893],u_xpb_out[47][893],u_xpb_out[48][893],u_xpb_out[49][893],u_xpb_out[50][893],u_xpb_out[51][893],u_xpb_out[52][893],u_xpb_out[53][893],u_xpb_out[54][893],u_xpb_out[55][893],u_xpb_out[56][893],u_xpb_out[57][893],u_xpb_out[58][893],u_xpb_out[59][893],u_xpb_out[60][893],u_xpb_out[61][893],u_xpb_out[62][893],u_xpb_out[63][893],u_xpb_out[64][893],u_xpb_out[65][893],u_xpb_out[66][893],u_xpb_out[67][893],u_xpb_out[68][893],u_xpb_out[69][893],u_xpb_out[70][893],u_xpb_out[71][893],u_xpb_out[72][893],u_xpb_out[73][893],u_xpb_out[74][893],u_xpb_out[75][893],u_xpb_out[76][893],u_xpb_out[77][893],u_xpb_out[78][893],u_xpb_out[79][893],u_xpb_out[80][893],u_xpb_out[81][893],u_xpb_out[82][893],u_xpb_out[83][893],u_xpb_out[84][893],u_xpb_out[85][893],u_xpb_out[86][893],u_xpb_out[87][893],u_xpb_out[88][893],u_xpb_out[89][893],u_xpb_out[90][893],u_xpb_out[91][893],u_xpb_out[92][893],u_xpb_out[93][893],u_xpb_out[94][893],u_xpb_out[95][893],u_xpb_out[96][893],u_xpb_out[97][893],u_xpb_out[98][893],u_xpb_out[99][893],u_xpb_out[100][893],u_xpb_out[101][893],u_xpb_out[102][893],u_xpb_out[103][893],u_xpb_out[104][893],u_xpb_out[105][893]};

assign col_out_894 = {u_xpb_out[0][894],u_xpb_out[1][894],u_xpb_out[2][894],u_xpb_out[3][894],u_xpb_out[4][894],u_xpb_out[5][894],u_xpb_out[6][894],u_xpb_out[7][894],u_xpb_out[8][894],u_xpb_out[9][894],u_xpb_out[10][894],u_xpb_out[11][894],u_xpb_out[12][894],u_xpb_out[13][894],u_xpb_out[14][894],u_xpb_out[15][894],u_xpb_out[16][894],u_xpb_out[17][894],u_xpb_out[18][894],u_xpb_out[19][894],u_xpb_out[20][894],u_xpb_out[21][894],u_xpb_out[22][894],u_xpb_out[23][894],u_xpb_out[24][894],u_xpb_out[25][894],u_xpb_out[26][894],u_xpb_out[27][894],u_xpb_out[28][894],u_xpb_out[29][894],u_xpb_out[30][894],u_xpb_out[31][894],u_xpb_out[32][894],u_xpb_out[33][894],u_xpb_out[34][894],u_xpb_out[35][894],u_xpb_out[36][894],u_xpb_out[37][894],u_xpb_out[38][894],u_xpb_out[39][894],u_xpb_out[40][894],u_xpb_out[41][894],u_xpb_out[42][894],u_xpb_out[43][894],u_xpb_out[44][894],u_xpb_out[45][894],u_xpb_out[46][894],u_xpb_out[47][894],u_xpb_out[48][894],u_xpb_out[49][894],u_xpb_out[50][894],u_xpb_out[51][894],u_xpb_out[52][894],u_xpb_out[53][894],u_xpb_out[54][894],u_xpb_out[55][894],u_xpb_out[56][894],u_xpb_out[57][894],u_xpb_out[58][894],u_xpb_out[59][894],u_xpb_out[60][894],u_xpb_out[61][894],u_xpb_out[62][894],u_xpb_out[63][894],u_xpb_out[64][894],u_xpb_out[65][894],u_xpb_out[66][894],u_xpb_out[67][894],u_xpb_out[68][894],u_xpb_out[69][894],u_xpb_out[70][894],u_xpb_out[71][894],u_xpb_out[72][894],u_xpb_out[73][894],u_xpb_out[74][894],u_xpb_out[75][894],u_xpb_out[76][894],u_xpb_out[77][894],u_xpb_out[78][894],u_xpb_out[79][894],u_xpb_out[80][894],u_xpb_out[81][894],u_xpb_out[82][894],u_xpb_out[83][894],u_xpb_out[84][894],u_xpb_out[85][894],u_xpb_out[86][894],u_xpb_out[87][894],u_xpb_out[88][894],u_xpb_out[89][894],u_xpb_out[90][894],u_xpb_out[91][894],u_xpb_out[92][894],u_xpb_out[93][894],u_xpb_out[94][894],u_xpb_out[95][894],u_xpb_out[96][894],u_xpb_out[97][894],u_xpb_out[98][894],u_xpb_out[99][894],u_xpb_out[100][894],u_xpb_out[101][894],u_xpb_out[102][894],u_xpb_out[103][894],u_xpb_out[104][894],u_xpb_out[105][894]};

assign col_out_895 = {u_xpb_out[0][895],u_xpb_out[1][895],u_xpb_out[2][895],u_xpb_out[3][895],u_xpb_out[4][895],u_xpb_out[5][895],u_xpb_out[6][895],u_xpb_out[7][895],u_xpb_out[8][895],u_xpb_out[9][895],u_xpb_out[10][895],u_xpb_out[11][895],u_xpb_out[12][895],u_xpb_out[13][895],u_xpb_out[14][895],u_xpb_out[15][895],u_xpb_out[16][895],u_xpb_out[17][895],u_xpb_out[18][895],u_xpb_out[19][895],u_xpb_out[20][895],u_xpb_out[21][895],u_xpb_out[22][895],u_xpb_out[23][895],u_xpb_out[24][895],u_xpb_out[25][895],u_xpb_out[26][895],u_xpb_out[27][895],u_xpb_out[28][895],u_xpb_out[29][895],u_xpb_out[30][895],u_xpb_out[31][895],u_xpb_out[32][895],u_xpb_out[33][895],u_xpb_out[34][895],u_xpb_out[35][895],u_xpb_out[36][895],u_xpb_out[37][895],u_xpb_out[38][895],u_xpb_out[39][895],u_xpb_out[40][895],u_xpb_out[41][895],u_xpb_out[42][895],u_xpb_out[43][895],u_xpb_out[44][895],u_xpb_out[45][895],u_xpb_out[46][895],u_xpb_out[47][895],u_xpb_out[48][895],u_xpb_out[49][895],u_xpb_out[50][895],u_xpb_out[51][895],u_xpb_out[52][895],u_xpb_out[53][895],u_xpb_out[54][895],u_xpb_out[55][895],u_xpb_out[56][895],u_xpb_out[57][895],u_xpb_out[58][895],u_xpb_out[59][895],u_xpb_out[60][895],u_xpb_out[61][895],u_xpb_out[62][895],u_xpb_out[63][895],u_xpb_out[64][895],u_xpb_out[65][895],u_xpb_out[66][895],u_xpb_out[67][895],u_xpb_out[68][895],u_xpb_out[69][895],u_xpb_out[70][895],u_xpb_out[71][895],u_xpb_out[72][895],u_xpb_out[73][895],u_xpb_out[74][895],u_xpb_out[75][895],u_xpb_out[76][895],u_xpb_out[77][895],u_xpb_out[78][895],u_xpb_out[79][895],u_xpb_out[80][895],u_xpb_out[81][895],u_xpb_out[82][895],u_xpb_out[83][895],u_xpb_out[84][895],u_xpb_out[85][895],u_xpb_out[86][895],u_xpb_out[87][895],u_xpb_out[88][895],u_xpb_out[89][895],u_xpb_out[90][895],u_xpb_out[91][895],u_xpb_out[92][895],u_xpb_out[93][895],u_xpb_out[94][895],u_xpb_out[95][895],u_xpb_out[96][895],u_xpb_out[97][895],u_xpb_out[98][895],u_xpb_out[99][895],u_xpb_out[100][895],u_xpb_out[101][895],u_xpb_out[102][895],u_xpb_out[103][895],u_xpb_out[104][895],u_xpb_out[105][895]};

assign col_out_896 = {u_xpb_out[0][896],u_xpb_out[1][896],u_xpb_out[2][896],u_xpb_out[3][896],u_xpb_out[4][896],u_xpb_out[5][896],u_xpb_out[6][896],u_xpb_out[7][896],u_xpb_out[8][896],u_xpb_out[9][896],u_xpb_out[10][896],u_xpb_out[11][896],u_xpb_out[12][896],u_xpb_out[13][896],u_xpb_out[14][896],u_xpb_out[15][896],u_xpb_out[16][896],u_xpb_out[17][896],u_xpb_out[18][896],u_xpb_out[19][896],u_xpb_out[20][896],u_xpb_out[21][896],u_xpb_out[22][896],u_xpb_out[23][896],u_xpb_out[24][896],u_xpb_out[25][896],u_xpb_out[26][896],u_xpb_out[27][896],u_xpb_out[28][896],u_xpb_out[29][896],u_xpb_out[30][896],u_xpb_out[31][896],u_xpb_out[32][896],u_xpb_out[33][896],u_xpb_out[34][896],u_xpb_out[35][896],u_xpb_out[36][896],u_xpb_out[37][896],u_xpb_out[38][896],u_xpb_out[39][896],u_xpb_out[40][896],u_xpb_out[41][896],u_xpb_out[42][896],u_xpb_out[43][896],u_xpb_out[44][896],u_xpb_out[45][896],u_xpb_out[46][896],u_xpb_out[47][896],u_xpb_out[48][896],u_xpb_out[49][896],u_xpb_out[50][896],u_xpb_out[51][896],u_xpb_out[52][896],u_xpb_out[53][896],u_xpb_out[54][896],u_xpb_out[55][896],u_xpb_out[56][896],u_xpb_out[57][896],u_xpb_out[58][896],u_xpb_out[59][896],u_xpb_out[60][896],u_xpb_out[61][896],u_xpb_out[62][896],u_xpb_out[63][896],u_xpb_out[64][896],u_xpb_out[65][896],u_xpb_out[66][896],u_xpb_out[67][896],u_xpb_out[68][896],u_xpb_out[69][896],u_xpb_out[70][896],u_xpb_out[71][896],u_xpb_out[72][896],u_xpb_out[73][896],u_xpb_out[74][896],u_xpb_out[75][896],u_xpb_out[76][896],u_xpb_out[77][896],u_xpb_out[78][896],u_xpb_out[79][896],u_xpb_out[80][896],u_xpb_out[81][896],u_xpb_out[82][896],u_xpb_out[83][896],u_xpb_out[84][896],u_xpb_out[85][896],u_xpb_out[86][896],u_xpb_out[87][896],u_xpb_out[88][896],u_xpb_out[89][896],u_xpb_out[90][896],u_xpb_out[91][896],u_xpb_out[92][896],u_xpb_out[93][896],u_xpb_out[94][896],u_xpb_out[95][896],u_xpb_out[96][896],u_xpb_out[97][896],u_xpb_out[98][896],u_xpb_out[99][896],u_xpb_out[100][896],u_xpb_out[101][896],u_xpb_out[102][896],u_xpb_out[103][896],u_xpb_out[104][896],u_xpb_out[105][896]};

assign col_out_897 = {u_xpb_out[0][897],u_xpb_out[1][897],u_xpb_out[2][897],u_xpb_out[3][897],u_xpb_out[4][897],u_xpb_out[5][897],u_xpb_out[6][897],u_xpb_out[7][897],u_xpb_out[8][897],u_xpb_out[9][897],u_xpb_out[10][897],u_xpb_out[11][897],u_xpb_out[12][897],u_xpb_out[13][897],u_xpb_out[14][897],u_xpb_out[15][897],u_xpb_out[16][897],u_xpb_out[17][897],u_xpb_out[18][897],u_xpb_out[19][897],u_xpb_out[20][897],u_xpb_out[21][897],u_xpb_out[22][897],u_xpb_out[23][897],u_xpb_out[24][897],u_xpb_out[25][897],u_xpb_out[26][897],u_xpb_out[27][897],u_xpb_out[28][897],u_xpb_out[29][897],u_xpb_out[30][897],u_xpb_out[31][897],u_xpb_out[32][897],u_xpb_out[33][897],u_xpb_out[34][897],u_xpb_out[35][897],u_xpb_out[36][897],u_xpb_out[37][897],u_xpb_out[38][897],u_xpb_out[39][897],u_xpb_out[40][897],u_xpb_out[41][897],u_xpb_out[42][897],u_xpb_out[43][897],u_xpb_out[44][897],u_xpb_out[45][897],u_xpb_out[46][897],u_xpb_out[47][897],u_xpb_out[48][897],u_xpb_out[49][897],u_xpb_out[50][897],u_xpb_out[51][897],u_xpb_out[52][897],u_xpb_out[53][897],u_xpb_out[54][897],u_xpb_out[55][897],u_xpb_out[56][897],u_xpb_out[57][897],u_xpb_out[58][897],u_xpb_out[59][897],u_xpb_out[60][897],u_xpb_out[61][897],u_xpb_out[62][897],u_xpb_out[63][897],u_xpb_out[64][897],u_xpb_out[65][897],u_xpb_out[66][897],u_xpb_out[67][897],u_xpb_out[68][897],u_xpb_out[69][897],u_xpb_out[70][897],u_xpb_out[71][897],u_xpb_out[72][897],u_xpb_out[73][897],u_xpb_out[74][897],u_xpb_out[75][897],u_xpb_out[76][897],u_xpb_out[77][897],u_xpb_out[78][897],u_xpb_out[79][897],u_xpb_out[80][897],u_xpb_out[81][897],u_xpb_out[82][897],u_xpb_out[83][897],u_xpb_out[84][897],u_xpb_out[85][897],u_xpb_out[86][897],u_xpb_out[87][897],u_xpb_out[88][897],u_xpb_out[89][897],u_xpb_out[90][897],u_xpb_out[91][897],u_xpb_out[92][897],u_xpb_out[93][897],u_xpb_out[94][897],u_xpb_out[95][897],u_xpb_out[96][897],u_xpb_out[97][897],u_xpb_out[98][897],u_xpb_out[99][897],u_xpb_out[100][897],u_xpb_out[101][897],u_xpb_out[102][897],u_xpb_out[103][897],u_xpb_out[104][897],u_xpb_out[105][897]};

assign col_out_898 = {u_xpb_out[0][898],u_xpb_out[1][898],u_xpb_out[2][898],u_xpb_out[3][898],u_xpb_out[4][898],u_xpb_out[5][898],u_xpb_out[6][898],u_xpb_out[7][898],u_xpb_out[8][898],u_xpb_out[9][898],u_xpb_out[10][898],u_xpb_out[11][898],u_xpb_out[12][898],u_xpb_out[13][898],u_xpb_out[14][898],u_xpb_out[15][898],u_xpb_out[16][898],u_xpb_out[17][898],u_xpb_out[18][898],u_xpb_out[19][898],u_xpb_out[20][898],u_xpb_out[21][898],u_xpb_out[22][898],u_xpb_out[23][898],u_xpb_out[24][898],u_xpb_out[25][898],u_xpb_out[26][898],u_xpb_out[27][898],u_xpb_out[28][898],u_xpb_out[29][898],u_xpb_out[30][898],u_xpb_out[31][898],u_xpb_out[32][898],u_xpb_out[33][898],u_xpb_out[34][898],u_xpb_out[35][898],u_xpb_out[36][898],u_xpb_out[37][898],u_xpb_out[38][898],u_xpb_out[39][898],u_xpb_out[40][898],u_xpb_out[41][898],u_xpb_out[42][898],u_xpb_out[43][898],u_xpb_out[44][898],u_xpb_out[45][898],u_xpb_out[46][898],u_xpb_out[47][898],u_xpb_out[48][898],u_xpb_out[49][898],u_xpb_out[50][898],u_xpb_out[51][898],u_xpb_out[52][898],u_xpb_out[53][898],u_xpb_out[54][898],u_xpb_out[55][898],u_xpb_out[56][898],u_xpb_out[57][898],u_xpb_out[58][898],u_xpb_out[59][898],u_xpb_out[60][898],u_xpb_out[61][898],u_xpb_out[62][898],u_xpb_out[63][898],u_xpb_out[64][898],u_xpb_out[65][898],u_xpb_out[66][898],u_xpb_out[67][898],u_xpb_out[68][898],u_xpb_out[69][898],u_xpb_out[70][898],u_xpb_out[71][898],u_xpb_out[72][898],u_xpb_out[73][898],u_xpb_out[74][898],u_xpb_out[75][898],u_xpb_out[76][898],u_xpb_out[77][898],u_xpb_out[78][898],u_xpb_out[79][898],u_xpb_out[80][898],u_xpb_out[81][898],u_xpb_out[82][898],u_xpb_out[83][898],u_xpb_out[84][898],u_xpb_out[85][898],u_xpb_out[86][898],u_xpb_out[87][898],u_xpb_out[88][898],u_xpb_out[89][898],u_xpb_out[90][898],u_xpb_out[91][898],u_xpb_out[92][898],u_xpb_out[93][898],u_xpb_out[94][898],u_xpb_out[95][898],u_xpb_out[96][898],u_xpb_out[97][898],u_xpb_out[98][898],u_xpb_out[99][898],u_xpb_out[100][898],u_xpb_out[101][898],u_xpb_out[102][898],u_xpb_out[103][898],u_xpb_out[104][898],u_xpb_out[105][898]};

assign col_out_899 = {u_xpb_out[0][899],u_xpb_out[1][899],u_xpb_out[2][899],u_xpb_out[3][899],u_xpb_out[4][899],u_xpb_out[5][899],u_xpb_out[6][899],u_xpb_out[7][899],u_xpb_out[8][899],u_xpb_out[9][899],u_xpb_out[10][899],u_xpb_out[11][899],u_xpb_out[12][899],u_xpb_out[13][899],u_xpb_out[14][899],u_xpb_out[15][899],u_xpb_out[16][899],u_xpb_out[17][899],u_xpb_out[18][899],u_xpb_out[19][899],u_xpb_out[20][899],u_xpb_out[21][899],u_xpb_out[22][899],u_xpb_out[23][899],u_xpb_out[24][899],u_xpb_out[25][899],u_xpb_out[26][899],u_xpb_out[27][899],u_xpb_out[28][899],u_xpb_out[29][899],u_xpb_out[30][899],u_xpb_out[31][899],u_xpb_out[32][899],u_xpb_out[33][899],u_xpb_out[34][899],u_xpb_out[35][899],u_xpb_out[36][899],u_xpb_out[37][899],u_xpb_out[38][899],u_xpb_out[39][899],u_xpb_out[40][899],u_xpb_out[41][899],u_xpb_out[42][899],u_xpb_out[43][899],u_xpb_out[44][899],u_xpb_out[45][899],u_xpb_out[46][899],u_xpb_out[47][899],u_xpb_out[48][899],u_xpb_out[49][899],u_xpb_out[50][899],u_xpb_out[51][899],u_xpb_out[52][899],u_xpb_out[53][899],u_xpb_out[54][899],u_xpb_out[55][899],u_xpb_out[56][899],u_xpb_out[57][899],u_xpb_out[58][899],u_xpb_out[59][899],u_xpb_out[60][899],u_xpb_out[61][899],u_xpb_out[62][899],u_xpb_out[63][899],u_xpb_out[64][899],u_xpb_out[65][899],u_xpb_out[66][899],u_xpb_out[67][899],u_xpb_out[68][899],u_xpb_out[69][899],u_xpb_out[70][899],u_xpb_out[71][899],u_xpb_out[72][899],u_xpb_out[73][899],u_xpb_out[74][899],u_xpb_out[75][899],u_xpb_out[76][899],u_xpb_out[77][899],u_xpb_out[78][899],u_xpb_out[79][899],u_xpb_out[80][899],u_xpb_out[81][899],u_xpb_out[82][899],u_xpb_out[83][899],u_xpb_out[84][899],u_xpb_out[85][899],u_xpb_out[86][899],u_xpb_out[87][899],u_xpb_out[88][899],u_xpb_out[89][899],u_xpb_out[90][899],u_xpb_out[91][899],u_xpb_out[92][899],u_xpb_out[93][899],u_xpb_out[94][899],u_xpb_out[95][899],u_xpb_out[96][899],u_xpb_out[97][899],u_xpb_out[98][899],u_xpb_out[99][899],u_xpb_out[100][899],u_xpb_out[101][899],u_xpb_out[102][899],u_xpb_out[103][899],u_xpb_out[104][899],u_xpb_out[105][899]};

assign col_out_900 = {u_xpb_out[0][900],u_xpb_out[1][900],u_xpb_out[2][900],u_xpb_out[3][900],u_xpb_out[4][900],u_xpb_out[5][900],u_xpb_out[6][900],u_xpb_out[7][900],u_xpb_out[8][900],u_xpb_out[9][900],u_xpb_out[10][900],u_xpb_out[11][900],u_xpb_out[12][900],u_xpb_out[13][900],u_xpb_out[14][900],u_xpb_out[15][900],u_xpb_out[16][900],u_xpb_out[17][900],u_xpb_out[18][900],u_xpb_out[19][900],u_xpb_out[20][900],u_xpb_out[21][900],u_xpb_out[22][900],u_xpb_out[23][900],u_xpb_out[24][900],u_xpb_out[25][900],u_xpb_out[26][900],u_xpb_out[27][900],u_xpb_out[28][900],u_xpb_out[29][900],u_xpb_out[30][900],u_xpb_out[31][900],u_xpb_out[32][900],u_xpb_out[33][900],u_xpb_out[34][900],u_xpb_out[35][900],u_xpb_out[36][900],u_xpb_out[37][900],u_xpb_out[38][900],u_xpb_out[39][900],u_xpb_out[40][900],u_xpb_out[41][900],u_xpb_out[42][900],u_xpb_out[43][900],u_xpb_out[44][900],u_xpb_out[45][900],u_xpb_out[46][900],u_xpb_out[47][900],u_xpb_out[48][900],u_xpb_out[49][900],u_xpb_out[50][900],u_xpb_out[51][900],u_xpb_out[52][900],u_xpb_out[53][900],u_xpb_out[54][900],u_xpb_out[55][900],u_xpb_out[56][900],u_xpb_out[57][900],u_xpb_out[58][900],u_xpb_out[59][900],u_xpb_out[60][900],u_xpb_out[61][900],u_xpb_out[62][900],u_xpb_out[63][900],u_xpb_out[64][900],u_xpb_out[65][900],u_xpb_out[66][900],u_xpb_out[67][900],u_xpb_out[68][900],u_xpb_out[69][900],u_xpb_out[70][900],u_xpb_out[71][900],u_xpb_out[72][900],u_xpb_out[73][900],u_xpb_out[74][900],u_xpb_out[75][900],u_xpb_out[76][900],u_xpb_out[77][900],u_xpb_out[78][900],u_xpb_out[79][900],u_xpb_out[80][900],u_xpb_out[81][900],u_xpb_out[82][900],u_xpb_out[83][900],u_xpb_out[84][900],u_xpb_out[85][900],u_xpb_out[86][900],u_xpb_out[87][900],u_xpb_out[88][900],u_xpb_out[89][900],u_xpb_out[90][900],u_xpb_out[91][900],u_xpb_out[92][900],u_xpb_out[93][900],u_xpb_out[94][900],u_xpb_out[95][900],u_xpb_out[96][900],u_xpb_out[97][900],u_xpb_out[98][900],u_xpb_out[99][900],u_xpb_out[100][900],u_xpb_out[101][900],u_xpb_out[102][900],u_xpb_out[103][900],u_xpb_out[104][900],u_xpb_out[105][900]};

assign col_out_901 = {u_xpb_out[0][901],u_xpb_out[1][901],u_xpb_out[2][901],u_xpb_out[3][901],u_xpb_out[4][901],u_xpb_out[5][901],u_xpb_out[6][901],u_xpb_out[7][901],u_xpb_out[8][901],u_xpb_out[9][901],u_xpb_out[10][901],u_xpb_out[11][901],u_xpb_out[12][901],u_xpb_out[13][901],u_xpb_out[14][901],u_xpb_out[15][901],u_xpb_out[16][901],u_xpb_out[17][901],u_xpb_out[18][901],u_xpb_out[19][901],u_xpb_out[20][901],u_xpb_out[21][901],u_xpb_out[22][901],u_xpb_out[23][901],u_xpb_out[24][901],u_xpb_out[25][901],u_xpb_out[26][901],u_xpb_out[27][901],u_xpb_out[28][901],u_xpb_out[29][901],u_xpb_out[30][901],u_xpb_out[31][901],u_xpb_out[32][901],u_xpb_out[33][901],u_xpb_out[34][901],u_xpb_out[35][901],u_xpb_out[36][901],u_xpb_out[37][901],u_xpb_out[38][901],u_xpb_out[39][901],u_xpb_out[40][901],u_xpb_out[41][901],u_xpb_out[42][901],u_xpb_out[43][901],u_xpb_out[44][901],u_xpb_out[45][901],u_xpb_out[46][901],u_xpb_out[47][901],u_xpb_out[48][901],u_xpb_out[49][901],u_xpb_out[50][901],u_xpb_out[51][901],u_xpb_out[52][901],u_xpb_out[53][901],u_xpb_out[54][901],u_xpb_out[55][901],u_xpb_out[56][901],u_xpb_out[57][901],u_xpb_out[58][901],u_xpb_out[59][901],u_xpb_out[60][901],u_xpb_out[61][901],u_xpb_out[62][901],u_xpb_out[63][901],u_xpb_out[64][901],u_xpb_out[65][901],u_xpb_out[66][901],u_xpb_out[67][901],u_xpb_out[68][901],u_xpb_out[69][901],u_xpb_out[70][901],u_xpb_out[71][901],u_xpb_out[72][901],u_xpb_out[73][901],u_xpb_out[74][901],u_xpb_out[75][901],u_xpb_out[76][901],u_xpb_out[77][901],u_xpb_out[78][901],u_xpb_out[79][901],u_xpb_out[80][901],u_xpb_out[81][901],u_xpb_out[82][901],u_xpb_out[83][901],u_xpb_out[84][901],u_xpb_out[85][901],u_xpb_out[86][901],u_xpb_out[87][901],u_xpb_out[88][901],u_xpb_out[89][901],u_xpb_out[90][901],u_xpb_out[91][901],u_xpb_out[92][901],u_xpb_out[93][901],u_xpb_out[94][901],u_xpb_out[95][901],u_xpb_out[96][901],u_xpb_out[97][901],u_xpb_out[98][901],u_xpb_out[99][901],u_xpb_out[100][901],u_xpb_out[101][901],u_xpb_out[102][901],u_xpb_out[103][901],u_xpb_out[104][901],u_xpb_out[105][901]};

assign col_out_902 = {u_xpb_out[0][902],u_xpb_out[1][902],u_xpb_out[2][902],u_xpb_out[3][902],u_xpb_out[4][902],u_xpb_out[5][902],u_xpb_out[6][902],u_xpb_out[7][902],u_xpb_out[8][902],u_xpb_out[9][902],u_xpb_out[10][902],u_xpb_out[11][902],u_xpb_out[12][902],u_xpb_out[13][902],u_xpb_out[14][902],u_xpb_out[15][902],u_xpb_out[16][902],u_xpb_out[17][902],u_xpb_out[18][902],u_xpb_out[19][902],u_xpb_out[20][902],u_xpb_out[21][902],u_xpb_out[22][902],u_xpb_out[23][902],u_xpb_out[24][902],u_xpb_out[25][902],u_xpb_out[26][902],u_xpb_out[27][902],u_xpb_out[28][902],u_xpb_out[29][902],u_xpb_out[30][902],u_xpb_out[31][902],u_xpb_out[32][902],u_xpb_out[33][902],u_xpb_out[34][902],u_xpb_out[35][902],u_xpb_out[36][902],u_xpb_out[37][902],u_xpb_out[38][902],u_xpb_out[39][902],u_xpb_out[40][902],u_xpb_out[41][902],u_xpb_out[42][902],u_xpb_out[43][902],u_xpb_out[44][902],u_xpb_out[45][902],u_xpb_out[46][902],u_xpb_out[47][902],u_xpb_out[48][902],u_xpb_out[49][902],u_xpb_out[50][902],u_xpb_out[51][902],u_xpb_out[52][902],u_xpb_out[53][902],u_xpb_out[54][902],u_xpb_out[55][902],u_xpb_out[56][902],u_xpb_out[57][902],u_xpb_out[58][902],u_xpb_out[59][902],u_xpb_out[60][902],u_xpb_out[61][902],u_xpb_out[62][902],u_xpb_out[63][902],u_xpb_out[64][902],u_xpb_out[65][902],u_xpb_out[66][902],u_xpb_out[67][902],u_xpb_out[68][902],u_xpb_out[69][902],u_xpb_out[70][902],u_xpb_out[71][902],u_xpb_out[72][902],u_xpb_out[73][902],u_xpb_out[74][902],u_xpb_out[75][902],u_xpb_out[76][902],u_xpb_out[77][902],u_xpb_out[78][902],u_xpb_out[79][902],u_xpb_out[80][902],u_xpb_out[81][902],u_xpb_out[82][902],u_xpb_out[83][902],u_xpb_out[84][902],u_xpb_out[85][902],u_xpb_out[86][902],u_xpb_out[87][902],u_xpb_out[88][902],u_xpb_out[89][902],u_xpb_out[90][902],u_xpb_out[91][902],u_xpb_out[92][902],u_xpb_out[93][902],u_xpb_out[94][902],u_xpb_out[95][902],u_xpb_out[96][902],u_xpb_out[97][902],u_xpb_out[98][902],u_xpb_out[99][902],u_xpb_out[100][902],u_xpb_out[101][902],u_xpb_out[102][902],u_xpb_out[103][902],u_xpb_out[104][902],u_xpb_out[105][902]};

assign col_out_903 = {u_xpb_out[0][903],u_xpb_out[1][903],u_xpb_out[2][903],u_xpb_out[3][903],u_xpb_out[4][903],u_xpb_out[5][903],u_xpb_out[6][903],u_xpb_out[7][903],u_xpb_out[8][903],u_xpb_out[9][903],u_xpb_out[10][903],u_xpb_out[11][903],u_xpb_out[12][903],u_xpb_out[13][903],u_xpb_out[14][903],u_xpb_out[15][903],u_xpb_out[16][903],u_xpb_out[17][903],u_xpb_out[18][903],u_xpb_out[19][903],u_xpb_out[20][903],u_xpb_out[21][903],u_xpb_out[22][903],u_xpb_out[23][903],u_xpb_out[24][903],u_xpb_out[25][903],u_xpb_out[26][903],u_xpb_out[27][903],u_xpb_out[28][903],u_xpb_out[29][903],u_xpb_out[30][903],u_xpb_out[31][903],u_xpb_out[32][903],u_xpb_out[33][903],u_xpb_out[34][903],u_xpb_out[35][903],u_xpb_out[36][903],u_xpb_out[37][903],u_xpb_out[38][903],u_xpb_out[39][903],u_xpb_out[40][903],u_xpb_out[41][903],u_xpb_out[42][903],u_xpb_out[43][903],u_xpb_out[44][903],u_xpb_out[45][903],u_xpb_out[46][903],u_xpb_out[47][903],u_xpb_out[48][903],u_xpb_out[49][903],u_xpb_out[50][903],u_xpb_out[51][903],u_xpb_out[52][903],u_xpb_out[53][903],u_xpb_out[54][903],u_xpb_out[55][903],u_xpb_out[56][903],u_xpb_out[57][903],u_xpb_out[58][903],u_xpb_out[59][903],u_xpb_out[60][903],u_xpb_out[61][903],u_xpb_out[62][903],u_xpb_out[63][903],u_xpb_out[64][903],u_xpb_out[65][903],u_xpb_out[66][903],u_xpb_out[67][903],u_xpb_out[68][903],u_xpb_out[69][903],u_xpb_out[70][903],u_xpb_out[71][903],u_xpb_out[72][903],u_xpb_out[73][903],u_xpb_out[74][903],u_xpb_out[75][903],u_xpb_out[76][903],u_xpb_out[77][903],u_xpb_out[78][903],u_xpb_out[79][903],u_xpb_out[80][903],u_xpb_out[81][903],u_xpb_out[82][903],u_xpb_out[83][903],u_xpb_out[84][903],u_xpb_out[85][903],u_xpb_out[86][903],u_xpb_out[87][903],u_xpb_out[88][903],u_xpb_out[89][903],u_xpb_out[90][903],u_xpb_out[91][903],u_xpb_out[92][903],u_xpb_out[93][903],u_xpb_out[94][903],u_xpb_out[95][903],u_xpb_out[96][903],u_xpb_out[97][903],u_xpb_out[98][903],u_xpb_out[99][903],u_xpb_out[100][903],u_xpb_out[101][903],u_xpb_out[102][903],u_xpb_out[103][903],u_xpb_out[104][903],u_xpb_out[105][903]};

assign col_out_904 = {u_xpb_out[0][904],u_xpb_out[1][904],u_xpb_out[2][904],u_xpb_out[3][904],u_xpb_out[4][904],u_xpb_out[5][904],u_xpb_out[6][904],u_xpb_out[7][904],u_xpb_out[8][904],u_xpb_out[9][904],u_xpb_out[10][904],u_xpb_out[11][904],u_xpb_out[12][904],u_xpb_out[13][904],u_xpb_out[14][904],u_xpb_out[15][904],u_xpb_out[16][904],u_xpb_out[17][904],u_xpb_out[18][904],u_xpb_out[19][904],u_xpb_out[20][904],u_xpb_out[21][904],u_xpb_out[22][904],u_xpb_out[23][904],u_xpb_out[24][904],u_xpb_out[25][904],u_xpb_out[26][904],u_xpb_out[27][904],u_xpb_out[28][904],u_xpb_out[29][904],u_xpb_out[30][904],u_xpb_out[31][904],u_xpb_out[32][904],u_xpb_out[33][904],u_xpb_out[34][904],u_xpb_out[35][904],u_xpb_out[36][904],u_xpb_out[37][904],u_xpb_out[38][904],u_xpb_out[39][904],u_xpb_out[40][904],u_xpb_out[41][904],u_xpb_out[42][904],u_xpb_out[43][904],u_xpb_out[44][904],u_xpb_out[45][904],u_xpb_out[46][904],u_xpb_out[47][904],u_xpb_out[48][904],u_xpb_out[49][904],u_xpb_out[50][904],u_xpb_out[51][904],u_xpb_out[52][904],u_xpb_out[53][904],u_xpb_out[54][904],u_xpb_out[55][904],u_xpb_out[56][904],u_xpb_out[57][904],u_xpb_out[58][904],u_xpb_out[59][904],u_xpb_out[60][904],u_xpb_out[61][904],u_xpb_out[62][904],u_xpb_out[63][904],u_xpb_out[64][904],u_xpb_out[65][904],u_xpb_out[66][904],u_xpb_out[67][904],u_xpb_out[68][904],u_xpb_out[69][904],u_xpb_out[70][904],u_xpb_out[71][904],u_xpb_out[72][904],u_xpb_out[73][904],u_xpb_out[74][904],u_xpb_out[75][904],u_xpb_out[76][904],u_xpb_out[77][904],u_xpb_out[78][904],u_xpb_out[79][904],u_xpb_out[80][904],u_xpb_out[81][904],u_xpb_out[82][904],u_xpb_out[83][904],u_xpb_out[84][904],u_xpb_out[85][904],u_xpb_out[86][904],u_xpb_out[87][904],u_xpb_out[88][904],u_xpb_out[89][904],u_xpb_out[90][904],u_xpb_out[91][904],u_xpb_out[92][904],u_xpb_out[93][904],u_xpb_out[94][904],u_xpb_out[95][904],u_xpb_out[96][904],u_xpb_out[97][904],u_xpb_out[98][904],u_xpb_out[99][904],u_xpb_out[100][904],u_xpb_out[101][904],u_xpb_out[102][904],u_xpb_out[103][904],u_xpb_out[104][904],u_xpb_out[105][904]};

assign col_out_905 = {u_xpb_out[0][905],u_xpb_out[1][905],u_xpb_out[2][905],u_xpb_out[3][905],u_xpb_out[4][905],u_xpb_out[5][905],u_xpb_out[6][905],u_xpb_out[7][905],u_xpb_out[8][905],u_xpb_out[9][905],u_xpb_out[10][905],u_xpb_out[11][905],u_xpb_out[12][905],u_xpb_out[13][905],u_xpb_out[14][905],u_xpb_out[15][905],u_xpb_out[16][905],u_xpb_out[17][905],u_xpb_out[18][905],u_xpb_out[19][905],u_xpb_out[20][905],u_xpb_out[21][905],u_xpb_out[22][905],u_xpb_out[23][905],u_xpb_out[24][905],u_xpb_out[25][905],u_xpb_out[26][905],u_xpb_out[27][905],u_xpb_out[28][905],u_xpb_out[29][905],u_xpb_out[30][905],u_xpb_out[31][905],u_xpb_out[32][905],u_xpb_out[33][905],u_xpb_out[34][905],u_xpb_out[35][905],u_xpb_out[36][905],u_xpb_out[37][905],u_xpb_out[38][905],u_xpb_out[39][905],u_xpb_out[40][905],u_xpb_out[41][905],u_xpb_out[42][905],u_xpb_out[43][905],u_xpb_out[44][905],u_xpb_out[45][905],u_xpb_out[46][905],u_xpb_out[47][905],u_xpb_out[48][905],u_xpb_out[49][905],u_xpb_out[50][905],u_xpb_out[51][905],u_xpb_out[52][905],u_xpb_out[53][905],u_xpb_out[54][905],u_xpb_out[55][905],u_xpb_out[56][905],u_xpb_out[57][905],u_xpb_out[58][905],u_xpb_out[59][905],u_xpb_out[60][905],u_xpb_out[61][905],u_xpb_out[62][905],u_xpb_out[63][905],u_xpb_out[64][905],u_xpb_out[65][905],u_xpb_out[66][905],u_xpb_out[67][905],u_xpb_out[68][905],u_xpb_out[69][905],u_xpb_out[70][905],u_xpb_out[71][905],u_xpb_out[72][905],u_xpb_out[73][905],u_xpb_out[74][905],u_xpb_out[75][905],u_xpb_out[76][905],u_xpb_out[77][905],u_xpb_out[78][905],u_xpb_out[79][905],u_xpb_out[80][905],u_xpb_out[81][905],u_xpb_out[82][905],u_xpb_out[83][905],u_xpb_out[84][905],u_xpb_out[85][905],u_xpb_out[86][905],u_xpb_out[87][905],u_xpb_out[88][905],u_xpb_out[89][905],u_xpb_out[90][905],u_xpb_out[91][905],u_xpb_out[92][905],u_xpb_out[93][905],u_xpb_out[94][905],u_xpb_out[95][905],u_xpb_out[96][905],u_xpb_out[97][905],u_xpb_out[98][905],u_xpb_out[99][905],u_xpb_out[100][905],u_xpb_out[101][905],u_xpb_out[102][905],u_xpb_out[103][905],u_xpb_out[104][905],u_xpb_out[105][905]};

assign col_out_906 = {u_xpb_out[0][906],u_xpb_out[1][906],u_xpb_out[2][906],u_xpb_out[3][906],u_xpb_out[4][906],u_xpb_out[5][906],u_xpb_out[6][906],u_xpb_out[7][906],u_xpb_out[8][906],u_xpb_out[9][906],u_xpb_out[10][906],u_xpb_out[11][906],u_xpb_out[12][906],u_xpb_out[13][906],u_xpb_out[14][906],u_xpb_out[15][906],u_xpb_out[16][906],u_xpb_out[17][906],u_xpb_out[18][906],u_xpb_out[19][906],u_xpb_out[20][906],u_xpb_out[21][906],u_xpb_out[22][906],u_xpb_out[23][906],u_xpb_out[24][906],u_xpb_out[25][906],u_xpb_out[26][906],u_xpb_out[27][906],u_xpb_out[28][906],u_xpb_out[29][906],u_xpb_out[30][906],u_xpb_out[31][906],u_xpb_out[32][906],u_xpb_out[33][906],u_xpb_out[34][906],u_xpb_out[35][906],u_xpb_out[36][906],u_xpb_out[37][906],u_xpb_out[38][906],u_xpb_out[39][906],u_xpb_out[40][906],u_xpb_out[41][906],u_xpb_out[42][906],u_xpb_out[43][906],u_xpb_out[44][906],u_xpb_out[45][906],u_xpb_out[46][906],u_xpb_out[47][906],u_xpb_out[48][906],u_xpb_out[49][906],u_xpb_out[50][906],u_xpb_out[51][906],u_xpb_out[52][906],u_xpb_out[53][906],u_xpb_out[54][906],u_xpb_out[55][906],u_xpb_out[56][906],u_xpb_out[57][906],u_xpb_out[58][906],u_xpb_out[59][906],u_xpb_out[60][906],u_xpb_out[61][906],u_xpb_out[62][906],u_xpb_out[63][906],u_xpb_out[64][906],u_xpb_out[65][906],u_xpb_out[66][906],u_xpb_out[67][906],u_xpb_out[68][906],u_xpb_out[69][906],u_xpb_out[70][906],u_xpb_out[71][906],u_xpb_out[72][906],u_xpb_out[73][906],u_xpb_out[74][906],u_xpb_out[75][906],u_xpb_out[76][906],u_xpb_out[77][906],u_xpb_out[78][906],u_xpb_out[79][906],u_xpb_out[80][906],u_xpb_out[81][906],u_xpb_out[82][906],u_xpb_out[83][906],u_xpb_out[84][906],u_xpb_out[85][906],u_xpb_out[86][906],u_xpb_out[87][906],u_xpb_out[88][906],u_xpb_out[89][906],u_xpb_out[90][906],u_xpb_out[91][906],u_xpb_out[92][906],u_xpb_out[93][906],u_xpb_out[94][906],u_xpb_out[95][906],u_xpb_out[96][906],u_xpb_out[97][906],u_xpb_out[98][906],u_xpb_out[99][906],u_xpb_out[100][906],u_xpb_out[101][906],u_xpb_out[102][906],u_xpb_out[103][906],u_xpb_out[104][906],u_xpb_out[105][906]};

assign col_out_907 = {u_xpb_out[0][907],u_xpb_out[1][907],u_xpb_out[2][907],u_xpb_out[3][907],u_xpb_out[4][907],u_xpb_out[5][907],u_xpb_out[6][907],u_xpb_out[7][907],u_xpb_out[8][907],u_xpb_out[9][907],u_xpb_out[10][907],u_xpb_out[11][907],u_xpb_out[12][907],u_xpb_out[13][907],u_xpb_out[14][907],u_xpb_out[15][907],u_xpb_out[16][907],u_xpb_out[17][907],u_xpb_out[18][907],u_xpb_out[19][907],u_xpb_out[20][907],u_xpb_out[21][907],u_xpb_out[22][907],u_xpb_out[23][907],u_xpb_out[24][907],u_xpb_out[25][907],u_xpb_out[26][907],u_xpb_out[27][907],u_xpb_out[28][907],u_xpb_out[29][907],u_xpb_out[30][907],u_xpb_out[31][907],u_xpb_out[32][907],u_xpb_out[33][907],u_xpb_out[34][907],u_xpb_out[35][907],u_xpb_out[36][907],u_xpb_out[37][907],u_xpb_out[38][907],u_xpb_out[39][907],u_xpb_out[40][907],u_xpb_out[41][907],u_xpb_out[42][907],u_xpb_out[43][907],u_xpb_out[44][907],u_xpb_out[45][907],u_xpb_out[46][907],u_xpb_out[47][907],u_xpb_out[48][907],u_xpb_out[49][907],u_xpb_out[50][907],u_xpb_out[51][907],u_xpb_out[52][907],u_xpb_out[53][907],u_xpb_out[54][907],u_xpb_out[55][907],u_xpb_out[56][907],u_xpb_out[57][907],u_xpb_out[58][907],u_xpb_out[59][907],u_xpb_out[60][907],u_xpb_out[61][907],u_xpb_out[62][907],u_xpb_out[63][907],u_xpb_out[64][907],u_xpb_out[65][907],u_xpb_out[66][907],u_xpb_out[67][907],u_xpb_out[68][907],u_xpb_out[69][907],u_xpb_out[70][907],u_xpb_out[71][907],u_xpb_out[72][907],u_xpb_out[73][907],u_xpb_out[74][907],u_xpb_out[75][907],u_xpb_out[76][907],u_xpb_out[77][907],u_xpb_out[78][907],u_xpb_out[79][907],u_xpb_out[80][907],u_xpb_out[81][907],u_xpb_out[82][907],u_xpb_out[83][907],u_xpb_out[84][907],u_xpb_out[85][907],u_xpb_out[86][907],u_xpb_out[87][907],u_xpb_out[88][907],u_xpb_out[89][907],u_xpb_out[90][907],u_xpb_out[91][907],u_xpb_out[92][907],u_xpb_out[93][907],u_xpb_out[94][907],u_xpb_out[95][907],u_xpb_out[96][907],u_xpb_out[97][907],u_xpb_out[98][907],u_xpb_out[99][907],u_xpb_out[100][907],u_xpb_out[101][907],u_xpb_out[102][907],u_xpb_out[103][907],u_xpb_out[104][907],u_xpb_out[105][907]};

assign col_out_908 = {u_xpb_out[0][908],u_xpb_out[1][908],u_xpb_out[2][908],u_xpb_out[3][908],u_xpb_out[4][908],u_xpb_out[5][908],u_xpb_out[6][908],u_xpb_out[7][908],u_xpb_out[8][908],u_xpb_out[9][908],u_xpb_out[10][908],u_xpb_out[11][908],u_xpb_out[12][908],u_xpb_out[13][908],u_xpb_out[14][908],u_xpb_out[15][908],u_xpb_out[16][908],u_xpb_out[17][908],u_xpb_out[18][908],u_xpb_out[19][908],u_xpb_out[20][908],u_xpb_out[21][908],u_xpb_out[22][908],u_xpb_out[23][908],u_xpb_out[24][908],u_xpb_out[25][908],u_xpb_out[26][908],u_xpb_out[27][908],u_xpb_out[28][908],u_xpb_out[29][908],u_xpb_out[30][908],u_xpb_out[31][908],u_xpb_out[32][908],u_xpb_out[33][908],u_xpb_out[34][908],u_xpb_out[35][908],u_xpb_out[36][908],u_xpb_out[37][908],u_xpb_out[38][908],u_xpb_out[39][908],u_xpb_out[40][908],u_xpb_out[41][908],u_xpb_out[42][908],u_xpb_out[43][908],u_xpb_out[44][908],u_xpb_out[45][908],u_xpb_out[46][908],u_xpb_out[47][908],u_xpb_out[48][908],u_xpb_out[49][908],u_xpb_out[50][908],u_xpb_out[51][908],u_xpb_out[52][908],u_xpb_out[53][908],u_xpb_out[54][908],u_xpb_out[55][908],u_xpb_out[56][908],u_xpb_out[57][908],u_xpb_out[58][908],u_xpb_out[59][908],u_xpb_out[60][908],u_xpb_out[61][908],u_xpb_out[62][908],u_xpb_out[63][908],u_xpb_out[64][908],u_xpb_out[65][908],u_xpb_out[66][908],u_xpb_out[67][908],u_xpb_out[68][908],u_xpb_out[69][908],u_xpb_out[70][908],u_xpb_out[71][908],u_xpb_out[72][908],u_xpb_out[73][908],u_xpb_out[74][908],u_xpb_out[75][908],u_xpb_out[76][908],u_xpb_out[77][908],u_xpb_out[78][908],u_xpb_out[79][908],u_xpb_out[80][908],u_xpb_out[81][908],u_xpb_out[82][908],u_xpb_out[83][908],u_xpb_out[84][908],u_xpb_out[85][908],u_xpb_out[86][908],u_xpb_out[87][908],u_xpb_out[88][908],u_xpb_out[89][908],u_xpb_out[90][908],u_xpb_out[91][908],u_xpb_out[92][908],u_xpb_out[93][908],u_xpb_out[94][908],u_xpb_out[95][908],u_xpb_out[96][908],u_xpb_out[97][908],u_xpb_out[98][908],u_xpb_out[99][908],u_xpb_out[100][908],u_xpb_out[101][908],u_xpb_out[102][908],u_xpb_out[103][908],u_xpb_out[104][908],u_xpb_out[105][908]};

assign col_out_909 = {u_xpb_out[0][909],u_xpb_out[1][909],u_xpb_out[2][909],u_xpb_out[3][909],u_xpb_out[4][909],u_xpb_out[5][909],u_xpb_out[6][909],u_xpb_out[7][909],u_xpb_out[8][909],u_xpb_out[9][909],u_xpb_out[10][909],u_xpb_out[11][909],u_xpb_out[12][909],u_xpb_out[13][909],u_xpb_out[14][909],u_xpb_out[15][909],u_xpb_out[16][909],u_xpb_out[17][909],u_xpb_out[18][909],u_xpb_out[19][909],u_xpb_out[20][909],u_xpb_out[21][909],u_xpb_out[22][909],u_xpb_out[23][909],u_xpb_out[24][909],u_xpb_out[25][909],u_xpb_out[26][909],u_xpb_out[27][909],u_xpb_out[28][909],u_xpb_out[29][909],u_xpb_out[30][909],u_xpb_out[31][909],u_xpb_out[32][909],u_xpb_out[33][909],u_xpb_out[34][909],u_xpb_out[35][909],u_xpb_out[36][909],u_xpb_out[37][909],u_xpb_out[38][909],u_xpb_out[39][909],u_xpb_out[40][909],u_xpb_out[41][909],u_xpb_out[42][909],u_xpb_out[43][909],u_xpb_out[44][909],u_xpb_out[45][909],u_xpb_out[46][909],u_xpb_out[47][909],u_xpb_out[48][909],u_xpb_out[49][909],u_xpb_out[50][909],u_xpb_out[51][909],u_xpb_out[52][909],u_xpb_out[53][909],u_xpb_out[54][909],u_xpb_out[55][909],u_xpb_out[56][909],u_xpb_out[57][909],u_xpb_out[58][909],u_xpb_out[59][909],u_xpb_out[60][909],u_xpb_out[61][909],u_xpb_out[62][909],u_xpb_out[63][909],u_xpb_out[64][909],u_xpb_out[65][909],u_xpb_out[66][909],u_xpb_out[67][909],u_xpb_out[68][909],u_xpb_out[69][909],u_xpb_out[70][909],u_xpb_out[71][909],u_xpb_out[72][909],u_xpb_out[73][909],u_xpb_out[74][909],u_xpb_out[75][909],u_xpb_out[76][909],u_xpb_out[77][909],u_xpb_out[78][909],u_xpb_out[79][909],u_xpb_out[80][909],u_xpb_out[81][909],u_xpb_out[82][909],u_xpb_out[83][909],u_xpb_out[84][909],u_xpb_out[85][909],u_xpb_out[86][909],u_xpb_out[87][909],u_xpb_out[88][909],u_xpb_out[89][909],u_xpb_out[90][909],u_xpb_out[91][909],u_xpb_out[92][909],u_xpb_out[93][909],u_xpb_out[94][909],u_xpb_out[95][909],u_xpb_out[96][909],u_xpb_out[97][909],u_xpb_out[98][909],u_xpb_out[99][909],u_xpb_out[100][909],u_xpb_out[101][909],u_xpb_out[102][909],u_xpb_out[103][909],u_xpb_out[104][909],u_xpb_out[105][909]};

assign col_out_910 = {u_xpb_out[0][910],u_xpb_out[1][910],u_xpb_out[2][910],u_xpb_out[3][910],u_xpb_out[4][910],u_xpb_out[5][910],u_xpb_out[6][910],u_xpb_out[7][910],u_xpb_out[8][910],u_xpb_out[9][910],u_xpb_out[10][910],u_xpb_out[11][910],u_xpb_out[12][910],u_xpb_out[13][910],u_xpb_out[14][910],u_xpb_out[15][910],u_xpb_out[16][910],u_xpb_out[17][910],u_xpb_out[18][910],u_xpb_out[19][910],u_xpb_out[20][910],u_xpb_out[21][910],u_xpb_out[22][910],u_xpb_out[23][910],u_xpb_out[24][910],u_xpb_out[25][910],u_xpb_out[26][910],u_xpb_out[27][910],u_xpb_out[28][910],u_xpb_out[29][910],u_xpb_out[30][910],u_xpb_out[31][910],u_xpb_out[32][910],u_xpb_out[33][910],u_xpb_out[34][910],u_xpb_out[35][910],u_xpb_out[36][910],u_xpb_out[37][910],u_xpb_out[38][910],u_xpb_out[39][910],u_xpb_out[40][910],u_xpb_out[41][910],u_xpb_out[42][910],u_xpb_out[43][910],u_xpb_out[44][910],u_xpb_out[45][910],u_xpb_out[46][910],u_xpb_out[47][910],u_xpb_out[48][910],u_xpb_out[49][910],u_xpb_out[50][910],u_xpb_out[51][910],u_xpb_out[52][910],u_xpb_out[53][910],u_xpb_out[54][910],u_xpb_out[55][910],u_xpb_out[56][910],u_xpb_out[57][910],u_xpb_out[58][910],u_xpb_out[59][910],u_xpb_out[60][910],u_xpb_out[61][910],u_xpb_out[62][910],u_xpb_out[63][910],u_xpb_out[64][910],u_xpb_out[65][910],u_xpb_out[66][910],u_xpb_out[67][910],u_xpb_out[68][910],u_xpb_out[69][910],u_xpb_out[70][910],u_xpb_out[71][910],u_xpb_out[72][910],u_xpb_out[73][910],u_xpb_out[74][910],u_xpb_out[75][910],u_xpb_out[76][910],u_xpb_out[77][910],u_xpb_out[78][910],u_xpb_out[79][910],u_xpb_out[80][910],u_xpb_out[81][910],u_xpb_out[82][910],u_xpb_out[83][910],u_xpb_out[84][910],u_xpb_out[85][910],u_xpb_out[86][910],u_xpb_out[87][910],u_xpb_out[88][910],u_xpb_out[89][910],u_xpb_out[90][910],u_xpb_out[91][910],u_xpb_out[92][910],u_xpb_out[93][910],u_xpb_out[94][910],u_xpb_out[95][910],u_xpb_out[96][910],u_xpb_out[97][910],u_xpb_out[98][910],u_xpb_out[99][910],u_xpb_out[100][910],u_xpb_out[101][910],u_xpb_out[102][910],u_xpb_out[103][910],u_xpb_out[104][910],u_xpb_out[105][910]};

assign col_out_911 = {u_xpb_out[0][911],u_xpb_out[1][911],u_xpb_out[2][911],u_xpb_out[3][911],u_xpb_out[4][911],u_xpb_out[5][911],u_xpb_out[6][911],u_xpb_out[7][911],u_xpb_out[8][911],u_xpb_out[9][911],u_xpb_out[10][911],u_xpb_out[11][911],u_xpb_out[12][911],u_xpb_out[13][911],u_xpb_out[14][911],u_xpb_out[15][911],u_xpb_out[16][911],u_xpb_out[17][911],u_xpb_out[18][911],u_xpb_out[19][911],u_xpb_out[20][911],u_xpb_out[21][911],u_xpb_out[22][911],u_xpb_out[23][911],u_xpb_out[24][911],u_xpb_out[25][911],u_xpb_out[26][911],u_xpb_out[27][911],u_xpb_out[28][911],u_xpb_out[29][911],u_xpb_out[30][911],u_xpb_out[31][911],u_xpb_out[32][911],u_xpb_out[33][911],u_xpb_out[34][911],u_xpb_out[35][911],u_xpb_out[36][911],u_xpb_out[37][911],u_xpb_out[38][911],u_xpb_out[39][911],u_xpb_out[40][911],u_xpb_out[41][911],u_xpb_out[42][911],u_xpb_out[43][911],u_xpb_out[44][911],u_xpb_out[45][911],u_xpb_out[46][911],u_xpb_out[47][911],u_xpb_out[48][911],u_xpb_out[49][911],u_xpb_out[50][911],u_xpb_out[51][911],u_xpb_out[52][911],u_xpb_out[53][911],u_xpb_out[54][911],u_xpb_out[55][911],u_xpb_out[56][911],u_xpb_out[57][911],u_xpb_out[58][911],u_xpb_out[59][911],u_xpb_out[60][911],u_xpb_out[61][911],u_xpb_out[62][911],u_xpb_out[63][911],u_xpb_out[64][911],u_xpb_out[65][911],u_xpb_out[66][911],u_xpb_out[67][911],u_xpb_out[68][911],u_xpb_out[69][911],u_xpb_out[70][911],u_xpb_out[71][911],u_xpb_out[72][911],u_xpb_out[73][911],u_xpb_out[74][911],u_xpb_out[75][911],u_xpb_out[76][911],u_xpb_out[77][911],u_xpb_out[78][911],u_xpb_out[79][911],u_xpb_out[80][911],u_xpb_out[81][911],u_xpb_out[82][911],u_xpb_out[83][911],u_xpb_out[84][911],u_xpb_out[85][911],u_xpb_out[86][911],u_xpb_out[87][911],u_xpb_out[88][911],u_xpb_out[89][911],u_xpb_out[90][911],u_xpb_out[91][911],u_xpb_out[92][911],u_xpb_out[93][911],u_xpb_out[94][911],u_xpb_out[95][911],u_xpb_out[96][911],u_xpb_out[97][911],u_xpb_out[98][911],u_xpb_out[99][911],u_xpb_out[100][911],u_xpb_out[101][911],u_xpb_out[102][911],u_xpb_out[103][911],u_xpb_out[104][911],u_xpb_out[105][911]};

assign col_out_912 = {u_xpb_out[0][912],u_xpb_out[1][912],u_xpb_out[2][912],u_xpb_out[3][912],u_xpb_out[4][912],u_xpb_out[5][912],u_xpb_out[6][912],u_xpb_out[7][912],u_xpb_out[8][912],u_xpb_out[9][912],u_xpb_out[10][912],u_xpb_out[11][912],u_xpb_out[12][912],u_xpb_out[13][912],u_xpb_out[14][912],u_xpb_out[15][912],u_xpb_out[16][912],u_xpb_out[17][912],u_xpb_out[18][912],u_xpb_out[19][912],u_xpb_out[20][912],u_xpb_out[21][912],u_xpb_out[22][912],u_xpb_out[23][912],u_xpb_out[24][912],u_xpb_out[25][912],u_xpb_out[26][912],u_xpb_out[27][912],u_xpb_out[28][912],u_xpb_out[29][912],u_xpb_out[30][912],u_xpb_out[31][912],u_xpb_out[32][912],u_xpb_out[33][912],u_xpb_out[34][912],u_xpb_out[35][912],u_xpb_out[36][912],u_xpb_out[37][912],u_xpb_out[38][912],u_xpb_out[39][912],u_xpb_out[40][912],u_xpb_out[41][912],u_xpb_out[42][912],u_xpb_out[43][912],u_xpb_out[44][912],u_xpb_out[45][912],u_xpb_out[46][912],u_xpb_out[47][912],u_xpb_out[48][912],u_xpb_out[49][912],u_xpb_out[50][912],u_xpb_out[51][912],u_xpb_out[52][912],u_xpb_out[53][912],u_xpb_out[54][912],u_xpb_out[55][912],u_xpb_out[56][912],u_xpb_out[57][912],u_xpb_out[58][912],u_xpb_out[59][912],u_xpb_out[60][912],u_xpb_out[61][912],u_xpb_out[62][912],u_xpb_out[63][912],u_xpb_out[64][912],u_xpb_out[65][912],u_xpb_out[66][912],u_xpb_out[67][912],u_xpb_out[68][912],u_xpb_out[69][912],u_xpb_out[70][912],u_xpb_out[71][912],u_xpb_out[72][912],u_xpb_out[73][912],u_xpb_out[74][912],u_xpb_out[75][912],u_xpb_out[76][912],u_xpb_out[77][912],u_xpb_out[78][912],u_xpb_out[79][912],u_xpb_out[80][912],u_xpb_out[81][912],u_xpb_out[82][912],u_xpb_out[83][912],u_xpb_out[84][912],u_xpb_out[85][912],u_xpb_out[86][912],u_xpb_out[87][912],u_xpb_out[88][912],u_xpb_out[89][912],u_xpb_out[90][912],u_xpb_out[91][912],u_xpb_out[92][912],u_xpb_out[93][912],u_xpb_out[94][912],u_xpb_out[95][912],u_xpb_out[96][912],u_xpb_out[97][912],u_xpb_out[98][912],u_xpb_out[99][912],u_xpb_out[100][912],u_xpb_out[101][912],u_xpb_out[102][912],u_xpb_out[103][912],u_xpb_out[104][912],u_xpb_out[105][912]};

assign col_out_913 = {u_xpb_out[0][913],u_xpb_out[1][913],u_xpb_out[2][913],u_xpb_out[3][913],u_xpb_out[4][913],u_xpb_out[5][913],u_xpb_out[6][913],u_xpb_out[7][913],u_xpb_out[8][913],u_xpb_out[9][913],u_xpb_out[10][913],u_xpb_out[11][913],u_xpb_out[12][913],u_xpb_out[13][913],u_xpb_out[14][913],u_xpb_out[15][913],u_xpb_out[16][913],u_xpb_out[17][913],u_xpb_out[18][913],u_xpb_out[19][913],u_xpb_out[20][913],u_xpb_out[21][913],u_xpb_out[22][913],u_xpb_out[23][913],u_xpb_out[24][913],u_xpb_out[25][913],u_xpb_out[26][913],u_xpb_out[27][913],u_xpb_out[28][913],u_xpb_out[29][913],u_xpb_out[30][913],u_xpb_out[31][913],u_xpb_out[32][913],u_xpb_out[33][913],u_xpb_out[34][913],u_xpb_out[35][913],u_xpb_out[36][913],u_xpb_out[37][913],u_xpb_out[38][913],u_xpb_out[39][913],u_xpb_out[40][913],u_xpb_out[41][913],u_xpb_out[42][913],u_xpb_out[43][913],u_xpb_out[44][913],u_xpb_out[45][913],u_xpb_out[46][913],u_xpb_out[47][913],u_xpb_out[48][913],u_xpb_out[49][913],u_xpb_out[50][913],u_xpb_out[51][913],u_xpb_out[52][913],u_xpb_out[53][913],u_xpb_out[54][913],u_xpb_out[55][913],u_xpb_out[56][913],u_xpb_out[57][913],u_xpb_out[58][913],u_xpb_out[59][913],u_xpb_out[60][913],u_xpb_out[61][913],u_xpb_out[62][913],u_xpb_out[63][913],u_xpb_out[64][913],u_xpb_out[65][913],u_xpb_out[66][913],u_xpb_out[67][913],u_xpb_out[68][913],u_xpb_out[69][913],u_xpb_out[70][913],u_xpb_out[71][913],u_xpb_out[72][913],u_xpb_out[73][913],u_xpb_out[74][913],u_xpb_out[75][913],u_xpb_out[76][913],u_xpb_out[77][913],u_xpb_out[78][913],u_xpb_out[79][913],u_xpb_out[80][913],u_xpb_out[81][913],u_xpb_out[82][913],u_xpb_out[83][913],u_xpb_out[84][913],u_xpb_out[85][913],u_xpb_out[86][913],u_xpb_out[87][913],u_xpb_out[88][913],u_xpb_out[89][913],u_xpb_out[90][913],u_xpb_out[91][913],u_xpb_out[92][913],u_xpb_out[93][913],u_xpb_out[94][913],u_xpb_out[95][913],u_xpb_out[96][913],u_xpb_out[97][913],u_xpb_out[98][913],u_xpb_out[99][913],u_xpb_out[100][913],u_xpb_out[101][913],u_xpb_out[102][913],u_xpb_out[103][913],u_xpb_out[104][913],u_xpb_out[105][913]};

assign col_out_914 = {u_xpb_out[0][914],u_xpb_out[1][914],u_xpb_out[2][914],u_xpb_out[3][914],u_xpb_out[4][914],u_xpb_out[5][914],u_xpb_out[6][914],u_xpb_out[7][914],u_xpb_out[8][914],u_xpb_out[9][914],u_xpb_out[10][914],u_xpb_out[11][914],u_xpb_out[12][914],u_xpb_out[13][914],u_xpb_out[14][914],u_xpb_out[15][914],u_xpb_out[16][914],u_xpb_out[17][914],u_xpb_out[18][914],u_xpb_out[19][914],u_xpb_out[20][914],u_xpb_out[21][914],u_xpb_out[22][914],u_xpb_out[23][914],u_xpb_out[24][914],u_xpb_out[25][914],u_xpb_out[26][914],u_xpb_out[27][914],u_xpb_out[28][914],u_xpb_out[29][914],u_xpb_out[30][914],u_xpb_out[31][914],u_xpb_out[32][914],u_xpb_out[33][914],u_xpb_out[34][914],u_xpb_out[35][914],u_xpb_out[36][914],u_xpb_out[37][914],u_xpb_out[38][914],u_xpb_out[39][914],u_xpb_out[40][914],u_xpb_out[41][914],u_xpb_out[42][914],u_xpb_out[43][914],u_xpb_out[44][914],u_xpb_out[45][914],u_xpb_out[46][914],u_xpb_out[47][914],u_xpb_out[48][914],u_xpb_out[49][914],u_xpb_out[50][914],u_xpb_out[51][914],u_xpb_out[52][914],u_xpb_out[53][914],u_xpb_out[54][914],u_xpb_out[55][914],u_xpb_out[56][914],u_xpb_out[57][914],u_xpb_out[58][914],u_xpb_out[59][914],u_xpb_out[60][914],u_xpb_out[61][914],u_xpb_out[62][914],u_xpb_out[63][914],u_xpb_out[64][914],u_xpb_out[65][914],u_xpb_out[66][914],u_xpb_out[67][914],u_xpb_out[68][914],u_xpb_out[69][914],u_xpb_out[70][914],u_xpb_out[71][914],u_xpb_out[72][914],u_xpb_out[73][914],u_xpb_out[74][914],u_xpb_out[75][914],u_xpb_out[76][914],u_xpb_out[77][914],u_xpb_out[78][914],u_xpb_out[79][914],u_xpb_out[80][914],u_xpb_out[81][914],u_xpb_out[82][914],u_xpb_out[83][914],u_xpb_out[84][914],u_xpb_out[85][914],u_xpb_out[86][914],u_xpb_out[87][914],u_xpb_out[88][914],u_xpb_out[89][914],u_xpb_out[90][914],u_xpb_out[91][914],u_xpb_out[92][914],u_xpb_out[93][914],u_xpb_out[94][914],u_xpb_out[95][914],u_xpb_out[96][914],u_xpb_out[97][914],u_xpb_out[98][914],u_xpb_out[99][914],u_xpb_out[100][914],u_xpb_out[101][914],u_xpb_out[102][914],u_xpb_out[103][914],u_xpb_out[104][914],u_xpb_out[105][914]};

assign col_out_915 = {u_xpb_out[0][915],u_xpb_out[1][915],u_xpb_out[2][915],u_xpb_out[3][915],u_xpb_out[4][915],u_xpb_out[5][915],u_xpb_out[6][915],u_xpb_out[7][915],u_xpb_out[8][915],u_xpb_out[9][915],u_xpb_out[10][915],u_xpb_out[11][915],u_xpb_out[12][915],u_xpb_out[13][915],u_xpb_out[14][915],u_xpb_out[15][915],u_xpb_out[16][915],u_xpb_out[17][915],u_xpb_out[18][915],u_xpb_out[19][915],u_xpb_out[20][915],u_xpb_out[21][915],u_xpb_out[22][915],u_xpb_out[23][915],u_xpb_out[24][915],u_xpb_out[25][915],u_xpb_out[26][915],u_xpb_out[27][915],u_xpb_out[28][915],u_xpb_out[29][915],u_xpb_out[30][915],u_xpb_out[31][915],u_xpb_out[32][915],u_xpb_out[33][915],u_xpb_out[34][915],u_xpb_out[35][915],u_xpb_out[36][915],u_xpb_out[37][915],u_xpb_out[38][915],u_xpb_out[39][915],u_xpb_out[40][915],u_xpb_out[41][915],u_xpb_out[42][915],u_xpb_out[43][915],u_xpb_out[44][915],u_xpb_out[45][915],u_xpb_out[46][915],u_xpb_out[47][915],u_xpb_out[48][915],u_xpb_out[49][915],u_xpb_out[50][915],u_xpb_out[51][915],u_xpb_out[52][915],u_xpb_out[53][915],u_xpb_out[54][915],u_xpb_out[55][915],u_xpb_out[56][915],u_xpb_out[57][915],u_xpb_out[58][915],u_xpb_out[59][915],u_xpb_out[60][915],u_xpb_out[61][915],u_xpb_out[62][915],u_xpb_out[63][915],u_xpb_out[64][915],u_xpb_out[65][915],u_xpb_out[66][915],u_xpb_out[67][915],u_xpb_out[68][915],u_xpb_out[69][915],u_xpb_out[70][915],u_xpb_out[71][915],u_xpb_out[72][915],u_xpb_out[73][915],u_xpb_out[74][915],u_xpb_out[75][915],u_xpb_out[76][915],u_xpb_out[77][915],u_xpb_out[78][915],u_xpb_out[79][915],u_xpb_out[80][915],u_xpb_out[81][915],u_xpb_out[82][915],u_xpb_out[83][915],u_xpb_out[84][915],u_xpb_out[85][915],u_xpb_out[86][915],u_xpb_out[87][915],u_xpb_out[88][915],u_xpb_out[89][915],u_xpb_out[90][915],u_xpb_out[91][915],u_xpb_out[92][915],u_xpb_out[93][915],u_xpb_out[94][915],u_xpb_out[95][915],u_xpb_out[96][915],u_xpb_out[97][915],u_xpb_out[98][915],u_xpb_out[99][915],u_xpb_out[100][915],u_xpb_out[101][915],u_xpb_out[102][915],u_xpb_out[103][915],u_xpb_out[104][915],u_xpb_out[105][915]};

assign col_out_916 = {u_xpb_out[0][916],u_xpb_out[1][916],u_xpb_out[2][916],u_xpb_out[3][916],u_xpb_out[4][916],u_xpb_out[5][916],u_xpb_out[6][916],u_xpb_out[7][916],u_xpb_out[8][916],u_xpb_out[9][916],u_xpb_out[10][916],u_xpb_out[11][916],u_xpb_out[12][916],u_xpb_out[13][916],u_xpb_out[14][916],u_xpb_out[15][916],u_xpb_out[16][916],u_xpb_out[17][916],u_xpb_out[18][916],u_xpb_out[19][916],u_xpb_out[20][916],u_xpb_out[21][916],u_xpb_out[22][916],u_xpb_out[23][916],u_xpb_out[24][916],u_xpb_out[25][916],u_xpb_out[26][916],u_xpb_out[27][916],u_xpb_out[28][916],u_xpb_out[29][916],u_xpb_out[30][916],u_xpb_out[31][916],u_xpb_out[32][916],u_xpb_out[33][916],u_xpb_out[34][916],u_xpb_out[35][916],u_xpb_out[36][916],u_xpb_out[37][916],u_xpb_out[38][916],u_xpb_out[39][916],u_xpb_out[40][916],u_xpb_out[41][916],u_xpb_out[42][916],u_xpb_out[43][916],u_xpb_out[44][916],u_xpb_out[45][916],u_xpb_out[46][916],u_xpb_out[47][916],u_xpb_out[48][916],u_xpb_out[49][916],u_xpb_out[50][916],u_xpb_out[51][916],u_xpb_out[52][916],u_xpb_out[53][916],u_xpb_out[54][916],u_xpb_out[55][916],u_xpb_out[56][916],u_xpb_out[57][916],u_xpb_out[58][916],u_xpb_out[59][916],u_xpb_out[60][916],u_xpb_out[61][916],u_xpb_out[62][916],u_xpb_out[63][916],u_xpb_out[64][916],u_xpb_out[65][916],u_xpb_out[66][916],u_xpb_out[67][916],u_xpb_out[68][916],u_xpb_out[69][916],u_xpb_out[70][916],u_xpb_out[71][916],u_xpb_out[72][916],u_xpb_out[73][916],u_xpb_out[74][916],u_xpb_out[75][916],u_xpb_out[76][916],u_xpb_out[77][916],u_xpb_out[78][916],u_xpb_out[79][916],u_xpb_out[80][916],u_xpb_out[81][916],u_xpb_out[82][916],u_xpb_out[83][916],u_xpb_out[84][916],u_xpb_out[85][916],u_xpb_out[86][916],u_xpb_out[87][916],u_xpb_out[88][916],u_xpb_out[89][916],u_xpb_out[90][916],u_xpb_out[91][916],u_xpb_out[92][916],u_xpb_out[93][916],u_xpb_out[94][916],u_xpb_out[95][916],u_xpb_out[96][916],u_xpb_out[97][916],u_xpb_out[98][916],u_xpb_out[99][916],u_xpb_out[100][916],u_xpb_out[101][916],u_xpb_out[102][916],u_xpb_out[103][916],u_xpb_out[104][916],u_xpb_out[105][916]};

assign col_out_917 = {u_xpb_out[0][917],u_xpb_out[1][917],u_xpb_out[2][917],u_xpb_out[3][917],u_xpb_out[4][917],u_xpb_out[5][917],u_xpb_out[6][917],u_xpb_out[7][917],u_xpb_out[8][917],u_xpb_out[9][917],u_xpb_out[10][917],u_xpb_out[11][917],u_xpb_out[12][917],u_xpb_out[13][917],u_xpb_out[14][917],u_xpb_out[15][917],u_xpb_out[16][917],u_xpb_out[17][917],u_xpb_out[18][917],u_xpb_out[19][917],u_xpb_out[20][917],u_xpb_out[21][917],u_xpb_out[22][917],u_xpb_out[23][917],u_xpb_out[24][917],u_xpb_out[25][917],u_xpb_out[26][917],u_xpb_out[27][917],u_xpb_out[28][917],u_xpb_out[29][917],u_xpb_out[30][917],u_xpb_out[31][917],u_xpb_out[32][917],u_xpb_out[33][917],u_xpb_out[34][917],u_xpb_out[35][917],u_xpb_out[36][917],u_xpb_out[37][917],u_xpb_out[38][917],u_xpb_out[39][917],u_xpb_out[40][917],u_xpb_out[41][917],u_xpb_out[42][917],u_xpb_out[43][917],u_xpb_out[44][917],u_xpb_out[45][917],u_xpb_out[46][917],u_xpb_out[47][917],u_xpb_out[48][917],u_xpb_out[49][917],u_xpb_out[50][917],u_xpb_out[51][917],u_xpb_out[52][917],u_xpb_out[53][917],u_xpb_out[54][917],u_xpb_out[55][917],u_xpb_out[56][917],u_xpb_out[57][917],u_xpb_out[58][917],u_xpb_out[59][917],u_xpb_out[60][917],u_xpb_out[61][917],u_xpb_out[62][917],u_xpb_out[63][917],u_xpb_out[64][917],u_xpb_out[65][917],u_xpb_out[66][917],u_xpb_out[67][917],u_xpb_out[68][917],u_xpb_out[69][917],u_xpb_out[70][917],u_xpb_out[71][917],u_xpb_out[72][917],u_xpb_out[73][917],u_xpb_out[74][917],u_xpb_out[75][917],u_xpb_out[76][917],u_xpb_out[77][917],u_xpb_out[78][917],u_xpb_out[79][917],u_xpb_out[80][917],u_xpb_out[81][917],u_xpb_out[82][917],u_xpb_out[83][917],u_xpb_out[84][917],u_xpb_out[85][917],u_xpb_out[86][917],u_xpb_out[87][917],u_xpb_out[88][917],u_xpb_out[89][917],u_xpb_out[90][917],u_xpb_out[91][917],u_xpb_out[92][917],u_xpb_out[93][917],u_xpb_out[94][917],u_xpb_out[95][917],u_xpb_out[96][917],u_xpb_out[97][917],u_xpb_out[98][917],u_xpb_out[99][917],u_xpb_out[100][917],u_xpb_out[101][917],u_xpb_out[102][917],u_xpb_out[103][917],u_xpb_out[104][917],u_xpb_out[105][917]};

assign col_out_918 = {u_xpb_out[0][918],u_xpb_out[1][918],u_xpb_out[2][918],u_xpb_out[3][918],u_xpb_out[4][918],u_xpb_out[5][918],u_xpb_out[6][918],u_xpb_out[7][918],u_xpb_out[8][918],u_xpb_out[9][918],u_xpb_out[10][918],u_xpb_out[11][918],u_xpb_out[12][918],u_xpb_out[13][918],u_xpb_out[14][918],u_xpb_out[15][918],u_xpb_out[16][918],u_xpb_out[17][918],u_xpb_out[18][918],u_xpb_out[19][918],u_xpb_out[20][918],u_xpb_out[21][918],u_xpb_out[22][918],u_xpb_out[23][918],u_xpb_out[24][918],u_xpb_out[25][918],u_xpb_out[26][918],u_xpb_out[27][918],u_xpb_out[28][918],u_xpb_out[29][918],u_xpb_out[30][918],u_xpb_out[31][918],u_xpb_out[32][918],u_xpb_out[33][918],u_xpb_out[34][918],u_xpb_out[35][918],u_xpb_out[36][918],u_xpb_out[37][918],u_xpb_out[38][918],u_xpb_out[39][918],u_xpb_out[40][918],u_xpb_out[41][918],u_xpb_out[42][918],u_xpb_out[43][918],u_xpb_out[44][918],u_xpb_out[45][918],u_xpb_out[46][918],u_xpb_out[47][918],u_xpb_out[48][918],u_xpb_out[49][918],u_xpb_out[50][918],u_xpb_out[51][918],u_xpb_out[52][918],u_xpb_out[53][918],u_xpb_out[54][918],u_xpb_out[55][918],u_xpb_out[56][918],u_xpb_out[57][918],u_xpb_out[58][918],u_xpb_out[59][918],u_xpb_out[60][918],u_xpb_out[61][918],u_xpb_out[62][918],u_xpb_out[63][918],u_xpb_out[64][918],u_xpb_out[65][918],u_xpb_out[66][918],u_xpb_out[67][918],u_xpb_out[68][918],u_xpb_out[69][918],u_xpb_out[70][918],u_xpb_out[71][918],u_xpb_out[72][918],u_xpb_out[73][918],u_xpb_out[74][918],u_xpb_out[75][918],u_xpb_out[76][918],u_xpb_out[77][918],u_xpb_out[78][918],u_xpb_out[79][918],u_xpb_out[80][918],u_xpb_out[81][918],u_xpb_out[82][918],u_xpb_out[83][918],u_xpb_out[84][918],u_xpb_out[85][918],u_xpb_out[86][918],u_xpb_out[87][918],u_xpb_out[88][918],u_xpb_out[89][918],u_xpb_out[90][918],u_xpb_out[91][918],u_xpb_out[92][918],u_xpb_out[93][918],u_xpb_out[94][918],u_xpb_out[95][918],u_xpb_out[96][918],u_xpb_out[97][918],u_xpb_out[98][918],u_xpb_out[99][918],u_xpb_out[100][918],u_xpb_out[101][918],u_xpb_out[102][918],u_xpb_out[103][918],u_xpb_out[104][918],u_xpb_out[105][918]};

assign col_out_919 = {u_xpb_out[0][919],u_xpb_out[1][919],u_xpb_out[2][919],u_xpb_out[3][919],u_xpb_out[4][919],u_xpb_out[5][919],u_xpb_out[6][919],u_xpb_out[7][919],u_xpb_out[8][919],u_xpb_out[9][919],u_xpb_out[10][919],u_xpb_out[11][919],u_xpb_out[12][919],u_xpb_out[13][919],u_xpb_out[14][919],u_xpb_out[15][919],u_xpb_out[16][919],u_xpb_out[17][919],u_xpb_out[18][919],u_xpb_out[19][919],u_xpb_out[20][919],u_xpb_out[21][919],u_xpb_out[22][919],u_xpb_out[23][919],u_xpb_out[24][919],u_xpb_out[25][919],u_xpb_out[26][919],u_xpb_out[27][919],u_xpb_out[28][919],u_xpb_out[29][919],u_xpb_out[30][919],u_xpb_out[31][919],u_xpb_out[32][919],u_xpb_out[33][919],u_xpb_out[34][919],u_xpb_out[35][919],u_xpb_out[36][919],u_xpb_out[37][919],u_xpb_out[38][919],u_xpb_out[39][919],u_xpb_out[40][919],u_xpb_out[41][919],u_xpb_out[42][919],u_xpb_out[43][919],u_xpb_out[44][919],u_xpb_out[45][919],u_xpb_out[46][919],u_xpb_out[47][919],u_xpb_out[48][919],u_xpb_out[49][919],u_xpb_out[50][919],u_xpb_out[51][919],u_xpb_out[52][919],u_xpb_out[53][919],u_xpb_out[54][919],u_xpb_out[55][919],u_xpb_out[56][919],u_xpb_out[57][919],u_xpb_out[58][919],u_xpb_out[59][919],u_xpb_out[60][919],u_xpb_out[61][919],u_xpb_out[62][919],u_xpb_out[63][919],u_xpb_out[64][919],u_xpb_out[65][919],u_xpb_out[66][919],u_xpb_out[67][919],u_xpb_out[68][919],u_xpb_out[69][919],u_xpb_out[70][919],u_xpb_out[71][919],u_xpb_out[72][919],u_xpb_out[73][919],u_xpb_out[74][919],u_xpb_out[75][919],u_xpb_out[76][919],u_xpb_out[77][919],u_xpb_out[78][919],u_xpb_out[79][919],u_xpb_out[80][919],u_xpb_out[81][919],u_xpb_out[82][919],u_xpb_out[83][919],u_xpb_out[84][919],u_xpb_out[85][919],u_xpb_out[86][919],u_xpb_out[87][919],u_xpb_out[88][919],u_xpb_out[89][919],u_xpb_out[90][919],u_xpb_out[91][919],u_xpb_out[92][919],u_xpb_out[93][919],u_xpb_out[94][919],u_xpb_out[95][919],u_xpb_out[96][919],u_xpb_out[97][919],u_xpb_out[98][919],u_xpb_out[99][919],u_xpb_out[100][919],u_xpb_out[101][919],u_xpb_out[102][919],u_xpb_out[103][919],u_xpb_out[104][919],u_xpb_out[105][919]};

assign col_out_920 = {u_xpb_out[0][920],u_xpb_out[1][920],u_xpb_out[2][920],u_xpb_out[3][920],u_xpb_out[4][920],u_xpb_out[5][920],u_xpb_out[6][920],u_xpb_out[7][920],u_xpb_out[8][920],u_xpb_out[9][920],u_xpb_out[10][920],u_xpb_out[11][920],u_xpb_out[12][920],u_xpb_out[13][920],u_xpb_out[14][920],u_xpb_out[15][920],u_xpb_out[16][920],u_xpb_out[17][920],u_xpb_out[18][920],u_xpb_out[19][920],u_xpb_out[20][920],u_xpb_out[21][920],u_xpb_out[22][920],u_xpb_out[23][920],u_xpb_out[24][920],u_xpb_out[25][920],u_xpb_out[26][920],u_xpb_out[27][920],u_xpb_out[28][920],u_xpb_out[29][920],u_xpb_out[30][920],u_xpb_out[31][920],u_xpb_out[32][920],u_xpb_out[33][920],u_xpb_out[34][920],u_xpb_out[35][920],u_xpb_out[36][920],u_xpb_out[37][920],u_xpb_out[38][920],u_xpb_out[39][920],u_xpb_out[40][920],u_xpb_out[41][920],u_xpb_out[42][920],u_xpb_out[43][920],u_xpb_out[44][920],u_xpb_out[45][920],u_xpb_out[46][920],u_xpb_out[47][920],u_xpb_out[48][920],u_xpb_out[49][920],u_xpb_out[50][920],u_xpb_out[51][920],u_xpb_out[52][920],u_xpb_out[53][920],u_xpb_out[54][920],u_xpb_out[55][920],u_xpb_out[56][920],u_xpb_out[57][920],u_xpb_out[58][920],u_xpb_out[59][920],u_xpb_out[60][920],u_xpb_out[61][920],u_xpb_out[62][920],u_xpb_out[63][920],u_xpb_out[64][920],u_xpb_out[65][920],u_xpb_out[66][920],u_xpb_out[67][920],u_xpb_out[68][920],u_xpb_out[69][920],u_xpb_out[70][920],u_xpb_out[71][920],u_xpb_out[72][920],u_xpb_out[73][920],u_xpb_out[74][920],u_xpb_out[75][920],u_xpb_out[76][920],u_xpb_out[77][920],u_xpb_out[78][920],u_xpb_out[79][920],u_xpb_out[80][920],u_xpb_out[81][920],u_xpb_out[82][920],u_xpb_out[83][920],u_xpb_out[84][920],u_xpb_out[85][920],u_xpb_out[86][920],u_xpb_out[87][920],u_xpb_out[88][920],u_xpb_out[89][920],u_xpb_out[90][920],u_xpb_out[91][920],u_xpb_out[92][920],u_xpb_out[93][920],u_xpb_out[94][920],u_xpb_out[95][920],u_xpb_out[96][920],u_xpb_out[97][920],u_xpb_out[98][920],u_xpb_out[99][920],u_xpb_out[100][920],u_xpb_out[101][920],u_xpb_out[102][920],u_xpb_out[103][920],u_xpb_out[104][920],u_xpb_out[105][920]};

assign col_out_921 = {u_xpb_out[0][921],u_xpb_out[1][921],u_xpb_out[2][921],u_xpb_out[3][921],u_xpb_out[4][921],u_xpb_out[5][921],u_xpb_out[6][921],u_xpb_out[7][921],u_xpb_out[8][921],u_xpb_out[9][921],u_xpb_out[10][921],u_xpb_out[11][921],u_xpb_out[12][921],u_xpb_out[13][921],u_xpb_out[14][921],u_xpb_out[15][921],u_xpb_out[16][921],u_xpb_out[17][921],u_xpb_out[18][921],u_xpb_out[19][921],u_xpb_out[20][921],u_xpb_out[21][921],u_xpb_out[22][921],u_xpb_out[23][921],u_xpb_out[24][921],u_xpb_out[25][921],u_xpb_out[26][921],u_xpb_out[27][921],u_xpb_out[28][921],u_xpb_out[29][921],u_xpb_out[30][921],u_xpb_out[31][921],u_xpb_out[32][921],u_xpb_out[33][921],u_xpb_out[34][921],u_xpb_out[35][921],u_xpb_out[36][921],u_xpb_out[37][921],u_xpb_out[38][921],u_xpb_out[39][921],u_xpb_out[40][921],u_xpb_out[41][921],u_xpb_out[42][921],u_xpb_out[43][921],u_xpb_out[44][921],u_xpb_out[45][921],u_xpb_out[46][921],u_xpb_out[47][921],u_xpb_out[48][921],u_xpb_out[49][921],u_xpb_out[50][921],u_xpb_out[51][921],u_xpb_out[52][921],u_xpb_out[53][921],u_xpb_out[54][921],u_xpb_out[55][921],u_xpb_out[56][921],u_xpb_out[57][921],u_xpb_out[58][921],u_xpb_out[59][921],u_xpb_out[60][921],u_xpb_out[61][921],u_xpb_out[62][921],u_xpb_out[63][921],u_xpb_out[64][921],u_xpb_out[65][921],u_xpb_out[66][921],u_xpb_out[67][921],u_xpb_out[68][921],u_xpb_out[69][921],u_xpb_out[70][921],u_xpb_out[71][921],u_xpb_out[72][921],u_xpb_out[73][921],u_xpb_out[74][921],u_xpb_out[75][921],u_xpb_out[76][921],u_xpb_out[77][921],u_xpb_out[78][921],u_xpb_out[79][921],u_xpb_out[80][921],u_xpb_out[81][921],u_xpb_out[82][921],u_xpb_out[83][921],u_xpb_out[84][921],u_xpb_out[85][921],u_xpb_out[86][921],u_xpb_out[87][921],u_xpb_out[88][921],u_xpb_out[89][921],u_xpb_out[90][921],u_xpb_out[91][921],u_xpb_out[92][921],u_xpb_out[93][921],u_xpb_out[94][921],u_xpb_out[95][921],u_xpb_out[96][921],u_xpb_out[97][921],u_xpb_out[98][921],u_xpb_out[99][921],u_xpb_out[100][921],u_xpb_out[101][921],u_xpb_out[102][921],u_xpb_out[103][921],u_xpb_out[104][921],u_xpb_out[105][921]};

assign col_out_922 = {u_xpb_out[0][922],u_xpb_out[1][922],u_xpb_out[2][922],u_xpb_out[3][922],u_xpb_out[4][922],u_xpb_out[5][922],u_xpb_out[6][922],u_xpb_out[7][922],u_xpb_out[8][922],u_xpb_out[9][922],u_xpb_out[10][922],u_xpb_out[11][922],u_xpb_out[12][922],u_xpb_out[13][922],u_xpb_out[14][922],u_xpb_out[15][922],u_xpb_out[16][922],u_xpb_out[17][922],u_xpb_out[18][922],u_xpb_out[19][922],u_xpb_out[20][922],u_xpb_out[21][922],u_xpb_out[22][922],u_xpb_out[23][922],u_xpb_out[24][922],u_xpb_out[25][922],u_xpb_out[26][922],u_xpb_out[27][922],u_xpb_out[28][922],u_xpb_out[29][922],u_xpb_out[30][922],u_xpb_out[31][922],u_xpb_out[32][922],u_xpb_out[33][922],u_xpb_out[34][922],u_xpb_out[35][922],u_xpb_out[36][922],u_xpb_out[37][922],u_xpb_out[38][922],u_xpb_out[39][922],u_xpb_out[40][922],u_xpb_out[41][922],u_xpb_out[42][922],u_xpb_out[43][922],u_xpb_out[44][922],u_xpb_out[45][922],u_xpb_out[46][922],u_xpb_out[47][922],u_xpb_out[48][922],u_xpb_out[49][922],u_xpb_out[50][922],u_xpb_out[51][922],u_xpb_out[52][922],u_xpb_out[53][922],u_xpb_out[54][922],u_xpb_out[55][922],u_xpb_out[56][922],u_xpb_out[57][922],u_xpb_out[58][922],u_xpb_out[59][922],u_xpb_out[60][922],u_xpb_out[61][922],u_xpb_out[62][922],u_xpb_out[63][922],u_xpb_out[64][922],u_xpb_out[65][922],u_xpb_out[66][922],u_xpb_out[67][922],u_xpb_out[68][922],u_xpb_out[69][922],u_xpb_out[70][922],u_xpb_out[71][922],u_xpb_out[72][922],u_xpb_out[73][922],u_xpb_out[74][922],u_xpb_out[75][922],u_xpb_out[76][922],u_xpb_out[77][922],u_xpb_out[78][922],u_xpb_out[79][922],u_xpb_out[80][922],u_xpb_out[81][922],u_xpb_out[82][922],u_xpb_out[83][922],u_xpb_out[84][922],u_xpb_out[85][922],u_xpb_out[86][922],u_xpb_out[87][922],u_xpb_out[88][922],u_xpb_out[89][922],u_xpb_out[90][922],u_xpb_out[91][922],u_xpb_out[92][922],u_xpb_out[93][922],u_xpb_out[94][922],u_xpb_out[95][922],u_xpb_out[96][922],u_xpb_out[97][922],u_xpb_out[98][922],u_xpb_out[99][922],u_xpb_out[100][922],u_xpb_out[101][922],u_xpb_out[102][922],u_xpb_out[103][922],u_xpb_out[104][922],u_xpb_out[105][922]};

assign col_out_923 = {u_xpb_out[0][923],u_xpb_out[1][923],u_xpb_out[2][923],u_xpb_out[3][923],u_xpb_out[4][923],u_xpb_out[5][923],u_xpb_out[6][923],u_xpb_out[7][923],u_xpb_out[8][923],u_xpb_out[9][923],u_xpb_out[10][923],u_xpb_out[11][923],u_xpb_out[12][923],u_xpb_out[13][923],u_xpb_out[14][923],u_xpb_out[15][923],u_xpb_out[16][923],u_xpb_out[17][923],u_xpb_out[18][923],u_xpb_out[19][923],u_xpb_out[20][923],u_xpb_out[21][923],u_xpb_out[22][923],u_xpb_out[23][923],u_xpb_out[24][923],u_xpb_out[25][923],u_xpb_out[26][923],u_xpb_out[27][923],u_xpb_out[28][923],u_xpb_out[29][923],u_xpb_out[30][923],u_xpb_out[31][923],u_xpb_out[32][923],u_xpb_out[33][923],u_xpb_out[34][923],u_xpb_out[35][923],u_xpb_out[36][923],u_xpb_out[37][923],u_xpb_out[38][923],u_xpb_out[39][923],u_xpb_out[40][923],u_xpb_out[41][923],u_xpb_out[42][923],u_xpb_out[43][923],u_xpb_out[44][923],u_xpb_out[45][923],u_xpb_out[46][923],u_xpb_out[47][923],u_xpb_out[48][923],u_xpb_out[49][923],u_xpb_out[50][923],u_xpb_out[51][923],u_xpb_out[52][923],u_xpb_out[53][923],u_xpb_out[54][923],u_xpb_out[55][923],u_xpb_out[56][923],u_xpb_out[57][923],u_xpb_out[58][923],u_xpb_out[59][923],u_xpb_out[60][923],u_xpb_out[61][923],u_xpb_out[62][923],u_xpb_out[63][923],u_xpb_out[64][923],u_xpb_out[65][923],u_xpb_out[66][923],u_xpb_out[67][923],u_xpb_out[68][923],u_xpb_out[69][923],u_xpb_out[70][923],u_xpb_out[71][923],u_xpb_out[72][923],u_xpb_out[73][923],u_xpb_out[74][923],u_xpb_out[75][923],u_xpb_out[76][923],u_xpb_out[77][923],u_xpb_out[78][923],u_xpb_out[79][923],u_xpb_out[80][923],u_xpb_out[81][923],u_xpb_out[82][923],u_xpb_out[83][923],u_xpb_out[84][923],u_xpb_out[85][923],u_xpb_out[86][923],u_xpb_out[87][923],u_xpb_out[88][923],u_xpb_out[89][923],u_xpb_out[90][923],u_xpb_out[91][923],u_xpb_out[92][923],u_xpb_out[93][923],u_xpb_out[94][923],u_xpb_out[95][923],u_xpb_out[96][923],u_xpb_out[97][923],u_xpb_out[98][923],u_xpb_out[99][923],u_xpb_out[100][923],u_xpb_out[101][923],u_xpb_out[102][923],u_xpb_out[103][923],u_xpb_out[104][923],u_xpb_out[105][923]};

assign col_out_924 = {u_xpb_out[0][924],u_xpb_out[1][924],u_xpb_out[2][924],u_xpb_out[3][924],u_xpb_out[4][924],u_xpb_out[5][924],u_xpb_out[6][924],u_xpb_out[7][924],u_xpb_out[8][924],u_xpb_out[9][924],u_xpb_out[10][924],u_xpb_out[11][924],u_xpb_out[12][924],u_xpb_out[13][924],u_xpb_out[14][924],u_xpb_out[15][924],u_xpb_out[16][924],u_xpb_out[17][924],u_xpb_out[18][924],u_xpb_out[19][924],u_xpb_out[20][924],u_xpb_out[21][924],u_xpb_out[22][924],u_xpb_out[23][924],u_xpb_out[24][924],u_xpb_out[25][924],u_xpb_out[26][924],u_xpb_out[27][924],u_xpb_out[28][924],u_xpb_out[29][924],u_xpb_out[30][924],u_xpb_out[31][924],u_xpb_out[32][924],u_xpb_out[33][924],u_xpb_out[34][924],u_xpb_out[35][924],u_xpb_out[36][924],u_xpb_out[37][924],u_xpb_out[38][924],u_xpb_out[39][924],u_xpb_out[40][924],u_xpb_out[41][924],u_xpb_out[42][924],u_xpb_out[43][924],u_xpb_out[44][924],u_xpb_out[45][924],u_xpb_out[46][924],u_xpb_out[47][924],u_xpb_out[48][924],u_xpb_out[49][924],u_xpb_out[50][924],u_xpb_out[51][924],u_xpb_out[52][924],u_xpb_out[53][924],u_xpb_out[54][924],u_xpb_out[55][924],u_xpb_out[56][924],u_xpb_out[57][924],u_xpb_out[58][924],u_xpb_out[59][924],u_xpb_out[60][924],u_xpb_out[61][924],u_xpb_out[62][924],u_xpb_out[63][924],u_xpb_out[64][924],u_xpb_out[65][924],u_xpb_out[66][924],u_xpb_out[67][924],u_xpb_out[68][924],u_xpb_out[69][924],u_xpb_out[70][924],u_xpb_out[71][924],u_xpb_out[72][924],u_xpb_out[73][924],u_xpb_out[74][924],u_xpb_out[75][924],u_xpb_out[76][924],u_xpb_out[77][924],u_xpb_out[78][924],u_xpb_out[79][924],u_xpb_out[80][924],u_xpb_out[81][924],u_xpb_out[82][924],u_xpb_out[83][924],u_xpb_out[84][924],u_xpb_out[85][924],u_xpb_out[86][924],u_xpb_out[87][924],u_xpb_out[88][924],u_xpb_out[89][924],u_xpb_out[90][924],u_xpb_out[91][924],u_xpb_out[92][924],u_xpb_out[93][924],u_xpb_out[94][924],u_xpb_out[95][924],u_xpb_out[96][924],u_xpb_out[97][924],u_xpb_out[98][924],u_xpb_out[99][924],u_xpb_out[100][924],u_xpb_out[101][924],u_xpb_out[102][924],u_xpb_out[103][924],u_xpb_out[104][924],u_xpb_out[105][924]};

assign col_out_925 = {u_xpb_out[0][925],u_xpb_out[1][925],u_xpb_out[2][925],u_xpb_out[3][925],u_xpb_out[4][925],u_xpb_out[5][925],u_xpb_out[6][925],u_xpb_out[7][925],u_xpb_out[8][925],u_xpb_out[9][925],u_xpb_out[10][925],u_xpb_out[11][925],u_xpb_out[12][925],u_xpb_out[13][925],u_xpb_out[14][925],u_xpb_out[15][925],u_xpb_out[16][925],u_xpb_out[17][925],u_xpb_out[18][925],u_xpb_out[19][925],u_xpb_out[20][925],u_xpb_out[21][925],u_xpb_out[22][925],u_xpb_out[23][925],u_xpb_out[24][925],u_xpb_out[25][925],u_xpb_out[26][925],u_xpb_out[27][925],u_xpb_out[28][925],u_xpb_out[29][925],u_xpb_out[30][925],u_xpb_out[31][925],u_xpb_out[32][925],u_xpb_out[33][925],u_xpb_out[34][925],u_xpb_out[35][925],u_xpb_out[36][925],u_xpb_out[37][925],u_xpb_out[38][925],u_xpb_out[39][925],u_xpb_out[40][925],u_xpb_out[41][925],u_xpb_out[42][925],u_xpb_out[43][925],u_xpb_out[44][925],u_xpb_out[45][925],u_xpb_out[46][925],u_xpb_out[47][925],u_xpb_out[48][925],u_xpb_out[49][925],u_xpb_out[50][925],u_xpb_out[51][925],u_xpb_out[52][925],u_xpb_out[53][925],u_xpb_out[54][925],u_xpb_out[55][925],u_xpb_out[56][925],u_xpb_out[57][925],u_xpb_out[58][925],u_xpb_out[59][925],u_xpb_out[60][925],u_xpb_out[61][925],u_xpb_out[62][925],u_xpb_out[63][925],u_xpb_out[64][925],u_xpb_out[65][925],u_xpb_out[66][925],u_xpb_out[67][925],u_xpb_out[68][925],u_xpb_out[69][925],u_xpb_out[70][925],u_xpb_out[71][925],u_xpb_out[72][925],u_xpb_out[73][925],u_xpb_out[74][925],u_xpb_out[75][925],u_xpb_out[76][925],u_xpb_out[77][925],u_xpb_out[78][925],u_xpb_out[79][925],u_xpb_out[80][925],u_xpb_out[81][925],u_xpb_out[82][925],u_xpb_out[83][925],u_xpb_out[84][925],u_xpb_out[85][925],u_xpb_out[86][925],u_xpb_out[87][925],u_xpb_out[88][925],u_xpb_out[89][925],u_xpb_out[90][925],u_xpb_out[91][925],u_xpb_out[92][925],u_xpb_out[93][925],u_xpb_out[94][925],u_xpb_out[95][925],u_xpb_out[96][925],u_xpb_out[97][925],u_xpb_out[98][925],u_xpb_out[99][925],u_xpb_out[100][925],u_xpb_out[101][925],u_xpb_out[102][925],u_xpb_out[103][925],u_xpb_out[104][925],u_xpb_out[105][925]};

assign col_out_926 = {u_xpb_out[0][926],u_xpb_out[1][926],u_xpb_out[2][926],u_xpb_out[3][926],u_xpb_out[4][926],u_xpb_out[5][926],u_xpb_out[6][926],u_xpb_out[7][926],u_xpb_out[8][926],u_xpb_out[9][926],u_xpb_out[10][926],u_xpb_out[11][926],u_xpb_out[12][926],u_xpb_out[13][926],u_xpb_out[14][926],u_xpb_out[15][926],u_xpb_out[16][926],u_xpb_out[17][926],u_xpb_out[18][926],u_xpb_out[19][926],u_xpb_out[20][926],u_xpb_out[21][926],u_xpb_out[22][926],u_xpb_out[23][926],u_xpb_out[24][926],u_xpb_out[25][926],u_xpb_out[26][926],u_xpb_out[27][926],u_xpb_out[28][926],u_xpb_out[29][926],u_xpb_out[30][926],u_xpb_out[31][926],u_xpb_out[32][926],u_xpb_out[33][926],u_xpb_out[34][926],u_xpb_out[35][926],u_xpb_out[36][926],u_xpb_out[37][926],u_xpb_out[38][926],u_xpb_out[39][926],u_xpb_out[40][926],u_xpb_out[41][926],u_xpb_out[42][926],u_xpb_out[43][926],u_xpb_out[44][926],u_xpb_out[45][926],u_xpb_out[46][926],u_xpb_out[47][926],u_xpb_out[48][926],u_xpb_out[49][926],u_xpb_out[50][926],u_xpb_out[51][926],u_xpb_out[52][926],u_xpb_out[53][926],u_xpb_out[54][926],u_xpb_out[55][926],u_xpb_out[56][926],u_xpb_out[57][926],u_xpb_out[58][926],u_xpb_out[59][926],u_xpb_out[60][926],u_xpb_out[61][926],u_xpb_out[62][926],u_xpb_out[63][926],u_xpb_out[64][926],u_xpb_out[65][926],u_xpb_out[66][926],u_xpb_out[67][926],u_xpb_out[68][926],u_xpb_out[69][926],u_xpb_out[70][926],u_xpb_out[71][926],u_xpb_out[72][926],u_xpb_out[73][926],u_xpb_out[74][926],u_xpb_out[75][926],u_xpb_out[76][926],u_xpb_out[77][926],u_xpb_out[78][926],u_xpb_out[79][926],u_xpb_out[80][926],u_xpb_out[81][926],u_xpb_out[82][926],u_xpb_out[83][926],u_xpb_out[84][926],u_xpb_out[85][926],u_xpb_out[86][926],u_xpb_out[87][926],u_xpb_out[88][926],u_xpb_out[89][926],u_xpb_out[90][926],u_xpb_out[91][926],u_xpb_out[92][926],u_xpb_out[93][926],u_xpb_out[94][926],u_xpb_out[95][926],u_xpb_out[96][926],u_xpb_out[97][926],u_xpb_out[98][926],u_xpb_out[99][926],u_xpb_out[100][926],u_xpb_out[101][926],u_xpb_out[102][926],u_xpb_out[103][926],u_xpb_out[104][926],u_xpb_out[105][926]};

assign col_out_927 = {u_xpb_out[0][927],u_xpb_out[1][927],u_xpb_out[2][927],u_xpb_out[3][927],u_xpb_out[4][927],u_xpb_out[5][927],u_xpb_out[6][927],u_xpb_out[7][927],u_xpb_out[8][927],u_xpb_out[9][927],u_xpb_out[10][927],u_xpb_out[11][927],u_xpb_out[12][927],u_xpb_out[13][927],u_xpb_out[14][927],u_xpb_out[15][927],u_xpb_out[16][927],u_xpb_out[17][927],u_xpb_out[18][927],u_xpb_out[19][927],u_xpb_out[20][927],u_xpb_out[21][927],u_xpb_out[22][927],u_xpb_out[23][927],u_xpb_out[24][927],u_xpb_out[25][927],u_xpb_out[26][927],u_xpb_out[27][927],u_xpb_out[28][927],u_xpb_out[29][927],u_xpb_out[30][927],u_xpb_out[31][927],u_xpb_out[32][927],u_xpb_out[33][927],u_xpb_out[34][927],u_xpb_out[35][927],u_xpb_out[36][927],u_xpb_out[37][927],u_xpb_out[38][927],u_xpb_out[39][927],u_xpb_out[40][927],u_xpb_out[41][927],u_xpb_out[42][927],u_xpb_out[43][927],u_xpb_out[44][927],u_xpb_out[45][927],u_xpb_out[46][927],u_xpb_out[47][927],u_xpb_out[48][927],u_xpb_out[49][927],u_xpb_out[50][927],u_xpb_out[51][927],u_xpb_out[52][927],u_xpb_out[53][927],u_xpb_out[54][927],u_xpb_out[55][927],u_xpb_out[56][927],u_xpb_out[57][927],u_xpb_out[58][927],u_xpb_out[59][927],u_xpb_out[60][927],u_xpb_out[61][927],u_xpb_out[62][927],u_xpb_out[63][927],u_xpb_out[64][927],u_xpb_out[65][927],u_xpb_out[66][927],u_xpb_out[67][927],u_xpb_out[68][927],u_xpb_out[69][927],u_xpb_out[70][927],u_xpb_out[71][927],u_xpb_out[72][927],u_xpb_out[73][927],u_xpb_out[74][927],u_xpb_out[75][927],u_xpb_out[76][927],u_xpb_out[77][927],u_xpb_out[78][927],u_xpb_out[79][927],u_xpb_out[80][927],u_xpb_out[81][927],u_xpb_out[82][927],u_xpb_out[83][927],u_xpb_out[84][927],u_xpb_out[85][927],u_xpb_out[86][927],u_xpb_out[87][927],u_xpb_out[88][927],u_xpb_out[89][927],u_xpb_out[90][927],u_xpb_out[91][927],u_xpb_out[92][927],u_xpb_out[93][927],u_xpb_out[94][927],u_xpb_out[95][927],u_xpb_out[96][927],u_xpb_out[97][927],u_xpb_out[98][927],u_xpb_out[99][927],u_xpb_out[100][927],u_xpb_out[101][927],u_xpb_out[102][927],u_xpb_out[103][927],u_xpb_out[104][927],u_xpb_out[105][927]};

assign col_out_928 = {u_xpb_out[0][928],u_xpb_out[1][928],u_xpb_out[2][928],u_xpb_out[3][928],u_xpb_out[4][928],u_xpb_out[5][928],u_xpb_out[6][928],u_xpb_out[7][928],u_xpb_out[8][928],u_xpb_out[9][928],u_xpb_out[10][928],u_xpb_out[11][928],u_xpb_out[12][928],u_xpb_out[13][928],u_xpb_out[14][928],u_xpb_out[15][928],u_xpb_out[16][928],u_xpb_out[17][928],u_xpb_out[18][928],u_xpb_out[19][928],u_xpb_out[20][928],u_xpb_out[21][928],u_xpb_out[22][928],u_xpb_out[23][928],u_xpb_out[24][928],u_xpb_out[25][928],u_xpb_out[26][928],u_xpb_out[27][928],u_xpb_out[28][928],u_xpb_out[29][928],u_xpb_out[30][928],u_xpb_out[31][928],u_xpb_out[32][928],u_xpb_out[33][928],u_xpb_out[34][928],u_xpb_out[35][928],u_xpb_out[36][928],u_xpb_out[37][928],u_xpb_out[38][928],u_xpb_out[39][928],u_xpb_out[40][928],u_xpb_out[41][928],u_xpb_out[42][928],u_xpb_out[43][928],u_xpb_out[44][928],u_xpb_out[45][928],u_xpb_out[46][928],u_xpb_out[47][928],u_xpb_out[48][928],u_xpb_out[49][928],u_xpb_out[50][928],u_xpb_out[51][928],u_xpb_out[52][928],u_xpb_out[53][928],u_xpb_out[54][928],u_xpb_out[55][928],u_xpb_out[56][928],u_xpb_out[57][928],u_xpb_out[58][928],u_xpb_out[59][928],u_xpb_out[60][928],u_xpb_out[61][928],u_xpb_out[62][928],u_xpb_out[63][928],u_xpb_out[64][928],u_xpb_out[65][928],u_xpb_out[66][928],u_xpb_out[67][928],u_xpb_out[68][928],u_xpb_out[69][928],u_xpb_out[70][928],u_xpb_out[71][928],u_xpb_out[72][928],u_xpb_out[73][928],u_xpb_out[74][928],u_xpb_out[75][928],u_xpb_out[76][928],u_xpb_out[77][928],u_xpb_out[78][928],u_xpb_out[79][928],u_xpb_out[80][928],u_xpb_out[81][928],u_xpb_out[82][928],u_xpb_out[83][928],u_xpb_out[84][928],u_xpb_out[85][928],u_xpb_out[86][928],u_xpb_out[87][928],u_xpb_out[88][928],u_xpb_out[89][928],u_xpb_out[90][928],u_xpb_out[91][928],u_xpb_out[92][928],u_xpb_out[93][928],u_xpb_out[94][928],u_xpb_out[95][928],u_xpb_out[96][928],u_xpb_out[97][928],u_xpb_out[98][928],u_xpb_out[99][928],u_xpb_out[100][928],u_xpb_out[101][928],u_xpb_out[102][928],u_xpb_out[103][928],u_xpb_out[104][928],u_xpb_out[105][928]};

assign col_out_929 = {u_xpb_out[0][929],u_xpb_out[1][929],u_xpb_out[2][929],u_xpb_out[3][929],u_xpb_out[4][929],u_xpb_out[5][929],u_xpb_out[6][929],u_xpb_out[7][929],u_xpb_out[8][929],u_xpb_out[9][929],u_xpb_out[10][929],u_xpb_out[11][929],u_xpb_out[12][929],u_xpb_out[13][929],u_xpb_out[14][929],u_xpb_out[15][929],u_xpb_out[16][929],u_xpb_out[17][929],u_xpb_out[18][929],u_xpb_out[19][929],u_xpb_out[20][929],u_xpb_out[21][929],u_xpb_out[22][929],u_xpb_out[23][929],u_xpb_out[24][929],u_xpb_out[25][929],u_xpb_out[26][929],u_xpb_out[27][929],u_xpb_out[28][929],u_xpb_out[29][929],u_xpb_out[30][929],u_xpb_out[31][929],u_xpb_out[32][929],u_xpb_out[33][929],u_xpb_out[34][929],u_xpb_out[35][929],u_xpb_out[36][929],u_xpb_out[37][929],u_xpb_out[38][929],u_xpb_out[39][929],u_xpb_out[40][929],u_xpb_out[41][929],u_xpb_out[42][929],u_xpb_out[43][929],u_xpb_out[44][929],u_xpb_out[45][929],u_xpb_out[46][929],u_xpb_out[47][929],u_xpb_out[48][929],u_xpb_out[49][929],u_xpb_out[50][929],u_xpb_out[51][929],u_xpb_out[52][929],u_xpb_out[53][929],u_xpb_out[54][929],u_xpb_out[55][929],u_xpb_out[56][929],u_xpb_out[57][929],u_xpb_out[58][929],u_xpb_out[59][929],u_xpb_out[60][929],u_xpb_out[61][929],u_xpb_out[62][929],u_xpb_out[63][929],u_xpb_out[64][929],u_xpb_out[65][929],u_xpb_out[66][929],u_xpb_out[67][929],u_xpb_out[68][929],u_xpb_out[69][929],u_xpb_out[70][929],u_xpb_out[71][929],u_xpb_out[72][929],u_xpb_out[73][929],u_xpb_out[74][929],u_xpb_out[75][929],u_xpb_out[76][929],u_xpb_out[77][929],u_xpb_out[78][929],u_xpb_out[79][929],u_xpb_out[80][929],u_xpb_out[81][929],u_xpb_out[82][929],u_xpb_out[83][929],u_xpb_out[84][929],u_xpb_out[85][929],u_xpb_out[86][929],u_xpb_out[87][929],u_xpb_out[88][929],u_xpb_out[89][929],u_xpb_out[90][929],u_xpb_out[91][929],u_xpb_out[92][929],u_xpb_out[93][929],u_xpb_out[94][929],u_xpb_out[95][929],u_xpb_out[96][929],u_xpb_out[97][929],u_xpb_out[98][929],u_xpb_out[99][929],u_xpb_out[100][929],u_xpb_out[101][929],u_xpb_out[102][929],u_xpb_out[103][929],u_xpb_out[104][929],u_xpb_out[105][929]};

assign col_out_930 = {u_xpb_out[0][930],u_xpb_out[1][930],u_xpb_out[2][930],u_xpb_out[3][930],u_xpb_out[4][930],u_xpb_out[5][930],u_xpb_out[6][930],u_xpb_out[7][930],u_xpb_out[8][930],u_xpb_out[9][930],u_xpb_out[10][930],u_xpb_out[11][930],u_xpb_out[12][930],u_xpb_out[13][930],u_xpb_out[14][930],u_xpb_out[15][930],u_xpb_out[16][930],u_xpb_out[17][930],u_xpb_out[18][930],u_xpb_out[19][930],u_xpb_out[20][930],u_xpb_out[21][930],u_xpb_out[22][930],u_xpb_out[23][930],u_xpb_out[24][930],u_xpb_out[25][930],u_xpb_out[26][930],u_xpb_out[27][930],u_xpb_out[28][930],u_xpb_out[29][930],u_xpb_out[30][930],u_xpb_out[31][930],u_xpb_out[32][930],u_xpb_out[33][930],u_xpb_out[34][930],u_xpb_out[35][930],u_xpb_out[36][930],u_xpb_out[37][930],u_xpb_out[38][930],u_xpb_out[39][930],u_xpb_out[40][930],u_xpb_out[41][930],u_xpb_out[42][930],u_xpb_out[43][930],u_xpb_out[44][930],u_xpb_out[45][930],u_xpb_out[46][930],u_xpb_out[47][930],u_xpb_out[48][930],u_xpb_out[49][930],u_xpb_out[50][930],u_xpb_out[51][930],u_xpb_out[52][930],u_xpb_out[53][930],u_xpb_out[54][930],u_xpb_out[55][930],u_xpb_out[56][930],u_xpb_out[57][930],u_xpb_out[58][930],u_xpb_out[59][930],u_xpb_out[60][930],u_xpb_out[61][930],u_xpb_out[62][930],u_xpb_out[63][930],u_xpb_out[64][930],u_xpb_out[65][930],u_xpb_out[66][930],u_xpb_out[67][930],u_xpb_out[68][930],u_xpb_out[69][930],u_xpb_out[70][930],u_xpb_out[71][930],u_xpb_out[72][930],u_xpb_out[73][930],u_xpb_out[74][930],u_xpb_out[75][930],u_xpb_out[76][930],u_xpb_out[77][930],u_xpb_out[78][930],u_xpb_out[79][930],u_xpb_out[80][930],u_xpb_out[81][930],u_xpb_out[82][930],u_xpb_out[83][930],u_xpb_out[84][930],u_xpb_out[85][930],u_xpb_out[86][930],u_xpb_out[87][930],u_xpb_out[88][930],u_xpb_out[89][930],u_xpb_out[90][930],u_xpb_out[91][930],u_xpb_out[92][930],u_xpb_out[93][930],u_xpb_out[94][930],u_xpb_out[95][930],u_xpb_out[96][930],u_xpb_out[97][930],u_xpb_out[98][930],u_xpb_out[99][930],u_xpb_out[100][930],u_xpb_out[101][930],u_xpb_out[102][930],u_xpb_out[103][930],u_xpb_out[104][930],u_xpb_out[105][930]};

assign col_out_931 = {u_xpb_out[0][931],u_xpb_out[1][931],u_xpb_out[2][931],u_xpb_out[3][931],u_xpb_out[4][931],u_xpb_out[5][931],u_xpb_out[6][931],u_xpb_out[7][931],u_xpb_out[8][931],u_xpb_out[9][931],u_xpb_out[10][931],u_xpb_out[11][931],u_xpb_out[12][931],u_xpb_out[13][931],u_xpb_out[14][931],u_xpb_out[15][931],u_xpb_out[16][931],u_xpb_out[17][931],u_xpb_out[18][931],u_xpb_out[19][931],u_xpb_out[20][931],u_xpb_out[21][931],u_xpb_out[22][931],u_xpb_out[23][931],u_xpb_out[24][931],u_xpb_out[25][931],u_xpb_out[26][931],u_xpb_out[27][931],u_xpb_out[28][931],u_xpb_out[29][931],u_xpb_out[30][931],u_xpb_out[31][931],u_xpb_out[32][931],u_xpb_out[33][931],u_xpb_out[34][931],u_xpb_out[35][931],u_xpb_out[36][931],u_xpb_out[37][931],u_xpb_out[38][931],u_xpb_out[39][931],u_xpb_out[40][931],u_xpb_out[41][931],u_xpb_out[42][931],u_xpb_out[43][931],u_xpb_out[44][931],u_xpb_out[45][931],u_xpb_out[46][931],u_xpb_out[47][931],u_xpb_out[48][931],u_xpb_out[49][931],u_xpb_out[50][931],u_xpb_out[51][931],u_xpb_out[52][931],u_xpb_out[53][931],u_xpb_out[54][931],u_xpb_out[55][931],u_xpb_out[56][931],u_xpb_out[57][931],u_xpb_out[58][931],u_xpb_out[59][931],u_xpb_out[60][931],u_xpb_out[61][931],u_xpb_out[62][931],u_xpb_out[63][931],u_xpb_out[64][931],u_xpb_out[65][931],u_xpb_out[66][931],u_xpb_out[67][931],u_xpb_out[68][931],u_xpb_out[69][931],u_xpb_out[70][931],u_xpb_out[71][931],u_xpb_out[72][931],u_xpb_out[73][931],u_xpb_out[74][931],u_xpb_out[75][931],u_xpb_out[76][931],u_xpb_out[77][931],u_xpb_out[78][931],u_xpb_out[79][931],u_xpb_out[80][931],u_xpb_out[81][931],u_xpb_out[82][931],u_xpb_out[83][931],u_xpb_out[84][931],u_xpb_out[85][931],u_xpb_out[86][931],u_xpb_out[87][931],u_xpb_out[88][931],u_xpb_out[89][931],u_xpb_out[90][931],u_xpb_out[91][931],u_xpb_out[92][931],u_xpb_out[93][931],u_xpb_out[94][931],u_xpb_out[95][931],u_xpb_out[96][931],u_xpb_out[97][931],u_xpb_out[98][931],u_xpb_out[99][931],u_xpb_out[100][931],u_xpb_out[101][931],u_xpb_out[102][931],u_xpb_out[103][931],u_xpb_out[104][931],u_xpb_out[105][931]};

assign col_out_932 = {u_xpb_out[0][932],u_xpb_out[1][932],u_xpb_out[2][932],u_xpb_out[3][932],u_xpb_out[4][932],u_xpb_out[5][932],u_xpb_out[6][932],u_xpb_out[7][932],u_xpb_out[8][932],u_xpb_out[9][932],u_xpb_out[10][932],u_xpb_out[11][932],u_xpb_out[12][932],u_xpb_out[13][932],u_xpb_out[14][932],u_xpb_out[15][932],u_xpb_out[16][932],u_xpb_out[17][932],u_xpb_out[18][932],u_xpb_out[19][932],u_xpb_out[20][932],u_xpb_out[21][932],u_xpb_out[22][932],u_xpb_out[23][932],u_xpb_out[24][932],u_xpb_out[25][932],u_xpb_out[26][932],u_xpb_out[27][932],u_xpb_out[28][932],u_xpb_out[29][932],u_xpb_out[30][932],u_xpb_out[31][932],u_xpb_out[32][932],u_xpb_out[33][932],u_xpb_out[34][932],u_xpb_out[35][932],u_xpb_out[36][932],u_xpb_out[37][932],u_xpb_out[38][932],u_xpb_out[39][932],u_xpb_out[40][932],u_xpb_out[41][932],u_xpb_out[42][932],u_xpb_out[43][932],u_xpb_out[44][932],u_xpb_out[45][932],u_xpb_out[46][932],u_xpb_out[47][932],u_xpb_out[48][932],u_xpb_out[49][932],u_xpb_out[50][932],u_xpb_out[51][932],u_xpb_out[52][932],u_xpb_out[53][932],u_xpb_out[54][932],u_xpb_out[55][932],u_xpb_out[56][932],u_xpb_out[57][932],u_xpb_out[58][932],u_xpb_out[59][932],u_xpb_out[60][932],u_xpb_out[61][932],u_xpb_out[62][932],u_xpb_out[63][932],u_xpb_out[64][932],u_xpb_out[65][932],u_xpb_out[66][932],u_xpb_out[67][932],u_xpb_out[68][932],u_xpb_out[69][932],u_xpb_out[70][932],u_xpb_out[71][932],u_xpb_out[72][932],u_xpb_out[73][932],u_xpb_out[74][932],u_xpb_out[75][932],u_xpb_out[76][932],u_xpb_out[77][932],u_xpb_out[78][932],u_xpb_out[79][932],u_xpb_out[80][932],u_xpb_out[81][932],u_xpb_out[82][932],u_xpb_out[83][932],u_xpb_out[84][932],u_xpb_out[85][932],u_xpb_out[86][932],u_xpb_out[87][932],u_xpb_out[88][932],u_xpb_out[89][932],u_xpb_out[90][932],u_xpb_out[91][932],u_xpb_out[92][932],u_xpb_out[93][932],u_xpb_out[94][932],u_xpb_out[95][932],u_xpb_out[96][932],u_xpb_out[97][932],u_xpb_out[98][932],u_xpb_out[99][932],u_xpb_out[100][932],u_xpb_out[101][932],u_xpb_out[102][932],u_xpb_out[103][932],u_xpb_out[104][932],u_xpb_out[105][932]};

assign col_out_933 = {u_xpb_out[0][933],u_xpb_out[1][933],u_xpb_out[2][933],u_xpb_out[3][933],u_xpb_out[4][933],u_xpb_out[5][933],u_xpb_out[6][933],u_xpb_out[7][933],u_xpb_out[8][933],u_xpb_out[9][933],u_xpb_out[10][933],u_xpb_out[11][933],u_xpb_out[12][933],u_xpb_out[13][933],u_xpb_out[14][933],u_xpb_out[15][933],u_xpb_out[16][933],u_xpb_out[17][933],u_xpb_out[18][933],u_xpb_out[19][933],u_xpb_out[20][933],u_xpb_out[21][933],u_xpb_out[22][933],u_xpb_out[23][933],u_xpb_out[24][933],u_xpb_out[25][933],u_xpb_out[26][933],u_xpb_out[27][933],u_xpb_out[28][933],u_xpb_out[29][933],u_xpb_out[30][933],u_xpb_out[31][933],u_xpb_out[32][933],u_xpb_out[33][933],u_xpb_out[34][933],u_xpb_out[35][933],u_xpb_out[36][933],u_xpb_out[37][933],u_xpb_out[38][933],u_xpb_out[39][933],u_xpb_out[40][933],u_xpb_out[41][933],u_xpb_out[42][933],u_xpb_out[43][933],u_xpb_out[44][933],u_xpb_out[45][933],u_xpb_out[46][933],u_xpb_out[47][933],u_xpb_out[48][933],u_xpb_out[49][933],u_xpb_out[50][933],u_xpb_out[51][933],u_xpb_out[52][933],u_xpb_out[53][933],u_xpb_out[54][933],u_xpb_out[55][933],u_xpb_out[56][933],u_xpb_out[57][933],u_xpb_out[58][933],u_xpb_out[59][933],u_xpb_out[60][933],u_xpb_out[61][933],u_xpb_out[62][933],u_xpb_out[63][933],u_xpb_out[64][933],u_xpb_out[65][933],u_xpb_out[66][933],u_xpb_out[67][933],u_xpb_out[68][933],u_xpb_out[69][933],u_xpb_out[70][933],u_xpb_out[71][933],u_xpb_out[72][933],u_xpb_out[73][933],u_xpb_out[74][933],u_xpb_out[75][933],u_xpb_out[76][933],u_xpb_out[77][933],u_xpb_out[78][933],u_xpb_out[79][933],u_xpb_out[80][933],u_xpb_out[81][933],u_xpb_out[82][933],u_xpb_out[83][933],u_xpb_out[84][933],u_xpb_out[85][933],u_xpb_out[86][933],u_xpb_out[87][933],u_xpb_out[88][933],u_xpb_out[89][933],u_xpb_out[90][933],u_xpb_out[91][933],u_xpb_out[92][933],u_xpb_out[93][933],u_xpb_out[94][933],u_xpb_out[95][933],u_xpb_out[96][933],u_xpb_out[97][933],u_xpb_out[98][933],u_xpb_out[99][933],u_xpb_out[100][933],u_xpb_out[101][933],u_xpb_out[102][933],u_xpb_out[103][933],u_xpb_out[104][933],u_xpb_out[105][933]};

assign col_out_934 = {u_xpb_out[0][934],u_xpb_out[1][934],u_xpb_out[2][934],u_xpb_out[3][934],u_xpb_out[4][934],u_xpb_out[5][934],u_xpb_out[6][934],u_xpb_out[7][934],u_xpb_out[8][934],u_xpb_out[9][934],u_xpb_out[10][934],u_xpb_out[11][934],u_xpb_out[12][934],u_xpb_out[13][934],u_xpb_out[14][934],u_xpb_out[15][934],u_xpb_out[16][934],u_xpb_out[17][934],u_xpb_out[18][934],u_xpb_out[19][934],u_xpb_out[20][934],u_xpb_out[21][934],u_xpb_out[22][934],u_xpb_out[23][934],u_xpb_out[24][934],u_xpb_out[25][934],u_xpb_out[26][934],u_xpb_out[27][934],u_xpb_out[28][934],u_xpb_out[29][934],u_xpb_out[30][934],u_xpb_out[31][934],u_xpb_out[32][934],u_xpb_out[33][934],u_xpb_out[34][934],u_xpb_out[35][934],u_xpb_out[36][934],u_xpb_out[37][934],u_xpb_out[38][934],u_xpb_out[39][934],u_xpb_out[40][934],u_xpb_out[41][934],u_xpb_out[42][934],u_xpb_out[43][934],u_xpb_out[44][934],u_xpb_out[45][934],u_xpb_out[46][934],u_xpb_out[47][934],u_xpb_out[48][934],u_xpb_out[49][934],u_xpb_out[50][934],u_xpb_out[51][934],u_xpb_out[52][934],u_xpb_out[53][934],u_xpb_out[54][934],u_xpb_out[55][934],u_xpb_out[56][934],u_xpb_out[57][934],u_xpb_out[58][934],u_xpb_out[59][934],u_xpb_out[60][934],u_xpb_out[61][934],u_xpb_out[62][934],u_xpb_out[63][934],u_xpb_out[64][934],u_xpb_out[65][934],u_xpb_out[66][934],u_xpb_out[67][934],u_xpb_out[68][934],u_xpb_out[69][934],u_xpb_out[70][934],u_xpb_out[71][934],u_xpb_out[72][934],u_xpb_out[73][934],u_xpb_out[74][934],u_xpb_out[75][934],u_xpb_out[76][934],u_xpb_out[77][934],u_xpb_out[78][934],u_xpb_out[79][934],u_xpb_out[80][934],u_xpb_out[81][934],u_xpb_out[82][934],u_xpb_out[83][934],u_xpb_out[84][934],u_xpb_out[85][934],u_xpb_out[86][934],u_xpb_out[87][934],u_xpb_out[88][934],u_xpb_out[89][934],u_xpb_out[90][934],u_xpb_out[91][934],u_xpb_out[92][934],u_xpb_out[93][934],u_xpb_out[94][934],u_xpb_out[95][934],u_xpb_out[96][934],u_xpb_out[97][934],u_xpb_out[98][934],u_xpb_out[99][934],u_xpb_out[100][934],u_xpb_out[101][934],u_xpb_out[102][934],u_xpb_out[103][934],u_xpb_out[104][934],u_xpb_out[105][934]};

assign col_out_935 = {u_xpb_out[0][935],u_xpb_out[1][935],u_xpb_out[2][935],u_xpb_out[3][935],u_xpb_out[4][935],u_xpb_out[5][935],u_xpb_out[6][935],u_xpb_out[7][935],u_xpb_out[8][935],u_xpb_out[9][935],u_xpb_out[10][935],u_xpb_out[11][935],u_xpb_out[12][935],u_xpb_out[13][935],u_xpb_out[14][935],u_xpb_out[15][935],u_xpb_out[16][935],u_xpb_out[17][935],u_xpb_out[18][935],u_xpb_out[19][935],u_xpb_out[20][935],u_xpb_out[21][935],u_xpb_out[22][935],u_xpb_out[23][935],u_xpb_out[24][935],u_xpb_out[25][935],u_xpb_out[26][935],u_xpb_out[27][935],u_xpb_out[28][935],u_xpb_out[29][935],u_xpb_out[30][935],u_xpb_out[31][935],u_xpb_out[32][935],u_xpb_out[33][935],u_xpb_out[34][935],u_xpb_out[35][935],u_xpb_out[36][935],u_xpb_out[37][935],u_xpb_out[38][935],u_xpb_out[39][935],u_xpb_out[40][935],u_xpb_out[41][935],u_xpb_out[42][935],u_xpb_out[43][935],u_xpb_out[44][935],u_xpb_out[45][935],u_xpb_out[46][935],u_xpb_out[47][935],u_xpb_out[48][935],u_xpb_out[49][935],u_xpb_out[50][935],u_xpb_out[51][935],u_xpb_out[52][935],u_xpb_out[53][935],u_xpb_out[54][935],u_xpb_out[55][935],u_xpb_out[56][935],u_xpb_out[57][935],u_xpb_out[58][935],u_xpb_out[59][935],u_xpb_out[60][935],u_xpb_out[61][935],u_xpb_out[62][935],u_xpb_out[63][935],u_xpb_out[64][935],u_xpb_out[65][935],u_xpb_out[66][935],u_xpb_out[67][935],u_xpb_out[68][935],u_xpb_out[69][935],u_xpb_out[70][935],u_xpb_out[71][935],u_xpb_out[72][935],u_xpb_out[73][935],u_xpb_out[74][935],u_xpb_out[75][935],u_xpb_out[76][935],u_xpb_out[77][935],u_xpb_out[78][935],u_xpb_out[79][935],u_xpb_out[80][935],u_xpb_out[81][935],u_xpb_out[82][935],u_xpb_out[83][935],u_xpb_out[84][935],u_xpb_out[85][935],u_xpb_out[86][935],u_xpb_out[87][935],u_xpb_out[88][935],u_xpb_out[89][935],u_xpb_out[90][935],u_xpb_out[91][935],u_xpb_out[92][935],u_xpb_out[93][935],u_xpb_out[94][935],u_xpb_out[95][935],u_xpb_out[96][935],u_xpb_out[97][935],u_xpb_out[98][935],u_xpb_out[99][935],u_xpb_out[100][935],u_xpb_out[101][935],u_xpb_out[102][935],u_xpb_out[103][935],u_xpb_out[104][935],u_xpb_out[105][935]};

assign col_out_936 = {u_xpb_out[0][936],u_xpb_out[1][936],u_xpb_out[2][936],u_xpb_out[3][936],u_xpb_out[4][936],u_xpb_out[5][936],u_xpb_out[6][936],u_xpb_out[7][936],u_xpb_out[8][936],u_xpb_out[9][936],u_xpb_out[10][936],u_xpb_out[11][936],u_xpb_out[12][936],u_xpb_out[13][936],u_xpb_out[14][936],u_xpb_out[15][936],u_xpb_out[16][936],u_xpb_out[17][936],u_xpb_out[18][936],u_xpb_out[19][936],u_xpb_out[20][936],u_xpb_out[21][936],u_xpb_out[22][936],u_xpb_out[23][936],u_xpb_out[24][936],u_xpb_out[25][936],u_xpb_out[26][936],u_xpb_out[27][936],u_xpb_out[28][936],u_xpb_out[29][936],u_xpb_out[30][936],u_xpb_out[31][936],u_xpb_out[32][936],u_xpb_out[33][936],u_xpb_out[34][936],u_xpb_out[35][936],u_xpb_out[36][936],u_xpb_out[37][936],u_xpb_out[38][936],u_xpb_out[39][936],u_xpb_out[40][936],u_xpb_out[41][936],u_xpb_out[42][936],u_xpb_out[43][936],u_xpb_out[44][936],u_xpb_out[45][936],u_xpb_out[46][936],u_xpb_out[47][936],u_xpb_out[48][936],u_xpb_out[49][936],u_xpb_out[50][936],u_xpb_out[51][936],u_xpb_out[52][936],u_xpb_out[53][936],u_xpb_out[54][936],u_xpb_out[55][936],u_xpb_out[56][936],u_xpb_out[57][936],u_xpb_out[58][936],u_xpb_out[59][936],u_xpb_out[60][936],u_xpb_out[61][936],u_xpb_out[62][936],u_xpb_out[63][936],u_xpb_out[64][936],u_xpb_out[65][936],u_xpb_out[66][936],u_xpb_out[67][936],u_xpb_out[68][936],u_xpb_out[69][936],u_xpb_out[70][936],u_xpb_out[71][936],u_xpb_out[72][936],u_xpb_out[73][936],u_xpb_out[74][936],u_xpb_out[75][936],u_xpb_out[76][936],u_xpb_out[77][936],u_xpb_out[78][936],u_xpb_out[79][936],u_xpb_out[80][936],u_xpb_out[81][936],u_xpb_out[82][936],u_xpb_out[83][936],u_xpb_out[84][936],u_xpb_out[85][936],u_xpb_out[86][936],u_xpb_out[87][936],u_xpb_out[88][936],u_xpb_out[89][936],u_xpb_out[90][936],u_xpb_out[91][936],u_xpb_out[92][936],u_xpb_out[93][936],u_xpb_out[94][936],u_xpb_out[95][936],u_xpb_out[96][936],u_xpb_out[97][936],u_xpb_out[98][936],u_xpb_out[99][936],u_xpb_out[100][936],u_xpb_out[101][936],u_xpb_out[102][936],u_xpb_out[103][936],u_xpb_out[104][936],u_xpb_out[105][936]};

assign col_out_937 = {u_xpb_out[0][937],u_xpb_out[1][937],u_xpb_out[2][937],u_xpb_out[3][937],u_xpb_out[4][937],u_xpb_out[5][937],u_xpb_out[6][937],u_xpb_out[7][937],u_xpb_out[8][937],u_xpb_out[9][937],u_xpb_out[10][937],u_xpb_out[11][937],u_xpb_out[12][937],u_xpb_out[13][937],u_xpb_out[14][937],u_xpb_out[15][937],u_xpb_out[16][937],u_xpb_out[17][937],u_xpb_out[18][937],u_xpb_out[19][937],u_xpb_out[20][937],u_xpb_out[21][937],u_xpb_out[22][937],u_xpb_out[23][937],u_xpb_out[24][937],u_xpb_out[25][937],u_xpb_out[26][937],u_xpb_out[27][937],u_xpb_out[28][937],u_xpb_out[29][937],u_xpb_out[30][937],u_xpb_out[31][937],u_xpb_out[32][937],u_xpb_out[33][937],u_xpb_out[34][937],u_xpb_out[35][937],u_xpb_out[36][937],u_xpb_out[37][937],u_xpb_out[38][937],u_xpb_out[39][937],u_xpb_out[40][937],u_xpb_out[41][937],u_xpb_out[42][937],u_xpb_out[43][937],u_xpb_out[44][937],u_xpb_out[45][937],u_xpb_out[46][937],u_xpb_out[47][937],u_xpb_out[48][937],u_xpb_out[49][937],u_xpb_out[50][937],u_xpb_out[51][937],u_xpb_out[52][937],u_xpb_out[53][937],u_xpb_out[54][937],u_xpb_out[55][937],u_xpb_out[56][937],u_xpb_out[57][937],u_xpb_out[58][937],u_xpb_out[59][937],u_xpb_out[60][937],u_xpb_out[61][937],u_xpb_out[62][937],u_xpb_out[63][937],u_xpb_out[64][937],u_xpb_out[65][937],u_xpb_out[66][937],u_xpb_out[67][937],u_xpb_out[68][937],u_xpb_out[69][937],u_xpb_out[70][937],u_xpb_out[71][937],u_xpb_out[72][937],u_xpb_out[73][937],u_xpb_out[74][937],u_xpb_out[75][937],u_xpb_out[76][937],u_xpb_out[77][937],u_xpb_out[78][937],u_xpb_out[79][937],u_xpb_out[80][937],u_xpb_out[81][937],u_xpb_out[82][937],u_xpb_out[83][937],u_xpb_out[84][937],u_xpb_out[85][937],u_xpb_out[86][937],u_xpb_out[87][937],u_xpb_out[88][937],u_xpb_out[89][937],u_xpb_out[90][937],u_xpb_out[91][937],u_xpb_out[92][937],u_xpb_out[93][937],u_xpb_out[94][937],u_xpb_out[95][937],u_xpb_out[96][937],u_xpb_out[97][937],u_xpb_out[98][937],u_xpb_out[99][937],u_xpb_out[100][937],u_xpb_out[101][937],u_xpb_out[102][937],u_xpb_out[103][937],u_xpb_out[104][937],u_xpb_out[105][937]};

assign col_out_938 = {u_xpb_out[0][938],u_xpb_out[1][938],u_xpb_out[2][938],u_xpb_out[3][938],u_xpb_out[4][938],u_xpb_out[5][938],u_xpb_out[6][938],u_xpb_out[7][938],u_xpb_out[8][938],u_xpb_out[9][938],u_xpb_out[10][938],u_xpb_out[11][938],u_xpb_out[12][938],u_xpb_out[13][938],u_xpb_out[14][938],u_xpb_out[15][938],u_xpb_out[16][938],u_xpb_out[17][938],u_xpb_out[18][938],u_xpb_out[19][938],u_xpb_out[20][938],u_xpb_out[21][938],u_xpb_out[22][938],u_xpb_out[23][938],u_xpb_out[24][938],u_xpb_out[25][938],u_xpb_out[26][938],u_xpb_out[27][938],u_xpb_out[28][938],u_xpb_out[29][938],u_xpb_out[30][938],u_xpb_out[31][938],u_xpb_out[32][938],u_xpb_out[33][938],u_xpb_out[34][938],u_xpb_out[35][938],u_xpb_out[36][938],u_xpb_out[37][938],u_xpb_out[38][938],u_xpb_out[39][938],u_xpb_out[40][938],u_xpb_out[41][938],u_xpb_out[42][938],u_xpb_out[43][938],u_xpb_out[44][938],u_xpb_out[45][938],u_xpb_out[46][938],u_xpb_out[47][938],u_xpb_out[48][938],u_xpb_out[49][938],u_xpb_out[50][938],u_xpb_out[51][938],u_xpb_out[52][938],u_xpb_out[53][938],u_xpb_out[54][938],u_xpb_out[55][938],u_xpb_out[56][938],u_xpb_out[57][938],u_xpb_out[58][938],u_xpb_out[59][938],u_xpb_out[60][938],u_xpb_out[61][938],u_xpb_out[62][938],u_xpb_out[63][938],u_xpb_out[64][938],u_xpb_out[65][938],u_xpb_out[66][938],u_xpb_out[67][938],u_xpb_out[68][938],u_xpb_out[69][938],u_xpb_out[70][938],u_xpb_out[71][938],u_xpb_out[72][938],u_xpb_out[73][938],u_xpb_out[74][938],u_xpb_out[75][938],u_xpb_out[76][938],u_xpb_out[77][938],u_xpb_out[78][938],u_xpb_out[79][938],u_xpb_out[80][938],u_xpb_out[81][938],u_xpb_out[82][938],u_xpb_out[83][938],u_xpb_out[84][938],u_xpb_out[85][938],u_xpb_out[86][938],u_xpb_out[87][938],u_xpb_out[88][938],u_xpb_out[89][938],u_xpb_out[90][938],u_xpb_out[91][938],u_xpb_out[92][938],u_xpb_out[93][938],u_xpb_out[94][938],u_xpb_out[95][938],u_xpb_out[96][938],u_xpb_out[97][938],u_xpb_out[98][938],u_xpb_out[99][938],u_xpb_out[100][938],u_xpb_out[101][938],u_xpb_out[102][938],u_xpb_out[103][938],u_xpb_out[104][938],u_xpb_out[105][938]};

assign col_out_939 = {u_xpb_out[0][939],u_xpb_out[1][939],u_xpb_out[2][939],u_xpb_out[3][939],u_xpb_out[4][939],u_xpb_out[5][939],u_xpb_out[6][939],u_xpb_out[7][939],u_xpb_out[8][939],u_xpb_out[9][939],u_xpb_out[10][939],u_xpb_out[11][939],u_xpb_out[12][939],u_xpb_out[13][939],u_xpb_out[14][939],u_xpb_out[15][939],u_xpb_out[16][939],u_xpb_out[17][939],u_xpb_out[18][939],u_xpb_out[19][939],u_xpb_out[20][939],u_xpb_out[21][939],u_xpb_out[22][939],u_xpb_out[23][939],u_xpb_out[24][939],u_xpb_out[25][939],u_xpb_out[26][939],u_xpb_out[27][939],u_xpb_out[28][939],u_xpb_out[29][939],u_xpb_out[30][939],u_xpb_out[31][939],u_xpb_out[32][939],u_xpb_out[33][939],u_xpb_out[34][939],u_xpb_out[35][939],u_xpb_out[36][939],u_xpb_out[37][939],u_xpb_out[38][939],u_xpb_out[39][939],u_xpb_out[40][939],u_xpb_out[41][939],u_xpb_out[42][939],u_xpb_out[43][939],u_xpb_out[44][939],u_xpb_out[45][939],u_xpb_out[46][939],u_xpb_out[47][939],u_xpb_out[48][939],u_xpb_out[49][939],u_xpb_out[50][939],u_xpb_out[51][939],u_xpb_out[52][939],u_xpb_out[53][939],u_xpb_out[54][939],u_xpb_out[55][939],u_xpb_out[56][939],u_xpb_out[57][939],u_xpb_out[58][939],u_xpb_out[59][939],u_xpb_out[60][939],u_xpb_out[61][939],u_xpb_out[62][939],u_xpb_out[63][939],u_xpb_out[64][939],u_xpb_out[65][939],u_xpb_out[66][939],u_xpb_out[67][939],u_xpb_out[68][939],u_xpb_out[69][939],u_xpb_out[70][939],u_xpb_out[71][939],u_xpb_out[72][939],u_xpb_out[73][939],u_xpb_out[74][939],u_xpb_out[75][939],u_xpb_out[76][939],u_xpb_out[77][939],u_xpb_out[78][939],u_xpb_out[79][939],u_xpb_out[80][939],u_xpb_out[81][939],u_xpb_out[82][939],u_xpb_out[83][939],u_xpb_out[84][939],u_xpb_out[85][939],u_xpb_out[86][939],u_xpb_out[87][939],u_xpb_out[88][939],u_xpb_out[89][939],u_xpb_out[90][939],u_xpb_out[91][939],u_xpb_out[92][939],u_xpb_out[93][939],u_xpb_out[94][939],u_xpb_out[95][939],u_xpb_out[96][939],u_xpb_out[97][939],u_xpb_out[98][939],u_xpb_out[99][939],u_xpb_out[100][939],u_xpb_out[101][939],u_xpb_out[102][939],u_xpb_out[103][939],u_xpb_out[104][939],u_xpb_out[105][939]};

assign col_out_940 = {u_xpb_out[0][940],u_xpb_out[1][940],u_xpb_out[2][940],u_xpb_out[3][940],u_xpb_out[4][940],u_xpb_out[5][940],u_xpb_out[6][940],u_xpb_out[7][940],u_xpb_out[8][940],u_xpb_out[9][940],u_xpb_out[10][940],u_xpb_out[11][940],u_xpb_out[12][940],u_xpb_out[13][940],u_xpb_out[14][940],u_xpb_out[15][940],u_xpb_out[16][940],u_xpb_out[17][940],u_xpb_out[18][940],u_xpb_out[19][940],u_xpb_out[20][940],u_xpb_out[21][940],u_xpb_out[22][940],u_xpb_out[23][940],u_xpb_out[24][940],u_xpb_out[25][940],u_xpb_out[26][940],u_xpb_out[27][940],u_xpb_out[28][940],u_xpb_out[29][940],u_xpb_out[30][940],u_xpb_out[31][940],u_xpb_out[32][940],u_xpb_out[33][940],u_xpb_out[34][940],u_xpb_out[35][940],u_xpb_out[36][940],u_xpb_out[37][940],u_xpb_out[38][940],u_xpb_out[39][940],u_xpb_out[40][940],u_xpb_out[41][940],u_xpb_out[42][940],u_xpb_out[43][940],u_xpb_out[44][940],u_xpb_out[45][940],u_xpb_out[46][940],u_xpb_out[47][940],u_xpb_out[48][940],u_xpb_out[49][940],u_xpb_out[50][940],u_xpb_out[51][940],u_xpb_out[52][940],u_xpb_out[53][940],u_xpb_out[54][940],u_xpb_out[55][940],u_xpb_out[56][940],u_xpb_out[57][940],u_xpb_out[58][940],u_xpb_out[59][940],u_xpb_out[60][940],u_xpb_out[61][940],u_xpb_out[62][940],u_xpb_out[63][940],u_xpb_out[64][940],u_xpb_out[65][940],u_xpb_out[66][940],u_xpb_out[67][940],u_xpb_out[68][940],u_xpb_out[69][940],u_xpb_out[70][940],u_xpb_out[71][940],u_xpb_out[72][940],u_xpb_out[73][940],u_xpb_out[74][940],u_xpb_out[75][940],u_xpb_out[76][940],u_xpb_out[77][940],u_xpb_out[78][940],u_xpb_out[79][940],u_xpb_out[80][940],u_xpb_out[81][940],u_xpb_out[82][940],u_xpb_out[83][940],u_xpb_out[84][940],u_xpb_out[85][940],u_xpb_out[86][940],u_xpb_out[87][940],u_xpb_out[88][940],u_xpb_out[89][940],u_xpb_out[90][940],u_xpb_out[91][940],u_xpb_out[92][940],u_xpb_out[93][940],u_xpb_out[94][940],u_xpb_out[95][940],u_xpb_out[96][940],u_xpb_out[97][940],u_xpb_out[98][940],u_xpb_out[99][940],u_xpb_out[100][940],u_xpb_out[101][940],u_xpb_out[102][940],u_xpb_out[103][940],u_xpb_out[104][940],u_xpb_out[105][940]};

assign col_out_941 = {u_xpb_out[0][941],u_xpb_out[1][941],u_xpb_out[2][941],u_xpb_out[3][941],u_xpb_out[4][941],u_xpb_out[5][941],u_xpb_out[6][941],u_xpb_out[7][941],u_xpb_out[8][941],u_xpb_out[9][941],u_xpb_out[10][941],u_xpb_out[11][941],u_xpb_out[12][941],u_xpb_out[13][941],u_xpb_out[14][941],u_xpb_out[15][941],u_xpb_out[16][941],u_xpb_out[17][941],u_xpb_out[18][941],u_xpb_out[19][941],u_xpb_out[20][941],u_xpb_out[21][941],u_xpb_out[22][941],u_xpb_out[23][941],u_xpb_out[24][941],u_xpb_out[25][941],u_xpb_out[26][941],u_xpb_out[27][941],u_xpb_out[28][941],u_xpb_out[29][941],u_xpb_out[30][941],u_xpb_out[31][941],u_xpb_out[32][941],u_xpb_out[33][941],u_xpb_out[34][941],u_xpb_out[35][941],u_xpb_out[36][941],u_xpb_out[37][941],u_xpb_out[38][941],u_xpb_out[39][941],u_xpb_out[40][941],u_xpb_out[41][941],u_xpb_out[42][941],u_xpb_out[43][941],u_xpb_out[44][941],u_xpb_out[45][941],u_xpb_out[46][941],u_xpb_out[47][941],u_xpb_out[48][941],u_xpb_out[49][941],u_xpb_out[50][941],u_xpb_out[51][941],u_xpb_out[52][941],u_xpb_out[53][941],u_xpb_out[54][941],u_xpb_out[55][941],u_xpb_out[56][941],u_xpb_out[57][941],u_xpb_out[58][941],u_xpb_out[59][941],u_xpb_out[60][941],u_xpb_out[61][941],u_xpb_out[62][941],u_xpb_out[63][941],u_xpb_out[64][941],u_xpb_out[65][941],u_xpb_out[66][941],u_xpb_out[67][941],u_xpb_out[68][941],u_xpb_out[69][941],u_xpb_out[70][941],u_xpb_out[71][941],u_xpb_out[72][941],u_xpb_out[73][941],u_xpb_out[74][941],u_xpb_out[75][941],u_xpb_out[76][941],u_xpb_out[77][941],u_xpb_out[78][941],u_xpb_out[79][941],u_xpb_out[80][941],u_xpb_out[81][941],u_xpb_out[82][941],u_xpb_out[83][941],u_xpb_out[84][941],u_xpb_out[85][941],u_xpb_out[86][941],u_xpb_out[87][941],u_xpb_out[88][941],u_xpb_out[89][941],u_xpb_out[90][941],u_xpb_out[91][941],u_xpb_out[92][941],u_xpb_out[93][941],u_xpb_out[94][941],u_xpb_out[95][941],u_xpb_out[96][941],u_xpb_out[97][941],u_xpb_out[98][941],u_xpb_out[99][941],u_xpb_out[100][941],u_xpb_out[101][941],u_xpb_out[102][941],u_xpb_out[103][941],u_xpb_out[104][941],u_xpb_out[105][941]};

assign col_out_942 = {u_xpb_out[0][942],u_xpb_out[1][942],u_xpb_out[2][942],u_xpb_out[3][942],u_xpb_out[4][942],u_xpb_out[5][942],u_xpb_out[6][942],u_xpb_out[7][942],u_xpb_out[8][942],u_xpb_out[9][942],u_xpb_out[10][942],u_xpb_out[11][942],u_xpb_out[12][942],u_xpb_out[13][942],u_xpb_out[14][942],u_xpb_out[15][942],u_xpb_out[16][942],u_xpb_out[17][942],u_xpb_out[18][942],u_xpb_out[19][942],u_xpb_out[20][942],u_xpb_out[21][942],u_xpb_out[22][942],u_xpb_out[23][942],u_xpb_out[24][942],u_xpb_out[25][942],u_xpb_out[26][942],u_xpb_out[27][942],u_xpb_out[28][942],u_xpb_out[29][942],u_xpb_out[30][942],u_xpb_out[31][942],u_xpb_out[32][942],u_xpb_out[33][942],u_xpb_out[34][942],u_xpb_out[35][942],u_xpb_out[36][942],u_xpb_out[37][942],u_xpb_out[38][942],u_xpb_out[39][942],u_xpb_out[40][942],u_xpb_out[41][942],u_xpb_out[42][942],u_xpb_out[43][942],u_xpb_out[44][942],u_xpb_out[45][942],u_xpb_out[46][942],u_xpb_out[47][942],u_xpb_out[48][942],u_xpb_out[49][942],u_xpb_out[50][942],u_xpb_out[51][942],u_xpb_out[52][942],u_xpb_out[53][942],u_xpb_out[54][942],u_xpb_out[55][942],u_xpb_out[56][942],u_xpb_out[57][942],u_xpb_out[58][942],u_xpb_out[59][942],u_xpb_out[60][942],u_xpb_out[61][942],u_xpb_out[62][942],u_xpb_out[63][942],u_xpb_out[64][942],u_xpb_out[65][942],u_xpb_out[66][942],u_xpb_out[67][942],u_xpb_out[68][942],u_xpb_out[69][942],u_xpb_out[70][942],u_xpb_out[71][942],u_xpb_out[72][942],u_xpb_out[73][942],u_xpb_out[74][942],u_xpb_out[75][942],u_xpb_out[76][942],u_xpb_out[77][942],u_xpb_out[78][942],u_xpb_out[79][942],u_xpb_out[80][942],u_xpb_out[81][942],u_xpb_out[82][942],u_xpb_out[83][942],u_xpb_out[84][942],u_xpb_out[85][942],u_xpb_out[86][942],u_xpb_out[87][942],u_xpb_out[88][942],u_xpb_out[89][942],u_xpb_out[90][942],u_xpb_out[91][942],u_xpb_out[92][942],u_xpb_out[93][942],u_xpb_out[94][942],u_xpb_out[95][942],u_xpb_out[96][942],u_xpb_out[97][942],u_xpb_out[98][942],u_xpb_out[99][942],u_xpb_out[100][942],u_xpb_out[101][942],u_xpb_out[102][942],u_xpb_out[103][942],u_xpb_out[104][942],u_xpb_out[105][942]};

assign col_out_943 = {u_xpb_out[0][943],u_xpb_out[1][943],u_xpb_out[2][943],u_xpb_out[3][943],u_xpb_out[4][943],u_xpb_out[5][943],u_xpb_out[6][943],u_xpb_out[7][943],u_xpb_out[8][943],u_xpb_out[9][943],u_xpb_out[10][943],u_xpb_out[11][943],u_xpb_out[12][943],u_xpb_out[13][943],u_xpb_out[14][943],u_xpb_out[15][943],u_xpb_out[16][943],u_xpb_out[17][943],u_xpb_out[18][943],u_xpb_out[19][943],u_xpb_out[20][943],u_xpb_out[21][943],u_xpb_out[22][943],u_xpb_out[23][943],u_xpb_out[24][943],u_xpb_out[25][943],u_xpb_out[26][943],u_xpb_out[27][943],u_xpb_out[28][943],u_xpb_out[29][943],u_xpb_out[30][943],u_xpb_out[31][943],u_xpb_out[32][943],u_xpb_out[33][943],u_xpb_out[34][943],u_xpb_out[35][943],u_xpb_out[36][943],u_xpb_out[37][943],u_xpb_out[38][943],u_xpb_out[39][943],u_xpb_out[40][943],u_xpb_out[41][943],u_xpb_out[42][943],u_xpb_out[43][943],u_xpb_out[44][943],u_xpb_out[45][943],u_xpb_out[46][943],u_xpb_out[47][943],u_xpb_out[48][943],u_xpb_out[49][943],u_xpb_out[50][943],u_xpb_out[51][943],u_xpb_out[52][943],u_xpb_out[53][943],u_xpb_out[54][943],u_xpb_out[55][943],u_xpb_out[56][943],u_xpb_out[57][943],u_xpb_out[58][943],u_xpb_out[59][943],u_xpb_out[60][943],u_xpb_out[61][943],u_xpb_out[62][943],u_xpb_out[63][943],u_xpb_out[64][943],u_xpb_out[65][943],u_xpb_out[66][943],u_xpb_out[67][943],u_xpb_out[68][943],u_xpb_out[69][943],u_xpb_out[70][943],u_xpb_out[71][943],u_xpb_out[72][943],u_xpb_out[73][943],u_xpb_out[74][943],u_xpb_out[75][943],u_xpb_out[76][943],u_xpb_out[77][943],u_xpb_out[78][943],u_xpb_out[79][943],u_xpb_out[80][943],u_xpb_out[81][943],u_xpb_out[82][943],u_xpb_out[83][943],u_xpb_out[84][943],u_xpb_out[85][943],u_xpb_out[86][943],u_xpb_out[87][943],u_xpb_out[88][943],u_xpb_out[89][943],u_xpb_out[90][943],u_xpb_out[91][943],u_xpb_out[92][943],u_xpb_out[93][943],u_xpb_out[94][943],u_xpb_out[95][943],u_xpb_out[96][943],u_xpb_out[97][943],u_xpb_out[98][943],u_xpb_out[99][943],u_xpb_out[100][943],u_xpb_out[101][943],u_xpb_out[102][943],u_xpb_out[103][943],u_xpb_out[104][943],u_xpb_out[105][943]};

assign col_out_944 = {u_xpb_out[0][944],u_xpb_out[1][944],u_xpb_out[2][944],u_xpb_out[3][944],u_xpb_out[4][944],u_xpb_out[5][944],u_xpb_out[6][944],u_xpb_out[7][944],u_xpb_out[8][944],u_xpb_out[9][944],u_xpb_out[10][944],u_xpb_out[11][944],u_xpb_out[12][944],u_xpb_out[13][944],u_xpb_out[14][944],u_xpb_out[15][944],u_xpb_out[16][944],u_xpb_out[17][944],u_xpb_out[18][944],u_xpb_out[19][944],u_xpb_out[20][944],u_xpb_out[21][944],u_xpb_out[22][944],u_xpb_out[23][944],u_xpb_out[24][944],u_xpb_out[25][944],u_xpb_out[26][944],u_xpb_out[27][944],u_xpb_out[28][944],u_xpb_out[29][944],u_xpb_out[30][944],u_xpb_out[31][944],u_xpb_out[32][944],u_xpb_out[33][944],u_xpb_out[34][944],u_xpb_out[35][944],u_xpb_out[36][944],u_xpb_out[37][944],u_xpb_out[38][944],u_xpb_out[39][944],u_xpb_out[40][944],u_xpb_out[41][944],u_xpb_out[42][944],u_xpb_out[43][944],u_xpb_out[44][944],u_xpb_out[45][944],u_xpb_out[46][944],u_xpb_out[47][944],u_xpb_out[48][944],u_xpb_out[49][944],u_xpb_out[50][944],u_xpb_out[51][944],u_xpb_out[52][944],u_xpb_out[53][944],u_xpb_out[54][944],u_xpb_out[55][944],u_xpb_out[56][944],u_xpb_out[57][944],u_xpb_out[58][944],u_xpb_out[59][944],u_xpb_out[60][944],u_xpb_out[61][944],u_xpb_out[62][944],u_xpb_out[63][944],u_xpb_out[64][944],u_xpb_out[65][944],u_xpb_out[66][944],u_xpb_out[67][944],u_xpb_out[68][944],u_xpb_out[69][944],u_xpb_out[70][944],u_xpb_out[71][944],u_xpb_out[72][944],u_xpb_out[73][944],u_xpb_out[74][944],u_xpb_out[75][944],u_xpb_out[76][944],u_xpb_out[77][944],u_xpb_out[78][944],u_xpb_out[79][944],u_xpb_out[80][944],u_xpb_out[81][944],u_xpb_out[82][944],u_xpb_out[83][944],u_xpb_out[84][944],u_xpb_out[85][944],u_xpb_out[86][944],u_xpb_out[87][944],u_xpb_out[88][944],u_xpb_out[89][944],u_xpb_out[90][944],u_xpb_out[91][944],u_xpb_out[92][944],u_xpb_out[93][944],u_xpb_out[94][944],u_xpb_out[95][944],u_xpb_out[96][944],u_xpb_out[97][944],u_xpb_out[98][944],u_xpb_out[99][944],u_xpb_out[100][944],u_xpb_out[101][944],u_xpb_out[102][944],u_xpb_out[103][944],u_xpb_out[104][944],u_xpb_out[105][944]};

assign col_out_945 = {u_xpb_out[0][945],u_xpb_out[1][945],u_xpb_out[2][945],u_xpb_out[3][945],u_xpb_out[4][945],u_xpb_out[5][945],u_xpb_out[6][945],u_xpb_out[7][945],u_xpb_out[8][945],u_xpb_out[9][945],u_xpb_out[10][945],u_xpb_out[11][945],u_xpb_out[12][945],u_xpb_out[13][945],u_xpb_out[14][945],u_xpb_out[15][945],u_xpb_out[16][945],u_xpb_out[17][945],u_xpb_out[18][945],u_xpb_out[19][945],u_xpb_out[20][945],u_xpb_out[21][945],u_xpb_out[22][945],u_xpb_out[23][945],u_xpb_out[24][945],u_xpb_out[25][945],u_xpb_out[26][945],u_xpb_out[27][945],u_xpb_out[28][945],u_xpb_out[29][945],u_xpb_out[30][945],u_xpb_out[31][945],u_xpb_out[32][945],u_xpb_out[33][945],u_xpb_out[34][945],u_xpb_out[35][945],u_xpb_out[36][945],u_xpb_out[37][945],u_xpb_out[38][945],u_xpb_out[39][945],u_xpb_out[40][945],u_xpb_out[41][945],u_xpb_out[42][945],u_xpb_out[43][945],u_xpb_out[44][945],u_xpb_out[45][945],u_xpb_out[46][945],u_xpb_out[47][945],u_xpb_out[48][945],u_xpb_out[49][945],u_xpb_out[50][945],u_xpb_out[51][945],u_xpb_out[52][945],u_xpb_out[53][945],u_xpb_out[54][945],u_xpb_out[55][945],u_xpb_out[56][945],u_xpb_out[57][945],u_xpb_out[58][945],u_xpb_out[59][945],u_xpb_out[60][945],u_xpb_out[61][945],u_xpb_out[62][945],u_xpb_out[63][945],u_xpb_out[64][945],u_xpb_out[65][945],u_xpb_out[66][945],u_xpb_out[67][945],u_xpb_out[68][945],u_xpb_out[69][945],u_xpb_out[70][945],u_xpb_out[71][945],u_xpb_out[72][945],u_xpb_out[73][945],u_xpb_out[74][945],u_xpb_out[75][945],u_xpb_out[76][945],u_xpb_out[77][945],u_xpb_out[78][945],u_xpb_out[79][945],u_xpb_out[80][945],u_xpb_out[81][945],u_xpb_out[82][945],u_xpb_out[83][945],u_xpb_out[84][945],u_xpb_out[85][945],u_xpb_out[86][945],u_xpb_out[87][945],u_xpb_out[88][945],u_xpb_out[89][945],u_xpb_out[90][945],u_xpb_out[91][945],u_xpb_out[92][945],u_xpb_out[93][945],u_xpb_out[94][945],u_xpb_out[95][945],u_xpb_out[96][945],u_xpb_out[97][945],u_xpb_out[98][945],u_xpb_out[99][945],u_xpb_out[100][945],u_xpb_out[101][945],u_xpb_out[102][945],u_xpb_out[103][945],u_xpb_out[104][945],u_xpb_out[105][945]};

assign col_out_946 = {u_xpb_out[0][946],u_xpb_out[1][946],u_xpb_out[2][946],u_xpb_out[3][946],u_xpb_out[4][946],u_xpb_out[5][946],u_xpb_out[6][946],u_xpb_out[7][946],u_xpb_out[8][946],u_xpb_out[9][946],u_xpb_out[10][946],u_xpb_out[11][946],u_xpb_out[12][946],u_xpb_out[13][946],u_xpb_out[14][946],u_xpb_out[15][946],u_xpb_out[16][946],u_xpb_out[17][946],u_xpb_out[18][946],u_xpb_out[19][946],u_xpb_out[20][946],u_xpb_out[21][946],u_xpb_out[22][946],u_xpb_out[23][946],u_xpb_out[24][946],u_xpb_out[25][946],u_xpb_out[26][946],u_xpb_out[27][946],u_xpb_out[28][946],u_xpb_out[29][946],u_xpb_out[30][946],u_xpb_out[31][946],u_xpb_out[32][946],u_xpb_out[33][946],u_xpb_out[34][946],u_xpb_out[35][946],u_xpb_out[36][946],u_xpb_out[37][946],u_xpb_out[38][946],u_xpb_out[39][946],u_xpb_out[40][946],u_xpb_out[41][946],u_xpb_out[42][946],u_xpb_out[43][946],u_xpb_out[44][946],u_xpb_out[45][946],u_xpb_out[46][946],u_xpb_out[47][946],u_xpb_out[48][946],u_xpb_out[49][946],u_xpb_out[50][946],u_xpb_out[51][946],u_xpb_out[52][946],u_xpb_out[53][946],u_xpb_out[54][946],u_xpb_out[55][946],u_xpb_out[56][946],u_xpb_out[57][946],u_xpb_out[58][946],u_xpb_out[59][946],u_xpb_out[60][946],u_xpb_out[61][946],u_xpb_out[62][946],u_xpb_out[63][946],u_xpb_out[64][946],u_xpb_out[65][946],u_xpb_out[66][946],u_xpb_out[67][946],u_xpb_out[68][946],u_xpb_out[69][946],u_xpb_out[70][946],u_xpb_out[71][946],u_xpb_out[72][946],u_xpb_out[73][946],u_xpb_out[74][946],u_xpb_out[75][946],u_xpb_out[76][946],u_xpb_out[77][946],u_xpb_out[78][946],u_xpb_out[79][946],u_xpb_out[80][946],u_xpb_out[81][946],u_xpb_out[82][946],u_xpb_out[83][946],u_xpb_out[84][946],u_xpb_out[85][946],u_xpb_out[86][946],u_xpb_out[87][946],u_xpb_out[88][946],u_xpb_out[89][946],u_xpb_out[90][946],u_xpb_out[91][946],u_xpb_out[92][946],u_xpb_out[93][946],u_xpb_out[94][946],u_xpb_out[95][946],u_xpb_out[96][946],u_xpb_out[97][946],u_xpb_out[98][946],u_xpb_out[99][946],u_xpb_out[100][946],u_xpb_out[101][946],u_xpb_out[102][946],u_xpb_out[103][946],u_xpb_out[104][946],u_xpb_out[105][946]};

assign col_out_947 = {u_xpb_out[0][947],u_xpb_out[1][947],u_xpb_out[2][947],u_xpb_out[3][947],u_xpb_out[4][947],u_xpb_out[5][947],u_xpb_out[6][947],u_xpb_out[7][947],u_xpb_out[8][947],u_xpb_out[9][947],u_xpb_out[10][947],u_xpb_out[11][947],u_xpb_out[12][947],u_xpb_out[13][947],u_xpb_out[14][947],u_xpb_out[15][947],u_xpb_out[16][947],u_xpb_out[17][947],u_xpb_out[18][947],u_xpb_out[19][947],u_xpb_out[20][947],u_xpb_out[21][947],u_xpb_out[22][947],u_xpb_out[23][947],u_xpb_out[24][947],u_xpb_out[25][947],u_xpb_out[26][947],u_xpb_out[27][947],u_xpb_out[28][947],u_xpb_out[29][947],u_xpb_out[30][947],u_xpb_out[31][947],u_xpb_out[32][947],u_xpb_out[33][947],u_xpb_out[34][947],u_xpb_out[35][947],u_xpb_out[36][947],u_xpb_out[37][947],u_xpb_out[38][947],u_xpb_out[39][947],u_xpb_out[40][947],u_xpb_out[41][947],u_xpb_out[42][947],u_xpb_out[43][947],u_xpb_out[44][947],u_xpb_out[45][947],u_xpb_out[46][947],u_xpb_out[47][947],u_xpb_out[48][947],u_xpb_out[49][947],u_xpb_out[50][947],u_xpb_out[51][947],u_xpb_out[52][947],u_xpb_out[53][947],u_xpb_out[54][947],u_xpb_out[55][947],u_xpb_out[56][947],u_xpb_out[57][947],u_xpb_out[58][947],u_xpb_out[59][947],u_xpb_out[60][947],u_xpb_out[61][947],u_xpb_out[62][947],u_xpb_out[63][947],u_xpb_out[64][947],u_xpb_out[65][947],u_xpb_out[66][947],u_xpb_out[67][947],u_xpb_out[68][947],u_xpb_out[69][947],u_xpb_out[70][947],u_xpb_out[71][947],u_xpb_out[72][947],u_xpb_out[73][947],u_xpb_out[74][947],u_xpb_out[75][947],u_xpb_out[76][947],u_xpb_out[77][947],u_xpb_out[78][947],u_xpb_out[79][947],u_xpb_out[80][947],u_xpb_out[81][947],u_xpb_out[82][947],u_xpb_out[83][947],u_xpb_out[84][947],u_xpb_out[85][947],u_xpb_out[86][947],u_xpb_out[87][947],u_xpb_out[88][947],u_xpb_out[89][947],u_xpb_out[90][947],u_xpb_out[91][947],u_xpb_out[92][947],u_xpb_out[93][947],u_xpb_out[94][947],u_xpb_out[95][947],u_xpb_out[96][947],u_xpb_out[97][947],u_xpb_out[98][947],u_xpb_out[99][947],u_xpb_out[100][947],u_xpb_out[101][947],u_xpb_out[102][947],u_xpb_out[103][947],u_xpb_out[104][947],u_xpb_out[105][947]};

assign col_out_948 = {u_xpb_out[0][948],u_xpb_out[1][948],u_xpb_out[2][948],u_xpb_out[3][948],u_xpb_out[4][948],u_xpb_out[5][948],u_xpb_out[6][948],u_xpb_out[7][948],u_xpb_out[8][948],u_xpb_out[9][948],u_xpb_out[10][948],u_xpb_out[11][948],u_xpb_out[12][948],u_xpb_out[13][948],u_xpb_out[14][948],u_xpb_out[15][948],u_xpb_out[16][948],u_xpb_out[17][948],u_xpb_out[18][948],u_xpb_out[19][948],u_xpb_out[20][948],u_xpb_out[21][948],u_xpb_out[22][948],u_xpb_out[23][948],u_xpb_out[24][948],u_xpb_out[25][948],u_xpb_out[26][948],u_xpb_out[27][948],u_xpb_out[28][948],u_xpb_out[29][948],u_xpb_out[30][948],u_xpb_out[31][948],u_xpb_out[32][948],u_xpb_out[33][948],u_xpb_out[34][948],u_xpb_out[35][948],u_xpb_out[36][948],u_xpb_out[37][948],u_xpb_out[38][948],u_xpb_out[39][948],u_xpb_out[40][948],u_xpb_out[41][948],u_xpb_out[42][948],u_xpb_out[43][948],u_xpb_out[44][948],u_xpb_out[45][948],u_xpb_out[46][948],u_xpb_out[47][948],u_xpb_out[48][948],u_xpb_out[49][948],u_xpb_out[50][948],u_xpb_out[51][948],u_xpb_out[52][948],u_xpb_out[53][948],u_xpb_out[54][948],u_xpb_out[55][948],u_xpb_out[56][948],u_xpb_out[57][948],u_xpb_out[58][948],u_xpb_out[59][948],u_xpb_out[60][948],u_xpb_out[61][948],u_xpb_out[62][948],u_xpb_out[63][948],u_xpb_out[64][948],u_xpb_out[65][948],u_xpb_out[66][948],u_xpb_out[67][948],u_xpb_out[68][948],u_xpb_out[69][948],u_xpb_out[70][948],u_xpb_out[71][948],u_xpb_out[72][948],u_xpb_out[73][948],u_xpb_out[74][948],u_xpb_out[75][948],u_xpb_out[76][948],u_xpb_out[77][948],u_xpb_out[78][948],u_xpb_out[79][948],u_xpb_out[80][948],u_xpb_out[81][948],u_xpb_out[82][948],u_xpb_out[83][948],u_xpb_out[84][948],u_xpb_out[85][948],u_xpb_out[86][948],u_xpb_out[87][948],u_xpb_out[88][948],u_xpb_out[89][948],u_xpb_out[90][948],u_xpb_out[91][948],u_xpb_out[92][948],u_xpb_out[93][948],u_xpb_out[94][948],u_xpb_out[95][948],u_xpb_out[96][948],u_xpb_out[97][948],u_xpb_out[98][948],u_xpb_out[99][948],u_xpb_out[100][948],u_xpb_out[101][948],u_xpb_out[102][948],u_xpb_out[103][948],u_xpb_out[104][948],u_xpb_out[105][948]};

assign col_out_949 = {u_xpb_out[0][949],u_xpb_out[1][949],u_xpb_out[2][949],u_xpb_out[3][949],u_xpb_out[4][949],u_xpb_out[5][949],u_xpb_out[6][949],u_xpb_out[7][949],u_xpb_out[8][949],u_xpb_out[9][949],u_xpb_out[10][949],u_xpb_out[11][949],u_xpb_out[12][949],u_xpb_out[13][949],u_xpb_out[14][949],u_xpb_out[15][949],u_xpb_out[16][949],u_xpb_out[17][949],u_xpb_out[18][949],u_xpb_out[19][949],u_xpb_out[20][949],u_xpb_out[21][949],u_xpb_out[22][949],u_xpb_out[23][949],u_xpb_out[24][949],u_xpb_out[25][949],u_xpb_out[26][949],u_xpb_out[27][949],u_xpb_out[28][949],u_xpb_out[29][949],u_xpb_out[30][949],u_xpb_out[31][949],u_xpb_out[32][949],u_xpb_out[33][949],u_xpb_out[34][949],u_xpb_out[35][949],u_xpb_out[36][949],u_xpb_out[37][949],u_xpb_out[38][949],u_xpb_out[39][949],u_xpb_out[40][949],u_xpb_out[41][949],u_xpb_out[42][949],u_xpb_out[43][949],u_xpb_out[44][949],u_xpb_out[45][949],u_xpb_out[46][949],u_xpb_out[47][949],u_xpb_out[48][949],u_xpb_out[49][949],u_xpb_out[50][949],u_xpb_out[51][949],u_xpb_out[52][949],u_xpb_out[53][949],u_xpb_out[54][949],u_xpb_out[55][949],u_xpb_out[56][949],u_xpb_out[57][949],u_xpb_out[58][949],u_xpb_out[59][949],u_xpb_out[60][949],u_xpb_out[61][949],u_xpb_out[62][949],u_xpb_out[63][949],u_xpb_out[64][949],u_xpb_out[65][949],u_xpb_out[66][949],u_xpb_out[67][949],u_xpb_out[68][949],u_xpb_out[69][949],u_xpb_out[70][949],u_xpb_out[71][949],u_xpb_out[72][949],u_xpb_out[73][949],u_xpb_out[74][949],u_xpb_out[75][949],u_xpb_out[76][949],u_xpb_out[77][949],u_xpb_out[78][949],u_xpb_out[79][949],u_xpb_out[80][949],u_xpb_out[81][949],u_xpb_out[82][949],u_xpb_out[83][949],u_xpb_out[84][949],u_xpb_out[85][949],u_xpb_out[86][949],u_xpb_out[87][949],u_xpb_out[88][949],u_xpb_out[89][949],u_xpb_out[90][949],u_xpb_out[91][949],u_xpb_out[92][949],u_xpb_out[93][949],u_xpb_out[94][949],u_xpb_out[95][949],u_xpb_out[96][949],u_xpb_out[97][949],u_xpb_out[98][949],u_xpb_out[99][949],u_xpb_out[100][949],u_xpb_out[101][949],u_xpb_out[102][949],u_xpb_out[103][949],u_xpb_out[104][949],u_xpb_out[105][949]};

assign col_out_950 = {u_xpb_out[0][950],u_xpb_out[1][950],u_xpb_out[2][950],u_xpb_out[3][950],u_xpb_out[4][950],u_xpb_out[5][950],u_xpb_out[6][950],u_xpb_out[7][950],u_xpb_out[8][950],u_xpb_out[9][950],u_xpb_out[10][950],u_xpb_out[11][950],u_xpb_out[12][950],u_xpb_out[13][950],u_xpb_out[14][950],u_xpb_out[15][950],u_xpb_out[16][950],u_xpb_out[17][950],u_xpb_out[18][950],u_xpb_out[19][950],u_xpb_out[20][950],u_xpb_out[21][950],u_xpb_out[22][950],u_xpb_out[23][950],u_xpb_out[24][950],u_xpb_out[25][950],u_xpb_out[26][950],u_xpb_out[27][950],u_xpb_out[28][950],u_xpb_out[29][950],u_xpb_out[30][950],u_xpb_out[31][950],u_xpb_out[32][950],u_xpb_out[33][950],u_xpb_out[34][950],u_xpb_out[35][950],u_xpb_out[36][950],u_xpb_out[37][950],u_xpb_out[38][950],u_xpb_out[39][950],u_xpb_out[40][950],u_xpb_out[41][950],u_xpb_out[42][950],u_xpb_out[43][950],u_xpb_out[44][950],u_xpb_out[45][950],u_xpb_out[46][950],u_xpb_out[47][950],u_xpb_out[48][950],u_xpb_out[49][950],u_xpb_out[50][950],u_xpb_out[51][950],u_xpb_out[52][950],u_xpb_out[53][950],u_xpb_out[54][950],u_xpb_out[55][950],u_xpb_out[56][950],u_xpb_out[57][950],u_xpb_out[58][950],u_xpb_out[59][950],u_xpb_out[60][950],u_xpb_out[61][950],u_xpb_out[62][950],u_xpb_out[63][950],u_xpb_out[64][950],u_xpb_out[65][950],u_xpb_out[66][950],u_xpb_out[67][950],u_xpb_out[68][950],u_xpb_out[69][950],u_xpb_out[70][950],u_xpb_out[71][950],u_xpb_out[72][950],u_xpb_out[73][950],u_xpb_out[74][950],u_xpb_out[75][950],u_xpb_out[76][950],u_xpb_out[77][950],u_xpb_out[78][950],u_xpb_out[79][950],u_xpb_out[80][950],u_xpb_out[81][950],u_xpb_out[82][950],u_xpb_out[83][950],u_xpb_out[84][950],u_xpb_out[85][950],u_xpb_out[86][950],u_xpb_out[87][950],u_xpb_out[88][950],u_xpb_out[89][950],u_xpb_out[90][950],u_xpb_out[91][950],u_xpb_out[92][950],u_xpb_out[93][950],u_xpb_out[94][950],u_xpb_out[95][950],u_xpb_out[96][950],u_xpb_out[97][950],u_xpb_out[98][950],u_xpb_out[99][950],u_xpb_out[100][950],u_xpb_out[101][950],u_xpb_out[102][950],u_xpb_out[103][950],u_xpb_out[104][950],u_xpb_out[105][950]};

assign col_out_951 = {u_xpb_out[0][951],u_xpb_out[1][951],u_xpb_out[2][951],u_xpb_out[3][951],u_xpb_out[4][951],u_xpb_out[5][951],u_xpb_out[6][951],u_xpb_out[7][951],u_xpb_out[8][951],u_xpb_out[9][951],u_xpb_out[10][951],u_xpb_out[11][951],u_xpb_out[12][951],u_xpb_out[13][951],u_xpb_out[14][951],u_xpb_out[15][951],u_xpb_out[16][951],u_xpb_out[17][951],u_xpb_out[18][951],u_xpb_out[19][951],u_xpb_out[20][951],u_xpb_out[21][951],u_xpb_out[22][951],u_xpb_out[23][951],u_xpb_out[24][951],u_xpb_out[25][951],u_xpb_out[26][951],u_xpb_out[27][951],u_xpb_out[28][951],u_xpb_out[29][951],u_xpb_out[30][951],u_xpb_out[31][951],u_xpb_out[32][951],u_xpb_out[33][951],u_xpb_out[34][951],u_xpb_out[35][951],u_xpb_out[36][951],u_xpb_out[37][951],u_xpb_out[38][951],u_xpb_out[39][951],u_xpb_out[40][951],u_xpb_out[41][951],u_xpb_out[42][951],u_xpb_out[43][951],u_xpb_out[44][951],u_xpb_out[45][951],u_xpb_out[46][951],u_xpb_out[47][951],u_xpb_out[48][951],u_xpb_out[49][951],u_xpb_out[50][951],u_xpb_out[51][951],u_xpb_out[52][951],u_xpb_out[53][951],u_xpb_out[54][951],u_xpb_out[55][951],u_xpb_out[56][951],u_xpb_out[57][951],u_xpb_out[58][951],u_xpb_out[59][951],u_xpb_out[60][951],u_xpb_out[61][951],u_xpb_out[62][951],u_xpb_out[63][951],u_xpb_out[64][951],u_xpb_out[65][951],u_xpb_out[66][951],u_xpb_out[67][951],u_xpb_out[68][951],u_xpb_out[69][951],u_xpb_out[70][951],u_xpb_out[71][951],u_xpb_out[72][951],u_xpb_out[73][951],u_xpb_out[74][951],u_xpb_out[75][951],u_xpb_out[76][951],u_xpb_out[77][951],u_xpb_out[78][951],u_xpb_out[79][951],u_xpb_out[80][951],u_xpb_out[81][951],u_xpb_out[82][951],u_xpb_out[83][951],u_xpb_out[84][951],u_xpb_out[85][951],u_xpb_out[86][951],u_xpb_out[87][951],u_xpb_out[88][951],u_xpb_out[89][951],u_xpb_out[90][951],u_xpb_out[91][951],u_xpb_out[92][951],u_xpb_out[93][951],u_xpb_out[94][951],u_xpb_out[95][951],u_xpb_out[96][951],u_xpb_out[97][951],u_xpb_out[98][951],u_xpb_out[99][951],u_xpb_out[100][951],u_xpb_out[101][951],u_xpb_out[102][951],u_xpb_out[103][951],u_xpb_out[104][951],u_xpb_out[105][951]};

assign col_out_952 = {u_xpb_out[0][952],u_xpb_out[1][952],u_xpb_out[2][952],u_xpb_out[3][952],u_xpb_out[4][952],u_xpb_out[5][952],u_xpb_out[6][952],u_xpb_out[7][952],u_xpb_out[8][952],u_xpb_out[9][952],u_xpb_out[10][952],u_xpb_out[11][952],u_xpb_out[12][952],u_xpb_out[13][952],u_xpb_out[14][952],u_xpb_out[15][952],u_xpb_out[16][952],u_xpb_out[17][952],u_xpb_out[18][952],u_xpb_out[19][952],u_xpb_out[20][952],u_xpb_out[21][952],u_xpb_out[22][952],u_xpb_out[23][952],u_xpb_out[24][952],u_xpb_out[25][952],u_xpb_out[26][952],u_xpb_out[27][952],u_xpb_out[28][952],u_xpb_out[29][952],u_xpb_out[30][952],u_xpb_out[31][952],u_xpb_out[32][952],u_xpb_out[33][952],u_xpb_out[34][952],u_xpb_out[35][952],u_xpb_out[36][952],u_xpb_out[37][952],u_xpb_out[38][952],u_xpb_out[39][952],u_xpb_out[40][952],u_xpb_out[41][952],u_xpb_out[42][952],u_xpb_out[43][952],u_xpb_out[44][952],u_xpb_out[45][952],u_xpb_out[46][952],u_xpb_out[47][952],u_xpb_out[48][952],u_xpb_out[49][952],u_xpb_out[50][952],u_xpb_out[51][952],u_xpb_out[52][952],u_xpb_out[53][952],u_xpb_out[54][952],u_xpb_out[55][952],u_xpb_out[56][952],u_xpb_out[57][952],u_xpb_out[58][952],u_xpb_out[59][952],u_xpb_out[60][952],u_xpb_out[61][952],u_xpb_out[62][952],u_xpb_out[63][952],u_xpb_out[64][952],u_xpb_out[65][952],u_xpb_out[66][952],u_xpb_out[67][952],u_xpb_out[68][952],u_xpb_out[69][952],u_xpb_out[70][952],u_xpb_out[71][952],u_xpb_out[72][952],u_xpb_out[73][952],u_xpb_out[74][952],u_xpb_out[75][952],u_xpb_out[76][952],u_xpb_out[77][952],u_xpb_out[78][952],u_xpb_out[79][952],u_xpb_out[80][952],u_xpb_out[81][952],u_xpb_out[82][952],u_xpb_out[83][952],u_xpb_out[84][952],u_xpb_out[85][952],u_xpb_out[86][952],u_xpb_out[87][952],u_xpb_out[88][952],u_xpb_out[89][952],u_xpb_out[90][952],u_xpb_out[91][952],u_xpb_out[92][952],u_xpb_out[93][952],u_xpb_out[94][952],u_xpb_out[95][952],u_xpb_out[96][952],u_xpb_out[97][952],u_xpb_out[98][952],u_xpb_out[99][952],u_xpb_out[100][952],u_xpb_out[101][952],u_xpb_out[102][952],u_xpb_out[103][952],u_xpb_out[104][952],u_xpb_out[105][952]};

assign col_out_953 = {u_xpb_out[0][953],u_xpb_out[1][953],u_xpb_out[2][953],u_xpb_out[3][953],u_xpb_out[4][953],u_xpb_out[5][953],u_xpb_out[6][953],u_xpb_out[7][953],u_xpb_out[8][953],u_xpb_out[9][953],u_xpb_out[10][953],u_xpb_out[11][953],u_xpb_out[12][953],u_xpb_out[13][953],u_xpb_out[14][953],u_xpb_out[15][953],u_xpb_out[16][953],u_xpb_out[17][953],u_xpb_out[18][953],u_xpb_out[19][953],u_xpb_out[20][953],u_xpb_out[21][953],u_xpb_out[22][953],u_xpb_out[23][953],u_xpb_out[24][953],u_xpb_out[25][953],u_xpb_out[26][953],u_xpb_out[27][953],u_xpb_out[28][953],u_xpb_out[29][953],u_xpb_out[30][953],u_xpb_out[31][953],u_xpb_out[32][953],u_xpb_out[33][953],u_xpb_out[34][953],u_xpb_out[35][953],u_xpb_out[36][953],u_xpb_out[37][953],u_xpb_out[38][953],u_xpb_out[39][953],u_xpb_out[40][953],u_xpb_out[41][953],u_xpb_out[42][953],u_xpb_out[43][953],u_xpb_out[44][953],u_xpb_out[45][953],u_xpb_out[46][953],u_xpb_out[47][953],u_xpb_out[48][953],u_xpb_out[49][953],u_xpb_out[50][953],u_xpb_out[51][953],u_xpb_out[52][953],u_xpb_out[53][953],u_xpb_out[54][953],u_xpb_out[55][953],u_xpb_out[56][953],u_xpb_out[57][953],u_xpb_out[58][953],u_xpb_out[59][953],u_xpb_out[60][953],u_xpb_out[61][953],u_xpb_out[62][953],u_xpb_out[63][953],u_xpb_out[64][953],u_xpb_out[65][953],u_xpb_out[66][953],u_xpb_out[67][953],u_xpb_out[68][953],u_xpb_out[69][953],u_xpb_out[70][953],u_xpb_out[71][953],u_xpb_out[72][953],u_xpb_out[73][953],u_xpb_out[74][953],u_xpb_out[75][953],u_xpb_out[76][953],u_xpb_out[77][953],u_xpb_out[78][953],u_xpb_out[79][953],u_xpb_out[80][953],u_xpb_out[81][953],u_xpb_out[82][953],u_xpb_out[83][953],u_xpb_out[84][953],u_xpb_out[85][953],u_xpb_out[86][953],u_xpb_out[87][953],u_xpb_out[88][953],u_xpb_out[89][953],u_xpb_out[90][953],u_xpb_out[91][953],u_xpb_out[92][953],u_xpb_out[93][953],u_xpb_out[94][953],u_xpb_out[95][953],u_xpb_out[96][953],u_xpb_out[97][953],u_xpb_out[98][953],u_xpb_out[99][953],u_xpb_out[100][953],u_xpb_out[101][953],u_xpb_out[102][953],u_xpb_out[103][953],u_xpb_out[104][953],u_xpb_out[105][953]};

assign col_out_954 = {u_xpb_out[0][954],u_xpb_out[1][954],u_xpb_out[2][954],u_xpb_out[3][954],u_xpb_out[4][954],u_xpb_out[5][954],u_xpb_out[6][954],u_xpb_out[7][954],u_xpb_out[8][954],u_xpb_out[9][954],u_xpb_out[10][954],u_xpb_out[11][954],u_xpb_out[12][954],u_xpb_out[13][954],u_xpb_out[14][954],u_xpb_out[15][954],u_xpb_out[16][954],u_xpb_out[17][954],u_xpb_out[18][954],u_xpb_out[19][954],u_xpb_out[20][954],u_xpb_out[21][954],u_xpb_out[22][954],u_xpb_out[23][954],u_xpb_out[24][954],u_xpb_out[25][954],u_xpb_out[26][954],u_xpb_out[27][954],u_xpb_out[28][954],u_xpb_out[29][954],u_xpb_out[30][954],u_xpb_out[31][954],u_xpb_out[32][954],u_xpb_out[33][954],u_xpb_out[34][954],u_xpb_out[35][954],u_xpb_out[36][954],u_xpb_out[37][954],u_xpb_out[38][954],u_xpb_out[39][954],u_xpb_out[40][954],u_xpb_out[41][954],u_xpb_out[42][954],u_xpb_out[43][954],u_xpb_out[44][954],u_xpb_out[45][954],u_xpb_out[46][954],u_xpb_out[47][954],u_xpb_out[48][954],u_xpb_out[49][954],u_xpb_out[50][954],u_xpb_out[51][954],u_xpb_out[52][954],u_xpb_out[53][954],u_xpb_out[54][954],u_xpb_out[55][954],u_xpb_out[56][954],u_xpb_out[57][954],u_xpb_out[58][954],u_xpb_out[59][954],u_xpb_out[60][954],u_xpb_out[61][954],u_xpb_out[62][954],u_xpb_out[63][954],u_xpb_out[64][954],u_xpb_out[65][954],u_xpb_out[66][954],u_xpb_out[67][954],u_xpb_out[68][954],u_xpb_out[69][954],u_xpb_out[70][954],u_xpb_out[71][954],u_xpb_out[72][954],u_xpb_out[73][954],u_xpb_out[74][954],u_xpb_out[75][954],u_xpb_out[76][954],u_xpb_out[77][954],u_xpb_out[78][954],u_xpb_out[79][954],u_xpb_out[80][954],u_xpb_out[81][954],u_xpb_out[82][954],u_xpb_out[83][954],u_xpb_out[84][954],u_xpb_out[85][954],u_xpb_out[86][954],u_xpb_out[87][954],u_xpb_out[88][954],u_xpb_out[89][954],u_xpb_out[90][954],u_xpb_out[91][954],u_xpb_out[92][954],u_xpb_out[93][954],u_xpb_out[94][954],u_xpb_out[95][954],u_xpb_out[96][954],u_xpb_out[97][954],u_xpb_out[98][954],u_xpb_out[99][954],u_xpb_out[100][954],u_xpb_out[101][954],u_xpb_out[102][954],u_xpb_out[103][954],u_xpb_out[104][954],u_xpb_out[105][954]};

assign col_out_955 = {u_xpb_out[0][955],u_xpb_out[1][955],u_xpb_out[2][955],u_xpb_out[3][955],u_xpb_out[4][955],u_xpb_out[5][955],u_xpb_out[6][955],u_xpb_out[7][955],u_xpb_out[8][955],u_xpb_out[9][955],u_xpb_out[10][955],u_xpb_out[11][955],u_xpb_out[12][955],u_xpb_out[13][955],u_xpb_out[14][955],u_xpb_out[15][955],u_xpb_out[16][955],u_xpb_out[17][955],u_xpb_out[18][955],u_xpb_out[19][955],u_xpb_out[20][955],u_xpb_out[21][955],u_xpb_out[22][955],u_xpb_out[23][955],u_xpb_out[24][955],u_xpb_out[25][955],u_xpb_out[26][955],u_xpb_out[27][955],u_xpb_out[28][955],u_xpb_out[29][955],u_xpb_out[30][955],u_xpb_out[31][955],u_xpb_out[32][955],u_xpb_out[33][955],u_xpb_out[34][955],u_xpb_out[35][955],u_xpb_out[36][955],u_xpb_out[37][955],u_xpb_out[38][955],u_xpb_out[39][955],u_xpb_out[40][955],u_xpb_out[41][955],u_xpb_out[42][955],u_xpb_out[43][955],u_xpb_out[44][955],u_xpb_out[45][955],u_xpb_out[46][955],u_xpb_out[47][955],u_xpb_out[48][955],u_xpb_out[49][955],u_xpb_out[50][955],u_xpb_out[51][955],u_xpb_out[52][955],u_xpb_out[53][955],u_xpb_out[54][955],u_xpb_out[55][955],u_xpb_out[56][955],u_xpb_out[57][955],u_xpb_out[58][955],u_xpb_out[59][955],u_xpb_out[60][955],u_xpb_out[61][955],u_xpb_out[62][955],u_xpb_out[63][955],u_xpb_out[64][955],u_xpb_out[65][955],u_xpb_out[66][955],u_xpb_out[67][955],u_xpb_out[68][955],u_xpb_out[69][955],u_xpb_out[70][955],u_xpb_out[71][955],u_xpb_out[72][955],u_xpb_out[73][955],u_xpb_out[74][955],u_xpb_out[75][955],u_xpb_out[76][955],u_xpb_out[77][955],u_xpb_out[78][955],u_xpb_out[79][955],u_xpb_out[80][955],u_xpb_out[81][955],u_xpb_out[82][955],u_xpb_out[83][955],u_xpb_out[84][955],u_xpb_out[85][955],u_xpb_out[86][955],u_xpb_out[87][955],u_xpb_out[88][955],u_xpb_out[89][955],u_xpb_out[90][955],u_xpb_out[91][955],u_xpb_out[92][955],u_xpb_out[93][955],u_xpb_out[94][955],u_xpb_out[95][955],u_xpb_out[96][955],u_xpb_out[97][955],u_xpb_out[98][955],u_xpb_out[99][955],u_xpb_out[100][955],u_xpb_out[101][955],u_xpb_out[102][955],u_xpb_out[103][955],u_xpb_out[104][955],u_xpb_out[105][955]};

assign col_out_956 = {u_xpb_out[0][956],u_xpb_out[1][956],u_xpb_out[2][956],u_xpb_out[3][956],u_xpb_out[4][956],u_xpb_out[5][956],u_xpb_out[6][956],u_xpb_out[7][956],u_xpb_out[8][956],u_xpb_out[9][956],u_xpb_out[10][956],u_xpb_out[11][956],u_xpb_out[12][956],u_xpb_out[13][956],u_xpb_out[14][956],u_xpb_out[15][956],u_xpb_out[16][956],u_xpb_out[17][956],u_xpb_out[18][956],u_xpb_out[19][956],u_xpb_out[20][956],u_xpb_out[21][956],u_xpb_out[22][956],u_xpb_out[23][956],u_xpb_out[24][956],u_xpb_out[25][956],u_xpb_out[26][956],u_xpb_out[27][956],u_xpb_out[28][956],u_xpb_out[29][956],u_xpb_out[30][956],u_xpb_out[31][956],u_xpb_out[32][956],u_xpb_out[33][956],u_xpb_out[34][956],u_xpb_out[35][956],u_xpb_out[36][956],u_xpb_out[37][956],u_xpb_out[38][956],u_xpb_out[39][956],u_xpb_out[40][956],u_xpb_out[41][956],u_xpb_out[42][956],u_xpb_out[43][956],u_xpb_out[44][956],u_xpb_out[45][956],u_xpb_out[46][956],u_xpb_out[47][956],u_xpb_out[48][956],u_xpb_out[49][956],u_xpb_out[50][956],u_xpb_out[51][956],u_xpb_out[52][956],u_xpb_out[53][956],u_xpb_out[54][956],u_xpb_out[55][956],u_xpb_out[56][956],u_xpb_out[57][956],u_xpb_out[58][956],u_xpb_out[59][956],u_xpb_out[60][956],u_xpb_out[61][956],u_xpb_out[62][956],u_xpb_out[63][956],u_xpb_out[64][956],u_xpb_out[65][956],u_xpb_out[66][956],u_xpb_out[67][956],u_xpb_out[68][956],u_xpb_out[69][956],u_xpb_out[70][956],u_xpb_out[71][956],u_xpb_out[72][956],u_xpb_out[73][956],u_xpb_out[74][956],u_xpb_out[75][956],u_xpb_out[76][956],u_xpb_out[77][956],u_xpb_out[78][956],u_xpb_out[79][956],u_xpb_out[80][956],u_xpb_out[81][956],u_xpb_out[82][956],u_xpb_out[83][956],u_xpb_out[84][956],u_xpb_out[85][956],u_xpb_out[86][956],u_xpb_out[87][956],u_xpb_out[88][956],u_xpb_out[89][956],u_xpb_out[90][956],u_xpb_out[91][956],u_xpb_out[92][956],u_xpb_out[93][956],u_xpb_out[94][956],u_xpb_out[95][956],u_xpb_out[96][956],u_xpb_out[97][956],u_xpb_out[98][956],u_xpb_out[99][956],u_xpb_out[100][956],u_xpb_out[101][956],u_xpb_out[102][956],u_xpb_out[103][956],u_xpb_out[104][956],u_xpb_out[105][956]};

assign col_out_957 = {u_xpb_out[0][957],u_xpb_out[1][957],u_xpb_out[2][957],u_xpb_out[3][957],u_xpb_out[4][957],u_xpb_out[5][957],u_xpb_out[6][957],u_xpb_out[7][957],u_xpb_out[8][957],u_xpb_out[9][957],u_xpb_out[10][957],u_xpb_out[11][957],u_xpb_out[12][957],u_xpb_out[13][957],u_xpb_out[14][957],u_xpb_out[15][957],u_xpb_out[16][957],u_xpb_out[17][957],u_xpb_out[18][957],u_xpb_out[19][957],u_xpb_out[20][957],u_xpb_out[21][957],u_xpb_out[22][957],u_xpb_out[23][957],u_xpb_out[24][957],u_xpb_out[25][957],u_xpb_out[26][957],u_xpb_out[27][957],u_xpb_out[28][957],u_xpb_out[29][957],u_xpb_out[30][957],u_xpb_out[31][957],u_xpb_out[32][957],u_xpb_out[33][957],u_xpb_out[34][957],u_xpb_out[35][957],u_xpb_out[36][957],u_xpb_out[37][957],u_xpb_out[38][957],u_xpb_out[39][957],u_xpb_out[40][957],u_xpb_out[41][957],u_xpb_out[42][957],u_xpb_out[43][957],u_xpb_out[44][957],u_xpb_out[45][957],u_xpb_out[46][957],u_xpb_out[47][957],u_xpb_out[48][957],u_xpb_out[49][957],u_xpb_out[50][957],u_xpb_out[51][957],u_xpb_out[52][957],u_xpb_out[53][957],u_xpb_out[54][957],u_xpb_out[55][957],u_xpb_out[56][957],u_xpb_out[57][957],u_xpb_out[58][957],u_xpb_out[59][957],u_xpb_out[60][957],u_xpb_out[61][957],u_xpb_out[62][957],u_xpb_out[63][957],u_xpb_out[64][957],u_xpb_out[65][957],u_xpb_out[66][957],u_xpb_out[67][957],u_xpb_out[68][957],u_xpb_out[69][957],u_xpb_out[70][957],u_xpb_out[71][957],u_xpb_out[72][957],u_xpb_out[73][957],u_xpb_out[74][957],u_xpb_out[75][957],u_xpb_out[76][957],u_xpb_out[77][957],u_xpb_out[78][957],u_xpb_out[79][957],u_xpb_out[80][957],u_xpb_out[81][957],u_xpb_out[82][957],u_xpb_out[83][957],u_xpb_out[84][957],u_xpb_out[85][957],u_xpb_out[86][957],u_xpb_out[87][957],u_xpb_out[88][957],u_xpb_out[89][957],u_xpb_out[90][957],u_xpb_out[91][957],u_xpb_out[92][957],u_xpb_out[93][957],u_xpb_out[94][957],u_xpb_out[95][957],u_xpb_out[96][957],u_xpb_out[97][957],u_xpb_out[98][957],u_xpb_out[99][957],u_xpb_out[100][957],u_xpb_out[101][957],u_xpb_out[102][957],u_xpb_out[103][957],u_xpb_out[104][957],u_xpb_out[105][957]};

assign col_out_958 = {u_xpb_out[0][958],u_xpb_out[1][958],u_xpb_out[2][958],u_xpb_out[3][958],u_xpb_out[4][958],u_xpb_out[5][958],u_xpb_out[6][958],u_xpb_out[7][958],u_xpb_out[8][958],u_xpb_out[9][958],u_xpb_out[10][958],u_xpb_out[11][958],u_xpb_out[12][958],u_xpb_out[13][958],u_xpb_out[14][958],u_xpb_out[15][958],u_xpb_out[16][958],u_xpb_out[17][958],u_xpb_out[18][958],u_xpb_out[19][958],u_xpb_out[20][958],u_xpb_out[21][958],u_xpb_out[22][958],u_xpb_out[23][958],u_xpb_out[24][958],u_xpb_out[25][958],u_xpb_out[26][958],u_xpb_out[27][958],u_xpb_out[28][958],u_xpb_out[29][958],u_xpb_out[30][958],u_xpb_out[31][958],u_xpb_out[32][958],u_xpb_out[33][958],u_xpb_out[34][958],u_xpb_out[35][958],u_xpb_out[36][958],u_xpb_out[37][958],u_xpb_out[38][958],u_xpb_out[39][958],u_xpb_out[40][958],u_xpb_out[41][958],u_xpb_out[42][958],u_xpb_out[43][958],u_xpb_out[44][958],u_xpb_out[45][958],u_xpb_out[46][958],u_xpb_out[47][958],u_xpb_out[48][958],u_xpb_out[49][958],u_xpb_out[50][958],u_xpb_out[51][958],u_xpb_out[52][958],u_xpb_out[53][958],u_xpb_out[54][958],u_xpb_out[55][958],u_xpb_out[56][958],u_xpb_out[57][958],u_xpb_out[58][958],u_xpb_out[59][958],u_xpb_out[60][958],u_xpb_out[61][958],u_xpb_out[62][958],u_xpb_out[63][958],u_xpb_out[64][958],u_xpb_out[65][958],u_xpb_out[66][958],u_xpb_out[67][958],u_xpb_out[68][958],u_xpb_out[69][958],u_xpb_out[70][958],u_xpb_out[71][958],u_xpb_out[72][958],u_xpb_out[73][958],u_xpb_out[74][958],u_xpb_out[75][958],u_xpb_out[76][958],u_xpb_out[77][958],u_xpb_out[78][958],u_xpb_out[79][958],u_xpb_out[80][958],u_xpb_out[81][958],u_xpb_out[82][958],u_xpb_out[83][958],u_xpb_out[84][958],u_xpb_out[85][958],u_xpb_out[86][958],u_xpb_out[87][958],u_xpb_out[88][958],u_xpb_out[89][958],u_xpb_out[90][958],u_xpb_out[91][958],u_xpb_out[92][958],u_xpb_out[93][958],u_xpb_out[94][958],u_xpb_out[95][958],u_xpb_out[96][958],u_xpb_out[97][958],u_xpb_out[98][958],u_xpb_out[99][958],u_xpb_out[100][958],u_xpb_out[101][958],u_xpb_out[102][958],u_xpb_out[103][958],u_xpb_out[104][958],u_xpb_out[105][958]};

assign col_out_959 = {u_xpb_out[0][959],u_xpb_out[1][959],u_xpb_out[2][959],u_xpb_out[3][959],u_xpb_out[4][959],u_xpb_out[5][959],u_xpb_out[6][959],u_xpb_out[7][959],u_xpb_out[8][959],u_xpb_out[9][959],u_xpb_out[10][959],u_xpb_out[11][959],u_xpb_out[12][959],u_xpb_out[13][959],u_xpb_out[14][959],u_xpb_out[15][959],u_xpb_out[16][959],u_xpb_out[17][959],u_xpb_out[18][959],u_xpb_out[19][959],u_xpb_out[20][959],u_xpb_out[21][959],u_xpb_out[22][959],u_xpb_out[23][959],u_xpb_out[24][959],u_xpb_out[25][959],u_xpb_out[26][959],u_xpb_out[27][959],u_xpb_out[28][959],u_xpb_out[29][959],u_xpb_out[30][959],u_xpb_out[31][959],u_xpb_out[32][959],u_xpb_out[33][959],u_xpb_out[34][959],u_xpb_out[35][959],u_xpb_out[36][959],u_xpb_out[37][959],u_xpb_out[38][959],u_xpb_out[39][959],u_xpb_out[40][959],u_xpb_out[41][959],u_xpb_out[42][959],u_xpb_out[43][959],u_xpb_out[44][959],u_xpb_out[45][959],u_xpb_out[46][959],u_xpb_out[47][959],u_xpb_out[48][959],u_xpb_out[49][959],u_xpb_out[50][959],u_xpb_out[51][959],u_xpb_out[52][959],u_xpb_out[53][959],u_xpb_out[54][959],u_xpb_out[55][959],u_xpb_out[56][959],u_xpb_out[57][959],u_xpb_out[58][959],u_xpb_out[59][959],u_xpb_out[60][959],u_xpb_out[61][959],u_xpb_out[62][959],u_xpb_out[63][959],u_xpb_out[64][959],u_xpb_out[65][959],u_xpb_out[66][959],u_xpb_out[67][959],u_xpb_out[68][959],u_xpb_out[69][959],u_xpb_out[70][959],u_xpb_out[71][959],u_xpb_out[72][959],u_xpb_out[73][959],u_xpb_out[74][959],u_xpb_out[75][959],u_xpb_out[76][959],u_xpb_out[77][959],u_xpb_out[78][959],u_xpb_out[79][959],u_xpb_out[80][959],u_xpb_out[81][959],u_xpb_out[82][959],u_xpb_out[83][959],u_xpb_out[84][959],u_xpb_out[85][959],u_xpb_out[86][959],u_xpb_out[87][959],u_xpb_out[88][959],u_xpb_out[89][959],u_xpb_out[90][959],u_xpb_out[91][959],u_xpb_out[92][959],u_xpb_out[93][959],u_xpb_out[94][959],u_xpb_out[95][959],u_xpb_out[96][959],u_xpb_out[97][959],u_xpb_out[98][959],u_xpb_out[99][959],u_xpb_out[100][959],u_xpb_out[101][959],u_xpb_out[102][959],u_xpb_out[103][959],u_xpb_out[104][959],u_xpb_out[105][959]};

assign col_out_960 = {u_xpb_out[0][960],u_xpb_out[1][960],u_xpb_out[2][960],u_xpb_out[3][960],u_xpb_out[4][960],u_xpb_out[5][960],u_xpb_out[6][960],u_xpb_out[7][960],u_xpb_out[8][960],u_xpb_out[9][960],u_xpb_out[10][960],u_xpb_out[11][960],u_xpb_out[12][960],u_xpb_out[13][960],u_xpb_out[14][960],u_xpb_out[15][960],u_xpb_out[16][960],u_xpb_out[17][960],u_xpb_out[18][960],u_xpb_out[19][960],u_xpb_out[20][960],u_xpb_out[21][960],u_xpb_out[22][960],u_xpb_out[23][960],u_xpb_out[24][960],u_xpb_out[25][960],u_xpb_out[26][960],u_xpb_out[27][960],u_xpb_out[28][960],u_xpb_out[29][960],u_xpb_out[30][960],u_xpb_out[31][960],u_xpb_out[32][960],u_xpb_out[33][960],u_xpb_out[34][960],u_xpb_out[35][960],u_xpb_out[36][960],u_xpb_out[37][960],u_xpb_out[38][960],u_xpb_out[39][960],u_xpb_out[40][960],u_xpb_out[41][960],u_xpb_out[42][960],u_xpb_out[43][960],u_xpb_out[44][960],u_xpb_out[45][960],u_xpb_out[46][960],u_xpb_out[47][960],u_xpb_out[48][960],u_xpb_out[49][960],u_xpb_out[50][960],u_xpb_out[51][960],u_xpb_out[52][960],u_xpb_out[53][960],u_xpb_out[54][960],u_xpb_out[55][960],u_xpb_out[56][960],u_xpb_out[57][960],u_xpb_out[58][960],u_xpb_out[59][960],u_xpb_out[60][960],u_xpb_out[61][960],u_xpb_out[62][960],u_xpb_out[63][960],u_xpb_out[64][960],u_xpb_out[65][960],u_xpb_out[66][960],u_xpb_out[67][960],u_xpb_out[68][960],u_xpb_out[69][960],u_xpb_out[70][960],u_xpb_out[71][960],u_xpb_out[72][960],u_xpb_out[73][960],u_xpb_out[74][960],u_xpb_out[75][960],u_xpb_out[76][960],u_xpb_out[77][960],u_xpb_out[78][960],u_xpb_out[79][960],u_xpb_out[80][960],u_xpb_out[81][960],u_xpb_out[82][960],u_xpb_out[83][960],u_xpb_out[84][960],u_xpb_out[85][960],u_xpb_out[86][960],u_xpb_out[87][960],u_xpb_out[88][960],u_xpb_out[89][960],u_xpb_out[90][960],u_xpb_out[91][960],u_xpb_out[92][960],u_xpb_out[93][960],u_xpb_out[94][960],u_xpb_out[95][960],u_xpb_out[96][960],u_xpb_out[97][960],u_xpb_out[98][960],u_xpb_out[99][960],u_xpb_out[100][960],u_xpb_out[101][960],u_xpb_out[102][960],u_xpb_out[103][960],u_xpb_out[104][960],u_xpb_out[105][960]};

assign col_out_961 = {u_xpb_out[0][961],u_xpb_out[1][961],u_xpb_out[2][961],u_xpb_out[3][961],u_xpb_out[4][961],u_xpb_out[5][961],u_xpb_out[6][961],u_xpb_out[7][961],u_xpb_out[8][961],u_xpb_out[9][961],u_xpb_out[10][961],u_xpb_out[11][961],u_xpb_out[12][961],u_xpb_out[13][961],u_xpb_out[14][961],u_xpb_out[15][961],u_xpb_out[16][961],u_xpb_out[17][961],u_xpb_out[18][961],u_xpb_out[19][961],u_xpb_out[20][961],u_xpb_out[21][961],u_xpb_out[22][961],u_xpb_out[23][961],u_xpb_out[24][961],u_xpb_out[25][961],u_xpb_out[26][961],u_xpb_out[27][961],u_xpb_out[28][961],u_xpb_out[29][961],u_xpb_out[30][961],u_xpb_out[31][961],u_xpb_out[32][961],u_xpb_out[33][961],u_xpb_out[34][961],u_xpb_out[35][961],u_xpb_out[36][961],u_xpb_out[37][961],u_xpb_out[38][961],u_xpb_out[39][961],u_xpb_out[40][961],u_xpb_out[41][961],u_xpb_out[42][961],u_xpb_out[43][961],u_xpb_out[44][961],u_xpb_out[45][961],u_xpb_out[46][961],u_xpb_out[47][961],u_xpb_out[48][961],u_xpb_out[49][961],u_xpb_out[50][961],u_xpb_out[51][961],u_xpb_out[52][961],u_xpb_out[53][961],u_xpb_out[54][961],u_xpb_out[55][961],u_xpb_out[56][961],u_xpb_out[57][961],u_xpb_out[58][961],u_xpb_out[59][961],u_xpb_out[60][961],u_xpb_out[61][961],u_xpb_out[62][961],u_xpb_out[63][961],u_xpb_out[64][961],u_xpb_out[65][961],u_xpb_out[66][961],u_xpb_out[67][961],u_xpb_out[68][961],u_xpb_out[69][961],u_xpb_out[70][961],u_xpb_out[71][961],u_xpb_out[72][961],u_xpb_out[73][961],u_xpb_out[74][961],u_xpb_out[75][961],u_xpb_out[76][961],u_xpb_out[77][961],u_xpb_out[78][961],u_xpb_out[79][961],u_xpb_out[80][961],u_xpb_out[81][961],u_xpb_out[82][961],u_xpb_out[83][961],u_xpb_out[84][961],u_xpb_out[85][961],u_xpb_out[86][961],u_xpb_out[87][961],u_xpb_out[88][961],u_xpb_out[89][961],u_xpb_out[90][961],u_xpb_out[91][961],u_xpb_out[92][961],u_xpb_out[93][961],u_xpb_out[94][961],u_xpb_out[95][961],u_xpb_out[96][961],u_xpb_out[97][961],u_xpb_out[98][961],u_xpb_out[99][961],u_xpb_out[100][961],u_xpb_out[101][961],u_xpb_out[102][961],u_xpb_out[103][961],u_xpb_out[104][961],u_xpb_out[105][961]};

assign col_out_962 = {u_xpb_out[0][962],u_xpb_out[1][962],u_xpb_out[2][962],u_xpb_out[3][962],u_xpb_out[4][962],u_xpb_out[5][962],u_xpb_out[6][962],u_xpb_out[7][962],u_xpb_out[8][962],u_xpb_out[9][962],u_xpb_out[10][962],u_xpb_out[11][962],u_xpb_out[12][962],u_xpb_out[13][962],u_xpb_out[14][962],u_xpb_out[15][962],u_xpb_out[16][962],u_xpb_out[17][962],u_xpb_out[18][962],u_xpb_out[19][962],u_xpb_out[20][962],u_xpb_out[21][962],u_xpb_out[22][962],u_xpb_out[23][962],u_xpb_out[24][962],u_xpb_out[25][962],u_xpb_out[26][962],u_xpb_out[27][962],u_xpb_out[28][962],u_xpb_out[29][962],u_xpb_out[30][962],u_xpb_out[31][962],u_xpb_out[32][962],u_xpb_out[33][962],u_xpb_out[34][962],u_xpb_out[35][962],u_xpb_out[36][962],u_xpb_out[37][962],u_xpb_out[38][962],u_xpb_out[39][962],u_xpb_out[40][962],u_xpb_out[41][962],u_xpb_out[42][962],u_xpb_out[43][962],u_xpb_out[44][962],u_xpb_out[45][962],u_xpb_out[46][962],u_xpb_out[47][962],u_xpb_out[48][962],u_xpb_out[49][962],u_xpb_out[50][962],u_xpb_out[51][962],u_xpb_out[52][962],u_xpb_out[53][962],u_xpb_out[54][962],u_xpb_out[55][962],u_xpb_out[56][962],u_xpb_out[57][962],u_xpb_out[58][962],u_xpb_out[59][962],u_xpb_out[60][962],u_xpb_out[61][962],u_xpb_out[62][962],u_xpb_out[63][962],u_xpb_out[64][962],u_xpb_out[65][962],u_xpb_out[66][962],u_xpb_out[67][962],u_xpb_out[68][962],u_xpb_out[69][962],u_xpb_out[70][962],u_xpb_out[71][962],u_xpb_out[72][962],u_xpb_out[73][962],u_xpb_out[74][962],u_xpb_out[75][962],u_xpb_out[76][962],u_xpb_out[77][962],u_xpb_out[78][962],u_xpb_out[79][962],u_xpb_out[80][962],u_xpb_out[81][962],u_xpb_out[82][962],u_xpb_out[83][962],u_xpb_out[84][962],u_xpb_out[85][962],u_xpb_out[86][962],u_xpb_out[87][962],u_xpb_out[88][962],u_xpb_out[89][962],u_xpb_out[90][962],u_xpb_out[91][962],u_xpb_out[92][962],u_xpb_out[93][962],u_xpb_out[94][962],u_xpb_out[95][962],u_xpb_out[96][962],u_xpb_out[97][962],u_xpb_out[98][962],u_xpb_out[99][962],u_xpb_out[100][962],u_xpb_out[101][962],u_xpb_out[102][962],u_xpb_out[103][962],u_xpb_out[104][962],u_xpb_out[105][962]};

assign col_out_963 = {u_xpb_out[0][963],u_xpb_out[1][963],u_xpb_out[2][963],u_xpb_out[3][963],u_xpb_out[4][963],u_xpb_out[5][963],u_xpb_out[6][963],u_xpb_out[7][963],u_xpb_out[8][963],u_xpb_out[9][963],u_xpb_out[10][963],u_xpb_out[11][963],u_xpb_out[12][963],u_xpb_out[13][963],u_xpb_out[14][963],u_xpb_out[15][963],u_xpb_out[16][963],u_xpb_out[17][963],u_xpb_out[18][963],u_xpb_out[19][963],u_xpb_out[20][963],u_xpb_out[21][963],u_xpb_out[22][963],u_xpb_out[23][963],u_xpb_out[24][963],u_xpb_out[25][963],u_xpb_out[26][963],u_xpb_out[27][963],u_xpb_out[28][963],u_xpb_out[29][963],u_xpb_out[30][963],u_xpb_out[31][963],u_xpb_out[32][963],u_xpb_out[33][963],u_xpb_out[34][963],u_xpb_out[35][963],u_xpb_out[36][963],u_xpb_out[37][963],u_xpb_out[38][963],u_xpb_out[39][963],u_xpb_out[40][963],u_xpb_out[41][963],u_xpb_out[42][963],u_xpb_out[43][963],u_xpb_out[44][963],u_xpb_out[45][963],u_xpb_out[46][963],u_xpb_out[47][963],u_xpb_out[48][963],u_xpb_out[49][963],u_xpb_out[50][963],u_xpb_out[51][963],u_xpb_out[52][963],u_xpb_out[53][963],u_xpb_out[54][963],u_xpb_out[55][963],u_xpb_out[56][963],u_xpb_out[57][963],u_xpb_out[58][963],u_xpb_out[59][963],u_xpb_out[60][963],u_xpb_out[61][963],u_xpb_out[62][963],u_xpb_out[63][963],u_xpb_out[64][963],u_xpb_out[65][963],u_xpb_out[66][963],u_xpb_out[67][963],u_xpb_out[68][963],u_xpb_out[69][963],u_xpb_out[70][963],u_xpb_out[71][963],u_xpb_out[72][963],u_xpb_out[73][963],u_xpb_out[74][963],u_xpb_out[75][963],u_xpb_out[76][963],u_xpb_out[77][963],u_xpb_out[78][963],u_xpb_out[79][963],u_xpb_out[80][963],u_xpb_out[81][963],u_xpb_out[82][963],u_xpb_out[83][963],u_xpb_out[84][963],u_xpb_out[85][963],u_xpb_out[86][963],u_xpb_out[87][963],u_xpb_out[88][963],u_xpb_out[89][963],u_xpb_out[90][963],u_xpb_out[91][963],u_xpb_out[92][963],u_xpb_out[93][963],u_xpb_out[94][963],u_xpb_out[95][963],u_xpb_out[96][963],u_xpb_out[97][963],u_xpb_out[98][963],u_xpb_out[99][963],u_xpb_out[100][963],u_xpb_out[101][963],u_xpb_out[102][963],u_xpb_out[103][963],u_xpb_out[104][963],u_xpb_out[105][963]};

assign col_out_964 = {u_xpb_out[0][964],u_xpb_out[1][964],u_xpb_out[2][964],u_xpb_out[3][964],u_xpb_out[4][964],u_xpb_out[5][964],u_xpb_out[6][964],u_xpb_out[7][964],u_xpb_out[8][964],u_xpb_out[9][964],u_xpb_out[10][964],u_xpb_out[11][964],u_xpb_out[12][964],u_xpb_out[13][964],u_xpb_out[14][964],u_xpb_out[15][964],u_xpb_out[16][964],u_xpb_out[17][964],u_xpb_out[18][964],u_xpb_out[19][964],u_xpb_out[20][964],u_xpb_out[21][964],u_xpb_out[22][964],u_xpb_out[23][964],u_xpb_out[24][964],u_xpb_out[25][964],u_xpb_out[26][964],u_xpb_out[27][964],u_xpb_out[28][964],u_xpb_out[29][964],u_xpb_out[30][964],u_xpb_out[31][964],u_xpb_out[32][964],u_xpb_out[33][964],u_xpb_out[34][964],u_xpb_out[35][964],u_xpb_out[36][964],u_xpb_out[37][964],u_xpb_out[38][964],u_xpb_out[39][964],u_xpb_out[40][964],u_xpb_out[41][964],u_xpb_out[42][964],u_xpb_out[43][964],u_xpb_out[44][964],u_xpb_out[45][964],u_xpb_out[46][964],u_xpb_out[47][964],u_xpb_out[48][964],u_xpb_out[49][964],u_xpb_out[50][964],u_xpb_out[51][964],u_xpb_out[52][964],u_xpb_out[53][964],u_xpb_out[54][964],u_xpb_out[55][964],u_xpb_out[56][964],u_xpb_out[57][964],u_xpb_out[58][964],u_xpb_out[59][964],u_xpb_out[60][964],u_xpb_out[61][964],u_xpb_out[62][964],u_xpb_out[63][964],u_xpb_out[64][964],u_xpb_out[65][964],u_xpb_out[66][964],u_xpb_out[67][964],u_xpb_out[68][964],u_xpb_out[69][964],u_xpb_out[70][964],u_xpb_out[71][964],u_xpb_out[72][964],u_xpb_out[73][964],u_xpb_out[74][964],u_xpb_out[75][964],u_xpb_out[76][964],u_xpb_out[77][964],u_xpb_out[78][964],u_xpb_out[79][964],u_xpb_out[80][964],u_xpb_out[81][964],u_xpb_out[82][964],u_xpb_out[83][964],u_xpb_out[84][964],u_xpb_out[85][964],u_xpb_out[86][964],u_xpb_out[87][964],u_xpb_out[88][964],u_xpb_out[89][964],u_xpb_out[90][964],u_xpb_out[91][964],u_xpb_out[92][964],u_xpb_out[93][964],u_xpb_out[94][964],u_xpb_out[95][964],u_xpb_out[96][964],u_xpb_out[97][964],u_xpb_out[98][964],u_xpb_out[99][964],u_xpb_out[100][964],u_xpb_out[101][964],u_xpb_out[102][964],u_xpb_out[103][964],u_xpb_out[104][964],u_xpb_out[105][964]};

assign col_out_965 = {u_xpb_out[0][965],u_xpb_out[1][965],u_xpb_out[2][965],u_xpb_out[3][965],u_xpb_out[4][965],u_xpb_out[5][965],u_xpb_out[6][965],u_xpb_out[7][965],u_xpb_out[8][965],u_xpb_out[9][965],u_xpb_out[10][965],u_xpb_out[11][965],u_xpb_out[12][965],u_xpb_out[13][965],u_xpb_out[14][965],u_xpb_out[15][965],u_xpb_out[16][965],u_xpb_out[17][965],u_xpb_out[18][965],u_xpb_out[19][965],u_xpb_out[20][965],u_xpb_out[21][965],u_xpb_out[22][965],u_xpb_out[23][965],u_xpb_out[24][965],u_xpb_out[25][965],u_xpb_out[26][965],u_xpb_out[27][965],u_xpb_out[28][965],u_xpb_out[29][965],u_xpb_out[30][965],u_xpb_out[31][965],u_xpb_out[32][965],u_xpb_out[33][965],u_xpb_out[34][965],u_xpb_out[35][965],u_xpb_out[36][965],u_xpb_out[37][965],u_xpb_out[38][965],u_xpb_out[39][965],u_xpb_out[40][965],u_xpb_out[41][965],u_xpb_out[42][965],u_xpb_out[43][965],u_xpb_out[44][965],u_xpb_out[45][965],u_xpb_out[46][965],u_xpb_out[47][965],u_xpb_out[48][965],u_xpb_out[49][965],u_xpb_out[50][965],u_xpb_out[51][965],u_xpb_out[52][965],u_xpb_out[53][965],u_xpb_out[54][965],u_xpb_out[55][965],u_xpb_out[56][965],u_xpb_out[57][965],u_xpb_out[58][965],u_xpb_out[59][965],u_xpb_out[60][965],u_xpb_out[61][965],u_xpb_out[62][965],u_xpb_out[63][965],u_xpb_out[64][965],u_xpb_out[65][965],u_xpb_out[66][965],u_xpb_out[67][965],u_xpb_out[68][965],u_xpb_out[69][965],u_xpb_out[70][965],u_xpb_out[71][965],u_xpb_out[72][965],u_xpb_out[73][965],u_xpb_out[74][965],u_xpb_out[75][965],u_xpb_out[76][965],u_xpb_out[77][965],u_xpb_out[78][965],u_xpb_out[79][965],u_xpb_out[80][965],u_xpb_out[81][965],u_xpb_out[82][965],u_xpb_out[83][965],u_xpb_out[84][965],u_xpb_out[85][965],u_xpb_out[86][965],u_xpb_out[87][965],u_xpb_out[88][965],u_xpb_out[89][965],u_xpb_out[90][965],u_xpb_out[91][965],u_xpb_out[92][965],u_xpb_out[93][965],u_xpb_out[94][965],u_xpb_out[95][965],u_xpb_out[96][965],u_xpb_out[97][965],u_xpb_out[98][965],u_xpb_out[99][965],u_xpb_out[100][965],u_xpb_out[101][965],u_xpb_out[102][965],u_xpb_out[103][965],u_xpb_out[104][965],u_xpb_out[105][965]};

assign col_out_966 = {u_xpb_out[0][966],u_xpb_out[1][966],u_xpb_out[2][966],u_xpb_out[3][966],u_xpb_out[4][966],u_xpb_out[5][966],u_xpb_out[6][966],u_xpb_out[7][966],u_xpb_out[8][966],u_xpb_out[9][966],u_xpb_out[10][966],u_xpb_out[11][966],u_xpb_out[12][966],u_xpb_out[13][966],u_xpb_out[14][966],u_xpb_out[15][966],u_xpb_out[16][966],u_xpb_out[17][966],u_xpb_out[18][966],u_xpb_out[19][966],u_xpb_out[20][966],u_xpb_out[21][966],u_xpb_out[22][966],u_xpb_out[23][966],u_xpb_out[24][966],u_xpb_out[25][966],u_xpb_out[26][966],u_xpb_out[27][966],u_xpb_out[28][966],u_xpb_out[29][966],u_xpb_out[30][966],u_xpb_out[31][966],u_xpb_out[32][966],u_xpb_out[33][966],u_xpb_out[34][966],u_xpb_out[35][966],u_xpb_out[36][966],u_xpb_out[37][966],u_xpb_out[38][966],u_xpb_out[39][966],u_xpb_out[40][966],u_xpb_out[41][966],u_xpb_out[42][966],u_xpb_out[43][966],u_xpb_out[44][966],u_xpb_out[45][966],u_xpb_out[46][966],u_xpb_out[47][966],u_xpb_out[48][966],u_xpb_out[49][966],u_xpb_out[50][966],u_xpb_out[51][966],u_xpb_out[52][966],u_xpb_out[53][966],u_xpb_out[54][966],u_xpb_out[55][966],u_xpb_out[56][966],u_xpb_out[57][966],u_xpb_out[58][966],u_xpb_out[59][966],u_xpb_out[60][966],u_xpb_out[61][966],u_xpb_out[62][966],u_xpb_out[63][966],u_xpb_out[64][966],u_xpb_out[65][966],u_xpb_out[66][966],u_xpb_out[67][966],u_xpb_out[68][966],u_xpb_out[69][966],u_xpb_out[70][966],u_xpb_out[71][966],u_xpb_out[72][966],u_xpb_out[73][966],u_xpb_out[74][966],u_xpb_out[75][966],u_xpb_out[76][966],u_xpb_out[77][966],u_xpb_out[78][966],u_xpb_out[79][966],u_xpb_out[80][966],u_xpb_out[81][966],u_xpb_out[82][966],u_xpb_out[83][966],u_xpb_out[84][966],u_xpb_out[85][966],u_xpb_out[86][966],u_xpb_out[87][966],u_xpb_out[88][966],u_xpb_out[89][966],u_xpb_out[90][966],u_xpb_out[91][966],u_xpb_out[92][966],u_xpb_out[93][966],u_xpb_out[94][966],u_xpb_out[95][966],u_xpb_out[96][966],u_xpb_out[97][966],u_xpb_out[98][966],u_xpb_out[99][966],u_xpb_out[100][966],u_xpb_out[101][966],u_xpb_out[102][966],u_xpb_out[103][966],u_xpb_out[104][966],u_xpb_out[105][966]};

assign col_out_967 = {u_xpb_out[0][967],u_xpb_out[1][967],u_xpb_out[2][967],u_xpb_out[3][967],u_xpb_out[4][967],u_xpb_out[5][967],u_xpb_out[6][967],u_xpb_out[7][967],u_xpb_out[8][967],u_xpb_out[9][967],u_xpb_out[10][967],u_xpb_out[11][967],u_xpb_out[12][967],u_xpb_out[13][967],u_xpb_out[14][967],u_xpb_out[15][967],u_xpb_out[16][967],u_xpb_out[17][967],u_xpb_out[18][967],u_xpb_out[19][967],u_xpb_out[20][967],u_xpb_out[21][967],u_xpb_out[22][967],u_xpb_out[23][967],u_xpb_out[24][967],u_xpb_out[25][967],u_xpb_out[26][967],u_xpb_out[27][967],u_xpb_out[28][967],u_xpb_out[29][967],u_xpb_out[30][967],u_xpb_out[31][967],u_xpb_out[32][967],u_xpb_out[33][967],u_xpb_out[34][967],u_xpb_out[35][967],u_xpb_out[36][967],u_xpb_out[37][967],u_xpb_out[38][967],u_xpb_out[39][967],u_xpb_out[40][967],u_xpb_out[41][967],u_xpb_out[42][967],u_xpb_out[43][967],u_xpb_out[44][967],u_xpb_out[45][967],u_xpb_out[46][967],u_xpb_out[47][967],u_xpb_out[48][967],u_xpb_out[49][967],u_xpb_out[50][967],u_xpb_out[51][967],u_xpb_out[52][967],u_xpb_out[53][967],u_xpb_out[54][967],u_xpb_out[55][967],u_xpb_out[56][967],u_xpb_out[57][967],u_xpb_out[58][967],u_xpb_out[59][967],u_xpb_out[60][967],u_xpb_out[61][967],u_xpb_out[62][967],u_xpb_out[63][967],u_xpb_out[64][967],u_xpb_out[65][967],u_xpb_out[66][967],u_xpb_out[67][967],u_xpb_out[68][967],u_xpb_out[69][967],u_xpb_out[70][967],u_xpb_out[71][967],u_xpb_out[72][967],u_xpb_out[73][967],u_xpb_out[74][967],u_xpb_out[75][967],u_xpb_out[76][967],u_xpb_out[77][967],u_xpb_out[78][967],u_xpb_out[79][967],u_xpb_out[80][967],u_xpb_out[81][967],u_xpb_out[82][967],u_xpb_out[83][967],u_xpb_out[84][967],u_xpb_out[85][967],u_xpb_out[86][967],u_xpb_out[87][967],u_xpb_out[88][967],u_xpb_out[89][967],u_xpb_out[90][967],u_xpb_out[91][967],u_xpb_out[92][967],u_xpb_out[93][967],u_xpb_out[94][967],u_xpb_out[95][967],u_xpb_out[96][967],u_xpb_out[97][967],u_xpb_out[98][967],u_xpb_out[99][967],u_xpb_out[100][967],u_xpb_out[101][967],u_xpb_out[102][967],u_xpb_out[103][967],u_xpb_out[104][967],u_xpb_out[105][967]};

assign col_out_968 = {u_xpb_out[0][968],u_xpb_out[1][968],u_xpb_out[2][968],u_xpb_out[3][968],u_xpb_out[4][968],u_xpb_out[5][968],u_xpb_out[6][968],u_xpb_out[7][968],u_xpb_out[8][968],u_xpb_out[9][968],u_xpb_out[10][968],u_xpb_out[11][968],u_xpb_out[12][968],u_xpb_out[13][968],u_xpb_out[14][968],u_xpb_out[15][968],u_xpb_out[16][968],u_xpb_out[17][968],u_xpb_out[18][968],u_xpb_out[19][968],u_xpb_out[20][968],u_xpb_out[21][968],u_xpb_out[22][968],u_xpb_out[23][968],u_xpb_out[24][968],u_xpb_out[25][968],u_xpb_out[26][968],u_xpb_out[27][968],u_xpb_out[28][968],u_xpb_out[29][968],u_xpb_out[30][968],u_xpb_out[31][968],u_xpb_out[32][968],u_xpb_out[33][968],u_xpb_out[34][968],u_xpb_out[35][968],u_xpb_out[36][968],u_xpb_out[37][968],u_xpb_out[38][968],u_xpb_out[39][968],u_xpb_out[40][968],u_xpb_out[41][968],u_xpb_out[42][968],u_xpb_out[43][968],u_xpb_out[44][968],u_xpb_out[45][968],u_xpb_out[46][968],u_xpb_out[47][968],u_xpb_out[48][968],u_xpb_out[49][968],u_xpb_out[50][968],u_xpb_out[51][968],u_xpb_out[52][968],u_xpb_out[53][968],u_xpb_out[54][968],u_xpb_out[55][968],u_xpb_out[56][968],u_xpb_out[57][968],u_xpb_out[58][968],u_xpb_out[59][968],u_xpb_out[60][968],u_xpb_out[61][968],u_xpb_out[62][968],u_xpb_out[63][968],u_xpb_out[64][968],u_xpb_out[65][968],u_xpb_out[66][968],u_xpb_out[67][968],u_xpb_out[68][968],u_xpb_out[69][968],u_xpb_out[70][968],u_xpb_out[71][968],u_xpb_out[72][968],u_xpb_out[73][968],u_xpb_out[74][968],u_xpb_out[75][968],u_xpb_out[76][968],u_xpb_out[77][968],u_xpb_out[78][968],u_xpb_out[79][968],u_xpb_out[80][968],u_xpb_out[81][968],u_xpb_out[82][968],u_xpb_out[83][968],u_xpb_out[84][968],u_xpb_out[85][968],u_xpb_out[86][968],u_xpb_out[87][968],u_xpb_out[88][968],u_xpb_out[89][968],u_xpb_out[90][968],u_xpb_out[91][968],u_xpb_out[92][968],u_xpb_out[93][968],u_xpb_out[94][968],u_xpb_out[95][968],u_xpb_out[96][968],u_xpb_out[97][968],u_xpb_out[98][968],u_xpb_out[99][968],u_xpb_out[100][968],u_xpb_out[101][968],u_xpb_out[102][968],u_xpb_out[103][968],u_xpb_out[104][968],u_xpb_out[105][968]};

assign col_out_969 = {u_xpb_out[0][969],u_xpb_out[1][969],u_xpb_out[2][969],u_xpb_out[3][969],u_xpb_out[4][969],u_xpb_out[5][969],u_xpb_out[6][969],u_xpb_out[7][969],u_xpb_out[8][969],u_xpb_out[9][969],u_xpb_out[10][969],u_xpb_out[11][969],u_xpb_out[12][969],u_xpb_out[13][969],u_xpb_out[14][969],u_xpb_out[15][969],u_xpb_out[16][969],u_xpb_out[17][969],u_xpb_out[18][969],u_xpb_out[19][969],u_xpb_out[20][969],u_xpb_out[21][969],u_xpb_out[22][969],u_xpb_out[23][969],u_xpb_out[24][969],u_xpb_out[25][969],u_xpb_out[26][969],u_xpb_out[27][969],u_xpb_out[28][969],u_xpb_out[29][969],u_xpb_out[30][969],u_xpb_out[31][969],u_xpb_out[32][969],u_xpb_out[33][969],u_xpb_out[34][969],u_xpb_out[35][969],u_xpb_out[36][969],u_xpb_out[37][969],u_xpb_out[38][969],u_xpb_out[39][969],u_xpb_out[40][969],u_xpb_out[41][969],u_xpb_out[42][969],u_xpb_out[43][969],u_xpb_out[44][969],u_xpb_out[45][969],u_xpb_out[46][969],u_xpb_out[47][969],u_xpb_out[48][969],u_xpb_out[49][969],u_xpb_out[50][969],u_xpb_out[51][969],u_xpb_out[52][969],u_xpb_out[53][969],u_xpb_out[54][969],u_xpb_out[55][969],u_xpb_out[56][969],u_xpb_out[57][969],u_xpb_out[58][969],u_xpb_out[59][969],u_xpb_out[60][969],u_xpb_out[61][969],u_xpb_out[62][969],u_xpb_out[63][969],u_xpb_out[64][969],u_xpb_out[65][969],u_xpb_out[66][969],u_xpb_out[67][969],u_xpb_out[68][969],u_xpb_out[69][969],u_xpb_out[70][969],u_xpb_out[71][969],u_xpb_out[72][969],u_xpb_out[73][969],u_xpb_out[74][969],u_xpb_out[75][969],u_xpb_out[76][969],u_xpb_out[77][969],u_xpb_out[78][969],u_xpb_out[79][969],u_xpb_out[80][969],u_xpb_out[81][969],u_xpb_out[82][969],u_xpb_out[83][969],u_xpb_out[84][969],u_xpb_out[85][969],u_xpb_out[86][969],u_xpb_out[87][969],u_xpb_out[88][969],u_xpb_out[89][969],u_xpb_out[90][969],u_xpb_out[91][969],u_xpb_out[92][969],u_xpb_out[93][969],u_xpb_out[94][969],u_xpb_out[95][969],u_xpb_out[96][969],u_xpb_out[97][969],u_xpb_out[98][969],u_xpb_out[99][969],u_xpb_out[100][969],u_xpb_out[101][969],u_xpb_out[102][969],u_xpb_out[103][969],u_xpb_out[104][969],u_xpb_out[105][969]};

assign col_out_970 = {u_xpb_out[0][970],u_xpb_out[1][970],u_xpb_out[2][970],u_xpb_out[3][970],u_xpb_out[4][970],u_xpb_out[5][970],u_xpb_out[6][970],u_xpb_out[7][970],u_xpb_out[8][970],u_xpb_out[9][970],u_xpb_out[10][970],u_xpb_out[11][970],u_xpb_out[12][970],u_xpb_out[13][970],u_xpb_out[14][970],u_xpb_out[15][970],u_xpb_out[16][970],u_xpb_out[17][970],u_xpb_out[18][970],u_xpb_out[19][970],u_xpb_out[20][970],u_xpb_out[21][970],u_xpb_out[22][970],u_xpb_out[23][970],u_xpb_out[24][970],u_xpb_out[25][970],u_xpb_out[26][970],u_xpb_out[27][970],u_xpb_out[28][970],u_xpb_out[29][970],u_xpb_out[30][970],u_xpb_out[31][970],u_xpb_out[32][970],u_xpb_out[33][970],u_xpb_out[34][970],u_xpb_out[35][970],u_xpb_out[36][970],u_xpb_out[37][970],u_xpb_out[38][970],u_xpb_out[39][970],u_xpb_out[40][970],u_xpb_out[41][970],u_xpb_out[42][970],u_xpb_out[43][970],u_xpb_out[44][970],u_xpb_out[45][970],u_xpb_out[46][970],u_xpb_out[47][970],u_xpb_out[48][970],u_xpb_out[49][970],u_xpb_out[50][970],u_xpb_out[51][970],u_xpb_out[52][970],u_xpb_out[53][970],u_xpb_out[54][970],u_xpb_out[55][970],u_xpb_out[56][970],u_xpb_out[57][970],u_xpb_out[58][970],u_xpb_out[59][970],u_xpb_out[60][970],u_xpb_out[61][970],u_xpb_out[62][970],u_xpb_out[63][970],u_xpb_out[64][970],u_xpb_out[65][970],u_xpb_out[66][970],u_xpb_out[67][970],u_xpb_out[68][970],u_xpb_out[69][970],u_xpb_out[70][970],u_xpb_out[71][970],u_xpb_out[72][970],u_xpb_out[73][970],u_xpb_out[74][970],u_xpb_out[75][970],u_xpb_out[76][970],u_xpb_out[77][970],u_xpb_out[78][970],u_xpb_out[79][970],u_xpb_out[80][970],u_xpb_out[81][970],u_xpb_out[82][970],u_xpb_out[83][970],u_xpb_out[84][970],u_xpb_out[85][970],u_xpb_out[86][970],u_xpb_out[87][970],u_xpb_out[88][970],u_xpb_out[89][970],u_xpb_out[90][970],u_xpb_out[91][970],u_xpb_out[92][970],u_xpb_out[93][970],u_xpb_out[94][970],u_xpb_out[95][970],u_xpb_out[96][970],u_xpb_out[97][970],u_xpb_out[98][970],u_xpb_out[99][970],u_xpb_out[100][970],u_xpb_out[101][970],u_xpb_out[102][970],u_xpb_out[103][970],u_xpb_out[104][970],u_xpb_out[105][970]};

assign col_out_971 = {u_xpb_out[0][971],u_xpb_out[1][971],u_xpb_out[2][971],u_xpb_out[3][971],u_xpb_out[4][971],u_xpb_out[5][971],u_xpb_out[6][971],u_xpb_out[7][971],u_xpb_out[8][971],u_xpb_out[9][971],u_xpb_out[10][971],u_xpb_out[11][971],u_xpb_out[12][971],u_xpb_out[13][971],u_xpb_out[14][971],u_xpb_out[15][971],u_xpb_out[16][971],u_xpb_out[17][971],u_xpb_out[18][971],u_xpb_out[19][971],u_xpb_out[20][971],u_xpb_out[21][971],u_xpb_out[22][971],u_xpb_out[23][971],u_xpb_out[24][971],u_xpb_out[25][971],u_xpb_out[26][971],u_xpb_out[27][971],u_xpb_out[28][971],u_xpb_out[29][971],u_xpb_out[30][971],u_xpb_out[31][971],u_xpb_out[32][971],u_xpb_out[33][971],u_xpb_out[34][971],u_xpb_out[35][971],u_xpb_out[36][971],u_xpb_out[37][971],u_xpb_out[38][971],u_xpb_out[39][971],u_xpb_out[40][971],u_xpb_out[41][971],u_xpb_out[42][971],u_xpb_out[43][971],u_xpb_out[44][971],u_xpb_out[45][971],u_xpb_out[46][971],u_xpb_out[47][971],u_xpb_out[48][971],u_xpb_out[49][971],u_xpb_out[50][971],u_xpb_out[51][971],u_xpb_out[52][971],u_xpb_out[53][971],u_xpb_out[54][971],u_xpb_out[55][971],u_xpb_out[56][971],u_xpb_out[57][971],u_xpb_out[58][971],u_xpb_out[59][971],u_xpb_out[60][971],u_xpb_out[61][971],u_xpb_out[62][971],u_xpb_out[63][971],u_xpb_out[64][971],u_xpb_out[65][971],u_xpb_out[66][971],u_xpb_out[67][971],u_xpb_out[68][971],u_xpb_out[69][971],u_xpb_out[70][971],u_xpb_out[71][971],u_xpb_out[72][971],u_xpb_out[73][971],u_xpb_out[74][971],u_xpb_out[75][971],u_xpb_out[76][971],u_xpb_out[77][971],u_xpb_out[78][971],u_xpb_out[79][971],u_xpb_out[80][971],u_xpb_out[81][971],u_xpb_out[82][971],u_xpb_out[83][971],u_xpb_out[84][971],u_xpb_out[85][971],u_xpb_out[86][971],u_xpb_out[87][971],u_xpb_out[88][971],u_xpb_out[89][971],u_xpb_out[90][971],u_xpb_out[91][971],u_xpb_out[92][971],u_xpb_out[93][971],u_xpb_out[94][971],u_xpb_out[95][971],u_xpb_out[96][971],u_xpb_out[97][971],u_xpb_out[98][971],u_xpb_out[99][971],u_xpb_out[100][971],u_xpb_out[101][971],u_xpb_out[102][971],u_xpb_out[103][971],u_xpb_out[104][971],u_xpb_out[105][971]};

assign col_out_972 = {u_xpb_out[0][972],u_xpb_out[1][972],u_xpb_out[2][972],u_xpb_out[3][972],u_xpb_out[4][972],u_xpb_out[5][972],u_xpb_out[6][972],u_xpb_out[7][972],u_xpb_out[8][972],u_xpb_out[9][972],u_xpb_out[10][972],u_xpb_out[11][972],u_xpb_out[12][972],u_xpb_out[13][972],u_xpb_out[14][972],u_xpb_out[15][972],u_xpb_out[16][972],u_xpb_out[17][972],u_xpb_out[18][972],u_xpb_out[19][972],u_xpb_out[20][972],u_xpb_out[21][972],u_xpb_out[22][972],u_xpb_out[23][972],u_xpb_out[24][972],u_xpb_out[25][972],u_xpb_out[26][972],u_xpb_out[27][972],u_xpb_out[28][972],u_xpb_out[29][972],u_xpb_out[30][972],u_xpb_out[31][972],u_xpb_out[32][972],u_xpb_out[33][972],u_xpb_out[34][972],u_xpb_out[35][972],u_xpb_out[36][972],u_xpb_out[37][972],u_xpb_out[38][972],u_xpb_out[39][972],u_xpb_out[40][972],u_xpb_out[41][972],u_xpb_out[42][972],u_xpb_out[43][972],u_xpb_out[44][972],u_xpb_out[45][972],u_xpb_out[46][972],u_xpb_out[47][972],u_xpb_out[48][972],u_xpb_out[49][972],u_xpb_out[50][972],u_xpb_out[51][972],u_xpb_out[52][972],u_xpb_out[53][972],u_xpb_out[54][972],u_xpb_out[55][972],u_xpb_out[56][972],u_xpb_out[57][972],u_xpb_out[58][972],u_xpb_out[59][972],u_xpb_out[60][972],u_xpb_out[61][972],u_xpb_out[62][972],u_xpb_out[63][972],u_xpb_out[64][972],u_xpb_out[65][972],u_xpb_out[66][972],u_xpb_out[67][972],u_xpb_out[68][972],u_xpb_out[69][972],u_xpb_out[70][972],u_xpb_out[71][972],u_xpb_out[72][972],u_xpb_out[73][972],u_xpb_out[74][972],u_xpb_out[75][972],u_xpb_out[76][972],u_xpb_out[77][972],u_xpb_out[78][972],u_xpb_out[79][972],u_xpb_out[80][972],u_xpb_out[81][972],u_xpb_out[82][972],u_xpb_out[83][972],u_xpb_out[84][972],u_xpb_out[85][972],u_xpb_out[86][972],u_xpb_out[87][972],u_xpb_out[88][972],u_xpb_out[89][972],u_xpb_out[90][972],u_xpb_out[91][972],u_xpb_out[92][972],u_xpb_out[93][972],u_xpb_out[94][972],u_xpb_out[95][972],u_xpb_out[96][972],u_xpb_out[97][972],u_xpb_out[98][972],u_xpb_out[99][972],u_xpb_out[100][972],u_xpb_out[101][972],u_xpb_out[102][972],u_xpb_out[103][972],u_xpb_out[104][972],u_xpb_out[105][972]};

assign col_out_973 = {u_xpb_out[0][973],u_xpb_out[1][973],u_xpb_out[2][973],u_xpb_out[3][973],u_xpb_out[4][973],u_xpb_out[5][973],u_xpb_out[6][973],u_xpb_out[7][973],u_xpb_out[8][973],u_xpb_out[9][973],u_xpb_out[10][973],u_xpb_out[11][973],u_xpb_out[12][973],u_xpb_out[13][973],u_xpb_out[14][973],u_xpb_out[15][973],u_xpb_out[16][973],u_xpb_out[17][973],u_xpb_out[18][973],u_xpb_out[19][973],u_xpb_out[20][973],u_xpb_out[21][973],u_xpb_out[22][973],u_xpb_out[23][973],u_xpb_out[24][973],u_xpb_out[25][973],u_xpb_out[26][973],u_xpb_out[27][973],u_xpb_out[28][973],u_xpb_out[29][973],u_xpb_out[30][973],u_xpb_out[31][973],u_xpb_out[32][973],u_xpb_out[33][973],u_xpb_out[34][973],u_xpb_out[35][973],u_xpb_out[36][973],u_xpb_out[37][973],u_xpb_out[38][973],u_xpb_out[39][973],u_xpb_out[40][973],u_xpb_out[41][973],u_xpb_out[42][973],u_xpb_out[43][973],u_xpb_out[44][973],u_xpb_out[45][973],u_xpb_out[46][973],u_xpb_out[47][973],u_xpb_out[48][973],u_xpb_out[49][973],u_xpb_out[50][973],u_xpb_out[51][973],u_xpb_out[52][973],u_xpb_out[53][973],u_xpb_out[54][973],u_xpb_out[55][973],u_xpb_out[56][973],u_xpb_out[57][973],u_xpb_out[58][973],u_xpb_out[59][973],u_xpb_out[60][973],u_xpb_out[61][973],u_xpb_out[62][973],u_xpb_out[63][973],u_xpb_out[64][973],u_xpb_out[65][973],u_xpb_out[66][973],u_xpb_out[67][973],u_xpb_out[68][973],u_xpb_out[69][973],u_xpb_out[70][973],u_xpb_out[71][973],u_xpb_out[72][973],u_xpb_out[73][973],u_xpb_out[74][973],u_xpb_out[75][973],u_xpb_out[76][973],u_xpb_out[77][973],u_xpb_out[78][973],u_xpb_out[79][973],u_xpb_out[80][973],u_xpb_out[81][973],u_xpb_out[82][973],u_xpb_out[83][973],u_xpb_out[84][973],u_xpb_out[85][973],u_xpb_out[86][973],u_xpb_out[87][973],u_xpb_out[88][973],u_xpb_out[89][973],u_xpb_out[90][973],u_xpb_out[91][973],u_xpb_out[92][973],u_xpb_out[93][973],u_xpb_out[94][973],u_xpb_out[95][973],u_xpb_out[96][973],u_xpb_out[97][973],u_xpb_out[98][973],u_xpb_out[99][973],u_xpb_out[100][973],u_xpb_out[101][973],u_xpb_out[102][973],u_xpb_out[103][973],u_xpb_out[104][973],u_xpb_out[105][973]};

assign col_out_974 = {u_xpb_out[0][974],u_xpb_out[1][974],u_xpb_out[2][974],u_xpb_out[3][974],u_xpb_out[4][974],u_xpb_out[5][974],u_xpb_out[6][974],u_xpb_out[7][974],u_xpb_out[8][974],u_xpb_out[9][974],u_xpb_out[10][974],u_xpb_out[11][974],u_xpb_out[12][974],u_xpb_out[13][974],u_xpb_out[14][974],u_xpb_out[15][974],u_xpb_out[16][974],u_xpb_out[17][974],u_xpb_out[18][974],u_xpb_out[19][974],u_xpb_out[20][974],u_xpb_out[21][974],u_xpb_out[22][974],u_xpb_out[23][974],u_xpb_out[24][974],u_xpb_out[25][974],u_xpb_out[26][974],u_xpb_out[27][974],u_xpb_out[28][974],u_xpb_out[29][974],u_xpb_out[30][974],u_xpb_out[31][974],u_xpb_out[32][974],u_xpb_out[33][974],u_xpb_out[34][974],u_xpb_out[35][974],u_xpb_out[36][974],u_xpb_out[37][974],u_xpb_out[38][974],u_xpb_out[39][974],u_xpb_out[40][974],u_xpb_out[41][974],u_xpb_out[42][974],u_xpb_out[43][974],u_xpb_out[44][974],u_xpb_out[45][974],u_xpb_out[46][974],u_xpb_out[47][974],u_xpb_out[48][974],u_xpb_out[49][974],u_xpb_out[50][974],u_xpb_out[51][974],u_xpb_out[52][974],u_xpb_out[53][974],u_xpb_out[54][974],u_xpb_out[55][974],u_xpb_out[56][974],u_xpb_out[57][974],u_xpb_out[58][974],u_xpb_out[59][974],u_xpb_out[60][974],u_xpb_out[61][974],u_xpb_out[62][974],u_xpb_out[63][974],u_xpb_out[64][974],u_xpb_out[65][974],u_xpb_out[66][974],u_xpb_out[67][974],u_xpb_out[68][974],u_xpb_out[69][974],u_xpb_out[70][974],u_xpb_out[71][974],u_xpb_out[72][974],u_xpb_out[73][974],u_xpb_out[74][974],u_xpb_out[75][974],u_xpb_out[76][974],u_xpb_out[77][974],u_xpb_out[78][974],u_xpb_out[79][974],u_xpb_out[80][974],u_xpb_out[81][974],u_xpb_out[82][974],u_xpb_out[83][974],u_xpb_out[84][974],u_xpb_out[85][974],u_xpb_out[86][974],u_xpb_out[87][974],u_xpb_out[88][974],u_xpb_out[89][974],u_xpb_out[90][974],u_xpb_out[91][974],u_xpb_out[92][974],u_xpb_out[93][974],u_xpb_out[94][974],u_xpb_out[95][974],u_xpb_out[96][974],u_xpb_out[97][974],u_xpb_out[98][974],u_xpb_out[99][974],u_xpb_out[100][974],u_xpb_out[101][974],u_xpb_out[102][974],u_xpb_out[103][974],u_xpb_out[104][974],u_xpb_out[105][974]};

assign col_out_975 = {u_xpb_out[0][975],u_xpb_out[1][975],u_xpb_out[2][975],u_xpb_out[3][975],u_xpb_out[4][975],u_xpb_out[5][975],u_xpb_out[6][975],u_xpb_out[7][975],u_xpb_out[8][975],u_xpb_out[9][975],u_xpb_out[10][975],u_xpb_out[11][975],u_xpb_out[12][975],u_xpb_out[13][975],u_xpb_out[14][975],u_xpb_out[15][975],u_xpb_out[16][975],u_xpb_out[17][975],u_xpb_out[18][975],u_xpb_out[19][975],u_xpb_out[20][975],u_xpb_out[21][975],u_xpb_out[22][975],u_xpb_out[23][975],u_xpb_out[24][975],u_xpb_out[25][975],u_xpb_out[26][975],u_xpb_out[27][975],u_xpb_out[28][975],u_xpb_out[29][975],u_xpb_out[30][975],u_xpb_out[31][975],u_xpb_out[32][975],u_xpb_out[33][975],u_xpb_out[34][975],u_xpb_out[35][975],u_xpb_out[36][975],u_xpb_out[37][975],u_xpb_out[38][975],u_xpb_out[39][975],u_xpb_out[40][975],u_xpb_out[41][975],u_xpb_out[42][975],u_xpb_out[43][975],u_xpb_out[44][975],u_xpb_out[45][975],u_xpb_out[46][975],u_xpb_out[47][975],u_xpb_out[48][975],u_xpb_out[49][975],u_xpb_out[50][975],u_xpb_out[51][975],u_xpb_out[52][975],u_xpb_out[53][975],u_xpb_out[54][975],u_xpb_out[55][975],u_xpb_out[56][975],u_xpb_out[57][975],u_xpb_out[58][975],u_xpb_out[59][975],u_xpb_out[60][975],u_xpb_out[61][975],u_xpb_out[62][975],u_xpb_out[63][975],u_xpb_out[64][975],u_xpb_out[65][975],u_xpb_out[66][975],u_xpb_out[67][975],u_xpb_out[68][975],u_xpb_out[69][975],u_xpb_out[70][975],u_xpb_out[71][975],u_xpb_out[72][975],u_xpb_out[73][975],u_xpb_out[74][975],u_xpb_out[75][975],u_xpb_out[76][975],u_xpb_out[77][975],u_xpb_out[78][975],u_xpb_out[79][975],u_xpb_out[80][975],u_xpb_out[81][975],u_xpb_out[82][975],u_xpb_out[83][975],u_xpb_out[84][975],u_xpb_out[85][975],u_xpb_out[86][975],u_xpb_out[87][975],u_xpb_out[88][975],u_xpb_out[89][975],u_xpb_out[90][975],u_xpb_out[91][975],u_xpb_out[92][975],u_xpb_out[93][975],u_xpb_out[94][975],u_xpb_out[95][975],u_xpb_out[96][975],u_xpb_out[97][975],u_xpb_out[98][975],u_xpb_out[99][975],u_xpb_out[100][975],u_xpb_out[101][975],u_xpb_out[102][975],u_xpb_out[103][975],u_xpb_out[104][975],u_xpb_out[105][975]};

assign col_out_976 = {u_xpb_out[0][976],u_xpb_out[1][976],u_xpb_out[2][976],u_xpb_out[3][976],u_xpb_out[4][976],u_xpb_out[5][976],u_xpb_out[6][976],u_xpb_out[7][976],u_xpb_out[8][976],u_xpb_out[9][976],u_xpb_out[10][976],u_xpb_out[11][976],u_xpb_out[12][976],u_xpb_out[13][976],u_xpb_out[14][976],u_xpb_out[15][976],u_xpb_out[16][976],u_xpb_out[17][976],u_xpb_out[18][976],u_xpb_out[19][976],u_xpb_out[20][976],u_xpb_out[21][976],u_xpb_out[22][976],u_xpb_out[23][976],u_xpb_out[24][976],u_xpb_out[25][976],u_xpb_out[26][976],u_xpb_out[27][976],u_xpb_out[28][976],u_xpb_out[29][976],u_xpb_out[30][976],u_xpb_out[31][976],u_xpb_out[32][976],u_xpb_out[33][976],u_xpb_out[34][976],u_xpb_out[35][976],u_xpb_out[36][976],u_xpb_out[37][976],u_xpb_out[38][976],u_xpb_out[39][976],u_xpb_out[40][976],u_xpb_out[41][976],u_xpb_out[42][976],u_xpb_out[43][976],u_xpb_out[44][976],u_xpb_out[45][976],u_xpb_out[46][976],u_xpb_out[47][976],u_xpb_out[48][976],u_xpb_out[49][976],u_xpb_out[50][976],u_xpb_out[51][976],u_xpb_out[52][976],u_xpb_out[53][976],u_xpb_out[54][976],u_xpb_out[55][976],u_xpb_out[56][976],u_xpb_out[57][976],u_xpb_out[58][976],u_xpb_out[59][976],u_xpb_out[60][976],u_xpb_out[61][976],u_xpb_out[62][976],u_xpb_out[63][976],u_xpb_out[64][976],u_xpb_out[65][976],u_xpb_out[66][976],u_xpb_out[67][976],u_xpb_out[68][976],u_xpb_out[69][976],u_xpb_out[70][976],u_xpb_out[71][976],u_xpb_out[72][976],u_xpb_out[73][976],u_xpb_out[74][976],u_xpb_out[75][976],u_xpb_out[76][976],u_xpb_out[77][976],u_xpb_out[78][976],u_xpb_out[79][976],u_xpb_out[80][976],u_xpb_out[81][976],u_xpb_out[82][976],u_xpb_out[83][976],u_xpb_out[84][976],u_xpb_out[85][976],u_xpb_out[86][976],u_xpb_out[87][976],u_xpb_out[88][976],u_xpb_out[89][976],u_xpb_out[90][976],u_xpb_out[91][976],u_xpb_out[92][976],u_xpb_out[93][976],u_xpb_out[94][976],u_xpb_out[95][976],u_xpb_out[96][976],u_xpb_out[97][976],u_xpb_out[98][976],u_xpb_out[99][976],u_xpb_out[100][976],u_xpb_out[101][976],u_xpb_out[102][976],u_xpb_out[103][976],u_xpb_out[104][976],u_xpb_out[105][976]};

assign col_out_977 = {u_xpb_out[0][977],u_xpb_out[1][977],u_xpb_out[2][977],u_xpb_out[3][977],u_xpb_out[4][977],u_xpb_out[5][977],u_xpb_out[6][977],u_xpb_out[7][977],u_xpb_out[8][977],u_xpb_out[9][977],u_xpb_out[10][977],u_xpb_out[11][977],u_xpb_out[12][977],u_xpb_out[13][977],u_xpb_out[14][977],u_xpb_out[15][977],u_xpb_out[16][977],u_xpb_out[17][977],u_xpb_out[18][977],u_xpb_out[19][977],u_xpb_out[20][977],u_xpb_out[21][977],u_xpb_out[22][977],u_xpb_out[23][977],u_xpb_out[24][977],u_xpb_out[25][977],u_xpb_out[26][977],u_xpb_out[27][977],u_xpb_out[28][977],u_xpb_out[29][977],u_xpb_out[30][977],u_xpb_out[31][977],u_xpb_out[32][977],u_xpb_out[33][977],u_xpb_out[34][977],u_xpb_out[35][977],u_xpb_out[36][977],u_xpb_out[37][977],u_xpb_out[38][977],u_xpb_out[39][977],u_xpb_out[40][977],u_xpb_out[41][977],u_xpb_out[42][977],u_xpb_out[43][977],u_xpb_out[44][977],u_xpb_out[45][977],u_xpb_out[46][977],u_xpb_out[47][977],u_xpb_out[48][977],u_xpb_out[49][977],u_xpb_out[50][977],u_xpb_out[51][977],u_xpb_out[52][977],u_xpb_out[53][977],u_xpb_out[54][977],u_xpb_out[55][977],u_xpb_out[56][977],u_xpb_out[57][977],u_xpb_out[58][977],u_xpb_out[59][977],u_xpb_out[60][977],u_xpb_out[61][977],u_xpb_out[62][977],u_xpb_out[63][977],u_xpb_out[64][977],u_xpb_out[65][977],u_xpb_out[66][977],u_xpb_out[67][977],u_xpb_out[68][977],u_xpb_out[69][977],u_xpb_out[70][977],u_xpb_out[71][977],u_xpb_out[72][977],u_xpb_out[73][977],u_xpb_out[74][977],u_xpb_out[75][977],u_xpb_out[76][977],u_xpb_out[77][977],u_xpb_out[78][977],u_xpb_out[79][977],u_xpb_out[80][977],u_xpb_out[81][977],u_xpb_out[82][977],u_xpb_out[83][977],u_xpb_out[84][977],u_xpb_out[85][977],u_xpb_out[86][977],u_xpb_out[87][977],u_xpb_out[88][977],u_xpb_out[89][977],u_xpb_out[90][977],u_xpb_out[91][977],u_xpb_out[92][977],u_xpb_out[93][977],u_xpb_out[94][977],u_xpb_out[95][977],u_xpb_out[96][977],u_xpb_out[97][977],u_xpb_out[98][977],u_xpb_out[99][977],u_xpb_out[100][977],u_xpb_out[101][977],u_xpb_out[102][977],u_xpb_out[103][977],u_xpb_out[104][977],u_xpb_out[105][977]};

assign col_out_978 = {u_xpb_out[0][978],u_xpb_out[1][978],u_xpb_out[2][978],u_xpb_out[3][978],u_xpb_out[4][978],u_xpb_out[5][978],u_xpb_out[6][978],u_xpb_out[7][978],u_xpb_out[8][978],u_xpb_out[9][978],u_xpb_out[10][978],u_xpb_out[11][978],u_xpb_out[12][978],u_xpb_out[13][978],u_xpb_out[14][978],u_xpb_out[15][978],u_xpb_out[16][978],u_xpb_out[17][978],u_xpb_out[18][978],u_xpb_out[19][978],u_xpb_out[20][978],u_xpb_out[21][978],u_xpb_out[22][978],u_xpb_out[23][978],u_xpb_out[24][978],u_xpb_out[25][978],u_xpb_out[26][978],u_xpb_out[27][978],u_xpb_out[28][978],u_xpb_out[29][978],u_xpb_out[30][978],u_xpb_out[31][978],u_xpb_out[32][978],u_xpb_out[33][978],u_xpb_out[34][978],u_xpb_out[35][978],u_xpb_out[36][978],u_xpb_out[37][978],u_xpb_out[38][978],u_xpb_out[39][978],u_xpb_out[40][978],u_xpb_out[41][978],u_xpb_out[42][978],u_xpb_out[43][978],u_xpb_out[44][978],u_xpb_out[45][978],u_xpb_out[46][978],u_xpb_out[47][978],u_xpb_out[48][978],u_xpb_out[49][978],u_xpb_out[50][978],u_xpb_out[51][978],u_xpb_out[52][978],u_xpb_out[53][978],u_xpb_out[54][978],u_xpb_out[55][978],u_xpb_out[56][978],u_xpb_out[57][978],u_xpb_out[58][978],u_xpb_out[59][978],u_xpb_out[60][978],u_xpb_out[61][978],u_xpb_out[62][978],u_xpb_out[63][978],u_xpb_out[64][978],u_xpb_out[65][978],u_xpb_out[66][978],u_xpb_out[67][978],u_xpb_out[68][978],u_xpb_out[69][978],u_xpb_out[70][978],u_xpb_out[71][978],u_xpb_out[72][978],u_xpb_out[73][978],u_xpb_out[74][978],u_xpb_out[75][978],u_xpb_out[76][978],u_xpb_out[77][978],u_xpb_out[78][978],u_xpb_out[79][978],u_xpb_out[80][978],u_xpb_out[81][978],u_xpb_out[82][978],u_xpb_out[83][978],u_xpb_out[84][978],u_xpb_out[85][978],u_xpb_out[86][978],u_xpb_out[87][978],u_xpb_out[88][978],u_xpb_out[89][978],u_xpb_out[90][978],u_xpb_out[91][978],u_xpb_out[92][978],u_xpb_out[93][978],u_xpb_out[94][978],u_xpb_out[95][978],u_xpb_out[96][978],u_xpb_out[97][978],u_xpb_out[98][978],u_xpb_out[99][978],u_xpb_out[100][978],u_xpb_out[101][978],u_xpb_out[102][978],u_xpb_out[103][978],u_xpb_out[104][978],u_xpb_out[105][978]};

assign col_out_979 = {u_xpb_out[0][979],u_xpb_out[1][979],u_xpb_out[2][979],u_xpb_out[3][979],u_xpb_out[4][979],u_xpb_out[5][979],u_xpb_out[6][979],u_xpb_out[7][979],u_xpb_out[8][979],u_xpb_out[9][979],u_xpb_out[10][979],u_xpb_out[11][979],u_xpb_out[12][979],u_xpb_out[13][979],u_xpb_out[14][979],u_xpb_out[15][979],u_xpb_out[16][979],u_xpb_out[17][979],u_xpb_out[18][979],u_xpb_out[19][979],u_xpb_out[20][979],u_xpb_out[21][979],u_xpb_out[22][979],u_xpb_out[23][979],u_xpb_out[24][979],u_xpb_out[25][979],u_xpb_out[26][979],u_xpb_out[27][979],u_xpb_out[28][979],u_xpb_out[29][979],u_xpb_out[30][979],u_xpb_out[31][979],u_xpb_out[32][979],u_xpb_out[33][979],u_xpb_out[34][979],u_xpb_out[35][979],u_xpb_out[36][979],u_xpb_out[37][979],u_xpb_out[38][979],u_xpb_out[39][979],u_xpb_out[40][979],u_xpb_out[41][979],u_xpb_out[42][979],u_xpb_out[43][979],u_xpb_out[44][979],u_xpb_out[45][979],u_xpb_out[46][979],u_xpb_out[47][979],u_xpb_out[48][979],u_xpb_out[49][979],u_xpb_out[50][979],u_xpb_out[51][979],u_xpb_out[52][979],u_xpb_out[53][979],u_xpb_out[54][979],u_xpb_out[55][979],u_xpb_out[56][979],u_xpb_out[57][979],u_xpb_out[58][979],u_xpb_out[59][979],u_xpb_out[60][979],u_xpb_out[61][979],u_xpb_out[62][979],u_xpb_out[63][979],u_xpb_out[64][979],u_xpb_out[65][979],u_xpb_out[66][979],u_xpb_out[67][979],u_xpb_out[68][979],u_xpb_out[69][979],u_xpb_out[70][979],u_xpb_out[71][979],u_xpb_out[72][979],u_xpb_out[73][979],u_xpb_out[74][979],u_xpb_out[75][979],u_xpb_out[76][979],u_xpb_out[77][979],u_xpb_out[78][979],u_xpb_out[79][979],u_xpb_out[80][979],u_xpb_out[81][979],u_xpb_out[82][979],u_xpb_out[83][979],u_xpb_out[84][979],u_xpb_out[85][979],u_xpb_out[86][979],u_xpb_out[87][979],u_xpb_out[88][979],u_xpb_out[89][979],u_xpb_out[90][979],u_xpb_out[91][979],u_xpb_out[92][979],u_xpb_out[93][979],u_xpb_out[94][979],u_xpb_out[95][979],u_xpb_out[96][979],u_xpb_out[97][979],u_xpb_out[98][979],u_xpb_out[99][979],u_xpb_out[100][979],u_xpb_out[101][979],u_xpb_out[102][979],u_xpb_out[103][979],u_xpb_out[104][979],u_xpb_out[105][979]};

assign col_out_980 = {u_xpb_out[0][980],u_xpb_out[1][980],u_xpb_out[2][980],u_xpb_out[3][980],u_xpb_out[4][980],u_xpb_out[5][980],u_xpb_out[6][980],u_xpb_out[7][980],u_xpb_out[8][980],u_xpb_out[9][980],u_xpb_out[10][980],u_xpb_out[11][980],u_xpb_out[12][980],u_xpb_out[13][980],u_xpb_out[14][980],u_xpb_out[15][980],u_xpb_out[16][980],u_xpb_out[17][980],u_xpb_out[18][980],u_xpb_out[19][980],u_xpb_out[20][980],u_xpb_out[21][980],u_xpb_out[22][980],u_xpb_out[23][980],u_xpb_out[24][980],u_xpb_out[25][980],u_xpb_out[26][980],u_xpb_out[27][980],u_xpb_out[28][980],u_xpb_out[29][980],u_xpb_out[30][980],u_xpb_out[31][980],u_xpb_out[32][980],u_xpb_out[33][980],u_xpb_out[34][980],u_xpb_out[35][980],u_xpb_out[36][980],u_xpb_out[37][980],u_xpb_out[38][980],u_xpb_out[39][980],u_xpb_out[40][980],u_xpb_out[41][980],u_xpb_out[42][980],u_xpb_out[43][980],u_xpb_out[44][980],u_xpb_out[45][980],u_xpb_out[46][980],u_xpb_out[47][980],u_xpb_out[48][980],u_xpb_out[49][980],u_xpb_out[50][980],u_xpb_out[51][980],u_xpb_out[52][980],u_xpb_out[53][980],u_xpb_out[54][980],u_xpb_out[55][980],u_xpb_out[56][980],u_xpb_out[57][980],u_xpb_out[58][980],u_xpb_out[59][980],u_xpb_out[60][980],u_xpb_out[61][980],u_xpb_out[62][980],u_xpb_out[63][980],u_xpb_out[64][980],u_xpb_out[65][980],u_xpb_out[66][980],u_xpb_out[67][980],u_xpb_out[68][980],u_xpb_out[69][980],u_xpb_out[70][980],u_xpb_out[71][980],u_xpb_out[72][980],u_xpb_out[73][980],u_xpb_out[74][980],u_xpb_out[75][980],u_xpb_out[76][980],u_xpb_out[77][980],u_xpb_out[78][980],u_xpb_out[79][980],u_xpb_out[80][980],u_xpb_out[81][980],u_xpb_out[82][980],u_xpb_out[83][980],u_xpb_out[84][980],u_xpb_out[85][980],u_xpb_out[86][980],u_xpb_out[87][980],u_xpb_out[88][980],u_xpb_out[89][980],u_xpb_out[90][980],u_xpb_out[91][980],u_xpb_out[92][980],u_xpb_out[93][980],u_xpb_out[94][980],u_xpb_out[95][980],u_xpb_out[96][980],u_xpb_out[97][980],u_xpb_out[98][980],u_xpb_out[99][980],u_xpb_out[100][980],u_xpb_out[101][980],u_xpb_out[102][980],u_xpb_out[103][980],u_xpb_out[104][980],u_xpb_out[105][980]};

assign col_out_981 = {u_xpb_out[0][981],u_xpb_out[1][981],u_xpb_out[2][981],u_xpb_out[3][981],u_xpb_out[4][981],u_xpb_out[5][981],u_xpb_out[6][981],u_xpb_out[7][981],u_xpb_out[8][981],u_xpb_out[9][981],u_xpb_out[10][981],u_xpb_out[11][981],u_xpb_out[12][981],u_xpb_out[13][981],u_xpb_out[14][981],u_xpb_out[15][981],u_xpb_out[16][981],u_xpb_out[17][981],u_xpb_out[18][981],u_xpb_out[19][981],u_xpb_out[20][981],u_xpb_out[21][981],u_xpb_out[22][981],u_xpb_out[23][981],u_xpb_out[24][981],u_xpb_out[25][981],u_xpb_out[26][981],u_xpb_out[27][981],u_xpb_out[28][981],u_xpb_out[29][981],u_xpb_out[30][981],u_xpb_out[31][981],u_xpb_out[32][981],u_xpb_out[33][981],u_xpb_out[34][981],u_xpb_out[35][981],u_xpb_out[36][981],u_xpb_out[37][981],u_xpb_out[38][981],u_xpb_out[39][981],u_xpb_out[40][981],u_xpb_out[41][981],u_xpb_out[42][981],u_xpb_out[43][981],u_xpb_out[44][981],u_xpb_out[45][981],u_xpb_out[46][981],u_xpb_out[47][981],u_xpb_out[48][981],u_xpb_out[49][981],u_xpb_out[50][981],u_xpb_out[51][981],u_xpb_out[52][981],u_xpb_out[53][981],u_xpb_out[54][981],u_xpb_out[55][981],u_xpb_out[56][981],u_xpb_out[57][981],u_xpb_out[58][981],u_xpb_out[59][981],u_xpb_out[60][981],u_xpb_out[61][981],u_xpb_out[62][981],u_xpb_out[63][981],u_xpb_out[64][981],u_xpb_out[65][981],u_xpb_out[66][981],u_xpb_out[67][981],u_xpb_out[68][981],u_xpb_out[69][981],u_xpb_out[70][981],u_xpb_out[71][981],u_xpb_out[72][981],u_xpb_out[73][981],u_xpb_out[74][981],u_xpb_out[75][981],u_xpb_out[76][981],u_xpb_out[77][981],u_xpb_out[78][981],u_xpb_out[79][981],u_xpb_out[80][981],u_xpb_out[81][981],u_xpb_out[82][981],u_xpb_out[83][981],u_xpb_out[84][981],u_xpb_out[85][981],u_xpb_out[86][981],u_xpb_out[87][981],u_xpb_out[88][981],u_xpb_out[89][981],u_xpb_out[90][981],u_xpb_out[91][981],u_xpb_out[92][981],u_xpb_out[93][981],u_xpb_out[94][981],u_xpb_out[95][981],u_xpb_out[96][981],u_xpb_out[97][981],u_xpb_out[98][981],u_xpb_out[99][981],u_xpb_out[100][981],u_xpb_out[101][981],u_xpb_out[102][981],u_xpb_out[103][981],u_xpb_out[104][981],u_xpb_out[105][981]};

assign col_out_982 = {u_xpb_out[0][982],u_xpb_out[1][982],u_xpb_out[2][982],u_xpb_out[3][982],u_xpb_out[4][982],u_xpb_out[5][982],u_xpb_out[6][982],u_xpb_out[7][982],u_xpb_out[8][982],u_xpb_out[9][982],u_xpb_out[10][982],u_xpb_out[11][982],u_xpb_out[12][982],u_xpb_out[13][982],u_xpb_out[14][982],u_xpb_out[15][982],u_xpb_out[16][982],u_xpb_out[17][982],u_xpb_out[18][982],u_xpb_out[19][982],u_xpb_out[20][982],u_xpb_out[21][982],u_xpb_out[22][982],u_xpb_out[23][982],u_xpb_out[24][982],u_xpb_out[25][982],u_xpb_out[26][982],u_xpb_out[27][982],u_xpb_out[28][982],u_xpb_out[29][982],u_xpb_out[30][982],u_xpb_out[31][982],u_xpb_out[32][982],u_xpb_out[33][982],u_xpb_out[34][982],u_xpb_out[35][982],u_xpb_out[36][982],u_xpb_out[37][982],u_xpb_out[38][982],u_xpb_out[39][982],u_xpb_out[40][982],u_xpb_out[41][982],u_xpb_out[42][982],u_xpb_out[43][982],u_xpb_out[44][982],u_xpb_out[45][982],u_xpb_out[46][982],u_xpb_out[47][982],u_xpb_out[48][982],u_xpb_out[49][982],u_xpb_out[50][982],u_xpb_out[51][982],u_xpb_out[52][982],u_xpb_out[53][982],u_xpb_out[54][982],u_xpb_out[55][982],u_xpb_out[56][982],u_xpb_out[57][982],u_xpb_out[58][982],u_xpb_out[59][982],u_xpb_out[60][982],u_xpb_out[61][982],u_xpb_out[62][982],u_xpb_out[63][982],u_xpb_out[64][982],u_xpb_out[65][982],u_xpb_out[66][982],u_xpb_out[67][982],u_xpb_out[68][982],u_xpb_out[69][982],u_xpb_out[70][982],u_xpb_out[71][982],u_xpb_out[72][982],u_xpb_out[73][982],u_xpb_out[74][982],u_xpb_out[75][982],u_xpb_out[76][982],u_xpb_out[77][982],u_xpb_out[78][982],u_xpb_out[79][982],u_xpb_out[80][982],u_xpb_out[81][982],u_xpb_out[82][982],u_xpb_out[83][982],u_xpb_out[84][982],u_xpb_out[85][982],u_xpb_out[86][982],u_xpb_out[87][982],u_xpb_out[88][982],u_xpb_out[89][982],u_xpb_out[90][982],u_xpb_out[91][982],u_xpb_out[92][982],u_xpb_out[93][982],u_xpb_out[94][982],u_xpb_out[95][982],u_xpb_out[96][982],u_xpb_out[97][982],u_xpb_out[98][982],u_xpb_out[99][982],u_xpb_out[100][982],u_xpb_out[101][982],u_xpb_out[102][982],u_xpb_out[103][982],u_xpb_out[104][982],u_xpb_out[105][982]};

assign col_out_983 = {u_xpb_out[0][983],u_xpb_out[1][983],u_xpb_out[2][983],u_xpb_out[3][983],u_xpb_out[4][983],u_xpb_out[5][983],u_xpb_out[6][983],u_xpb_out[7][983],u_xpb_out[8][983],u_xpb_out[9][983],u_xpb_out[10][983],u_xpb_out[11][983],u_xpb_out[12][983],u_xpb_out[13][983],u_xpb_out[14][983],u_xpb_out[15][983],u_xpb_out[16][983],u_xpb_out[17][983],u_xpb_out[18][983],u_xpb_out[19][983],u_xpb_out[20][983],u_xpb_out[21][983],u_xpb_out[22][983],u_xpb_out[23][983],u_xpb_out[24][983],u_xpb_out[25][983],u_xpb_out[26][983],u_xpb_out[27][983],u_xpb_out[28][983],u_xpb_out[29][983],u_xpb_out[30][983],u_xpb_out[31][983],u_xpb_out[32][983],u_xpb_out[33][983],u_xpb_out[34][983],u_xpb_out[35][983],u_xpb_out[36][983],u_xpb_out[37][983],u_xpb_out[38][983],u_xpb_out[39][983],u_xpb_out[40][983],u_xpb_out[41][983],u_xpb_out[42][983],u_xpb_out[43][983],u_xpb_out[44][983],u_xpb_out[45][983],u_xpb_out[46][983],u_xpb_out[47][983],u_xpb_out[48][983],u_xpb_out[49][983],u_xpb_out[50][983],u_xpb_out[51][983],u_xpb_out[52][983],u_xpb_out[53][983],u_xpb_out[54][983],u_xpb_out[55][983],u_xpb_out[56][983],u_xpb_out[57][983],u_xpb_out[58][983],u_xpb_out[59][983],u_xpb_out[60][983],u_xpb_out[61][983],u_xpb_out[62][983],u_xpb_out[63][983],u_xpb_out[64][983],u_xpb_out[65][983],u_xpb_out[66][983],u_xpb_out[67][983],u_xpb_out[68][983],u_xpb_out[69][983],u_xpb_out[70][983],u_xpb_out[71][983],u_xpb_out[72][983],u_xpb_out[73][983],u_xpb_out[74][983],u_xpb_out[75][983],u_xpb_out[76][983],u_xpb_out[77][983],u_xpb_out[78][983],u_xpb_out[79][983],u_xpb_out[80][983],u_xpb_out[81][983],u_xpb_out[82][983],u_xpb_out[83][983],u_xpb_out[84][983],u_xpb_out[85][983],u_xpb_out[86][983],u_xpb_out[87][983],u_xpb_out[88][983],u_xpb_out[89][983],u_xpb_out[90][983],u_xpb_out[91][983],u_xpb_out[92][983],u_xpb_out[93][983],u_xpb_out[94][983],u_xpb_out[95][983],u_xpb_out[96][983],u_xpb_out[97][983],u_xpb_out[98][983],u_xpb_out[99][983],u_xpb_out[100][983],u_xpb_out[101][983],u_xpb_out[102][983],u_xpb_out[103][983],u_xpb_out[104][983],u_xpb_out[105][983]};

assign col_out_984 = {u_xpb_out[0][984],u_xpb_out[1][984],u_xpb_out[2][984],u_xpb_out[3][984],u_xpb_out[4][984],u_xpb_out[5][984],u_xpb_out[6][984],u_xpb_out[7][984],u_xpb_out[8][984],u_xpb_out[9][984],u_xpb_out[10][984],u_xpb_out[11][984],u_xpb_out[12][984],u_xpb_out[13][984],u_xpb_out[14][984],u_xpb_out[15][984],u_xpb_out[16][984],u_xpb_out[17][984],u_xpb_out[18][984],u_xpb_out[19][984],u_xpb_out[20][984],u_xpb_out[21][984],u_xpb_out[22][984],u_xpb_out[23][984],u_xpb_out[24][984],u_xpb_out[25][984],u_xpb_out[26][984],u_xpb_out[27][984],u_xpb_out[28][984],u_xpb_out[29][984],u_xpb_out[30][984],u_xpb_out[31][984],u_xpb_out[32][984],u_xpb_out[33][984],u_xpb_out[34][984],u_xpb_out[35][984],u_xpb_out[36][984],u_xpb_out[37][984],u_xpb_out[38][984],u_xpb_out[39][984],u_xpb_out[40][984],u_xpb_out[41][984],u_xpb_out[42][984],u_xpb_out[43][984],u_xpb_out[44][984],u_xpb_out[45][984],u_xpb_out[46][984],u_xpb_out[47][984],u_xpb_out[48][984],u_xpb_out[49][984],u_xpb_out[50][984],u_xpb_out[51][984],u_xpb_out[52][984],u_xpb_out[53][984],u_xpb_out[54][984],u_xpb_out[55][984],u_xpb_out[56][984],u_xpb_out[57][984],u_xpb_out[58][984],u_xpb_out[59][984],u_xpb_out[60][984],u_xpb_out[61][984],u_xpb_out[62][984],u_xpb_out[63][984],u_xpb_out[64][984],u_xpb_out[65][984],u_xpb_out[66][984],u_xpb_out[67][984],u_xpb_out[68][984],u_xpb_out[69][984],u_xpb_out[70][984],u_xpb_out[71][984],u_xpb_out[72][984],u_xpb_out[73][984],u_xpb_out[74][984],u_xpb_out[75][984],u_xpb_out[76][984],u_xpb_out[77][984],u_xpb_out[78][984],u_xpb_out[79][984],u_xpb_out[80][984],u_xpb_out[81][984],u_xpb_out[82][984],u_xpb_out[83][984],u_xpb_out[84][984],u_xpb_out[85][984],u_xpb_out[86][984],u_xpb_out[87][984],u_xpb_out[88][984],u_xpb_out[89][984],u_xpb_out[90][984],u_xpb_out[91][984],u_xpb_out[92][984],u_xpb_out[93][984],u_xpb_out[94][984],u_xpb_out[95][984],u_xpb_out[96][984],u_xpb_out[97][984],u_xpb_out[98][984],u_xpb_out[99][984],u_xpb_out[100][984],u_xpb_out[101][984],u_xpb_out[102][984],u_xpb_out[103][984],u_xpb_out[104][984],u_xpb_out[105][984]};

assign col_out_985 = {u_xpb_out[0][985],u_xpb_out[1][985],u_xpb_out[2][985],u_xpb_out[3][985],u_xpb_out[4][985],u_xpb_out[5][985],u_xpb_out[6][985],u_xpb_out[7][985],u_xpb_out[8][985],u_xpb_out[9][985],u_xpb_out[10][985],u_xpb_out[11][985],u_xpb_out[12][985],u_xpb_out[13][985],u_xpb_out[14][985],u_xpb_out[15][985],u_xpb_out[16][985],u_xpb_out[17][985],u_xpb_out[18][985],u_xpb_out[19][985],u_xpb_out[20][985],u_xpb_out[21][985],u_xpb_out[22][985],u_xpb_out[23][985],u_xpb_out[24][985],u_xpb_out[25][985],u_xpb_out[26][985],u_xpb_out[27][985],u_xpb_out[28][985],u_xpb_out[29][985],u_xpb_out[30][985],u_xpb_out[31][985],u_xpb_out[32][985],u_xpb_out[33][985],u_xpb_out[34][985],u_xpb_out[35][985],u_xpb_out[36][985],u_xpb_out[37][985],u_xpb_out[38][985],u_xpb_out[39][985],u_xpb_out[40][985],u_xpb_out[41][985],u_xpb_out[42][985],u_xpb_out[43][985],u_xpb_out[44][985],u_xpb_out[45][985],u_xpb_out[46][985],u_xpb_out[47][985],u_xpb_out[48][985],u_xpb_out[49][985],u_xpb_out[50][985],u_xpb_out[51][985],u_xpb_out[52][985],u_xpb_out[53][985],u_xpb_out[54][985],u_xpb_out[55][985],u_xpb_out[56][985],u_xpb_out[57][985],u_xpb_out[58][985],u_xpb_out[59][985],u_xpb_out[60][985],u_xpb_out[61][985],u_xpb_out[62][985],u_xpb_out[63][985],u_xpb_out[64][985],u_xpb_out[65][985],u_xpb_out[66][985],u_xpb_out[67][985],u_xpb_out[68][985],u_xpb_out[69][985],u_xpb_out[70][985],u_xpb_out[71][985],u_xpb_out[72][985],u_xpb_out[73][985],u_xpb_out[74][985],u_xpb_out[75][985],u_xpb_out[76][985],u_xpb_out[77][985],u_xpb_out[78][985],u_xpb_out[79][985],u_xpb_out[80][985],u_xpb_out[81][985],u_xpb_out[82][985],u_xpb_out[83][985],u_xpb_out[84][985],u_xpb_out[85][985],u_xpb_out[86][985],u_xpb_out[87][985],u_xpb_out[88][985],u_xpb_out[89][985],u_xpb_out[90][985],u_xpb_out[91][985],u_xpb_out[92][985],u_xpb_out[93][985],u_xpb_out[94][985],u_xpb_out[95][985],u_xpb_out[96][985],u_xpb_out[97][985],u_xpb_out[98][985],u_xpb_out[99][985],u_xpb_out[100][985],u_xpb_out[101][985],u_xpb_out[102][985],u_xpb_out[103][985],u_xpb_out[104][985],u_xpb_out[105][985]};

assign col_out_986 = {u_xpb_out[0][986],u_xpb_out[1][986],u_xpb_out[2][986],u_xpb_out[3][986],u_xpb_out[4][986],u_xpb_out[5][986],u_xpb_out[6][986],u_xpb_out[7][986],u_xpb_out[8][986],u_xpb_out[9][986],u_xpb_out[10][986],u_xpb_out[11][986],u_xpb_out[12][986],u_xpb_out[13][986],u_xpb_out[14][986],u_xpb_out[15][986],u_xpb_out[16][986],u_xpb_out[17][986],u_xpb_out[18][986],u_xpb_out[19][986],u_xpb_out[20][986],u_xpb_out[21][986],u_xpb_out[22][986],u_xpb_out[23][986],u_xpb_out[24][986],u_xpb_out[25][986],u_xpb_out[26][986],u_xpb_out[27][986],u_xpb_out[28][986],u_xpb_out[29][986],u_xpb_out[30][986],u_xpb_out[31][986],u_xpb_out[32][986],u_xpb_out[33][986],u_xpb_out[34][986],u_xpb_out[35][986],u_xpb_out[36][986],u_xpb_out[37][986],u_xpb_out[38][986],u_xpb_out[39][986],u_xpb_out[40][986],u_xpb_out[41][986],u_xpb_out[42][986],u_xpb_out[43][986],u_xpb_out[44][986],u_xpb_out[45][986],u_xpb_out[46][986],u_xpb_out[47][986],u_xpb_out[48][986],u_xpb_out[49][986],u_xpb_out[50][986],u_xpb_out[51][986],u_xpb_out[52][986],u_xpb_out[53][986],u_xpb_out[54][986],u_xpb_out[55][986],u_xpb_out[56][986],u_xpb_out[57][986],u_xpb_out[58][986],u_xpb_out[59][986],u_xpb_out[60][986],u_xpb_out[61][986],u_xpb_out[62][986],u_xpb_out[63][986],u_xpb_out[64][986],u_xpb_out[65][986],u_xpb_out[66][986],u_xpb_out[67][986],u_xpb_out[68][986],u_xpb_out[69][986],u_xpb_out[70][986],u_xpb_out[71][986],u_xpb_out[72][986],u_xpb_out[73][986],u_xpb_out[74][986],u_xpb_out[75][986],u_xpb_out[76][986],u_xpb_out[77][986],u_xpb_out[78][986],u_xpb_out[79][986],u_xpb_out[80][986],u_xpb_out[81][986],u_xpb_out[82][986],u_xpb_out[83][986],u_xpb_out[84][986],u_xpb_out[85][986],u_xpb_out[86][986],u_xpb_out[87][986],u_xpb_out[88][986],u_xpb_out[89][986],u_xpb_out[90][986],u_xpb_out[91][986],u_xpb_out[92][986],u_xpb_out[93][986],u_xpb_out[94][986],u_xpb_out[95][986],u_xpb_out[96][986],u_xpb_out[97][986],u_xpb_out[98][986],u_xpb_out[99][986],u_xpb_out[100][986],u_xpb_out[101][986],u_xpb_out[102][986],u_xpb_out[103][986],u_xpb_out[104][986],u_xpb_out[105][986]};

assign col_out_987 = {u_xpb_out[0][987],u_xpb_out[1][987],u_xpb_out[2][987],u_xpb_out[3][987],u_xpb_out[4][987],u_xpb_out[5][987],u_xpb_out[6][987],u_xpb_out[7][987],u_xpb_out[8][987],u_xpb_out[9][987],u_xpb_out[10][987],u_xpb_out[11][987],u_xpb_out[12][987],u_xpb_out[13][987],u_xpb_out[14][987],u_xpb_out[15][987],u_xpb_out[16][987],u_xpb_out[17][987],u_xpb_out[18][987],u_xpb_out[19][987],u_xpb_out[20][987],u_xpb_out[21][987],u_xpb_out[22][987],u_xpb_out[23][987],u_xpb_out[24][987],u_xpb_out[25][987],u_xpb_out[26][987],u_xpb_out[27][987],u_xpb_out[28][987],u_xpb_out[29][987],u_xpb_out[30][987],u_xpb_out[31][987],u_xpb_out[32][987],u_xpb_out[33][987],u_xpb_out[34][987],u_xpb_out[35][987],u_xpb_out[36][987],u_xpb_out[37][987],u_xpb_out[38][987],u_xpb_out[39][987],u_xpb_out[40][987],u_xpb_out[41][987],u_xpb_out[42][987],u_xpb_out[43][987],u_xpb_out[44][987],u_xpb_out[45][987],u_xpb_out[46][987],u_xpb_out[47][987],u_xpb_out[48][987],u_xpb_out[49][987],u_xpb_out[50][987],u_xpb_out[51][987],u_xpb_out[52][987],u_xpb_out[53][987],u_xpb_out[54][987],u_xpb_out[55][987],u_xpb_out[56][987],u_xpb_out[57][987],u_xpb_out[58][987],u_xpb_out[59][987],u_xpb_out[60][987],u_xpb_out[61][987],u_xpb_out[62][987],u_xpb_out[63][987],u_xpb_out[64][987],u_xpb_out[65][987],u_xpb_out[66][987],u_xpb_out[67][987],u_xpb_out[68][987],u_xpb_out[69][987],u_xpb_out[70][987],u_xpb_out[71][987],u_xpb_out[72][987],u_xpb_out[73][987],u_xpb_out[74][987],u_xpb_out[75][987],u_xpb_out[76][987],u_xpb_out[77][987],u_xpb_out[78][987],u_xpb_out[79][987],u_xpb_out[80][987],u_xpb_out[81][987],u_xpb_out[82][987],u_xpb_out[83][987],u_xpb_out[84][987],u_xpb_out[85][987],u_xpb_out[86][987],u_xpb_out[87][987],u_xpb_out[88][987],u_xpb_out[89][987],u_xpb_out[90][987],u_xpb_out[91][987],u_xpb_out[92][987],u_xpb_out[93][987],u_xpb_out[94][987],u_xpb_out[95][987],u_xpb_out[96][987],u_xpb_out[97][987],u_xpb_out[98][987],u_xpb_out[99][987],u_xpb_out[100][987],u_xpb_out[101][987],u_xpb_out[102][987],u_xpb_out[103][987],u_xpb_out[104][987],u_xpb_out[105][987]};

assign col_out_988 = {u_xpb_out[0][988],u_xpb_out[1][988],u_xpb_out[2][988],u_xpb_out[3][988],u_xpb_out[4][988],u_xpb_out[5][988],u_xpb_out[6][988],u_xpb_out[7][988],u_xpb_out[8][988],u_xpb_out[9][988],u_xpb_out[10][988],u_xpb_out[11][988],u_xpb_out[12][988],u_xpb_out[13][988],u_xpb_out[14][988],u_xpb_out[15][988],u_xpb_out[16][988],u_xpb_out[17][988],u_xpb_out[18][988],u_xpb_out[19][988],u_xpb_out[20][988],u_xpb_out[21][988],u_xpb_out[22][988],u_xpb_out[23][988],u_xpb_out[24][988],u_xpb_out[25][988],u_xpb_out[26][988],u_xpb_out[27][988],u_xpb_out[28][988],u_xpb_out[29][988],u_xpb_out[30][988],u_xpb_out[31][988],u_xpb_out[32][988],u_xpb_out[33][988],u_xpb_out[34][988],u_xpb_out[35][988],u_xpb_out[36][988],u_xpb_out[37][988],u_xpb_out[38][988],u_xpb_out[39][988],u_xpb_out[40][988],u_xpb_out[41][988],u_xpb_out[42][988],u_xpb_out[43][988],u_xpb_out[44][988],u_xpb_out[45][988],u_xpb_out[46][988],u_xpb_out[47][988],u_xpb_out[48][988],u_xpb_out[49][988],u_xpb_out[50][988],u_xpb_out[51][988],u_xpb_out[52][988],u_xpb_out[53][988],u_xpb_out[54][988],u_xpb_out[55][988],u_xpb_out[56][988],u_xpb_out[57][988],u_xpb_out[58][988],u_xpb_out[59][988],u_xpb_out[60][988],u_xpb_out[61][988],u_xpb_out[62][988],u_xpb_out[63][988],u_xpb_out[64][988],u_xpb_out[65][988],u_xpb_out[66][988],u_xpb_out[67][988],u_xpb_out[68][988],u_xpb_out[69][988],u_xpb_out[70][988],u_xpb_out[71][988],u_xpb_out[72][988],u_xpb_out[73][988],u_xpb_out[74][988],u_xpb_out[75][988],u_xpb_out[76][988],u_xpb_out[77][988],u_xpb_out[78][988],u_xpb_out[79][988],u_xpb_out[80][988],u_xpb_out[81][988],u_xpb_out[82][988],u_xpb_out[83][988],u_xpb_out[84][988],u_xpb_out[85][988],u_xpb_out[86][988],u_xpb_out[87][988],u_xpb_out[88][988],u_xpb_out[89][988],u_xpb_out[90][988],u_xpb_out[91][988],u_xpb_out[92][988],u_xpb_out[93][988],u_xpb_out[94][988],u_xpb_out[95][988],u_xpb_out[96][988],u_xpb_out[97][988],u_xpb_out[98][988],u_xpb_out[99][988],u_xpb_out[100][988],u_xpb_out[101][988],u_xpb_out[102][988],u_xpb_out[103][988],u_xpb_out[104][988],u_xpb_out[105][988]};

assign col_out_989 = {u_xpb_out[0][989],u_xpb_out[1][989],u_xpb_out[2][989],u_xpb_out[3][989],u_xpb_out[4][989],u_xpb_out[5][989],u_xpb_out[6][989],u_xpb_out[7][989],u_xpb_out[8][989],u_xpb_out[9][989],u_xpb_out[10][989],u_xpb_out[11][989],u_xpb_out[12][989],u_xpb_out[13][989],u_xpb_out[14][989],u_xpb_out[15][989],u_xpb_out[16][989],u_xpb_out[17][989],u_xpb_out[18][989],u_xpb_out[19][989],u_xpb_out[20][989],u_xpb_out[21][989],u_xpb_out[22][989],u_xpb_out[23][989],u_xpb_out[24][989],u_xpb_out[25][989],u_xpb_out[26][989],u_xpb_out[27][989],u_xpb_out[28][989],u_xpb_out[29][989],u_xpb_out[30][989],u_xpb_out[31][989],u_xpb_out[32][989],u_xpb_out[33][989],u_xpb_out[34][989],u_xpb_out[35][989],u_xpb_out[36][989],u_xpb_out[37][989],u_xpb_out[38][989],u_xpb_out[39][989],u_xpb_out[40][989],u_xpb_out[41][989],u_xpb_out[42][989],u_xpb_out[43][989],u_xpb_out[44][989],u_xpb_out[45][989],u_xpb_out[46][989],u_xpb_out[47][989],u_xpb_out[48][989],u_xpb_out[49][989],u_xpb_out[50][989],u_xpb_out[51][989],u_xpb_out[52][989],u_xpb_out[53][989],u_xpb_out[54][989],u_xpb_out[55][989],u_xpb_out[56][989],u_xpb_out[57][989],u_xpb_out[58][989],u_xpb_out[59][989],u_xpb_out[60][989],u_xpb_out[61][989],u_xpb_out[62][989],u_xpb_out[63][989],u_xpb_out[64][989],u_xpb_out[65][989],u_xpb_out[66][989],u_xpb_out[67][989],u_xpb_out[68][989],u_xpb_out[69][989],u_xpb_out[70][989],u_xpb_out[71][989],u_xpb_out[72][989],u_xpb_out[73][989],u_xpb_out[74][989],u_xpb_out[75][989],u_xpb_out[76][989],u_xpb_out[77][989],u_xpb_out[78][989],u_xpb_out[79][989],u_xpb_out[80][989],u_xpb_out[81][989],u_xpb_out[82][989],u_xpb_out[83][989],u_xpb_out[84][989],u_xpb_out[85][989],u_xpb_out[86][989],u_xpb_out[87][989],u_xpb_out[88][989],u_xpb_out[89][989],u_xpb_out[90][989],u_xpb_out[91][989],u_xpb_out[92][989],u_xpb_out[93][989],u_xpb_out[94][989],u_xpb_out[95][989],u_xpb_out[96][989],u_xpb_out[97][989],u_xpb_out[98][989],u_xpb_out[99][989],u_xpb_out[100][989],u_xpb_out[101][989],u_xpb_out[102][989],u_xpb_out[103][989],u_xpb_out[104][989],u_xpb_out[105][989]};

assign col_out_990 = {u_xpb_out[0][990],u_xpb_out[1][990],u_xpb_out[2][990],u_xpb_out[3][990],u_xpb_out[4][990],u_xpb_out[5][990],u_xpb_out[6][990],u_xpb_out[7][990],u_xpb_out[8][990],u_xpb_out[9][990],u_xpb_out[10][990],u_xpb_out[11][990],u_xpb_out[12][990],u_xpb_out[13][990],u_xpb_out[14][990],u_xpb_out[15][990],u_xpb_out[16][990],u_xpb_out[17][990],u_xpb_out[18][990],u_xpb_out[19][990],u_xpb_out[20][990],u_xpb_out[21][990],u_xpb_out[22][990],u_xpb_out[23][990],u_xpb_out[24][990],u_xpb_out[25][990],u_xpb_out[26][990],u_xpb_out[27][990],u_xpb_out[28][990],u_xpb_out[29][990],u_xpb_out[30][990],u_xpb_out[31][990],u_xpb_out[32][990],u_xpb_out[33][990],u_xpb_out[34][990],u_xpb_out[35][990],u_xpb_out[36][990],u_xpb_out[37][990],u_xpb_out[38][990],u_xpb_out[39][990],u_xpb_out[40][990],u_xpb_out[41][990],u_xpb_out[42][990],u_xpb_out[43][990],u_xpb_out[44][990],u_xpb_out[45][990],u_xpb_out[46][990],u_xpb_out[47][990],u_xpb_out[48][990],u_xpb_out[49][990],u_xpb_out[50][990],u_xpb_out[51][990],u_xpb_out[52][990],u_xpb_out[53][990],u_xpb_out[54][990],u_xpb_out[55][990],u_xpb_out[56][990],u_xpb_out[57][990],u_xpb_out[58][990],u_xpb_out[59][990],u_xpb_out[60][990],u_xpb_out[61][990],u_xpb_out[62][990],u_xpb_out[63][990],u_xpb_out[64][990],u_xpb_out[65][990],u_xpb_out[66][990],u_xpb_out[67][990],u_xpb_out[68][990],u_xpb_out[69][990],u_xpb_out[70][990],u_xpb_out[71][990],u_xpb_out[72][990],u_xpb_out[73][990],u_xpb_out[74][990],u_xpb_out[75][990],u_xpb_out[76][990],u_xpb_out[77][990],u_xpb_out[78][990],u_xpb_out[79][990],u_xpb_out[80][990],u_xpb_out[81][990],u_xpb_out[82][990],u_xpb_out[83][990],u_xpb_out[84][990],u_xpb_out[85][990],u_xpb_out[86][990],u_xpb_out[87][990],u_xpb_out[88][990],u_xpb_out[89][990],u_xpb_out[90][990],u_xpb_out[91][990],u_xpb_out[92][990],u_xpb_out[93][990],u_xpb_out[94][990],u_xpb_out[95][990],u_xpb_out[96][990],u_xpb_out[97][990],u_xpb_out[98][990],u_xpb_out[99][990],u_xpb_out[100][990],u_xpb_out[101][990],u_xpb_out[102][990],u_xpb_out[103][990],u_xpb_out[104][990],u_xpb_out[105][990]};

assign col_out_991 = {u_xpb_out[0][991],u_xpb_out[1][991],u_xpb_out[2][991],u_xpb_out[3][991],u_xpb_out[4][991],u_xpb_out[5][991],u_xpb_out[6][991],u_xpb_out[7][991],u_xpb_out[8][991],u_xpb_out[9][991],u_xpb_out[10][991],u_xpb_out[11][991],u_xpb_out[12][991],u_xpb_out[13][991],u_xpb_out[14][991],u_xpb_out[15][991],u_xpb_out[16][991],u_xpb_out[17][991],u_xpb_out[18][991],u_xpb_out[19][991],u_xpb_out[20][991],u_xpb_out[21][991],u_xpb_out[22][991],u_xpb_out[23][991],u_xpb_out[24][991],u_xpb_out[25][991],u_xpb_out[26][991],u_xpb_out[27][991],u_xpb_out[28][991],u_xpb_out[29][991],u_xpb_out[30][991],u_xpb_out[31][991],u_xpb_out[32][991],u_xpb_out[33][991],u_xpb_out[34][991],u_xpb_out[35][991],u_xpb_out[36][991],u_xpb_out[37][991],u_xpb_out[38][991],u_xpb_out[39][991],u_xpb_out[40][991],u_xpb_out[41][991],u_xpb_out[42][991],u_xpb_out[43][991],u_xpb_out[44][991],u_xpb_out[45][991],u_xpb_out[46][991],u_xpb_out[47][991],u_xpb_out[48][991],u_xpb_out[49][991],u_xpb_out[50][991],u_xpb_out[51][991],u_xpb_out[52][991],u_xpb_out[53][991],u_xpb_out[54][991],u_xpb_out[55][991],u_xpb_out[56][991],u_xpb_out[57][991],u_xpb_out[58][991],u_xpb_out[59][991],u_xpb_out[60][991],u_xpb_out[61][991],u_xpb_out[62][991],u_xpb_out[63][991],u_xpb_out[64][991],u_xpb_out[65][991],u_xpb_out[66][991],u_xpb_out[67][991],u_xpb_out[68][991],u_xpb_out[69][991],u_xpb_out[70][991],u_xpb_out[71][991],u_xpb_out[72][991],u_xpb_out[73][991],u_xpb_out[74][991],u_xpb_out[75][991],u_xpb_out[76][991],u_xpb_out[77][991],u_xpb_out[78][991],u_xpb_out[79][991],u_xpb_out[80][991],u_xpb_out[81][991],u_xpb_out[82][991],u_xpb_out[83][991],u_xpb_out[84][991],u_xpb_out[85][991],u_xpb_out[86][991],u_xpb_out[87][991],u_xpb_out[88][991],u_xpb_out[89][991],u_xpb_out[90][991],u_xpb_out[91][991],u_xpb_out[92][991],u_xpb_out[93][991],u_xpb_out[94][991],u_xpb_out[95][991],u_xpb_out[96][991],u_xpb_out[97][991],u_xpb_out[98][991],u_xpb_out[99][991],u_xpb_out[100][991],u_xpb_out[101][991],u_xpb_out[102][991],u_xpb_out[103][991],u_xpb_out[104][991],u_xpb_out[105][991]};

assign col_out_992 = {u_xpb_out[0][992],u_xpb_out[1][992],u_xpb_out[2][992],u_xpb_out[3][992],u_xpb_out[4][992],u_xpb_out[5][992],u_xpb_out[6][992],u_xpb_out[7][992],u_xpb_out[8][992],u_xpb_out[9][992],u_xpb_out[10][992],u_xpb_out[11][992],u_xpb_out[12][992],u_xpb_out[13][992],u_xpb_out[14][992],u_xpb_out[15][992],u_xpb_out[16][992],u_xpb_out[17][992],u_xpb_out[18][992],u_xpb_out[19][992],u_xpb_out[20][992],u_xpb_out[21][992],u_xpb_out[22][992],u_xpb_out[23][992],u_xpb_out[24][992],u_xpb_out[25][992],u_xpb_out[26][992],u_xpb_out[27][992],u_xpb_out[28][992],u_xpb_out[29][992],u_xpb_out[30][992],u_xpb_out[31][992],u_xpb_out[32][992],u_xpb_out[33][992],u_xpb_out[34][992],u_xpb_out[35][992],u_xpb_out[36][992],u_xpb_out[37][992],u_xpb_out[38][992],u_xpb_out[39][992],u_xpb_out[40][992],u_xpb_out[41][992],u_xpb_out[42][992],u_xpb_out[43][992],u_xpb_out[44][992],u_xpb_out[45][992],u_xpb_out[46][992],u_xpb_out[47][992],u_xpb_out[48][992],u_xpb_out[49][992],u_xpb_out[50][992],u_xpb_out[51][992],u_xpb_out[52][992],u_xpb_out[53][992],u_xpb_out[54][992],u_xpb_out[55][992],u_xpb_out[56][992],u_xpb_out[57][992],u_xpb_out[58][992],u_xpb_out[59][992],u_xpb_out[60][992],u_xpb_out[61][992],u_xpb_out[62][992],u_xpb_out[63][992],u_xpb_out[64][992],u_xpb_out[65][992],u_xpb_out[66][992],u_xpb_out[67][992],u_xpb_out[68][992],u_xpb_out[69][992],u_xpb_out[70][992],u_xpb_out[71][992],u_xpb_out[72][992],u_xpb_out[73][992],u_xpb_out[74][992],u_xpb_out[75][992],u_xpb_out[76][992],u_xpb_out[77][992],u_xpb_out[78][992],u_xpb_out[79][992],u_xpb_out[80][992],u_xpb_out[81][992],u_xpb_out[82][992],u_xpb_out[83][992],u_xpb_out[84][992],u_xpb_out[85][992],u_xpb_out[86][992],u_xpb_out[87][992],u_xpb_out[88][992],u_xpb_out[89][992],u_xpb_out[90][992],u_xpb_out[91][992],u_xpb_out[92][992],u_xpb_out[93][992],u_xpb_out[94][992],u_xpb_out[95][992],u_xpb_out[96][992],u_xpb_out[97][992],u_xpb_out[98][992],u_xpb_out[99][992],u_xpb_out[100][992],u_xpb_out[101][992],u_xpb_out[102][992],u_xpb_out[103][992],u_xpb_out[104][992],u_xpb_out[105][992]};

assign col_out_993 = {u_xpb_out[0][993],u_xpb_out[1][993],u_xpb_out[2][993],u_xpb_out[3][993],u_xpb_out[4][993],u_xpb_out[5][993],u_xpb_out[6][993],u_xpb_out[7][993],u_xpb_out[8][993],u_xpb_out[9][993],u_xpb_out[10][993],u_xpb_out[11][993],u_xpb_out[12][993],u_xpb_out[13][993],u_xpb_out[14][993],u_xpb_out[15][993],u_xpb_out[16][993],u_xpb_out[17][993],u_xpb_out[18][993],u_xpb_out[19][993],u_xpb_out[20][993],u_xpb_out[21][993],u_xpb_out[22][993],u_xpb_out[23][993],u_xpb_out[24][993],u_xpb_out[25][993],u_xpb_out[26][993],u_xpb_out[27][993],u_xpb_out[28][993],u_xpb_out[29][993],u_xpb_out[30][993],u_xpb_out[31][993],u_xpb_out[32][993],u_xpb_out[33][993],u_xpb_out[34][993],u_xpb_out[35][993],u_xpb_out[36][993],u_xpb_out[37][993],u_xpb_out[38][993],u_xpb_out[39][993],u_xpb_out[40][993],u_xpb_out[41][993],u_xpb_out[42][993],u_xpb_out[43][993],u_xpb_out[44][993],u_xpb_out[45][993],u_xpb_out[46][993],u_xpb_out[47][993],u_xpb_out[48][993],u_xpb_out[49][993],u_xpb_out[50][993],u_xpb_out[51][993],u_xpb_out[52][993],u_xpb_out[53][993],u_xpb_out[54][993],u_xpb_out[55][993],u_xpb_out[56][993],u_xpb_out[57][993],u_xpb_out[58][993],u_xpb_out[59][993],u_xpb_out[60][993],u_xpb_out[61][993],u_xpb_out[62][993],u_xpb_out[63][993],u_xpb_out[64][993],u_xpb_out[65][993],u_xpb_out[66][993],u_xpb_out[67][993],u_xpb_out[68][993],u_xpb_out[69][993],u_xpb_out[70][993],u_xpb_out[71][993],u_xpb_out[72][993],u_xpb_out[73][993],u_xpb_out[74][993],u_xpb_out[75][993],u_xpb_out[76][993],u_xpb_out[77][993],u_xpb_out[78][993],u_xpb_out[79][993],u_xpb_out[80][993],u_xpb_out[81][993],u_xpb_out[82][993],u_xpb_out[83][993],u_xpb_out[84][993],u_xpb_out[85][993],u_xpb_out[86][993],u_xpb_out[87][993],u_xpb_out[88][993],u_xpb_out[89][993],u_xpb_out[90][993],u_xpb_out[91][993],u_xpb_out[92][993],u_xpb_out[93][993],u_xpb_out[94][993],u_xpb_out[95][993],u_xpb_out[96][993],u_xpb_out[97][993],u_xpb_out[98][993],u_xpb_out[99][993],u_xpb_out[100][993],u_xpb_out[101][993],u_xpb_out[102][993],u_xpb_out[103][993],u_xpb_out[104][993],u_xpb_out[105][993]};

assign col_out_994 = {u_xpb_out[0][994],u_xpb_out[1][994],u_xpb_out[2][994],u_xpb_out[3][994],u_xpb_out[4][994],u_xpb_out[5][994],u_xpb_out[6][994],u_xpb_out[7][994],u_xpb_out[8][994],u_xpb_out[9][994],u_xpb_out[10][994],u_xpb_out[11][994],u_xpb_out[12][994],u_xpb_out[13][994],u_xpb_out[14][994],u_xpb_out[15][994],u_xpb_out[16][994],u_xpb_out[17][994],u_xpb_out[18][994],u_xpb_out[19][994],u_xpb_out[20][994],u_xpb_out[21][994],u_xpb_out[22][994],u_xpb_out[23][994],u_xpb_out[24][994],u_xpb_out[25][994],u_xpb_out[26][994],u_xpb_out[27][994],u_xpb_out[28][994],u_xpb_out[29][994],u_xpb_out[30][994],u_xpb_out[31][994],u_xpb_out[32][994],u_xpb_out[33][994],u_xpb_out[34][994],u_xpb_out[35][994],u_xpb_out[36][994],u_xpb_out[37][994],u_xpb_out[38][994],u_xpb_out[39][994],u_xpb_out[40][994],u_xpb_out[41][994],u_xpb_out[42][994],u_xpb_out[43][994],u_xpb_out[44][994],u_xpb_out[45][994],u_xpb_out[46][994],u_xpb_out[47][994],u_xpb_out[48][994],u_xpb_out[49][994],u_xpb_out[50][994],u_xpb_out[51][994],u_xpb_out[52][994],u_xpb_out[53][994],u_xpb_out[54][994],u_xpb_out[55][994],u_xpb_out[56][994],u_xpb_out[57][994],u_xpb_out[58][994],u_xpb_out[59][994],u_xpb_out[60][994],u_xpb_out[61][994],u_xpb_out[62][994],u_xpb_out[63][994],u_xpb_out[64][994],u_xpb_out[65][994],u_xpb_out[66][994],u_xpb_out[67][994],u_xpb_out[68][994],u_xpb_out[69][994],u_xpb_out[70][994],u_xpb_out[71][994],u_xpb_out[72][994],u_xpb_out[73][994],u_xpb_out[74][994],u_xpb_out[75][994],u_xpb_out[76][994],u_xpb_out[77][994],u_xpb_out[78][994],u_xpb_out[79][994],u_xpb_out[80][994],u_xpb_out[81][994],u_xpb_out[82][994],u_xpb_out[83][994],u_xpb_out[84][994],u_xpb_out[85][994],u_xpb_out[86][994],u_xpb_out[87][994],u_xpb_out[88][994],u_xpb_out[89][994],u_xpb_out[90][994],u_xpb_out[91][994],u_xpb_out[92][994],u_xpb_out[93][994],u_xpb_out[94][994],u_xpb_out[95][994],u_xpb_out[96][994],u_xpb_out[97][994],u_xpb_out[98][994],u_xpb_out[99][994],u_xpb_out[100][994],u_xpb_out[101][994],u_xpb_out[102][994],u_xpb_out[103][994],u_xpb_out[104][994],u_xpb_out[105][994]};

assign col_out_995 = {u_xpb_out[0][995],u_xpb_out[1][995],u_xpb_out[2][995],u_xpb_out[3][995],u_xpb_out[4][995],u_xpb_out[5][995],u_xpb_out[6][995],u_xpb_out[7][995],u_xpb_out[8][995],u_xpb_out[9][995],u_xpb_out[10][995],u_xpb_out[11][995],u_xpb_out[12][995],u_xpb_out[13][995],u_xpb_out[14][995],u_xpb_out[15][995],u_xpb_out[16][995],u_xpb_out[17][995],u_xpb_out[18][995],u_xpb_out[19][995],u_xpb_out[20][995],u_xpb_out[21][995],u_xpb_out[22][995],u_xpb_out[23][995],u_xpb_out[24][995],u_xpb_out[25][995],u_xpb_out[26][995],u_xpb_out[27][995],u_xpb_out[28][995],u_xpb_out[29][995],u_xpb_out[30][995],u_xpb_out[31][995],u_xpb_out[32][995],u_xpb_out[33][995],u_xpb_out[34][995],u_xpb_out[35][995],u_xpb_out[36][995],u_xpb_out[37][995],u_xpb_out[38][995],u_xpb_out[39][995],u_xpb_out[40][995],u_xpb_out[41][995],u_xpb_out[42][995],u_xpb_out[43][995],u_xpb_out[44][995],u_xpb_out[45][995],u_xpb_out[46][995],u_xpb_out[47][995],u_xpb_out[48][995],u_xpb_out[49][995],u_xpb_out[50][995],u_xpb_out[51][995],u_xpb_out[52][995],u_xpb_out[53][995],u_xpb_out[54][995],u_xpb_out[55][995],u_xpb_out[56][995],u_xpb_out[57][995],u_xpb_out[58][995],u_xpb_out[59][995],u_xpb_out[60][995],u_xpb_out[61][995],u_xpb_out[62][995],u_xpb_out[63][995],u_xpb_out[64][995],u_xpb_out[65][995],u_xpb_out[66][995],u_xpb_out[67][995],u_xpb_out[68][995],u_xpb_out[69][995],u_xpb_out[70][995],u_xpb_out[71][995],u_xpb_out[72][995],u_xpb_out[73][995],u_xpb_out[74][995],u_xpb_out[75][995],u_xpb_out[76][995],u_xpb_out[77][995],u_xpb_out[78][995],u_xpb_out[79][995],u_xpb_out[80][995],u_xpb_out[81][995],u_xpb_out[82][995],u_xpb_out[83][995],u_xpb_out[84][995],u_xpb_out[85][995],u_xpb_out[86][995],u_xpb_out[87][995],u_xpb_out[88][995],u_xpb_out[89][995],u_xpb_out[90][995],u_xpb_out[91][995],u_xpb_out[92][995],u_xpb_out[93][995],u_xpb_out[94][995],u_xpb_out[95][995],u_xpb_out[96][995],u_xpb_out[97][995],u_xpb_out[98][995],u_xpb_out[99][995],u_xpb_out[100][995],u_xpb_out[101][995],u_xpb_out[102][995],u_xpb_out[103][995],u_xpb_out[104][995],u_xpb_out[105][995]};

assign col_out_996 = {u_xpb_out[0][996],u_xpb_out[1][996],u_xpb_out[2][996],u_xpb_out[3][996],u_xpb_out[4][996],u_xpb_out[5][996],u_xpb_out[6][996],u_xpb_out[7][996],u_xpb_out[8][996],u_xpb_out[9][996],u_xpb_out[10][996],u_xpb_out[11][996],u_xpb_out[12][996],u_xpb_out[13][996],u_xpb_out[14][996],u_xpb_out[15][996],u_xpb_out[16][996],u_xpb_out[17][996],u_xpb_out[18][996],u_xpb_out[19][996],u_xpb_out[20][996],u_xpb_out[21][996],u_xpb_out[22][996],u_xpb_out[23][996],u_xpb_out[24][996],u_xpb_out[25][996],u_xpb_out[26][996],u_xpb_out[27][996],u_xpb_out[28][996],u_xpb_out[29][996],u_xpb_out[30][996],u_xpb_out[31][996],u_xpb_out[32][996],u_xpb_out[33][996],u_xpb_out[34][996],u_xpb_out[35][996],u_xpb_out[36][996],u_xpb_out[37][996],u_xpb_out[38][996],u_xpb_out[39][996],u_xpb_out[40][996],u_xpb_out[41][996],u_xpb_out[42][996],u_xpb_out[43][996],u_xpb_out[44][996],u_xpb_out[45][996],u_xpb_out[46][996],u_xpb_out[47][996],u_xpb_out[48][996],u_xpb_out[49][996],u_xpb_out[50][996],u_xpb_out[51][996],u_xpb_out[52][996],u_xpb_out[53][996],u_xpb_out[54][996],u_xpb_out[55][996],u_xpb_out[56][996],u_xpb_out[57][996],u_xpb_out[58][996],u_xpb_out[59][996],u_xpb_out[60][996],u_xpb_out[61][996],u_xpb_out[62][996],u_xpb_out[63][996],u_xpb_out[64][996],u_xpb_out[65][996],u_xpb_out[66][996],u_xpb_out[67][996],u_xpb_out[68][996],u_xpb_out[69][996],u_xpb_out[70][996],u_xpb_out[71][996],u_xpb_out[72][996],u_xpb_out[73][996],u_xpb_out[74][996],u_xpb_out[75][996],u_xpb_out[76][996],u_xpb_out[77][996],u_xpb_out[78][996],u_xpb_out[79][996],u_xpb_out[80][996],u_xpb_out[81][996],u_xpb_out[82][996],u_xpb_out[83][996],u_xpb_out[84][996],u_xpb_out[85][996],u_xpb_out[86][996],u_xpb_out[87][996],u_xpb_out[88][996],u_xpb_out[89][996],u_xpb_out[90][996],u_xpb_out[91][996],u_xpb_out[92][996],u_xpb_out[93][996],u_xpb_out[94][996],u_xpb_out[95][996],u_xpb_out[96][996],u_xpb_out[97][996],u_xpb_out[98][996],u_xpb_out[99][996],u_xpb_out[100][996],u_xpb_out[101][996],u_xpb_out[102][996],u_xpb_out[103][996],u_xpb_out[104][996],u_xpb_out[105][996]};

assign col_out_997 = {u_xpb_out[0][997],u_xpb_out[1][997],u_xpb_out[2][997],u_xpb_out[3][997],u_xpb_out[4][997],u_xpb_out[5][997],u_xpb_out[6][997],u_xpb_out[7][997],u_xpb_out[8][997],u_xpb_out[9][997],u_xpb_out[10][997],u_xpb_out[11][997],u_xpb_out[12][997],u_xpb_out[13][997],u_xpb_out[14][997],u_xpb_out[15][997],u_xpb_out[16][997],u_xpb_out[17][997],u_xpb_out[18][997],u_xpb_out[19][997],u_xpb_out[20][997],u_xpb_out[21][997],u_xpb_out[22][997],u_xpb_out[23][997],u_xpb_out[24][997],u_xpb_out[25][997],u_xpb_out[26][997],u_xpb_out[27][997],u_xpb_out[28][997],u_xpb_out[29][997],u_xpb_out[30][997],u_xpb_out[31][997],u_xpb_out[32][997],u_xpb_out[33][997],u_xpb_out[34][997],u_xpb_out[35][997],u_xpb_out[36][997],u_xpb_out[37][997],u_xpb_out[38][997],u_xpb_out[39][997],u_xpb_out[40][997],u_xpb_out[41][997],u_xpb_out[42][997],u_xpb_out[43][997],u_xpb_out[44][997],u_xpb_out[45][997],u_xpb_out[46][997],u_xpb_out[47][997],u_xpb_out[48][997],u_xpb_out[49][997],u_xpb_out[50][997],u_xpb_out[51][997],u_xpb_out[52][997],u_xpb_out[53][997],u_xpb_out[54][997],u_xpb_out[55][997],u_xpb_out[56][997],u_xpb_out[57][997],u_xpb_out[58][997],u_xpb_out[59][997],u_xpb_out[60][997],u_xpb_out[61][997],u_xpb_out[62][997],u_xpb_out[63][997],u_xpb_out[64][997],u_xpb_out[65][997],u_xpb_out[66][997],u_xpb_out[67][997],u_xpb_out[68][997],u_xpb_out[69][997],u_xpb_out[70][997],u_xpb_out[71][997],u_xpb_out[72][997],u_xpb_out[73][997],u_xpb_out[74][997],u_xpb_out[75][997],u_xpb_out[76][997],u_xpb_out[77][997],u_xpb_out[78][997],u_xpb_out[79][997],u_xpb_out[80][997],u_xpb_out[81][997],u_xpb_out[82][997],u_xpb_out[83][997],u_xpb_out[84][997],u_xpb_out[85][997],u_xpb_out[86][997],u_xpb_out[87][997],u_xpb_out[88][997],u_xpb_out[89][997],u_xpb_out[90][997],u_xpb_out[91][997],u_xpb_out[92][997],u_xpb_out[93][997],u_xpb_out[94][997],u_xpb_out[95][997],u_xpb_out[96][997],u_xpb_out[97][997],u_xpb_out[98][997],u_xpb_out[99][997],u_xpb_out[100][997],u_xpb_out[101][997],u_xpb_out[102][997],u_xpb_out[103][997],u_xpb_out[104][997],u_xpb_out[105][997]};

assign col_out_998 = {u_xpb_out[0][998],u_xpb_out[1][998],u_xpb_out[2][998],u_xpb_out[3][998],u_xpb_out[4][998],u_xpb_out[5][998],u_xpb_out[6][998],u_xpb_out[7][998],u_xpb_out[8][998],u_xpb_out[9][998],u_xpb_out[10][998],u_xpb_out[11][998],u_xpb_out[12][998],u_xpb_out[13][998],u_xpb_out[14][998],u_xpb_out[15][998],u_xpb_out[16][998],u_xpb_out[17][998],u_xpb_out[18][998],u_xpb_out[19][998],u_xpb_out[20][998],u_xpb_out[21][998],u_xpb_out[22][998],u_xpb_out[23][998],u_xpb_out[24][998],u_xpb_out[25][998],u_xpb_out[26][998],u_xpb_out[27][998],u_xpb_out[28][998],u_xpb_out[29][998],u_xpb_out[30][998],u_xpb_out[31][998],u_xpb_out[32][998],u_xpb_out[33][998],u_xpb_out[34][998],u_xpb_out[35][998],u_xpb_out[36][998],u_xpb_out[37][998],u_xpb_out[38][998],u_xpb_out[39][998],u_xpb_out[40][998],u_xpb_out[41][998],u_xpb_out[42][998],u_xpb_out[43][998],u_xpb_out[44][998],u_xpb_out[45][998],u_xpb_out[46][998],u_xpb_out[47][998],u_xpb_out[48][998],u_xpb_out[49][998],u_xpb_out[50][998],u_xpb_out[51][998],u_xpb_out[52][998],u_xpb_out[53][998],u_xpb_out[54][998],u_xpb_out[55][998],u_xpb_out[56][998],u_xpb_out[57][998],u_xpb_out[58][998],u_xpb_out[59][998],u_xpb_out[60][998],u_xpb_out[61][998],u_xpb_out[62][998],u_xpb_out[63][998],u_xpb_out[64][998],u_xpb_out[65][998],u_xpb_out[66][998],u_xpb_out[67][998],u_xpb_out[68][998],u_xpb_out[69][998],u_xpb_out[70][998],u_xpb_out[71][998],u_xpb_out[72][998],u_xpb_out[73][998],u_xpb_out[74][998],u_xpb_out[75][998],u_xpb_out[76][998],u_xpb_out[77][998],u_xpb_out[78][998],u_xpb_out[79][998],u_xpb_out[80][998],u_xpb_out[81][998],u_xpb_out[82][998],u_xpb_out[83][998],u_xpb_out[84][998],u_xpb_out[85][998],u_xpb_out[86][998],u_xpb_out[87][998],u_xpb_out[88][998],u_xpb_out[89][998],u_xpb_out[90][998],u_xpb_out[91][998],u_xpb_out[92][998],u_xpb_out[93][998],u_xpb_out[94][998],u_xpb_out[95][998],u_xpb_out[96][998],u_xpb_out[97][998],u_xpb_out[98][998],u_xpb_out[99][998],u_xpb_out[100][998],u_xpb_out[101][998],u_xpb_out[102][998],u_xpb_out[103][998],u_xpb_out[104][998],u_xpb_out[105][998]};

assign col_out_999 = {u_xpb_out[0][999],u_xpb_out[1][999],u_xpb_out[2][999],u_xpb_out[3][999],u_xpb_out[4][999],u_xpb_out[5][999],u_xpb_out[6][999],u_xpb_out[7][999],u_xpb_out[8][999],u_xpb_out[9][999],u_xpb_out[10][999],u_xpb_out[11][999],u_xpb_out[12][999],u_xpb_out[13][999],u_xpb_out[14][999],u_xpb_out[15][999],u_xpb_out[16][999],u_xpb_out[17][999],u_xpb_out[18][999],u_xpb_out[19][999],u_xpb_out[20][999],u_xpb_out[21][999],u_xpb_out[22][999],u_xpb_out[23][999],u_xpb_out[24][999],u_xpb_out[25][999],u_xpb_out[26][999],u_xpb_out[27][999],u_xpb_out[28][999],u_xpb_out[29][999],u_xpb_out[30][999],u_xpb_out[31][999],u_xpb_out[32][999],u_xpb_out[33][999],u_xpb_out[34][999],u_xpb_out[35][999],u_xpb_out[36][999],u_xpb_out[37][999],u_xpb_out[38][999],u_xpb_out[39][999],u_xpb_out[40][999],u_xpb_out[41][999],u_xpb_out[42][999],u_xpb_out[43][999],u_xpb_out[44][999],u_xpb_out[45][999],u_xpb_out[46][999],u_xpb_out[47][999],u_xpb_out[48][999],u_xpb_out[49][999],u_xpb_out[50][999],u_xpb_out[51][999],u_xpb_out[52][999],u_xpb_out[53][999],u_xpb_out[54][999],u_xpb_out[55][999],u_xpb_out[56][999],u_xpb_out[57][999],u_xpb_out[58][999],u_xpb_out[59][999],u_xpb_out[60][999],u_xpb_out[61][999],u_xpb_out[62][999],u_xpb_out[63][999],u_xpb_out[64][999],u_xpb_out[65][999],u_xpb_out[66][999],u_xpb_out[67][999],u_xpb_out[68][999],u_xpb_out[69][999],u_xpb_out[70][999],u_xpb_out[71][999],u_xpb_out[72][999],u_xpb_out[73][999],u_xpb_out[74][999],u_xpb_out[75][999],u_xpb_out[76][999],u_xpb_out[77][999],u_xpb_out[78][999],u_xpb_out[79][999],u_xpb_out[80][999],u_xpb_out[81][999],u_xpb_out[82][999],u_xpb_out[83][999],u_xpb_out[84][999],u_xpb_out[85][999],u_xpb_out[86][999],u_xpb_out[87][999],u_xpb_out[88][999],u_xpb_out[89][999],u_xpb_out[90][999],u_xpb_out[91][999],u_xpb_out[92][999],u_xpb_out[93][999],u_xpb_out[94][999],u_xpb_out[95][999],u_xpb_out[96][999],u_xpb_out[97][999],u_xpb_out[98][999],u_xpb_out[99][999],u_xpb_out[100][999],u_xpb_out[101][999],u_xpb_out[102][999],u_xpb_out[103][999],u_xpb_out[104][999],u_xpb_out[105][999]};

assign col_out_1000 = {u_xpb_out[0][1000],u_xpb_out[1][1000],u_xpb_out[2][1000],u_xpb_out[3][1000],u_xpb_out[4][1000],u_xpb_out[5][1000],u_xpb_out[6][1000],u_xpb_out[7][1000],u_xpb_out[8][1000],u_xpb_out[9][1000],u_xpb_out[10][1000],u_xpb_out[11][1000],u_xpb_out[12][1000],u_xpb_out[13][1000],u_xpb_out[14][1000],u_xpb_out[15][1000],u_xpb_out[16][1000],u_xpb_out[17][1000],u_xpb_out[18][1000],u_xpb_out[19][1000],u_xpb_out[20][1000],u_xpb_out[21][1000],u_xpb_out[22][1000],u_xpb_out[23][1000],u_xpb_out[24][1000],u_xpb_out[25][1000],u_xpb_out[26][1000],u_xpb_out[27][1000],u_xpb_out[28][1000],u_xpb_out[29][1000],u_xpb_out[30][1000],u_xpb_out[31][1000],u_xpb_out[32][1000],u_xpb_out[33][1000],u_xpb_out[34][1000],u_xpb_out[35][1000],u_xpb_out[36][1000],u_xpb_out[37][1000],u_xpb_out[38][1000],u_xpb_out[39][1000],u_xpb_out[40][1000],u_xpb_out[41][1000],u_xpb_out[42][1000],u_xpb_out[43][1000],u_xpb_out[44][1000],u_xpb_out[45][1000],u_xpb_out[46][1000],u_xpb_out[47][1000],u_xpb_out[48][1000],u_xpb_out[49][1000],u_xpb_out[50][1000],u_xpb_out[51][1000],u_xpb_out[52][1000],u_xpb_out[53][1000],u_xpb_out[54][1000],u_xpb_out[55][1000],u_xpb_out[56][1000],u_xpb_out[57][1000],u_xpb_out[58][1000],u_xpb_out[59][1000],u_xpb_out[60][1000],u_xpb_out[61][1000],u_xpb_out[62][1000],u_xpb_out[63][1000],u_xpb_out[64][1000],u_xpb_out[65][1000],u_xpb_out[66][1000],u_xpb_out[67][1000],u_xpb_out[68][1000],u_xpb_out[69][1000],u_xpb_out[70][1000],u_xpb_out[71][1000],u_xpb_out[72][1000],u_xpb_out[73][1000],u_xpb_out[74][1000],u_xpb_out[75][1000],u_xpb_out[76][1000],u_xpb_out[77][1000],u_xpb_out[78][1000],u_xpb_out[79][1000],u_xpb_out[80][1000],u_xpb_out[81][1000],u_xpb_out[82][1000],u_xpb_out[83][1000],u_xpb_out[84][1000],u_xpb_out[85][1000],u_xpb_out[86][1000],u_xpb_out[87][1000],u_xpb_out[88][1000],u_xpb_out[89][1000],u_xpb_out[90][1000],u_xpb_out[91][1000],u_xpb_out[92][1000],u_xpb_out[93][1000],u_xpb_out[94][1000],u_xpb_out[95][1000],u_xpb_out[96][1000],u_xpb_out[97][1000],u_xpb_out[98][1000],u_xpb_out[99][1000],u_xpb_out[100][1000],u_xpb_out[101][1000],u_xpb_out[102][1000],u_xpb_out[103][1000],u_xpb_out[104][1000],u_xpb_out[105][1000]};

assign col_out_1001 = {u_xpb_out[0][1001],u_xpb_out[1][1001],u_xpb_out[2][1001],u_xpb_out[3][1001],u_xpb_out[4][1001],u_xpb_out[5][1001],u_xpb_out[6][1001],u_xpb_out[7][1001],u_xpb_out[8][1001],u_xpb_out[9][1001],u_xpb_out[10][1001],u_xpb_out[11][1001],u_xpb_out[12][1001],u_xpb_out[13][1001],u_xpb_out[14][1001],u_xpb_out[15][1001],u_xpb_out[16][1001],u_xpb_out[17][1001],u_xpb_out[18][1001],u_xpb_out[19][1001],u_xpb_out[20][1001],u_xpb_out[21][1001],u_xpb_out[22][1001],u_xpb_out[23][1001],u_xpb_out[24][1001],u_xpb_out[25][1001],u_xpb_out[26][1001],u_xpb_out[27][1001],u_xpb_out[28][1001],u_xpb_out[29][1001],u_xpb_out[30][1001],u_xpb_out[31][1001],u_xpb_out[32][1001],u_xpb_out[33][1001],u_xpb_out[34][1001],u_xpb_out[35][1001],u_xpb_out[36][1001],u_xpb_out[37][1001],u_xpb_out[38][1001],u_xpb_out[39][1001],u_xpb_out[40][1001],u_xpb_out[41][1001],u_xpb_out[42][1001],u_xpb_out[43][1001],u_xpb_out[44][1001],u_xpb_out[45][1001],u_xpb_out[46][1001],u_xpb_out[47][1001],u_xpb_out[48][1001],u_xpb_out[49][1001],u_xpb_out[50][1001],u_xpb_out[51][1001],u_xpb_out[52][1001],u_xpb_out[53][1001],u_xpb_out[54][1001],u_xpb_out[55][1001],u_xpb_out[56][1001],u_xpb_out[57][1001],u_xpb_out[58][1001],u_xpb_out[59][1001],u_xpb_out[60][1001],u_xpb_out[61][1001],u_xpb_out[62][1001],u_xpb_out[63][1001],u_xpb_out[64][1001],u_xpb_out[65][1001],u_xpb_out[66][1001],u_xpb_out[67][1001],u_xpb_out[68][1001],u_xpb_out[69][1001],u_xpb_out[70][1001],u_xpb_out[71][1001],u_xpb_out[72][1001],u_xpb_out[73][1001],u_xpb_out[74][1001],u_xpb_out[75][1001],u_xpb_out[76][1001],u_xpb_out[77][1001],u_xpb_out[78][1001],u_xpb_out[79][1001],u_xpb_out[80][1001],u_xpb_out[81][1001],u_xpb_out[82][1001],u_xpb_out[83][1001],u_xpb_out[84][1001],u_xpb_out[85][1001],u_xpb_out[86][1001],u_xpb_out[87][1001],u_xpb_out[88][1001],u_xpb_out[89][1001],u_xpb_out[90][1001],u_xpb_out[91][1001],u_xpb_out[92][1001],u_xpb_out[93][1001],u_xpb_out[94][1001],u_xpb_out[95][1001],u_xpb_out[96][1001],u_xpb_out[97][1001],u_xpb_out[98][1001],u_xpb_out[99][1001],u_xpb_out[100][1001],u_xpb_out[101][1001],u_xpb_out[102][1001],u_xpb_out[103][1001],u_xpb_out[104][1001],u_xpb_out[105][1001]};

assign col_out_1002 = {u_xpb_out[0][1002],u_xpb_out[1][1002],u_xpb_out[2][1002],u_xpb_out[3][1002],u_xpb_out[4][1002],u_xpb_out[5][1002],u_xpb_out[6][1002],u_xpb_out[7][1002],u_xpb_out[8][1002],u_xpb_out[9][1002],u_xpb_out[10][1002],u_xpb_out[11][1002],u_xpb_out[12][1002],u_xpb_out[13][1002],u_xpb_out[14][1002],u_xpb_out[15][1002],u_xpb_out[16][1002],u_xpb_out[17][1002],u_xpb_out[18][1002],u_xpb_out[19][1002],u_xpb_out[20][1002],u_xpb_out[21][1002],u_xpb_out[22][1002],u_xpb_out[23][1002],u_xpb_out[24][1002],u_xpb_out[25][1002],u_xpb_out[26][1002],u_xpb_out[27][1002],u_xpb_out[28][1002],u_xpb_out[29][1002],u_xpb_out[30][1002],u_xpb_out[31][1002],u_xpb_out[32][1002],u_xpb_out[33][1002],u_xpb_out[34][1002],u_xpb_out[35][1002],u_xpb_out[36][1002],u_xpb_out[37][1002],u_xpb_out[38][1002],u_xpb_out[39][1002],u_xpb_out[40][1002],u_xpb_out[41][1002],u_xpb_out[42][1002],u_xpb_out[43][1002],u_xpb_out[44][1002],u_xpb_out[45][1002],u_xpb_out[46][1002],u_xpb_out[47][1002],u_xpb_out[48][1002],u_xpb_out[49][1002],u_xpb_out[50][1002],u_xpb_out[51][1002],u_xpb_out[52][1002],u_xpb_out[53][1002],u_xpb_out[54][1002],u_xpb_out[55][1002],u_xpb_out[56][1002],u_xpb_out[57][1002],u_xpb_out[58][1002],u_xpb_out[59][1002],u_xpb_out[60][1002],u_xpb_out[61][1002],u_xpb_out[62][1002],u_xpb_out[63][1002],u_xpb_out[64][1002],u_xpb_out[65][1002],u_xpb_out[66][1002],u_xpb_out[67][1002],u_xpb_out[68][1002],u_xpb_out[69][1002],u_xpb_out[70][1002],u_xpb_out[71][1002],u_xpb_out[72][1002],u_xpb_out[73][1002],u_xpb_out[74][1002],u_xpb_out[75][1002],u_xpb_out[76][1002],u_xpb_out[77][1002],u_xpb_out[78][1002],u_xpb_out[79][1002],u_xpb_out[80][1002],u_xpb_out[81][1002],u_xpb_out[82][1002],u_xpb_out[83][1002],u_xpb_out[84][1002],u_xpb_out[85][1002],u_xpb_out[86][1002],u_xpb_out[87][1002],u_xpb_out[88][1002],u_xpb_out[89][1002],u_xpb_out[90][1002],u_xpb_out[91][1002],u_xpb_out[92][1002],u_xpb_out[93][1002],u_xpb_out[94][1002],u_xpb_out[95][1002],u_xpb_out[96][1002],u_xpb_out[97][1002],u_xpb_out[98][1002],u_xpb_out[99][1002],u_xpb_out[100][1002],u_xpb_out[101][1002],u_xpb_out[102][1002],u_xpb_out[103][1002],u_xpb_out[104][1002],u_xpb_out[105][1002]};

assign col_out_1003 = {u_xpb_out[0][1003],u_xpb_out[1][1003],u_xpb_out[2][1003],u_xpb_out[3][1003],u_xpb_out[4][1003],u_xpb_out[5][1003],u_xpb_out[6][1003],u_xpb_out[7][1003],u_xpb_out[8][1003],u_xpb_out[9][1003],u_xpb_out[10][1003],u_xpb_out[11][1003],u_xpb_out[12][1003],u_xpb_out[13][1003],u_xpb_out[14][1003],u_xpb_out[15][1003],u_xpb_out[16][1003],u_xpb_out[17][1003],u_xpb_out[18][1003],u_xpb_out[19][1003],u_xpb_out[20][1003],u_xpb_out[21][1003],u_xpb_out[22][1003],u_xpb_out[23][1003],u_xpb_out[24][1003],u_xpb_out[25][1003],u_xpb_out[26][1003],u_xpb_out[27][1003],u_xpb_out[28][1003],u_xpb_out[29][1003],u_xpb_out[30][1003],u_xpb_out[31][1003],u_xpb_out[32][1003],u_xpb_out[33][1003],u_xpb_out[34][1003],u_xpb_out[35][1003],u_xpb_out[36][1003],u_xpb_out[37][1003],u_xpb_out[38][1003],u_xpb_out[39][1003],u_xpb_out[40][1003],u_xpb_out[41][1003],u_xpb_out[42][1003],u_xpb_out[43][1003],u_xpb_out[44][1003],u_xpb_out[45][1003],u_xpb_out[46][1003],u_xpb_out[47][1003],u_xpb_out[48][1003],u_xpb_out[49][1003],u_xpb_out[50][1003],u_xpb_out[51][1003],u_xpb_out[52][1003],u_xpb_out[53][1003],u_xpb_out[54][1003],u_xpb_out[55][1003],u_xpb_out[56][1003],u_xpb_out[57][1003],u_xpb_out[58][1003],u_xpb_out[59][1003],u_xpb_out[60][1003],u_xpb_out[61][1003],u_xpb_out[62][1003],u_xpb_out[63][1003],u_xpb_out[64][1003],u_xpb_out[65][1003],u_xpb_out[66][1003],u_xpb_out[67][1003],u_xpb_out[68][1003],u_xpb_out[69][1003],u_xpb_out[70][1003],u_xpb_out[71][1003],u_xpb_out[72][1003],u_xpb_out[73][1003],u_xpb_out[74][1003],u_xpb_out[75][1003],u_xpb_out[76][1003],u_xpb_out[77][1003],u_xpb_out[78][1003],u_xpb_out[79][1003],u_xpb_out[80][1003],u_xpb_out[81][1003],u_xpb_out[82][1003],u_xpb_out[83][1003],u_xpb_out[84][1003],u_xpb_out[85][1003],u_xpb_out[86][1003],u_xpb_out[87][1003],u_xpb_out[88][1003],u_xpb_out[89][1003],u_xpb_out[90][1003],u_xpb_out[91][1003],u_xpb_out[92][1003],u_xpb_out[93][1003],u_xpb_out[94][1003],u_xpb_out[95][1003],u_xpb_out[96][1003],u_xpb_out[97][1003],u_xpb_out[98][1003],u_xpb_out[99][1003],u_xpb_out[100][1003],u_xpb_out[101][1003],u_xpb_out[102][1003],u_xpb_out[103][1003],u_xpb_out[104][1003],u_xpb_out[105][1003]};

assign col_out_1004 = {u_xpb_out[0][1004],u_xpb_out[1][1004],u_xpb_out[2][1004],u_xpb_out[3][1004],u_xpb_out[4][1004],u_xpb_out[5][1004],u_xpb_out[6][1004],u_xpb_out[7][1004],u_xpb_out[8][1004],u_xpb_out[9][1004],u_xpb_out[10][1004],u_xpb_out[11][1004],u_xpb_out[12][1004],u_xpb_out[13][1004],u_xpb_out[14][1004],u_xpb_out[15][1004],u_xpb_out[16][1004],u_xpb_out[17][1004],u_xpb_out[18][1004],u_xpb_out[19][1004],u_xpb_out[20][1004],u_xpb_out[21][1004],u_xpb_out[22][1004],u_xpb_out[23][1004],u_xpb_out[24][1004],u_xpb_out[25][1004],u_xpb_out[26][1004],u_xpb_out[27][1004],u_xpb_out[28][1004],u_xpb_out[29][1004],u_xpb_out[30][1004],u_xpb_out[31][1004],u_xpb_out[32][1004],u_xpb_out[33][1004],u_xpb_out[34][1004],u_xpb_out[35][1004],u_xpb_out[36][1004],u_xpb_out[37][1004],u_xpb_out[38][1004],u_xpb_out[39][1004],u_xpb_out[40][1004],u_xpb_out[41][1004],u_xpb_out[42][1004],u_xpb_out[43][1004],u_xpb_out[44][1004],u_xpb_out[45][1004],u_xpb_out[46][1004],u_xpb_out[47][1004],u_xpb_out[48][1004],u_xpb_out[49][1004],u_xpb_out[50][1004],u_xpb_out[51][1004],u_xpb_out[52][1004],u_xpb_out[53][1004],u_xpb_out[54][1004],u_xpb_out[55][1004],u_xpb_out[56][1004],u_xpb_out[57][1004],u_xpb_out[58][1004],u_xpb_out[59][1004],u_xpb_out[60][1004],u_xpb_out[61][1004],u_xpb_out[62][1004],u_xpb_out[63][1004],u_xpb_out[64][1004],u_xpb_out[65][1004],u_xpb_out[66][1004],u_xpb_out[67][1004],u_xpb_out[68][1004],u_xpb_out[69][1004],u_xpb_out[70][1004],u_xpb_out[71][1004],u_xpb_out[72][1004],u_xpb_out[73][1004],u_xpb_out[74][1004],u_xpb_out[75][1004],u_xpb_out[76][1004],u_xpb_out[77][1004],u_xpb_out[78][1004],u_xpb_out[79][1004],u_xpb_out[80][1004],u_xpb_out[81][1004],u_xpb_out[82][1004],u_xpb_out[83][1004],u_xpb_out[84][1004],u_xpb_out[85][1004],u_xpb_out[86][1004],u_xpb_out[87][1004],u_xpb_out[88][1004],u_xpb_out[89][1004],u_xpb_out[90][1004],u_xpb_out[91][1004],u_xpb_out[92][1004],u_xpb_out[93][1004],u_xpb_out[94][1004],u_xpb_out[95][1004],u_xpb_out[96][1004],u_xpb_out[97][1004],u_xpb_out[98][1004],u_xpb_out[99][1004],u_xpb_out[100][1004],u_xpb_out[101][1004],u_xpb_out[102][1004],u_xpb_out[103][1004],u_xpb_out[104][1004],u_xpb_out[105][1004]};

assign col_out_1005 = {u_xpb_out[0][1005],u_xpb_out[1][1005],u_xpb_out[2][1005],u_xpb_out[3][1005],u_xpb_out[4][1005],u_xpb_out[5][1005],u_xpb_out[6][1005],u_xpb_out[7][1005],u_xpb_out[8][1005],u_xpb_out[9][1005],u_xpb_out[10][1005],u_xpb_out[11][1005],u_xpb_out[12][1005],u_xpb_out[13][1005],u_xpb_out[14][1005],u_xpb_out[15][1005],u_xpb_out[16][1005],u_xpb_out[17][1005],u_xpb_out[18][1005],u_xpb_out[19][1005],u_xpb_out[20][1005],u_xpb_out[21][1005],u_xpb_out[22][1005],u_xpb_out[23][1005],u_xpb_out[24][1005],u_xpb_out[25][1005],u_xpb_out[26][1005],u_xpb_out[27][1005],u_xpb_out[28][1005],u_xpb_out[29][1005],u_xpb_out[30][1005],u_xpb_out[31][1005],u_xpb_out[32][1005],u_xpb_out[33][1005],u_xpb_out[34][1005],u_xpb_out[35][1005],u_xpb_out[36][1005],u_xpb_out[37][1005],u_xpb_out[38][1005],u_xpb_out[39][1005],u_xpb_out[40][1005],u_xpb_out[41][1005],u_xpb_out[42][1005],u_xpb_out[43][1005],u_xpb_out[44][1005],u_xpb_out[45][1005],u_xpb_out[46][1005],u_xpb_out[47][1005],u_xpb_out[48][1005],u_xpb_out[49][1005],u_xpb_out[50][1005],u_xpb_out[51][1005],u_xpb_out[52][1005],u_xpb_out[53][1005],u_xpb_out[54][1005],u_xpb_out[55][1005],u_xpb_out[56][1005],u_xpb_out[57][1005],u_xpb_out[58][1005],u_xpb_out[59][1005],u_xpb_out[60][1005],u_xpb_out[61][1005],u_xpb_out[62][1005],u_xpb_out[63][1005],u_xpb_out[64][1005],u_xpb_out[65][1005],u_xpb_out[66][1005],u_xpb_out[67][1005],u_xpb_out[68][1005],u_xpb_out[69][1005],u_xpb_out[70][1005],u_xpb_out[71][1005],u_xpb_out[72][1005],u_xpb_out[73][1005],u_xpb_out[74][1005],u_xpb_out[75][1005],u_xpb_out[76][1005],u_xpb_out[77][1005],u_xpb_out[78][1005],u_xpb_out[79][1005],u_xpb_out[80][1005],u_xpb_out[81][1005],u_xpb_out[82][1005],u_xpb_out[83][1005],u_xpb_out[84][1005],u_xpb_out[85][1005],u_xpb_out[86][1005],u_xpb_out[87][1005],u_xpb_out[88][1005],u_xpb_out[89][1005],u_xpb_out[90][1005],u_xpb_out[91][1005],u_xpb_out[92][1005],u_xpb_out[93][1005],u_xpb_out[94][1005],u_xpb_out[95][1005],u_xpb_out[96][1005],u_xpb_out[97][1005],u_xpb_out[98][1005],u_xpb_out[99][1005],u_xpb_out[100][1005],u_xpb_out[101][1005],u_xpb_out[102][1005],u_xpb_out[103][1005],u_xpb_out[104][1005],u_xpb_out[105][1005]};

assign col_out_1006 = {u_xpb_out[0][1006],u_xpb_out[1][1006],u_xpb_out[2][1006],u_xpb_out[3][1006],u_xpb_out[4][1006],u_xpb_out[5][1006],u_xpb_out[6][1006],u_xpb_out[7][1006],u_xpb_out[8][1006],u_xpb_out[9][1006],u_xpb_out[10][1006],u_xpb_out[11][1006],u_xpb_out[12][1006],u_xpb_out[13][1006],u_xpb_out[14][1006],u_xpb_out[15][1006],u_xpb_out[16][1006],u_xpb_out[17][1006],u_xpb_out[18][1006],u_xpb_out[19][1006],u_xpb_out[20][1006],u_xpb_out[21][1006],u_xpb_out[22][1006],u_xpb_out[23][1006],u_xpb_out[24][1006],u_xpb_out[25][1006],u_xpb_out[26][1006],u_xpb_out[27][1006],u_xpb_out[28][1006],u_xpb_out[29][1006],u_xpb_out[30][1006],u_xpb_out[31][1006],u_xpb_out[32][1006],u_xpb_out[33][1006],u_xpb_out[34][1006],u_xpb_out[35][1006],u_xpb_out[36][1006],u_xpb_out[37][1006],u_xpb_out[38][1006],u_xpb_out[39][1006],u_xpb_out[40][1006],u_xpb_out[41][1006],u_xpb_out[42][1006],u_xpb_out[43][1006],u_xpb_out[44][1006],u_xpb_out[45][1006],u_xpb_out[46][1006],u_xpb_out[47][1006],u_xpb_out[48][1006],u_xpb_out[49][1006],u_xpb_out[50][1006],u_xpb_out[51][1006],u_xpb_out[52][1006],u_xpb_out[53][1006],u_xpb_out[54][1006],u_xpb_out[55][1006],u_xpb_out[56][1006],u_xpb_out[57][1006],u_xpb_out[58][1006],u_xpb_out[59][1006],u_xpb_out[60][1006],u_xpb_out[61][1006],u_xpb_out[62][1006],u_xpb_out[63][1006],u_xpb_out[64][1006],u_xpb_out[65][1006],u_xpb_out[66][1006],u_xpb_out[67][1006],u_xpb_out[68][1006],u_xpb_out[69][1006],u_xpb_out[70][1006],u_xpb_out[71][1006],u_xpb_out[72][1006],u_xpb_out[73][1006],u_xpb_out[74][1006],u_xpb_out[75][1006],u_xpb_out[76][1006],u_xpb_out[77][1006],u_xpb_out[78][1006],u_xpb_out[79][1006],u_xpb_out[80][1006],u_xpb_out[81][1006],u_xpb_out[82][1006],u_xpb_out[83][1006],u_xpb_out[84][1006],u_xpb_out[85][1006],u_xpb_out[86][1006],u_xpb_out[87][1006],u_xpb_out[88][1006],u_xpb_out[89][1006],u_xpb_out[90][1006],u_xpb_out[91][1006],u_xpb_out[92][1006],u_xpb_out[93][1006],u_xpb_out[94][1006],u_xpb_out[95][1006],u_xpb_out[96][1006],u_xpb_out[97][1006],u_xpb_out[98][1006],u_xpb_out[99][1006],u_xpb_out[100][1006],u_xpb_out[101][1006],u_xpb_out[102][1006],u_xpb_out[103][1006],u_xpb_out[104][1006],u_xpb_out[105][1006]};

assign col_out_1007 = {u_xpb_out[0][1007],u_xpb_out[1][1007],u_xpb_out[2][1007],u_xpb_out[3][1007],u_xpb_out[4][1007],u_xpb_out[5][1007],u_xpb_out[6][1007],u_xpb_out[7][1007],u_xpb_out[8][1007],u_xpb_out[9][1007],u_xpb_out[10][1007],u_xpb_out[11][1007],u_xpb_out[12][1007],u_xpb_out[13][1007],u_xpb_out[14][1007],u_xpb_out[15][1007],u_xpb_out[16][1007],u_xpb_out[17][1007],u_xpb_out[18][1007],u_xpb_out[19][1007],u_xpb_out[20][1007],u_xpb_out[21][1007],u_xpb_out[22][1007],u_xpb_out[23][1007],u_xpb_out[24][1007],u_xpb_out[25][1007],u_xpb_out[26][1007],u_xpb_out[27][1007],u_xpb_out[28][1007],u_xpb_out[29][1007],u_xpb_out[30][1007],u_xpb_out[31][1007],u_xpb_out[32][1007],u_xpb_out[33][1007],u_xpb_out[34][1007],u_xpb_out[35][1007],u_xpb_out[36][1007],u_xpb_out[37][1007],u_xpb_out[38][1007],u_xpb_out[39][1007],u_xpb_out[40][1007],u_xpb_out[41][1007],u_xpb_out[42][1007],u_xpb_out[43][1007],u_xpb_out[44][1007],u_xpb_out[45][1007],u_xpb_out[46][1007],u_xpb_out[47][1007],u_xpb_out[48][1007],u_xpb_out[49][1007],u_xpb_out[50][1007],u_xpb_out[51][1007],u_xpb_out[52][1007],u_xpb_out[53][1007],u_xpb_out[54][1007],u_xpb_out[55][1007],u_xpb_out[56][1007],u_xpb_out[57][1007],u_xpb_out[58][1007],u_xpb_out[59][1007],u_xpb_out[60][1007],u_xpb_out[61][1007],u_xpb_out[62][1007],u_xpb_out[63][1007],u_xpb_out[64][1007],u_xpb_out[65][1007],u_xpb_out[66][1007],u_xpb_out[67][1007],u_xpb_out[68][1007],u_xpb_out[69][1007],u_xpb_out[70][1007],u_xpb_out[71][1007],u_xpb_out[72][1007],u_xpb_out[73][1007],u_xpb_out[74][1007],u_xpb_out[75][1007],u_xpb_out[76][1007],u_xpb_out[77][1007],u_xpb_out[78][1007],u_xpb_out[79][1007],u_xpb_out[80][1007],u_xpb_out[81][1007],u_xpb_out[82][1007],u_xpb_out[83][1007],u_xpb_out[84][1007],u_xpb_out[85][1007],u_xpb_out[86][1007],u_xpb_out[87][1007],u_xpb_out[88][1007],u_xpb_out[89][1007],u_xpb_out[90][1007],u_xpb_out[91][1007],u_xpb_out[92][1007],u_xpb_out[93][1007],u_xpb_out[94][1007],u_xpb_out[95][1007],u_xpb_out[96][1007],u_xpb_out[97][1007],u_xpb_out[98][1007],u_xpb_out[99][1007],u_xpb_out[100][1007],u_xpb_out[101][1007],u_xpb_out[102][1007],u_xpb_out[103][1007],u_xpb_out[104][1007],u_xpb_out[105][1007]};

assign col_out_1008 = {u_xpb_out[0][1008],u_xpb_out[1][1008],u_xpb_out[2][1008],u_xpb_out[3][1008],u_xpb_out[4][1008],u_xpb_out[5][1008],u_xpb_out[6][1008],u_xpb_out[7][1008],u_xpb_out[8][1008],u_xpb_out[9][1008],u_xpb_out[10][1008],u_xpb_out[11][1008],u_xpb_out[12][1008],u_xpb_out[13][1008],u_xpb_out[14][1008],u_xpb_out[15][1008],u_xpb_out[16][1008],u_xpb_out[17][1008],u_xpb_out[18][1008],u_xpb_out[19][1008],u_xpb_out[20][1008],u_xpb_out[21][1008],u_xpb_out[22][1008],u_xpb_out[23][1008],u_xpb_out[24][1008],u_xpb_out[25][1008],u_xpb_out[26][1008],u_xpb_out[27][1008],u_xpb_out[28][1008],u_xpb_out[29][1008],u_xpb_out[30][1008],u_xpb_out[31][1008],u_xpb_out[32][1008],u_xpb_out[33][1008],u_xpb_out[34][1008],u_xpb_out[35][1008],u_xpb_out[36][1008],u_xpb_out[37][1008],u_xpb_out[38][1008],u_xpb_out[39][1008],u_xpb_out[40][1008],u_xpb_out[41][1008],u_xpb_out[42][1008],u_xpb_out[43][1008],u_xpb_out[44][1008],u_xpb_out[45][1008],u_xpb_out[46][1008],u_xpb_out[47][1008],u_xpb_out[48][1008],u_xpb_out[49][1008],u_xpb_out[50][1008],u_xpb_out[51][1008],u_xpb_out[52][1008],u_xpb_out[53][1008],u_xpb_out[54][1008],u_xpb_out[55][1008],u_xpb_out[56][1008],u_xpb_out[57][1008],u_xpb_out[58][1008],u_xpb_out[59][1008],u_xpb_out[60][1008],u_xpb_out[61][1008],u_xpb_out[62][1008],u_xpb_out[63][1008],u_xpb_out[64][1008],u_xpb_out[65][1008],u_xpb_out[66][1008],u_xpb_out[67][1008],u_xpb_out[68][1008],u_xpb_out[69][1008],u_xpb_out[70][1008],u_xpb_out[71][1008],u_xpb_out[72][1008],u_xpb_out[73][1008],u_xpb_out[74][1008],u_xpb_out[75][1008],u_xpb_out[76][1008],u_xpb_out[77][1008],u_xpb_out[78][1008],u_xpb_out[79][1008],u_xpb_out[80][1008],u_xpb_out[81][1008],u_xpb_out[82][1008],u_xpb_out[83][1008],u_xpb_out[84][1008],u_xpb_out[85][1008],u_xpb_out[86][1008],u_xpb_out[87][1008],u_xpb_out[88][1008],u_xpb_out[89][1008],u_xpb_out[90][1008],u_xpb_out[91][1008],u_xpb_out[92][1008],u_xpb_out[93][1008],u_xpb_out[94][1008],u_xpb_out[95][1008],u_xpb_out[96][1008],u_xpb_out[97][1008],u_xpb_out[98][1008],u_xpb_out[99][1008],u_xpb_out[100][1008],u_xpb_out[101][1008],u_xpb_out[102][1008],u_xpb_out[103][1008],u_xpb_out[104][1008],u_xpb_out[105][1008]};

assign col_out_1009 = {u_xpb_out[0][1009],u_xpb_out[1][1009],u_xpb_out[2][1009],u_xpb_out[3][1009],u_xpb_out[4][1009],u_xpb_out[5][1009],u_xpb_out[6][1009],u_xpb_out[7][1009],u_xpb_out[8][1009],u_xpb_out[9][1009],u_xpb_out[10][1009],u_xpb_out[11][1009],u_xpb_out[12][1009],u_xpb_out[13][1009],u_xpb_out[14][1009],u_xpb_out[15][1009],u_xpb_out[16][1009],u_xpb_out[17][1009],u_xpb_out[18][1009],u_xpb_out[19][1009],u_xpb_out[20][1009],u_xpb_out[21][1009],u_xpb_out[22][1009],u_xpb_out[23][1009],u_xpb_out[24][1009],u_xpb_out[25][1009],u_xpb_out[26][1009],u_xpb_out[27][1009],u_xpb_out[28][1009],u_xpb_out[29][1009],u_xpb_out[30][1009],u_xpb_out[31][1009],u_xpb_out[32][1009],u_xpb_out[33][1009],u_xpb_out[34][1009],u_xpb_out[35][1009],u_xpb_out[36][1009],u_xpb_out[37][1009],u_xpb_out[38][1009],u_xpb_out[39][1009],u_xpb_out[40][1009],u_xpb_out[41][1009],u_xpb_out[42][1009],u_xpb_out[43][1009],u_xpb_out[44][1009],u_xpb_out[45][1009],u_xpb_out[46][1009],u_xpb_out[47][1009],u_xpb_out[48][1009],u_xpb_out[49][1009],u_xpb_out[50][1009],u_xpb_out[51][1009],u_xpb_out[52][1009],u_xpb_out[53][1009],u_xpb_out[54][1009],u_xpb_out[55][1009],u_xpb_out[56][1009],u_xpb_out[57][1009],u_xpb_out[58][1009],u_xpb_out[59][1009],u_xpb_out[60][1009],u_xpb_out[61][1009],u_xpb_out[62][1009],u_xpb_out[63][1009],u_xpb_out[64][1009],u_xpb_out[65][1009],u_xpb_out[66][1009],u_xpb_out[67][1009],u_xpb_out[68][1009],u_xpb_out[69][1009],u_xpb_out[70][1009],u_xpb_out[71][1009],u_xpb_out[72][1009],u_xpb_out[73][1009],u_xpb_out[74][1009],u_xpb_out[75][1009],u_xpb_out[76][1009],u_xpb_out[77][1009],u_xpb_out[78][1009],u_xpb_out[79][1009],u_xpb_out[80][1009],u_xpb_out[81][1009],u_xpb_out[82][1009],u_xpb_out[83][1009],u_xpb_out[84][1009],u_xpb_out[85][1009],u_xpb_out[86][1009],u_xpb_out[87][1009],u_xpb_out[88][1009],u_xpb_out[89][1009],u_xpb_out[90][1009],u_xpb_out[91][1009],u_xpb_out[92][1009],u_xpb_out[93][1009],u_xpb_out[94][1009],u_xpb_out[95][1009],u_xpb_out[96][1009],u_xpb_out[97][1009],u_xpb_out[98][1009],u_xpb_out[99][1009],u_xpb_out[100][1009],u_xpb_out[101][1009],u_xpb_out[102][1009],u_xpb_out[103][1009],u_xpb_out[104][1009],u_xpb_out[105][1009]};

assign col_out_1010 = {u_xpb_out[0][1010],u_xpb_out[1][1010],u_xpb_out[2][1010],u_xpb_out[3][1010],u_xpb_out[4][1010],u_xpb_out[5][1010],u_xpb_out[6][1010],u_xpb_out[7][1010],u_xpb_out[8][1010],u_xpb_out[9][1010],u_xpb_out[10][1010],u_xpb_out[11][1010],u_xpb_out[12][1010],u_xpb_out[13][1010],u_xpb_out[14][1010],u_xpb_out[15][1010],u_xpb_out[16][1010],u_xpb_out[17][1010],u_xpb_out[18][1010],u_xpb_out[19][1010],u_xpb_out[20][1010],u_xpb_out[21][1010],u_xpb_out[22][1010],u_xpb_out[23][1010],u_xpb_out[24][1010],u_xpb_out[25][1010],u_xpb_out[26][1010],u_xpb_out[27][1010],u_xpb_out[28][1010],u_xpb_out[29][1010],u_xpb_out[30][1010],u_xpb_out[31][1010],u_xpb_out[32][1010],u_xpb_out[33][1010],u_xpb_out[34][1010],u_xpb_out[35][1010],u_xpb_out[36][1010],u_xpb_out[37][1010],u_xpb_out[38][1010],u_xpb_out[39][1010],u_xpb_out[40][1010],u_xpb_out[41][1010],u_xpb_out[42][1010],u_xpb_out[43][1010],u_xpb_out[44][1010],u_xpb_out[45][1010],u_xpb_out[46][1010],u_xpb_out[47][1010],u_xpb_out[48][1010],u_xpb_out[49][1010],u_xpb_out[50][1010],u_xpb_out[51][1010],u_xpb_out[52][1010],u_xpb_out[53][1010],u_xpb_out[54][1010],u_xpb_out[55][1010],u_xpb_out[56][1010],u_xpb_out[57][1010],u_xpb_out[58][1010],u_xpb_out[59][1010],u_xpb_out[60][1010],u_xpb_out[61][1010],u_xpb_out[62][1010],u_xpb_out[63][1010],u_xpb_out[64][1010],u_xpb_out[65][1010],u_xpb_out[66][1010],u_xpb_out[67][1010],u_xpb_out[68][1010],u_xpb_out[69][1010],u_xpb_out[70][1010],u_xpb_out[71][1010],u_xpb_out[72][1010],u_xpb_out[73][1010],u_xpb_out[74][1010],u_xpb_out[75][1010],u_xpb_out[76][1010],u_xpb_out[77][1010],u_xpb_out[78][1010],u_xpb_out[79][1010],u_xpb_out[80][1010],u_xpb_out[81][1010],u_xpb_out[82][1010],u_xpb_out[83][1010],u_xpb_out[84][1010],u_xpb_out[85][1010],u_xpb_out[86][1010],u_xpb_out[87][1010],u_xpb_out[88][1010],u_xpb_out[89][1010],u_xpb_out[90][1010],u_xpb_out[91][1010],u_xpb_out[92][1010],u_xpb_out[93][1010],u_xpb_out[94][1010],u_xpb_out[95][1010],u_xpb_out[96][1010],u_xpb_out[97][1010],u_xpb_out[98][1010],u_xpb_out[99][1010],u_xpb_out[100][1010],u_xpb_out[101][1010],u_xpb_out[102][1010],u_xpb_out[103][1010],u_xpb_out[104][1010],u_xpb_out[105][1010]};

assign col_out_1011 = {u_xpb_out[0][1011],u_xpb_out[1][1011],u_xpb_out[2][1011],u_xpb_out[3][1011],u_xpb_out[4][1011],u_xpb_out[5][1011],u_xpb_out[6][1011],u_xpb_out[7][1011],u_xpb_out[8][1011],u_xpb_out[9][1011],u_xpb_out[10][1011],u_xpb_out[11][1011],u_xpb_out[12][1011],u_xpb_out[13][1011],u_xpb_out[14][1011],u_xpb_out[15][1011],u_xpb_out[16][1011],u_xpb_out[17][1011],u_xpb_out[18][1011],u_xpb_out[19][1011],u_xpb_out[20][1011],u_xpb_out[21][1011],u_xpb_out[22][1011],u_xpb_out[23][1011],u_xpb_out[24][1011],u_xpb_out[25][1011],u_xpb_out[26][1011],u_xpb_out[27][1011],u_xpb_out[28][1011],u_xpb_out[29][1011],u_xpb_out[30][1011],u_xpb_out[31][1011],u_xpb_out[32][1011],u_xpb_out[33][1011],u_xpb_out[34][1011],u_xpb_out[35][1011],u_xpb_out[36][1011],u_xpb_out[37][1011],u_xpb_out[38][1011],u_xpb_out[39][1011],u_xpb_out[40][1011],u_xpb_out[41][1011],u_xpb_out[42][1011],u_xpb_out[43][1011],u_xpb_out[44][1011],u_xpb_out[45][1011],u_xpb_out[46][1011],u_xpb_out[47][1011],u_xpb_out[48][1011],u_xpb_out[49][1011],u_xpb_out[50][1011],u_xpb_out[51][1011],u_xpb_out[52][1011],u_xpb_out[53][1011],u_xpb_out[54][1011],u_xpb_out[55][1011],u_xpb_out[56][1011],u_xpb_out[57][1011],u_xpb_out[58][1011],u_xpb_out[59][1011],u_xpb_out[60][1011],u_xpb_out[61][1011],u_xpb_out[62][1011],u_xpb_out[63][1011],u_xpb_out[64][1011],u_xpb_out[65][1011],u_xpb_out[66][1011],u_xpb_out[67][1011],u_xpb_out[68][1011],u_xpb_out[69][1011],u_xpb_out[70][1011],u_xpb_out[71][1011],u_xpb_out[72][1011],u_xpb_out[73][1011],u_xpb_out[74][1011],u_xpb_out[75][1011],u_xpb_out[76][1011],u_xpb_out[77][1011],u_xpb_out[78][1011],u_xpb_out[79][1011],u_xpb_out[80][1011],u_xpb_out[81][1011],u_xpb_out[82][1011],u_xpb_out[83][1011],u_xpb_out[84][1011],u_xpb_out[85][1011],u_xpb_out[86][1011],u_xpb_out[87][1011],u_xpb_out[88][1011],u_xpb_out[89][1011],u_xpb_out[90][1011],u_xpb_out[91][1011],u_xpb_out[92][1011],u_xpb_out[93][1011],u_xpb_out[94][1011],u_xpb_out[95][1011],u_xpb_out[96][1011],u_xpb_out[97][1011],u_xpb_out[98][1011],u_xpb_out[99][1011],u_xpb_out[100][1011],u_xpb_out[101][1011],u_xpb_out[102][1011],u_xpb_out[103][1011],u_xpb_out[104][1011],u_xpb_out[105][1011]};

assign col_out_1012 = {u_xpb_out[0][1012],u_xpb_out[1][1012],u_xpb_out[2][1012],u_xpb_out[3][1012],u_xpb_out[4][1012],u_xpb_out[5][1012],u_xpb_out[6][1012],u_xpb_out[7][1012],u_xpb_out[8][1012],u_xpb_out[9][1012],u_xpb_out[10][1012],u_xpb_out[11][1012],u_xpb_out[12][1012],u_xpb_out[13][1012],u_xpb_out[14][1012],u_xpb_out[15][1012],u_xpb_out[16][1012],u_xpb_out[17][1012],u_xpb_out[18][1012],u_xpb_out[19][1012],u_xpb_out[20][1012],u_xpb_out[21][1012],u_xpb_out[22][1012],u_xpb_out[23][1012],u_xpb_out[24][1012],u_xpb_out[25][1012],u_xpb_out[26][1012],u_xpb_out[27][1012],u_xpb_out[28][1012],u_xpb_out[29][1012],u_xpb_out[30][1012],u_xpb_out[31][1012],u_xpb_out[32][1012],u_xpb_out[33][1012],u_xpb_out[34][1012],u_xpb_out[35][1012],u_xpb_out[36][1012],u_xpb_out[37][1012],u_xpb_out[38][1012],u_xpb_out[39][1012],u_xpb_out[40][1012],u_xpb_out[41][1012],u_xpb_out[42][1012],u_xpb_out[43][1012],u_xpb_out[44][1012],u_xpb_out[45][1012],u_xpb_out[46][1012],u_xpb_out[47][1012],u_xpb_out[48][1012],u_xpb_out[49][1012],u_xpb_out[50][1012],u_xpb_out[51][1012],u_xpb_out[52][1012],u_xpb_out[53][1012],u_xpb_out[54][1012],u_xpb_out[55][1012],u_xpb_out[56][1012],u_xpb_out[57][1012],u_xpb_out[58][1012],u_xpb_out[59][1012],u_xpb_out[60][1012],u_xpb_out[61][1012],u_xpb_out[62][1012],u_xpb_out[63][1012],u_xpb_out[64][1012],u_xpb_out[65][1012],u_xpb_out[66][1012],u_xpb_out[67][1012],u_xpb_out[68][1012],u_xpb_out[69][1012],u_xpb_out[70][1012],u_xpb_out[71][1012],u_xpb_out[72][1012],u_xpb_out[73][1012],u_xpb_out[74][1012],u_xpb_out[75][1012],u_xpb_out[76][1012],u_xpb_out[77][1012],u_xpb_out[78][1012],u_xpb_out[79][1012],u_xpb_out[80][1012],u_xpb_out[81][1012],u_xpb_out[82][1012],u_xpb_out[83][1012],u_xpb_out[84][1012],u_xpb_out[85][1012],u_xpb_out[86][1012],u_xpb_out[87][1012],u_xpb_out[88][1012],u_xpb_out[89][1012],u_xpb_out[90][1012],u_xpb_out[91][1012],u_xpb_out[92][1012],u_xpb_out[93][1012],u_xpb_out[94][1012],u_xpb_out[95][1012],u_xpb_out[96][1012],u_xpb_out[97][1012],u_xpb_out[98][1012],u_xpb_out[99][1012],u_xpb_out[100][1012],u_xpb_out[101][1012],u_xpb_out[102][1012],u_xpb_out[103][1012],u_xpb_out[104][1012],u_xpb_out[105][1012]};

assign col_out_1013 = {u_xpb_out[0][1013],u_xpb_out[1][1013],u_xpb_out[2][1013],u_xpb_out[3][1013],u_xpb_out[4][1013],u_xpb_out[5][1013],u_xpb_out[6][1013],u_xpb_out[7][1013],u_xpb_out[8][1013],u_xpb_out[9][1013],u_xpb_out[10][1013],u_xpb_out[11][1013],u_xpb_out[12][1013],u_xpb_out[13][1013],u_xpb_out[14][1013],u_xpb_out[15][1013],u_xpb_out[16][1013],u_xpb_out[17][1013],u_xpb_out[18][1013],u_xpb_out[19][1013],u_xpb_out[20][1013],u_xpb_out[21][1013],u_xpb_out[22][1013],u_xpb_out[23][1013],u_xpb_out[24][1013],u_xpb_out[25][1013],u_xpb_out[26][1013],u_xpb_out[27][1013],u_xpb_out[28][1013],u_xpb_out[29][1013],u_xpb_out[30][1013],u_xpb_out[31][1013],u_xpb_out[32][1013],u_xpb_out[33][1013],u_xpb_out[34][1013],u_xpb_out[35][1013],u_xpb_out[36][1013],u_xpb_out[37][1013],u_xpb_out[38][1013],u_xpb_out[39][1013],u_xpb_out[40][1013],u_xpb_out[41][1013],u_xpb_out[42][1013],u_xpb_out[43][1013],u_xpb_out[44][1013],u_xpb_out[45][1013],u_xpb_out[46][1013],u_xpb_out[47][1013],u_xpb_out[48][1013],u_xpb_out[49][1013],u_xpb_out[50][1013],u_xpb_out[51][1013],u_xpb_out[52][1013],u_xpb_out[53][1013],u_xpb_out[54][1013],u_xpb_out[55][1013],u_xpb_out[56][1013],u_xpb_out[57][1013],u_xpb_out[58][1013],u_xpb_out[59][1013],u_xpb_out[60][1013],u_xpb_out[61][1013],u_xpb_out[62][1013],u_xpb_out[63][1013],u_xpb_out[64][1013],u_xpb_out[65][1013],u_xpb_out[66][1013],u_xpb_out[67][1013],u_xpb_out[68][1013],u_xpb_out[69][1013],u_xpb_out[70][1013],u_xpb_out[71][1013],u_xpb_out[72][1013],u_xpb_out[73][1013],u_xpb_out[74][1013],u_xpb_out[75][1013],u_xpb_out[76][1013],u_xpb_out[77][1013],u_xpb_out[78][1013],u_xpb_out[79][1013],u_xpb_out[80][1013],u_xpb_out[81][1013],u_xpb_out[82][1013],u_xpb_out[83][1013],u_xpb_out[84][1013],u_xpb_out[85][1013],u_xpb_out[86][1013],u_xpb_out[87][1013],u_xpb_out[88][1013],u_xpb_out[89][1013],u_xpb_out[90][1013],u_xpb_out[91][1013],u_xpb_out[92][1013],u_xpb_out[93][1013],u_xpb_out[94][1013],u_xpb_out[95][1013],u_xpb_out[96][1013],u_xpb_out[97][1013],u_xpb_out[98][1013],u_xpb_out[99][1013],u_xpb_out[100][1013],u_xpb_out[101][1013],u_xpb_out[102][1013],u_xpb_out[103][1013],u_xpb_out[104][1013],u_xpb_out[105][1013]};

assign col_out_1014 = {u_xpb_out[0][1014],u_xpb_out[1][1014],u_xpb_out[2][1014],u_xpb_out[3][1014],u_xpb_out[4][1014],u_xpb_out[5][1014],u_xpb_out[6][1014],u_xpb_out[7][1014],u_xpb_out[8][1014],u_xpb_out[9][1014],u_xpb_out[10][1014],u_xpb_out[11][1014],u_xpb_out[12][1014],u_xpb_out[13][1014],u_xpb_out[14][1014],u_xpb_out[15][1014],u_xpb_out[16][1014],u_xpb_out[17][1014],u_xpb_out[18][1014],u_xpb_out[19][1014],u_xpb_out[20][1014],u_xpb_out[21][1014],u_xpb_out[22][1014],u_xpb_out[23][1014],u_xpb_out[24][1014],u_xpb_out[25][1014],u_xpb_out[26][1014],u_xpb_out[27][1014],u_xpb_out[28][1014],u_xpb_out[29][1014],u_xpb_out[30][1014],u_xpb_out[31][1014],u_xpb_out[32][1014],u_xpb_out[33][1014],u_xpb_out[34][1014],u_xpb_out[35][1014],u_xpb_out[36][1014],u_xpb_out[37][1014],u_xpb_out[38][1014],u_xpb_out[39][1014],u_xpb_out[40][1014],u_xpb_out[41][1014],u_xpb_out[42][1014],u_xpb_out[43][1014],u_xpb_out[44][1014],u_xpb_out[45][1014],u_xpb_out[46][1014],u_xpb_out[47][1014],u_xpb_out[48][1014],u_xpb_out[49][1014],u_xpb_out[50][1014],u_xpb_out[51][1014],u_xpb_out[52][1014],u_xpb_out[53][1014],u_xpb_out[54][1014],u_xpb_out[55][1014],u_xpb_out[56][1014],u_xpb_out[57][1014],u_xpb_out[58][1014],u_xpb_out[59][1014],u_xpb_out[60][1014],u_xpb_out[61][1014],u_xpb_out[62][1014],u_xpb_out[63][1014],u_xpb_out[64][1014],u_xpb_out[65][1014],u_xpb_out[66][1014],u_xpb_out[67][1014],u_xpb_out[68][1014],u_xpb_out[69][1014],u_xpb_out[70][1014],u_xpb_out[71][1014],u_xpb_out[72][1014],u_xpb_out[73][1014],u_xpb_out[74][1014],u_xpb_out[75][1014],u_xpb_out[76][1014],u_xpb_out[77][1014],u_xpb_out[78][1014],u_xpb_out[79][1014],u_xpb_out[80][1014],u_xpb_out[81][1014],u_xpb_out[82][1014],u_xpb_out[83][1014],u_xpb_out[84][1014],u_xpb_out[85][1014],u_xpb_out[86][1014],u_xpb_out[87][1014],u_xpb_out[88][1014],u_xpb_out[89][1014],u_xpb_out[90][1014],u_xpb_out[91][1014],u_xpb_out[92][1014],u_xpb_out[93][1014],u_xpb_out[94][1014],u_xpb_out[95][1014],u_xpb_out[96][1014],u_xpb_out[97][1014],u_xpb_out[98][1014],u_xpb_out[99][1014],u_xpb_out[100][1014],u_xpb_out[101][1014],u_xpb_out[102][1014],u_xpb_out[103][1014],u_xpb_out[104][1014],u_xpb_out[105][1014]};

assign col_out_1015 = {u_xpb_out[0][1015],u_xpb_out[1][1015],u_xpb_out[2][1015],u_xpb_out[3][1015],u_xpb_out[4][1015],u_xpb_out[5][1015],u_xpb_out[6][1015],u_xpb_out[7][1015],u_xpb_out[8][1015],u_xpb_out[9][1015],u_xpb_out[10][1015],u_xpb_out[11][1015],u_xpb_out[12][1015],u_xpb_out[13][1015],u_xpb_out[14][1015],u_xpb_out[15][1015],u_xpb_out[16][1015],u_xpb_out[17][1015],u_xpb_out[18][1015],u_xpb_out[19][1015],u_xpb_out[20][1015],u_xpb_out[21][1015],u_xpb_out[22][1015],u_xpb_out[23][1015],u_xpb_out[24][1015],u_xpb_out[25][1015],u_xpb_out[26][1015],u_xpb_out[27][1015],u_xpb_out[28][1015],u_xpb_out[29][1015],u_xpb_out[30][1015],u_xpb_out[31][1015],u_xpb_out[32][1015],u_xpb_out[33][1015],u_xpb_out[34][1015],u_xpb_out[35][1015],u_xpb_out[36][1015],u_xpb_out[37][1015],u_xpb_out[38][1015],u_xpb_out[39][1015],u_xpb_out[40][1015],u_xpb_out[41][1015],u_xpb_out[42][1015],u_xpb_out[43][1015],u_xpb_out[44][1015],u_xpb_out[45][1015],u_xpb_out[46][1015],u_xpb_out[47][1015],u_xpb_out[48][1015],u_xpb_out[49][1015],u_xpb_out[50][1015],u_xpb_out[51][1015],u_xpb_out[52][1015],u_xpb_out[53][1015],u_xpb_out[54][1015],u_xpb_out[55][1015],u_xpb_out[56][1015],u_xpb_out[57][1015],u_xpb_out[58][1015],u_xpb_out[59][1015],u_xpb_out[60][1015],u_xpb_out[61][1015],u_xpb_out[62][1015],u_xpb_out[63][1015],u_xpb_out[64][1015],u_xpb_out[65][1015],u_xpb_out[66][1015],u_xpb_out[67][1015],u_xpb_out[68][1015],u_xpb_out[69][1015],u_xpb_out[70][1015],u_xpb_out[71][1015],u_xpb_out[72][1015],u_xpb_out[73][1015],u_xpb_out[74][1015],u_xpb_out[75][1015],u_xpb_out[76][1015],u_xpb_out[77][1015],u_xpb_out[78][1015],u_xpb_out[79][1015],u_xpb_out[80][1015],u_xpb_out[81][1015],u_xpb_out[82][1015],u_xpb_out[83][1015],u_xpb_out[84][1015],u_xpb_out[85][1015],u_xpb_out[86][1015],u_xpb_out[87][1015],u_xpb_out[88][1015],u_xpb_out[89][1015],u_xpb_out[90][1015],u_xpb_out[91][1015],u_xpb_out[92][1015],u_xpb_out[93][1015],u_xpb_out[94][1015],u_xpb_out[95][1015],u_xpb_out[96][1015],u_xpb_out[97][1015],u_xpb_out[98][1015],u_xpb_out[99][1015],u_xpb_out[100][1015],u_xpb_out[101][1015],u_xpb_out[102][1015],u_xpb_out[103][1015],u_xpb_out[104][1015],u_xpb_out[105][1015]};

assign col_out_1016 = {u_xpb_out[0][1016],u_xpb_out[1][1016],u_xpb_out[2][1016],u_xpb_out[3][1016],u_xpb_out[4][1016],u_xpb_out[5][1016],u_xpb_out[6][1016],u_xpb_out[7][1016],u_xpb_out[8][1016],u_xpb_out[9][1016],u_xpb_out[10][1016],u_xpb_out[11][1016],u_xpb_out[12][1016],u_xpb_out[13][1016],u_xpb_out[14][1016],u_xpb_out[15][1016],u_xpb_out[16][1016],u_xpb_out[17][1016],u_xpb_out[18][1016],u_xpb_out[19][1016],u_xpb_out[20][1016],u_xpb_out[21][1016],u_xpb_out[22][1016],u_xpb_out[23][1016],u_xpb_out[24][1016],u_xpb_out[25][1016],u_xpb_out[26][1016],u_xpb_out[27][1016],u_xpb_out[28][1016],u_xpb_out[29][1016],u_xpb_out[30][1016],u_xpb_out[31][1016],u_xpb_out[32][1016],u_xpb_out[33][1016],u_xpb_out[34][1016],u_xpb_out[35][1016],u_xpb_out[36][1016],u_xpb_out[37][1016],u_xpb_out[38][1016],u_xpb_out[39][1016],u_xpb_out[40][1016],u_xpb_out[41][1016],u_xpb_out[42][1016],u_xpb_out[43][1016],u_xpb_out[44][1016],u_xpb_out[45][1016],u_xpb_out[46][1016],u_xpb_out[47][1016],u_xpb_out[48][1016],u_xpb_out[49][1016],u_xpb_out[50][1016],u_xpb_out[51][1016],u_xpb_out[52][1016],u_xpb_out[53][1016],u_xpb_out[54][1016],u_xpb_out[55][1016],u_xpb_out[56][1016],u_xpb_out[57][1016],u_xpb_out[58][1016],u_xpb_out[59][1016],u_xpb_out[60][1016],u_xpb_out[61][1016],u_xpb_out[62][1016],u_xpb_out[63][1016],u_xpb_out[64][1016],u_xpb_out[65][1016],u_xpb_out[66][1016],u_xpb_out[67][1016],u_xpb_out[68][1016],u_xpb_out[69][1016],u_xpb_out[70][1016],u_xpb_out[71][1016],u_xpb_out[72][1016],u_xpb_out[73][1016],u_xpb_out[74][1016],u_xpb_out[75][1016],u_xpb_out[76][1016],u_xpb_out[77][1016],u_xpb_out[78][1016],u_xpb_out[79][1016],u_xpb_out[80][1016],u_xpb_out[81][1016],u_xpb_out[82][1016],u_xpb_out[83][1016],u_xpb_out[84][1016],u_xpb_out[85][1016],u_xpb_out[86][1016],u_xpb_out[87][1016],u_xpb_out[88][1016],u_xpb_out[89][1016],u_xpb_out[90][1016],u_xpb_out[91][1016],u_xpb_out[92][1016],u_xpb_out[93][1016],u_xpb_out[94][1016],u_xpb_out[95][1016],u_xpb_out[96][1016],u_xpb_out[97][1016],u_xpb_out[98][1016],u_xpb_out[99][1016],u_xpb_out[100][1016],u_xpb_out[101][1016],u_xpb_out[102][1016],u_xpb_out[103][1016],u_xpb_out[104][1016],u_xpb_out[105][1016]};

assign col_out_1017 = {u_xpb_out[0][1017],u_xpb_out[1][1017],u_xpb_out[2][1017],u_xpb_out[3][1017],u_xpb_out[4][1017],u_xpb_out[5][1017],u_xpb_out[6][1017],u_xpb_out[7][1017],u_xpb_out[8][1017],u_xpb_out[9][1017],u_xpb_out[10][1017],u_xpb_out[11][1017],u_xpb_out[12][1017],u_xpb_out[13][1017],u_xpb_out[14][1017],u_xpb_out[15][1017],u_xpb_out[16][1017],u_xpb_out[17][1017],u_xpb_out[18][1017],u_xpb_out[19][1017],u_xpb_out[20][1017],u_xpb_out[21][1017],u_xpb_out[22][1017],u_xpb_out[23][1017],u_xpb_out[24][1017],u_xpb_out[25][1017],u_xpb_out[26][1017],u_xpb_out[27][1017],u_xpb_out[28][1017],u_xpb_out[29][1017],u_xpb_out[30][1017],u_xpb_out[31][1017],u_xpb_out[32][1017],u_xpb_out[33][1017],u_xpb_out[34][1017],u_xpb_out[35][1017],u_xpb_out[36][1017],u_xpb_out[37][1017],u_xpb_out[38][1017],u_xpb_out[39][1017],u_xpb_out[40][1017],u_xpb_out[41][1017],u_xpb_out[42][1017],u_xpb_out[43][1017],u_xpb_out[44][1017],u_xpb_out[45][1017],u_xpb_out[46][1017],u_xpb_out[47][1017],u_xpb_out[48][1017],u_xpb_out[49][1017],u_xpb_out[50][1017],u_xpb_out[51][1017],u_xpb_out[52][1017],u_xpb_out[53][1017],u_xpb_out[54][1017],u_xpb_out[55][1017],u_xpb_out[56][1017],u_xpb_out[57][1017],u_xpb_out[58][1017],u_xpb_out[59][1017],u_xpb_out[60][1017],u_xpb_out[61][1017],u_xpb_out[62][1017],u_xpb_out[63][1017],u_xpb_out[64][1017],u_xpb_out[65][1017],u_xpb_out[66][1017],u_xpb_out[67][1017],u_xpb_out[68][1017],u_xpb_out[69][1017],u_xpb_out[70][1017],u_xpb_out[71][1017],u_xpb_out[72][1017],u_xpb_out[73][1017],u_xpb_out[74][1017],u_xpb_out[75][1017],u_xpb_out[76][1017],u_xpb_out[77][1017],u_xpb_out[78][1017],u_xpb_out[79][1017],u_xpb_out[80][1017],u_xpb_out[81][1017],u_xpb_out[82][1017],u_xpb_out[83][1017],u_xpb_out[84][1017],u_xpb_out[85][1017],u_xpb_out[86][1017],u_xpb_out[87][1017],u_xpb_out[88][1017],u_xpb_out[89][1017],u_xpb_out[90][1017],u_xpb_out[91][1017],u_xpb_out[92][1017],u_xpb_out[93][1017],u_xpb_out[94][1017],u_xpb_out[95][1017],u_xpb_out[96][1017],u_xpb_out[97][1017],u_xpb_out[98][1017],u_xpb_out[99][1017],u_xpb_out[100][1017],u_xpb_out[101][1017],u_xpb_out[102][1017],u_xpb_out[103][1017],u_xpb_out[104][1017],u_xpb_out[105][1017]};

assign col_out_1018 = {u_xpb_out[0][1018],u_xpb_out[1][1018],u_xpb_out[2][1018],u_xpb_out[3][1018],u_xpb_out[4][1018],u_xpb_out[5][1018],u_xpb_out[6][1018],u_xpb_out[7][1018],u_xpb_out[8][1018],u_xpb_out[9][1018],u_xpb_out[10][1018],u_xpb_out[11][1018],u_xpb_out[12][1018],u_xpb_out[13][1018],u_xpb_out[14][1018],u_xpb_out[15][1018],u_xpb_out[16][1018],u_xpb_out[17][1018],u_xpb_out[18][1018],u_xpb_out[19][1018],u_xpb_out[20][1018],u_xpb_out[21][1018],u_xpb_out[22][1018],u_xpb_out[23][1018],u_xpb_out[24][1018],u_xpb_out[25][1018],u_xpb_out[26][1018],u_xpb_out[27][1018],u_xpb_out[28][1018],u_xpb_out[29][1018],u_xpb_out[30][1018],u_xpb_out[31][1018],u_xpb_out[32][1018],u_xpb_out[33][1018],u_xpb_out[34][1018],u_xpb_out[35][1018],u_xpb_out[36][1018],u_xpb_out[37][1018],u_xpb_out[38][1018],u_xpb_out[39][1018],u_xpb_out[40][1018],u_xpb_out[41][1018],u_xpb_out[42][1018],u_xpb_out[43][1018],u_xpb_out[44][1018],u_xpb_out[45][1018],u_xpb_out[46][1018],u_xpb_out[47][1018],u_xpb_out[48][1018],u_xpb_out[49][1018],u_xpb_out[50][1018],u_xpb_out[51][1018],u_xpb_out[52][1018],u_xpb_out[53][1018],u_xpb_out[54][1018],u_xpb_out[55][1018],u_xpb_out[56][1018],u_xpb_out[57][1018],u_xpb_out[58][1018],u_xpb_out[59][1018],u_xpb_out[60][1018],u_xpb_out[61][1018],u_xpb_out[62][1018],u_xpb_out[63][1018],u_xpb_out[64][1018],u_xpb_out[65][1018],u_xpb_out[66][1018],u_xpb_out[67][1018],u_xpb_out[68][1018],u_xpb_out[69][1018],u_xpb_out[70][1018],u_xpb_out[71][1018],u_xpb_out[72][1018],u_xpb_out[73][1018],u_xpb_out[74][1018],u_xpb_out[75][1018],u_xpb_out[76][1018],u_xpb_out[77][1018],u_xpb_out[78][1018],u_xpb_out[79][1018],u_xpb_out[80][1018],u_xpb_out[81][1018],u_xpb_out[82][1018],u_xpb_out[83][1018],u_xpb_out[84][1018],u_xpb_out[85][1018],u_xpb_out[86][1018],u_xpb_out[87][1018],u_xpb_out[88][1018],u_xpb_out[89][1018],u_xpb_out[90][1018],u_xpb_out[91][1018],u_xpb_out[92][1018],u_xpb_out[93][1018],u_xpb_out[94][1018],u_xpb_out[95][1018],u_xpb_out[96][1018],u_xpb_out[97][1018],u_xpb_out[98][1018],u_xpb_out[99][1018],u_xpb_out[100][1018],u_xpb_out[101][1018],u_xpb_out[102][1018],u_xpb_out[103][1018],u_xpb_out[104][1018],u_xpb_out[105][1018]};

assign col_out_1019 = {u_xpb_out[0][1019],u_xpb_out[1][1019],u_xpb_out[2][1019],u_xpb_out[3][1019],u_xpb_out[4][1019],u_xpb_out[5][1019],u_xpb_out[6][1019],u_xpb_out[7][1019],u_xpb_out[8][1019],u_xpb_out[9][1019],u_xpb_out[10][1019],u_xpb_out[11][1019],u_xpb_out[12][1019],u_xpb_out[13][1019],u_xpb_out[14][1019],u_xpb_out[15][1019],u_xpb_out[16][1019],u_xpb_out[17][1019],u_xpb_out[18][1019],u_xpb_out[19][1019],u_xpb_out[20][1019],u_xpb_out[21][1019],u_xpb_out[22][1019],u_xpb_out[23][1019],u_xpb_out[24][1019],u_xpb_out[25][1019],u_xpb_out[26][1019],u_xpb_out[27][1019],u_xpb_out[28][1019],u_xpb_out[29][1019],u_xpb_out[30][1019],u_xpb_out[31][1019],u_xpb_out[32][1019],u_xpb_out[33][1019],u_xpb_out[34][1019],u_xpb_out[35][1019],u_xpb_out[36][1019],u_xpb_out[37][1019],u_xpb_out[38][1019],u_xpb_out[39][1019],u_xpb_out[40][1019],u_xpb_out[41][1019],u_xpb_out[42][1019],u_xpb_out[43][1019],u_xpb_out[44][1019],u_xpb_out[45][1019],u_xpb_out[46][1019],u_xpb_out[47][1019],u_xpb_out[48][1019],u_xpb_out[49][1019],u_xpb_out[50][1019],u_xpb_out[51][1019],u_xpb_out[52][1019],u_xpb_out[53][1019],u_xpb_out[54][1019],u_xpb_out[55][1019],u_xpb_out[56][1019],u_xpb_out[57][1019],u_xpb_out[58][1019],u_xpb_out[59][1019],u_xpb_out[60][1019],u_xpb_out[61][1019],u_xpb_out[62][1019],u_xpb_out[63][1019],u_xpb_out[64][1019],u_xpb_out[65][1019],u_xpb_out[66][1019],u_xpb_out[67][1019],u_xpb_out[68][1019],u_xpb_out[69][1019],u_xpb_out[70][1019],u_xpb_out[71][1019],u_xpb_out[72][1019],u_xpb_out[73][1019],u_xpb_out[74][1019],u_xpb_out[75][1019],u_xpb_out[76][1019],u_xpb_out[77][1019],u_xpb_out[78][1019],u_xpb_out[79][1019],u_xpb_out[80][1019],u_xpb_out[81][1019],u_xpb_out[82][1019],u_xpb_out[83][1019],u_xpb_out[84][1019],u_xpb_out[85][1019],u_xpb_out[86][1019],u_xpb_out[87][1019],u_xpb_out[88][1019],u_xpb_out[89][1019],u_xpb_out[90][1019],u_xpb_out[91][1019],u_xpb_out[92][1019],u_xpb_out[93][1019],u_xpb_out[94][1019],u_xpb_out[95][1019],u_xpb_out[96][1019],u_xpb_out[97][1019],u_xpb_out[98][1019],u_xpb_out[99][1019],u_xpb_out[100][1019],u_xpb_out[101][1019],u_xpb_out[102][1019],u_xpb_out[103][1019],u_xpb_out[104][1019],u_xpb_out[105][1019]};

assign col_out_1020 = {u_xpb_out[0][1020],u_xpb_out[1][1020],u_xpb_out[2][1020],u_xpb_out[3][1020],u_xpb_out[4][1020],u_xpb_out[5][1020],u_xpb_out[6][1020],u_xpb_out[7][1020],u_xpb_out[8][1020],u_xpb_out[9][1020],u_xpb_out[10][1020],u_xpb_out[11][1020],u_xpb_out[12][1020],u_xpb_out[13][1020],u_xpb_out[14][1020],u_xpb_out[15][1020],u_xpb_out[16][1020],u_xpb_out[17][1020],u_xpb_out[18][1020],u_xpb_out[19][1020],u_xpb_out[20][1020],u_xpb_out[21][1020],u_xpb_out[22][1020],u_xpb_out[23][1020],u_xpb_out[24][1020],u_xpb_out[25][1020],u_xpb_out[26][1020],u_xpb_out[27][1020],u_xpb_out[28][1020],u_xpb_out[29][1020],u_xpb_out[30][1020],u_xpb_out[31][1020],u_xpb_out[32][1020],u_xpb_out[33][1020],u_xpb_out[34][1020],u_xpb_out[35][1020],u_xpb_out[36][1020],u_xpb_out[37][1020],u_xpb_out[38][1020],u_xpb_out[39][1020],u_xpb_out[40][1020],u_xpb_out[41][1020],u_xpb_out[42][1020],u_xpb_out[43][1020],u_xpb_out[44][1020],u_xpb_out[45][1020],u_xpb_out[46][1020],u_xpb_out[47][1020],u_xpb_out[48][1020],u_xpb_out[49][1020],u_xpb_out[50][1020],u_xpb_out[51][1020],u_xpb_out[52][1020],u_xpb_out[53][1020],u_xpb_out[54][1020],u_xpb_out[55][1020],u_xpb_out[56][1020],u_xpb_out[57][1020],u_xpb_out[58][1020],u_xpb_out[59][1020],u_xpb_out[60][1020],u_xpb_out[61][1020],u_xpb_out[62][1020],u_xpb_out[63][1020],u_xpb_out[64][1020],u_xpb_out[65][1020],u_xpb_out[66][1020],u_xpb_out[67][1020],u_xpb_out[68][1020],u_xpb_out[69][1020],u_xpb_out[70][1020],u_xpb_out[71][1020],u_xpb_out[72][1020],u_xpb_out[73][1020],u_xpb_out[74][1020],u_xpb_out[75][1020],u_xpb_out[76][1020],u_xpb_out[77][1020],u_xpb_out[78][1020],u_xpb_out[79][1020],u_xpb_out[80][1020],u_xpb_out[81][1020],u_xpb_out[82][1020],u_xpb_out[83][1020],u_xpb_out[84][1020],u_xpb_out[85][1020],u_xpb_out[86][1020],u_xpb_out[87][1020],u_xpb_out[88][1020],u_xpb_out[89][1020],u_xpb_out[90][1020],u_xpb_out[91][1020],u_xpb_out[92][1020],u_xpb_out[93][1020],u_xpb_out[94][1020],u_xpb_out[95][1020],u_xpb_out[96][1020],u_xpb_out[97][1020],u_xpb_out[98][1020],u_xpb_out[99][1020],u_xpb_out[100][1020],u_xpb_out[101][1020],u_xpb_out[102][1020],u_xpb_out[103][1020],u_xpb_out[104][1020],u_xpb_out[105][1020]};

assign col_out_1021 = {u_xpb_out[0][1021],u_xpb_out[1][1021],u_xpb_out[2][1021],u_xpb_out[3][1021],u_xpb_out[4][1021],u_xpb_out[5][1021],u_xpb_out[6][1021],u_xpb_out[7][1021],u_xpb_out[8][1021],u_xpb_out[9][1021],u_xpb_out[10][1021],u_xpb_out[11][1021],u_xpb_out[12][1021],u_xpb_out[13][1021],u_xpb_out[14][1021],u_xpb_out[15][1021],u_xpb_out[16][1021],u_xpb_out[17][1021],u_xpb_out[18][1021],u_xpb_out[19][1021],u_xpb_out[20][1021],u_xpb_out[21][1021],u_xpb_out[22][1021],u_xpb_out[23][1021],u_xpb_out[24][1021],u_xpb_out[25][1021],u_xpb_out[26][1021],u_xpb_out[27][1021],u_xpb_out[28][1021],u_xpb_out[29][1021],u_xpb_out[30][1021],u_xpb_out[31][1021],u_xpb_out[32][1021],u_xpb_out[33][1021],u_xpb_out[34][1021],u_xpb_out[35][1021],u_xpb_out[36][1021],u_xpb_out[37][1021],u_xpb_out[38][1021],u_xpb_out[39][1021],u_xpb_out[40][1021],u_xpb_out[41][1021],u_xpb_out[42][1021],u_xpb_out[43][1021],u_xpb_out[44][1021],u_xpb_out[45][1021],u_xpb_out[46][1021],u_xpb_out[47][1021],u_xpb_out[48][1021],u_xpb_out[49][1021],u_xpb_out[50][1021],u_xpb_out[51][1021],u_xpb_out[52][1021],u_xpb_out[53][1021],u_xpb_out[54][1021],u_xpb_out[55][1021],u_xpb_out[56][1021],u_xpb_out[57][1021],u_xpb_out[58][1021],u_xpb_out[59][1021],u_xpb_out[60][1021],u_xpb_out[61][1021],u_xpb_out[62][1021],u_xpb_out[63][1021],u_xpb_out[64][1021],u_xpb_out[65][1021],u_xpb_out[66][1021],u_xpb_out[67][1021],u_xpb_out[68][1021],u_xpb_out[69][1021],u_xpb_out[70][1021],u_xpb_out[71][1021],u_xpb_out[72][1021],u_xpb_out[73][1021],u_xpb_out[74][1021],u_xpb_out[75][1021],u_xpb_out[76][1021],u_xpb_out[77][1021],u_xpb_out[78][1021],u_xpb_out[79][1021],u_xpb_out[80][1021],u_xpb_out[81][1021],u_xpb_out[82][1021],u_xpb_out[83][1021],u_xpb_out[84][1021],u_xpb_out[85][1021],u_xpb_out[86][1021],u_xpb_out[87][1021],u_xpb_out[88][1021],u_xpb_out[89][1021],u_xpb_out[90][1021],u_xpb_out[91][1021],u_xpb_out[92][1021],u_xpb_out[93][1021],u_xpb_out[94][1021],u_xpb_out[95][1021],u_xpb_out[96][1021],u_xpb_out[97][1021],u_xpb_out[98][1021],u_xpb_out[99][1021],u_xpb_out[100][1021],u_xpb_out[101][1021],u_xpb_out[102][1021],u_xpb_out[103][1021],u_xpb_out[104][1021],u_xpb_out[105][1021]};

assign col_out_1022 = {u_xpb_out[0][1022],u_xpb_out[1][1022],u_xpb_out[2][1022],u_xpb_out[3][1022],u_xpb_out[4][1022],u_xpb_out[5][1022],u_xpb_out[6][1022],u_xpb_out[7][1022],u_xpb_out[8][1022],u_xpb_out[9][1022],u_xpb_out[10][1022],u_xpb_out[11][1022],u_xpb_out[12][1022],u_xpb_out[13][1022],u_xpb_out[14][1022],u_xpb_out[15][1022],u_xpb_out[16][1022],u_xpb_out[17][1022],u_xpb_out[18][1022],u_xpb_out[19][1022],u_xpb_out[20][1022],u_xpb_out[21][1022],u_xpb_out[22][1022],u_xpb_out[23][1022],u_xpb_out[24][1022],u_xpb_out[25][1022],u_xpb_out[26][1022],u_xpb_out[27][1022],u_xpb_out[28][1022],u_xpb_out[29][1022],u_xpb_out[30][1022],u_xpb_out[31][1022],u_xpb_out[32][1022],u_xpb_out[33][1022],u_xpb_out[34][1022],u_xpb_out[35][1022],u_xpb_out[36][1022],u_xpb_out[37][1022],u_xpb_out[38][1022],u_xpb_out[39][1022],u_xpb_out[40][1022],u_xpb_out[41][1022],u_xpb_out[42][1022],u_xpb_out[43][1022],u_xpb_out[44][1022],u_xpb_out[45][1022],u_xpb_out[46][1022],u_xpb_out[47][1022],u_xpb_out[48][1022],u_xpb_out[49][1022],u_xpb_out[50][1022],u_xpb_out[51][1022],u_xpb_out[52][1022],u_xpb_out[53][1022],u_xpb_out[54][1022],u_xpb_out[55][1022],u_xpb_out[56][1022],u_xpb_out[57][1022],u_xpb_out[58][1022],u_xpb_out[59][1022],u_xpb_out[60][1022],u_xpb_out[61][1022],u_xpb_out[62][1022],u_xpb_out[63][1022],u_xpb_out[64][1022],u_xpb_out[65][1022],u_xpb_out[66][1022],u_xpb_out[67][1022],u_xpb_out[68][1022],u_xpb_out[69][1022],u_xpb_out[70][1022],u_xpb_out[71][1022],u_xpb_out[72][1022],u_xpb_out[73][1022],u_xpb_out[74][1022],u_xpb_out[75][1022],u_xpb_out[76][1022],u_xpb_out[77][1022],u_xpb_out[78][1022],u_xpb_out[79][1022],u_xpb_out[80][1022],u_xpb_out[81][1022],u_xpb_out[82][1022],u_xpb_out[83][1022],u_xpb_out[84][1022],u_xpb_out[85][1022],u_xpb_out[86][1022],u_xpb_out[87][1022],u_xpb_out[88][1022],u_xpb_out[89][1022],u_xpb_out[90][1022],u_xpb_out[91][1022],u_xpb_out[92][1022],u_xpb_out[93][1022],u_xpb_out[94][1022],u_xpb_out[95][1022],u_xpb_out[96][1022],u_xpb_out[97][1022],u_xpb_out[98][1022],u_xpb_out[99][1022],u_xpb_out[100][1022],u_xpb_out[101][1022],u_xpb_out[102][1022],u_xpb_out[103][1022],u_xpb_out[104][1022],u_xpb_out[105][1022]};

assign col_out_1023 = {u_xpb_out[0][1023],u_xpb_out[1][1023],u_xpb_out[2][1023],u_xpb_out[3][1023],u_xpb_out[4][1023],u_xpb_out[5][1023],u_xpb_out[6][1023],u_xpb_out[7][1023],u_xpb_out[8][1023],u_xpb_out[9][1023],u_xpb_out[10][1023],u_xpb_out[11][1023],u_xpb_out[12][1023],u_xpb_out[13][1023],u_xpb_out[14][1023],u_xpb_out[15][1023],u_xpb_out[16][1023],u_xpb_out[17][1023],u_xpb_out[18][1023],u_xpb_out[19][1023],u_xpb_out[20][1023],u_xpb_out[21][1023],u_xpb_out[22][1023],u_xpb_out[23][1023],u_xpb_out[24][1023],u_xpb_out[25][1023],u_xpb_out[26][1023],u_xpb_out[27][1023],u_xpb_out[28][1023],u_xpb_out[29][1023],u_xpb_out[30][1023],u_xpb_out[31][1023],u_xpb_out[32][1023],u_xpb_out[33][1023],u_xpb_out[34][1023],u_xpb_out[35][1023],u_xpb_out[36][1023],u_xpb_out[37][1023],u_xpb_out[38][1023],u_xpb_out[39][1023],u_xpb_out[40][1023],u_xpb_out[41][1023],u_xpb_out[42][1023],u_xpb_out[43][1023],u_xpb_out[44][1023],u_xpb_out[45][1023],u_xpb_out[46][1023],u_xpb_out[47][1023],u_xpb_out[48][1023],u_xpb_out[49][1023],u_xpb_out[50][1023],u_xpb_out[51][1023],u_xpb_out[52][1023],u_xpb_out[53][1023],u_xpb_out[54][1023],u_xpb_out[55][1023],u_xpb_out[56][1023],u_xpb_out[57][1023],u_xpb_out[58][1023],u_xpb_out[59][1023],u_xpb_out[60][1023],u_xpb_out[61][1023],u_xpb_out[62][1023],u_xpb_out[63][1023],u_xpb_out[64][1023],u_xpb_out[65][1023],u_xpb_out[66][1023],u_xpb_out[67][1023],u_xpb_out[68][1023],u_xpb_out[69][1023],u_xpb_out[70][1023],u_xpb_out[71][1023],u_xpb_out[72][1023],u_xpb_out[73][1023],u_xpb_out[74][1023],u_xpb_out[75][1023],u_xpb_out[76][1023],u_xpb_out[77][1023],u_xpb_out[78][1023],u_xpb_out[79][1023],u_xpb_out[80][1023],u_xpb_out[81][1023],u_xpb_out[82][1023],u_xpb_out[83][1023],u_xpb_out[84][1023],u_xpb_out[85][1023],u_xpb_out[86][1023],u_xpb_out[87][1023],u_xpb_out[88][1023],u_xpb_out[89][1023],u_xpb_out[90][1023],u_xpb_out[91][1023],u_xpb_out[92][1023],u_xpb_out[93][1023],u_xpb_out[94][1023],u_xpb_out[95][1023],u_xpb_out[96][1023],u_xpb_out[97][1023],u_xpb_out[98][1023],u_xpb_out[99][1023],u_xpb_out[100][1023],u_xpb_out[101][1023],u_xpb_out[102][1023],u_xpb_out[103][1023],u_xpb_out[104][1023],u_xpb_out[105][1023]};



endmodule



module compressor_array_152_48_1027
(
    input  [151:0] col_in_0,
    input  [151:0] col_in_1,
    input  [151:0] col_in_2,
    input  [151:0] col_in_3,
    input  [151:0] col_in_4,
    input  [151:0] col_in_5,
    input  [151:0] col_in_6,
    input  [151:0] col_in_7,
    input  [151:0] col_in_8,
    input  [151:0] col_in_9,
    input  [151:0] col_in_10,
    input  [151:0] col_in_11,
    input  [151:0] col_in_12,
    input  [151:0] col_in_13,
    input  [151:0] col_in_14,
    input  [151:0] col_in_15,
    input  [151:0] col_in_16,
    input  [151:0] col_in_17,
    input  [151:0] col_in_18,
    input  [151:0] col_in_19,
    input  [151:0] col_in_20,
    input  [151:0] col_in_21,
    input  [151:0] col_in_22,
    input  [151:0] col_in_23,
    input  [151:0] col_in_24,
    input  [151:0] col_in_25,
    input  [151:0] col_in_26,
    input  [151:0] col_in_27,
    input  [151:0] col_in_28,
    input  [151:0] col_in_29,
    input  [151:0] col_in_30,
    input  [151:0] col_in_31,
    input  [151:0] col_in_32,
    input  [151:0] col_in_33,
    input  [151:0] col_in_34,
    input  [151:0] col_in_35,
    input  [151:0] col_in_36,
    input  [151:0] col_in_37,
    input  [151:0] col_in_38,
    input  [151:0] col_in_39,
    input  [151:0] col_in_40,
    input  [151:0] col_in_41,
    input  [151:0] col_in_42,
    input  [151:0] col_in_43,
    input  [151:0] col_in_44,
    input  [151:0] col_in_45,
    input  [151:0] col_in_46,
    input  [151:0] col_in_47,
    input  [151:0] col_in_48,
    input  [151:0] col_in_49,
    input  [151:0] col_in_50,
    input  [151:0] col_in_51,
    input  [151:0] col_in_52,
    input  [151:0] col_in_53,
    input  [151:0] col_in_54,
    input  [151:0] col_in_55,
    input  [151:0] col_in_56,
    input  [151:0] col_in_57,
    input  [151:0] col_in_58,
    input  [151:0] col_in_59,
    input  [151:0] col_in_60,
    input  [151:0] col_in_61,
    input  [151:0] col_in_62,
    input  [151:0] col_in_63,
    input  [151:0] col_in_64,
    input  [151:0] col_in_65,
    input  [151:0] col_in_66,
    input  [151:0] col_in_67,
    input  [151:0] col_in_68,
    input  [151:0] col_in_69,
    input  [151:0] col_in_70,
    input  [151:0] col_in_71,
    input  [151:0] col_in_72,
    input  [151:0] col_in_73,
    input  [151:0] col_in_74,
    input  [151:0] col_in_75,
    input  [151:0] col_in_76,
    input  [151:0] col_in_77,
    input  [151:0] col_in_78,
    input  [151:0] col_in_79,
    input  [151:0] col_in_80,
    input  [151:0] col_in_81,
    input  [151:0] col_in_82,
    input  [151:0] col_in_83,
    input  [151:0] col_in_84,
    input  [151:0] col_in_85,
    input  [151:0] col_in_86,
    input  [151:0] col_in_87,
    input  [151:0] col_in_88,
    input  [151:0] col_in_89,
    input  [151:0] col_in_90,
    input  [151:0] col_in_91,
    input  [151:0] col_in_92,
    input  [151:0] col_in_93,
    input  [151:0] col_in_94,
    input  [151:0] col_in_95,
    input  [151:0] col_in_96,
    input  [151:0] col_in_97,
    input  [151:0] col_in_98,
    input  [151:0] col_in_99,
    input  [151:0] col_in_100,
    input  [151:0] col_in_101,
    input  [151:0] col_in_102,
    input  [151:0] col_in_103,
    input  [151:0] col_in_104,
    input  [151:0] col_in_105,
    input  [151:0] col_in_106,
    input  [151:0] col_in_107,
    input  [151:0] col_in_108,
    input  [151:0] col_in_109,
    input  [151:0] col_in_110,
    input  [151:0] col_in_111,
    input  [151:0] col_in_112,
    input  [151:0] col_in_113,
    input  [151:0] col_in_114,
    input  [151:0] col_in_115,
    input  [151:0] col_in_116,
    input  [151:0] col_in_117,
    input  [151:0] col_in_118,
    input  [151:0] col_in_119,
    input  [151:0] col_in_120,
    input  [151:0] col_in_121,
    input  [151:0] col_in_122,
    input  [151:0] col_in_123,
    input  [151:0] col_in_124,
    input  [151:0] col_in_125,
    input  [151:0] col_in_126,
    input  [151:0] col_in_127,
    input  [151:0] col_in_128,
    input  [151:0] col_in_129,
    input  [151:0] col_in_130,
    input  [151:0] col_in_131,
    input  [151:0] col_in_132,
    input  [151:0] col_in_133,
    input  [151:0] col_in_134,
    input  [151:0] col_in_135,
    input  [151:0] col_in_136,
    input  [151:0] col_in_137,
    input  [151:0] col_in_138,
    input  [151:0] col_in_139,
    input  [151:0] col_in_140,
    input  [151:0] col_in_141,
    input  [151:0] col_in_142,
    input  [151:0] col_in_143,
    input  [151:0] col_in_144,
    input  [151:0] col_in_145,
    input  [151:0] col_in_146,
    input  [151:0] col_in_147,
    input  [151:0] col_in_148,
    input  [151:0] col_in_149,
    input  [151:0] col_in_150,
    input  [151:0] col_in_151,
    input  [151:0] col_in_152,
    input  [151:0] col_in_153,
    input  [151:0] col_in_154,
    input  [151:0] col_in_155,
    input  [151:0] col_in_156,
    input  [151:0] col_in_157,
    input  [151:0] col_in_158,
    input  [151:0] col_in_159,
    input  [151:0] col_in_160,
    input  [151:0] col_in_161,
    input  [151:0] col_in_162,
    input  [151:0] col_in_163,
    input  [151:0] col_in_164,
    input  [151:0] col_in_165,
    input  [151:0] col_in_166,
    input  [151:0] col_in_167,
    input  [151:0] col_in_168,
    input  [151:0] col_in_169,
    input  [151:0] col_in_170,
    input  [151:0] col_in_171,
    input  [151:0] col_in_172,
    input  [151:0] col_in_173,
    input  [151:0] col_in_174,
    input  [151:0] col_in_175,
    input  [151:0] col_in_176,
    input  [151:0] col_in_177,
    input  [151:0] col_in_178,
    input  [151:0] col_in_179,
    input  [151:0] col_in_180,
    input  [151:0] col_in_181,
    input  [151:0] col_in_182,
    input  [151:0] col_in_183,
    input  [151:0] col_in_184,
    input  [151:0] col_in_185,
    input  [151:0] col_in_186,
    input  [151:0] col_in_187,
    input  [151:0] col_in_188,
    input  [151:0] col_in_189,
    input  [151:0] col_in_190,
    input  [151:0] col_in_191,
    input  [151:0] col_in_192,
    input  [151:0] col_in_193,
    input  [151:0] col_in_194,
    input  [151:0] col_in_195,
    input  [151:0] col_in_196,
    input  [151:0] col_in_197,
    input  [151:0] col_in_198,
    input  [151:0] col_in_199,
    input  [151:0] col_in_200,
    input  [151:0] col_in_201,
    input  [151:0] col_in_202,
    input  [151:0] col_in_203,
    input  [151:0] col_in_204,
    input  [151:0] col_in_205,
    input  [151:0] col_in_206,
    input  [151:0] col_in_207,
    input  [151:0] col_in_208,
    input  [151:0] col_in_209,
    input  [151:0] col_in_210,
    input  [151:0] col_in_211,
    input  [151:0] col_in_212,
    input  [151:0] col_in_213,
    input  [151:0] col_in_214,
    input  [151:0] col_in_215,
    input  [151:0] col_in_216,
    input  [151:0] col_in_217,
    input  [151:0] col_in_218,
    input  [151:0] col_in_219,
    input  [151:0] col_in_220,
    input  [151:0] col_in_221,
    input  [151:0] col_in_222,
    input  [151:0] col_in_223,
    input  [151:0] col_in_224,
    input  [151:0] col_in_225,
    input  [151:0] col_in_226,
    input  [151:0] col_in_227,
    input  [151:0] col_in_228,
    input  [151:0] col_in_229,
    input  [151:0] col_in_230,
    input  [151:0] col_in_231,
    input  [151:0] col_in_232,
    input  [151:0] col_in_233,
    input  [151:0] col_in_234,
    input  [151:0] col_in_235,
    input  [151:0] col_in_236,
    input  [151:0] col_in_237,
    input  [151:0] col_in_238,
    input  [151:0] col_in_239,
    input  [151:0] col_in_240,
    input  [151:0] col_in_241,
    input  [151:0] col_in_242,
    input  [151:0] col_in_243,
    input  [151:0] col_in_244,
    input  [151:0] col_in_245,
    input  [151:0] col_in_246,
    input  [151:0] col_in_247,
    input  [151:0] col_in_248,
    input  [151:0] col_in_249,
    input  [151:0] col_in_250,
    input  [151:0] col_in_251,
    input  [151:0] col_in_252,
    input  [151:0] col_in_253,
    input  [151:0] col_in_254,
    input  [151:0] col_in_255,
    input  [151:0] col_in_256,
    input  [151:0] col_in_257,
    input  [151:0] col_in_258,
    input  [151:0] col_in_259,
    input  [151:0] col_in_260,
    input  [151:0] col_in_261,
    input  [151:0] col_in_262,
    input  [151:0] col_in_263,
    input  [151:0] col_in_264,
    input  [151:0] col_in_265,
    input  [151:0] col_in_266,
    input  [151:0] col_in_267,
    input  [151:0] col_in_268,
    input  [151:0] col_in_269,
    input  [151:0] col_in_270,
    input  [151:0] col_in_271,
    input  [151:0] col_in_272,
    input  [151:0] col_in_273,
    input  [151:0] col_in_274,
    input  [151:0] col_in_275,
    input  [151:0] col_in_276,
    input  [151:0] col_in_277,
    input  [151:0] col_in_278,
    input  [151:0] col_in_279,
    input  [151:0] col_in_280,
    input  [151:0] col_in_281,
    input  [151:0] col_in_282,
    input  [151:0] col_in_283,
    input  [151:0] col_in_284,
    input  [151:0] col_in_285,
    input  [151:0] col_in_286,
    input  [151:0] col_in_287,
    input  [151:0] col_in_288,
    input  [151:0] col_in_289,
    input  [151:0] col_in_290,
    input  [151:0] col_in_291,
    input  [151:0] col_in_292,
    input  [151:0] col_in_293,
    input  [151:0] col_in_294,
    input  [151:0] col_in_295,
    input  [151:0] col_in_296,
    input  [151:0] col_in_297,
    input  [151:0] col_in_298,
    input  [151:0] col_in_299,
    input  [151:0] col_in_300,
    input  [151:0] col_in_301,
    input  [151:0] col_in_302,
    input  [151:0] col_in_303,
    input  [151:0] col_in_304,
    input  [151:0] col_in_305,
    input  [151:0] col_in_306,
    input  [151:0] col_in_307,
    input  [151:0] col_in_308,
    input  [151:0] col_in_309,
    input  [151:0] col_in_310,
    input  [151:0] col_in_311,
    input  [151:0] col_in_312,
    input  [151:0] col_in_313,
    input  [151:0] col_in_314,
    input  [151:0] col_in_315,
    input  [151:0] col_in_316,
    input  [151:0] col_in_317,
    input  [151:0] col_in_318,
    input  [151:0] col_in_319,
    input  [151:0] col_in_320,
    input  [151:0] col_in_321,
    input  [151:0] col_in_322,
    input  [151:0] col_in_323,
    input  [151:0] col_in_324,
    input  [151:0] col_in_325,
    input  [151:0] col_in_326,
    input  [151:0] col_in_327,
    input  [151:0] col_in_328,
    input  [151:0] col_in_329,
    input  [151:0] col_in_330,
    input  [151:0] col_in_331,
    input  [151:0] col_in_332,
    input  [151:0] col_in_333,
    input  [151:0] col_in_334,
    input  [151:0] col_in_335,
    input  [151:0] col_in_336,
    input  [151:0] col_in_337,
    input  [151:0] col_in_338,
    input  [151:0] col_in_339,
    input  [151:0] col_in_340,
    input  [151:0] col_in_341,
    input  [151:0] col_in_342,
    input  [151:0] col_in_343,
    input  [151:0] col_in_344,
    input  [151:0] col_in_345,
    input  [151:0] col_in_346,
    input  [151:0] col_in_347,
    input  [151:0] col_in_348,
    input  [151:0] col_in_349,
    input  [151:0] col_in_350,
    input  [151:0] col_in_351,
    input  [151:0] col_in_352,
    input  [151:0] col_in_353,
    input  [151:0] col_in_354,
    input  [151:0] col_in_355,
    input  [151:0] col_in_356,
    input  [151:0] col_in_357,
    input  [151:0] col_in_358,
    input  [151:0] col_in_359,
    input  [151:0] col_in_360,
    input  [151:0] col_in_361,
    input  [151:0] col_in_362,
    input  [151:0] col_in_363,
    input  [151:0] col_in_364,
    input  [151:0] col_in_365,
    input  [151:0] col_in_366,
    input  [151:0] col_in_367,
    input  [151:0] col_in_368,
    input  [151:0] col_in_369,
    input  [151:0] col_in_370,
    input  [151:0] col_in_371,
    input  [151:0] col_in_372,
    input  [151:0] col_in_373,
    input  [151:0] col_in_374,
    input  [151:0] col_in_375,
    input  [151:0] col_in_376,
    input  [151:0] col_in_377,
    input  [151:0] col_in_378,
    input  [151:0] col_in_379,
    input  [151:0] col_in_380,
    input  [151:0] col_in_381,
    input  [151:0] col_in_382,
    input  [151:0] col_in_383,
    input  [151:0] col_in_384,
    input  [151:0] col_in_385,
    input  [151:0] col_in_386,
    input  [151:0] col_in_387,
    input  [151:0] col_in_388,
    input  [151:0] col_in_389,
    input  [151:0] col_in_390,
    input  [151:0] col_in_391,
    input  [151:0] col_in_392,
    input  [151:0] col_in_393,
    input  [151:0] col_in_394,
    input  [151:0] col_in_395,
    input  [151:0] col_in_396,
    input  [151:0] col_in_397,
    input  [151:0] col_in_398,
    input  [151:0] col_in_399,
    input  [151:0] col_in_400,
    input  [151:0] col_in_401,
    input  [151:0] col_in_402,
    input  [151:0] col_in_403,
    input  [151:0] col_in_404,
    input  [151:0] col_in_405,
    input  [151:0] col_in_406,
    input  [151:0] col_in_407,
    input  [151:0] col_in_408,
    input  [151:0] col_in_409,
    input  [151:0] col_in_410,
    input  [151:0] col_in_411,
    input  [151:0] col_in_412,
    input  [151:0] col_in_413,
    input  [151:0] col_in_414,
    input  [151:0] col_in_415,
    input  [151:0] col_in_416,
    input  [151:0] col_in_417,
    input  [151:0] col_in_418,
    input  [151:0] col_in_419,
    input  [151:0] col_in_420,
    input  [151:0] col_in_421,
    input  [151:0] col_in_422,
    input  [151:0] col_in_423,
    input  [151:0] col_in_424,
    input  [151:0] col_in_425,
    input  [151:0] col_in_426,
    input  [151:0] col_in_427,
    input  [151:0] col_in_428,
    input  [151:0] col_in_429,
    input  [151:0] col_in_430,
    input  [151:0] col_in_431,
    input  [151:0] col_in_432,
    input  [151:0] col_in_433,
    input  [151:0] col_in_434,
    input  [151:0] col_in_435,
    input  [151:0] col_in_436,
    input  [151:0] col_in_437,
    input  [151:0] col_in_438,
    input  [151:0] col_in_439,
    input  [151:0] col_in_440,
    input  [151:0] col_in_441,
    input  [151:0] col_in_442,
    input  [151:0] col_in_443,
    input  [151:0] col_in_444,
    input  [151:0] col_in_445,
    input  [151:0] col_in_446,
    input  [151:0] col_in_447,
    input  [151:0] col_in_448,
    input  [151:0] col_in_449,
    input  [151:0] col_in_450,
    input  [151:0] col_in_451,
    input  [151:0] col_in_452,
    input  [151:0] col_in_453,
    input  [151:0] col_in_454,
    input  [151:0] col_in_455,
    input  [151:0] col_in_456,
    input  [151:0] col_in_457,
    input  [151:0] col_in_458,
    input  [151:0] col_in_459,
    input  [151:0] col_in_460,
    input  [151:0] col_in_461,
    input  [151:0] col_in_462,
    input  [151:0] col_in_463,
    input  [151:0] col_in_464,
    input  [151:0] col_in_465,
    input  [151:0] col_in_466,
    input  [151:0] col_in_467,
    input  [151:0] col_in_468,
    input  [151:0] col_in_469,
    input  [151:0] col_in_470,
    input  [151:0] col_in_471,
    input  [151:0] col_in_472,
    input  [151:0] col_in_473,
    input  [151:0] col_in_474,
    input  [151:0] col_in_475,
    input  [151:0] col_in_476,
    input  [151:0] col_in_477,
    input  [151:0] col_in_478,
    input  [151:0] col_in_479,
    input  [151:0] col_in_480,
    input  [151:0] col_in_481,
    input  [151:0] col_in_482,
    input  [151:0] col_in_483,
    input  [151:0] col_in_484,
    input  [151:0] col_in_485,
    input  [151:0] col_in_486,
    input  [151:0] col_in_487,
    input  [151:0] col_in_488,
    input  [151:0] col_in_489,
    input  [151:0] col_in_490,
    input  [151:0] col_in_491,
    input  [151:0] col_in_492,
    input  [151:0] col_in_493,
    input  [151:0] col_in_494,
    input  [151:0] col_in_495,
    input  [151:0] col_in_496,
    input  [151:0] col_in_497,
    input  [151:0] col_in_498,
    input  [151:0] col_in_499,
    input  [151:0] col_in_500,
    input  [151:0] col_in_501,
    input  [151:0] col_in_502,
    input  [151:0] col_in_503,
    input  [151:0] col_in_504,
    input  [151:0] col_in_505,
    input  [151:0] col_in_506,
    input  [151:0] col_in_507,
    input  [151:0] col_in_508,
    input  [151:0] col_in_509,
    input  [151:0] col_in_510,
    input  [151:0] col_in_511,
    input  [151:0] col_in_512,
    input  [151:0] col_in_513,
    input  [151:0] col_in_514,
    input  [151:0] col_in_515,
    input  [151:0] col_in_516,
    input  [151:0] col_in_517,
    input  [151:0] col_in_518,
    input  [151:0] col_in_519,
    input  [151:0] col_in_520,
    input  [151:0] col_in_521,
    input  [151:0] col_in_522,
    input  [151:0] col_in_523,
    input  [151:0] col_in_524,
    input  [151:0] col_in_525,
    input  [151:0] col_in_526,
    input  [151:0] col_in_527,
    input  [151:0] col_in_528,
    input  [151:0] col_in_529,
    input  [151:0] col_in_530,
    input  [151:0] col_in_531,
    input  [151:0] col_in_532,
    input  [151:0] col_in_533,
    input  [151:0] col_in_534,
    input  [151:0] col_in_535,
    input  [151:0] col_in_536,
    input  [151:0] col_in_537,
    input  [151:0] col_in_538,
    input  [151:0] col_in_539,
    input  [151:0] col_in_540,
    input  [151:0] col_in_541,
    input  [151:0] col_in_542,
    input  [151:0] col_in_543,
    input  [151:0] col_in_544,
    input  [151:0] col_in_545,
    input  [151:0] col_in_546,
    input  [151:0] col_in_547,
    input  [151:0] col_in_548,
    input  [151:0] col_in_549,
    input  [151:0] col_in_550,
    input  [151:0] col_in_551,
    input  [151:0] col_in_552,
    input  [151:0] col_in_553,
    input  [151:0] col_in_554,
    input  [151:0] col_in_555,
    input  [151:0] col_in_556,
    input  [151:0] col_in_557,
    input  [151:0] col_in_558,
    input  [151:0] col_in_559,
    input  [151:0] col_in_560,
    input  [151:0] col_in_561,
    input  [151:0] col_in_562,
    input  [151:0] col_in_563,
    input  [151:0] col_in_564,
    input  [151:0] col_in_565,
    input  [151:0] col_in_566,
    input  [151:0] col_in_567,
    input  [151:0] col_in_568,
    input  [151:0] col_in_569,
    input  [151:0] col_in_570,
    input  [151:0] col_in_571,
    input  [151:0] col_in_572,
    input  [151:0] col_in_573,
    input  [151:0] col_in_574,
    input  [151:0] col_in_575,
    input  [151:0] col_in_576,
    input  [151:0] col_in_577,
    input  [151:0] col_in_578,
    input  [151:0] col_in_579,
    input  [151:0] col_in_580,
    input  [151:0] col_in_581,
    input  [151:0] col_in_582,
    input  [151:0] col_in_583,
    input  [151:0] col_in_584,
    input  [151:0] col_in_585,
    input  [151:0] col_in_586,
    input  [151:0] col_in_587,
    input  [151:0] col_in_588,
    input  [151:0] col_in_589,
    input  [151:0] col_in_590,
    input  [151:0] col_in_591,
    input  [151:0] col_in_592,
    input  [151:0] col_in_593,
    input  [151:0] col_in_594,
    input  [151:0] col_in_595,
    input  [151:0] col_in_596,
    input  [151:0] col_in_597,
    input  [151:0] col_in_598,
    input  [151:0] col_in_599,
    input  [151:0] col_in_600,
    input  [151:0] col_in_601,
    input  [151:0] col_in_602,
    input  [151:0] col_in_603,
    input  [151:0] col_in_604,
    input  [151:0] col_in_605,
    input  [151:0] col_in_606,
    input  [151:0] col_in_607,
    input  [151:0] col_in_608,
    input  [151:0] col_in_609,
    input  [151:0] col_in_610,
    input  [151:0] col_in_611,
    input  [151:0] col_in_612,
    input  [151:0] col_in_613,
    input  [151:0] col_in_614,
    input  [151:0] col_in_615,
    input  [151:0] col_in_616,
    input  [151:0] col_in_617,
    input  [151:0] col_in_618,
    input  [151:0] col_in_619,
    input  [151:0] col_in_620,
    input  [151:0] col_in_621,
    input  [151:0] col_in_622,
    input  [151:0] col_in_623,
    input  [151:0] col_in_624,
    input  [151:0] col_in_625,
    input  [151:0] col_in_626,
    input  [151:0] col_in_627,
    input  [151:0] col_in_628,
    input  [151:0] col_in_629,
    input  [151:0] col_in_630,
    input  [151:0] col_in_631,
    input  [151:0] col_in_632,
    input  [151:0] col_in_633,
    input  [151:0] col_in_634,
    input  [151:0] col_in_635,
    input  [151:0] col_in_636,
    input  [151:0] col_in_637,
    input  [151:0] col_in_638,
    input  [151:0] col_in_639,
    input  [151:0] col_in_640,
    input  [151:0] col_in_641,
    input  [151:0] col_in_642,
    input  [151:0] col_in_643,
    input  [151:0] col_in_644,
    input  [151:0] col_in_645,
    input  [151:0] col_in_646,
    input  [151:0] col_in_647,
    input  [151:0] col_in_648,
    input  [151:0] col_in_649,
    input  [151:0] col_in_650,
    input  [151:0] col_in_651,
    input  [151:0] col_in_652,
    input  [151:0] col_in_653,
    input  [151:0] col_in_654,
    input  [151:0] col_in_655,
    input  [151:0] col_in_656,
    input  [151:0] col_in_657,
    input  [151:0] col_in_658,
    input  [151:0] col_in_659,
    input  [151:0] col_in_660,
    input  [151:0] col_in_661,
    input  [151:0] col_in_662,
    input  [151:0] col_in_663,
    input  [151:0] col_in_664,
    input  [151:0] col_in_665,
    input  [151:0] col_in_666,
    input  [151:0] col_in_667,
    input  [151:0] col_in_668,
    input  [151:0] col_in_669,
    input  [151:0] col_in_670,
    input  [151:0] col_in_671,
    input  [151:0] col_in_672,
    input  [151:0] col_in_673,
    input  [151:0] col_in_674,
    input  [151:0] col_in_675,
    input  [151:0] col_in_676,
    input  [151:0] col_in_677,
    input  [151:0] col_in_678,
    input  [151:0] col_in_679,
    input  [151:0] col_in_680,
    input  [151:0] col_in_681,
    input  [151:0] col_in_682,
    input  [151:0] col_in_683,
    input  [151:0] col_in_684,
    input  [151:0] col_in_685,
    input  [151:0] col_in_686,
    input  [151:0] col_in_687,
    input  [151:0] col_in_688,
    input  [151:0] col_in_689,
    input  [151:0] col_in_690,
    input  [151:0] col_in_691,
    input  [151:0] col_in_692,
    input  [151:0] col_in_693,
    input  [151:0] col_in_694,
    input  [151:0] col_in_695,
    input  [151:0] col_in_696,
    input  [151:0] col_in_697,
    input  [151:0] col_in_698,
    input  [151:0] col_in_699,
    input  [151:0] col_in_700,
    input  [151:0] col_in_701,
    input  [151:0] col_in_702,
    input  [151:0] col_in_703,
    input  [151:0] col_in_704,
    input  [151:0] col_in_705,
    input  [151:0] col_in_706,
    input  [151:0] col_in_707,
    input  [151:0] col_in_708,
    input  [151:0] col_in_709,
    input  [151:0] col_in_710,
    input  [151:0] col_in_711,
    input  [151:0] col_in_712,
    input  [151:0] col_in_713,
    input  [151:0] col_in_714,
    input  [151:0] col_in_715,
    input  [151:0] col_in_716,
    input  [151:0] col_in_717,
    input  [151:0] col_in_718,
    input  [151:0] col_in_719,
    input  [151:0] col_in_720,
    input  [151:0] col_in_721,
    input  [151:0] col_in_722,
    input  [151:0] col_in_723,
    input  [151:0] col_in_724,
    input  [151:0] col_in_725,
    input  [151:0] col_in_726,
    input  [151:0] col_in_727,
    input  [151:0] col_in_728,
    input  [151:0] col_in_729,
    input  [151:0] col_in_730,
    input  [151:0] col_in_731,
    input  [151:0] col_in_732,
    input  [151:0] col_in_733,
    input  [151:0] col_in_734,
    input  [151:0] col_in_735,
    input  [151:0] col_in_736,
    input  [151:0] col_in_737,
    input  [151:0] col_in_738,
    input  [151:0] col_in_739,
    input  [151:0] col_in_740,
    input  [151:0] col_in_741,
    input  [151:0] col_in_742,
    input  [151:0] col_in_743,
    input  [151:0] col_in_744,
    input  [151:0] col_in_745,
    input  [151:0] col_in_746,
    input  [151:0] col_in_747,
    input  [151:0] col_in_748,
    input  [151:0] col_in_749,
    input  [151:0] col_in_750,
    input  [151:0] col_in_751,
    input  [151:0] col_in_752,
    input  [151:0] col_in_753,
    input  [151:0] col_in_754,
    input  [151:0] col_in_755,
    input  [151:0] col_in_756,
    input  [151:0] col_in_757,
    input  [151:0] col_in_758,
    input  [151:0] col_in_759,
    input  [151:0] col_in_760,
    input  [151:0] col_in_761,
    input  [151:0] col_in_762,
    input  [151:0] col_in_763,
    input  [151:0] col_in_764,
    input  [151:0] col_in_765,
    input  [151:0] col_in_766,
    input  [151:0] col_in_767,
    input  [151:0] col_in_768,
    input  [151:0] col_in_769,
    input  [151:0] col_in_770,
    input  [151:0] col_in_771,
    input  [151:0] col_in_772,
    input  [151:0] col_in_773,
    input  [151:0] col_in_774,
    input  [151:0] col_in_775,
    input  [151:0] col_in_776,
    input  [151:0] col_in_777,
    input  [151:0] col_in_778,
    input  [151:0] col_in_779,
    input  [151:0] col_in_780,
    input  [151:0] col_in_781,
    input  [151:0] col_in_782,
    input  [151:0] col_in_783,
    input  [151:0] col_in_784,
    input  [151:0] col_in_785,
    input  [151:0] col_in_786,
    input  [151:0] col_in_787,
    input  [151:0] col_in_788,
    input  [151:0] col_in_789,
    input  [151:0] col_in_790,
    input  [151:0] col_in_791,
    input  [151:0] col_in_792,
    input  [151:0] col_in_793,
    input  [151:0] col_in_794,
    input  [151:0] col_in_795,
    input  [151:0] col_in_796,
    input  [151:0] col_in_797,
    input  [151:0] col_in_798,
    input  [151:0] col_in_799,
    input  [151:0] col_in_800,
    input  [151:0] col_in_801,
    input  [151:0] col_in_802,
    input  [151:0] col_in_803,
    input  [151:0] col_in_804,
    input  [151:0] col_in_805,
    input  [151:0] col_in_806,
    input  [151:0] col_in_807,
    input  [151:0] col_in_808,
    input  [151:0] col_in_809,
    input  [151:0] col_in_810,
    input  [151:0] col_in_811,
    input  [151:0] col_in_812,
    input  [151:0] col_in_813,
    input  [151:0] col_in_814,
    input  [151:0] col_in_815,
    input  [151:0] col_in_816,
    input  [151:0] col_in_817,
    input  [151:0] col_in_818,
    input  [151:0] col_in_819,
    input  [151:0] col_in_820,
    input  [151:0] col_in_821,
    input  [151:0] col_in_822,
    input  [151:0] col_in_823,
    input  [151:0] col_in_824,
    input  [151:0] col_in_825,
    input  [151:0] col_in_826,
    input  [151:0] col_in_827,
    input  [151:0] col_in_828,
    input  [151:0] col_in_829,
    input  [151:0] col_in_830,
    input  [151:0] col_in_831,
    input  [151:0] col_in_832,
    input  [151:0] col_in_833,
    input  [151:0] col_in_834,
    input  [151:0] col_in_835,
    input  [151:0] col_in_836,
    input  [151:0] col_in_837,
    input  [151:0] col_in_838,
    input  [151:0] col_in_839,
    input  [151:0] col_in_840,
    input  [151:0] col_in_841,
    input  [151:0] col_in_842,
    input  [151:0] col_in_843,
    input  [151:0] col_in_844,
    input  [151:0] col_in_845,
    input  [151:0] col_in_846,
    input  [151:0] col_in_847,
    input  [151:0] col_in_848,
    input  [151:0] col_in_849,
    input  [151:0] col_in_850,
    input  [151:0] col_in_851,
    input  [151:0] col_in_852,
    input  [151:0] col_in_853,
    input  [151:0] col_in_854,
    input  [151:0] col_in_855,
    input  [151:0] col_in_856,
    input  [151:0] col_in_857,
    input  [151:0] col_in_858,
    input  [151:0] col_in_859,
    input  [151:0] col_in_860,
    input  [151:0] col_in_861,
    input  [151:0] col_in_862,
    input  [151:0] col_in_863,
    input  [151:0] col_in_864,
    input  [151:0] col_in_865,
    input  [151:0] col_in_866,
    input  [151:0] col_in_867,
    input  [151:0] col_in_868,
    input  [151:0] col_in_869,
    input  [151:0] col_in_870,
    input  [151:0] col_in_871,
    input  [151:0] col_in_872,
    input  [151:0] col_in_873,
    input  [151:0] col_in_874,
    input  [151:0] col_in_875,
    input  [151:0] col_in_876,
    input  [151:0] col_in_877,
    input  [151:0] col_in_878,
    input  [151:0] col_in_879,
    input  [151:0] col_in_880,
    input  [151:0] col_in_881,
    input  [151:0] col_in_882,
    input  [151:0] col_in_883,
    input  [151:0] col_in_884,
    input  [151:0] col_in_885,
    input  [151:0] col_in_886,
    input  [151:0] col_in_887,
    input  [151:0] col_in_888,
    input  [151:0] col_in_889,
    input  [151:0] col_in_890,
    input  [151:0] col_in_891,
    input  [151:0] col_in_892,
    input  [151:0] col_in_893,
    input  [151:0] col_in_894,
    input  [151:0] col_in_895,
    input  [151:0] col_in_896,
    input  [151:0] col_in_897,
    input  [151:0] col_in_898,
    input  [151:0] col_in_899,
    input  [151:0] col_in_900,
    input  [151:0] col_in_901,
    input  [151:0] col_in_902,
    input  [151:0] col_in_903,
    input  [151:0] col_in_904,
    input  [151:0] col_in_905,
    input  [151:0] col_in_906,
    input  [151:0] col_in_907,
    input  [151:0] col_in_908,
    input  [151:0] col_in_909,
    input  [151:0] col_in_910,
    input  [151:0] col_in_911,
    input  [151:0] col_in_912,
    input  [151:0] col_in_913,
    input  [151:0] col_in_914,
    input  [151:0] col_in_915,
    input  [151:0] col_in_916,
    input  [151:0] col_in_917,
    input  [151:0] col_in_918,
    input  [151:0] col_in_919,
    input  [151:0] col_in_920,
    input  [151:0] col_in_921,
    input  [151:0] col_in_922,
    input  [151:0] col_in_923,
    input  [151:0] col_in_924,
    input  [151:0] col_in_925,
    input  [151:0] col_in_926,
    input  [151:0] col_in_927,
    input  [151:0] col_in_928,
    input  [151:0] col_in_929,
    input  [151:0] col_in_930,
    input  [151:0] col_in_931,
    input  [151:0] col_in_932,
    input  [151:0] col_in_933,
    input  [151:0] col_in_934,
    input  [151:0] col_in_935,
    input  [151:0] col_in_936,
    input  [151:0] col_in_937,
    input  [151:0] col_in_938,
    input  [151:0] col_in_939,
    input  [151:0] col_in_940,
    input  [151:0] col_in_941,
    input  [151:0] col_in_942,
    input  [151:0] col_in_943,
    input  [151:0] col_in_944,
    input  [151:0] col_in_945,
    input  [151:0] col_in_946,
    input  [151:0] col_in_947,
    input  [151:0] col_in_948,
    input  [151:0] col_in_949,
    input  [151:0] col_in_950,
    input  [151:0] col_in_951,
    input  [151:0] col_in_952,
    input  [151:0] col_in_953,
    input  [151:0] col_in_954,
    input  [151:0] col_in_955,
    input  [151:0] col_in_956,
    input  [151:0] col_in_957,
    input  [151:0] col_in_958,
    input  [151:0] col_in_959,
    input  [151:0] col_in_960,
    input  [151:0] col_in_961,
    input  [151:0] col_in_962,
    input  [151:0] col_in_963,
    input  [151:0] col_in_964,
    input  [151:0] col_in_965,
    input  [151:0] col_in_966,
    input  [151:0] col_in_967,
    input  [151:0] col_in_968,
    input  [151:0] col_in_969,
    input  [151:0] col_in_970,
    input  [151:0] col_in_971,
    input  [151:0] col_in_972,
    input  [151:0] col_in_973,
    input  [151:0] col_in_974,
    input  [151:0] col_in_975,
    input  [151:0] col_in_976,
    input  [151:0] col_in_977,
    input  [151:0] col_in_978,
    input  [151:0] col_in_979,
    input  [151:0] col_in_980,
    input  [151:0] col_in_981,
    input  [151:0] col_in_982,
    input  [151:0] col_in_983,
    input  [151:0] col_in_984,
    input  [151:0] col_in_985,
    input  [151:0] col_in_986,
    input  [151:0] col_in_987,
    input  [151:0] col_in_988,
    input  [151:0] col_in_989,
    input  [151:0] col_in_990,
    input  [151:0] col_in_991,
    input  [151:0] col_in_992,
    input  [151:0] col_in_993,
    input  [151:0] col_in_994,
    input  [151:0] col_in_995,
    input  [151:0] col_in_996,
    input  [151:0] col_in_997,
    input  [151:0] col_in_998,
    input  [151:0] col_in_999,
    input  [151:0] col_in_1000,
    input  [151:0] col_in_1001,
    input  [151:0] col_in_1002,
    input  [151:0] col_in_1003,
    input  [151:0] col_in_1004,
    input  [151:0] col_in_1005,
    input  [151:0] col_in_1006,
    input  [151:0] col_in_1007,
    input  [151:0] col_in_1008,
    input  [151:0] col_in_1009,
    input  [151:0] col_in_1010,
    input  [151:0] col_in_1011,
    input  [151:0] col_in_1012,
    input  [151:0] col_in_1013,
    input  [151:0] col_in_1014,
    input  [151:0] col_in_1015,
    input  [151:0] col_in_1016,
    input  [151:0] col_in_1017,
    input  [151:0] col_in_1018,
    input  [151:0] col_in_1019,
    input  [151:0] col_in_1020,
    input  [151:0] col_in_1021,
    input  [151:0] col_in_1022,
    input  [151:0] col_in_1023,
    input  [151:0] col_in_1024,
    input  [151:0] col_in_1025,
    input  [151:0] col_in_1026,

    output [47:0] col_out_0,
    output [47:0] col_out_1,
    output [47:0] col_out_2,
    output [47:0] col_out_3,
    output [47:0] col_out_4,
    output [47:0] col_out_5,
    output [47:0] col_out_6,
    output [47:0] col_out_7,
    output [47:0] col_out_8,
    output [47:0] col_out_9,
    output [47:0] col_out_10,
    output [47:0] col_out_11,
    output [47:0] col_out_12,
    output [47:0] col_out_13,
    output [47:0] col_out_14,
    output [47:0] col_out_15,
    output [47:0] col_out_16,
    output [47:0] col_out_17,
    output [47:0] col_out_18,
    output [47:0] col_out_19,
    output [47:0] col_out_20,
    output [47:0] col_out_21,
    output [47:0] col_out_22,
    output [47:0] col_out_23,
    output [47:0] col_out_24,
    output [47:0] col_out_25,
    output [47:0] col_out_26,
    output [47:0] col_out_27,
    output [47:0] col_out_28,
    output [47:0] col_out_29,
    output [47:0] col_out_30,
    output [47:0] col_out_31,
    output [47:0] col_out_32,
    output [47:0] col_out_33,
    output [47:0] col_out_34,
    output [47:0] col_out_35,
    output [47:0] col_out_36,
    output [47:0] col_out_37,
    output [47:0] col_out_38,
    output [47:0] col_out_39,
    output [47:0] col_out_40,
    output [47:0] col_out_41,
    output [47:0] col_out_42,
    output [47:0] col_out_43,
    output [47:0] col_out_44,
    output [47:0] col_out_45,
    output [47:0] col_out_46,
    output [47:0] col_out_47,
    output [47:0] col_out_48,
    output [47:0] col_out_49,
    output [47:0] col_out_50,
    output [47:0] col_out_51,
    output [47:0] col_out_52,
    output [47:0] col_out_53,
    output [47:0] col_out_54,
    output [47:0] col_out_55,
    output [47:0] col_out_56,
    output [47:0] col_out_57,
    output [47:0] col_out_58,
    output [47:0] col_out_59,
    output [47:0] col_out_60,
    output [47:0] col_out_61,
    output [47:0] col_out_62,
    output [47:0] col_out_63,
    output [47:0] col_out_64,
    output [47:0] col_out_65,
    output [47:0] col_out_66,
    output [47:0] col_out_67,
    output [47:0] col_out_68,
    output [47:0] col_out_69,
    output [47:0] col_out_70,
    output [47:0] col_out_71,
    output [47:0] col_out_72,
    output [47:0] col_out_73,
    output [47:0] col_out_74,
    output [47:0] col_out_75,
    output [47:0] col_out_76,
    output [47:0] col_out_77,
    output [47:0] col_out_78,
    output [47:0] col_out_79,
    output [47:0] col_out_80,
    output [47:0] col_out_81,
    output [47:0] col_out_82,
    output [47:0] col_out_83,
    output [47:0] col_out_84,
    output [47:0] col_out_85,
    output [47:0] col_out_86,
    output [47:0] col_out_87,
    output [47:0] col_out_88,
    output [47:0] col_out_89,
    output [47:0] col_out_90,
    output [47:0] col_out_91,
    output [47:0] col_out_92,
    output [47:0] col_out_93,
    output [47:0] col_out_94,
    output [47:0] col_out_95,
    output [47:0] col_out_96,
    output [47:0] col_out_97,
    output [47:0] col_out_98,
    output [47:0] col_out_99,
    output [47:0] col_out_100,
    output [47:0] col_out_101,
    output [47:0] col_out_102,
    output [47:0] col_out_103,
    output [47:0] col_out_104,
    output [47:0] col_out_105,
    output [47:0] col_out_106,
    output [47:0] col_out_107,
    output [47:0] col_out_108,
    output [47:0] col_out_109,
    output [47:0] col_out_110,
    output [47:0] col_out_111,
    output [47:0] col_out_112,
    output [47:0] col_out_113,
    output [47:0] col_out_114,
    output [47:0] col_out_115,
    output [47:0] col_out_116,
    output [47:0] col_out_117,
    output [47:0] col_out_118,
    output [47:0] col_out_119,
    output [47:0] col_out_120,
    output [47:0] col_out_121,
    output [47:0] col_out_122,
    output [47:0] col_out_123,
    output [47:0] col_out_124,
    output [47:0] col_out_125,
    output [47:0] col_out_126,
    output [47:0] col_out_127,
    output [47:0] col_out_128,
    output [47:0] col_out_129,
    output [47:0] col_out_130,
    output [47:0] col_out_131,
    output [47:0] col_out_132,
    output [47:0] col_out_133,
    output [47:0] col_out_134,
    output [47:0] col_out_135,
    output [47:0] col_out_136,
    output [47:0] col_out_137,
    output [47:0] col_out_138,
    output [47:0] col_out_139,
    output [47:0] col_out_140,
    output [47:0] col_out_141,
    output [47:0] col_out_142,
    output [47:0] col_out_143,
    output [47:0] col_out_144,
    output [47:0] col_out_145,
    output [47:0] col_out_146,
    output [47:0] col_out_147,
    output [47:0] col_out_148,
    output [47:0] col_out_149,
    output [47:0] col_out_150,
    output [47:0] col_out_151,
    output [47:0] col_out_152,
    output [47:0] col_out_153,
    output [47:0] col_out_154,
    output [47:0] col_out_155,
    output [47:0] col_out_156,
    output [47:0] col_out_157,
    output [47:0] col_out_158,
    output [47:0] col_out_159,
    output [47:0] col_out_160,
    output [47:0] col_out_161,
    output [47:0] col_out_162,
    output [47:0] col_out_163,
    output [47:0] col_out_164,
    output [47:0] col_out_165,
    output [47:0] col_out_166,
    output [47:0] col_out_167,
    output [47:0] col_out_168,
    output [47:0] col_out_169,
    output [47:0] col_out_170,
    output [47:0] col_out_171,
    output [47:0] col_out_172,
    output [47:0] col_out_173,
    output [47:0] col_out_174,
    output [47:0] col_out_175,
    output [47:0] col_out_176,
    output [47:0] col_out_177,
    output [47:0] col_out_178,
    output [47:0] col_out_179,
    output [47:0] col_out_180,
    output [47:0] col_out_181,
    output [47:0] col_out_182,
    output [47:0] col_out_183,
    output [47:0] col_out_184,
    output [47:0] col_out_185,
    output [47:0] col_out_186,
    output [47:0] col_out_187,
    output [47:0] col_out_188,
    output [47:0] col_out_189,
    output [47:0] col_out_190,
    output [47:0] col_out_191,
    output [47:0] col_out_192,
    output [47:0] col_out_193,
    output [47:0] col_out_194,
    output [47:0] col_out_195,
    output [47:0] col_out_196,
    output [47:0] col_out_197,
    output [47:0] col_out_198,
    output [47:0] col_out_199,
    output [47:0] col_out_200,
    output [47:0] col_out_201,
    output [47:0] col_out_202,
    output [47:0] col_out_203,
    output [47:0] col_out_204,
    output [47:0] col_out_205,
    output [47:0] col_out_206,
    output [47:0] col_out_207,
    output [47:0] col_out_208,
    output [47:0] col_out_209,
    output [47:0] col_out_210,
    output [47:0] col_out_211,
    output [47:0] col_out_212,
    output [47:0] col_out_213,
    output [47:0] col_out_214,
    output [47:0] col_out_215,
    output [47:0] col_out_216,
    output [47:0] col_out_217,
    output [47:0] col_out_218,
    output [47:0] col_out_219,
    output [47:0] col_out_220,
    output [47:0] col_out_221,
    output [47:0] col_out_222,
    output [47:0] col_out_223,
    output [47:0] col_out_224,
    output [47:0] col_out_225,
    output [47:0] col_out_226,
    output [47:0] col_out_227,
    output [47:0] col_out_228,
    output [47:0] col_out_229,
    output [47:0] col_out_230,
    output [47:0] col_out_231,
    output [47:0] col_out_232,
    output [47:0] col_out_233,
    output [47:0] col_out_234,
    output [47:0] col_out_235,
    output [47:0] col_out_236,
    output [47:0] col_out_237,
    output [47:0] col_out_238,
    output [47:0] col_out_239,
    output [47:0] col_out_240,
    output [47:0] col_out_241,
    output [47:0] col_out_242,
    output [47:0] col_out_243,
    output [47:0] col_out_244,
    output [47:0] col_out_245,
    output [47:0] col_out_246,
    output [47:0] col_out_247,
    output [47:0] col_out_248,
    output [47:0] col_out_249,
    output [47:0] col_out_250,
    output [47:0] col_out_251,
    output [47:0] col_out_252,
    output [47:0] col_out_253,
    output [47:0] col_out_254,
    output [47:0] col_out_255,
    output [47:0] col_out_256,
    output [47:0] col_out_257,
    output [47:0] col_out_258,
    output [47:0] col_out_259,
    output [47:0] col_out_260,
    output [47:0] col_out_261,
    output [47:0] col_out_262,
    output [47:0] col_out_263,
    output [47:0] col_out_264,
    output [47:0] col_out_265,
    output [47:0] col_out_266,
    output [47:0] col_out_267,
    output [47:0] col_out_268,
    output [47:0] col_out_269,
    output [47:0] col_out_270,
    output [47:0] col_out_271,
    output [47:0] col_out_272,
    output [47:0] col_out_273,
    output [47:0] col_out_274,
    output [47:0] col_out_275,
    output [47:0] col_out_276,
    output [47:0] col_out_277,
    output [47:0] col_out_278,
    output [47:0] col_out_279,
    output [47:0] col_out_280,
    output [47:0] col_out_281,
    output [47:0] col_out_282,
    output [47:0] col_out_283,
    output [47:0] col_out_284,
    output [47:0] col_out_285,
    output [47:0] col_out_286,
    output [47:0] col_out_287,
    output [47:0] col_out_288,
    output [47:0] col_out_289,
    output [47:0] col_out_290,
    output [47:0] col_out_291,
    output [47:0] col_out_292,
    output [47:0] col_out_293,
    output [47:0] col_out_294,
    output [47:0] col_out_295,
    output [47:0] col_out_296,
    output [47:0] col_out_297,
    output [47:0] col_out_298,
    output [47:0] col_out_299,
    output [47:0] col_out_300,
    output [47:0] col_out_301,
    output [47:0] col_out_302,
    output [47:0] col_out_303,
    output [47:0] col_out_304,
    output [47:0] col_out_305,
    output [47:0] col_out_306,
    output [47:0] col_out_307,
    output [47:0] col_out_308,
    output [47:0] col_out_309,
    output [47:0] col_out_310,
    output [47:0] col_out_311,
    output [47:0] col_out_312,
    output [47:0] col_out_313,
    output [47:0] col_out_314,
    output [47:0] col_out_315,
    output [47:0] col_out_316,
    output [47:0] col_out_317,
    output [47:0] col_out_318,
    output [47:0] col_out_319,
    output [47:0] col_out_320,
    output [47:0] col_out_321,
    output [47:0] col_out_322,
    output [47:0] col_out_323,
    output [47:0] col_out_324,
    output [47:0] col_out_325,
    output [47:0] col_out_326,
    output [47:0] col_out_327,
    output [47:0] col_out_328,
    output [47:0] col_out_329,
    output [47:0] col_out_330,
    output [47:0] col_out_331,
    output [47:0] col_out_332,
    output [47:0] col_out_333,
    output [47:0] col_out_334,
    output [47:0] col_out_335,
    output [47:0] col_out_336,
    output [47:0] col_out_337,
    output [47:0] col_out_338,
    output [47:0] col_out_339,
    output [47:0] col_out_340,
    output [47:0] col_out_341,
    output [47:0] col_out_342,
    output [47:0] col_out_343,
    output [47:0] col_out_344,
    output [47:0] col_out_345,
    output [47:0] col_out_346,
    output [47:0] col_out_347,
    output [47:0] col_out_348,
    output [47:0] col_out_349,
    output [47:0] col_out_350,
    output [47:0] col_out_351,
    output [47:0] col_out_352,
    output [47:0] col_out_353,
    output [47:0] col_out_354,
    output [47:0] col_out_355,
    output [47:0] col_out_356,
    output [47:0] col_out_357,
    output [47:0] col_out_358,
    output [47:0] col_out_359,
    output [47:0] col_out_360,
    output [47:0] col_out_361,
    output [47:0] col_out_362,
    output [47:0] col_out_363,
    output [47:0] col_out_364,
    output [47:0] col_out_365,
    output [47:0] col_out_366,
    output [47:0] col_out_367,
    output [47:0] col_out_368,
    output [47:0] col_out_369,
    output [47:0] col_out_370,
    output [47:0] col_out_371,
    output [47:0] col_out_372,
    output [47:0] col_out_373,
    output [47:0] col_out_374,
    output [47:0] col_out_375,
    output [47:0] col_out_376,
    output [47:0] col_out_377,
    output [47:0] col_out_378,
    output [47:0] col_out_379,
    output [47:0] col_out_380,
    output [47:0] col_out_381,
    output [47:0] col_out_382,
    output [47:0] col_out_383,
    output [47:0] col_out_384,
    output [47:0] col_out_385,
    output [47:0] col_out_386,
    output [47:0] col_out_387,
    output [47:0] col_out_388,
    output [47:0] col_out_389,
    output [47:0] col_out_390,
    output [47:0] col_out_391,
    output [47:0] col_out_392,
    output [47:0] col_out_393,
    output [47:0] col_out_394,
    output [47:0] col_out_395,
    output [47:0] col_out_396,
    output [47:0] col_out_397,
    output [47:0] col_out_398,
    output [47:0] col_out_399,
    output [47:0] col_out_400,
    output [47:0] col_out_401,
    output [47:0] col_out_402,
    output [47:0] col_out_403,
    output [47:0] col_out_404,
    output [47:0] col_out_405,
    output [47:0] col_out_406,
    output [47:0] col_out_407,
    output [47:0] col_out_408,
    output [47:0] col_out_409,
    output [47:0] col_out_410,
    output [47:0] col_out_411,
    output [47:0] col_out_412,
    output [47:0] col_out_413,
    output [47:0] col_out_414,
    output [47:0] col_out_415,
    output [47:0] col_out_416,
    output [47:0] col_out_417,
    output [47:0] col_out_418,
    output [47:0] col_out_419,
    output [47:0] col_out_420,
    output [47:0] col_out_421,
    output [47:0] col_out_422,
    output [47:0] col_out_423,
    output [47:0] col_out_424,
    output [47:0] col_out_425,
    output [47:0] col_out_426,
    output [47:0] col_out_427,
    output [47:0] col_out_428,
    output [47:0] col_out_429,
    output [47:0] col_out_430,
    output [47:0] col_out_431,
    output [47:0] col_out_432,
    output [47:0] col_out_433,
    output [47:0] col_out_434,
    output [47:0] col_out_435,
    output [47:0] col_out_436,
    output [47:0] col_out_437,
    output [47:0] col_out_438,
    output [47:0] col_out_439,
    output [47:0] col_out_440,
    output [47:0] col_out_441,
    output [47:0] col_out_442,
    output [47:0] col_out_443,
    output [47:0] col_out_444,
    output [47:0] col_out_445,
    output [47:0] col_out_446,
    output [47:0] col_out_447,
    output [47:0] col_out_448,
    output [47:0] col_out_449,
    output [47:0] col_out_450,
    output [47:0] col_out_451,
    output [47:0] col_out_452,
    output [47:0] col_out_453,
    output [47:0] col_out_454,
    output [47:0] col_out_455,
    output [47:0] col_out_456,
    output [47:0] col_out_457,
    output [47:0] col_out_458,
    output [47:0] col_out_459,
    output [47:0] col_out_460,
    output [47:0] col_out_461,
    output [47:0] col_out_462,
    output [47:0] col_out_463,
    output [47:0] col_out_464,
    output [47:0] col_out_465,
    output [47:0] col_out_466,
    output [47:0] col_out_467,
    output [47:0] col_out_468,
    output [47:0] col_out_469,
    output [47:0] col_out_470,
    output [47:0] col_out_471,
    output [47:0] col_out_472,
    output [47:0] col_out_473,
    output [47:0] col_out_474,
    output [47:0] col_out_475,
    output [47:0] col_out_476,
    output [47:0] col_out_477,
    output [47:0] col_out_478,
    output [47:0] col_out_479,
    output [47:0] col_out_480,
    output [47:0] col_out_481,
    output [47:0] col_out_482,
    output [47:0] col_out_483,
    output [47:0] col_out_484,
    output [47:0] col_out_485,
    output [47:0] col_out_486,
    output [47:0] col_out_487,
    output [47:0] col_out_488,
    output [47:0] col_out_489,
    output [47:0] col_out_490,
    output [47:0] col_out_491,
    output [47:0] col_out_492,
    output [47:0] col_out_493,
    output [47:0] col_out_494,
    output [47:0] col_out_495,
    output [47:0] col_out_496,
    output [47:0] col_out_497,
    output [47:0] col_out_498,
    output [47:0] col_out_499,
    output [47:0] col_out_500,
    output [47:0] col_out_501,
    output [47:0] col_out_502,
    output [47:0] col_out_503,
    output [47:0] col_out_504,
    output [47:0] col_out_505,
    output [47:0] col_out_506,
    output [47:0] col_out_507,
    output [47:0] col_out_508,
    output [47:0] col_out_509,
    output [47:0] col_out_510,
    output [47:0] col_out_511,
    output [47:0] col_out_512,
    output [47:0] col_out_513,
    output [47:0] col_out_514,
    output [47:0] col_out_515,
    output [47:0] col_out_516,
    output [47:0] col_out_517,
    output [47:0] col_out_518,
    output [47:0] col_out_519,
    output [47:0] col_out_520,
    output [47:0] col_out_521,
    output [47:0] col_out_522,
    output [47:0] col_out_523,
    output [47:0] col_out_524,
    output [47:0] col_out_525,
    output [47:0] col_out_526,
    output [47:0] col_out_527,
    output [47:0] col_out_528,
    output [47:0] col_out_529,
    output [47:0] col_out_530,
    output [47:0] col_out_531,
    output [47:0] col_out_532,
    output [47:0] col_out_533,
    output [47:0] col_out_534,
    output [47:0] col_out_535,
    output [47:0] col_out_536,
    output [47:0] col_out_537,
    output [47:0] col_out_538,
    output [47:0] col_out_539,
    output [47:0] col_out_540,
    output [47:0] col_out_541,
    output [47:0] col_out_542,
    output [47:0] col_out_543,
    output [47:0] col_out_544,
    output [47:0] col_out_545,
    output [47:0] col_out_546,
    output [47:0] col_out_547,
    output [47:0] col_out_548,
    output [47:0] col_out_549,
    output [47:0] col_out_550,
    output [47:0] col_out_551,
    output [47:0] col_out_552,
    output [47:0] col_out_553,
    output [47:0] col_out_554,
    output [47:0] col_out_555,
    output [47:0] col_out_556,
    output [47:0] col_out_557,
    output [47:0] col_out_558,
    output [47:0] col_out_559,
    output [47:0] col_out_560,
    output [47:0] col_out_561,
    output [47:0] col_out_562,
    output [47:0] col_out_563,
    output [47:0] col_out_564,
    output [47:0] col_out_565,
    output [47:0] col_out_566,
    output [47:0] col_out_567,
    output [47:0] col_out_568,
    output [47:0] col_out_569,
    output [47:0] col_out_570,
    output [47:0] col_out_571,
    output [47:0] col_out_572,
    output [47:0] col_out_573,
    output [47:0] col_out_574,
    output [47:0] col_out_575,
    output [47:0] col_out_576,
    output [47:0] col_out_577,
    output [47:0] col_out_578,
    output [47:0] col_out_579,
    output [47:0] col_out_580,
    output [47:0] col_out_581,
    output [47:0] col_out_582,
    output [47:0] col_out_583,
    output [47:0] col_out_584,
    output [47:0] col_out_585,
    output [47:0] col_out_586,
    output [47:0] col_out_587,
    output [47:0] col_out_588,
    output [47:0] col_out_589,
    output [47:0] col_out_590,
    output [47:0] col_out_591,
    output [47:0] col_out_592,
    output [47:0] col_out_593,
    output [47:0] col_out_594,
    output [47:0] col_out_595,
    output [47:0] col_out_596,
    output [47:0] col_out_597,
    output [47:0] col_out_598,
    output [47:0] col_out_599,
    output [47:0] col_out_600,
    output [47:0] col_out_601,
    output [47:0] col_out_602,
    output [47:0] col_out_603,
    output [47:0] col_out_604,
    output [47:0] col_out_605,
    output [47:0] col_out_606,
    output [47:0] col_out_607,
    output [47:0] col_out_608,
    output [47:0] col_out_609,
    output [47:0] col_out_610,
    output [47:0] col_out_611,
    output [47:0] col_out_612,
    output [47:0] col_out_613,
    output [47:0] col_out_614,
    output [47:0] col_out_615,
    output [47:0] col_out_616,
    output [47:0] col_out_617,
    output [47:0] col_out_618,
    output [47:0] col_out_619,
    output [47:0] col_out_620,
    output [47:0] col_out_621,
    output [47:0] col_out_622,
    output [47:0] col_out_623,
    output [47:0] col_out_624,
    output [47:0] col_out_625,
    output [47:0] col_out_626,
    output [47:0] col_out_627,
    output [47:0] col_out_628,
    output [47:0] col_out_629,
    output [47:0] col_out_630,
    output [47:0] col_out_631,
    output [47:0] col_out_632,
    output [47:0] col_out_633,
    output [47:0] col_out_634,
    output [47:0] col_out_635,
    output [47:0] col_out_636,
    output [47:0] col_out_637,
    output [47:0] col_out_638,
    output [47:0] col_out_639,
    output [47:0] col_out_640,
    output [47:0] col_out_641,
    output [47:0] col_out_642,
    output [47:0] col_out_643,
    output [47:0] col_out_644,
    output [47:0] col_out_645,
    output [47:0] col_out_646,
    output [47:0] col_out_647,
    output [47:0] col_out_648,
    output [47:0] col_out_649,
    output [47:0] col_out_650,
    output [47:0] col_out_651,
    output [47:0] col_out_652,
    output [47:0] col_out_653,
    output [47:0] col_out_654,
    output [47:0] col_out_655,
    output [47:0] col_out_656,
    output [47:0] col_out_657,
    output [47:0] col_out_658,
    output [47:0] col_out_659,
    output [47:0] col_out_660,
    output [47:0] col_out_661,
    output [47:0] col_out_662,
    output [47:0] col_out_663,
    output [47:0] col_out_664,
    output [47:0] col_out_665,
    output [47:0] col_out_666,
    output [47:0] col_out_667,
    output [47:0] col_out_668,
    output [47:0] col_out_669,
    output [47:0] col_out_670,
    output [47:0] col_out_671,
    output [47:0] col_out_672,
    output [47:0] col_out_673,
    output [47:0] col_out_674,
    output [47:0] col_out_675,
    output [47:0] col_out_676,
    output [47:0] col_out_677,
    output [47:0] col_out_678,
    output [47:0] col_out_679,
    output [47:0] col_out_680,
    output [47:0] col_out_681,
    output [47:0] col_out_682,
    output [47:0] col_out_683,
    output [47:0] col_out_684,
    output [47:0] col_out_685,
    output [47:0] col_out_686,
    output [47:0] col_out_687,
    output [47:0] col_out_688,
    output [47:0] col_out_689,
    output [47:0] col_out_690,
    output [47:0] col_out_691,
    output [47:0] col_out_692,
    output [47:0] col_out_693,
    output [47:0] col_out_694,
    output [47:0] col_out_695,
    output [47:0] col_out_696,
    output [47:0] col_out_697,
    output [47:0] col_out_698,
    output [47:0] col_out_699,
    output [47:0] col_out_700,
    output [47:0] col_out_701,
    output [47:0] col_out_702,
    output [47:0] col_out_703,
    output [47:0] col_out_704,
    output [47:0] col_out_705,
    output [47:0] col_out_706,
    output [47:0] col_out_707,
    output [47:0] col_out_708,
    output [47:0] col_out_709,
    output [47:0] col_out_710,
    output [47:0] col_out_711,
    output [47:0] col_out_712,
    output [47:0] col_out_713,
    output [47:0] col_out_714,
    output [47:0] col_out_715,
    output [47:0] col_out_716,
    output [47:0] col_out_717,
    output [47:0] col_out_718,
    output [47:0] col_out_719,
    output [47:0] col_out_720,
    output [47:0] col_out_721,
    output [47:0] col_out_722,
    output [47:0] col_out_723,
    output [47:0] col_out_724,
    output [47:0] col_out_725,
    output [47:0] col_out_726,
    output [47:0] col_out_727,
    output [47:0] col_out_728,
    output [47:0] col_out_729,
    output [47:0] col_out_730,
    output [47:0] col_out_731,
    output [47:0] col_out_732,
    output [47:0] col_out_733,
    output [47:0] col_out_734,
    output [47:0] col_out_735,
    output [47:0] col_out_736,
    output [47:0] col_out_737,
    output [47:0] col_out_738,
    output [47:0] col_out_739,
    output [47:0] col_out_740,
    output [47:0] col_out_741,
    output [47:0] col_out_742,
    output [47:0] col_out_743,
    output [47:0] col_out_744,
    output [47:0] col_out_745,
    output [47:0] col_out_746,
    output [47:0] col_out_747,
    output [47:0] col_out_748,
    output [47:0] col_out_749,
    output [47:0] col_out_750,
    output [47:0] col_out_751,
    output [47:0] col_out_752,
    output [47:0] col_out_753,
    output [47:0] col_out_754,
    output [47:0] col_out_755,
    output [47:0] col_out_756,
    output [47:0] col_out_757,
    output [47:0] col_out_758,
    output [47:0] col_out_759,
    output [47:0] col_out_760,
    output [47:0] col_out_761,
    output [47:0] col_out_762,
    output [47:0] col_out_763,
    output [47:0] col_out_764,
    output [47:0] col_out_765,
    output [47:0] col_out_766,
    output [47:0] col_out_767,
    output [47:0] col_out_768,
    output [47:0] col_out_769,
    output [47:0] col_out_770,
    output [47:0] col_out_771,
    output [47:0] col_out_772,
    output [47:0] col_out_773,
    output [47:0] col_out_774,
    output [47:0] col_out_775,
    output [47:0] col_out_776,
    output [47:0] col_out_777,
    output [47:0] col_out_778,
    output [47:0] col_out_779,
    output [47:0] col_out_780,
    output [47:0] col_out_781,
    output [47:0] col_out_782,
    output [47:0] col_out_783,
    output [47:0] col_out_784,
    output [47:0] col_out_785,
    output [47:0] col_out_786,
    output [47:0] col_out_787,
    output [47:0] col_out_788,
    output [47:0] col_out_789,
    output [47:0] col_out_790,
    output [47:0] col_out_791,
    output [47:0] col_out_792,
    output [47:0] col_out_793,
    output [47:0] col_out_794,
    output [47:0] col_out_795,
    output [47:0] col_out_796,
    output [47:0] col_out_797,
    output [47:0] col_out_798,
    output [47:0] col_out_799,
    output [47:0] col_out_800,
    output [47:0] col_out_801,
    output [47:0] col_out_802,
    output [47:0] col_out_803,
    output [47:0] col_out_804,
    output [47:0] col_out_805,
    output [47:0] col_out_806,
    output [47:0] col_out_807,
    output [47:0] col_out_808,
    output [47:0] col_out_809,
    output [47:0] col_out_810,
    output [47:0] col_out_811,
    output [47:0] col_out_812,
    output [47:0] col_out_813,
    output [47:0] col_out_814,
    output [47:0] col_out_815,
    output [47:0] col_out_816,
    output [47:0] col_out_817,
    output [47:0] col_out_818,
    output [47:0] col_out_819,
    output [47:0] col_out_820,
    output [47:0] col_out_821,
    output [47:0] col_out_822,
    output [47:0] col_out_823,
    output [47:0] col_out_824,
    output [47:0] col_out_825,
    output [47:0] col_out_826,
    output [47:0] col_out_827,
    output [47:0] col_out_828,
    output [47:0] col_out_829,
    output [47:0] col_out_830,
    output [47:0] col_out_831,
    output [47:0] col_out_832,
    output [47:0] col_out_833,
    output [47:0] col_out_834,
    output [47:0] col_out_835,
    output [47:0] col_out_836,
    output [47:0] col_out_837,
    output [47:0] col_out_838,
    output [47:0] col_out_839,
    output [47:0] col_out_840,
    output [47:0] col_out_841,
    output [47:0] col_out_842,
    output [47:0] col_out_843,
    output [47:0] col_out_844,
    output [47:0] col_out_845,
    output [47:0] col_out_846,
    output [47:0] col_out_847,
    output [47:0] col_out_848,
    output [47:0] col_out_849,
    output [47:0] col_out_850,
    output [47:0] col_out_851,
    output [47:0] col_out_852,
    output [47:0] col_out_853,
    output [47:0] col_out_854,
    output [47:0] col_out_855,
    output [47:0] col_out_856,
    output [47:0] col_out_857,
    output [47:0] col_out_858,
    output [47:0] col_out_859,
    output [47:0] col_out_860,
    output [47:0] col_out_861,
    output [47:0] col_out_862,
    output [47:0] col_out_863,
    output [47:0] col_out_864,
    output [47:0] col_out_865,
    output [47:0] col_out_866,
    output [47:0] col_out_867,
    output [47:0] col_out_868,
    output [47:0] col_out_869,
    output [47:0] col_out_870,
    output [47:0] col_out_871,
    output [47:0] col_out_872,
    output [47:0] col_out_873,
    output [47:0] col_out_874,
    output [47:0] col_out_875,
    output [47:0] col_out_876,
    output [47:0] col_out_877,
    output [47:0] col_out_878,
    output [47:0] col_out_879,
    output [47:0] col_out_880,
    output [47:0] col_out_881,
    output [47:0] col_out_882,
    output [47:0] col_out_883,
    output [47:0] col_out_884,
    output [47:0] col_out_885,
    output [47:0] col_out_886,
    output [47:0] col_out_887,
    output [47:0] col_out_888,
    output [47:0] col_out_889,
    output [47:0] col_out_890,
    output [47:0] col_out_891,
    output [47:0] col_out_892,
    output [47:0] col_out_893,
    output [47:0] col_out_894,
    output [47:0] col_out_895,
    output [47:0] col_out_896,
    output [47:0] col_out_897,
    output [47:0] col_out_898,
    output [47:0] col_out_899,
    output [47:0] col_out_900,
    output [47:0] col_out_901,
    output [47:0] col_out_902,
    output [47:0] col_out_903,
    output [47:0] col_out_904,
    output [47:0] col_out_905,
    output [47:0] col_out_906,
    output [47:0] col_out_907,
    output [47:0] col_out_908,
    output [47:0] col_out_909,
    output [47:0] col_out_910,
    output [47:0] col_out_911,
    output [47:0] col_out_912,
    output [47:0] col_out_913,
    output [47:0] col_out_914,
    output [47:0] col_out_915,
    output [47:0] col_out_916,
    output [47:0] col_out_917,
    output [47:0] col_out_918,
    output [47:0] col_out_919,
    output [47:0] col_out_920,
    output [47:0] col_out_921,
    output [47:0] col_out_922,
    output [47:0] col_out_923,
    output [47:0] col_out_924,
    output [47:0] col_out_925,
    output [47:0] col_out_926,
    output [47:0] col_out_927,
    output [47:0] col_out_928,
    output [47:0] col_out_929,
    output [47:0] col_out_930,
    output [47:0] col_out_931,
    output [47:0] col_out_932,
    output [47:0] col_out_933,
    output [47:0] col_out_934,
    output [47:0] col_out_935,
    output [47:0] col_out_936,
    output [47:0] col_out_937,
    output [47:0] col_out_938,
    output [47:0] col_out_939,
    output [47:0] col_out_940,
    output [47:0] col_out_941,
    output [47:0] col_out_942,
    output [47:0] col_out_943,
    output [47:0] col_out_944,
    output [47:0] col_out_945,
    output [47:0] col_out_946,
    output [47:0] col_out_947,
    output [47:0] col_out_948,
    output [47:0] col_out_949,
    output [47:0] col_out_950,
    output [47:0] col_out_951,
    output [47:0] col_out_952,
    output [47:0] col_out_953,
    output [47:0] col_out_954,
    output [47:0] col_out_955,
    output [47:0] col_out_956,
    output [47:0] col_out_957,
    output [47:0] col_out_958,
    output [47:0] col_out_959,
    output [47:0] col_out_960,
    output [47:0] col_out_961,
    output [47:0] col_out_962,
    output [47:0] col_out_963,
    output [47:0] col_out_964,
    output [47:0] col_out_965,
    output [47:0] col_out_966,
    output [47:0] col_out_967,
    output [47:0] col_out_968,
    output [47:0] col_out_969,
    output [47:0] col_out_970,
    output [47:0] col_out_971,
    output [47:0] col_out_972,
    output [47:0] col_out_973,
    output [47:0] col_out_974,
    output [47:0] col_out_975,
    output [47:0] col_out_976,
    output [47:0] col_out_977,
    output [47:0] col_out_978,
    output [47:0] col_out_979,
    output [47:0] col_out_980,
    output [47:0] col_out_981,
    output [47:0] col_out_982,
    output [47:0] col_out_983,
    output [47:0] col_out_984,
    output [47:0] col_out_985,
    output [47:0] col_out_986,
    output [47:0] col_out_987,
    output [47:0] col_out_988,
    output [47:0] col_out_989,
    output [47:0] col_out_990,
    output [47:0] col_out_991,
    output [47:0] col_out_992,
    output [47:0] col_out_993,
    output [47:0] col_out_994,
    output [47:0] col_out_995,
    output [47:0] col_out_996,
    output [47:0] col_out_997,
    output [47:0] col_out_998,
    output [47:0] col_out_999,
    output [47:0] col_out_1000,
    output [47:0] col_out_1001,
    output [47:0] col_out_1002,
    output [47:0] col_out_1003,
    output [47:0] col_out_1004,
    output [47:0] col_out_1005,
    output [47:0] col_out_1006,
    output [47:0] col_out_1007,
    output [47:0] col_out_1008,
    output [47:0] col_out_1009,
    output [47:0] col_out_1010,
    output [47:0] col_out_1011,
    output [47:0] col_out_1012,
    output [47:0] col_out_1013,
    output [47:0] col_out_1014,
    output [47:0] col_out_1015,
    output [47:0] col_out_1016,
    output [47:0] col_out_1017,
    output [47:0] col_out_1018,
    output [47:0] col_out_1019,
    output [47:0] col_out_1020,
    output [47:0] col_out_1021,
    output [47:0] col_out_1022,
    output [47:0] col_out_1023,
    output [47:0] col_out_1024,
    output [47:0] col_out_1025,
    output [47:0] col_out_1026,
    output [47:0] col_out_1027,
    output [47:0] col_out_1028,
    output [47:0] col_out_1029
);



//--compressor_array input and output----------------------

wire [161:0] u_ca_in_0;
wire [161:0] u_ca_in_1;
wire [161:0] u_ca_in_2;
wire [161:0] u_ca_in_3;
wire [161:0] u_ca_in_4;
wire [161:0] u_ca_in_5;
wire [161:0] u_ca_in_6;
wire [161:0] u_ca_in_7;
wire [161:0] u_ca_in_8;
wire [161:0] u_ca_in_9;
wire [161:0] u_ca_in_10;
wire [161:0] u_ca_in_11;
wire [161:0] u_ca_in_12;
wire [161:0] u_ca_in_13;
wire [161:0] u_ca_in_14;
wire [161:0] u_ca_in_15;
wire [161:0] u_ca_in_16;
wire [161:0] u_ca_in_17;
wire [161:0] u_ca_in_18;
wire [161:0] u_ca_in_19;
wire [161:0] u_ca_in_20;
wire [161:0] u_ca_in_21;
wire [161:0] u_ca_in_22;
wire [161:0] u_ca_in_23;
wire [161:0] u_ca_in_24;
wire [161:0] u_ca_in_25;
wire [161:0] u_ca_in_26;
wire [161:0] u_ca_in_27;
wire [161:0] u_ca_in_28;
wire [161:0] u_ca_in_29;
wire [161:0] u_ca_in_30;
wire [161:0] u_ca_in_31;
wire [161:0] u_ca_in_32;
wire [161:0] u_ca_in_33;
wire [161:0] u_ca_in_34;
wire [161:0] u_ca_in_35;
wire [161:0] u_ca_in_36;
wire [161:0] u_ca_in_37;
wire [161:0] u_ca_in_38;
wire [161:0] u_ca_in_39;
wire [161:0] u_ca_in_40;
wire [161:0] u_ca_in_41;
wire [161:0] u_ca_in_42;
wire [161:0] u_ca_in_43;
wire [161:0] u_ca_in_44;
wire [161:0] u_ca_in_45;
wire [161:0] u_ca_in_46;
wire [161:0] u_ca_in_47;
wire [161:0] u_ca_in_48;
wire [161:0] u_ca_in_49;
wire [161:0] u_ca_in_50;
wire [161:0] u_ca_in_51;
wire [161:0] u_ca_in_52;
wire [161:0] u_ca_in_53;
wire [161:0] u_ca_in_54;
wire [161:0] u_ca_in_55;
wire [161:0] u_ca_in_56;
wire [161:0] u_ca_in_57;
wire [161:0] u_ca_in_58;
wire [161:0] u_ca_in_59;
wire [161:0] u_ca_in_60;
wire [161:0] u_ca_in_61;
wire [161:0] u_ca_in_62;
wire [161:0] u_ca_in_63;
wire [161:0] u_ca_in_64;
wire [161:0] u_ca_in_65;
wire [161:0] u_ca_in_66;
wire [161:0] u_ca_in_67;
wire [161:0] u_ca_in_68;
wire [161:0] u_ca_in_69;
wire [161:0] u_ca_in_70;
wire [161:0] u_ca_in_71;
wire [161:0] u_ca_in_72;
wire [161:0] u_ca_in_73;
wire [161:0] u_ca_in_74;
wire [161:0] u_ca_in_75;
wire [161:0] u_ca_in_76;
wire [161:0] u_ca_in_77;
wire [161:0] u_ca_in_78;
wire [161:0] u_ca_in_79;
wire [161:0] u_ca_in_80;
wire [161:0] u_ca_in_81;
wire [161:0] u_ca_in_82;
wire [161:0] u_ca_in_83;
wire [161:0] u_ca_in_84;
wire [161:0] u_ca_in_85;
wire [161:0] u_ca_in_86;
wire [161:0] u_ca_in_87;
wire [161:0] u_ca_in_88;
wire [161:0] u_ca_in_89;
wire [161:0] u_ca_in_90;
wire [161:0] u_ca_in_91;
wire [161:0] u_ca_in_92;
wire [161:0] u_ca_in_93;
wire [161:0] u_ca_in_94;
wire [161:0] u_ca_in_95;
wire [161:0] u_ca_in_96;
wire [161:0] u_ca_in_97;
wire [161:0] u_ca_in_98;
wire [161:0] u_ca_in_99;
wire [161:0] u_ca_in_100;
wire [161:0] u_ca_in_101;
wire [161:0] u_ca_in_102;
wire [161:0] u_ca_in_103;
wire [161:0] u_ca_in_104;
wire [161:0] u_ca_in_105;
wire [161:0] u_ca_in_106;
wire [161:0] u_ca_in_107;
wire [161:0] u_ca_in_108;
wire [161:0] u_ca_in_109;
wire [161:0] u_ca_in_110;
wire [161:0] u_ca_in_111;
wire [161:0] u_ca_in_112;
wire [161:0] u_ca_in_113;
wire [161:0] u_ca_in_114;
wire [161:0] u_ca_in_115;
wire [161:0] u_ca_in_116;
wire [161:0] u_ca_in_117;
wire [161:0] u_ca_in_118;
wire [161:0] u_ca_in_119;
wire [161:0] u_ca_in_120;
wire [161:0] u_ca_in_121;
wire [161:0] u_ca_in_122;
wire [161:0] u_ca_in_123;
wire [161:0] u_ca_in_124;
wire [161:0] u_ca_in_125;
wire [161:0] u_ca_in_126;
wire [161:0] u_ca_in_127;
wire [161:0] u_ca_in_128;
wire [161:0] u_ca_in_129;
wire [161:0] u_ca_in_130;
wire [161:0] u_ca_in_131;
wire [161:0] u_ca_in_132;
wire [161:0] u_ca_in_133;
wire [161:0] u_ca_in_134;
wire [161:0] u_ca_in_135;
wire [161:0] u_ca_in_136;
wire [161:0] u_ca_in_137;
wire [161:0] u_ca_in_138;
wire [161:0] u_ca_in_139;
wire [161:0] u_ca_in_140;
wire [161:0] u_ca_in_141;
wire [161:0] u_ca_in_142;
wire [161:0] u_ca_in_143;
wire [161:0] u_ca_in_144;
wire [161:0] u_ca_in_145;
wire [161:0] u_ca_in_146;
wire [161:0] u_ca_in_147;
wire [161:0] u_ca_in_148;
wire [161:0] u_ca_in_149;
wire [161:0] u_ca_in_150;
wire [161:0] u_ca_in_151;
wire [161:0] u_ca_in_152;
wire [161:0] u_ca_in_153;
wire [161:0] u_ca_in_154;
wire [161:0] u_ca_in_155;
wire [161:0] u_ca_in_156;
wire [161:0] u_ca_in_157;
wire [161:0] u_ca_in_158;
wire [161:0] u_ca_in_159;
wire [161:0] u_ca_in_160;
wire [161:0] u_ca_in_161;
wire [161:0] u_ca_in_162;
wire [161:0] u_ca_in_163;
wire [161:0] u_ca_in_164;
wire [161:0] u_ca_in_165;
wire [161:0] u_ca_in_166;
wire [161:0] u_ca_in_167;
wire [161:0] u_ca_in_168;
wire [161:0] u_ca_in_169;
wire [161:0] u_ca_in_170;
wire [161:0] u_ca_in_171;
wire [161:0] u_ca_in_172;
wire [161:0] u_ca_in_173;
wire [161:0] u_ca_in_174;
wire [161:0] u_ca_in_175;
wire [161:0] u_ca_in_176;
wire [161:0] u_ca_in_177;
wire [161:0] u_ca_in_178;
wire [161:0] u_ca_in_179;
wire [161:0] u_ca_in_180;
wire [161:0] u_ca_in_181;
wire [161:0] u_ca_in_182;
wire [161:0] u_ca_in_183;
wire [161:0] u_ca_in_184;
wire [161:0] u_ca_in_185;
wire [161:0] u_ca_in_186;
wire [161:0] u_ca_in_187;
wire [161:0] u_ca_in_188;
wire [161:0] u_ca_in_189;
wire [161:0] u_ca_in_190;
wire [161:0] u_ca_in_191;
wire [161:0] u_ca_in_192;
wire [161:0] u_ca_in_193;
wire [161:0] u_ca_in_194;
wire [161:0] u_ca_in_195;
wire [161:0] u_ca_in_196;
wire [161:0] u_ca_in_197;
wire [161:0] u_ca_in_198;
wire [161:0] u_ca_in_199;
wire [161:0] u_ca_in_200;
wire [161:0] u_ca_in_201;
wire [161:0] u_ca_in_202;
wire [161:0] u_ca_in_203;
wire [161:0] u_ca_in_204;
wire [161:0] u_ca_in_205;
wire [161:0] u_ca_in_206;
wire [161:0] u_ca_in_207;
wire [161:0] u_ca_in_208;
wire [161:0] u_ca_in_209;
wire [161:0] u_ca_in_210;
wire [161:0] u_ca_in_211;
wire [161:0] u_ca_in_212;
wire [161:0] u_ca_in_213;
wire [161:0] u_ca_in_214;
wire [161:0] u_ca_in_215;
wire [161:0] u_ca_in_216;
wire [161:0] u_ca_in_217;
wire [161:0] u_ca_in_218;
wire [161:0] u_ca_in_219;
wire [161:0] u_ca_in_220;
wire [161:0] u_ca_in_221;
wire [161:0] u_ca_in_222;
wire [161:0] u_ca_in_223;
wire [161:0] u_ca_in_224;
wire [161:0] u_ca_in_225;
wire [161:0] u_ca_in_226;
wire [161:0] u_ca_in_227;
wire [161:0] u_ca_in_228;
wire [161:0] u_ca_in_229;
wire [161:0] u_ca_in_230;
wire [161:0] u_ca_in_231;
wire [161:0] u_ca_in_232;
wire [161:0] u_ca_in_233;
wire [161:0] u_ca_in_234;
wire [161:0] u_ca_in_235;
wire [161:0] u_ca_in_236;
wire [161:0] u_ca_in_237;
wire [161:0] u_ca_in_238;
wire [161:0] u_ca_in_239;
wire [161:0] u_ca_in_240;
wire [161:0] u_ca_in_241;
wire [161:0] u_ca_in_242;
wire [161:0] u_ca_in_243;
wire [161:0] u_ca_in_244;
wire [161:0] u_ca_in_245;
wire [161:0] u_ca_in_246;
wire [161:0] u_ca_in_247;
wire [161:0] u_ca_in_248;
wire [161:0] u_ca_in_249;
wire [161:0] u_ca_in_250;
wire [161:0] u_ca_in_251;
wire [161:0] u_ca_in_252;
wire [161:0] u_ca_in_253;
wire [161:0] u_ca_in_254;
wire [161:0] u_ca_in_255;
wire [161:0] u_ca_in_256;
wire [161:0] u_ca_in_257;
wire [161:0] u_ca_in_258;
wire [161:0] u_ca_in_259;
wire [161:0] u_ca_in_260;
wire [161:0] u_ca_in_261;
wire [161:0] u_ca_in_262;
wire [161:0] u_ca_in_263;
wire [161:0] u_ca_in_264;
wire [161:0] u_ca_in_265;
wire [161:0] u_ca_in_266;
wire [161:0] u_ca_in_267;
wire [161:0] u_ca_in_268;
wire [161:0] u_ca_in_269;
wire [161:0] u_ca_in_270;
wire [161:0] u_ca_in_271;
wire [161:0] u_ca_in_272;
wire [161:0] u_ca_in_273;
wire [161:0] u_ca_in_274;
wire [161:0] u_ca_in_275;
wire [161:0] u_ca_in_276;
wire [161:0] u_ca_in_277;
wire [161:0] u_ca_in_278;
wire [161:0] u_ca_in_279;
wire [161:0] u_ca_in_280;
wire [161:0] u_ca_in_281;
wire [161:0] u_ca_in_282;
wire [161:0] u_ca_in_283;
wire [161:0] u_ca_in_284;
wire [161:0] u_ca_in_285;
wire [161:0] u_ca_in_286;
wire [161:0] u_ca_in_287;
wire [161:0] u_ca_in_288;
wire [161:0] u_ca_in_289;
wire [161:0] u_ca_in_290;
wire [161:0] u_ca_in_291;
wire [161:0] u_ca_in_292;
wire [161:0] u_ca_in_293;
wire [161:0] u_ca_in_294;
wire [161:0] u_ca_in_295;
wire [161:0] u_ca_in_296;
wire [161:0] u_ca_in_297;
wire [161:0] u_ca_in_298;
wire [161:0] u_ca_in_299;
wire [161:0] u_ca_in_300;
wire [161:0] u_ca_in_301;
wire [161:0] u_ca_in_302;
wire [161:0] u_ca_in_303;
wire [161:0] u_ca_in_304;
wire [161:0] u_ca_in_305;
wire [161:0] u_ca_in_306;
wire [161:0] u_ca_in_307;
wire [161:0] u_ca_in_308;
wire [161:0] u_ca_in_309;
wire [161:0] u_ca_in_310;
wire [161:0] u_ca_in_311;
wire [161:0] u_ca_in_312;
wire [161:0] u_ca_in_313;
wire [161:0] u_ca_in_314;
wire [161:0] u_ca_in_315;
wire [161:0] u_ca_in_316;
wire [161:0] u_ca_in_317;
wire [161:0] u_ca_in_318;
wire [161:0] u_ca_in_319;
wire [161:0] u_ca_in_320;
wire [161:0] u_ca_in_321;
wire [161:0] u_ca_in_322;
wire [161:0] u_ca_in_323;
wire [161:0] u_ca_in_324;
wire [161:0] u_ca_in_325;
wire [161:0] u_ca_in_326;
wire [161:0] u_ca_in_327;
wire [161:0] u_ca_in_328;
wire [161:0] u_ca_in_329;
wire [161:0] u_ca_in_330;
wire [161:0] u_ca_in_331;
wire [161:0] u_ca_in_332;
wire [161:0] u_ca_in_333;
wire [161:0] u_ca_in_334;
wire [161:0] u_ca_in_335;
wire [161:0] u_ca_in_336;
wire [161:0] u_ca_in_337;
wire [161:0] u_ca_in_338;
wire [161:0] u_ca_in_339;
wire [161:0] u_ca_in_340;
wire [161:0] u_ca_in_341;
wire [161:0] u_ca_in_342;
wire [161:0] u_ca_in_343;
wire [161:0] u_ca_in_344;
wire [161:0] u_ca_in_345;
wire [161:0] u_ca_in_346;
wire [161:0] u_ca_in_347;
wire [161:0] u_ca_in_348;
wire [161:0] u_ca_in_349;
wire [161:0] u_ca_in_350;
wire [161:0] u_ca_in_351;
wire [161:0] u_ca_in_352;
wire [161:0] u_ca_in_353;
wire [161:0] u_ca_in_354;
wire [161:0] u_ca_in_355;
wire [161:0] u_ca_in_356;
wire [161:0] u_ca_in_357;
wire [161:0] u_ca_in_358;
wire [161:0] u_ca_in_359;
wire [161:0] u_ca_in_360;
wire [161:0] u_ca_in_361;
wire [161:0] u_ca_in_362;
wire [161:0] u_ca_in_363;
wire [161:0] u_ca_in_364;
wire [161:0] u_ca_in_365;
wire [161:0] u_ca_in_366;
wire [161:0] u_ca_in_367;
wire [161:0] u_ca_in_368;
wire [161:0] u_ca_in_369;
wire [161:0] u_ca_in_370;
wire [161:0] u_ca_in_371;
wire [161:0] u_ca_in_372;
wire [161:0] u_ca_in_373;
wire [161:0] u_ca_in_374;
wire [161:0] u_ca_in_375;
wire [161:0] u_ca_in_376;
wire [161:0] u_ca_in_377;
wire [161:0] u_ca_in_378;
wire [161:0] u_ca_in_379;
wire [161:0] u_ca_in_380;
wire [161:0] u_ca_in_381;
wire [161:0] u_ca_in_382;
wire [161:0] u_ca_in_383;
wire [161:0] u_ca_in_384;
wire [161:0] u_ca_in_385;
wire [161:0] u_ca_in_386;
wire [161:0] u_ca_in_387;
wire [161:0] u_ca_in_388;
wire [161:0] u_ca_in_389;
wire [161:0] u_ca_in_390;
wire [161:0] u_ca_in_391;
wire [161:0] u_ca_in_392;
wire [161:0] u_ca_in_393;
wire [161:0] u_ca_in_394;
wire [161:0] u_ca_in_395;
wire [161:0] u_ca_in_396;
wire [161:0] u_ca_in_397;
wire [161:0] u_ca_in_398;
wire [161:0] u_ca_in_399;
wire [161:0] u_ca_in_400;
wire [161:0] u_ca_in_401;
wire [161:0] u_ca_in_402;
wire [161:0] u_ca_in_403;
wire [161:0] u_ca_in_404;
wire [161:0] u_ca_in_405;
wire [161:0] u_ca_in_406;
wire [161:0] u_ca_in_407;
wire [161:0] u_ca_in_408;
wire [161:0] u_ca_in_409;
wire [161:0] u_ca_in_410;
wire [161:0] u_ca_in_411;
wire [161:0] u_ca_in_412;
wire [161:0] u_ca_in_413;
wire [161:0] u_ca_in_414;
wire [161:0] u_ca_in_415;
wire [161:0] u_ca_in_416;
wire [161:0] u_ca_in_417;
wire [161:0] u_ca_in_418;
wire [161:0] u_ca_in_419;
wire [161:0] u_ca_in_420;
wire [161:0] u_ca_in_421;
wire [161:0] u_ca_in_422;
wire [161:0] u_ca_in_423;
wire [161:0] u_ca_in_424;
wire [161:0] u_ca_in_425;
wire [161:0] u_ca_in_426;
wire [161:0] u_ca_in_427;
wire [161:0] u_ca_in_428;
wire [161:0] u_ca_in_429;
wire [161:0] u_ca_in_430;
wire [161:0] u_ca_in_431;
wire [161:0] u_ca_in_432;
wire [161:0] u_ca_in_433;
wire [161:0] u_ca_in_434;
wire [161:0] u_ca_in_435;
wire [161:0] u_ca_in_436;
wire [161:0] u_ca_in_437;
wire [161:0] u_ca_in_438;
wire [161:0] u_ca_in_439;
wire [161:0] u_ca_in_440;
wire [161:0] u_ca_in_441;
wire [161:0] u_ca_in_442;
wire [161:0] u_ca_in_443;
wire [161:0] u_ca_in_444;
wire [161:0] u_ca_in_445;
wire [161:0] u_ca_in_446;
wire [161:0] u_ca_in_447;
wire [161:0] u_ca_in_448;
wire [161:0] u_ca_in_449;
wire [161:0] u_ca_in_450;
wire [161:0] u_ca_in_451;
wire [161:0] u_ca_in_452;
wire [161:0] u_ca_in_453;
wire [161:0] u_ca_in_454;
wire [161:0] u_ca_in_455;
wire [161:0] u_ca_in_456;
wire [161:0] u_ca_in_457;
wire [161:0] u_ca_in_458;
wire [161:0] u_ca_in_459;
wire [161:0] u_ca_in_460;
wire [161:0] u_ca_in_461;
wire [161:0] u_ca_in_462;
wire [161:0] u_ca_in_463;
wire [161:0] u_ca_in_464;
wire [161:0] u_ca_in_465;
wire [161:0] u_ca_in_466;
wire [161:0] u_ca_in_467;
wire [161:0] u_ca_in_468;
wire [161:0] u_ca_in_469;
wire [161:0] u_ca_in_470;
wire [161:0] u_ca_in_471;
wire [161:0] u_ca_in_472;
wire [161:0] u_ca_in_473;
wire [161:0] u_ca_in_474;
wire [161:0] u_ca_in_475;
wire [161:0] u_ca_in_476;
wire [161:0] u_ca_in_477;
wire [161:0] u_ca_in_478;
wire [161:0] u_ca_in_479;
wire [161:0] u_ca_in_480;
wire [161:0] u_ca_in_481;
wire [161:0] u_ca_in_482;
wire [161:0] u_ca_in_483;
wire [161:0] u_ca_in_484;
wire [161:0] u_ca_in_485;
wire [161:0] u_ca_in_486;
wire [161:0] u_ca_in_487;
wire [161:0] u_ca_in_488;
wire [161:0] u_ca_in_489;
wire [161:0] u_ca_in_490;
wire [161:0] u_ca_in_491;
wire [161:0] u_ca_in_492;
wire [161:0] u_ca_in_493;
wire [161:0] u_ca_in_494;
wire [161:0] u_ca_in_495;
wire [161:0] u_ca_in_496;
wire [161:0] u_ca_in_497;
wire [161:0] u_ca_in_498;
wire [161:0] u_ca_in_499;
wire [161:0] u_ca_in_500;
wire [161:0] u_ca_in_501;
wire [161:0] u_ca_in_502;
wire [161:0] u_ca_in_503;
wire [161:0] u_ca_in_504;
wire [161:0] u_ca_in_505;
wire [161:0] u_ca_in_506;
wire [161:0] u_ca_in_507;
wire [161:0] u_ca_in_508;
wire [161:0] u_ca_in_509;
wire [161:0] u_ca_in_510;
wire [161:0] u_ca_in_511;
wire [161:0] u_ca_in_512;
wire [161:0] u_ca_in_513;
wire [161:0] u_ca_in_514;
wire [161:0] u_ca_in_515;
wire [161:0] u_ca_in_516;
wire [161:0] u_ca_in_517;
wire [161:0] u_ca_in_518;
wire [161:0] u_ca_in_519;
wire [161:0] u_ca_in_520;
wire [161:0] u_ca_in_521;
wire [161:0] u_ca_in_522;
wire [161:0] u_ca_in_523;
wire [161:0] u_ca_in_524;
wire [161:0] u_ca_in_525;
wire [161:0] u_ca_in_526;
wire [161:0] u_ca_in_527;
wire [161:0] u_ca_in_528;
wire [161:0] u_ca_in_529;
wire [161:0] u_ca_in_530;
wire [161:0] u_ca_in_531;
wire [161:0] u_ca_in_532;
wire [161:0] u_ca_in_533;
wire [161:0] u_ca_in_534;
wire [161:0] u_ca_in_535;
wire [161:0] u_ca_in_536;
wire [161:0] u_ca_in_537;
wire [161:0] u_ca_in_538;
wire [161:0] u_ca_in_539;
wire [161:0] u_ca_in_540;
wire [161:0] u_ca_in_541;
wire [161:0] u_ca_in_542;
wire [161:0] u_ca_in_543;
wire [161:0] u_ca_in_544;
wire [161:0] u_ca_in_545;
wire [161:0] u_ca_in_546;
wire [161:0] u_ca_in_547;
wire [161:0] u_ca_in_548;
wire [161:0] u_ca_in_549;
wire [161:0] u_ca_in_550;
wire [161:0] u_ca_in_551;
wire [161:0] u_ca_in_552;
wire [161:0] u_ca_in_553;
wire [161:0] u_ca_in_554;
wire [161:0] u_ca_in_555;
wire [161:0] u_ca_in_556;
wire [161:0] u_ca_in_557;
wire [161:0] u_ca_in_558;
wire [161:0] u_ca_in_559;
wire [161:0] u_ca_in_560;
wire [161:0] u_ca_in_561;
wire [161:0] u_ca_in_562;
wire [161:0] u_ca_in_563;
wire [161:0] u_ca_in_564;
wire [161:0] u_ca_in_565;
wire [161:0] u_ca_in_566;
wire [161:0] u_ca_in_567;
wire [161:0] u_ca_in_568;
wire [161:0] u_ca_in_569;
wire [161:0] u_ca_in_570;
wire [161:0] u_ca_in_571;
wire [161:0] u_ca_in_572;
wire [161:0] u_ca_in_573;
wire [161:0] u_ca_in_574;
wire [161:0] u_ca_in_575;
wire [161:0] u_ca_in_576;
wire [161:0] u_ca_in_577;
wire [161:0] u_ca_in_578;
wire [161:0] u_ca_in_579;
wire [161:0] u_ca_in_580;
wire [161:0] u_ca_in_581;
wire [161:0] u_ca_in_582;
wire [161:0] u_ca_in_583;
wire [161:0] u_ca_in_584;
wire [161:0] u_ca_in_585;
wire [161:0] u_ca_in_586;
wire [161:0] u_ca_in_587;
wire [161:0] u_ca_in_588;
wire [161:0] u_ca_in_589;
wire [161:0] u_ca_in_590;
wire [161:0] u_ca_in_591;
wire [161:0] u_ca_in_592;
wire [161:0] u_ca_in_593;
wire [161:0] u_ca_in_594;
wire [161:0] u_ca_in_595;
wire [161:0] u_ca_in_596;
wire [161:0] u_ca_in_597;
wire [161:0] u_ca_in_598;
wire [161:0] u_ca_in_599;
wire [161:0] u_ca_in_600;
wire [161:0] u_ca_in_601;
wire [161:0] u_ca_in_602;
wire [161:0] u_ca_in_603;
wire [161:0] u_ca_in_604;
wire [161:0] u_ca_in_605;
wire [161:0] u_ca_in_606;
wire [161:0] u_ca_in_607;
wire [161:0] u_ca_in_608;
wire [161:0] u_ca_in_609;
wire [161:0] u_ca_in_610;
wire [161:0] u_ca_in_611;
wire [161:0] u_ca_in_612;
wire [161:0] u_ca_in_613;
wire [161:0] u_ca_in_614;
wire [161:0] u_ca_in_615;
wire [161:0] u_ca_in_616;
wire [161:0] u_ca_in_617;
wire [161:0] u_ca_in_618;
wire [161:0] u_ca_in_619;
wire [161:0] u_ca_in_620;
wire [161:0] u_ca_in_621;
wire [161:0] u_ca_in_622;
wire [161:0] u_ca_in_623;
wire [161:0] u_ca_in_624;
wire [161:0] u_ca_in_625;
wire [161:0] u_ca_in_626;
wire [161:0] u_ca_in_627;
wire [161:0] u_ca_in_628;
wire [161:0] u_ca_in_629;
wire [161:0] u_ca_in_630;
wire [161:0] u_ca_in_631;
wire [161:0] u_ca_in_632;
wire [161:0] u_ca_in_633;
wire [161:0] u_ca_in_634;
wire [161:0] u_ca_in_635;
wire [161:0] u_ca_in_636;
wire [161:0] u_ca_in_637;
wire [161:0] u_ca_in_638;
wire [161:0] u_ca_in_639;
wire [161:0] u_ca_in_640;
wire [161:0] u_ca_in_641;
wire [161:0] u_ca_in_642;
wire [161:0] u_ca_in_643;
wire [161:0] u_ca_in_644;
wire [161:0] u_ca_in_645;
wire [161:0] u_ca_in_646;
wire [161:0] u_ca_in_647;
wire [161:0] u_ca_in_648;
wire [161:0] u_ca_in_649;
wire [161:0] u_ca_in_650;
wire [161:0] u_ca_in_651;
wire [161:0] u_ca_in_652;
wire [161:0] u_ca_in_653;
wire [161:0] u_ca_in_654;
wire [161:0] u_ca_in_655;
wire [161:0] u_ca_in_656;
wire [161:0] u_ca_in_657;
wire [161:0] u_ca_in_658;
wire [161:0] u_ca_in_659;
wire [161:0] u_ca_in_660;
wire [161:0] u_ca_in_661;
wire [161:0] u_ca_in_662;
wire [161:0] u_ca_in_663;
wire [161:0] u_ca_in_664;
wire [161:0] u_ca_in_665;
wire [161:0] u_ca_in_666;
wire [161:0] u_ca_in_667;
wire [161:0] u_ca_in_668;
wire [161:0] u_ca_in_669;
wire [161:0] u_ca_in_670;
wire [161:0] u_ca_in_671;
wire [161:0] u_ca_in_672;
wire [161:0] u_ca_in_673;
wire [161:0] u_ca_in_674;
wire [161:0] u_ca_in_675;
wire [161:0] u_ca_in_676;
wire [161:0] u_ca_in_677;
wire [161:0] u_ca_in_678;
wire [161:0] u_ca_in_679;
wire [161:0] u_ca_in_680;
wire [161:0] u_ca_in_681;
wire [161:0] u_ca_in_682;
wire [161:0] u_ca_in_683;
wire [161:0] u_ca_in_684;
wire [161:0] u_ca_in_685;
wire [161:0] u_ca_in_686;
wire [161:0] u_ca_in_687;
wire [161:0] u_ca_in_688;
wire [161:0] u_ca_in_689;
wire [161:0] u_ca_in_690;
wire [161:0] u_ca_in_691;
wire [161:0] u_ca_in_692;
wire [161:0] u_ca_in_693;
wire [161:0] u_ca_in_694;
wire [161:0] u_ca_in_695;
wire [161:0] u_ca_in_696;
wire [161:0] u_ca_in_697;
wire [161:0] u_ca_in_698;
wire [161:0] u_ca_in_699;
wire [161:0] u_ca_in_700;
wire [161:0] u_ca_in_701;
wire [161:0] u_ca_in_702;
wire [161:0] u_ca_in_703;
wire [161:0] u_ca_in_704;
wire [161:0] u_ca_in_705;
wire [161:0] u_ca_in_706;
wire [161:0] u_ca_in_707;
wire [161:0] u_ca_in_708;
wire [161:0] u_ca_in_709;
wire [161:0] u_ca_in_710;
wire [161:0] u_ca_in_711;
wire [161:0] u_ca_in_712;
wire [161:0] u_ca_in_713;
wire [161:0] u_ca_in_714;
wire [161:0] u_ca_in_715;
wire [161:0] u_ca_in_716;
wire [161:0] u_ca_in_717;
wire [161:0] u_ca_in_718;
wire [161:0] u_ca_in_719;
wire [161:0] u_ca_in_720;
wire [161:0] u_ca_in_721;
wire [161:0] u_ca_in_722;
wire [161:0] u_ca_in_723;
wire [161:0] u_ca_in_724;
wire [161:0] u_ca_in_725;
wire [161:0] u_ca_in_726;
wire [161:0] u_ca_in_727;
wire [161:0] u_ca_in_728;
wire [161:0] u_ca_in_729;
wire [161:0] u_ca_in_730;
wire [161:0] u_ca_in_731;
wire [161:0] u_ca_in_732;
wire [161:0] u_ca_in_733;
wire [161:0] u_ca_in_734;
wire [161:0] u_ca_in_735;
wire [161:0] u_ca_in_736;
wire [161:0] u_ca_in_737;
wire [161:0] u_ca_in_738;
wire [161:0] u_ca_in_739;
wire [161:0] u_ca_in_740;
wire [161:0] u_ca_in_741;
wire [161:0] u_ca_in_742;
wire [161:0] u_ca_in_743;
wire [161:0] u_ca_in_744;
wire [161:0] u_ca_in_745;
wire [161:0] u_ca_in_746;
wire [161:0] u_ca_in_747;
wire [161:0] u_ca_in_748;
wire [161:0] u_ca_in_749;
wire [161:0] u_ca_in_750;
wire [161:0] u_ca_in_751;
wire [161:0] u_ca_in_752;
wire [161:0] u_ca_in_753;
wire [161:0] u_ca_in_754;
wire [161:0] u_ca_in_755;
wire [161:0] u_ca_in_756;
wire [161:0] u_ca_in_757;
wire [161:0] u_ca_in_758;
wire [161:0] u_ca_in_759;
wire [161:0] u_ca_in_760;
wire [161:0] u_ca_in_761;
wire [161:0] u_ca_in_762;
wire [161:0] u_ca_in_763;
wire [161:0] u_ca_in_764;
wire [161:0] u_ca_in_765;
wire [161:0] u_ca_in_766;
wire [161:0] u_ca_in_767;
wire [161:0] u_ca_in_768;
wire [161:0] u_ca_in_769;
wire [161:0] u_ca_in_770;
wire [161:0] u_ca_in_771;
wire [161:0] u_ca_in_772;
wire [161:0] u_ca_in_773;
wire [161:0] u_ca_in_774;
wire [161:0] u_ca_in_775;
wire [161:0] u_ca_in_776;
wire [161:0] u_ca_in_777;
wire [161:0] u_ca_in_778;
wire [161:0] u_ca_in_779;
wire [161:0] u_ca_in_780;
wire [161:0] u_ca_in_781;
wire [161:0] u_ca_in_782;
wire [161:0] u_ca_in_783;
wire [161:0] u_ca_in_784;
wire [161:0] u_ca_in_785;
wire [161:0] u_ca_in_786;
wire [161:0] u_ca_in_787;
wire [161:0] u_ca_in_788;
wire [161:0] u_ca_in_789;
wire [161:0] u_ca_in_790;
wire [161:0] u_ca_in_791;
wire [161:0] u_ca_in_792;
wire [161:0] u_ca_in_793;
wire [161:0] u_ca_in_794;
wire [161:0] u_ca_in_795;
wire [161:0] u_ca_in_796;
wire [161:0] u_ca_in_797;
wire [161:0] u_ca_in_798;
wire [161:0] u_ca_in_799;
wire [161:0] u_ca_in_800;
wire [161:0] u_ca_in_801;
wire [161:0] u_ca_in_802;
wire [161:0] u_ca_in_803;
wire [161:0] u_ca_in_804;
wire [161:0] u_ca_in_805;
wire [161:0] u_ca_in_806;
wire [161:0] u_ca_in_807;
wire [161:0] u_ca_in_808;
wire [161:0] u_ca_in_809;
wire [161:0] u_ca_in_810;
wire [161:0] u_ca_in_811;
wire [161:0] u_ca_in_812;
wire [161:0] u_ca_in_813;
wire [161:0] u_ca_in_814;
wire [161:0] u_ca_in_815;
wire [161:0] u_ca_in_816;
wire [161:0] u_ca_in_817;
wire [161:0] u_ca_in_818;
wire [161:0] u_ca_in_819;
wire [161:0] u_ca_in_820;
wire [161:0] u_ca_in_821;
wire [161:0] u_ca_in_822;
wire [161:0] u_ca_in_823;
wire [161:0] u_ca_in_824;
wire [161:0] u_ca_in_825;
wire [161:0] u_ca_in_826;
wire [161:0] u_ca_in_827;
wire [161:0] u_ca_in_828;
wire [161:0] u_ca_in_829;
wire [161:0] u_ca_in_830;
wire [161:0] u_ca_in_831;
wire [161:0] u_ca_in_832;
wire [161:0] u_ca_in_833;
wire [161:0] u_ca_in_834;
wire [161:0] u_ca_in_835;
wire [161:0] u_ca_in_836;
wire [161:0] u_ca_in_837;
wire [161:0] u_ca_in_838;
wire [161:0] u_ca_in_839;
wire [161:0] u_ca_in_840;
wire [161:0] u_ca_in_841;
wire [161:0] u_ca_in_842;
wire [161:0] u_ca_in_843;
wire [161:0] u_ca_in_844;
wire [161:0] u_ca_in_845;
wire [161:0] u_ca_in_846;
wire [161:0] u_ca_in_847;
wire [161:0] u_ca_in_848;
wire [161:0] u_ca_in_849;
wire [161:0] u_ca_in_850;
wire [161:0] u_ca_in_851;
wire [161:0] u_ca_in_852;
wire [161:0] u_ca_in_853;
wire [161:0] u_ca_in_854;
wire [161:0] u_ca_in_855;
wire [161:0] u_ca_in_856;
wire [161:0] u_ca_in_857;
wire [161:0] u_ca_in_858;
wire [161:0] u_ca_in_859;
wire [161:0] u_ca_in_860;
wire [161:0] u_ca_in_861;
wire [161:0] u_ca_in_862;
wire [161:0] u_ca_in_863;
wire [161:0] u_ca_in_864;
wire [161:0] u_ca_in_865;
wire [161:0] u_ca_in_866;
wire [161:0] u_ca_in_867;
wire [161:0] u_ca_in_868;
wire [161:0] u_ca_in_869;
wire [161:0] u_ca_in_870;
wire [161:0] u_ca_in_871;
wire [161:0] u_ca_in_872;
wire [161:0] u_ca_in_873;
wire [161:0] u_ca_in_874;
wire [161:0] u_ca_in_875;
wire [161:0] u_ca_in_876;
wire [161:0] u_ca_in_877;
wire [161:0] u_ca_in_878;
wire [161:0] u_ca_in_879;
wire [161:0] u_ca_in_880;
wire [161:0] u_ca_in_881;
wire [161:0] u_ca_in_882;
wire [161:0] u_ca_in_883;
wire [161:0] u_ca_in_884;
wire [161:0] u_ca_in_885;
wire [161:0] u_ca_in_886;
wire [161:0] u_ca_in_887;
wire [161:0] u_ca_in_888;
wire [161:0] u_ca_in_889;
wire [161:0] u_ca_in_890;
wire [161:0] u_ca_in_891;
wire [161:0] u_ca_in_892;
wire [161:0] u_ca_in_893;
wire [161:0] u_ca_in_894;
wire [161:0] u_ca_in_895;
wire [161:0] u_ca_in_896;
wire [161:0] u_ca_in_897;
wire [161:0] u_ca_in_898;
wire [161:0] u_ca_in_899;
wire [161:0] u_ca_in_900;
wire [161:0] u_ca_in_901;
wire [161:0] u_ca_in_902;
wire [161:0] u_ca_in_903;
wire [161:0] u_ca_in_904;
wire [161:0] u_ca_in_905;
wire [161:0] u_ca_in_906;
wire [161:0] u_ca_in_907;
wire [161:0] u_ca_in_908;
wire [161:0] u_ca_in_909;
wire [161:0] u_ca_in_910;
wire [161:0] u_ca_in_911;
wire [161:0] u_ca_in_912;
wire [161:0] u_ca_in_913;
wire [161:0] u_ca_in_914;
wire [161:0] u_ca_in_915;
wire [161:0] u_ca_in_916;
wire [161:0] u_ca_in_917;
wire [161:0] u_ca_in_918;
wire [161:0] u_ca_in_919;
wire [161:0] u_ca_in_920;
wire [161:0] u_ca_in_921;
wire [161:0] u_ca_in_922;
wire [161:0] u_ca_in_923;
wire [161:0] u_ca_in_924;
wire [161:0] u_ca_in_925;
wire [161:0] u_ca_in_926;
wire [161:0] u_ca_in_927;
wire [161:0] u_ca_in_928;
wire [161:0] u_ca_in_929;
wire [161:0] u_ca_in_930;
wire [161:0] u_ca_in_931;
wire [161:0] u_ca_in_932;
wire [161:0] u_ca_in_933;
wire [161:0] u_ca_in_934;
wire [161:0] u_ca_in_935;
wire [161:0] u_ca_in_936;
wire [161:0] u_ca_in_937;
wire [161:0] u_ca_in_938;
wire [161:0] u_ca_in_939;
wire [161:0] u_ca_in_940;
wire [161:0] u_ca_in_941;
wire [161:0] u_ca_in_942;
wire [161:0] u_ca_in_943;
wire [161:0] u_ca_in_944;
wire [161:0] u_ca_in_945;
wire [161:0] u_ca_in_946;
wire [161:0] u_ca_in_947;
wire [161:0] u_ca_in_948;
wire [161:0] u_ca_in_949;
wire [161:0] u_ca_in_950;
wire [161:0] u_ca_in_951;
wire [161:0] u_ca_in_952;
wire [161:0] u_ca_in_953;
wire [161:0] u_ca_in_954;
wire [161:0] u_ca_in_955;
wire [161:0] u_ca_in_956;
wire [161:0] u_ca_in_957;
wire [161:0] u_ca_in_958;
wire [161:0] u_ca_in_959;
wire [161:0] u_ca_in_960;
wire [161:0] u_ca_in_961;
wire [161:0] u_ca_in_962;
wire [161:0] u_ca_in_963;
wire [161:0] u_ca_in_964;
wire [161:0] u_ca_in_965;
wire [161:0] u_ca_in_966;
wire [161:0] u_ca_in_967;
wire [161:0] u_ca_in_968;
wire [161:0] u_ca_in_969;
wire [161:0] u_ca_in_970;
wire [161:0] u_ca_in_971;
wire [161:0] u_ca_in_972;
wire [161:0] u_ca_in_973;
wire [161:0] u_ca_in_974;
wire [161:0] u_ca_in_975;
wire [161:0] u_ca_in_976;
wire [161:0] u_ca_in_977;
wire [161:0] u_ca_in_978;
wire [161:0] u_ca_in_979;
wire [161:0] u_ca_in_980;
wire [161:0] u_ca_in_981;
wire [161:0] u_ca_in_982;
wire [161:0] u_ca_in_983;
wire [161:0] u_ca_in_984;
wire [161:0] u_ca_in_985;
wire [161:0] u_ca_in_986;
wire [161:0] u_ca_in_987;
wire [161:0] u_ca_in_988;
wire [161:0] u_ca_in_989;
wire [161:0] u_ca_in_990;
wire [161:0] u_ca_in_991;
wire [161:0] u_ca_in_992;
wire [161:0] u_ca_in_993;
wire [161:0] u_ca_in_994;
wire [161:0] u_ca_in_995;
wire [161:0] u_ca_in_996;
wire [161:0] u_ca_in_997;
wire [161:0] u_ca_in_998;
wire [161:0] u_ca_in_999;
wire [161:0] u_ca_in_1000;
wire [161:0] u_ca_in_1001;
wire [161:0] u_ca_in_1002;
wire [161:0] u_ca_in_1003;
wire [161:0] u_ca_in_1004;
wire [161:0] u_ca_in_1005;
wire [161:0] u_ca_in_1006;
wire [161:0] u_ca_in_1007;
wire [161:0] u_ca_in_1008;
wire [161:0] u_ca_in_1009;
wire [161:0] u_ca_in_1010;
wire [161:0] u_ca_in_1011;
wire [161:0] u_ca_in_1012;
wire [161:0] u_ca_in_1013;
wire [161:0] u_ca_in_1014;
wire [161:0] u_ca_in_1015;
wire [161:0] u_ca_in_1016;
wire [161:0] u_ca_in_1017;
wire [161:0] u_ca_in_1018;
wire [161:0] u_ca_in_1019;
wire [161:0] u_ca_in_1020;
wire [161:0] u_ca_in_1021;
wire [161:0] u_ca_in_1022;
wire [161:0] u_ca_in_1023;
wire [161:0] u_ca_in_1024;
wire [161:0] u_ca_in_1025;
wire [161:0] u_ca_in_1026;
wire [47:0] u_ca_out_0;
wire [47:0] u_ca_out_1;
wire [47:0] u_ca_out_2;
wire [47:0] u_ca_out_3;
wire [47:0] u_ca_out_4;
wire [47:0] u_ca_out_5;
wire [47:0] u_ca_out_6;
wire [47:0] u_ca_out_7;
wire [47:0] u_ca_out_8;
wire [47:0] u_ca_out_9;
wire [47:0] u_ca_out_10;
wire [47:0] u_ca_out_11;
wire [47:0] u_ca_out_12;
wire [47:0] u_ca_out_13;
wire [47:0] u_ca_out_14;
wire [47:0] u_ca_out_15;
wire [47:0] u_ca_out_16;
wire [47:0] u_ca_out_17;
wire [47:0] u_ca_out_18;
wire [47:0] u_ca_out_19;
wire [47:0] u_ca_out_20;
wire [47:0] u_ca_out_21;
wire [47:0] u_ca_out_22;
wire [47:0] u_ca_out_23;
wire [47:0] u_ca_out_24;
wire [47:0] u_ca_out_25;
wire [47:0] u_ca_out_26;
wire [47:0] u_ca_out_27;
wire [47:0] u_ca_out_28;
wire [47:0] u_ca_out_29;
wire [47:0] u_ca_out_30;
wire [47:0] u_ca_out_31;
wire [47:0] u_ca_out_32;
wire [47:0] u_ca_out_33;
wire [47:0] u_ca_out_34;
wire [47:0] u_ca_out_35;
wire [47:0] u_ca_out_36;
wire [47:0] u_ca_out_37;
wire [47:0] u_ca_out_38;
wire [47:0] u_ca_out_39;
wire [47:0] u_ca_out_40;
wire [47:0] u_ca_out_41;
wire [47:0] u_ca_out_42;
wire [47:0] u_ca_out_43;
wire [47:0] u_ca_out_44;
wire [47:0] u_ca_out_45;
wire [47:0] u_ca_out_46;
wire [47:0] u_ca_out_47;
wire [47:0] u_ca_out_48;
wire [47:0] u_ca_out_49;
wire [47:0] u_ca_out_50;
wire [47:0] u_ca_out_51;
wire [47:0] u_ca_out_52;
wire [47:0] u_ca_out_53;
wire [47:0] u_ca_out_54;
wire [47:0] u_ca_out_55;
wire [47:0] u_ca_out_56;
wire [47:0] u_ca_out_57;
wire [47:0] u_ca_out_58;
wire [47:0] u_ca_out_59;
wire [47:0] u_ca_out_60;
wire [47:0] u_ca_out_61;
wire [47:0] u_ca_out_62;
wire [47:0] u_ca_out_63;
wire [47:0] u_ca_out_64;
wire [47:0] u_ca_out_65;
wire [47:0] u_ca_out_66;
wire [47:0] u_ca_out_67;
wire [47:0] u_ca_out_68;
wire [47:0] u_ca_out_69;
wire [47:0] u_ca_out_70;
wire [47:0] u_ca_out_71;
wire [47:0] u_ca_out_72;
wire [47:0] u_ca_out_73;
wire [47:0] u_ca_out_74;
wire [47:0] u_ca_out_75;
wire [47:0] u_ca_out_76;
wire [47:0] u_ca_out_77;
wire [47:0] u_ca_out_78;
wire [47:0] u_ca_out_79;
wire [47:0] u_ca_out_80;
wire [47:0] u_ca_out_81;
wire [47:0] u_ca_out_82;
wire [47:0] u_ca_out_83;
wire [47:0] u_ca_out_84;
wire [47:0] u_ca_out_85;
wire [47:0] u_ca_out_86;
wire [47:0] u_ca_out_87;
wire [47:0] u_ca_out_88;
wire [47:0] u_ca_out_89;
wire [47:0] u_ca_out_90;
wire [47:0] u_ca_out_91;
wire [47:0] u_ca_out_92;
wire [47:0] u_ca_out_93;
wire [47:0] u_ca_out_94;
wire [47:0] u_ca_out_95;
wire [47:0] u_ca_out_96;
wire [47:0] u_ca_out_97;
wire [47:0] u_ca_out_98;
wire [47:0] u_ca_out_99;
wire [47:0] u_ca_out_100;
wire [47:0] u_ca_out_101;
wire [47:0] u_ca_out_102;
wire [47:0] u_ca_out_103;
wire [47:0] u_ca_out_104;
wire [47:0] u_ca_out_105;
wire [47:0] u_ca_out_106;
wire [47:0] u_ca_out_107;
wire [47:0] u_ca_out_108;
wire [47:0] u_ca_out_109;
wire [47:0] u_ca_out_110;
wire [47:0] u_ca_out_111;
wire [47:0] u_ca_out_112;
wire [47:0] u_ca_out_113;
wire [47:0] u_ca_out_114;
wire [47:0] u_ca_out_115;
wire [47:0] u_ca_out_116;
wire [47:0] u_ca_out_117;
wire [47:0] u_ca_out_118;
wire [47:0] u_ca_out_119;
wire [47:0] u_ca_out_120;
wire [47:0] u_ca_out_121;
wire [47:0] u_ca_out_122;
wire [47:0] u_ca_out_123;
wire [47:0] u_ca_out_124;
wire [47:0] u_ca_out_125;
wire [47:0] u_ca_out_126;
wire [47:0] u_ca_out_127;
wire [47:0] u_ca_out_128;
wire [47:0] u_ca_out_129;
wire [47:0] u_ca_out_130;
wire [47:0] u_ca_out_131;
wire [47:0] u_ca_out_132;
wire [47:0] u_ca_out_133;
wire [47:0] u_ca_out_134;
wire [47:0] u_ca_out_135;
wire [47:0] u_ca_out_136;
wire [47:0] u_ca_out_137;
wire [47:0] u_ca_out_138;
wire [47:0] u_ca_out_139;
wire [47:0] u_ca_out_140;
wire [47:0] u_ca_out_141;
wire [47:0] u_ca_out_142;
wire [47:0] u_ca_out_143;
wire [47:0] u_ca_out_144;
wire [47:0] u_ca_out_145;
wire [47:0] u_ca_out_146;
wire [47:0] u_ca_out_147;
wire [47:0] u_ca_out_148;
wire [47:0] u_ca_out_149;
wire [47:0] u_ca_out_150;
wire [47:0] u_ca_out_151;
wire [47:0] u_ca_out_152;
wire [47:0] u_ca_out_153;
wire [47:0] u_ca_out_154;
wire [47:0] u_ca_out_155;
wire [47:0] u_ca_out_156;
wire [47:0] u_ca_out_157;
wire [47:0] u_ca_out_158;
wire [47:0] u_ca_out_159;
wire [47:0] u_ca_out_160;
wire [47:0] u_ca_out_161;
wire [47:0] u_ca_out_162;
wire [47:0] u_ca_out_163;
wire [47:0] u_ca_out_164;
wire [47:0] u_ca_out_165;
wire [47:0] u_ca_out_166;
wire [47:0] u_ca_out_167;
wire [47:0] u_ca_out_168;
wire [47:0] u_ca_out_169;
wire [47:0] u_ca_out_170;
wire [47:0] u_ca_out_171;
wire [47:0] u_ca_out_172;
wire [47:0] u_ca_out_173;
wire [47:0] u_ca_out_174;
wire [47:0] u_ca_out_175;
wire [47:0] u_ca_out_176;
wire [47:0] u_ca_out_177;
wire [47:0] u_ca_out_178;
wire [47:0] u_ca_out_179;
wire [47:0] u_ca_out_180;
wire [47:0] u_ca_out_181;
wire [47:0] u_ca_out_182;
wire [47:0] u_ca_out_183;
wire [47:0] u_ca_out_184;
wire [47:0] u_ca_out_185;
wire [47:0] u_ca_out_186;
wire [47:0] u_ca_out_187;
wire [47:0] u_ca_out_188;
wire [47:0] u_ca_out_189;
wire [47:0] u_ca_out_190;
wire [47:0] u_ca_out_191;
wire [47:0] u_ca_out_192;
wire [47:0] u_ca_out_193;
wire [47:0] u_ca_out_194;
wire [47:0] u_ca_out_195;
wire [47:0] u_ca_out_196;
wire [47:0] u_ca_out_197;
wire [47:0] u_ca_out_198;
wire [47:0] u_ca_out_199;
wire [47:0] u_ca_out_200;
wire [47:0] u_ca_out_201;
wire [47:0] u_ca_out_202;
wire [47:0] u_ca_out_203;
wire [47:0] u_ca_out_204;
wire [47:0] u_ca_out_205;
wire [47:0] u_ca_out_206;
wire [47:0] u_ca_out_207;
wire [47:0] u_ca_out_208;
wire [47:0] u_ca_out_209;
wire [47:0] u_ca_out_210;
wire [47:0] u_ca_out_211;
wire [47:0] u_ca_out_212;
wire [47:0] u_ca_out_213;
wire [47:0] u_ca_out_214;
wire [47:0] u_ca_out_215;
wire [47:0] u_ca_out_216;
wire [47:0] u_ca_out_217;
wire [47:0] u_ca_out_218;
wire [47:0] u_ca_out_219;
wire [47:0] u_ca_out_220;
wire [47:0] u_ca_out_221;
wire [47:0] u_ca_out_222;
wire [47:0] u_ca_out_223;
wire [47:0] u_ca_out_224;
wire [47:0] u_ca_out_225;
wire [47:0] u_ca_out_226;
wire [47:0] u_ca_out_227;
wire [47:0] u_ca_out_228;
wire [47:0] u_ca_out_229;
wire [47:0] u_ca_out_230;
wire [47:0] u_ca_out_231;
wire [47:0] u_ca_out_232;
wire [47:0] u_ca_out_233;
wire [47:0] u_ca_out_234;
wire [47:0] u_ca_out_235;
wire [47:0] u_ca_out_236;
wire [47:0] u_ca_out_237;
wire [47:0] u_ca_out_238;
wire [47:0] u_ca_out_239;
wire [47:0] u_ca_out_240;
wire [47:0] u_ca_out_241;
wire [47:0] u_ca_out_242;
wire [47:0] u_ca_out_243;
wire [47:0] u_ca_out_244;
wire [47:0] u_ca_out_245;
wire [47:0] u_ca_out_246;
wire [47:0] u_ca_out_247;
wire [47:0] u_ca_out_248;
wire [47:0] u_ca_out_249;
wire [47:0] u_ca_out_250;
wire [47:0] u_ca_out_251;
wire [47:0] u_ca_out_252;
wire [47:0] u_ca_out_253;
wire [47:0] u_ca_out_254;
wire [47:0] u_ca_out_255;
wire [47:0] u_ca_out_256;
wire [47:0] u_ca_out_257;
wire [47:0] u_ca_out_258;
wire [47:0] u_ca_out_259;
wire [47:0] u_ca_out_260;
wire [47:0] u_ca_out_261;
wire [47:0] u_ca_out_262;
wire [47:0] u_ca_out_263;
wire [47:0] u_ca_out_264;
wire [47:0] u_ca_out_265;
wire [47:0] u_ca_out_266;
wire [47:0] u_ca_out_267;
wire [47:0] u_ca_out_268;
wire [47:0] u_ca_out_269;
wire [47:0] u_ca_out_270;
wire [47:0] u_ca_out_271;
wire [47:0] u_ca_out_272;
wire [47:0] u_ca_out_273;
wire [47:0] u_ca_out_274;
wire [47:0] u_ca_out_275;
wire [47:0] u_ca_out_276;
wire [47:0] u_ca_out_277;
wire [47:0] u_ca_out_278;
wire [47:0] u_ca_out_279;
wire [47:0] u_ca_out_280;
wire [47:0] u_ca_out_281;
wire [47:0] u_ca_out_282;
wire [47:0] u_ca_out_283;
wire [47:0] u_ca_out_284;
wire [47:0] u_ca_out_285;
wire [47:0] u_ca_out_286;
wire [47:0] u_ca_out_287;
wire [47:0] u_ca_out_288;
wire [47:0] u_ca_out_289;
wire [47:0] u_ca_out_290;
wire [47:0] u_ca_out_291;
wire [47:0] u_ca_out_292;
wire [47:0] u_ca_out_293;
wire [47:0] u_ca_out_294;
wire [47:0] u_ca_out_295;
wire [47:0] u_ca_out_296;
wire [47:0] u_ca_out_297;
wire [47:0] u_ca_out_298;
wire [47:0] u_ca_out_299;
wire [47:0] u_ca_out_300;
wire [47:0] u_ca_out_301;
wire [47:0] u_ca_out_302;
wire [47:0] u_ca_out_303;
wire [47:0] u_ca_out_304;
wire [47:0] u_ca_out_305;
wire [47:0] u_ca_out_306;
wire [47:0] u_ca_out_307;
wire [47:0] u_ca_out_308;
wire [47:0] u_ca_out_309;
wire [47:0] u_ca_out_310;
wire [47:0] u_ca_out_311;
wire [47:0] u_ca_out_312;
wire [47:0] u_ca_out_313;
wire [47:0] u_ca_out_314;
wire [47:0] u_ca_out_315;
wire [47:0] u_ca_out_316;
wire [47:0] u_ca_out_317;
wire [47:0] u_ca_out_318;
wire [47:0] u_ca_out_319;
wire [47:0] u_ca_out_320;
wire [47:0] u_ca_out_321;
wire [47:0] u_ca_out_322;
wire [47:0] u_ca_out_323;
wire [47:0] u_ca_out_324;
wire [47:0] u_ca_out_325;
wire [47:0] u_ca_out_326;
wire [47:0] u_ca_out_327;
wire [47:0] u_ca_out_328;
wire [47:0] u_ca_out_329;
wire [47:0] u_ca_out_330;
wire [47:0] u_ca_out_331;
wire [47:0] u_ca_out_332;
wire [47:0] u_ca_out_333;
wire [47:0] u_ca_out_334;
wire [47:0] u_ca_out_335;
wire [47:0] u_ca_out_336;
wire [47:0] u_ca_out_337;
wire [47:0] u_ca_out_338;
wire [47:0] u_ca_out_339;
wire [47:0] u_ca_out_340;
wire [47:0] u_ca_out_341;
wire [47:0] u_ca_out_342;
wire [47:0] u_ca_out_343;
wire [47:0] u_ca_out_344;
wire [47:0] u_ca_out_345;
wire [47:0] u_ca_out_346;
wire [47:0] u_ca_out_347;
wire [47:0] u_ca_out_348;
wire [47:0] u_ca_out_349;
wire [47:0] u_ca_out_350;
wire [47:0] u_ca_out_351;
wire [47:0] u_ca_out_352;
wire [47:0] u_ca_out_353;
wire [47:0] u_ca_out_354;
wire [47:0] u_ca_out_355;
wire [47:0] u_ca_out_356;
wire [47:0] u_ca_out_357;
wire [47:0] u_ca_out_358;
wire [47:0] u_ca_out_359;
wire [47:0] u_ca_out_360;
wire [47:0] u_ca_out_361;
wire [47:0] u_ca_out_362;
wire [47:0] u_ca_out_363;
wire [47:0] u_ca_out_364;
wire [47:0] u_ca_out_365;
wire [47:0] u_ca_out_366;
wire [47:0] u_ca_out_367;
wire [47:0] u_ca_out_368;
wire [47:0] u_ca_out_369;
wire [47:0] u_ca_out_370;
wire [47:0] u_ca_out_371;
wire [47:0] u_ca_out_372;
wire [47:0] u_ca_out_373;
wire [47:0] u_ca_out_374;
wire [47:0] u_ca_out_375;
wire [47:0] u_ca_out_376;
wire [47:0] u_ca_out_377;
wire [47:0] u_ca_out_378;
wire [47:0] u_ca_out_379;
wire [47:0] u_ca_out_380;
wire [47:0] u_ca_out_381;
wire [47:0] u_ca_out_382;
wire [47:0] u_ca_out_383;
wire [47:0] u_ca_out_384;
wire [47:0] u_ca_out_385;
wire [47:0] u_ca_out_386;
wire [47:0] u_ca_out_387;
wire [47:0] u_ca_out_388;
wire [47:0] u_ca_out_389;
wire [47:0] u_ca_out_390;
wire [47:0] u_ca_out_391;
wire [47:0] u_ca_out_392;
wire [47:0] u_ca_out_393;
wire [47:0] u_ca_out_394;
wire [47:0] u_ca_out_395;
wire [47:0] u_ca_out_396;
wire [47:0] u_ca_out_397;
wire [47:0] u_ca_out_398;
wire [47:0] u_ca_out_399;
wire [47:0] u_ca_out_400;
wire [47:0] u_ca_out_401;
wire [47:0] u_ca_out_402;
wire [47:0] u_ca_out_403;
wire [47:0] u_ca_out_404;
wire [47:0] u_ca_out_405;
wire [47:0] u_ca_out_406;
wire [47:0] u_ca_out_407;
wire [47:0] u_ca_out_408;
wire [47:0] u_ca_out_409;
wire [47:0] u_ca_out_410;
wire [47:0] u_ca_out_411;
wire [47:0] u_ca_out_412;
wire [47:0] u_ca_out_413;
wire [47:0] u_ca_out_414;
wire [47:0] u_ca_out_415;
wire [47:0] u_ca_out_416;
wire [47:0] u_ca_out_417;
wire [47:0] u_ca_out_418;
wire [47:0] u_ca_out_419;
wire [47:0] u_ca_out_420;
wire [47:0] u_ca_out_421;
wire [47:0] u_ca_out_422;
wire [47:0] u_ca_out_423;
wire [47:0] u_ca_out_424;
wire [47:0] u_ca_out_425;
wire [47:0] u_ca_out_426;
wire [47:0] u_ca_out_427;
wire [47:0] u_ca_out_428;
wire [47:0] u_ca_out_429;
wire [47:0] u_ca_out_430;
wire [47:0] u_ca_out_431;
wire [47:0] u_ca_out_432;
wire [47:0] u_ca_out_433;
wire [47:0] u_ca_out_434;
wire [47:0] u_ca_out_435;
wire [47:0] u_ca_out_436;
wire [47:0] u_ca_out_437;
wire [47:0] u_ca_out_438;
wire [47:0] u_ca_out_439;
wire [47:0] u_ca_out_440;
wire [47:0] u_ca_out_441;
wire [47:0] u_ca_out_442;
wire [47:0] u_ca_out_443;
wire [47:0] u_ca_out_444;
wire [47:0] u_ca_out_445;
wire [47:0] u_ca_out_446;
wire [47:0] u_ca_out_447;
wire [47:0] u_ca_out_448;
wire [47:0] u_ca_out_449;
wire [47:0] u_ca_out_450;
wire [47:0] u_ca_out_451;
wire [47:0] u_ca_out_452;
wire [47:0] u_ca_out_453;
wire [47:0] u_ca_out_454;
wire [47:0] u_ca_out_455;
wire [47:0] u_ca_out_456;
wire [47:0] u_ca_out_457;
wire [47:0] u_ca_out_458;
wire [47:0] u_ca_out_459;
wire [47:0] u_ca_out_460;
wire [47:0] u_ca_out_461;
wire [47:0] u_ca_out_462;
wire [47:0] u_ca_out_463;
wire [47:0] u_ca_out_464;
wire [47:0] u_ca_out_465;
wire [47:0] u_ca_out_466;
wire [47:0] u_ca_out_467;
wire [47:0] u_ca_out_468;
wire [47:0] u_ca_out_469;
wire [47:0] u_ca_out_470;
wire [47:0] u_ca_out_471;
wire [47:0] u_ca_out_472;
wire [47:0] u_ca_out_473;
wire [47:0] u_ca_out_474;
wire [47:0] u_ca_out_475;
wire [47:0] u_ca_out_476;
wire [47:0] u_ca_out_477;
wire [47:0] u_ca_out_478;
wire [47:0] u_ca_out_479;
wire [47:0] u_ca_out_480;
wire [47:0] u_ca_out_481;
wire [47:0] u_ca_out_482;
wire [47:0] u_ca_out_483;
wire [47:0] u_ca_out_484;
wire [47:0] u_ca_out_485;
wire [47:0] u_ca_out_486;
wire [47:0] u_ca_out_487;
wire [47:0] u_ca_out_488;
wire [47:0] u_ca_out_489;
wire [47:0] u_ca_out_490;
wire [47:0] u_ca_out_491;
wire [47:0] u_ca_out_492;
wire [47:0] u_ca_out_493;
wire [47:0] u_ca_out_494;
wire [47:0] u_ca_out_495;
wire [47:0] u_ca_out_496;
wire [47:0] u_ca_out_497;
wire [47:0] u_ca_out_498;
wire [47:0] u_ca_out_499;
wire [47:0] u_ca_out_500;
wire [47:0] u_ca_out_501;
wire [47:0] u_ca_out_502;
wire [47:0] u_ca_out_503;
wire [47:0] u_ca_out_504;
wire [47:0] u_ca_out_505;
wire [47:0] u_ca_out_506;
wire [47:0] u_ca_out_507;
wire [47:0] u_ca_out_508;
wire [47:0] u_ca_out_509;
wire [47:0] u_ca_out_510;
wire [47:0] u_ca_out_511;
wire [47:0] u_ca_out_512;
wire [47:0] u_ca_out_513;
wire [47:0] u_ca_out_514;
wire [47:0] u_ca_out_515;
wire [47:0] u_ca_out_516;
wire [47:0] u_ca_out_517;
wire [47:0] u_ca_out_518;
wire [47:0] u_ca_out_519;
wire [47:0] u_ca_out_520;
wire [47:0] u_ca_out_521;
wire [47:0] u_ca_out_522;
wire [47:0] u_ca_out_523;
wire [47:0] u_ca_out_524;
wire [47:0] u_ca_out_525;
wire [47:0] u_ca_out_526;
wire [47:0] u_ca_out_527;
wire [47:0] u_ca_out_528;
wire [47:0] u_ca_out_529;
wire [47:0] u_ca_out_530;
wire [47:0] u_ca_out_531;
wire [47:0] u_ca_out_532;
wire [47:0] u_ca_out_533;
wire [47:0] u_ca_out_534;
wire [47:0] u_ca_out_535;
wire [47:0] u_ca_out_536;
wire [47:0] u_ca_out_537;
wire [47:0] u_ca_out_538;
wire [47:0] u_ca_out_539;
wire [47:0] u_ca_out_540;
wire [47:0] u_ca_out_541;
wire [47:0] u_ca_out_542;
wire [47:0] u_ca_out_543;
wire [47:0] u_ca_out_544;
wire [47:0] u_ca_out_545;
wire [47:0] u_ca_out_546;
wire [47:0] u_ca_out_547;
wire [47:0] u_ca_out_548;
wire [47:0] u_ca_out_549;
wire [47:0] u_ca_out_550;
wire [47:0] u_ca_out_551;
wire [47:0] u_ca_out_552;
wire [47:0] u_ca_out_553;
wire [47:0] u_ca_out_554;
wire [47:0] u_ca_out_555;
wire [47:0] u_ca_out_556;
wire [47:0] u_ca_out_557;
wire [47:0] u_ca_out_558;
wire [47:0] u_ca_out_559;
wire [47:0] u_ca_out_560;
wire [47:0] u_ca_out_561;
wire [47:0] u_ca_out_562;
wire [47:0] u_ca_out_563;
wire [47:0] u_ca_out_564;
wire [47:0] u_ca_out_565;
wire [47:0] u_ca_out_566;
wire [47:0] u_ca_out_567;
wire [47:0] u_ca_out_568;
wire [47:0] u_ca_out_569;
wire [47:0] u_ca_out_570;
wire [47:0] u_ca_out_571;
wire [47:0] u_ca_out_572;
wire [47:0] u_ca_out_573;
wire [47:0] u_ca_out_574;
wire [47:0] u_ca_out_575;
wire [47:0] u_ca_out_576;
wire [47:0] u_ca_out_577;
wire [47:0] u_ca_out_578;
wire [47:0] u_ca_out_579;
wire [47:0] u_ca_out_580;
wire [47:0] u_ca_out_581;
wire [47:0] u_ca_out_582;
wire [47:0] u_ca_out_583;
wire [47:0] u_ca_out_584;
wire [47:0] u_ca_out_585;
wire [47:0] u_ca_out_586;
wire [47:0] u_ca_out_587;
wire [47:0] u_ca_out_588;
wire [47:0] u_ca_out_589;
wire [47:0] u_ca_out_590;
wire [47:0] u_ca_out_591;
wire [47:0] u_ca_out_592;
wire [47:0] u_ca_out_593;
wire [47:0] u_ca_out_594;
wire [47:0] u_ca_out_595;
wire [47:0] u_ca_out_596;
wire [47:0] u_ca_out_597;
wire [47:0] u_ca_out_598;
wire [47:0] u_ca_out_599;
wire [47:0] u_ca_out_600;
wire [47:0] u_ca_out_601;
wire [47:0] u_ca_out_602;
wire [47:0] u_ca_out_603;
wire [47:0] u_ca_out_604;
wire [47:0] u_ca_out_605;
wire [47:0] u_ca_out_606;
wire [47:0] u_ca_out_607;
wire [47:0] u_ca_out_608;
wire [47:0] u_ca_out_609;
wire [47:0] u_ca_out_610;
wire [47:0] u_ca_out_611;
wire [47:0] u_ca_out_612;
wire [47:0] u_ca_out_613;
wire [47:0] u_ca_out_614;
wire [47:0] u_ca_out_615;
wire [47:0] u_ca_out_616;
wire [47:0] u_ca_out_617;
wire [47:0] u_ca_out_618;
wire [47:0] u_ca_out_619;
wire [47:0] u_ca_out_620;
wire [47:0] u_ca_out_621;
wire [47:0] u_ca_out_622;
wire [47:0] u_ca_out_623;
wire [47:0] u_ca_out_624;
wire [47:0] u_ca_out_625;
wire [47:0] u_ca_out_626;
wire [47:0] u_ca_out_627;
wire [47:0] u_ca_out_628;
wire [47:0] u_ca_out_629;
wire [47:0] u_ca_out_630;
wire [47:0] u_ca_out_631;
wire [47:0] u_ca_out_632;
wire [47:0] u_ca_out_633;
wire [47:0] u_ca_out_634;
wire [47:0] u_ca_out_635;
wire [47:0] u_ca_out_636;
wire [47:0] u_ca_out_637;
wire [47:0] u_ca_out_638;
wire [47:0] u_ca_out_639;
wire [47:0] u_ca_out_640;
wire [47:0] u_ca_out_641;
wire [47:0] u_ca_out_642;
wire [47:0] u_ca_out_643;
wire [47:0] u_ca_out_644;
wire [47:0] u_ca_out_645;
wire [47:0] u_ca_out_646;
wire [47:0] u_ca_out_647;
wire [47:0] u_ca_out_648;
wire [47:0] u_ca_out_649;
wire [47:0] u_ca_out_650;
wire [47:0] u_ca_out_651;
wire [47:0] u_ca_out_652;
wire [47:0] u_ca_out_653;
wire [47:0] u_ca_out_654;
wire [47:0] u_ca_out_655;
wire [47:0] u_ca_out_656;
wire [47:0] u_ca_out_657;
wire [47:0] u_ca_out_658;
wire [47:0] u_ca_out_659;
wire [47:0] u_ca_out_660;
wire [47:0] u_ca_out_661;
wire [47:0] u_ca_out_662;
wire [47:0] u_ca_out_663;
wire [47:0] u_ca_out_664;
wire [47:0] u_ca_out_665;
wire [47:0] u_ca_out_666;
wire [47:0] u_ca_out_667;
wire [47:0] u_ca_out_668;
wire [47:0] u_ca_out_669;
wire [47:0] u_ca_out_670;
wire [47:0] u_ca_out_671;
wire [47:0] u_ca_out_672;
wire [47:0] u_ca_out_673;
wire [47:0] u_ca_out_674;
wire [47:0] u_ca_out_675;
wire [47:0] u_ca_out_676;
wire [47:0] u_ca_out_677;
wire [47:0] u_ca_out_678;
wire [47:0] u_ca_out_679;
wire [47:0] u_ca_out_680;
wire [47:0] u_ca_out_681;
wire [47:0] u_ca_out_682;
wire [47:0] u_ca_out_683;
wire [47:0] u_ca_out_684;
wire [47:0] u_ca_out_685;
wire [47:0] u_ca_out_686;
wire [47:0] u_ca_out_687;
wire [47:0] u_ca_out_688;
wire [47:0] u_ca_out_689;
wire [47:0] u_ca_out_690;
wire [47:0] u_ca_out_691;
wire [47:0] u_ca_out_692;
wire [47:0] u_ca_out_693;
wire [47:0] u_ca_out_694;
wire [47:0] u_ca_out_695;
wire [47:0] u_ca_out_696;
wire [47:0] u_ca_out_697;
wire [47:0] u_ca_out_698;
wire [47:0] u_ca_out_699;
wire [47:0] u_ca_out_700;
wire [47:0] u_ca_out_701;
wire [47:0] u_ca_out_702;
wire [47:0] u_ca_out_703;
wire [47:0] u_ca_out_704;
wire [47:0] u_ca_out_705;
wire [47:0] u_ca_out_706;
wire [47:0] u_ca_out_707;
wire [47:0] u_ca_out_708;
wire [47:0] u_ca_out_709;
wire [47:0] u_ca_out_710;
wire [47:0] u_ca_out_711;
wire [47:0] u_ca_out_712;
wire [47:0] u_ca_out_713;
wire [47:0] u_ca_out_714;
wire [47:0] u_ca_out_715;
wire [47:0] u_ca_out_716;
wire [47:0] u_ca_out_717;
wire [47:0] u_ca_out_718;
wire [47:0] u_ca_out_719;
wire [47:0] u_ca_out_720;
wire [47:0] u_ca_out_721;
wire [47:0] u_ca_out_722;
wire [47:0] u_ca_out_723;
wire [47:0] u_ca_out_724;
wire [47:0] u_ca_out_725;
wire [47:0] u_ca_out_726;
wire [47:0] u_ca_out_727;
wire [47:0] u_ca_out_728;
wire [47:0] u_ca_out_729;
wire [47:0] u_ca_out_730;
wire [47:0] u_ca_out_731;
wire [47:0] u_ca_out_732;
wire [47:0] u_ca_out_733;
wire [47:0] u_ca_out_734;
wire [47:0] u_ca_out_735;
wire [47:0] u_ca_out_736;
wire [47:0] u_ca_out_737;
wire [47:0] u_ca_out_738;
wire [47:0] u_ca_out_739;
wire [47:0] u_ca_out_740;
wire [47:0] u_ca_out_741;
wire [47:0] u_ca_out_742;
wire [47:0] u_ca_out_743;
wire [47:0] u_ca_out_744;
wire [47:0] u_ca_out_745;
wire [47:0] u_ca_out_746;
wire [47:0] u_ca_out_747;
wire [47:0] u_ca_out_748;
wire [47:0] u_ca_out_749;
wire [47:0] u_ca_out_750;
wire [47:0] u_ca_out_751;
wire [47:0] u_ca_out_752;
wire [47:0] u_ca_out_753;
wire [47:0] u_ca_out_754;
wire [47:0] u_ca_out_755;
wire [47:0] u_ca_out_756;
wire [47:0] u_ca_out_757;
wire [47:0] u_ca_out_758;
wire [47:0] u_ca_out_759;
wire [47:0] u_ca_out_760;
wire [47:0] u_ca_out_761;
wire [47:0] u_ca_out_762;
wire [47:0] u_ca_out_763;
wire [47:0] u_ca_out_764;
wire [47:0] u_ca_out_765;
wire [47:0] u_ca_out_766;
wire [47:0] u_ca_out_767;
wire [47:0] u_ca_out_768;
wire [47:0] u_ca_out_769;
wire [47:0] u_ca_out_770;
wire [47:0] u_ca_out_771;
wire [47:0] u_ca_out_772;
wire [47:0] u_ca_out_773;
wire [47:0] u_ca_out_774;
wire [47:0] u_ca_out_775;
wire [47:0] u_ca_out_776;
wire [47:0] u_ca_out_777;
wire [47:0] u_ca_out_778;
wire [47:0] u_ca_out_779;
wire [47:0] u_ca_out_780;
wire [47:0] u_ca_out_781;
wire [47:0] u_ca_out_782;
wire [47:0] u_ca_out_783;
wire [47:0] u_ca_out_784;
wire [47:0] u_ca_out_785;
wire [47:0] u_ca_out_786;
wire [47:0] u_ca_out_787;
wire [47:0] u_ca_out_788;
wire [47:0] u_ca_out_789;
wire [47:0] u_ca_out_790;
wire [47:0] u_ca_out_791;
wire [47:0] u_ca_out_792;
wire [47:0] u_ca_out_793;
wire [47:0] u_ca_out_794;
wire [47:0] u_ca_out_795;
wire [47:0] u_ca_out_796;
wire [47:0] u_ca_out_797;
wire [47:0] u_ca_out_798;
wire [47:0] u_ca_out_799;
wire [47:0] u_ca_out_800;
wire [47:0] u_ca_out_801;
wire [47:0] u_ca_out_802;
wire [47:0] u_ca_out_803;
wire [47:0] u_ca_out_804;
wire [47:0] u_ca_out_805;
wire [47:0] u_ca_out_806;
wire [47:0] u_ca_out_807;
wire [47:0] u_ca_out_808;
wire [47:0] u_ca_out_809;
wire [47:0] u_ca_out_810;
wire [47:0] u_ca_out_811;
wire [47:0] u_ca_out_812;
wire [47:0] u_ca_out_813;
wire [47:0] u_ca_out_814;
wire [47:0] u_ca_out_815;
wire [47:0] u_ca_out_816;
wire [47:0] u_ca_out_817;
wire [47:0] u_ca_out_818;
wire [47:0] u_ca_out_819;
wire [47:0] u_ca_out_820;
wire [47:0] u_ca_out_821;
wire [47:0] u_ca_out_822;
wire [47:0] u_ca_out_823;
wire [47:0] u_ca_out_824;
wire [47:0] u_ca_out_825;
wire [47:0] u_ca_out_826;
wire [47:0] u_ca_out_827;
wire [47:0] u_ca_out_828;
wire [47:0] u_ca_out_829;
wire [47:0] u_ca_out_830;
wire [47:0] u_ca_out_831;
wire [47:0] u_ca_out_832;
wire [47:0] u_ca_out_833;
wire [47:0] u_ca_out_834;
wire [47:0] u_ca_out_835;
wire [47:0] u_ca_out_836;
wire [47:0] u_ca_out_837;
wire [47:0] u_ca_out_838;
wire [47:0] u_ca_out_839;
wire [47:0] u_ca_out_840;
wire [47:0] u_ca_out_841;
wire [47:0] u_ca_out_842;
wire [47:0] u_ca_out_843;
wire [47:0] u_ca_out_844;
wire [47:0] u_ca_out_845;
wire [47:0] u_ca_out_846;
wire [47:0] u_ca_out_847;
wire [47:0] u_ca_out_848;
wire [47:0] u_ca_out_849;
wire [47:0] u_ca_out_850;
wire [47:0] u_ca_out_851;
wire [47:0] u_ca_out_852;
wire [47:0] u_ca_out_853;
wire [47:0] u_ca_out_854;
wire [47:0] u_ca_out_855;
wire [47:0] u_ca_out_856;
wire [47:0] u_ca_out_857;
wire [47:0] u_ca_out_858;
wire [47:0] u_ca_out_859;
wire [47:0] u_ca_out_860;
wire [47:0] u_ca_out_861;
wire [47:0] u_ca_out_862;
wire [47:0] u_ca_out_863;
wire [47:0] u_ca_out_864;
wire [47:0] u_ca_out_865;
wire [47:0] u_ca_out_866;
wire [47:0] u_ca_out_867;
wire [47:0] u_ca_out_868;
wire [47:0] u_ca_out_869;
wire [47:0] u_ca_out_870;
wire [47:0] u_ca_out_871;
wire [47:0] u_ca_out_872;
wire [47:0] u_ca_out_873;
wire [47:0] u_ca_out_874;
wire [47:0] u_ca_out_875;
wire [47:0] u_ca_out_876;
wire [47:0] u_ca_out_877;
wire [47:0] u_ca_out_878;
wire [47:0] u_ca_out_879;
wire [47:0] u_ca_out_880;
wire [47:0] u_ca_out_881;
wire [47:0] u_ca_out_882;
wire [47:0] u_ca_out_883;
wire [47:0] u_ca_out_884;
wire [47:0] u_ca_out_885;
wire [47:0] u_ca_out_886;
wire [47:0] u_ca_out_887;
wire [47:0] u_ca_out_888;
wire [47:0] u_ca_out_889;
wire [47:0] u_ca_out_890;
wire [47:0] u_ca_out_891;
wire [47:0] u_ca_out_892;
wire [47:0] u_ca_out_893;
wire [47:0] u_ca_out_894;
wire [47:0] u_ca_out_895;
wire [47:0] u_ca_out_896;
wire [47:0] u_ca_out_897;
wire [47:0] u_ca_out_898;
wire [47:0] u_ca_out_899;
wire [47:0] u_ca_out_900;
wire [47:0] u_ca_out_901;
wire [47:0] u_ca_out_902;
wire [47:0] u_ca_out_903;
wire [47:0] u_ca_out_904;
wire [47:0] u_ca_out_905;
wire [47:0] u_ca_out_906;
wire [47:0] u_ca_out_907;
wire [47:0] u_ca_out_908;
wire [47:0] u_ca_out_909;
wire [47:0] u_ca_out_910;
wire [47:0] u_ca_out_911;
wire [47:0] u_ca_out_912;
wire [47:0] u_ca_out_913;
wire [47:0] u_ca_out_914;
wire [47:0] u_ca_out_915;
wire [47:0] u_ca_out_916;
wire [47:0] u_ca_out_917;
wire [47:0] u_ca_out_918;
wire [47:0] u_ca_out_919;
wire [47:0] u_ca_out_920;
wire [47:0] u_ca_out_921;
wire [47:0] u_ca_out_922;
wire [47:0] u_ca_out_923;
wire [47:0] u_ca_out_924;
wire [47:0] u_ca_out_925;
wire [47:0] u_ca_out_926;
wire [47:0] u_ca_out_927;
wire [47:0] u_ca_out_928;
wire [47:0] u_ca_out_929;
wire [47:0] u_ca_out_930;
wire [47:0] u_ca_out_931;
wire [47:0] u_ca_out_932;
wire [47:0] u_ca_out_933;
wire [47:0] u_ca_out_934;
wire [47:0] u_ca_out_935;
wire [47:0] u_ca_out_936;
wire [47:0] u_ca_out_937;
wire [47:0] u_ca_out_938;
wire [47:0] u_ca_out_939;
wire [47:0] u_ca_out_940;
wire [47:0] u_ca_out_941;
wire [47:0] u_ca_out_942;
wire [47:0] u_ca_out_943;
wire [47:0] u_ca_out_944;
wire [47:0] u_ca_out_945;
wire [47:0] u_ca_out_946;
wire [47:0] u_ca_out_947;
wire [47:0] u_ca_out_948;
wire [47:0] u_ca_out_949;
wire [47:0] u_ca_out_950;
wire [47:0] u_ca_out_951;
wire [47:0] u_ca_out_952;
wire [47:0] u_ca_out_953;
wire [47:0] u_ca_out_954;
wire [47:0] u_ca_out_955;
wire [47:0] u_ca_out_956;
wire [47:0] u_ca_out_957;
wire [47:0] u_ca_out_958;
wire [47:0] u_ca_out_959;
wire [47:0] u_ca_out_960;
wire [47:0] u_ca_out_961;
wire [47:0] u_ca_out_962;
wire [47:0] u_ca_out_963;
wire [47:0] u_ca_out_964;
wire [47:0] u_ca_out_965;
wire [47:0] u_ca_out_966;
wire [47:0] u_ca_out_967;
wire [47:0] u_ca_out_968;
wire [47:0] u_ca_out_969;
wire [47:0] u_ca_out_970;
wire [47:0] u_ca_out_971;
wire [47:0] u_ca_out_972;
wire [47:0] u_ca_out_973;
wire [47:0] u_ca_out_974;
wire [47:0] u_ca_out_975;
wire [47:0] u_ca_out_976;
wire [47:0] u_ca_out_977;
wire [47:0] u_ca_out_978;
wire [47:0] u_ca_out_979;
wire [47:0] u_ca_out_980;
wire [47:0] u_ca_out_981;
wire [47:0] u_ca_out_982;
wire [47:0] u_ca_out_983;
wire [47:0] u_ca_out_984;
wire [47:0] u_ca_out_985;
wire [47:0] u_ca_out_986;
wire [47:0] u_ca_out_987;
wire [47:0] u_ca_out_988;
wire [47:0] u_ca_out_989;
wire [47:0] u_ca_out_990;
wire [47:0] u_ca_out_991;
wire [47:0] u_ca_out_992;
wire [47:0] u_ca_out_993;
wire [47:0] u_ca_out_994;
wire [47:0] u_ca_out_995;
wire [47:0] u_ca_out_996;
wire [47:0] u_ca_out_997;
wire [47:0] u_ca_out_998;
wire [47:0] u_ca_out_999;
wire [47:0] u_ca_out_1000;
wire [47:0] u_ca_out_1001;
wire [47:0] u_ca_out_1002;
wire [47:0] u_ca_out_1003;
wire [47:0] u_ca_out_1004;
wire [47:0] u_ca_out_1005;
wire [47:0] u_ca_out_1006;
wire [47:0] u_ca_out_1007;
wire [47:0] u_ca_out_1008;
wire [47:0] u_ca_out_1009;
wire [47:0] u_ca_out_1010;
wire [47:0] u_ca_out_1011;
wire [47:0] u_ca_out_1012;
wire [47:0] u_ca_out_1013;
wire [47:0] u_ca_out_1014;
wire [47:0] u_ca_out_1015;
wire [47:0] u_ca_out_1016;
wire [47:0] u_ca_out_1017;
wire [47:0] u_ca_out_1018;
wire [47:0] u_ca_out_1019;
wire [47:0] u_ca_out_1020;
wire [47:0] u_ca_out_1021;
wire [47:0] u_ca_out_1022;
wire [47:0] u_ca_out_1023;
wire [47:0] u_ca_out_1024;
wire [47:0] u_ca_out_1025;
wire [47:0] u_ca_out_1026;

assign u_ca_in_0 = {{10{1'b0}}, col_in_0};
assign u_ca_in_1 = {{10{1'b0}}, col_in_1};
assign u_ca_in_2 = {{10{1'b0}}, col_in_2};
assign u_ca_in_3 = {{10{1'b0}}, col_in_3};
assign u_ca_in_4 = {{10{1'b0}}, col_in_4};
assign u_ca_in_5 = {{10{1'b0}}, col_in_5};
assign u_ca_in_6 = {{10{1'b0}}, col_in_6};
assign u_ca_in_7 = {{10{1'b0}}, col_in_7};
assign u_ca_in_8 = {{10{1'b0}}, col_in_8};
assign u_ca_in_9 = {{10{1'b0}}, col_in_9};
assign u_ca_in_10 = {{10{1'b0}}, col_in_10};
assign u_ca_in_11 = {{10{1'b0}}, col_in_11};
assign u_ca_in_12 = {{10{1'b0}}, col_in_12};
assign u_ca_in_13 = {{10{1'b0}}, col_in_13};
assign u_ca_in_14 = {{10{1'b0}}, col_in_14};
assign u_ca_in_15 = {{10{1'b0}}, col_in_15};
assign u_ca_in_16 = {{10{1'b0}}, col_in_16};
assign u_ca_in_17 = {{10{1'b0}}, col_in_17};
assign u_ca_in_18 = {{10{1'b0}}, col_in_18};
assign u_ca_in_19 = {{10{1'b0}}, col_in_19};
assign u_ca_in_20 = {{10{1'b0}}, col_in_20};
assign u_ca_in_21 = {{10{1'b0}}, col_in_21};
assign u_ca_in_22 = {{10{1'b0}}, col_in_22};
assign u_ca_in_23 = {{10{1'b0}}, col_in_23};
assign u_ca_in_24 = {{10{1'b0}}, col_in_24};
assign u_ca_in_25 = {{10{1'b0}}, col_in_25};
assign u_ca_in_26 = {{10{1'b0}}, col_in_26};
assign u_ca_in_27 = {{10{1'b0}}, col_in_27};
assign u_ca_in_28 = {{10{1'b0}}, col_in_28};
assign u_ca_in_29 = {{10{1'b0}}, col_in_29};
assign u_ca_in_30 = {{10{1'b0}}, col_in_30};
assign u_ca_in_31 = {{10{1'b0}}, col_in_31};
assign u_ca_in_32 = {{10{1'b0}}, col_in_32};
assign u_ca_in_33 = {{10{1'b0}}, col_in_33};
assign u_ca_in_34 = {{10{1'b0}}, col_in_34};
assign u_ca_in_35 = {{10{1'b0}}, col_in_35};
assign u_ca_in_36 = {{10{1'b0}}, col_in_36};
assign u_ca_in_37 = {{10{1'b0}}, col_in_37};
assign u_ca_in_38 = {{10{1'b0}}, col_in_38};
assign u_ca_in_39 = {{10{1'b0}}, col_in_39};
assign u_ca_in_40 = {{10{1'b0}}, col_in_40};
assign u_ca_in_41 = {{10{1'b0}}, col_in_41};
assign u_ca_in_42 = {{10{1'b0}}, col_in_42};
assign u_ca_in_43 = {{10{1'b0}}, col_in_43};
assign u_ca_in_44 = {{10{1'b0}}, col_in_44};
assign u_ca_in_45 = {{10{1'b0}}, col_in_45};
assign u_ca_in_46 = {{10{1'b0}}, col_in_46};
assign u_ca_in_47 = {{10{1'b0}}, col_in_47};
assign u_ca_in_48 = {{10{1'b0}}, col_in_48};
assign u_ca_in_49 = {{10{1'b0}}, col_in_49};
assign u_ca_in_50 = {{10{1'b0}}, col_in_50};
assign u_ca_in_51 = {{10{1'b0}}, col_in_51};
assign u_ca_in_52 = {{10{1'b0}}, col_in_52};
assign u_ca_in_53 = {{10{1'b0}}, col_in_53};
assign u_ca_in_54 = {{10{1'b0}}, col_in_54};
assign u_ca_in_55 = {{10{1'b0}}, col_in_55};
assign u_ca_in_56 = {{10{1'b0}}, col_in_56};
assign u_ca_in_57 = {{10{1'b0}}, col_in_57};
assign u_ca_in_58 = {{10{1'b0}}, col_in_58};
assign u_ca_in_59 = {{10{1'b0}}, col_in_59};
assign u_ca_in_60 = {{10{1'b0}}, col_in_60};
assign u_ca_in_61 = {{10{1'b0}}, col_in_61};
assign u_ca_in_62 = {{10{1'b0}}, col_in_62};
assign u_ca_in_63 = {{10{1'b0}}, col_in_63};
assign u_ca_in_64 = {{10{1'b0}}, col_in_64};
assign u_ca_in_65 = {{10{1'b0}}, col_in_65};
assign u_ca_in_66 = {{10{1'b0}}, col_in_66};
assign u_ca_in_67 = {{10{1'b0}}, col_in_67};
assign u_ca_in_68 = {{10{1'b0}}, col_in_68};
assign u_ca_in_69 = {{10{1'b0}}, col_in_69};
assign u_ca_in_70 = {{10{1'b0}}, col_in_70};
assign u_ca_in_71 = {{10{1'b0}}, col_in_71};
assign u_ca_in_72 = {{10{1'b0}}, col_in_72};
assign u_ca_in_73 = {{10{1'b0}}, col_in_73};
assign u_ca_in_74 = {{10{1'b0}}, col_in_74};
assign u_ca_in_75 = {{10{1'b0}}, col_in_75};
assign u_ca_in_76 = {{10{1'b0}}, col_in_76};
assign u_ca_in_77 = {{10{1'b0}}, col_in_77};
assign u_ca_in_78 = {{10{1'b0}}, col_in_78};
assign u_ca_in_79 = {{10{1'b0}}, col_in_79};
assign u_ca_in_80 = {{10{1'b0}}, col_in_80};
assign u_ca_in_81 = {{10{1'b0}}, col_in_81};
assign u_ca_in_82 = {{10{1'b0}}, col_in_82};
assign u_ca_in_83 = {{10{1'b0}}, col_in_83};
assign u_ca_in_84 = {{10{1'b0}}, col_in_84};
assign u_ca_in_85 = {{10{1'b0}}, col_in_85};
assign u_ca_in_86 = {{10{1'b0}}, col_in_86};
assign u_ca_in_87 = {{10{1'b0}}, col_in_87};
assign u_ca_in_88 = {{10{1'b0}}, col_in_88};
assign u_ca_in_89 = {{10{1'b0}}, col_in_89};
assign u_ca_in_90 = {{10{1'b0}}, col_in_90};
assign u_ca_in_91 = {{10{1'b0}}, col_in_91};
assign u_ca_in_92 = {{10{1'b0}}, col_in_92};
assign u_ca_in_93 = {{10{1'b0}}, col_in_93};
assign u_ca_in_94 = {{10{1'b0}}, col_in_94};
assign u_ca_in_95 = {{10{1'b0}}, col_in_95};
assign u_ca_in_96 = {{10{1'b0}}, col_in_96};
assign u_ca_in_97 = {{10{1'b0}}, col_in_97};
assign u_ca_in_98 = {{10{1'b0}}, col_in_98};
assign u_ca_in_99 = {{10{1'b0}}, col_in_99};
assign u_ca_in_100 = {{10{1'b0}}, col_in_100};
assign u_ca_in_101 = {{10{1'b0}}, col_in_101};
assign u_ca_in_102 = {{10{1'b0}}, col_in_102};
assign u_ca_in_103 = {{10{1'b0}}, col_in_103};
assign u_ca_in_104 = {{10{1'b0}}, col_in_104};
assign u_ca_in_105 = {{10{1'b0}}, col_in_105};
assign u_ca_in_106 = {{10{1'b0}}, col_in_106};
assign u_ca_in_107 = {{10{1'b0}}, col_in_107};
assign u_ca_in_108 = {{10{1'b0}}, col_in_108};
assign u_ca_in_109 = {{10{1'b0}}, col_in_109};
assign u_ca_in_110 = {{10{1'b0}}, col_in_110};
assign u_ca_in_111 = {{10{1'b0}}, col_in_111};
assign u_ca_in_112 = {{10{1'b0}}, col_in_112};
assign u_ca_in_113 = {{10{1'b0}}, col_in_113};
assign u_ca_in_114 = {{10{1'b0}}, col_in_114};
assign u_ca_in_115 = {{10{1'b0}}, col_in_115};
assign u_ca_in_116 = {{10{1'b0}}, col_in_116};
assign u_ca_in_117 = {{10{1'b0}}, col_in_117};
assign u_ca_in_118 = {{10{1'b0}}, col_in_118};
assign u_ca_in_119 = {{10{1'b0}}, col_in_119};
assign u_ca_in_120 = {{10{1'b0}}, col_in_120};
assign u_ca_in_121 = {{10{1'b0}}, col_in_121};
assign u_ca_in_122 = {{10{1'b0}}, col_in_122};
assign u_ca_in_123 = {{10{1'b0}}, col_in_123};
assign u_ca_in_124 = {{10{1'b0}}, col_in_124};
assign u_ca_in_125 = {{10{1'b0}}, col_in_125};
assign u_ca_in_126 = {{10{1'b0}}, col_in_126};
assign u_ca_in_127 = {{10{1'b0}}, col_in_127};
assign u_ca_in_128 = {{10{1'b0}}, col_in_128};
assign u_ca_in_129 = {{10{1'b0}}, col_in_129};
assign u_ca_in_130 = {{10{1'b0}}, col_in_130};
assign u_ca_in_131 = {{10{1'b0}}, col_in_131};
assign u_ca_in_132 = {{10{1'b0}}, col_in_132};
assign u_ca_in_133 = {{10{1'b0}}, col_in_133};
assign u_ca_in_134 = {{10{1'b0}}, col_in_134};
assign u_ca_in_135 = {{10{1'b0}}, col_in_135};
assign u_ca_in_136 = {{10{1'b0}}, col_in_136};
assign u_ca_in_137 = {{10{1'b0}}, col_in_137};
assign u_ca_in_138 = {{10{1'b0}}, col_in_138};
assign u_ca_in_139 = {{10{1'b0}}, col_in_139};
assign u_ca_in_140 = {{10{1'b0}}, col_in_140};
assign u_ca_in_141 = {{10{1'b0}}, col_in_141};
assign u_ca_in_142 = {{10{1'b0}}, col_in_142};
assign u_ca_in_143 = {{10{1'b0}}, col_in_143};
assign u_ca_in_144 = {{10{1'b0}}, col_in_144};
assign u_ca_in_145 = {{10{1'b0}}, col_in_145};
assign u_ca_in_146 = {{10{1'b0}}, col_in_146};
assign u_ca_in_147 = {{10{1'b0}}, col_in_147};
assign u_ca_in_148 = {{10{1'b0}}, col_in_148};
assign u_ca_in_149 = {{10{1'b0}}, col_in_149};
assign u_ca_in_150 = {{10{1'b0}}, col_in_150};
assign u_ca_in_151 = {{10{1'b0}}, col_in_151};
assign u_ca_in_152 = {{10{1'b0}}, col_in_152};
assign u_ca_in_153 = {{10{1'b0}}, col_in_153};
assign u_ca_in_154 = {{10{1'b0}}, col_in_154};
assign u_ca_in_155 = {{10{1'b0}}, col_in_155};
assign u_ca_in_156 = {{10{1'b0}}, col_in_156};
assign u_ca_in_157 = {{10{1'b0}}, col_in_157};
assign u_ca_in_158 = {{10{1'b0}}, col_in_158};
assign u_ca_in_159 = {{10{1'b0}}, col_in_159};
assign u_ca_in_160 = {{10{1'b0}}, col_in_160};
assign u_ca_in_161 = {{10{1'b0}}, col_in_161};
assign u_ca_in_162 = {{10{1'b0}}, col_in_162};
assign u_ca_in_163 = {{10{1'b0}}, col_in_163};
assign u_ca_in_164 = {{10{1'b0}}, col_in_164};
assign u_ca_in_165 = {{10{1'b0}}, col_in_165};
assign u_ca_in_166 = {{10{1'b0}}, col_in_166};
assign u_ca_in_167 = {{10{1'b0}}, col_in_167};
assign u_ca_in_168 = {{10{1'b0}}, col_in_168};
assign u_ca_in_169 = {{10{1'b0}}, col_in_169};
assign u_ca_in_170 = {{10{1'b0}}, col_in_170};
assign u_ca_in_171 = {{10{1'b0}}, col_in_171};
assign u_ca_in_172 = {{10{1'b0}}, col_in_172};
assign u_ca_in_173 = {{10{1'b0}}, col_in_173};
assign u_ca_in_174 = {{10{1'b0}}, col_in_174};
assign u_ca_in_175 = {{10{1'b0}}, col_in_175};
assign u_ca_in_176 = {{10{1'b0}}, col_in_176};
assign u_ca_in_177 = {{10{1'b0}}, col_in_177};
assign u_ca_in_178 = {{10{1'b0}}, col_in_178};
assign u_ca_in_179 = {{10{1'b0}}, col_in_179};
assign u_ca_in_180 = {{10{1'b0}}, col_in_180};
assign u_ca_in_181 = {{10{1'b0}}, col_in_181};
assign u_ca_in_182 = {{10{1'b0}}, col_in_182};
assign u_ca_in_183 = {{10{1'b0}}, col_in_183};
assign u_ca_in_184 = {{10{1'b0}}, col_in_184};
assign u_ca_in_185 = {{10{1'b0}}, col_in_185};
assign u_ca_in_186 = {{10{1'b0}}, col_in_186};
assign u_ca_in_187 = {{10{1'b0}}, col_in_187};
assign u_ca_in_188 = {{10{1'b0}}, col_in_188};
assign u_ca_in_189 = {{10{1'b0}}, col_in_189};
assign u_ca_in_190 = {{10{1'b0}}, col_in_190};
assign u_ca_in_191 = {{10{1'b0}}, col_in_191};
assign u_ca_in_192 = {{10{1'b0}}, col_in_192};
assign u_ca_in_193 = {{10{1'b0}}, col_in_193};
assign u_ca_in_194 = {{10{1'b0}}, col_in_194};
assign u_ca_in_195 = {{10{1'b0}}, col_in_195};
assign u_ca_in_196 = {{10{1'b0}}, col_in_196};
assign u_ca_in_197 = {{10{1'b0}}, col_in_197};
assign u_ca_in_198 = {{10{1'b0}}, col_in_198};
assign u_ca_in_199 = {{10{1'b0}}, col_in_199};
assign u_ca_in_200 = {{10{1'b0}}, col_in_200};
assign u_ca_in_201 = {{10{1'b0}}, col_in_201};
assign u_ca_in_202 = {{10{1'b0}}, col_in_202};
assign u_ca_in_203 = {{10{1'b0}}, col_in_203};
assign u_ca_in_204 = {{10{1'b0}}, col_in_204};
assign u_ca_in_205 = {{10{1'b0}}, col_in_205};
assign u_ca_in_206 = {{10{1'b0}}, col_in_206};
assign u_ca_in_207 = {{10{1'b0}}, col_in_207};
assign u_ca_in_208 = {{10{1'b0}}, col_in_208};
assign u_ca_in_209 = {{10{1'b0}}, col_in_209};
assign u_ca_in_210 = {{10{1'b0}}, col_in_210};
assign u_ca_in_211 = {{10{1'b0}}, col_in_211};
assign u_ca_in_212 = {{10{1'b0}}, col_in_212};
assign u_ca_in_213 = {{10{1'b0}}, col_in_213};
assign u_ca_in_214 = {{10{1'b0}}, col_in_214};
assign u_ca_in_215 = {{10{1'b0}}, col_in_215};
assign u_ca_in_216 = {{10{1'b0}}, col_in_216};
assign u_ca_in_217 = {{10{1'b0}}, col_in_217};
assign u_ca_in_218 = {{10{1'b0}}, col_in_218};
assign u_ca_in_219 = {{10{1'b0}}, col_in_219};
assign u_ca_in_220 = {{10{1'b0}}, col_in_220};
assign u_ca_in_221 = {{10{1'b0}}, col_in_221};
assign u_ca_in_222 = {{10{1'b0}}, col_in_222};
assign u_ca_in_223 = {{10{1'b0}}, col_in_223};
assign u_ca_in_224 = {{10{1'b0}}, col_in_224};
assign u_ca_in_225 = {{10{1'b0}}, col_in_225};
assign u_ca_in_226 = {{10{1'b0}}, col_in_226};
assign u_ca_in_227 = {{10{1'b0}}, col_in_227};
assign u_ca_in_228 = {{10{1'b0}}, col_in_228};
assign u_ca_in_229 = {{10{1'b0}}, col_in_229};
assign u_ca_in_230 = {{10{1'b0}}, col_in_230};
assign u_ca_in_231 = {{10{1'b0}}, col_in_231};
assign u_ca_in_232 = {{10{1'b0}}, col_in_232};
assign u_ca_in_233 = {{10{1'b0}}, col_in_233};
assign u_ca_in_234 = {{10{1'b0}}, col_in_234};
assign u_ca_in_235 = {{10{1'b0}}, col_in_235};
assign u_ca_in_236 = {{10{1'b0}}, col_in_236};
assign u_ca_in_237 = {{10{1'b0}}, col_in_237};
assign u_ca_in_238 = {{10{1'b0}}, col_in_238};
assign u_ca_in_239 = {{10{1'b0}}, col_in_239};
assign u_ca_in_240 = {{10{1'b0}}, col_in_240};
assign u_ca_in_241 = {{10{1'b0}}, col_in_241};
assign u_ca_in_242 = {{10{1'b0}}, col_in_242};
assign u_ca_in_243 = {{10{1'b0}}, col_in_243};
assign u_ca_in_244 = {{10{1'b0}}, col_in_244};
assign u_ca_in_245 = {{10{1'b0}}, col_in_245};
assign u_ca_in_246 = {{10{1'b0}}, col_in_246};
assign u_ca_in_247 = {{10{1'b0}}, col_in_247};
assign u_ca_in_248 = {{10{1'b0}}, col_in_248};
assign u_ca_in_249 = {{10{1'b0}}, col_in_249};
assign u_ca_in_250 = {{10{1'b0}}, col_in_250};
assign u_ca_in_251 = {{10{1'b0}}, col_in_251};
assign u_ca_in_252 = {{10{1'b0}}, col_in_252};
assign u_ca_in_253 = {{10{1'b0}}, col_in_253};
assign u_ca_in_254 = {{10{1'b0}}, col_in_254};
assign u_ca_in_255 = {{10{1'b0}}, col_in_255};
assign u_ca_in_256 = {{10{1'b0}}, col_in_256};
assign u_ca_in_257 = {{10{1'b0}}, col_in_257};
assign u_ca_in_258 = {{10{1'b0}}, col_in_258};
assign u_ca_in_259 = {{10{1'b0}}, col_in_259};
assign u_ca_in_260 = {{10{1'b0}}, col_in_260};
assign u_ca_in_261 = {{10{1'b0}}, col_in_261};
assign u_ca_in_262 = {{10{1'b0}}, col_in_262};
assign u_ca_in_263 = {{10{1'b0}}, col_in_263};
assign u_ca_in_264 = {{10{1'b0}}, col_in_264};
assign u_ca_in_265 = {{10{1'b0}}, col_in_265};
assign u_ca_in_266 = {{10{1'b0}}, col_in_266};
assign u_ca_in_267 = {{10{1'b0}}, col_in_267};
assign u_ca_in_268 = {{10{1'b0}}, col_in_268};
assign u_ca_in_269 = {{10{1'b0}}, col_in_269};
assign u_ca_in_270 = {{10{1'b0}}, col_in_270};
assign u_ca_in_271 = {{10{1'b0}}, col_in_271};
assign u_ca_in_272 = {{10{1'b0}}, col_in_272};
assign u_ca_in_273 = {{10{1'b0}}, col_in_273};
assign u_ca_in_274 = {{10{1'b0}}, col_in_274};
assign u_ca_in_275 = {{10{1'b0}}, col_in_275};
assign u_ca_in_276 = {{10{1'b0}}, col_in_276};
assign u_ca_in_277 = {{10{1'b0}}, col_in_277};
assign u_ca_in_278 = {{10{1'b0}}, col_in_278};
assign u_ca_in_279 = {{10{1'b0}}, col_in_279};
assign u_ca_in_280 = {{10{1'b0}}, col_in_280};
assign u_ca_in_281 = {{10{1'b0}}, col_in_281};
assign u_ca_in_282 = {{10{1'b0}}, col_in_282};
assign u_ca_in_283 = {{10{1'b0}}, col_in_283};
assign u_ca_in_284 = {{10{1'b0}}, col_in_284};
assign u_ca_in_285 = {{10{1'b0}}, col_in_285};
assign u_ca_in_286 = {{10{1'b0}}, col_in_286};
assign u_ca_in_287 = {{10{1'b0}}, col_in_287};
assign u_ca_in_288 = {{10{1'b0}}, col_in_288};
assign u_ca_in_289 = {{10{1'b0}}, col_in_289};
assign u_ca_in_290 = {{10{1'b0}}, col_in_290};
assign u_ca_in_291 = {{10{1'b0}}, col_in_291};
assign u_ca_in_292 = {{10{1'b0}}, col_in_292};
assign u_ca_in_293 = {{10{1'b0}}, col_in_293};
assign u_ca_in_294 = {{10{1'b0}}, col_in_294};
assign u_ca_in_295 = {{10{1'b0}}, col_in_295};
assign u_ca_in_296 = {{10{1'b0}}, col_in_296};
assign u_ca_in_297 = {{10{1'b0}}, col_in_297};
assign u_ca_in_298 = {{10{1'b0}}, col_in_298};
assign u_ca_in_299 = {{10{1'b0}}, col_in_299};
assign u_ca_in_300 = {{10{1'b0}}, col_in_300};
assign u_ca_in_301 = {{10{1'b0}}, col_in_301};
assign u_ca_in_302 = {{10{1'b0}}, col_in_302};
assign u_ca_in_303 = {{10{1'b0}}, col_in_303};
assign u_ca_in_304 = {{10{1'b0}}, col_in_304};
assign u_ca_in_305 = {{10{1'b0}}, col_in_305};
assign u_ca_in_306 = {{10{1'b0}}, col_in_306};
assign u_ca_in_307 = {{10{1'b0}}, col_in_307};
assign u_ca_in_308 = {{10{1'b0}}, col_in_308};
assign u_ca_in_309 = {{10{1'b0}}, col_in_309};
assign u_ca_in_310 = {{10{1'b0}}, col_in_310};
assign u_ca_in_311 = {{10{1'b0}}, col_in_311};
assign u_ca_in_312 = {{10{1'b0}}, col_in_312};
assign u_ca_in_313 = {{10{1'b0}}, col_in_313};
assign u_ca_in_314 = {{10{1'b0}}, col_in_314};
assign u_ca_in_315 = {{10{1'b0}}, col_in_315};
assign u_ca_in_316 = {{10{1'b0}}, col_in_316};
assign u_ca_in_317 = {{10{1'b0}}, col_in_317};
assign u_ca_in_318 = {{10{1'b0}}, col_in_318};
assign u_ca_in_319 = {{10{1'b0}}, col_in_319};
assign u_ca_in_320 = {{10{1'b0}}, col_in_320};
assign u_ca_in_321 = {{10{1'b0}}, col_in_321};
assign u_ca_in_322 = {{10{1'b0}}, col_in_322};
assign u_ca_in_323 = {{10{1'b0}}, col_in_323};
assign u_ca_in_324 = {{10{1'b0}}, col_in_324};
assign u_ca_in_325 = {{10{1'b0}}, col_in_325};
assign u_ca_in_326 = {{10{1'b0}}, col_in_326};
assign u_ca_in_327 = {{10{1'b0}}, col_in_327};
assign u_ca_in_328 = {{10{1'b0}}, col_in_328};
assign u_ca_in_329 = {{10{1'b0}}, col_in_329};
assign u_ca_in_330 = {{10{1'b0}}, col_in_330};
assign u_ca_in_331 = {{10{1'b0}}, col_in_331};
assign u_ca_in_332 = {{10{1'b0}}, col_in_332};
assign u_ca_in_333 = {{10{1'b0}}, col_in_333};
assign u_ca_in_334 = {{10{1'b0}}, col_in_334};
assign u_ca_in_335 = {{10{1'b0}}, col_in_335};
assign u_ca_in_336 = {{10{1'b0}}, col_in_336};
assign u_ca_in_337 = {{10{1'b0}}, col_in_337};
assign u_ca_in_338 = {{10{1'b0}}, col_in_338};
assign u_ca_in_339 = {{10{1'b0}}, col_in_339};
assign u_ca_in_340 = {{10{1'b0}}, col_in_340};
assign u_ca_in_341 = {{10{1'b0}}, col_in_341};
assign u_ca_in_342 = {{10{1'b0}}, col_in_342};
assign u_ca_in_343 = {{10{1'b0}}, col_in_343};
assign u_ca_in_344 = {{10{1'b0}}, col_in_344};
assign u_ca_in_345 = {{10{1'b0}}, col_in_345};
assign u_ca_in_346 = {{10{1'b0}}, col_in_346};
assign u_ca_in_347 = {{10{1'b0}}, col_in_347};
assign u_ca_in_348 = {{10{1'b0}}, col_in_348};
assign u_ca_in_349 = {{10{1'b0}}, col_in_349};
assign u_ca_in_350 = {{10{1'b0}}, col_in_350};
assign u_ca_in_351 = {{10{1'b0}}, col_in_351};
assign u_ca_in_352 = {{10{1'b0}}, col_in_352};
assign u_ca_in_353 = {{10{1'b0}}, col_in_353};
assign u_ca_in_354 = {{10{1'b0}}, col_in_354};
assign u_ca_in_355 = {{10{1'b0}}, col_in_355};
assign u_ca_in_356 = {{10{1'b0}}, col_in_356};
assign u_ca_in_357 = {{10{1'b0}}, col_in_357};
assign u_ca_in_358 = {{10{1'b0}}, col_in_358};
assign u_ca_in_359 = {{10{1'b0}}, col_in_359};
assign u_ca_in_360 = {{10{1'b0}}, col_in_360};
assign u_ca_in_361 = {{10{1'b0}}, col_in_361};
assign u_ca_in_362 = {{10{1'b0}}, col_in_362};
assign u_ca_in_363 = {{10{1'b0}}, col_in_363};
assign u_ca_in_364 = {{10{1'b0}}, col_in_364};
assign u_ca_in_365 = {{10{1'b0}}, col_in_365};
assign u_ca_in_366 = {{10{1'b0}}, col_in_366};
assign u_ca_in_367 = {{10{1'b0}}, col_in_367};
assign u_ca_in_368 = {{10{1'b0}}, col_in_368};
assign u_ca_in_369 = {{10{1'b0}}, col_in_369};
assign u_ca_in_370 = {{10{1'b0}}, col_in_370};
assign u_ca_in_371 = {{10{1'b0}}, col_in_371};
assign u_ca_in_372 = {{10{1'b0}}, col_in_372};
assign u_ca_in_373 = {{10{1'b0}}, col_in_373};
assign u_ca_in_374 = {{10{1'b0}}, col_in_374};
assign u_ca_in_375 = {{10{1'b0}}, col_in_375};
assign u_ca_in_376 = {{10{1'b0}}, col_in_376};
assign u_ca_in_377 = {{10{1'b0}}, col_in_377};
assign u_ca_in_378 = {{10{1'b0}}, col_in_378};
assign u_ca_in_379 = {{10{1'b0}}, col_in_379};
assign u_ca_in_380 = {{10{1'b0}}, col_in_380};
assign u_ca_in_381 = {{10{1'b0}}, col_in_381};
assign u_ca_in_382 = {{10{1'b0}}, col_in_382};
assign u_ca_in_383 = {{10{1'b0}}, col_in_383};
assign u_ca_in_384 = {{10{1'b0}}, col_in_384};
assign u_ca_in_385 = {{10{1'b0}}, col_in_385};
assign u_ca_in_386 = {{10{1'b0}}, col_in_386};
assign u_ca_in_387 = {{10{1'b0}}, col_in_387};
assign u_ca_in_388 = {{10{1'b0}}, col_in_388};
assign u_ca_in_389 = {{10{1'b0}}, col_in_389};
assign u_ca_in_390 = {{10{1'b0}}, col_in_390};
assign u_ca_in_391 = {{10{1'b0}}, col_in_391};
assign u_ca_in_392 = {{10{1'b0}}, col_in_392};
assign u_ca_in_393 = {{10{1'b0}}, col_in_393};
assign u_ca_in_394 = {{10{1'b0}}, col_in_394};
assign u_ca_in_395 = {{10{1'b0}}, col_in_395};
assign u_ca_in_396 = {{10{1'b0}}, col_in_396};
assign u_ca_in_397 = {{10{1'b0}}, col_in_397};
assign u_ca_in_398 = {{10{1'b0}}, col_in_398};
assign u_ca_in_399 = {{10{1'b0}}, col_in_399};
assign u_ca_in_400 = {{10{1'b0}}, col_in_400};
assign u_ca_in_401 = {{10{1'b0}}, col_in_401};
assign u_ca_in_402 = {{10{1'b0}}, col_in_402};
assign u_ca_in_403 = {{10{1'b0}}, col_in_403};
assign u_ca_in_404 = {{10{1'b0}}, col_in_404};
assign u_ca_in_405 = {{10{1'b0}}, col_in_405};
assign u_ca_in_406 = {{10{1'b0}}, col_in_406};
assign u_ca_in_407 = {{10{1'b0}}, col_in_407};
assign u_ca_in_408 = {{10{1'b0}}, col_in_408};
assign u_ca_in_409 = {{10{1'b0}}, col_in_409};
assign u_ca_in_410 = {{10{1'b0}}, col_in_410};
assign u_ca_in_411 = {{10{1'b0}}, col_in_411};
assign u_ca_in_412 = {{10{1'b0}}, col_in_412};
assign u_ca_in_413 = {{10{1'b0}}, col_in_413};
assign u_ca_in_414 = {{10{1'b0}}, col_in_414};
assign u_ca_in_415 = {{10{1'b0}}, col_in_415};
assign u_ca_in_416 = {{10{1'b0}}, col_in_416};
assign u_ca_in_417 = {{10{1'b0}}, col_in_417};
assign u_ca_in_418 = {{10{1'b0}}, col_in_418};
assign u_ca_in_419 = {{10{1'b0}}, col_in_419};
assign u_ca_in_420 = {{10{1'b0}}, col_in_420};
assign u_ca_in_421 = {{10{1'b0}}, col_in_421};
assign u_ca_in_422 = {{10{1'b0}}, col_in_422};
assign u_ca_in_423 = {{10{1'b0}}, col_in_423};
assign u_ca_in_424 = {{10{1'b0}}, col_in_424};
assign u_ca_in_425 = {{10{1'b0}}, col_in_425};
assign u_ca_in_426 = {{10{1'b0}}, col_in_426};
assign u_ca_in_427 = {{10{1'b0}}, col_in_427};
assign u_ca_in_428 = {{10{1'b0}}, col_in_428};
assign u_ca_in_429 = {{10{1'b0}}, col_in_429};
assign u_ca_in_430 = {{10{1'b0}}, col_in_430};
assign u_ca_in_431 = {{10{1'b0}}, col_in_431};
assign u_ca_in_432 = {{10{1'b0}}, col_in_432};
assign u_ca_in_433 = {{10{1'b0}}, col_in_433};
assign u_ca_in_434 = {{10{1'b0}}, col_in_434};
assign u_ca_in_435 = {{10{1'b0}}, col_in_435};
assign u_ca_in_436 = {{10{1'b0}}, col_in_436};
assign u_ca_in_437 = {{10{1'b0}}, col_in_437};
assign u_ca_in_438 = {{10{1'b0}}, col_in_438};
assign u_ca_in_439 = {{10{1'b0}}, col_in_439};
assign u_ca_in_440 = {{10{1'b0}}, col_in_440};
assign u_ca_in_441 = {{10{1'b0}}, col_in_441};
assign u_ca_in_442 = {{10{1'b0}}, col_in_442};
assign u_ca_in_443 = {{10{1'b0}}, col_in_443};
assign u_ca_in_444 = {{10{1'b0}}, col_in_444};
assign u_ca_in_445 = {{10{1'b0}}, col_in_445};
assign u_ca_in_446 = {{10{1'b0}}, col_in_446};
assign u_ca_in_447 = {{10{1'b0}}, col_in_447};
assign u_ca_in_448 = {{10{1'b0}}, col_in_448};
assign u_ca_in_449 = {{10{1'b0}}, col_in_449};
assign u_ca_in_450 = {{10{1'b0}}, col_in_450};
assign u_ca_in_451 = {{10{1'b0}}, col_in_451};
assign u_ca_in_452 = {{10{1'b0}}, col_in_452};
assign u_ca_in_453 = {{10{1'b0}}, col_in_453};
assign u_ca_in_454 = {{10{1'b0}}, col_in_454};
assign u_ca_in_455 = {{10{1'b0}}, col_in_455};
assign u_ca_in_456 = {{10{1'b0}}, col_in_456};
assign u_ca_in_457 = {{10{1'b0}}, col_in_457};
assign u_ca_in_458 = {{10{1'b0}}, col_in_458};
assign u_ca_in_459 = {{10{1'b0}}, col_in_459};
assign u_ca_in_460 = {{10{1'b0}}, col_in_460};
assign u_ca_in_461 = {{10{1'b0}}, col_in_461};
assign u_ca_in_462 = {{10{1'b0}}, col_in_462};
assign u_ca_in_463 = {{10{1'b0}}, col_in_463};
assign u_ca_in_464 = {{10{1'b0}}, col_in_464};
assign u_ca_in_465 = {{10{1'b0}}, col_in_465};
assign u_ca_in_466 = {{10{1'b0}}, col_in_466};
assign u_ca_in_467 = {{10{1'b0}}, col_in_467};
assign u_ca_in_468 = {{10{1'b0}}, col_in_468};
assign u_ca_in_469 = {{10{1'b0}}, col_in_469};
assign u_ca_in_470 = {{10{1'b0}}, col_in_470};
assign u_ca_in_471 = {{10{1'b0}}, col_in_471};
assign u_ca_in_472 = {{10{1'b0}}, col_in_472};
assign u_ca_in_473 = {{10{1'b0}}, col_in_473};
assign u_ca_in_474 = {{10{1'b0}}, col_in_474};
assign u_ca_in_475 = {{10{1'b0}}, col_in_475};
assign u_ca_in_476 = {{10{1'b0}}, col_in_476};
assign u_ca_in_477 = {{10{1'b0}}, col_in_477};
assign u_ca_in_478 = {{10{1'b0}}, col_in_478};
assign u_ca_in_479 = {{10{1'b0}}, col_in_479};
assign u_ca_in_480 = {{10{1'b0}}, col_in_480};
assign u_ca_in_481 = {{10{1'b0}}, col_in_481};
assign u_ca_in_482 = {{10{1'b0}}, col_in_482};
assign u_ca_in_483 = {{10{1'b0}}, col_in_483};
assign u_ca_in_484 = {{10{1'b0}}, col_in_484};
assign u_ca_in_485 = {{10{1'b0}}, col_in_485};
assign u_ca_in_486 = {{10{1'b0}}, col_in_486};
assign u_ca_in_487 = {{10{1'b0}}, col_in_487};
assign u_ca_in_488 = {{10{1'b0}}, col_in_488};
assign u_ca_in_489 = {{10{1'b0}}, col_in_489};
assign u_ca_in_490 = {{10{1'b0}}, col_in_490};
assign u_ca_in_491 = {{10{1'b0}}, col_in_491};
assign u_ca_in_492 = {{10{1'b0}}, col_in_492};
assign u_ca_in_493 = {{10{1'b0}}, col_in_493};
assign u_ca_in_494 = {{10{1'b0}}, col_in_494};
assign u_ca_in_495 = {{10{1'b0}}, col_in_495};
assign u_ca_in_496 = {{10{1'b0}}, col_in_496};
assign u_ca_in_497 = {{10{1'b0}}, col_in_497};
assign u_ca_in_498 = {{10{1'b0}}, col_in_498};
assign u_ca_in_499 = {{10{1'b0}}, col_in_499};
assign u_ca_in_500 = {{10{1'b0}}, col_in_500};
assign u_ca_in_501 = {{10{1'b0}}, col_in_501};
assign u_ca_in_502 = {{10{1'b0}}, col_in_502};
assign u_ca_in_503 = {{10{1'b0}}, col_in_503};
assign u_ca_in_504 = {{10{1'b0}}, col_in_504};
assign u_ca_in_505 = {{10{1'b0}}, col_in_505};
assign u_ca_in_506 = {{10{1'b0}}, col_in_506};
assign u_ca_in_507 = {{10{1'b0}}, col_in_507};
assign u_ca_in_508 = {{10{1'b0}}, col_in_508};
assign u_ca_in_509 = {{10{1'b0}}, col_in_509};
assign u_ca_in_510 = {{10{1'b0}}, col_in_510};
assign u_ca_in_511 = {{10{1'b0}}, col_in_511};
assign u_ca_in_512 = {{10{1'b0}}, col_in_512};
assign u_ca_in_513 = {{10{1'b0}}, col_in_513};
assign u_ca_in_514 = {{10{1'b0}}, col_in_514};
assign u_ca_in_515 = {{10{1'b0}}, col_in_515};
assign u_ca_in_516 = {{10{1'b0}}, col_in_516};
assign u_ca_in_517 = {{10{1'b0}}, col_in_517};
assign u_ca_in_518 = {{10{1'b0}}, col_in_518};
assign u_ca_in_519 = {{10{1'b0}}, col_in_519};
assign u_ca_in_520 = {{10{1'b0}}, col_in_520};
assign u_ca_in_521 = {{10{1'b0}}, col_in_521};
assign u_ca_in_522 = {{10{1'b0}}, col_in_522};
assign u_ca_in_523 = {{10{1'b0}}, col_in_523};
assign u_ca_in_524 = {{10{1'b0}}, col_in_524};
assign u_ca_in_525 = {{10{1'b0}}, col_in_525};
assign u_ca_in_526 = {{10{1'b0}}, col_in_526};
assign u_ca_in_527 = {{10{1'b0}}, col_in_527};
assign u_ca_in_528 = {{10{1'b0}}, col_in_528};
assign u_ca_in_529 = {{10{1'b0}}, col_in_529};
assign u_ca_in_530 = {{10{1'b0}}, col_in_530};
assign u_ca_in_531 = {{10{1'b0}}, col_in_531};
assign u_ca_in_532 = {{10{1'b0}}, col_in_532};
assign u_ca_in_533 = {{10{1'b0}}, col_in_533};
assign u_ca_in_534 = {{10{1'b0}}, col_in_534};
assign u_ca_in_535 = {{10{1'b0}}, col_in_535};
assign u_ca_in_536 = {{10{1'b0}}, col_in_536};
assign u_ca_in_537 = {{10{1'b0}}, col_in_537};
assign u_ca_in_538 = {{10{1'b0}}, col_in_538};
assign u_ca_in_539 = {{10{1'b0}}, col_in_539};
assign u_ca_in_540 = {{10{1'b0}}, col_in_540};
assign u_ca_in_541 = {{10{1'b0}}, col_in_541};
assign u_ca_in_542 = {{10{1'b0}}, col_in_542};
assign u_ca_in_543 = {{10{1'b0}}, col_in_543};
assign u_ca_in_544 = {{10{1'b0}}, col_in_544};
assign u_ca_in_545 = {{10{1'b0}}, col_in_545};
assign u_ca_in_546 = {{10{1'b0}}, col_in_546};
assign u_ca_in_547 = {{10{1'b0}}, col_in_547};
assign u_ca_in_548 = {{10{1'b0}}, col_in_548};
assign u_ca_in_549 = {{10{1'b0}}, col_in_549};
assign u_ca_in_550 = {{10{1'b0}}, col_in_550};
assign u_ca_in_551 = {{10{1'b0}}, col_in_551};
assign u_ca_in_552 = {{10{1'b0}}, col_in_552};
assign u_ca_in_553 = {{10{1'b0}}, col_in_553};
assign u_ca_in_554 = {{10{1'b0}}, col_in_554};
assign u_ca_in_555 = {{10{1'b0}}, col_in_555};
assign u_ca_in_556 = {{10{1'b0}}, col_in_556};
assign u_ca_in_557 = {{10{1'b0}}, col_in_557};
assign u_ca_in_558 = {{10{1'b0}}, col_in_558};
assign u_ca_in_559 = {{10{1'b0}}, col_in_559};
assign u_ca_in_560 = {{10{1'b0}}, col_in_560};
assign u_ca_in_561 = {{10{1'b0}}, col_in_561};
assign u_ca_in_562 = {{10{1'b0}}, col_in_562};
assign u_ca_in_563 = {{10{1'b0}}, col_in_563};
assign u_ca_in_564 = {{10{1'b0}}, col_in_564};
assign u_ca_in_565 = {{10{1'b0}}, col_in_565};
assign u_ca_in_566 = {{10{1'b0}}, col_in_566};
assign u_ca_in_567 = {{10{1'b0}}, col_in_567};
assign u_ca_in_568 = {{10{1'b0}}, col_in_568};
assign u_ca_in_569 = {{10{1'b0}}, col_in_569};
assign u_ca_in_570 = {{10{1'b0}}, col_in_570};
assign u_ca_in_571 = {{10{1'b0}}, col_in_571};
assign u_ca_in_572 = {{10{1'b0}}, col_in_572};
assign u_ca_in_573 = {{10{1'b0}}, col_in_573};
assign u_ca_in_574 = {{10{1'b0}}, col_in_574};
assign u_ca_in_575 = {{10{1'b0}}, col_in_575};
assign u_ca_in_576 = {{10{1'b0}}, col_in_576};
assign u_ca_in_577 = {{10{1'b0}}, col_in_577};
assign u_ca_in_578 = {{10{1'b0}}, col_in_578};
assign u_ca_in_579 = {{10{1'b0}}, col_in_579};
assign u_ca_in_580 = {{10{1'b0}}, col_in_580};
assign u_ca_in_581 = {{10{1'b0}}, col_in_581};
assign u_ca_in_582 = {{10{1'b0}}, col_in_582};
assign u_ca_in_583 = {{10{1'b0}}, col_in_583};
assign u_ca_in_584 = {{10{1'b0}}, col_in_584};
assign u_ca_in_585 = {{10{1'b0}}, col_in_585};
assign u_ca_in_586 = {{10{1'b0}}, col_in_586};
assign u_ca_in_587 = {{10{1'b0}}, col_in_587};
assign u_ca_in_588 = {{10{1'b0}}, col_in_588};
assign u_ca_in_589 = {{10{1'b0}}, col_in_589};
assign u_ca_in_590 = {{10{1'b0}}, col_in_590};
assign u_ca_in_591 = {{10{1'b0}}, col_in_591};
assign u_ca_in_592 = {{10{1'b0}}, col_in_592};
assign u_ca_in_593 = {{10{1'b0}}, col_in_593};
assign u_ca_in_594 = {{10{1'b0}}, col_in_594};
assign u_ca_in_595 = {{10{1'b0}}, col_in_595};
assign u_ca_in_596 = {{10{1'b0}}, col_in_596};
assign u_ca_in_597 = {{10{1'b0}}, col_in_597};
assign u_ca_in_598 = {{10{1'b0}}, col_in_598};
assign u_ca_in_599 = {{10{1'b0}}, col_in_599};
assign u_ca_in_600 = {{10{1'b0}}, col_in_600};
assign u_ca_in_601 = {{10{1'b0}}, col_in_601};
assign u_ca_in_602 = {{10{1'b0}}, col_in_602};
assign u_ca_in_603 = {{10{1'b0}}, col_in_603};
assign u_ca_in_604 = {{10{1'b0}}, col_in_604};
assign u_ca_in_605 = {{10{1'b0}}, col_in_605};
assign u_ca_in_606 = {{10{1'b0}}, col_in_606};
assign u_ca_in_607 = {{10{1'b0}}, col_in_607};
assign u_ca_in_608 = {{10{1'b0}}, col_in_608};
assign u_ca_in_609 = {{10{1'b0}}, col_in_609};
assign u_ca_in_610 = {{10{1'b0}}, col_in_610};
assign u_ca_in_611 = {{10{1'b0}}, col_in_611};
assign u_ca_in_612 = {{10{1'b0}}, col_in_612};
assign u_ca_in_613 = {{10{1'b0}}, col_in_613};
assign u_ca_in_614 = {{10{1'b0}}, col_in_614};
assign u_ca_in_615 = {{10{1'b0}}, col_in_615};
assign u_ca_in_616 = {{10{1'b0}}, col_in_616};
assign u_ca_in_617 = {{10{1'b0}}, col_in_617};
assign u_ca_in_618 = {{10{1'b0}}, col_in_618};
assign u_ca_in_619 = {{10{1'b0}}, col_in_619};
assign u_ca_in_620 = {{10{1'b0}}, col_in_620};
assign u_ca_in_621 = {{10{1'b0}}, col_in_621};
assign u_ca_in_622 = {{10{1'b0}}, col_in_622};
assign u_ca_in_623 = {{10{1'b0}}, col_in_623};
assign u_ca_in_624 = {{10{1'b0}}, col_in_624};
assign u_ca_in_625 = {{10{1'b0}}, col_in_625};
assign u_ca_in_626 = {{10{1'b0}}, col_in_626};
assign u_ca_in_627 = {{10{1'b0}}, col_in_627};
assign u_ca_in_628 = {{10{1'b0}}, col_in_628};
assign u_ca_in_629 = {{10{1'b0}}, col_in_629};
assign u_ca_in_630 = {{10{1'b0}}, col_in_630};
assign u_ca_in_631 = {{10{1'b0}}, col_in_631};
assign u_ca_in_632 = {{10{1'b0}}, col_in_632};
assign u_ca_in_633 = {{10{1'b0}}, col_in_633};
assign u_ca_in_634 = {{10{1'b0}}, col_in_634};
assign u_ca_in_635 = {{10{1'b0}}, col_in_635};
assign u_ca_in_636 = {{10{1'b0}}, col_in_636};
assign u_ca_in_637 = {{10{1'b0}}, col_in_637};
assign u_ca_in_638 = {{10{1'b0}}, col_in_638};
assign u_ca_in_639 = {{10{1'b0}}, col_in_639};
assign u_ca_in_640 = {{10{1'b0}}, col_in_640};
assign u_ca_in_641 = {{10{1'b0}}, col_in_641};
assign u_ca_in_642 = {{10{1'b0}}, col_in_642};
assign u_ca_in_643 = {{10{1'b0}}, col_in_643};
assign u_ca_in_644 = {{10{1'b0}}, col_in_644};
assign u_ca_in_645 = {{10{1'b0}}, col_in_645};
assign u_ca_in_646 = {{10{1'b0}}, col_in_646};
assign u_ca_in_647 = {{10{1'b0}}, col_in_647};
assign u_ca_in_648 = {{10{1'b0}}, col_in_648};
assign u_ca_in_649 = {{10{1'b0}}, col_in_649};
assign u_ca_in_650 = {{10{1'b0}}, col_in_650};
assign u_ca_in_651 = {{10{1'b0}}, col_in_651};
assign u_ca_in_652 = {{10{1'b0}}, col_in_652};
assign u_ca_in_653 = {{10{1'b0}}, col_in_653};
assign u_ca_in_654 = {{10{1'b0}}, col_in_654};
assign u_ca_in_655 = {{10{1'b0}}, col_in_655};
assign u_ca_in_656 = {{10{1'b0}}, col_in_656};
assign u_ca_in_657 = {{10{1'b0}}, col_in_657};
assign u_ca_in_658 = {{10{1'b0}}, col_in_658};
assign u_ca_in_659 = {{10{1'b0}}, col_in_659};
assign u_ca_in_660 = {{10{1'b0}}, col_in_660};
assign u_ca_in_661 = {{10{1'b0}}, col_in_661};
assign u_ca_in_662 = {{10{1'b0}}, col_in_662};
assign u_ca_in_663 = {{10{1'b0}}, col_in_663};
assign u_ca_in_664 = {{10{1'b0}}, col_in_664};
assign u_ca_in_665 = {{10{1'b0}}, col_in_665};
assign u_ca_in_666 = {{10{1'b0}}, col_in_666};
assign u_ca_in_667 = {{10{1'b0}}, col_in_667};
assign u_ca_in_668 = {{10{1'b0}}, col_in_668};
assign u_ca_in_669 = {{10{1'b0}}, col_in_669};
assign u_ca_in_670 = {{10{1'b0}}, col_in_670};
assign u_ca_in_671 = {{10{1'b0}}, col_in_671};
assign u_ca_in_672 = {{10{1'b0}}, col_in_672};
assign u_ca_in_673 = {{10{1'b0}}, col_in_673};
assign u_ca_in_674 = {{10{1'b0}}, col_in_674};
assign u_ca_in_675 = {{10{1'b0}}, col_in_675};
assign u_ca_in_676 = {{10{1'b0}}, col_in_676};
assign u_ca_in_677 = {{10{1'b0}}, col_in_677};
assign u_ca_in_678 = {{10{1'b0}}, col_in_678};
assign u_ca_in_679 = {{10{1'b0}}, col_in_679};
assign u_ca_in_680 = {{10{1'b0}}, col_in_680};
assign u_ca_in_681 = {{10{1'b0}}, col_in_681};
assign u_ca_in_682 = {{10{1'b0}}, col_in_682};
assign u_ca_in_683 = {{10{1'b0}}, col_in_683};
assign u_ca_in_684 = {{10{1'b0}}, col_in_684};
assign u_ca_in_685 = {{10{1'b0}}, col_in_685};
assign u_ca_in_686 = {{10{1'b0}}, col_in_686};
assign u_ca_in_687 = {{10{1'b0}}, col_in_687};
assign u_ca_in_688 = {{10{1'b0}}, col_in_688};
assign u_ca_in_689 = {{10{1'b0}}, col_in_689};
assign u_ca_in_690 = {{10{1'b0}}, col_in_690};
assign u_ca_in_691 = {{10{1'b0}}, col_in_691};
assign u_ca_in_692 = {{10{1'b0}}, col_in_692};
assign u_ca_in_693 = {{10{1'b0}}, col_in_693};
assign u_ca_in_694 = {{10{1'b0}}, col_in_694};
assign u_ca_in_695 = {{10{1'b0}}, col_in_695};
assign u_ca_in_696 = {{10{1'b0}}, col_in_696};
assign u_ca_in_697 = {{10{1'b0}}, col_in_697};
assign u_ca_in_698 = {{10{1'b0}}, col_in_698};
assign u_ca_in_699 = {{10{1'b0}}, col_in_699};
assign u_ca_in_700 = {{10{1'b0}}, col_in_700};
assign u_ca_in_701 = {{10{1'b0}}, col_in_701};
assign u_ca_in_702 = {{10{1'b0}}, col_in_702};
assign u_ca_in_703 = {{10{1'b0}}, col_in_703};
assign u_ca_in_704 = {{10{1'b0}}, col_in_704};
assign u_ca_in_705 = {{10{1'b0}}, col_in_705};
assign u_ca_in_706 = {{10{1'b0}}, col_in_706};
assign u_ca_in_707 = {{10{1'b0}}, col_in_707};
assign u_ca_in_708 = {{10{1'b0}}, col_in_708};
assign u_ca_in_709 = {{10{1'b0}}, col_in_709};
assign u_ca_in_710 = {{10{1'b0}}, col_in_710};
assign u_ca_in_711 = {{10{1'b0}}, col_in_711};
assign u_ca_in_712 = {{10{1'b0}}, col_in_712};
assign u_ca_in_713 = {{10{1'b0}}, col_in_713};
assign u_ca_in_714 = {{10{1'b0}}, col_in_714};
assign u_ca_in_715 = {{10{1'b0}}, col_in_715};
assign u_ca_in_716 = {{10{1'b0}}, col_in_716};
assign u_ca_in_717 = {{10{1'b0}}, col_in_717};
assign u_ca_in_718 = {{10{1'b0}}, col_in_718};
assign u_ca_in_719 = {{10{1'b0}}, col_in_719};
assign u_ca_in_720 = {{10{1'b0}}, col_in_720};
assign u_ca_in_721 = {{10{1'b0}}, col_in_721};
assign u_ca_in_722 = {{10{1'b0}}, col_in_722};
assign u_ca_in_723 = {{10{1'b0}}, col_in_723};
assign u_ca_in_724 = {{10{1'b0}}, col_in_724};
assign u_ca_in_725 = {{10{1'b0}}, col_in_725};
assign u_ca_in_726 = {{10{1'b0}}, col_in_726};
assign u_ca_in_727 = {{10{1'b0}}, col_in_727};
assign u_ca_in_728 = {{10{1'b0}}, col_in_728};
assign u_ca_in_729 = {{10{1'b0}}, col_in_729};
assign u_ca_in_730 = {{10{1'b0}}, col_in_730};
assign u_ca_in_731 = {{10{1'b0}}, col_in_731};
assign u_ca_in_732 = {{10{1'b0}}, col_in_732};
assign u_ca_in_733 = {{10{1'b0}}, col_in_733};
assign u_ca_in_734 = {{10{1'b0}}, col_in_734};
assign u_ca_in_735 = {{10{1'b0}}, col_in_735};
assign u_ca_in_736 = {{10{1'b0}}, col_in_736};
assign u_ca_in_737 = {{10{1'b0}}, col_in_737};
assign u_ca_in_738 = {{10{1'b0}}, col_in_738};
assign u_ca_in_739 = {{10{1'b0}}, col_in_739};
assign u_ca_in_740 = {{10{1'b0}}, col_in_740};
assign u_ca_in_741 = {{10{1'b0}}, col_in_741};
assign u_ca_in_742 = {{10{1'b0}}, col_in_742};
assign u_ca_in_743 = {{10{1'b0}}, col_in_743};
assign u_ca_in_744 = {{10{1'b0}}, col_in_744};
assign u_ca_in_745 = {{10{1'b0}}, col_in_745};
assign u_ca_in_746 = {{10{1'b0}}, col_in_746};
assign u_ca_in_747 = {{10{1'b0}}, col_in_747};
assign u_ca_in_748 = {{10{1'b0}}, col_in_748};
assign u_ca_in_749 = {{10{1'b0}}, col_in_749};
assign u_ca_in_750 = {{10{1'b0}}, col_in_750};
assign u_ca_in_751 = {{10{1'b0}}, col_in_751};
assign u_ca_in_752 = {{10{1'b0}}, col_in_752};
assign u_ca_in_753 = {{10{1'b0}}, col_in_753};
assign u_ca_in_754 = {{10{1'b0}}, col_in_754};
assign u_ca_in_755 = {{10{1'b0}}, col_in_755};
assign u_ca_in_756 = {{10{1'b0}}, col_in_756};
assign u_ca_in_757 = {{10{1'b0}}, col_in_757};
assign u_ca_in_758 = {{10{1'b0}}, col_in_758};
assign u_ca_in_759 = {{10{1'b0}}, col_in_759};
assign u_ca_in_760 = {{10{1'b0}}, col_in_760};
assign u_ca_in_761 = {{10{1'b0}}, col_in_761};
assign u_ca_in_762 = {{10{1'b0}}, col_in_762};
assign u_ca_in_763 = {{10{1'b0}}, col_in_763};
assign u_ca_in_764 = {{10{1'b0}}, col_in_764};
assign u_ca_in_765 = {{10{1'b0}}, col_in_765};
assign u_ca_in_766 = {{10{1'b0}}, col_in_766};
assign u_ca_in_767 = {{10{1'b0}}, col_in_767};
assign u_ca_in_768 = {{10{1'b0}}, col_in_768};
assign u_ca_in_769 = {{10{1'b0}}, col_in_769};
assign u_ca_in_770 = {{10{1'b0}}, col_in_770};
assign u_ca_in_771 = {{10{1'b0}}, col_in_771};
assign u_ca_in_772 = {{10{1'b0}}, col_in_772};
assign u_ca_in_773 = {{10{1'b0}}, col_in_773};
assign u_ca_in_774 = {{10{1'b0}}, col_in_774};
assign u_ca_in_775 = {{10{1'b0}}, col_in_775};
assign u_ca_in_776 = {{10{1'b0}}, col_in_776};
assign u_ca_in_777 = {{10{1'b0}}, col_in_777};
assign u_ca_in_778 = {{10{1'b0}}, col_in_778};
assign u_ca_in_779 = {{10{1'b0}}, col_in_779};
assign u_ca_in_780 = {{10{1'b0}}, col_in_780};
assign u_ca_in_781 = {{10{1'b0}}, col_in_781};
assign u_ca_in_782 = {{10{1'b0}}, col_in_782};
assign u_ca_in_783 = {{10{1'b0}}, col_in_783};
assign u_ca_in_784 = {{10{1'b0}}, col_in_784};
assign u_ca_in_785 = {{10{1'b0}}, col_in_785};
assign u_ca_in_786 = {{10{1'b0}}, col_in_786};
assign u_ca_in_787 = {{10{1'b0}}, col_in_787};
assign u_ca_in_788 = {{10{1'b0}}, col_in_788};
assign u_ca_in_789 = {{10{1'b0}}, col_in_789};
assign u_ca_in_790 = {{10{1'b0}}, col_in_790};
assign u_ca_in_791 = {{10{1'b0}}, col_in_791};
assign u_ca_in_792 = {{10{1'b0}}, col_in_792};
assign u_ca_in_793 = {{10{1'b0}}, col_in_793};
assign u_ca_in_794 = {{10{1'b0}}, col_in_794};
assign u_ca_in_795 = {{10{1'b0}}, col_in_795};
assign u_ca_in_796 = {{10{1'b0}}, col_in_796};
assign u_ca_in_797 = {{10{1'b0}}, col_in_797};
assign u_ca_in_798 = {{10{1'b0}}, col_in_798};
assign u_ca_in_799 = {{10{1'b0}}, col_in_799};
assign u_ca_in_800 = {{10{1'b0}}, col_in_800};
assign u_ca_in_801 = {{10{1'b0}}, col_in_801};
assign u_ca_in_802 = {{10{1'b0}}, col_in_802};
assign u_ca_in_803 = {{10{1'b0}}, col_in_803};
assign u_ca_in_804 = {{10{1'b0}}, col_in_804};
assign u_ca_in_805 = {{10{1'b0}}, col_in_805};
assign u_ca_in_806 = {{10{1'b0}}, col_in_806};
assign u_ca_in_807 = {{10{1'b0}}, col_in_807};
assign u_ca_in_808 = {{10{1'b0}}, col_in_808};
assign u_ca_in_809 = {{10{1'b0}}, col_in_809};
assign u_ca_in_810 = {{10{1'b0}}, col_in_810};
assign u_ca_in_811 = {{10{1'b0}}, col_in_811};
assign u_ca_in_812 = {{10{1'b0}}, col_in_812};
assign u_ca_in_813 = {{10{1'b0}}, col_in_813};
assign u_ca_in_814 = {{10{1'b0}}, col_in_814};
assign u_ca_in_815 = {{10{1'b0}}, col_in_815};
assign u_ca_in_816 = {{10{1'b0}}, col_in_816};
assign u_ca_in_817 = {{10{1'b0}}, col_in_817};
assign u_ca_in_818 = {{10{1'b0}}, col_in_818};
assign u_ca_in_819 = {{10{1'b0}}, col_in_819};
assign u_ca_in_820 = {{10{1'b0}}, col_in_820};
assign u_ca_in_821 = {{10{1'b0}}, col_in_821};
assign u_ca_in_822 = {{10{1'b0}}, col_in_822};
assign u_ca_in_823 = {{10{1'b0}}, col_in_823};
assign u_ca_in_824 = {{10{1'b0}}, col_in_824};
assign u_ca_in_825 = {{10{1'b0}}, col_in_825};
assign u_ca_in_826 = {{10{1'b0}}, col_in_826};
assign u_ca_in_827 = {{10{1'b0}}, col_in_827};
assign u_ca_in_828 = {{10{1'b0}}, col_in_828};
assign u_ca_in_829 = {{10{1'b0}}, col_in_829};
assign u_ca_in_830 = {{10{1'b0}}, col_in_830};
assign u_ca_in_831 = {{10{1'b0}}, col_in_831};
assign u_ca_in_832 = {{10{1'b0}}, col_in_832};
assign u_ca_in_833 = {{10{1'b0}}, col_in_833};
assign u_ca_in_834 = {{10{1'b0}}, col_in_834};
assign u_ca_in_835 = {{10{1'b0}}, col_in_835};
assign u_ca_in_836 = {{10{1'b0}}, col_in_836};
assign u_ca_in_837 = {{10{1'b0}}, col_in_837};
assign u_ca_in_838 = {{10{1'b0}}, col_in_838};
assign u_ca_in_839 = {{10{1'b0}}, col_in_839};
assign u_ca_in_840 = {{10{1'b0}}, col_in_840};
assign u_ca_in_841 = {{10{1'b0}}, col_in_841};
assign u_ca_in_842 = {{10{1'b0}}, col_in_842};
assign u_ca_in_843 = {{10{1'b0}}, col_in_843};
assign u_ca_in_844 = {{10{1'b0}}, col_in_844};
assign u_ca_in_845 = {{10{1'b0}}, col_in_845};
assign u_ca_in_846 = {{10{1'b0}}, col_in_846};
assign u_ca_in_847 = {{10{1'b0}}, col_in_847};
assign u_ca_in_848 = {{10{1'b0}}, col_in_848};
assign u_ca_in_849 = {{10{1'b0}}, col_in_849};
assign u_ca_in_850 = {{10{1'b0}}, col_in_850};
assign u_ca_in_851 = {{10{1'b0}}, col_in_851};
assign u_ca_in_852 = {{10{1'b0}}, col_in_852};
assign u_ca_in_853 = {{10{1'b0}}, col_in_853};
assign u_ca_in_854 = {{10{1'b0}}, col_in_854};
assign u_ca_in_855 = {{10{1'b0}}, col_in_855};
assign u_ca_in_856 = {{10{1'b0}}, col_in_856};
assign u_ca_in_857 = {{10{1'b0}}, col_in_857};
assign u_ca_in_858 = {{10{1'b0}}, col_in_858};
assign u_ca_in_859 = {{10{1'b0}}, col_in_859};
assign u_ca_in_860 = {{10{1'b0}}, col_in_860};
assign u_ca_in_861 = {{10{1'b0}}, col_in_861};
assign u_ca_in_862 = {{10{1'b0}}, col_in_862};
assign u_ca_in_863 = {{10{1'b0}}, col_in_863};
assign u_ca_in_864 = {{10{1'b0}}, col_in_864};
assign u_ca_in_865 = {{10{1'b0}}, col_in_865};
assign u_ca_in_866 = {{10{1'b0}}, col_in_866};
assign u_ca_in_867 = {{10{1'b0}}, col_in_867};
assign u_ca_in_868 = {{10{1'b0}}, col_in_868};
assign u_ca_in_869 = {{10{1'b0}}, col_in_869};
assign u_ca_in_870 = {{10{1'b0}}, col_in_870};
assign u_ca_in_871 = {{10{1'b0}}, col_in_871};
assign u_ca_in_872 = {{10{1'b0}}, col_in_872};
assign u_ca_in_873 = {{10{1'b0}}, col_in_873};
assign u_ca_in_874 = {{10{1'b0}}, col_in_874};
assign u_ca_in_875 = {{10{1'b0}}, col_in_875};
assign u_ca_in_876 = {{10{1'b0}}, col_in_876};
assign u_ca_in_877 = {{10{1'b0}}, col_in_877};
assign u_ca_in_878 = {{10{1'b0}}, col_in_878};
assign u_ca_in_879 = {{10{1'b0}}, col_in_879};
assign u_ca_in_880 = {{10{1'b0}}, col_in_880};
assign u_ca_in_881 = {{10{1'b0}}, col_in_881};
assign u_ca_in_882 = {{10{1'b0}}, col_in_882};
assign u_ca_in_883 = {{10{1'b0}}, col_in_883};
assign u_ca_in_884 = {{10{1'b0}}, col_in_884};
assign u_ca_in_885 = {{10{1'b0}}, col_in_885};
assign u_ca_in_886 = {{10{1'b0}}, col_in_886};
assign u_ca_in_887 = {{10{1'b0}}, col_in_887};
assign u_ca_in_888 = {{10{1'b0}}, col_in_888};
assign u_ca_in_889 = {{10{1'b0}}, col_in_889};
assign u_ca_in_890 = {{10{1'b0}}, col_in_890};
assign u_ca_in_891 = {{10{1'b0}}, col_in_891};
assign u_ca_in_892 = {{10{1'b0}}, col_in_892};
assign u_ca_in_893 = {{10{1'b0}}, col_in_893};
assign u_ca_in_894 = {{10{1'b0}}, col_in_894};
assign u_ca_in_895 = {{10{1'b0}}, col_in_895};
assign u_ca_in_896 = {{10{1'b0}}, col_in_896};
assign u_ca_in_897 = {{10{1'b0}}, col_in_897};
assign u_ca_in_898 = {{10{1'b0}}, col_in_898};
assign u_ca_in_899 = {{10{1'b0}}, col_in_899};
assign u_ca_in_900 = {{10{1'b0}}, col_in_900};
assign u_ca_in_901 = {{10{1'b0}}, col_in_901};
assign u_ca_in_902 = {{10{1'b0}}, col_in_902};
assign u_ca_in_903 = {{10{1'b0}}, col_in_903};
assign u_ca_in_904 = {{10{1'b0}}, col_in_904};
assign u_ca_in_905 = {{10{1'b0}}, col_in_905};
assign u_ca_in_906 = {{10{1'b0}}, col_in_906};
assign u_ca_in_907 = {{10{1'b0}}, col_in_907};
assign u_ca_in_908 = {{10{1'b0}}, col_in_908};
assign u_ca_in_909 = {{10{1'b0}}, col_in_909};
assign u_ca_in_910 = {{10{1'b0}}, col_in_910};
assign u_ca_in_911 = {{10{1'b0}}, col_in_911};
assign u_ca_in_912 = {{10{1'b0}}, col_in_912};
assign u_ca_in_913 = {{10{1'b0}}, col_in_913};
assign u_ca_in_914 = {{10{1'b0}}, col_in_914};
assign u_ca_in_915 = {{10{1'b0}}, col_in_915};
assign u_ca_in_916 = {{10{1'b0}}, col_in_916};
assign u_ca_in_917 = {{10{1'b0}}, col_in_917};
assign u_ca_in_918 = {{10{1'b0}}, col_in_918};
assign u_ca_in_919 = {{10{1'b0}}, col_in_919};
assign u_ca_in_920 = {{10{1'b0}}, col_in_920};
assign u_ca_in_921 = {{10{1'b0}}, col_in_921};
assign u_ca_in_922 = {{10{1'b0}}, col_in_922};
assign u_ca_in_923 = {{10{1'b0}}, col_in_923};
assign u_ca_in_924 = {{10{1'b0}}, col_in_924};
assign u_ca_in_925 = {{10{1'b0}}, col_in_925};
assign u_ca_in_926 = {{10{1'b0}}, col_in_926};
assign u_ca_in_927 = {{10{1'b0}}, col_in_927};
assign u_ca_in_928 = {{10{1'b0}}, col_in_928};
assign u_ca_in_929 = {{10{1'b0}}, col_in_929};
assign u_ca_in_930 = {{10{1'b0}}, col_in_930};
assign u_ca_in_931 = {{10{1'b0}}, col_in_931};
assign u_ca_in_932 = {{10{1'b0}}, col_in_932};
assign u_ca_in_933 = {{10{1'b0}}, col_in_933};
assign u_ca_in_934 = {{10{1'b0}}, col_in_934};
assign u_ca_in_935 = {{10{1'b0}}, col_in_935};
assign u_ca_in_936 = {{10{1'b0}}, col_in_936};
assign u_ca_in_937 = {{10{1'b0}}, col_in_937};
assign u_ca_in_938 = {{10{1'b0}}, col_in_938};
assign u_ca_in_939 = {{10{1'b0}}, col_in_939};
assign u_ca_in_940 = {{10{1'b0}}, col_in_940};
assign u_ca_in_941 = {{10{1'b0}}, col_in_941};
assign u_ca_in_942 = {{10{1'b0}}, col_in_942};
assign u_ca_in_943 = {{10{1'b0}}, col_in_943};
assign u_ca_in_944 = {{10{1'b0}}, col_in_944};
assign u_ca_in_945 = {{10{1'b0}}, col_in_945};
assign u_ca_in_946 = {{10{1'b0}}, col_in_946};
assign u_ca_in_947 = {{10{1'b0}}, col_in_947};
assign u_ca_in_948 = {{10{1'b0}}, col_in_948};
assign u_ca_in_949 = {{10{1'b0}}, col_in_949};
assign u_ca_in_950 = {{10{1'b0}}, col_in_950};
assign u_ca_in_951 = {{10{1'b0}}, col_in_951};
assign u_ca_in_952 = {{10{1'b0}}, col_in_952};
assign u_ca_in_953 = {{10{1'b0}}, col_in_953};
assign u_ca_in_954 = {{10{1'b0}}, col_in_954};
assign u_ca_in_955 = {{10{1'b0}}, col_in_955};
assign u_ca_in_956 = {{10{1'b0}}, col_in_956};
assign u_ca_in_957 = {{10{1'b0}}, col_in_957};
assign u_ca_in_958 = {{10{1'b0}}, col_in_958};
assign u_ca_in_959 = {{10{1'b0}}, col_in_959};
assign u_ca_in_960 = {{10{1'b0}}, col_in_960};
assign u_ca_in_961 = {{10{1'b0}}, col_in_961};
assign u_ca_in_962 = {{10{1'b0}}, col_in_962};
assign u_ca_in_963 = {{10{1'b0}}, col_in_963};
assign u_ca_in_964 = {{10{1'b0}}, col_in_964};
assign u_ca_in_965 = {{10{1'b0}}, col_in_965};
assign u_ca_in_966 = {{10{1'b0}}, col_in_966};
assign u_ca_in_967 = {{10{1'b0}}, col_in_967};
assign u_ca_in_968 = {{10{1'b0}}, col_in_968};
assign u_ca_in_969 = {{10{1'b0}}, col_in_969};
assign u_ca_in_970 = {{10{1'b0}}, col_in_970};
assign u_ca_in_971 = {{10{1'b0}}, col_in_971};
assign u_ca_in_972 = {{10{1'b0}}, col_in_972};
assign u_ca_in_973 = {{10{1'b0}}, col_in_973};
assign u_ca_in_974 = {{10{1'b0}}, col_in_974};
assign u_ca_in_975 = {{10{1'b0}}, col_in_975};
assign u_ca_in_976 = {{10{1'b0}}, col_in_976};
assign u_ca_in_977 = {{10{1'b0}}, col_in_977};
assign u_ca_in_978 = {{10{1'b0}}, col_in_978};
assign u_ca_in_979 = {{10{1'b0}}, col_in_979};
assign u_ca_in_980 = {{10{1'b0}}, col_in_980};
assign u_ca_in_981 = {{10{1'b0}}, col_in_981};
assign u_ca_in_982 = {{10{1'b0}}, col_in_982};
assign u_ca_in_983 = {{10{1'b0}}, col_in_983};
assign u_ca_in_984 = {{10{1'b0}}, col_in_984};
assign u_ca_in_985 = {{10{1'b0}}, col_in_985};
assign u_ca_in_986 = {{10{1'b0}}, col_in_986};
assign u_ca_in_987 = {{10{1'b0}}, col_in_987};
assign u_ca_in_988 = {{10{1'b0}}, col_in_988};
assign u_ca_in_989 = {{10{1'b0}}, col_in_989};
assign u_ca_in_990 = {{10{1'b0}}, col_in_990};
assign u_ca_in_991 = {{10{1'b0}}, col_in_991};
assign u_ca_in_992 = {{10{1'b0}}, col_in_992};
assign u_ca_in_993 = {{10{1'b0}}, col_in_993};
assign u_ca_in_994 = {{10{1'b0}}, col_in_994};
assign u_ca_in_995 = {{10{1'b0}}, col_in_995};
assign u_ca_in_996 = {{10{1'b0}}, col_in_996};
assign u_ca_in_997 = {{10{1'b0}}, col_in_997};
assign u_ca_in_998 = {{10{1'b0}}, col_in_998};
assign u_ca_in_999 = {{10{1'b0}}, col_in_999};
assign u_ca_in_1000 = {{10{1'b0}}, col_in_1000};
assign u_ca_in_1001 = {{10{1'b0}}, col_in_1001};
assign u_ca_in_1002 = {{10{1'b0}}, col_in_1002};
assign u_ca_in_1003 = {{10{1'b0}}, col_in_1003};
assign u_ca_in_1004 = {{10{1'b0}}, col_in_1004};
assign u_ca_in_1005 = {{10{1'b0}}, col_in_1005};
assign u_ca_in_1006 = {{10{1'b0}}, col_in_1006};
assign u_ca_in_1007 = {{10{1'b0}}, col_in_1007};
assign u_ca_in_1008 = {{10{1'b0}}, col_in_1008};
assign u_ca_in_1009 = {{10{1'b0}}, col_in_1009};
assign u_ca_in_1010 = {{10{1'b0}}, col_in_1010};
assign u_ca_in_1011 = {{10{1'b0}}, col_in_1011};
assign u_ca_in_1012 = {{10{1'b0}}, col_in_1012};
assign u_ca_in_1013 = {{10{1'b0}}, col_in_1013};
assign u_ca_in_1014 = {{10{1'b0}}, col_in_1014};
assign u_ca_in_1015 = {{10{1'b0}}, col_in_1015};
assign u_ca_in_1016 = {{10{1'b0}}, col_in_1016};
assign u_ca_in_1017 = {{10{1'b0}}, col_in_1017};
assign u_ca_in_1018 = {{10{1'b0}}, col_in_1018};
assign u_ca_in_1019 = {{10{1'b0}}, col_in_1019};
assign u_ca_in_1020 = {{10{1'b0}}, col_in_1020};
assign u_ca_in_1021 = {{10{1'b0}}, col_in_1021};
assign u_ca_in_1022 = {{10{1'b0}}, col_in_1022};
assign u_ca_in_1023 = {{10{1'b0}}, col_in_1023};
assign u_ca_in_1024 = {{10{1'b0}}, col_in_1024};
assign u_ca_in_1025 = {{10{1'b0}}, col_in_1025};
assign u_ca_in_1026 = {{10{1'b0}}, col_in_1026};

//---------------------------------------------------------



//--compressor_array---------------------------------------
compressor_162_48 u_ca_162_48_0(.d_in(u_ca_in_0), .d_out(u_ca_out_0));
compressor_162_48 u_ca_162_48_1(.d_in(u_ca_in_1), .d_out(u_ca_out_1));
compressor_162_48 u_ca_162_48_2(.d_in(u_ca_in_2), .d_out(u_ca_out_2));
compressor_162_48 u_ca_162_48_3(.d_in(u_ca_in_3), .d_out(u_ca_out_3));
compressor_162_48 u_ca_162_48_4(.d_in(u_ca_in_4), .d_out(u_ca_out_4));
compressor_162_48 u_ca_162_48_5(.d_in(u_ca_in_5), .d_out(u_ca_out_5));
compressor_162_48 u_ca_162_48_6(.d_in(u_ca_in_6), .d_out(u_ca_out_6));
compressor_162_48 u_ca_162_48_7(.d_in(u_ca_in_7), .d_out(u_ca_out_7));
compressor_162_48 u_ca_162_48_8(.d_in(u_ca_in_8), .d_out(u_ca_out_8));
compressor_162_48 u_ca_162_48_9(.d_in(u_ca_in_9), .d_out(u_ca_out_9));
compressor_162_48 u_ca_162_48_10(.d_in(u_ca_in_10), .d_out(u_ca_out_10));
compressor_162_48 u_ca_162_48_11(.d_in(u_ca_in_11), .d_out(u_ca_out_11));
compressor_162_48 u_ca_162_48_12(.d_in(u_ca_in_12), .d_out(u_ca_out_12));
compressor_162_48 u_ca_162_48_13(.d_in(u_ca_in_13), .d_out(u_ca_out_13));
compressor_162_48 u_ca_162_48_14(.d_in(u_ca_in_14), .d_out(u_ca_out_14));
compressor_162_48 u_ca_162_48_15(.d_in(u_ca_in_15), .d_out(u_ca_out_15));
compressor_162_48 u_ca_162_48_16(.d_in(u_ca_in_16), .d_out(u_ca_out_16));
compressor_162_48 u_ca_162_48_17(.d_in(u_ca_in_17), .d_out(u_ca_out_17));
compressor_162_48 u_ca_162_48_18(.d_in(u_ca_in_18), .d_out(u_ca_out_18));
compressor_162_48 u_ca_162_48_19(.d_in(u_ca_in_19), .d_out(u_ca_out_19));
compressor_162_48 u_ca_162_48_20(.d_in(u_ca_in_20), .d_out(u_ca_out_20));
compressor_162_48 u_ca_162_48_21(.d_in(u_ca_in_21), .d_out(u_ca_out_21));
compressor_162_48 u_ca_162_48_22(.d_in(u_ca_in_22), .d_out(u_ca_out_22));
compressor_162_48 u_ca_162_48_23(.d_in(u_ca_in_23), .d_out(u_ca_out_23));
compressor_162_48 u_ca_162_48_24(.d_in(u_ca_in_24), .d_out(u_ca_out_24));
compressor_162_48 u_ca_162_48_25(.d_in(u_ca_in_25), .d_out(u_ca_out_25));
compressor_162_48 u_ca_162_48_26(.d_in(u_ca_in_26), .d_out(u_ca_out_26));
compressor_162_48 u_ca_162_48_27(.d_in(u_ca_in_27), .d_out(u_ca_out_27));
compressor_162_48 u_ca_162_48_28(.d_in(u_ca_in_28), .d_out(u_ca_out_28));
compressor_162_48 u_ca_162_48_29(.d_in(u_ca_in_29), .d_out(u_ca_out_29));
compressor_162_48 u_ca_162_48_30(.d_in(u_ca_in_30), .d_out(u_ca_out_30));
compressor_162_48 u_ca_162_48_31(.d_in(u_ca_in_31), .d_out(u_ca_out_31));
compressor_162_48 u_ca_162_48_32(.d_in(u_ca_in_32), .d_out(u_ca_out_32));
compressor_162_48 u_ca_162_48_33(.d_in(u_ca_in_33), .d_out(u_ca_out_33));
compressor_162_48 u_ca_162_48_34(.d_in(u_ca_in_34), .d_out(u_ca_out_34));
compressor_162_48 u_ca_162_48_35(.d_in(u_ca_in_35), .d_out(u_ca_out_35));
compressor_162_48 u_ca_162_48_36(.d_in(u_ca_in_36), .d_out(u_ca_out_36));
compressor_162_48 u_ca_162_48_37(.d_in(u_ca_in_37), .d_out(u_ca_out_37));
compressor_162_48 u_ca_162_48_38(.d_in(u_ca_in_38), .d_out(u_ca_out_38));
compressor_162_48 u_ca_162_48_39(.d_in(u_ca_in_39), .d_out(u_ca_out_39));
compressor_162_48 u_ca_162_48_40(.d_in(u_ca_in_40), .d_out(u_ca_out_40));
compressor_162_48 u_ca_162_48_41(.d_in(u_ca_in_41), .d_out(u_ca_out_41));
compressor_162_48 u_ca_162_48_42(.d_in(u_ca_in_42), .d_out(u_ca_out_42));
compressor_162_48 u_ca_162_48_43(.d_in(u_ca_in_43), .d_out(u_ca_out_43));
compressor_162_48 u_ca_162_48_44(.d_in(u_ca_in_44), .d_out(u_ca_out_44));
compressor_162_48 u_ca_162_48_45(.d_in(u_ca_in_45), .d_out(u_ca_out_45));
compressor_162_48 u_ca_162_48_46(.d_in(u_ca_in_46), .d_out(u_ca_out_46));
compressor_162_48 u_ca_162_48_47(.d_in(u_ca_in_47), .d_out(u_ca_out_47));
compressor_162_48 u_ca_162_48_48(.d_in(u_ca_in_48), .d_out(u_ca_out_48));
compressor_162_48 u_ca_162_48_49(.d_in(u_ca_in_49), .d_out(u_ca_out_49));
compressor_162_48 u_ca_162_48_50(.d_in(u_ca_in_50), .d_out(u_ca_out_50));
compressor_162_48 u_ca_162_48_51(.d_in(u_ca_in_51), .d_out(u_ca_out_51));
compressor_162_48 u_ca_162_48_52(.d_in(u_ca_in_52), .d_out(u_ca_out_52));
compressor_162_48 u_ca_162_48_53(.d_in(u_ca_in_53), .d_out(u_ca_out_53));
compressor_162_48 u_ca_162_48_54(.d_in(u_ca_in_54), .d_out(u_ca_out_54));
compressor_162_48 u_ca_162_48_55(.d_in(u_ca_in_55), .d_out(u_ca_out_55));
compressor_162_48 u_ca_162_48_56(.d_in(u_ca_in_56), .d_out(u_ca_out_56));
compressor_162_48 u_ca_162_48_57(.d_in(u_ca_in_57), .d_out(u_ca_out_57));
compressor_162_48 u_ca_162_48_58(.d_in(u_ca_in_58), .d_out(u_ca_out_58));
compressor_162_48 u_ca_162_48_59(.d_in(u_ca_in_59), .d_out(u_ca_out_59));
compressor_162_48 u_ca_162_48_60(.d_in(u_ca_in_60), .d_out(u_ca_out_60));
compressor_162_48 u_ca_162_48_61(.d_in(u_ca_in_61), .d_out(u_ca_out_61));
compressor_162_48 u_ca_162_48_62(.d_in(u_ca_in_62), .d_out(u_ca_out_62));
compressor_162_48 u_ca_162_48_63(.d_in(u_ca_in_63), .d_out(u_ca_out_63));
compressor_162_48 u_ca_162_48_64(.d_in(u_ca_in_64), .d_out(u_ca_out_64));
compressor_162_48 u_ca_162_48_65(.d_in(u_ca_in_65), .d_out(u_ca_out_65));
compressor_162_48 u_ca_162_48_66(.d_in(u_ca_in_66), .d_out(u_ca_out_66));
compressor_162_48 u_ca_162_48_67(.d_in(u_ca_in_67), .d_out(u_ca_out_67));
compressor_162_48 u_ca_162_48_68(.d_in(u_ca_in_68), .d_out(u_ca_out_68));
compressor_162_48 u_ca_162_48_69(.d_in(u_ca_in_69), .d_out(u_ca_out_69));
compressor_162_48 u_ca_162_48_70(.d_in(u_ca_in_70), .d_out(u_ca_out_70));
compressor_162_48 u_ca_162_48_71(.d_in(u_ca_in_71), .d_out(u_ca_out_71));
compressor_162_48 u_ca_162_48_72(.d_in(u_ca_in_72), .d_out(u_ca_out_72));
compressor_162_48 u_ca_162_48_73(.d_in(u_ca_in_73), .d_out(u_ca_out_73));
compressor_162_48 u_ca_162_48_74(.d_in(u_ca_in_74), .d_out(u_ca_out_74));
compressor_162_48 u_ca_162_48_75(.d_in(u_ca_in_75), .d_out(u_ca_out_75));
compressor_162_48 u_ca_162_48_76(.d_in(u_ca_in_76), .d_out(u_ca_out_76));
compressor_162_48 u_ca_162_48_77(.d_in(u_ca_in_77), .d_out(u_ca_out_77));
compressor_162_48 u_ca_162_48_78(.d_in(u_ca_in_78), .d_out(u_ca_out_78));
compressor_162_48 u_ca_162_48_79(.d_in(u_ca_in_79), .d_out(u_ca_out_79));
compressor_162_48 u_ca_162_48_80(.d_in(u_ca_in_80), .d_out(u_ca_out_80));
compressor_162_48 u_ca_162_48_81(.d_in(u_ca_in_81), .d_out(u_ca_out_81));
compressor_162_48 u_ca_162_48_82(.d_in(u_ca_in_82), .d_out(u_ca_out_82));
compressor_162_48 u_ca_162_48_83(.d_in(u_ca_in_83), .d_out(u_ca_out_83));
compressor_162_48 u_ca_162_48_84(.d_in(u_ca_in_84), .d_out(u_ca_out_84));
compressor_162_48 u_ca_162_48_85(.d_in(u_ca_in_85), .d_out(u_ca_out_85));
compressor_162_48 u_ca_162_48_86(.d_in(u_ca_in_86), .d_out(u_ca_out_86));
compressor_162_48 u_ca_162_48_87(.d_in(u_ca_in_87), .d_out(u_ca_out_87));
compressor_162_48 u_ca_162_48_88(.d_in(u_ca_in_88), .d_out(u_ca_out_88));
compressor_162_48 u_ca_162_48_89(.d_in(u_ca_in_89), .d_out(u_ca_out_89));
compressor_162_48 u_ca_162_48_90(.d_in(u_ca_in_90), .d_out(u_ca_out_90));
compressor_162_48 u_ca_162_48_91(.d_in(u_ca_in_91), .d_out(u_ca_out_91));
compressor_162_48 u_ca_162_48_92(.d_in(u_ca_in_92), .d_out(u_ca_out_92));
compressor_162_48 u_ca_162_48_93(.d_in(u_ca_in_93), .d_out(u_ca_out_93));
compressor_162_48 u_ca_162_48_94(.d_in(u_ca_in_94), .d_out(u_ca_out_94));
compressor_162_48 u_ca_162_48_95(.d_in(u_ca_in_95), .d_out(u_ca_out_95));
compressor_162_48 u_ca_162_48_96(.d_in(u_ca_in_96), .d_out(u_ca_out_96));
compressor_162_48 u_ca_162_48_97(.d_in(u_ca_in_97), .d_out(u_ca_out_97));
compressor_162_48 u_ca_162_48_98(.d_in(u_ca_in_98), .d_out(u_ca_out_98));
compressor_162_48 u_ca_162_48_99(.d_in(u_ca_in_99), .d_out(u_ca_out_99));
compressor_162_48 u_ca_162_48_100(.d_in(u_ca_in_100), .d_out(u_ca_out_100));
compressor_162_48 u_ca_162_48_101(.d_in(u_ca_in_101), .d_out(u_ca_out_101));
compressor_162_48 u_ca_162_48_102(.d_in(u_ca_in_102), .d_out(u_ca_out_102));
compressor_162_48 u_ca_162_48_103(.d_in(u_ca_in_103), .d_out(u_ca_out_103));
compressor_162_48 u_ca_162_48_104(.d_in(u_ca_in_104), .d_out(u_ca_out_104));
compressor_162_48 u_ca_162_48_105(.d_in(u_ca_in_105), .d_out(u_ca_out_105));
compressor_162_48 u_ca_162_48_106(.d_in(u_ca_in_106), .d_out(u_ca_out_106));
compressor_162_48 u_ca_162_48_107(.d_in(u_ca_in_107), .d_out(u_ca_out_107));
compressor_162_48 u_ca_162_48_108(.d_in(u_ca_in_108), .d_out(u_ca_out_108));
compressor_162_48 u_ca_162_48_109(.d_in(u_ca_in_109), .d_out(u_ca_out_109));
compressor_162_48 u_ca_162_48_110(.d_in(u_ca_in_110), .d_out(u_ca_out_110));
compressor_162_48 u_ca_162_48_111(.d_in(u_ca_in_111), .d_out(u_ca_out_111));
compressor_162_48 u_ca_162_48_112(.d_in(u_ca_in_112), .d_out(u_ca_out_112));
compressor_162_48 u_ca_162_48_113(.d_in(u_ca_in_113), .d_out(u_ca_out_113));
compressor_162_48 u_ca_162_48_114(.d_in(u_ca_in_114), .d_out(u_ca_out_114));
compressor_162_48 u_ca_162_48_115(.d_in(u_ca_in_115), .d_out(u_ca_out_115));
compressor_162_48 u_ca_162_48_116(.d_in(u_ca_in_116), .d_out(u_ca_out_116));
compressor_162_48 u_ca_162_48_117(.d_in(u_ca_in_117), .d_out(u_ca_out_117));
compressor_162_48 u_ca_162_48_118(.d_in(u_ca_in_118), .d_out(u_ca_out_118));
compressor_162_48 u_ca_162_48_119(.d_in(u_ca_in_119), .d_out(u_ca_out_119));
compressor_162_48 u_ca_162_48_120(.d_in(u_ca_in_120), .d_out(u_ca_out_120));
compressor_162_48 u_ca_162_48_121(.d_in(u_ca_in_121), .d_out(u_ca_out_121));
compressor_162_48 u_ca_162_48_122(.d_in(u_ca_in_122), .d_out(u_ca_out_122));
compressor_162_48 u_ca_162_48_123(.d_in(u_ca_in_123), .d_out(u_ca_out_123));
compressor_162_48 u_ca_162_48_124(.d_in(u_ca_in_124), .d_out(u_ca_out_124));
compressor_162_48 u_ca_162_48_125(.d_in(u_ca_in_125), .d_out(u_ca_out_125));
compressor_162_48 u_ca_162_48_126(.d_in(u_ca_in_126), .d_out(u_ca_out_126));
compressor_162_48 u_ca_162_48_127(.d_in(u_ca_in_127), .d_out(u_ca_out_127));
compressor_162_48 u_ca_162_48_128(.d_in(u_ca_in_128), .d_out(u_ca_out_128));
compressor_162_48 u_ca_162_48_129(.d_in(u_ca_in_129), .d_out(u_ca_out_129));
compressor_162_48 u_ca_162_48_130(.d_in(u_ca_in_130), .d_out(u_ca_out_130));
compressor_162_48 u_ca_162_48_131(.d_in(u_ca_in_131), .d_out(u_ca_out_131));
compressor_162_48 u_ca_162_48_132(.d_in(u_ca_in_132), .d_out(u_ca_out_132));
compressor_162_48 u_ca_162_48_133(.d_in(u_ca_in_133), .d_out(u_ca_out_133));
compressor_162_48 u_ca_162_48_134(.d_in(u_ca_in_134), .d_out(u_ca_out_134));
compressor_162_48 u_ca_162_48_135(.d_in(u_ca_in_135), .d_out(u_ca_out_135));
compressor_162_48 u_ca_162_48_136(.d_in(u_ca_in_136), .d_out(u_ca_out_136));
compressor_162_48 u_ca_162_48_137(.d_in(u_ca_in_137), .d_out(u_ca_out_137));
compressor_162_48 u_ca_162_48_138(.d_in(u_ca_in_138), .d_out(u_ca_out_138));
compressor_162_48 u_ca_162_48_139(.d_in(u_ca_in_139), .d_out(u_ca_out_139));
compressor_162_48 u_ca_162_48_140(.d_in(u_ca_in_140), .d_out(u_ca_out_140));
compressor_162_48 u_ca_162_48_141(.d_in(u_ca_in_141), .d_out(u_ca_out_141));
compressor_162_48 u_ca_162_48_142(.d_in(u_ca_in_142), .d_out(u_ca_out_142));
compressor_162_48 u_ca_162_48_143(.d_in(u_ca_in_143), .d_out(u_ca_out_143));
compressor_162_48 u_ca_162_48_144(.d_in(u_ca_in_144), .d_out(u_ca_out_144));
compressor_162_48 u_ca_162_48_145(.d_in(u_ca_in_145), .d_out(u_ca_out_145));
compressor_162_48 u_ca_162_48_146(.d_in(u_ca_in_146), .d_out(u_ca_out_146));
compressor_162_48 u_ca_162_48_147(.d_in(u_ca_in_147), .d_out(u_ca_out_147));
compressor_162_48 u_ca_162_48_148(.d_in(u_ca_in_148), .d_out(u_ca_out_148));
compressor_162_48 u_ca_162_48_149(.d_in(u_ca_in_149), .d_out(u_ca_out_149));
compressor_162_48 u_ca_162_48_150(.d_in(u_ca_in_150), .d_out(u_ca_out_150));
compressor_162_48 u_ca_162_48_151(.d_in(u_ca_in_151), .d_out(u_ca_out_151));
compressor_162_48 u_ca_162_48_152(.d_in(u_ca_in_152), .d_out(u_ca_out_152));
compressor_162_48 u_ca_162_48_153(.d_in(u_ca_in_153), .d_out(u_ca_out_153));
compressor_162_48 u_ca_162_48_154(.d_in(u_ca_in_154), .d_out(u_ca_out_154));
compressor_162_48 u_ca_162_48_155(.d_in(u_ca_in_155), .d_out(u_ca_out_155));
compressor_162_48 u_ca_162_48_156(.d_in(u_ca_in_156), .d_out(u_ca_out_156));
compressor_162_48 u_ca_162_48_157(.d_in(u_ca_in_157), .d_out(u_ca_out_157));
compressor_162_48 u_ca_162_48_158(.d_in(u_ca_in_158), .d_out(u_ca_out_158));
compressor_162_48 u_ca_162_48_159(.d_in(u_ca_in_159), .d_out(u_ca_out_159));
compressor_162_48 u_ca_162_48_160(.d_in(u_ca_in_160), .d_out(u_ca_out_160));
compressor_162_48 u_ca_162_48_161(.d_in(u_ca_in_161), .d_out(u_ca_out_161));
compressor_162_48 u_ca_162_48_162(.d_in(u_ca_in_162), .d_out(u_ca_out_162));
compressor_162_48 u_ca_162_48_163(.d_in(u_ca_in_163), .d_out(u_ca_out_163));
compressor_162_48 u_ca_162_48_164(.d_in(u_ca_in_164), .d_out(u_ca_out_164));
compressor_162_48 u_ca_162_48_165(.d_in(u_ca_in_165), .d_out(u_ca_out_165));
compressor_162_48 u_ca_162_48_166(.d_in(u_ca_in_166), .d_out(u_ca_out_166));
compressor_162_48 u_ca_162_48_167(.d_in(u_ca_in_167), .d_out(u_ca_out_167));
compressor_162_48 u_ca_162_48_168(.d_in(u_ca_in_168), .d_out(u_ca_out_168));
compressor_162_48 u_ca_162_48_169(.d_in(u_ca_in_169), .d_out(u_ca_out_169));
compressor_162_48 u_ca_162_48_170(.d_in(u_ca_in_170), .d_out(u_ca_out_170));
compressor_162_48 u_ca_162_48_171(.d_in(u_ca_in_171), .d_out(u_ca_out_171));
compressor_162_48 u_ca_162_48_172(.d_in(u_ca_in_172), .d_out(u_ca_out_172));
compressor_162_48 u_ca_162_48_173(.d_in(u_ca_in_173), .d_out(u_ca_out_173));
compressor_162_48 u_ca_162_48_174(.d_in(u_ca_in_174), .d_out(u_ca_out_174));
compressor_162_48 u_ca_162_48_175(.d_in(u_ca_in_175), .d_out(u_ca_out_175));
compressor_162_48 u_ca_162_48_176(.d_in(u_ca_in_176), .d_out(u_ca_out_176));
compressor_162_48 u_ca_162_48_177(.d_in(u_ca_in_177), .d_out(u_ca_out_177));
compressor_162_48 u_ca_162_48_178(.d_in(u_ca_in_178), .d_out(u_ca_out_178));
compressor_162_48 u_ca_162_48_179(.d_in(u_ca_in_179), .d_out(u_ca_out_179));
compressor_162_48 u_ca_162_48_180(.d_in(u_ca_in_180), .d_out(u_ca_out_180));
compressor_162_48 u_ca_162_48_181(.d_in(u_ca_in_181), .d_out(u_ca_out_181));
compressor_162_48 u_ca_162_48_182(.d_in(u_ca_in_182), .d_out(u_ca_out_182));
compressor_162_48 u_ca_162_48_183(.d_in(u_ca_in_183), .d_out(u_ca_out_183));
compressor_162_48 u_ca_162_48_184(.d_in(u_ca_in_184), .d_out(u_ca_out_184));
compressor_162_48 u_ca_162_48_185(.d_in(u_ca_in_185), .d_out(u_ca_out_185));
compressor_162_48 u_ca_162_48_186(.d_in(u_ca_in_186), .d_out(u_ca_out_186));
compressor_162_48 u_ca_162_48_187(.d_in(u_ca_in_187), .d_out(u_ca_out_187));
compressor_162_48 u_ca_162_48_188(.d_in(u_ca_in_188), .d_out(u_ca_out_188));
compressor_162_48 u_ca_162_48_189(.d_in(u_ca_in_189), .d_out(u_ca_out_189));
compressor_162_48 u_ca_162_48_190(.d_in(u_ca_in_190), .d_out(u_ca_out_190));
compressor_162_48 u_ca_162_48_191(.d_in(u_ca_in_191), .d_out(u_ca_out_191));
compressor_162_48 u_ca_162_48_192(.d_in(u_ca_in_192), .d_out(u_ca_out_192));
compressor_162_48 u_ca_162_48_193(.d_in(u_ca_in_193), .d_out(u_ca_out_193));
compressor_162_48 u_ca_162_48_194(.d_in(u_ca_in_194), .d_out(u_ca_out_194));
compressor_162_48 u_ca_162_48_195(.d_in(u_ca_in_195), .d_out(u_ca_out_195));
compressor_162_48 u_ca_162_48_196(.d_in(u_ca_in_196), .d_out(u_ca_out_196));
compressor_162_48 u_ca_162_48_197(.d_in(u_ca_in_197), .d_out(u_ca_out_197));
compressor_162_48 u_ca_162_48_198(.d_in(u_ca_in_198), .d_out(u_ca_out_198));
compressor_162_48 u_ca_162_48_199(.d_in(u_ca_in_199), .d_out(u_ca_out_199));
compressor_162_48 u_ca_162_48_200(.d_in(u_ca_in_200), .d_out(u_ca_out_200));
compressor_162_48 u_ca_162_48_201(.d_in(u_ca_in_201), .d_out(u_ca_out_201));
compressor_162_48 u_ca_162_48_202(.d_in(u_ca_in_202), .d_out(u_ca_out_202));
compressor_162_48 u_ca_162_48_203(.d_in(u_ca_in_203), .d_out(u_ca_out_203));
compressor_162_48 u_ca_162_48_204(.d_in(u_ca_in_204), .d_out(u_ca_out_204));
compressor_162_48 u_ca_162_48_205(.d_in(u_ca_in_205), .d_out(u_ca_out_205));
compressor_162_48 u_ca_162_48_206(.d_in(u_ca_in_206), .d_out(u_ca_out_206));
compressor_162_48 u_ca_162_48_207(.d_in(u_ca_in_207), .d_out(u_ca_out_207));
compressor_162_48 u_ca_162_48_208(.d_in(u_ca_in_208), .d_out(u_ca_out_208));
compressor_162_48 u_ca_162_48_209(.d_in(u_ca_in_209), .d_out(u_ca_out_209));
compressor_162_48 u_ca_162_48_210(.d_in(u_ca_in_210), .d_out(u_ca_out_210));
compressor_162_48 u_ca_162_48_211(.d_in(u_ca_in_211), .d_out(u_ca_out_211));
compressor_162_48 u_ca_162_48_212(.d_in(u_ca_in_212), .d_out(u_ca_out_212));
compressor_162_48 u_ca_162_48_213(.d_in(u_ca_in_213), .d_out(u_ca_out_213));
compressor_162_48 u_ca_162_48_214(.d_in(u_ca_in_214), .d_out(u_ca_out_214));
compressor_162_48 u_ca_162_48_215(.d_in(u_ca_in_215), .d_out(u_ca_out_215));
compressor_162_48 u_ca_162_48_216(.d_in(u_ca_in_216), .d_out(u_ca_out_216));
compressor_162_48 u_ca_162_48_217(.d_in(u_ca_in_217), .d_out(u_ca_out_217));
compressor_162_48 u_ca_162_48_218(.d_in(u_ca_in_218), .d_out(u_ca_out_218));
compressor_162_48 u_ca_162_48_219(.d_in(u_ca_in_219), .d_out(u_ca_out_219));
compressor_162_48 u_ca_162_48_220(.d_in(u_ca_in_220), .d_out(u_ca_out_220));
compressor_162_48 u_ca_162_48_221(.d_in(u_ca_in_221), .d_out(u_ca_out_221));
compressor_162_48 u_ca_162_48_222(.d_in(u_ca_in_222), .d_out(u_ca_out_222));
compressor_162_48 u_ca_162_48_223(.d_in(u_ca_in_223), .d_out(u_ca_out_223));
compressor_162_48 u_ca_162_48_224(.d_in(u_ca_in_224), .d_out(u_ca_out_224));
compressor_162_48 u_ca_162_48_225(.d_in(u_ca_in_225), .d_out(u_ca_out_225));
compressor_162_48 u_ca_162_48_226(.d_in(u_ca_in_226), .d_out(u_ca_out_226));
compressor_162_48 u_ca_162_48_227(.d_in(u_ca_in_227), .d_out(u_ca_out_227));
compressor_162_48 u_ca_162_48_228(.d_in(u_ca_in_228), .d_out(u_ca_out_228));
compressor_162_48 u_ca_162_48_229(.d_in(u_ca_in_229), .d_out(u_ca_out_229));
compressor_162_48 u_ca_162_48_230(.d_in(u_ca_in_230), .d_out(u_ca_out_230));
compressor_162_48 u_ca_162_48_231(.d_in(u_ca_in_231), .d_out(u_ca_out_231));
compressor_162_48 u_ca_162_48_232(.d_in(u_ca_in_232), .d_out(u_ca_out_232));
compressor_162_48 u_ca_162_48_233(.d_in(u_ca_in_233), .d_out(u_ca_out_233));
compressor_162_48 u_ca_162_48_234(.d_in(u_ca_in_234), .d_out(u_ca_out_234));
compressor_162_48 u_ca_162_48_235(.d_in(u_ca_in_235), .d_out(u_ca_out_235));
compressor_162_48 u_ca_162_48_236(.d_in(u_ca_in_236), .d_out(u_ca_out_236));
compressor_162_48 u_ca_162_48_237(.d_in(u_ca_in_237), .d_out(u_ca_out_237));
compressor_162_48 u_ca_162_48_238(.d_in(u_ca_in_238), .d_out(u_ca_out_238));
compressor_162_48 u_ca_162_48_239(.d_in(u_ca_in_239), .d_out(u_ca_out_239));
compressor_162_48 u_ca_162_48_240(.d_in(u_ca_in_240), .d_out(u_ca_out_240));
compressor_162_48 u_ca_162_48_241(.d_in(u_ca_in_241), .d_out(u_ca_out_241));
compressor_162_48 u_ca_162_48_242(.d_in(u_ca_in_242), .d_out(u_ca_out_242));
compressor_162_48 u_ca_162_48_243(.d_in(u_ca_in_243), .d_out(u_ca_out_243));
compressor_162_48 u_ca_162_48_244(.d_in(u_ca_in_244), .d_out(u_ca_out_244));
compressor_162_48 u_ca_162_48_245(.d_in(u_ca_in_245), .d_out(u_ca_out_245));
compressor_162_48 u_ca_162_48_246(.d_in(u_ca_in_246), .d_out(u_ca_out_246));
compressor_162_48 u_ca_162_48_247(.d_in(u_ca_in_247), .d_out(u_ca_out_247));
compressor_162_48 u_ca_162_48_248(.d_in(u_ca_in_248), .d_out(u_ca_out_248));
compressor_162_48 u_ca_162_48_249(.d_in(u_ca_in_249), .d_out(u_ca_out_249));
compressor_162_48 u_ca_162_48_250(.d_in(u_ca_in_250), .d_out(u_ca_out_250));
compressor_162_48 u_ca_162_48_251(.d_in(u_ca_in_251), .d_out(u_ca_out_251));
compressor_162_48 u_ca_162_48_252(.d_in(u_ca_in_252), .d_out(u_ca_out_252));
compressor_162_48 u_ca_162_48_253(.d_in(u_ca_in_253), .d_out(u_ca_out_253));
compressor_162_48 u_ca_162_48_254(.d_in(u_ca_in_254), .d_out(u_ca_out_254));
compressor_162_48 u_ca_162_48_255(.d_in(u_ca_in_255), .d_out(u_ca_out_255));
compressor_162_48 u_ca_162_48_256(.d_in(u_ca_in_256), .d_out(u_ca_out_256));
compressor_162_48 u_ca_162_48_257(.d_in(u_ca_in_257), .d_out(u_ca_out_257));
compressor_162_48 u_ca_162_48_258(.d_in(u_ca_in_258), .d_out(u_ca_out_258));
compressor_162_48 u_ca_162_48_259(.d_in(u_ca_in_259), .d_out(u_ca_out_259));
compressor_162_48 u_ca_162_48_260(.d_in(u_ca_in_260), .d_out(u_ca_out_260));
compressor_162_48 u_ca_162_48_261(.d_in(u_ca_in_261), .d_out(u_ca_out_261));
compressor_162_48 u_ca_162_48_262(.d_in(u_ca_in_262), .d_out(u_ca_out_262));
compressor_162_48 u_ca_162_48_263(.d_in(u_ca_in_263), .d_out(u_ca_out_263));
compressor_162_48 u_ca_162_48_264(.d_in(u_ca_in_264), .d_out(u_ca_out_264));
compressor_162_48 u_ca_162_48_265(.d_in(u_ca_in_265), .d_out(u_ca_out_265));
compressor_162_48 u_ca_162_48_266(.d_in(u_ca_in_266), .d_out(u_ca_out_266));
compressor_162_48 u_ca_162_48_267(.d_in(u_ca_in_267), .d_out(u_ca_out_267));
compressor_162_48 u_ca_162_48_268(.d_in(u_ca_in_268), .d_out(u_ca_out_268));
compressor_162_48 u_ca_162_48_269(.d_in(u_ca_in_269), .d_out(u_ca_out_269));
compressor_162_48 u_ca_162_48_270(.d_in(u_ca_in_270), .d_out(u_ca_out_270));
compressor_162_48 u_ca_162_48_271(.d_in(u_ca_in_271), .d_out(u_ca_out_271));
compressor_162_48 u_ca_162_48_272(.d_in(u_ca_in_272), .d_out(u_ca_out_272));
compressor_162_48 u_ca_162_48_273(.d_in(u_ca_in_273), .d_out(u_ca_out_273));
compressor_162_48 u_ca_162_48_274(.d_in(u_ca_in_274), .d_out(u_ca_out_274));
compressor_162_48 u_ca_162_48_275(.d_in(u_ca_in_275), .d_out(u_ca_out_275));
compressor_162_48 u_ca_162_48_276(.d_in(u_ca_in_276), .d_out(u_ca_out_276));
compressor_162_48 u_ca_162_48_277(.d_in(u_ca_in_277), .d_out(u_ca_out_277));
compressor_162_48 u_ca_162_48_278(.d_in(u_ca_in_278), .d_out(u_ca_out_278));
compressor_162_48 u_ca_162_48_279(.d_in(u_ca_in_279), .d_out(u_ca_out_279));
compressor_162_48 u_ca_162_48_280(.d_in(u_ca_in_280), .d_out(u_ca_out_280));
compressor_162_48 u_ca_162_48_281(.d_in(u_ca_in_281), .d_out(u_ca_out_281));
compressor_162_48 u_ca_162_48_282(.d_in(u_ca_in_282), .d_out(u_ca_out_282));
compressor_162_48 u_ca_162_48_283(.d_in(u_ca_in_283), .d_out(u_ca_out_283));
compressor_162_48 u_ca_162_48_284(.d_in(u_ca_in_284), .d_out(u_ca_out_284));
compressor_162_48 u_ca_162_48_285(.d_in(u_ca_in_285), .d_out(u_ca_out_285));
compressor_162_48 u_ca_162_48_286(.d_in(u_ca_in_286), .d_out(u_ca_out_286));
compressor_162_48 u_ca_162_48_287(.d_in(u_ca_in_287), .d_out(u_ca_out_287));
compressor_162_48 u_ca_162_48_288(.d_in(u_ca_in_288), .d_out(u_ca_out_288));
compressor_162_48 u_ca_162_48_289(.d_in(u_ca_in_289), .d_out(u_ca_out_289));
compressor_162_48 u_ca_162_48_290(.d_in(u_ca_in_290), .d_out(u_ca_out_290));
compressor_162_48 u_ca_162_48_291(.d_in(u_ca_in_291), .d_out(u_ca_out_291));
compressor_162_48 u_ca_162_48_292(.d_in(u_ca_in_292), .d_out(u_ca_out_292));
compressor_162_48 u_ca_162_48_293(.d_in(u_ca_in_293), .d_out(u_ca_out_293));
compressor_162_48 u_ca_162_48_294(.d_in(u_ca_in_294), .d_out(u_ca_out_294));
compressor_162_48 u_ca_162_48_295(.d_in(u_ca_in_295), .d_out(u_ca_out_295));
compressor_162_48 u_ca_162_48_296(.d_in(u_ca_in_296), .d_out(u_ca_out_296));
compressor_162_48 u_ca_162_48_297(.d_in(u_ca_in_297), .d_out(u_ca_out_297));
compressor_162_48 u_ca_162_48_298(.d_in(u_ca_in_298), .d_out(u_ca_out_298));
compressor_162_48 u_ca_162_48_299(.d_in(u_ca_in_299), .d_out(u_ca_out_299));
compressor_162_48 u_ca_162_48_300(.d_in(u_ca_in_300), .d_out(u_ca_out_300));
compressor_162_48 u_ca_162_48_301(.d_in(u_ca_in_301), .d_out(u_ca_out_301));
compressor_162_48 u_ca_162_48_302(.d_in(u_ca_in_302), .d_out(u_ca_out_302));
compressor_162_48 u_ca_162_48_303(.d_in(u_ca_in_303), .d_out(u_ca_out_303));
compressor_162_48 u_ca_162_48_304(.d_in(u_ca_in_304), .d_out(u_ca_out_304));
compressor_162_48 u_ca_162_48_305(.d_in(u_ca_in_305), .d_out(u_ca_out_305));
compressor_162_48 u_ca_162_48_306(.d_in(u_ca_in_306), .d_out(u_ca_out_306));
compressor_162_48 u_ca_162_48_307(.d_in(u_ca_in_307), .d_out(u_ca_out_307));
compressor_162_48 u_ca_162_48_308(.d_in(u_ca_in_308), .d_out(u_ca_out_308));
compressor_162_48 u_ca_162_48_309(.d_in(u_ca_in_309), .d_out(u_ca_out_309));
compressor_162_48 u_ca_162_48_310(.d_in(u_ca_in_310), .d_out(u_ca_out_310));
compressor_162_48 u_ca_162_48_311(.d_in(u_ca_in_311), .d_out(u_ca_out_311));
compressor_162_48 u_ca_162_48_312(.d_in(u_ca_in_312), .d_out(u_ca_out_312));
compressor_162_48 u_ca_162_48_313(.d_in(u_ca_in_313), .d_out(u_ca_out_313));
compressor_162_48 u_ca_162_48_314(.d_in(u_ca_in_314), .d_out(u_ca_out_314));
compressor_162_48 u_ca_162_48_315(.d_in(u_ca_in_315), .d_out(u_ca_out_315));
compressor_162_48 u_ca_162_48_316(.d_in(u_ca_in_316), .d_out(u_ca_out_316));
compressor_162_48 u_ca_162_48_317(.d_in(u_ca_in_317), .d_out(u_ca_out_317));
compressor_162_48 u_ca_162_48_318(.d_in(u_ca_in_318), .d_out(u_ca_out_318));
compressor_162_48 u_ca_162_48_319(.d_in(u_ca_in_319), .d_out(u_ca_out_319));
compressor_162_48 u_ca_162_48_320(.d_in(u_ca_in_320), .d_out(u_ca_out_320));
compressor_162_48 u_ca_162_48_321(.d_in(u_ca_in_321), .d_out(u_ca_out_321));
compressor_162_48 u_ca_162_48_322(.d_in(u_ca_in_322), .d_out(u_ca_out_322));
compressor_162_48 u_ca_162_48_323(.d_in(u_ca_in_323), .d_out(u_ca_out_323));
compressor_162_48 u_ca_162_48_324(.d_in(u_ca_in_324), .d_out(u_ca_out_324));
compressor_162_48 u_ca_162_48_325(.d_in(u_ca_in_325), .d_out(u_ca_out_325));
compressor_162_48 u_ca_162_48_326(.d_in(u_ca_in_326), .d_out(u_ca_out_326));
compressor_162_48 u_ca_162_48_327(.d_in(u_ca_in_327), .d_out(u_ca_out_327));
compressor_162_48 u_ca_162_48_328(.d_in(u_ca_in_328), .d_out(u_ca_out_328));
compressor_162_48 u_ca_162_48_329(.d_in(u_ca_in_329), .d_out(u_ca_out_329));
compressor_162_48 u_ca_162_48_330(.d_in(u_ca_in_330), .d_out(u_ca_out_330));
compressor_162_48 u_ca_162_48_331(.d_in(u_ca_in_331), .d_out(u_ca_out_331));
compressor_162_48 u_ca_162_48_332(.d_in(u_ca_in_332), .d_out(u_ca_out_332));
compressor_162_48 u_ca_162_48_333(.d_in(u_ca_in_333), .d_out(u_ca_out_333));
compressor_162_48 u_ca_162_48_334(.d_in(u_ca_in_334), .d_out(u_ca_out_334));
compressor_162_48 u_ca_162_48_335(.d_in(u_ca_in_335), .d_out(u_ca_out_335));
compressor_162_48 u_ca_162_48_336(.d_in(u_ca_in_336), .d_out(u_ca_out_336));
compressor_162_48 u_ca_162_48_337(.d_in(u_ca_in_337), .d_out(u_ca_out_337));
compressor_162_48 u_ca_162_48_338(.d_in(u_ca_in_338), .d_out(u_ca_out_338));
compressor_162_48 u_ca_162_48_339(.d_in(u_ca_in_339), .d_out(u_ca_out_339));
compressor_162_48 u_ca_162_48_340(.d_in(u_ca_in_340), .d_out(u_ca_out_340));
compressor_162_48 u_ca_162_48_341(.d_in(u_ca_in_341), .d_out(u_ca_out_341));
compressor_162_48 u_ca_162_48_342(.d_in(u_ca_in_342), .d_out(u_ca_out_342));
compressor_162_48 u_ca_162_48_343(.d_in(u_ca_in_343), .d_out(u_ca_out_343));
compressor_162_48 u_ca_162_48_344(.d_in(u_ca_in_344), .d_out(u_ca_out_344));
compressor_162_48 u_ca_162_48_345(.d_in(u_ca_in_345), .d_out(u_ca_out_345));
compressor_162_48 u_ca_162_48_346(.d_in(u_ca_in_346), .d_out(u_ca_out_346));
compressor_162_48 u_ca_162_48_347(.d_in(u_ca_in_347), .d_out(u_ca_out_347));
compressor_162_48 u_ca_162_48_348(.d_in(u_ca_in_348), .d_out(u_ca_out_348));
compressor_162_48 u_ca_162_48_349(.d_in(u_ca_in_349), .d_out(u_ca_out_349));
compressor_162_48 u_ca_162_48_350(.d_in(u_ca_in_350), .d_out(u_ca_out_350));
compressor_162_48 u_ca_162_48_351(.d_in(u_ca_in_351), .d_out(u_ca_out_351));
compressor_162_48 u_ca_162_48_352(.d_in(u_ca_in_352), .d_out(u_ca_out_352));
compressor_162_48 u_ca_162_48_353(.d_in(u_ca_in_353), .d_out(u_ca_out_353));
compressor_162_48 u_ca_162_48_354(.d_in(u_ca_in_354), .d_out(u_ca_out_354));
compressor_162_48 u_ca_162_48_355(.d_in(u_ca_in_355), .d_out(u_ca_out_355));
compressor_162_48 u_ca_162_48_356(.d_in(u_ca_in_356), .d_out(u_ca_out_356));
compressor_162_48 u_ca_162_48_357(.d_in(u_ca_in_357), .d_out(u_ca_out_357));
compressor_162_48 u_ca_162_48_358(.d_in(u_ca_in_358), .d_out(u_ca_out_358));
compressor_162_48 u_ca_162_48_359(.d_in(u_ca_in_359), .d_out(u_ca_out_359));
compressor_162_48 u_ca_162_48_360(.d_in(u_ca_in_360), .d_out(u_ca_out_360));
compressor_162_48 u_ca_162_48_361(.d_in(u_ca_in_361), .d_out(u_ca_out_361));
compressor_162_48 u_ca_162_48_362(.d_in(u_ca_in_362), .d_out(u_ca_out_362));
compressor_162_48 u_ca_162_48_363(.d_in(u_ca_in_363), .d_out(u_ca_out_363));
compressor_162_48 u_ca_162_48_364(.d_in(u_ca_in_364), .d_out(u_ca_out_364));
compressor_162_48 u_ca_162_48_365(.d_in(u_ca_in_365), .d_out(u_ca_out_365));
compressor_162_48 u_ca_162_48_366(.d_in(u_ca_in_366), .d_out(u_ca_out_366));
compressor_162_48 u_ca_162_48_367(.d_in(u_ca_in_367), .d_out(u_ca_out_367));
compressor_162_48 u_ca_162_48_368(.d_in(u_ca_in_368), .d_out(u_ca_out_368));
compressor_162_48 u_ca_162_48_369(.d_in(u_ca_in_369), .d_out(u_ca_out_369));
compressor_162_48 u_ca_162_48_370(.d_in(u_ca_in_370), .d_out(u_ca_out_370));
compressor_162_48 u_ca_162_48_371(.d_in(u_ca_in_371), .d_out(u_ca_out_371));
compressor_162_48 u_ca_162_48_372(.d_in(u_ca_in_372), .d_out(u_ca_out_372));
compressor_162_48 u_ca_162_48_373(.d_in(u_ca_in_373), .d_out(u_ca_out_373));
compressor_162_48 u_ca_162_48_374(.d_in(u_ca_in_374), .d_out(u_ca_out_374));
compressor_162_48 u_ca_162_48_375(.d_in(u_ca_in_375), .d_out(u_ca_out_375));
compressor_162_48 u_ca_162_48_376(.d_in(u_ca_in_376), .d_out(u_ca_out_376));
compressor_162_48 u_ca_162_48_377(.d_in(u_ca_in_377), .d_out(u_ca_out_377));
compressor_162_48 u_ca_162_48_378(.d_in(u_ca_in_378), .d_out(u_ca_out_378));
compressor_162_48 u_ca_162_48_379(.d_in(u_ca_in_379), .d_out(u_ca_out_379));
compressor_162_48 u_ca_162_48_380(.d_in(u_ca_in_380), .d_out(u_ca_out_380));
compressor_162_48 u_ca_162_48_381(.d_in(u_ca_in_381), .d_out(u_ca_out_381));
compressor_162_48 u_ca_162_48_382(.d_in(u_ca_in_382), .d_out(u_ca_out_382));
compressor_162_48 u_ca_162_48_383(.d_in(u_ca_in_383), .d_out(u_ca_out_383));
compressor_162_48 u_ca_162_48_384(.d_in(u_ca_in_384), .d_out(u_ca_out_384));
compressor_162_48 u_ca_162_48_385(.d_in(u_ca_in_385), .d_out(u_ca_out_385));
compressor_162_48 u_ca_162_48_386(.d_in(u_ca_in_386), .d_out(u_ca_out_386));
compressor_162_48 u_ca_162_48_387(.d_in(u_ca_in_387), .d_out(u_ca_out_387));
compressor_162_48 u_ca_162_48_388(.d_in(u_ca_in_388), .d_out(u_ca_out_388));
compressor_162_48 u_ca_162_48_389(.d_in(u_ca_in_389), .d_out(u_ca_out_389));
compressor_162_48 u_ca_162_48_390(.d_in(u_ca_in_390), .d_out(u_ca_out_390));
compressor_162_48 u_ca_162_48_391(.d_in(u_ca_in_391), .d_out(u_ca_out_391));
compressor_162_48 u_ca_162_48_392(.d_in(u_ca_in_392), .d_out(u_ca_out_392));
compressor_162_48 u_ca_162_48_393(.d_in(u_ca_in_393), .d_out(u_ca_out_393));
compressor_162_48 u_ca_162_48_394(.d_in(u_ca_in_394), .d_out(u_ca_out_394));
compressor_162_48 u_ca_162_48_395(.d_in(u_ca_in_395), .d_out(u_ca_out_395));
compressor_162_48 u_ca_162_48_396(.d_in(u_ca_in_396), .d_out(u_ca_out_396));
compressor_162_48 u_ca_162_48_397(.d_in(u_ca_in_397), .d_out(u_ca_out_397));
compressor_162_48 u_ca_162_48_398(.d_in(u_ca_in_398), .d_out(u_ca_out_398));
compressor_162_48 u_ca_162_48_399(.d_in(u_ca_in_399), .d_out(u_ca_out_399));
compressor_162_48 u_ca_162_48_400(.d_in(u_ca_in_400), .d_out(u_ca_out_400));
compressor_162_48 u_ca_162_48_401(.d_in(u_ca_in_401), .d_out(u_ca_out_401));
compressor_162_48 u_ca_162_48_402(.d_in(u_ca_in_402), .d_out(u_ca_out_402));
compressor_162_48 u_ca_162_48_403(.d_in(u_ca_in_403), .d_out(u_ca_out_403));
compressor_162_48 u_ca_162_48_404(.d_in(u_ca_in_404), .d_out(u_ca_out_404));
compressor_162_48 u_ca_162_48_405(.d_in(u_ca_in_405), .d_out(u_ca_out_405));
compressor_162_48 u_ca_162_48_406(.d_in(u_ca_in_406), .d_out(u_ca_out_406));
compressor_162_48 u_ca_162_48_407(.d_in(u_ca_in_407), .d_out(u_ca_out_407));
compressor_162_48 u_ca_162_48_408(.d_in(u_ca_in_408), .d_out(u_ca_out_408));
compressor_162_48 u_ca_162_48_409(.d_in(u_ca_in_409), .d_out(u_ca_out_409));
compressor_162_48 u_ca_162_48_410(.d_in(u_ca_in_410), .d_out(u_ca_out_410));
compressor_162_48 u_ca_162_48_411(.d_in(u_ca_in_411), .d_out(u_ca_out_411));
compressor_162_48 u_ca_162_48_412(.d_in(u_ca_in_412), .d_out(u_ca_out_412));
compressor_162_48 u_ca_162_48_413(.d_in(u_ca_in_413), .d_out(u_ca_out_413));
compressor_162_48 u_ca_162_48_414(.d_in(u_ca_in_414), .d_out(u_ca_out_414));
compressor_162_48 u_ca_162_48_415(.d_in(u_ca_in_415), .d_out(u_ca_out_415));
compressor_162_48 u_ca_162_48_416(.d_in(u_ca_in_416), .d_out(u_ca_out_416));
compressor_162_48 u_ca_162_48_417(.d_in(u_ca_in_417), .d_out(u_ca_out_417));
compressor_162_48 u_ca_162_48_418(.d_in(u_ca_in_418), .d_out(u_ca_out_418));
compressor_162_48 u_ca_162_48_419(.d_in(u_ca_in_419), .d_out(u_ca_out_419));
compressor_162_48 u_ca_162_48_420(.d_in(u_ca_in_420), .d_out(u_ca_out_420));
compressor_162_48 u_ca_162_48_421(.d_in(u_ca_in_421), .d_out(u_ca_out_421));
compressor_162_48 u_ca_162_48_422(.d_in(u_ca_in_422), .d_out(u_ca_out_422));
compressor_162_48 u_ca_162_48_423(.d_in(u_ca_in_423), .d_out(u_ca_out_423));
compressor_162_48 u_ca_162_48_424(.d_in(u_ca_in_424), .d_out(u_ca_out_424));
compressor_162_48 u_ca_162_48_425(.d_in(u_ca_in_425), .d_out(u_ca_out_425));
compressor_162_48 u_ca_162_48_426(.d_in(u_ca_in_426), .d_out(u_ca_out_426));
compressor_162_48 u_ca_162_48_427(.d_in(u_ca_in_427), .d_out(u_ca_out_427));
compressor_162_48 u_ca_162_48_428(.d_in(u_ca_in_428), .d_out(u_ca_out_428));
compressor_162_48 u_ca_162_48_429(.d_in(u_ca_in_429), .d_out(u_ca_out_429));
compressor_162_48 u_ca_162_48_430(.d_in(u_ca_in_430), .d_out(u_ca_out_430));
compressor_162_48 u_ca_162_48_431(.d_in(u_ca_in_431), .d_out(u_ca_out_431));
compressor_162_48 u_ca_162_48_432(.d_in(u_ca_in_432), .d_out(u_ca_out_432));
compressor_162_48 u_ca_162_48_433(.d_in(u_ca_in_433), .d_out(u_ca_out_433));
compressor_162_48 u_ca_162_48_434(.d_in(u_ca_in_434), .d_out(u_ca_out_434));
compressor_162_48 u_ca_162_48_435(.d_in(u_ca_in_435), .d_out(u_ca_out_435));
compressor_162_48 u_ca_162_48_436(.d_in(u_ca_in_436), .d_out(u_ca_out_436));
compressor_162_48 u_ca_162_48_437(.d_in(u_ca_in_437), .d_out(u_ca_out_437));
compressor_162_48 u_ca_162_48_438(.d_in(u_ca_in_438), .d_out(u_ca_out_438));
compressor_162_48 u_ca_162_48_439(.d_in(u_ca_in_439), .d_out(u_ca_out_439));
compressor_162_48 u_ca_162_48_440(.d_in(u_ca_in_440), .d_out(u_ca_out_440));
compressor_162_48 u_ca_162_48_441(.d_in(u_ca_in_441), .d_out(u_ca_out_441));
compressor_162_48 u_ca_162_48_442(.d_in(u_ca_in_442), .d_out(u_ca_out_442));
compressor_162_48 u_ca_162_48_443(.d_in(u_ca_in_443), .d_out(u_ca_out_443));
compressor_162_48 u_ca_162_48_444(.d_in(u_ca_in_444), .d_out(u_ca_out_444));
compressor_162_48 u_ca_162_48_445(.d_in(u_ca_in_445), .d_out(u_ca_out_445));
compressor_162_48 u_ca_162_48_446(.d_in(u_ca_in_446), .d_out(u_ca_out_446));
compressor_162_48 u_ca_162_48_447(.d_in(u_ca_in_447), .d_out(u_ca_out_447));
compressor_162_48 u_ca_162_48_448(.d_in(u_ca_in_448), .d_out(u_ca_out_448));
compressor_162_48 u_ca_162_48_449(.d_in(u_ca_in_449), .d_out(u_ca_out_449));
compressor_162_48 u_ca_162_48_450(.d_in(u_ca_in_450), .d_out(u_ca_out_450));
compressor_162_48 u_ca_162_48_451(.d_in(u_ca_in_451), .d_out(u_ca_out_451));
compressor_162_48 u_ca_162_48_452(.d_in(u_ca_in_452), .d_out(u_ca_out_452));
compressor_162_48 u_ca_162_48_453(.d_in(u_ca_in_453), .d_out(u_ca_out_453));
compressor_162_48 u_ca_162_48_454(.d_in(u_ca_in_454), .d_out(u_ca_out_454));
compressor_162_48 u_ca_162_48_455(.d_in(u_ca_in_455), .d_out(u_ca_out_455));
compressor_162_48 u_ca_162_48_456(.d_in(u_ca_in_456), .d_out(u_ca_out_456));
compressor_162_48 u_ca_162_48_457(.d_in(u_ca_in_457), .d_out(u_ca_out_457));
compressor_162_48 u_ca_162_48_458(.d_in(u_ca_in_458), .d_out(u_ca_out_458));
compressor_162_48 u_ca_162_48_459(.d_in(u_ca_in_459), .d_out(u_ca_out_459));
compressor_162_48 u_ca_162_48_460(.d_in(u_ca_in_460), .d_out(u_ca_out_460));
compressor_162_48 u_ca_162_48_461(.d_in(u_ca_in_461), .d_out(u_ca_out_461));
compressor_162_48 u_ca_162_48_462(.d_in(u_ca_in_462), .d_out(u_ca_out_462));
compressor_162_48 u_ca_162_48_463(.d_in(u_ca_in_463), .d_out(u_ca_out_463));
compressor_162_48 u_ca_162_48_464(.d_in(u_ca_in_464), .d_out(u_ca_out_464));
compressor_162_48 u_ca_162_48_465(.d_in(u_ca_in_465), .d_out(u_ca_out_465));
compressor_162_48 u_ca_162_48_466(.d_in(u_ca_in_466), .d_out(u_ca_out_466));
compressor_162_48 u_ca_162_48_467(.d_in(u_ca_in_467), .d_out(u_ca_out_467));
compressor_162_48 u_ca_162_48_468(.d_in(u_ca_in_468), .d_out(u_ca_out_468));
compressor_162_48 u_ca_162_48_469(.d_in(u_ca_in_469), .d_out(u_ca_out_469));
compressor_162_48 u_ca_162_48_470(.d_in(u_ca_in_470), .d_out(u_ca_out_470));
compressor_162_48 u_ca_162_48_471(.d_in(u_ca_in_471), .d_out(u_ca_out_471));
compressor_162_48 u_ca_162_48_472(.d_in(u_ca_in_472), .d_out(u_ca_out_472));
compressor_162_48 u_ca_162_48_473(.d_in(u_ca_in_473), .d_out(u_ca_out_473));
compressor_162_48 u_ca_162_48_474(.d_in(u_ca_in_474), .d_out(u_ca_out_474));
compressor_162_48 u_ca_162_48_475(.d_in(u_ca_in_475), .d_out(u_ca_out_475));
compressor_162_48 u_ca_162_48_476(.d_in(u_ca_in_476), .d_out(u_ca_out_476));
compressor_162_48 u_ca_162_48_477(.d_in(u_ca_in_477), .d_out(u_ca_out_477));
compressor_162_48 u_ca_162_48_478(.d_in(u_ca_in_478), .d_out(u_ca_out_478));
compressor_162_48 u_ca_162_48_479(.d_in(u_ca_in_479), .d_out(u_ca_out_479));
compressor_162_48 u_ca_162_48_480(.d_in(u_ca_in_480), .d_out(u_ca_out_480));
compressor_162_48 u_ca_162_48_481(.d_in(u_ca_in_481), .d_out(u_ca_out_481));
compressor_162_48 u_ca_162_48_482(.d_in(u_ca_in_482), .d_out(u_ca_out_482));
compressor_162_48 u_ca_162_48_483(.d_in(u_ca_in_483), .d_out(u_ca_out_483));
compressor_162_48 u_ca_162_48_484(.d_in(u_ca_in_484), .d_out(u_ca_out_484));
compressor_162_48 u_ca_162_48_485(.d_in(u_ca_in_485), .d_out(u_ca_out_485));
compressor_162_48 u_ca_162_48_486(.d_in(u_ca_in_486), .d_out(u_ca_out_486));
compressor_162_48 u_ca_162_48_487(.d_in(u_ca_in_487), .d_out(u_ca_out_487));
compressor_162_48 u_ca_162_48_488(.d_in(u_ca_in_488), .d_out(u_ca_out_488));
compressor_162_48 u_ca_162_48_489(.d_in(u_ca_in_489), .d_out(u_ca_out_489));
compressor_162_48 u_ca_162_48_490(.d_in(u_ca_in_490), .d_out(u_ca_out_490));
compressor_162_48 u_ca_162_48_491(.d_in(u_ca_in_491), .d_out(u_ca_out_491));
compressor_162_48 u_ca_162_48_492(.d_in(u_ca_in_492), .d_out(u_ca_out_492));
compressor_162_48 u_ca_162_48_493(.d_in(u_ca_in_493), .d_out(u_ca_out_493));
compressor_162_48 u_ca_162_48_494(.d_in(u_ca_in_494), .d_out(u_ca_out_494));
compressor_162_48 u_ca_162_48_495(.d_in(u_ca_in_495), .d_out(u_ca_out_495));
compressor_162_48 u_ca_162_48_496(.d_in(u_ca_in_496), .d_out(u_ca_out_496));
compressor_162_48 u_ca_162_48_497(.d_in(u_ca_in_497), .d_out(u_ca_out_497));
compressor_162_48 u_ca_162_48_498(.d_in(u_ca_in_498), .d_out(u_ca_out_498));
compressor_162_48 u_ca_162_48_499(.d_in(u_ca_in_499), .d_out(u_ca_out_499));
compressor_162_48 u_ca_162_48_500(.d_in(u_ca_in_500), .d_out(u_ca_out_500));
compressor_162_48 u_ca_162_48_501(.d_in(u_ca_in_501), .d_out(u_ca_out_501));
compressor_162_48 u_ca_162_48_502(.d_in(u_ca_in_502), .d_out(u_ca_out_502));
compressor_162_48 u_ca_162_48_503(.d_in(u_ca_in_503), .d_out(u_ca_out_503));
compressor_162_48 u_ca_162_48_504(.d_in(u_ca_in_504), .d_out(u_ca_out_504));
compressor_162_48 u_ca_162_48_505(.d_in(u_ca_in_505), .d_out(u_ca_out_505));
compressor_162_48 u_ca_162_48_506(.d_in(u_ca_in_506), .d_out(u_ca_out_506));
compressor_162_48 u_ca_162_48_507(.d_in(u_ca_in_507), .d_out(u_ca_out_507));
compressor_162_48 u_ca_162_48_508(.d_in(u_ca_in_508), .d_out(u_ca_out_508));
compressor_162_48 u_ca_162_48_509(.d_in(u_ca_in_509), .d_out(u_ca_out_509));
compressor_162_48 u_ca_162_48_510(.d_in(u_ca_in_510), .d_out(u_ca_out_510));
compressor_162_48 u_ca_162_48_511(.d_in(u_ca_in_511), .d_out(u_ca_out_511));
compressor_162_48 u_ca_162_48_512(.d_in(u_ca_in_512), .d_out(u_ca_out_512));
compressor_162_48 u_ca_162_48_513(.d_in(u_ca_in_513), .d_out(u_ca_out_513));
compressor_162_48 u_ca_162_48_514(.d_in(u_ca_in_514), .d_out(u_ca_out_514));
compressor_162_48 u_ca_162_48_515(.d_in(u_ca_in_515), .d_out(u_ca_out_515));
compressor_162_48 u_ca_162_48_516(.d_in(u_ca_in_516), .d_out(u_ca_out_516));
compressor_162_48 u_ca_162_48_517(.d_in(u_ca_in_517), .d_out(u_ca_out_517));
compressor_162_48 u_ca_162_48_518(.d_in(u_ca_in_518), .d_out(u_ca_out_518));
compressor_162_48 u_ca_162_48_519(.d_in(u_ca_in_519), .d_out(u_ca_out_519));
compressor_162_48 u_ca_162_48_520(.d_in(u_ca_in_520), .d_out(u_ca_out_520));
compressor_162_48 u_ca_162_48_521(.d_in(u_ca_in_521), .d_out(u_ca_out_521));
compressor_162_48 u_ca_162_48_522(.d_in(u_ca_in_522), .d_out(u_ca_out_522));
compressor_162_48 u_ca_162_48_523(.d_in(u_ca_in_523), .d_out(u_ca_out_523));
compressor_162_48 u_ca_162_48_524(.d_in(u_ca_in_524), .d_out(u_ca_out_524));
compressor_162_48 u_ca_162_48_525(.d_in(u_ca_in_525), .d_out(u_ca_out_525));
compressor_162_48 u_ca_162_48_526(.d_in(u_ca_in_526), .d_out(u_ca_out_526));
compressor_162_48 u_ca_162_48_527(.d_in(u_ca_in_527), .d_out(u_ca_out_527));
compressor_162_48 u_ca_162_48_528(.d_in(u_ca_in_528), .d_out(u_ca_out_528));
compressor_162_48 u_ca_162_48_529(.d_in(u_ca_in_529), .d_out(u_ca_out_529));
compressor_162_48 u_ca_162_48_530(.d_in(u_ca_in_530), .d_out(u_ca_out_530));
compressor_162_48 u_ca_162_48_531(.d_in(u_ca_in_531), .d_out(u_ca_out_531));
compressor_162_48 u_ca_162_48_532(.d_in(u_ca_in_532), .d_out(u_ca_out_532));
compressor_162_48 u_ca_162_48_533(.d_in(u_ca_in_533), .d_out(u_ca_out_533));
compressor_162_48 u_ca_162_48_534(.d_in(u_ca_in_534), .d_out(u_ca_out_534));
compressor_162_48 u_ca_162_48_535(.d_in(u_ca_in_535), .d_out(u_ca_out_535));
compressor_162_48 u_ca_162_48_536(.d_in(u_ca_in_536), .d_out(u_ca_out_536));
compressor_162_48 u_ca_162_48_537(.d_in(u_ca_in_537), .d_out(u_ca_out_537));
compressor_162_48 u_ca_162_48_538(.d_in(u_ca_in_538), .d_out(u_ca_out_538));
compressor_162_48 u_ca_162_48_539(.d_in(u_ca_in_539), .d_out(u_ca_out_539));
compressor_162_48 u_ca_162_48_540(.d_in(u_ca_in_540), .d_out(u_ca_out_540));
compressor_162_48 u_ca_162_48_541(.d_in(u_ca_in_541), .d_out(u_ca_out_541));
compressor_162_48 u_ca_162_48_542(.d_in(u_ca_in_542), .d_out(u_ca_out_542));
compressor_162_48 u_ca_162_48_543(.d_in(u_ca_in_543), .d_out(u_ca_out_543));
compressor_162_48 u_ca_162_48_544(.d_in(u_ca_in_544), .d_out(u_ca_out_544));
compressor_162_48 u_ca_162_48_545(.d_in(u_ca_in_545), .d_out(u_ca_out_545));
compressor_162_48 u_ca_162_48_546(.d_in(u_ca_in_546), .d_out(u_ca_out_546));
compressor_162_48 u_ca_162_48_547(.d_in(u_ca_in_547), .d_out(u_ca_out_547));
compressor_162_48 u_ca_162_48_548(.d_in(u_ca_in_548), .d_out(u_ca_out_548));
compressor_162_48 u_ca_162_48_549(.d_in(u_ca_in_549), .d_out(u_ca_out_549));
compressor_162_48 u_ca_162_48_550(.d_in(u_ca_in_550), .d_out(u_ca_out_550));
compressor_162_48 u_ca_162_48_551(.d_in(u_ca_in_551), .d_out(u_ca_out_551));
compressor_162_48 u_ca_162_48_552(.d_in(u_ca_in_552), .d_out(u_ca_out_552));
compressor_162_48 u_ca_162_48_553(.d_in(u_ca_in_553), .d_out(u_ca_out_553));
compressor_162_48 u_ca_162_48_554(.d_in(u_ca_in_554), .d_out(u_ca_out_554));
compressor_162_48 u_ca_162_48_555(.d_in(u_ca_in_555), .d_out(u_ca_out_555));
compressor_162_48 u_ca_162_48_556(.d_in(u_ca_in_556), .d_out(u_ca_out_556));
compressor_162_48 u_ca_162_48_557(.d_in(u_ca_in_557), .d_out(u_ca_out_557));
compressor_162_48 u_ca_162_48_558(.d_in(u_ca_in_558), .d_out(u_ca_out_558));
compressor_162_48 u_ca_162_48_559(.d_in(u_ca_in_559), .d_out(u_ca_out_559));
compressor_162_48 u_ca_162_48_560(.d_in(u_ca_in_560), .d_out(u_ca_out_560));
compressor_162_48 u_ca_162_48_561(.d_in(u_ca_in_561), .d_out(u_ca_out_561));
compressor_162_48 u_ca_162_48_562(.d_in(u_ca_in_562), .d_out(u_ca_out_562));
compressor_162_48 u_ca_162_48_563(.d_in(u_ca_in_563), .d_out(u_ca_out_563));
compressor_162_48 u_ca_162_48_564(.d_in(u_ca_in_564), .d_out(u_ca_out_564));
compressor_162_48 u_ca_162_48_565(.d_in(u_ca_in_565), .d_out(u_ca_out_565));
compressor_162_48 u_ca_162_48_566(.d_in(u_ca_in_566), .d_out(u_ca_out_566));
compressor_162_48 u_ca_162_48_567(.d_in(u_ca_in_567), .d_out(u_ca_out_567));
compressor_162_48 u_ca_162_48_568(.d_in(u_ca_in_568), .d_out(u_ca_out_568));
compressor_162_48 u_ca_162_48_569(.d_in(u_ca_in_569), .d_out(u_ca_out_569));
compressor_162_48 u_ca_162_48_570(.d_in(u_ca_in_570), .d_out(u_ca_out_570));
compressor_162_48 u_ca_162_48_571(.d_in(u_ca_in_571), .d_out(u_ca_out_571));
compressor_162_48 u_ca_162_48_572(.d_in(u_ca_in_572), .d_out(u_ca_out_572));
compressor_162_48 u_ca_162_48_573(.d_in(u_ca_in_573), .d_out(u_ca_out_573));
compressor_162_48 u_ca_162_48_574(.d_in(u_ca_in_574), .d_out(u_ca_out_574));
compressor_162_48 u_ca_162_48_575(.d_in(u_ca_in_575), .d_out(u_ca_out_575));
compressor_162_48 u_ca_162_48_576(.d_in(u_ca_in_576), .d_out(u_ca_out_576));
compressor_162_48 u_ca_162_48_577(.d_in(u_ca_in_577), .d_out(u_ca_out_577));
compressor_162_48 u_ca_162_48_578(.d_in(u_ca_in_578), .d_out(u_ca_out_578));
compressor_162_48 u_ca_162_48_579(.d_in(u_ca_in_579), .d_out(u_ca_out_579));
compressor_162_48 u_ca_162_48_580(.d_in(u_ca_in_580), .d_out(u_ca_out_580));
compressor_162_48 u_ca_162_48_581(.d_in(u_ca_in_581), .d_out(u_ca_out_581));
compressor_162_48 u_ca_162_48_582(.d_in(u_ca_in_582), .d_out(u_ca_out_582));
compressor_162_48 u_ca_162_48_583(.d_in(u_ca_in_583), .d_out(u_ca_out_583));
compressor_162_48 u_ca_162_48_584(.d_in(u_ca_in_584), .d_out(u_ca_out_584));
compressor_162_48 u_ca_162_48_585(.d_in(u_ca_in_585), .d_out(u_ca_out_585));
compressor_162_48 u_ca_162_48_586(.d_in(u_ca_in_586), .d_out(u_ca_out_586));
compressor_162_48 u_ca_162_48_587(.d_in(u_ca_in_587), .d_out(u_ca_out_587));
compressor_162_48 u_ca_162_48_588(.d_in(u_ca_in_588), .d_out(u_ca_out_588));
compressor_162_48 u_ca_162_48_589(.d_in(u_ca_in_589), .d_out(u_ca_out_589));
compressor_162_48 u_ca_162_48_590(.d_in(u_ca_in_590), .d_out(u_ca_out_590));
compressor_162_48 u_ca_162_48_591(.d_in(u_ca_in_591), .d_out(u_ca_out_591));
compressor_162_48 u_ca_162_48_592(.d_in(u_ca_in_592), .d_out(u_ca_out_592));
compressor_162_48 u_ca_162_48_593(.d_in(u_ca_in_593), .d_out(u_ca_out_593));
compressor_162_48 u_ca_162_48_594(.d_in(u_ca_in_594), .d_out(u_ca_out_594));
compressor_162_48 u_ca_162_48_595(.d_in(u_ca_in_595), .d_out(u_ca_out_595));
compressor_162_48 u_ca_162_48_596(.d_in(u_ca_in_596), .d_out(u_ca_out_596));
compressor_162_48 u_ca_162_48_597(.d_in(u_ca_in_597), .d_out(u_ca_out_597));
compressor_162_48 u_ca_162_48_598(.d_in(u_ca_in_598), .d_out(u_ca_out_598));
compressor_162_48 u_ca_162_48_599(.d_in(u_ca_in_599), .d_out(u_ca_out_599));
compressor_162_48 u_ca_162_48_600(.d_in(u_ca_in_600), .d_out(u_ca_out_600));
compressor_162_48 u_ca_162_48_601(.d_in(u_ca_in_601), .d_out(u_ca_out_601));
compressor_162_48 u_ca_162_48_602(.d_in(u_ca_in_602), .d_out(u_ca_out_602));
compressor_162_48 u_ca_162_48_603(.d_in(u_ca_in_603), .d_out(u_ca_out_603));
compressor_162_48 u_ca_162_48_604(.d_in(u_ca_in_604), .d_out(u_ca_out_604));
compressor_162_48 u_ca_162_48_605(.d_in(u_ca_in_605), .d_out(u_ca_out_605));
compressor_162_48 u_ca_162_48_606(.d_in(u_ca_in_606), .d_out(u_ca_out_606));
compressor_162_48 u_ca_162_48_607(.d_in(u_ca_in_607), .d_out(u_ca_out_607));
compressor_162_48 u_ca_162_48_608(.d_in(u_ca_in_608), .d_out(u_ca_out_608));
compressor_162_48 u_ca_162_48_609(.d_in(u_ca_in_609), .d_out(u_ca_out_609));
compressor_162_48 u_ca_162_48_610(.d_in(u_ca_in_610), .d_out(u_ca_out_610));
compressor_162_48 u_ca_162_48_611(.d_in(u_ca_in_611), .d_out(u_ca_out_611));
compressor_162_48 u_ca_162_48_612(.d_in(u_ca_in_612), .d_out(u_ca_out_612));
compressor_162_48 u_ca_162_48_613(.d_in(u_ca_in_613), .d_out(u_ca_out_613));
compressor_162_48 u_ca_162_48_614(.d_in(u_ca_in_614), .d_out(u_ca_out_614));
compressor_162_48 u_ca_162_48_615(.d_in(u_ca_in_615), .d_out(u_ca_out_615));
compressor_162_48 u_ca_162_48_616(.d_in(u_ca_in_616), .d_out(u_ca_out_616));
compressor_162_48 u_ca_162_48_617(.d_in(u_ca_in_617), .d_out(u_ca_out_617));
compressor_162_48 u_ca_162_48_618(.d_in(u_ca_in_618), .d_out(u_ca_out_618));
compressor_162_48 u_ca_162_48_619(.d_in(u_ca_in_619), .d_out(u_ca_out_619));
compressor_162_48 u_ca_162_48_620(.d_in(u_ca_in_620), .d_out(u_ca_out_620));
compressor_162_48 u_ca_162_48_621(.d_in(u_ca_in_621), .d_out(u_ca_out_621));
compressor_162_48 u_ca_162_48_622(.d_in(u_ca_in_622), .d_out(u_ca_out_622));
compressor_162_48 u_ca_162_48_623(.d_in(u_ca_in_623), .d_out(u_ca_out_623));
compressor_162_48 u_ca_162_48_624(.d_in(u_ca_in_624), .d_out(u_ca_out_624));
compressor_162_48 u_ca_162_48_625(.d_in(u_ca_in_625), .d_out(u_ca_out_625));
compressor_162_48 u_ca_162_48_626(.d_in(u_ca_in_626), .d_out(u_ca_out_626));
compressor_162_48 u_ca_162_48_627(.d_in(u_ca_in_627), .d_out(u_ca_out_627));
compressor_162_48 u_ca_162_48_628(.d_in(u_ca_in_628), .d_out(u_ca_out_628));
compressor_162_48 u_ca_162_48_629(.d_in(u_ca_in_629), .d_out(u_ca_out_629));
compressor_162_48 u_ca_162_48_630(.d_in(u_ca_in_630), .d_out(u_ca_out_630));
compressor_162_48 u_ca_162_48_631(.d_in(u_ca_in_631), .d_out(u_ca_out_631));
compressor_162_48 u_ca_162_48_632(.d_in(u_ca_in_632), .d_out(u_ca_out_632));
compressor_162_48 u_ca_162_48_633(.d_in(u_ca_in_633), .d_out(u_ca_out_633));
compressor_162_48 u_ca_162_48_634(.d_in(u_ca_in_634), .d_out(u_ca_out_634));
compressor_162_48 u_ca_162_48_635(.d_in(u_ca_in_635), .d_out(u_ca_out_635));
compressor_162_48 u_ca_162_48_636(.d_in(u_ca_in_636), .d_out(u_ca_out_636));
compressor_162_48 u_ca_162_48_637(.d_in(u_ca_in_637), .d_out(u_ca_out_637));
compressor_162_48 u_ca_162_48_638(.d_in(u_ca_in_638), .d_out(u_ca_out_638));
compressor_162_48 u_ca_162_48_639(.d_in(u_ca_in_639), .d_out(u_ca_out_639));
compressor_162_48 u_ca_162_48_640(.d_in(u_ca_in_640), .d_out(u_ca_out_640));
compressor_162_48 u_ca_162_48_641(.d_in(u_ca_in_641), .d_out(u_ca_out_641));
compressor_162_48 u_ca_162_48_642(.d_in(u_ca_in_642), .d_out(u_ca_out_642));
compressor_162_48 u_ca_162_48_643(.d_in(u_ca_in_643), .d_out(u_ca_out_643));
compressor_162_48 u_ca_162_48_644(.d_in(u_ca_in_644), .d_out(u_ca_out_644));
compressor_162_48 u_ca_162_48_645(.d_in(u_ca_in_645), .d_out(u_ca_out_645));
compressor_162_48 u_ca_162_48_646(.d_in(u_ca_in_646), .d_out(u_ca_out_646));
compressor_162_48 u_ca_162_48_647(.d_in(u_ca_in_647), .d_out(u_ca_out_647));
compressor_162_48 u_ca_162_48_648(.d_in(u_ca_in_648), .d_out(u_ca_out_648));
compressor_162_48 u_ca_162_48_649(.d_in(u_ca_in_649), .d_out(u_ca_out_649));
compressor_162_48 u_ca_162_48_650(.d_in(u_ca_in_650), .d_out(u_ca_out_650));
compressor_162_48 u_ca_162_48_651(.d_in(u_ca_in_651), .d_out(u_ca_out_651));
compressor_162_48 u_ca_162_48_652(.d_in(u_ca_in_652), .d_out(u_ca_out_652));
compressor_162_48 u_ca_162_48_653(.d_in(u_ca_in_653), .d_out(u_ca_out_653));
compressor_162_48 u_ca_162_48_654(.d_in(u_ca_in_654), .d_out(u_ca_out_654));
compressor_162_48 u_ca_162_48_655(.d_in(u_ca_in_655), .d_out(u_ca_out_655));
compressor_162_48 u_ca_162_48_656(.d_in(u_ca_in_656), .d_out(u_ca_out_656));
compressor_162_48 u_ca_162_48_657(.d_in(u_ca_in_657), .d_out(u_ca_out_657));
compressor_162_48 u_ca_162_48_658(.d_in(u_ca_in_658), .d_out(u_ca_out_658));
compressor_162_48 u_ca_162_48_659(.d_in(u_ca_in_659), .d_out(u_ca_out_659));
compressor_162_48 u_ca_162_48_660(.d_in(u_ca_in_660), .d_out(u_ca_out_660));
compressor_162_48 u_ca_162_48_661(.d_in(u_ca_in_661), .d_out(u_ca_out_661));
compressor_162_48 u_ca_162_48_662(.d_in(u_ca_in_662), .d_out(u_ca_out_662));
compressor_162_48 u_ca_162_48_663(.d_in(u_ca_in_663), .d_out(u_ca_out_663));
compressor_162_48 u_ca_162_48_664(.d_in(u_ca_in_664), .d_out(u_ca_out_664));
compressor_162_48 u_ca_162_48_665(.d_in(u_ca_in_665), .d_out(u_ca_out_665));
compressor_162_48 u_ca_162_48_666(.d_in(u_ca_in_666), .d_out(u_ca_out_666));
compressor_162_48 u_ca_162_48_667(.d_in(u_ca_in_667), .d_out(u_ca_out_667));
compressor_162_48 u_ca_162_48_668(.d_in(u_ca_in_668), .d_out(u_ca_out_668));
compressor_162_48 u_ca_162_48_669(.d_in(u_ca_in_669), .d_out(u_ca_out_669));
compressor_162_48 u_ca_162_48_670(.d_in(u_ca_in_670), .d_out(u_ca_out_670));
compressor_162_48 u_ca_162_48_671(.d_in(u_ca_in_671), .d_out(u_ca_out_671));
compressor_162_48 u_ca_162_48_672(.d_in(u_ca_in_672), .d_out(u_ca_out_672));
compressor_162_48 u_ca_162_48_673(.d_in(u_ca_in_673), .d_out(u_ca_out_673));
compressor_162_48 u_ca_162_48_674(.d_in(u_ca_in_674), .d_out(u_ca_out_674));
compressor_162_48 u_ca_162_48_675(.d_in(u_ca_in_675), .d_out(u_ca_out_675));
compressor_162_48 u_ca_162_48_676(.d_in(u_ca_in_676), .d_out(u_ca_out_676));
compressor_162_48 u_ca_162_48_677(.d_in(u_ca_in_677), .d_out(u_ca_out_677));
compressor_162_48 u_ca_162_48_678(.d_in(u_ca_in_678), .d_out(u_ca_out_678));
compressor_162_48 u_ca_162_48_679(.d_in(u_ca_in_679), .d_out(u_ca_out_679));
compressor_162_48 u_ca_162_48_680(.d_in(u_ca_in_680), .d_out(u_ca_out_680));
compressor_162_48 u_ca_162_48_681(.d_in(u_ca_in_681), .d_out(u_ca_out_681));
compressor_162_48 u_ca_162_48_682(.d_in(u_ca_in_682), .d_out(u_ca_out_682));
compressor_162_48 u_ca_162_48_683(.d_in(u_ca_in_683), .d_out(u_ca_out_683));
compressor_162_48 u_ca_162_48_684(.d_in(u_ca_in_684), .d_out(u_ca_out_684));
compressor_162_48 u_ca_162_48_685(.d_in(u_ca_in_685), .d_out(u_ca_out_685));
compressor_162_48 u_ca_162_48_686(.d_in(u_ca_in_686), .d_out(u_ca_out_686));
compressor_162_48 u_ca_162_48_687(.d_in(u_ca_in_687), .d_out(u_ca_out_687));
compressor_162_48 u_ca_162_48_688(.d_in(u_ca_in_688), .d_out(u_ca_out_688));
compressor_162_48 u_ca_162_48_689(.d_in(u_ca_in_689), .d_out(u_ca_out_689));
compressor_162_48 u_ca_162_48_690(.d_in(u_ca_in_690), .d_out(u_ca_out_690));
compressor_162_48 u_ca_162_48_691(.d_in(u_ca_in_691), .d_out(u_ca_out_691));
compressor_162_48 u_ca_162_48_692(.d_in(u_ca_in_692), .d_out(u_ca_out_692));
compressor_162_48 u_ca_162_48_693(.d_in(u_ca_in_693), .d_out(u_ca_out_693));
compressor_162_48 u_ca_162_48_694(.d_in(u_ca_in_694), .d_out(u_ca_out_694));
compressor_162_48 u_ca_162_48_695(.d_in(u_ca_in_695), .d_out(u_ca_out_695));
compressor_162_48 u_ca_162_48_696(.d_in(u_ca_in_696), .d_out(u_ca_out_696));
compressor_162_48 u_ca_162_48_697(.d_in(u_ca_in_697), .d_out(u_ca_out_697));
compressor_162_48 u_ca_162_48_698(.d_in(u_ca_in_698), .d_out(u_ca_out_698));
compressor_162_48 u_ca_162_48_699(.d_in(u_ca_in_699), .d_out(u_ca_out_699));
compressor_162_48 u_ca_162_48_700(.d_in(u_ca_in_700), .d_out(u_ca_out_700));
compressor_162_48 u_ca_162_48_701(.d_in(u_ca_in_701), .d_out(u_ca_out_701));
compressor_162_48 u_ca_162_48_702(.d_in(u_ca_in_702), .d_out(u_ca_out_702));
compressor_162_48 u_ca_162_48_703(.d_in(u_ca_in_703), .d_out(u_ca_out_703));
compressor_162_48 u_ca_162_48_704(.d_in(u_ca_in_704), .d_out(u_ca_out_704));
compressor_162_48 u_ca_162_48_705(.d_in(u_ca_in_705), .d_out(u_ca_out_705));
compressor_162_48 u_ca_162_48_706(.d_in(u_ca_in_706), .d_out(u_ca_out_706));
compressor_162_48 u_ca_162_48_707(.d_in(u_ca_in_707), .d_out(u_ca_out_707));
compressor_162_48 u_ca_162_48_708(.d_in(u_ca_in_708), .d_out(u_ca_out_708));
compressor_162_48 u_ca_162_48_709(.d_in(u_ca_in_709), .d_out(u_ca_out_709));
compressor_162_48 u_ca_162_48_710(.d_in(u_ca_in_710), .d_out(u_ca_out_710));
compressor_162_48 u_ca_162_48_711(.d_in(u_ca_in_711), .d_out(u_ca_out_711));
compressor_162_48 u_ca_162_48_712(.d_in(u_ca_in_712), .d_out(u_ca_out_712));
compressor_162_48 u_ca_162_48_713(.d_in(u_ca_in_713), .d_out(u_ca_out_713));
compressor_162_48 u_ca_162_48_714(.d_in(u_ca_in_714), .d_out(u_ca_out_714));
compressor_162_48 u_ca_162_48_715(.d_in(u_ca_in_715), .d_out(u_ca_out_715));
compressor_162_48 u_ca_162_48_716(.d_in(u_ca_in_716), .d_out(u_ca_out_716));
compressor_162_48 u_ca_162_48_717(.d_in(u_ca_in_717), .d_out(u_ca_out_717));
compressor_162_48 u_ca_162_48_718(.d_in(u_ca_in_718), .d_out(u_ca_out_718));
compressor_162_48 u_ca_162_48_719(.d_in(u_ca_in_719), .d_out(u_ca_out_719));
compressor_162_48 u_ca_162_48_720(.d_in(u_ca_in_720), .d_out(u_ca_out_720));
compressor_162_48 u_ca_162_48_721(.d_in(u_ca_in_721), .d_out(u_ca_out_721));
compressor_162_48 u_ca_162_48_722(.d_in(u_ca_in_722), .d_out(u_ca_out_722));
compressor_162_48 u_ca_162_48_723(.d_in(u_ca_in_723), .d_out(u_ca_out_723));
compressor_162_48 u_ca_162_48_724(.d_in(u_ca_in_724), .d_out(u_ca_out_724));
compressor_162_48 u_ca_162_48_725(.d_in(u_ca_in_725), .d_out(u_ca_out_725));
compressor_162_48 u_ca_162_48_726(.d_in(u_ca_in_726), .d_out(u_ca_out_726));
compressor_162_48 u_ca_162_48_727(.d_in(u_ca_in_727), .d_out(u_ca_out_727));
compressor_162_48 u_ca_162_48_728(.d_in(u_ca_in_728), .d_out(u_ca_out_728));
compressor_162_48 u_ca_162_48_729(.d_in(u_ca_in_729), .d_out(u_ca_out_729));
compressor_162_48 u_ca_162_48_730(.d_in(u_ca_in_730), .d_out(u_ca_out_730));
compressor_162_48 u_ca_162_48_731(.d_in(u_ca_in_731), .d_out(u_ca_out_731));
compressor_162_48 u_ca_162_48_732(.d_in(u_ca_in_732), .d_out(u_ca_out_732));
compressor_162_48 u_ca_162_48_733(.d_in(u_ca_in_733), .d_out(u_ca_out_733));
compressor_162_48 u_ca_162_48_734(.d_in(u_ca_in_734), .d_out(u_ca_out_734));
compressor_162_48 u_ca_162_48_735(.d_in(u_ca_in_735), .d_out(u_ca_out_735));
compressor_162_48 u_ca_162_48_736(.d_in(u_ca_in_736), .d_out(u_ca_out_736));
compressor_162_48 u_ca_162_48_737(.d_in(u_ca_in_737), .d_out(u_ca_out_737));
compressor_162_48 u_ca_162_48_738(.d_in(u_ca_in_738), .d_out(u_ca_out_738));
compressor_162_48 u_ca_162_48_739(.d_in(u_ca_in_739), .d_out(u_ca_out_739));
compressor_162_48 u_ca_162_48_740(.d_in(u_ca_in_740), .d_out(u_ca_out_740));
compressor_162_48 u_ca_162_48_741(.d_in(u_ca_in_741), .d_out(u_ca_out_741));
compressor_162_48 u_ca_162_48_742(.d_in(u_ca_in_742), .d_out(u_ca_out_742));
compressor_162_48 u_ca_162_48_743(.d_in(u_ca_in_743), .d_out(u_ca_out_743));
compressor_162_48 u_ca_162_48_744(.d_in(u_ca_in_744), .d_out(u_ca_out_744));
compressor_162_48 u_ca_162_48_745(.d_in(u_ca_in_745), .d_out(u_ca_out_745));
compressor_162_48 u_ca_162_48_746(.d_in(u_ca_in_746), .d_out(u_ca_out_746));
compressor_162_48 u_ca_162_48_747(.d_in(u_ca_in_747), .d_out(u_ca_out_747));
compressor_162_48 u_ca_162_48_748(.d_in(u_ca_in_748), .d_out(u_ca_out_748));
compressor_162_48 u_ca_162_48_749(.d_in(u_ca_in_749), .d_out(u_ca_out_749));
compressor_162_48 u_ca_162_48_750(.d_in(u_ca_in_750), .d_out(u_ca_out_750));
compressor_162_48 u_ca_162_48_751(.d_in(u_ca_in_751), .d_out(u_ca_out_751));
compressor_162_48 u_ca_162_48_752(.d_in(u_ca_in_752), .d_out(u_ca_out_752));
compressor_162_48 u_ca_162_48_753(.d_in(u_ca_in_753), .d_out(u_ca_out_753));
compressor_162_48 u_ca_162_48_754(.d_in(u_ca_in_754), .d_out(u_ca_out_754));
compressor_162_48 u_ca_162_48_755(.d_in(u_ca_in_755), .d_out(u_ca_out_755));
compressor_162_48 u_ca_162_48_756(.d_in(u_ca_in_756), .d_out(u_ca_out_756));
compressor_162_48 u_ca_162_48_757(.d_in(u_ca_in_757), .d_out(u_ca_out_757));
compressor_162_48 u_ca_162_48_758(.d_in(u_ca_in_758), .d_out(u_ca_out_758));
compressor_162_48 u_ca_162_48_759(.d_in(u_ca_in_759), .d_out(u_ca_out_759));
compressor_162_48 u_ca_162_48_760(.d_in(u_ca_in_760), .d_out(u_ca_out_760));
compressor_162_48 u_ca_162_48_761(.d_in(u_ca_in_761), .d_out(u_ca_out_761));
compressor_162_48 u_ca_162_48_762(.d_in(u_ca_in_762), .d_out(u_ca_out_762));
compressor_162_48 u_ca_162_48_763(.d_in(u_ca_in_763), .d_out(u_ca_out_763));
compressor_162_48 u_ca_162_48_764(.d_in(u_ca_in_764), .d_out(u_ca_out_764));
compressor_162_48 u_ca_162_48_765(.d_in(u_ca_in_765), .d_out(u_ca_out_765));
compressor_162_48 u_ca_162_48_766(.d_in(u_ca_in_766), .d_out(u_ca_out_766));
compressor_162_48 u_ca_162_48_767(.d_in(u_ca_in_767), .d_out(u_ca_out_767));
compressor_162_48 u_ca_162_48_768(.d_in(u_ca_in_768), .d_out(u_ca_out_768));
compressor_162_48 u_ca_162_48_769(.d_in(u_ca_in_769), .d_out(u_ca_out_769));
compressor_162_48 u_ca_162_48_770(.d_in(u_ca_in_770), .d_out(u_ca_out_770));
compressor_162_48 u_ca_162_48_771(.d_in(u_ca_in_771), .d_out(u_ca_out_771));
compressor_162_48 u_ca_162_48_772(.d_in(u_ca_in_772), .d_out(u_ca_out_772));
compressor_162_48 u_ca_162_48_773(.d_in(u_ca_in_773), .d_out(u_ca_out_773));
compressor_162_48 u_ca_162_48_774(.d_in(u_ca_in_774), .d_out(u_ca_out_774));
compressor_162_48 u_ca_162_48_775(.d_in(u_ca_in_775), .d_out(u_ca_out_775));
compressor_162_48 u_ca_162_48_776(.d_in(u_ca_in_776), .d_out(u_ca_out_776));
compressor_162_48 u_ca_162_48_777(.d_in(u_ca_in_777), .d_out(u_ca_out_777));
compressor_162_48 u_ca_162_48_778(.d_in(u_ca_in_778), .d_out(u_ca_out_778));
compressor_162_48 u_ca_162_48_779(.d_in(u_ca_in_779), .d_out(u_ca_out_779));
compressor_162_48 u_ca_162_48_780(.d_in(u_ca_in_780), .d_out(u_ca_out_780));
compressor_162_48 u_ca_162_48_781(.d_in(u_ca_in_781), .d_out(u_ca_out_781));
compressor_162_48 u_ca_162_48_782(.d_in(u_ca_in_782), .d_out(u_ca_out_782));
compressor_162_48 u_ca_162_48_783(.d_in(u_ca_in_783), .d_out(u_ca_out_783));
compressor_162_48 u_ca_162_48_784(.d_in(u_ca_in_784), .d_out(u_ca_out_784));
compressor_162_48 u_ca_162_48_785(.d_in(u_ca_in_785), .d_out(u_ca_out_785));
compressor_162_48 u_ca_162_48_786(.d_in(u_ca_in_786), .d_out(u_ca_out_786));
compressor_162_48 u_ca_162_48_787(.d_in(u_ca_in_787), .d_out(u_ca_out_787));
compressor_162_48 u_ca_162_48_788(.d_in(u_ca_in_788), .d_out(u_ca_out_788));
compressor_162_48 u_ca_162_48_789(.d_in(u_ca_in_789), .d_out(u_ca_out_789));
compressor_162_48 u_ca_162_48_790(.d_in(u_ca_in_790), .d_out(u_ca_out_790));
compressor_162_48 u_ca_162_48_791(.d_in(u_ca_in_791), .d_out(u_ca_out_791));
compressor_162_48 u_ca_162_48_792(.d_in(u_ca_in_792), .d_out(u_ca_out_792));
compressor_162_48 u_ca_162_48_793(.d_in(u_ca_in_793), .d_out(u_ca_out_793));
compressor_162_48 u_ca_162_48_794(.d_in(u_ca_in_794), .d_out(u_ca_out_794));
compressor_162_48 u_ca_162_48_795(.d_in(u_ca_in_795), .d_out(u_ca_out_795));
compressor_162_48 u_ca_162_48_796(.d_in(u_ca_in_796), .d_out(u_ca_out_796));
compressor_162_48 u_ca_162_48_797(.d_in(u_ca_in_797), .d_out(u_ca_out_797));
compressor_162_48 u_ca_162_48_798(.d_in(u_ca_in_798), .d_out(u_ca_out_798));
compressor_162_48 u_ca_162_48_799(.d_in(u_ca_in_799), .d_out(u_ca_out_799));
compressor_162_48 u_ca_162_48_800(.d_in(u_ca_in_800), .d_out(u_ca_out_800));
compressor_162_48 u_ca_162_48_801(.d_in(u_ca_in_801), .d_out(u_ca_out_801));
compressor_162_48 u_ca_162_48_802(.d_in(u_ca_in_802), .d_out(u_ca_out_802));
compressor_162_48 u_ca_162_48_803(.d_in(u_ca_in_803), .d_out(u_ca_out_803));
compressor_162_48 u_ca_162_48_804(.d_in(u_ca_in_804), .d_out(u_ca_out_804));
compressor_162_48 u_ca_162_48_805(.d_in(u_ca_in_805), .d_out(u_ca_out_805));
compressor_162_48 u_ca_162_48_806(.d_in(u_ca_in_806), .d_out(u_ca_out_806));
compressor_162_48 u_ca_162_48_807(.d_in(u_ca_in_807), .d_out(u_ca_out_807));
compressor_162_48 u_ca_162_48_808(.d_in(u_ca_in_808), .d_out(u_ca_out_808));
compressor_162_48 u_ca_162_48_809(.d_in(u_ca_in_809), .d_out(u_ca_out_809));
compressor_162_48 u_ca_162_48_810(.d_in(u_ca_in_810), .d_out(u_ca_out_810));
compressor_162_48 u_ca_162_48_811(.d_in(u_ca_in_811), .d_out(u_ca_out_811));
compressor_162_48 u_ca_162_48_812(.d_in(u_ca_in_812), .d_out(u_ca_out_812));
compressor_162_48 u_ca_162_48_813(.d_in(u_ca_in_813), .d_out(u_ca_out_813));
compressor_162_48 u_ca_162_48_814(.d_in(u_ca_in_814), .d_out(u_ca_out_814));
compressor_162_48 u_ca_162_48_815(.d_in(u_ca_in_815), .d_out(u_ca_out_815));
compressor_162_48 u_ca_162_48_816(.d_in(u_ca_in_816), .d_out(u_ca_out_816));
compressor_162_48 u_ca_162_48_817(.d_in(u_ca_in_817), .d_out(u_ca_out_817));
compressor_162_48 u_ca_162_48_818(.d_in(u_ca_in_818), .d_out(u_ca_out_818));
compressor_162_48 u_ca_162_48_819(.d_in(u_ca_in_819), .d_out(u_ca_out_819));
compressor_162_48 u_ca_162_48_820(.d_in(u_ca_in_820), .d_out(u_ca_out_820));
compressor_162_48 u_ca_162_48_821(.d_in(u_ca_in_821), .d_out(u_ca_out_821));
compressor_162_48 u_ca_162_48_822(.d_in(u_ca_in_822), .d_out(u_ca_out_822));
compressor_162_48 u_ca_162_48_823(.d_in(u_ca_in_823), .d_out(u_ca_out_823));
compressor_162_48 u_ca_162_48_824(.d_in(u_ca_in_824), .d_out(u_ca_out_824));
compressor_162_48 u_ca_162_48_825(.d_in(u_ca_in_825), .d_out(u_ca_out_825));
compressor_162_48 u_ca_162_48_826(.d_in(u_ca_in_826), .d_out(u_ca_out_826));
compressor_162_48 u_ca_162_48_827(.d_in(u_ca_in_827), .d_out(u_ca_out_827));
compressor_162_48 u_ca_162_48_828(.d_in(u_ca_in_828), .d_out(u_ca_out_828));
compressor_162_48 u_ca_162_48_829(.d_in(u_ca_in_829), .d_out(u_ca_out_829));
compressor_162_48 u_ca_162_48_830(.d_in(u_ca_in_830), .d_out(u_ca_out_830));
compressor_162_48 u_ca_162_48_831(.d_in(u_ca_in_831), .d_out(u_ca_out_831));
compressor_162_48 u_ca_162_48_832(.d_in(u_ca_in_832), .d_out(u_ca_out_832));
compressor_162_48 u_ca_162_48_833(.d_in(u_ca_in_833), .d_out(u_ca_out_833));
compressor_162_48 u_ca_162_48_834(.d_in(u_ca_in_834), .d_out(u_ca_out_834));
compressor_162_48 u_ca_162_48_835(.d_in(u_ca_in_835), .d_out(u_ca_out_835));
compressor_162_48 u_ca_162_48_836(.d_in(u_ca_in_836), .d_out(u_ca_out_836));
compressor_162_48 u_ca_162_48_837(.d_in(u_ca_in_837), .d_out(u_ca_out_837));
compressor_162_48 u_ca_162_48_838(.d_in(u_ca_in_838), .d_out(u_ca_out_838));
compressor_162_48 u_ca_162_48_839(.d_in(u_ca_in_839), .d_out(u_ca_out_839));
compressor_162_48 u_ca_162_48_840(.d_in(u_ca_in_840), .d_out(u_ca_out_840));
compressor_162_48 u_ca_162_48_841(.d_in(u_ca_in_841), .d_out(u_ca_out_841));
compressor_162_48 u_ca_162_48_842(.d_in(u_ca_in_842), .d_out(u_ca_out_842));
compressor_162_48 u_ca_162_48_843(.d_in(u_ca_in_843), .d_out(u_ca_out_843));
compressor_162_48 u_ca_162_48_844(.d_in(u_ca_in_844), .d_out(u_ca_out_844));
compressor_162_48 u_ca_162_48_845(.d_in(u_ca_in_845), .d_out(u_ca_out_845));
compressor_162_48 u_ca_162_48_846(.d_in(u_ca_in_846), .d_out(u_ca_out_846));
compressor_162_48 u_ca_162_48_847(.d_in(u_ca_in_847), .d_out(u_ca_out_847));
compressor_162_48 u_ca_162_48_848(.d_in(u_ca_in_848), .d_out(u_ca_out_848));
compressor_162_48 u_ca_162_48_849(.d_in(u_ca_in_849), .d_out(u_ca_out_849));
compressor_162_48 u_ca_162_48_850(.d_in(u_ca_in_850), .d_out(u_ca_out_850));
compressor_162_48 u_ca_162_48_851(.d_in(u_ca_in_851), .d_out(u_ca_out_851));
compressor_162_48 u_ca_162_48_852(.d_in(u_ca_in_852), .d_out(u_ca_out_852));
compressor_162_48 u_ca_162_48_853(.d_in(u_ca_in_853), .d_out(u_ca_out_853));
compressor_162_48 u_ca_162_48_854(.d_in(u_ca_in_854), .d_out(u_ca_out_854));
compressor_162_48 u_ca_162_48_855(.d_in(u_ca_in_855), .d_out(u_ca_out_855));
compressor_162_48 u_ca_162_48_856(.d_in(u_ca_in_856), .d_out(u_ca_out_856));
compressor_162_48 u_ca_162_48_857(.d_in(u_ca_in_857), .d_out(u_ca_out_857));
compressor_162_48 u_ca_162_48_858(.d_in(u_ca_in_858), .d_out(u_ca_out_858));
compressor_162_48 u_ca_162_48_859(.d_in(u_ca_in_859), .d_out(u_ca_out_859));
compressor_162_48 u_ca_162_48_860(.d_in(u_ca_in_860), .d_out(u_ca_out_860));
compressor_162_48 u_ca_162_48_861(.d_in(u_ca_in_861), .d_out(u_ca_out_861));
compressor_162_48 u_ca_162_48_862(.d_in(u_ca_in_862), .d_out(u_ca_out_862));
compressor_162_48 u_ca_162_48_863(.d_in(u_ca_in_863), .d_out(u_ca_out_863));
compressor_162_48 u_ca_162_48_864(.d_in(u_ca_in_864), .d_out(u_ca_out_864));
compressor_162_48 u_ca_162_48_865(.d_in(u_ca_in_865), .d_out(u_ca_out_865));
compressor_162_48 u_ca_162_48_866(.d_in(u_ca_in_866), .d_out(u_ca_out_866));
compressor_162_48 u_ca_162_48_867(.d_in(u_ca_in_867), .d_out(u_ca_out_867));
compressor_162_48 u_ca_162_48_868(.d_in(u_ca_in_868), .d_out(u_ca_out_868));
compressor_162_48 u_ca_162_48_869(.d_in(u_ca_in_869), .d_out(u_ca_out_869));
compressor_162_48 u_ca_162_48_870(.d_in(u_ca_in_870), .d_out(u_ca_out_870));
compressor_162_48 u_ca_162_48_871(.d_in(u_ca_in_871), .d_out(u_ca_out_871));
compressor_162_48 u_ca_162_48_872(.d_in(u_ca_in_872), .d_out(u_ca_out_872));
compressor_162_48 u_ca_162_48_873(.d_in(u_ca_in_873), .d_out(u_ca_out_873));
compressor_162_48 u_ca_162_48_874(.d_in(u_ca_in_874), .d_out(u_ca_out_874));
compressor_162_48 u_ca_162_48_875(.d_in(u_ca_in_875), .d_out(u_ca_out_875));
compressor_162_48 u_ca_162_48_876(.d_in(u_ca_in_876), .d_out(u_ca_out_876));
compressor_162_48 u_ca_162_48_877(.d_in(u_ca_in_877), .d_out(u_ca_out_877));
compressor_162_48 u_ca_162_48_878(.d_in(u_ca_in_878), .d_out(u_ca_out_878));
compressor_162_48 u_ca_162_48_879(.d_in(u_ca_in_879), .d_out(u_ca_out_879));
compressor_162_48 u_ca_162_48_880(.d_in(u_ca_in_880), .d_out(u_ca_out_880));
compressor_162_48 u_ca_162_48_881(.d_in(u_ca_in_881), .d_out(u_ca_out_881));
compressor_162_48 u_ca_162_48_882(.d_in(u_ca_in_882), .d_out(u_ca_out_882));
compressor_162_48 u_ca_162_48_883(.d_in(u_ca_in_883), .d_out(u_ca_out_883));
compressor_162_48 u_ca_162_48_884(.d_in(u_ca_in_884), .d_out(u_ca_out_884));
compressor_162_48 u_ca_162_48_885(.d_in(u_ca_in_885), .d_out(u_ca_out_885));
compressor_162_48 u_ca_162_48_886(.d_in(u_ca_in_886), .d_out(u_ca_out_886));
compressor_162_48 u_ca_162_48_887(.d_in(u_ca_in_887), .d_out(u_ca_out_887));
compressor_162_48 u_ca_162_48_888(.d_in(u_ca_in_888), .d_out(u_ca_out_888));
compressor_162_48 u_ca_162_48_889(.d_in(u_ca_in_889), .d_out(u_ca_out_889));
compressor_162_48 u_ca_162_48_890(.d_in(u_ca_in_890), .d_out(u_ca_out_890));
compressor_162_48 u_ca_162_48_891(.d_in(u_ca_in_891), .d_out(u_ca_out_891));
compressor_162_48 u_ca_162_48_892(.d_in(u_ca_in_892), .d_out(u_ca_out_892));
compressor_162_48 u_ca_162_48_893(.d_in(u_ca_in_893), .d_out(u_ca_out_893));
compressor_162_48 u_ca_162_48_894(.d_in(u_ca_in_894), .d_out(u_ca_out_894));
compressor_162_48 u_ca_162_48_895(.d_in(u_ca_in_895), .d_out(u_ca_out_895));
compressor_162_48 u_ca_162_48_896(.d_in(u_ca_in_896), .d_out(u_ca_out_896));
compressor_162_48 u_ca_162_48_897(.d_in(u_ca_in_897), .d_out(u_ca_out_897));
compressor_162_48 u_ca_162_48_898(.d_in(u_ca_in_898), .d_out(u_ca_out_898));
compressor_162_48 u_ca_162_48_899(.d_in(u_ca_in_899), .d_out(u_ca_out_899));
compressor_162_48 u_ca_162_48_900(.d_in(u_ca_in_900), .d_out(u_ca_out_900));
compressor_162_48 u_ca_162_48_901(.d_in(u_ca_in_901), .d_out(u_ca_out_901));
compressor_162_48 u_ca_162_48_902(.d_in(u_ca_in_902), .d_out(u_ca_out_902));
compressor_162_48 u_ca_162_48_903(.d_in(u_ca_in_903), .d_out(u_ca_out_903));
compressor_162_48 u_ca_162_48_904(.d_in(u_ca_in_904), .d_out(u_ca_out_904));
compressor_162_48 u_ca_162_48_905(.d_in(u_ca_in_905), .d_out(u_ca_out_905));
compressor_162_48 u_ca_162_48_906(.d_in(u_ca_in_906), .d_out(u_ca_out_906));
compressor_162_48 u_ca_162_48_907(.d_in(u_ca_in_907), .d_out(u_ca_out_907));
compressor_162_48 u_ca_162_48_908(.d_in(u_ca_in_908), .d_out(u_ca_out_908));
compressor_162_48 u_ca_162_48_909(.d_in(u_ca_in_909), .d_out(u_ca_out_909));
compressor_162_48 u_ca_162_48_910(.d_in(u_ca_in_910), .d_out(u_ca_out_910));
compressor_162_48 u_ca_162_48_911(.d_in(u_ca_in_911), .d_out(u_ca_out_911));
compressor_162_48 u_ca_162_48_912(.d_in(u_ca_in_912), .d_out(u_ca_out_912));
compressor_162_48 u_ca_162_48_913(.d_in(u_ca_in_913), .d_out(u_ca_out_913));
compressor_162_48 u_ca_162_48_914(.d_in(u_ca_in_914), .d_out(u_ca_out_914));
compressor_162_48 u_ca_162_48_915(.d_in(u_ca_in_915), .d_out(u_ca_out_915));
compressor_162_48 u_ca_162_48_916(.d_in(u_ca_in_916), .d_out(u_ca_out_916));
compressor_162_48 u_ca_162_48_917(.d_in(u_ca_in_917), .d_out(u_ca_out_917));
compressor_162_48 u_ca_162_48_918(.d_in(u_ca_in_918), .d_out(u_ca_out_918));
compressor_162_48 u_ca_162_48_919(.d_in(u_ca_in_919), .d_out(u_ca_out_919));
compressor_162_48 u_ca_162_48_920(.d_in(u_ca_in_920), .d_out(u_ca_out_920));
compressor_162_48 u_ca_162_48_921(.d_in(u_ca_in_921), .d_out(u_ca_out_921));
compressor_162_48 u_ca_162_48_922(.d_in(u_ca_in_922), .d_out(u_ca_out_922));
compressor_162_48 u_ca_162_48_923(.d_in(u_ca_in_923), .d_out(u_ca_out_923));
compressor_162_48 u_ca_162_48_924(.d_in(u_ca_in_924), .d_out(u_ca_out_924));
compressor_162_48 u_ca_162_48_925(.d_in(u_ca_in_925), .d_out(u_ca_out_925));
compressor_162_48 u_ca_162_48_926(.d_in(u_ca_in_926), .d_out(u_ca_out_926));
compressor_162_48 u_ca_162_48_927(.d_in(u_ca_in_927), .d_out(u_ca_out_927));
compressor_162_48 u_ca_162_48_928(.d_in(u_ca_in_928), .d_out(u_ca_out_928));
compressor_162_48 u_ca_162_48_929(.d_in(u_ca_in_929), .d_out(u_ca_out_929));
compressor_162_48 u_ca_162_48_930(.d_in(u_ca_in_930), .d_out(u_ca_out_930));
compressor_162_48 u_ca_162_48_931(.d_in(u_ca_in_931), .d_out(u_ca_out_931));
compressor_162_48 u_ca_162_48_932(.d_in(u_ca_in_932), .d_out(u_ca_out_932));
compressor_162_48 u_ca_162_48_933(.d_in(u_ca_in_933), .d_out(u_ca_out_933));
compressor_162_48 u_ca_162_48_934(.d_in(u_ca_in_934), .d_out(u_ca_out_934));
compressor_162_48 u_ca_162_48_935(.d_in(u_ca_in_935), .d_out(u_ca_out_935));
compressor_162_48 u_ca_162_48_936(.d_in(u_ca_in_936), .d_out(u_ca_out_936));
compressor_162_48 u_ca_162_48_937(.d_in(u_ca_in_937), .d_out(u_ca_out_937));
compressor_162_48 u_ca_162_48_938(.d_in(u_ca_in_938), .d_out(u_ca_out_938));
compressor_162_48 u_ca_162_48_939(.d_in(u_ca_in_939), .d_out(u_ca_out_939));
compressor_162_48 u_ca_162_48_940(.d_in(u_ca_in_940), .d_out(u_ca_out_940));
compressor_162_48 u_ca_162_48_941(.d_in(u_ca_in_941), .d_out(u_ca_out_941));
compressor_162_48 u_ca_162_48_942(.d_in(u_ca_in_942), .d_out(u_ca_out_942));
compressor_162_48 u_ca_162_48_943(.d_in(u_ca_in_943), .d_out(u_ca_out_943));
compressor_162_48 u_ca_162_48_944(.d_in(u_ca_in_944), .d_out(u_ca_out_944));
compressor_162_48 u_ca_162_48_945(.d_in(u_ca_in_945), .d_out(u_ca_out_945));
compressor_162_48 u_ca_162_48_946(.d_in(u_ca_in_946), .d_out(u_ca_out_946));
compressor_162_48 u_ca_162_48_947(.d_in(u_ca_in_947), .d_out(u_ca_out_947));
compressor_162_48 u_ca_162_48_948(.d_in(u_ca_in_948), .d_out(u_ca_out_948));
compressor_162_48 u_ca_162_48_949(.d_in(u_ca_in_949), .d_out(u_ca_out_949));
compressor_162_48 u_ca_162_48_950(.d_in(u_ca_in_950), .d_out(u_ca_out_950));
compressor_162_48 u_ca_162_48_951(.d_in(u_ca_in_951), .d_out(u_ca_out_951));
compressor_162_48 u_ca_162_48_952(.d_in(u_ca_in_952), .d_out(u_ca_out_952));
compressor_162_48 u_ca_162_48_953(.d_in(u_ca_in_953), .d_out(u_ca_out_953));
compressor_162_48 u_ca_162_48_954(.d_in(u_ca_in_954), .d_out(u_ca_out_954));
compressor_162_48 u_ca_162_48_955(.d_in(u_ca_in_955), .d_out(u_ca_out_955));
compressor_162_48 u_ca_162_48_956(.d_in(u_ca_in_956), .d_out(u_ca_out_956));
compressor_162_48 u_ca_162_48_957(.d_in(u_ca_in_957), .d_out(u_ca_out_957));
compressor_162_48 u_ca_162_48_958(.d_in(u_ca_in_958), .d_out(u_ca_out_958));
compressor_162_48 u_ca_162_48_959(.d_in(u_ca_in_959), .d_out(u_ca_out_959));
compressor_162_48 u_ca_162_48_960(.d_in(u_ca_in_960), .d_out(u_ca_out_960));
compressor_162_48 u_ca_162_48_961(.d_in(u_ca_in_961), .d_out(u_ca_out_961));
compressor_162_48 u_ca_162_48_962(.d_in(u_ca_in_962), .d_out(u_ca_out_962));
compressor_162_48 u_ca_162_48_963(.d_in(u_ca_in_963), .d_out(u_ca_out_963));
compressor_162_48 u_ca_162_48_964(.d_in(u_ca_in_964), .d_out(u_ca_out_964));
compressor_162_48 u_ca_162_48_965(.d_in(u_ca_in_965), .d_out(u_ca_out_965));
compressor_162_48 u_ca_162_48_966(.d_in(u_ca_in_966), .d_out(u_ca_out_966));
compressor_162_48 u_ca_162_48_967(.d_in(u_ca_in_967), .d_out(u_ca_out_967));
compressor_162_48 u_ca_162_48_968(.d_in(u_ca_in_968), .d_out(u_ca_out_968));
compressor_162_48 u_ca_162_48_969(.d_in(u_ca_in_969), .d_out(u_ca_out_969));
compressor_162_48 u_ca_162_48_970(.d_in(u_ca_in_970), .d_out(u_ca_out_970));
compressor_162_48 u_ca_162_48_971(.d_in(u_ca_in_971), .d_out(u_ca_out_971));
compressor_162_48 u_ca_162_48_972(.d_in(u_ca_in_972), .d_out(u_ca_out_972));
compressor_162_48 u_ca_162_48_973(.d_in(u_ca_in_973), .d_out(u_ca_out_973));
compressor_162_48 u_ca_162_48_974(.d_in(u_ca_in_974), .d_out(u_ca_out_974));
compressor_162_48 u_ca_162_48_975(.d_in(u_ca_in_975), .d_out(u_ca_out_975));
compressor_162_48 u_ca_162_48_976(.d_in(u_ca_in_976), .d_out(u_ca_out_976));
compressor_162_48 u_ca_162_48_977(.d_in(u_ca_in_977), .d_out(u_ca_out_977));
compressor_162_48 u_ca_162_48_978(.d_in(u_ca_in_978), .d_out(u_ca_out_978));
compressor_162_48 u_ca_162_48_979(.d_in(u_ca_in_979), .d_out(u_ca_out_979));
compressor_162_48 u_ca_162_48_980(.d_in(u_ca_in_980), .d_out(u_ca_out_980));
compressor_162_48 u_ca_162_48_981(.d_in(u_ca_in_981), .d_out(u_ca_out_981));
compressor_162_48 u_ca_162_48_982(.d_in(u_ca_in_982), .d_out(u_ca_out_982));
compressor_162_48 u_ca_162_48_983(.d_in(u_ca_in_983), .d_out(u_ca_out_983));
compressor_162_48 u_ca_162_48_984(.d_in(u_ca_in_984), .d_out(u_ca_out_984));
compressor_162_48 u_ca_162_48_985(.d_in(u_ca_in_985), .d_out(u_ca_out_985));
compressor_162_48 u_ca_162_48_986(.d_in(u_ca_in_986), .d_out(u_ca_out_986));
compressor_162_48 u_ca_162_48_987(.d_in(u_ca_in_987), .d_out(u_ca_out_987));
compressor_162_48 u_ca_162_48_988(.d_in(u_ca_in_988), .d_out(u_ca_out_988));
compressor_162_48 u_ca_162_48_989(.d_in(u_ca_in_989), .d_out(u_ca_out_989));
compressor_162_48 u_ca_162_48_990(.d_in(u_ca_in_990), .d_out(u_ca_out_990));
compressor_162_48 u_ca_162_48_991(.d_in(u_ca_in_991), .d_out(u_ca_out_991));
compressor_162_48 u_ca_162_48_992(.d_in(u_ca_in_992), .d_out(u_ca_out_992));
compressor_162_48 u_ca_162_48_993(.d_in(u_ca_in_993), .d_out(u_ca_out_993));
compressor_162_48 u_ca_162_48_994(.d_in(u_ca_in_994), .d_out(u_ca_out_994));
compressor_162_48 u_ca_162_48_995(.d_in(u_ca_in_995), .d_out(u_ca_out_995));
compressor_162_48 u_ca_162_48_996(.d_in(u_ca_in_996), .d_out(u_ca_out_996));
compressor_162_48 u_ca_162_48_997(.d_in(u_ca_in_997), .d_out(u_ca_out_997));
compressor_162_48 u_ca_162_48_998(.d_in(u_ca_in_998), .d_out(u_ca_out_998));
compressor_162_48 u_ca_162_48_999(.d_in(u_ca_in_999), .d_out(u_ca_out_999));
compressor_162_48 u_ca_162_48_1000(.d_in(u_ca_in_1000), .d_out(u_ca_out_1000));
compressor_162_48 u_ca_162_48_1001(.d_in(u_ca_in_1001), .d_out(u_ca_out_1001));
compressor_162_48 u_ca_162_48_1002(.d_in(u_ca_in_1002), .d_out(u_ca_out_1002));
compressor_162_48 u_ca_162_48_1003(.d_in(u_ca_in_1003), .d_out(u_ca_out_1003));
compressor_162_48 u_ca_162_48_1004(.d_in(u_ca_in_1004), .d_out(u_ca_out_1004));
compressor_162_48 u_ca_162_48_1005(.d_in(u_ca_in_1005), .d_out(u_ca_out_1005));
compressor_162_48 u_ca_162_48_1006(.d_in(u_ca_in_1006), .d_out(u_ca_out_1006));
compressor_162_48 u_ca_162_48_1007(.d_in(u_ca_in_1007), .d_out(u_ca_out_1007));
compressor_162_48 u_ca_162_48_1008(.d_in(u_ca_in_1008), .d_out(u_ca_out_1008));
compressor_162_48 u_ca_162_48_1009(.d_in(u_ca_in_1009), .d_out(u_ca_out_1009));
compressor_162_48 u_ca_162_48_1010(.d_in(u_ca_in_1010), .d_out(u_ca_out_1010));
compressor_162_48 u_ca_162_48_1011(.d_in(u_ca_in_1011), .d_out(u_ca_out_1011));
compressor_162_48 u_ca_162_48_1012(.d_in(u_ca_in_1012), .d_out(u_ca_out_1012));
compressor_162_48 u_ca_162_48_1013(.d_in(u_ca_in_1013), .d_out(u_ca_out_1013));
compressor_162_48 u_ca_162_48_1014(.d_in(u_ca_in_1014), .d_out(u_ca_out_1014));
compressor_162_48 u_ca_162_48_1015(.d_in(u_ca_in_1015), .d_out(u_ca_out_1015));
compressor_162_48 u_ca_162_48_1016(.d_in(u_ca_in_1016), .d_out(u_ca_out_1016));
compressor_162_48 u_ca_162_48_1017(.d_in(u_ca_in_1017), .d_out(u_ca_out_1017));
compressor_162_48 u_ca_162_48_1018(.d_in(u_ca_in_1018), .d_out(u_ca_out_1018));
compressor_162_48 u_ca_162_48_1019(.d_in(u_ca_in_1019), .d_out(u_ca_out_1019));
compressor_162_48 u_ca_162_48_1020(.d_in(u_ca_in_1020), .d_out(u_ca_out_1020));
compressor_162_48 u_ca_162_48_1021(.d_in(u_ca_in_1021), .d_out(u_ca_out_1021));
compressor_162_48 u_ca_162_48_1022(.d_in(u_ca_in_1022), .d_out(u_ca_out_1022));
compressor_162_48 u_ca_162_48_1023(.d_in(u_ca_in_1023), .d_out(u_ca_out_1023));
compressor_162_48 u_ca_162_48_1024(.d_in(u_ca_in_1024), .d_out(u_ca_out_1024));
compressor_162_48 u_ca_162_48_1025(.d_in(u_ca_in_1025), .d_out(u_ca_out_1025));
compressor_162_48 u_ca_162_48_1026(.d_in(u_ca_in_1026), .d_out(u_ca_out_1026));

//---------------------------------------------------------



//--output-------------------------------------------------

assign col_out_0 = {{42{1'b0}}, u_ca_out_0[5:0]};
assign col_out_1 = {{24{1'b0}}, u_ca_out_1[5:0], u_ca_out_0[23:6]};
assign col_out_2 = {{6{1'b0}}, u_ca_out_2[5:0], u_ca_out_1[23:6], u_ca_out_0[41:24]};
assign col_out_3 = {u_ca_out_3[5:0],u_ca_out_2[23:6], u_ca_out_1[41:24], u_ca_out_0[47:42]};
assign col_out_4 = {u_ca_out_4[5:0],u_ca_out_3[23:6], u_ca_out_2[41:24], u_ca_out_1[47:42]};
assign col_out_5 = {u_ca_out_5[5:0],u_ca_out_4[23:6], u_ca_out_3[41:24], u_ca_out_2[47:42]};
assign col_out_6 = {u_ca_out_6[5:0],u_ca_out_5[23:6], u_ca_out_4[41:24], u_ca_out_3[47:42]};
assign col_out_7 = {u_ca_out_7[5:0],u_ca_out_6[23:6], u_ca_out_5[41:24], u_ca_out_4[47:42]};
assign col_out_8 = {u_ca_out_8[5:0],u_ca_out_7[23:6], u_ca_out_6[41:24], u_ca_out_5[47:42]};
assign col_out_9 = {u_ca_out_9[5:0],u_ca_out_8[23:6], u_ca_out_7[41:24], u_ca_out_6[47:42]};
assign col_out_10 = {u_ca_out_10[5:0],u_ca_out_9[23:6], u_ca_out_8[41:24], u_ca_out_7[47:42]};
assign col_out_11 = {u_ca_out_11[5:0],u_ca_out_10[23:6], u_ca_out_9[41:24], u_ca_out_8[47:42]};
assign col_out_12 = {u_ca_out_12[5:0],u_ca_out_11[23:6], u_ca_out_10[41:24], u_ca_out_9[47:42]};
assign col_out_13 = {u_ca_out_13[5:0],u_ca_out_12[23:6], u_ca_out_11[41:24], u_ca_out_10[47:42]};
assign col_out_14 = {u_ca_out_14[5:0],u_ca_out_13[23:6], u_ca_out_12[41:24], u_ca_out_11[47:42]};
assign col_out_15 = {u_ca_out_15[5:0],u_ca_out_14[23:6], u_ca_out_13[41:24], u_ca_out_12[47:42]};
assign col_out_16 = {u_ca_out_16[5:0],u_ca_out_15[23:6], u_ca_out_14[41:24], u_ca_out_13[47:42]};
assign col_out_17 = {u_ca_out_17[5:0],u_ca_out_16[23:6], u_ca_out_15[41:24], u_ca_out_14[47:42]};
assign col_out_18 = {u_ca_out_18[5:0],u_ca_out_17[23:6], u_ca_out_16[41:24], u_ca_out_15[47:42]};
assign col_out_19 = {u_ca_out_19[5:0],u_ca_out_18[23:6], u_ca_out_17[41:24], u_ca_out_16[47:42]};
assign col_out_20 = {u_ca_out_20[5:0],u_ca_out_19[23:6], u_ca_out_18[41:24], u_ca_out_17[47:42]};
assign col_out_21 = {u_ca_out_21[5:0],u_ca_out_20[23:6], u_ca_out_19[41:24], u_ca_out_18[47:42]};
assign col_out_22 = {u_ca_out_22[5:0],u_ca_out_21[23:6], u_ca_out_20[41:24], u_ca_out_19[47:42]};
assign col_out_23 = {u_ca_out_23[5:0],u_ca_out_22[23:6], u_ca_out_21[41:24], u_ca_out_20[47:42]};
assign col_out_24 = {u_ca_out_24[5:0],u_ca_out_23[23:6], u_ca_out_22[41:24], u_ca_out_21[47:42]};
assign col_out_25 = {u_ca_out_25[5:0],u_ca_out_24[23:6], u_ca_out_23[41:24], u_ca_out_22[47:42]};
assign col_out_26 = {u_ca_out_26[5:0],u_ca_out_25[23:6], u_ca_out_24[41:24], u_ca_out_23[47:42]};
assign col_out_27 = {u_ca_out_27[5:0],u_ca_out_26[23:6], u_ca_out_25[41:24], u_ca_out_24[47:42]};
assign col_out_28 = {u_ca_out_28[5:0],u_ca_out_27[23:6], u_ca_out_26[41:24], u_ca_out_25[47:42]};
assign col_out_29 = {u_ca_out_29[5:0],u_ca_out_28[23:6], u_ca_out_27[41:24], u_ca_out_26[47:42]};
assign col_out_30 = {u_ca_out_30[5:0],u_ca_out_29[23:6], u_ca_out_28[41:24], u_ca_out_27[47:42]};
assign col_out_31 = {u_ca_out_31[5:0],u_ca_out_30[23:6], u_ca_out_29[41:24], u_ca_out_28[47:42]};
assign col_out_32 = {u_ca_out_32[5:0],u_ca_out_31[23:6], u_ca_out_30[41:24], u_ca_out_29[47:42]};
assign col_out_33 = {u_ca_out_33[5:0],u_ca_out_32[23:6], u_ca_out_31[41:24], u_ca_out_30[47:42]};
assign col_out_34 = {u_ca_out_34[5:0],u_ca_out_33[23:6], u_ca_out_32[41:24], u_ca_out_31[47:42]};
assign col_out_35 = {u_ca_out_35[5:0],u_ca_out_34[23:6], u_ca_out_33[41:24], u_ca_out_32[47:42]};
assign col_out_36 = {u_ca_out_36[5:0],u_ca_out_35[23:6], u_ca_out_34[41:24], u_ca_out_33[47:42]};
assign col_out_37 = {u_ca_out_37[5:0],u_ca_out_36[23:6], u_ca_out_35[41:24], u_ca_out_34[47:42]};
assign col_out_38 = {u_ca_out_38[5:0],u_ca_out_37[23:6], u_ca_out_36[41:24], u_ca_out_35[47:42]};
assign col_out_39 = {u_ca_out_39[5:0],u_ca_out_38[23:6], u_ca_out_37[41:24], u_ca_out_36[47:42]};
assign col_out_40 = {u_ca_out_40[5:0],u_ca_out_39[23:6], u_ca_out_38[41:24], u_ca_out_37[47:42]};
assign col_out_41 = {u_ca_out_41[5:0],u_ca_out_40[23:6], u_ca_out_39[41:24], u_ca_out_38[47:42]};
assign col_out_42 = {u_ca_out_42[5:0],u_ca_out_41[23:6], u_ca_out_40[41:24], u_ca_out_39[47:42]};
assign col_out_43 = {u_ca_out_43[5:0],u_ca_out_42[23:6], u_ca_out_41[41:24], u_ca_out_40[47:42]};
assign col_out_44 = {u_ca_out_44[5:0],u_ca_out_43[23:6], u_ca_out_42[41:24], u_ca_out_41[47:42]};
assign col_out_45 = {u_ca_out_45[5:0],u_ca_out_44[23:6], u_ca_out_43[41:24], u_ca_out_42[47:42]};
assign col_out_46 = {u_ca_out_46[5:0],u_ca_out_45[23:6], u_ca_out_44[41:24], u_ca_out_43[47:42]};
assign col_out_47 = {u_ca_out_47[5:0],u_ca_out_46[23:6], u_ca_out_45[41:24], u_ca_out_44[47:42]};
assign col_out_48 = {u_ca_out_48[5:0],u_ca_out_47[23:6], u_ca_out_46[41:24], u_ca_out_45[47:42]};
assign col_out_49 = {u_ca_out_49[5:0],u_ca_out_48[23:6], u_ca_out_47[41:24], u_ca_out_46[47:42]};
assign col_out_50 = {u_ca_out_50[5:0],u_ca_out_49[23:6], u_ca_out_48[41:24], u_ca_out_47[47:42]};
assign col_out_51 = {u_ca_out_51[5:0],u_ca_out_50[23:6], u_ca_out_49[41:24], u_ca_out_48[47:42]};
assign col_out_52 = {u_ca_out_52[5:0],u_ca_out_51[23:6], u_ca_out_50[41:24], u_ca_out_49[47:42]};
assign col_out_53 = {u_ca_out_53[5:0],u_ca_out_52[23:6], u_ca_out_51[41:24], u_ca_out_50[47:42]};
assign col_out_54 = {u_ca_out_54[5:0],u_ca_out_53[23:6], u_ca_out_52[41:24], u_ca_out_51[47:42]};
assign col_out_55 = {u_ca_out_55[5:0],u_ca_out_54[23:6], u_ca_out_53[41:24], u_ca_out_52[47:42]};
assign col_out_56 = {u_ca_out_56[5:0],u_ca_out_55[23:6], u_ca_out_54[41:24], u_ca_out_53[47:42]};
assign col_out_57 = {u_ca_out_57[5:0],u_ca_out_56[23:6], u_ca_out_55[41:24], u_ca_out_54[47:42]};
assign col_out_58 = {u_ca_out_58[5:0],u_ca_out_57[23:6], u_ca_out_56[41:24], u_ca_out_55[47:42]};
assign col_out_59 = {u_ca_out_59[5:0],u_ca_out_58[23:6], u_ca_out_57[41:24], u_ca_out_56[47:42]};
assign col_out_60 = {u_ca_out_60[5:0],u_ca_out_59[23:6], u_ca_out_58[41:24], u_ca_out_57[47:42]};
assign col_out_61 = {u_ca_out_61[5:0],u_ca_out_60[23:6], u_ca_out_59[41:24], u_ca_out_58[47:42]};
assign col_out_62 = {u_ca_out_62[5:0],u_ca_out_61[23:6], u_ca_out_60[41:24], u_ca_out_59[47:42]};
assign col_out_63 = {u_ca_out_63[5:0],u_ca_out_62[23:6], u_ca_out_61[41:24], u_ca_out_60[47:42]};
assign col_out_64 = {u_ca_out_64[5:0],u_ca_out_63[23:6], u_ca_out_62[41:24], u_ca_out_61[47:42]};
assign col_out_65 = {u_ca_out_65[5:0],u_ca_out_64[23:6], u_ca_out_63[41:24], u_ca_out_62[47:42]};
assign col_out_66 = {u_ca_out_66[5:0],u_ca_out_65[23:6], u_ca_out_64[41:24], u_ca_out_63[47:42]};
assign col_out_67 = {u_ca_out_67[5:0],u_ca_out_66[23:6], u_ca_out_65[41:24], u_ca_out_64[47:42]};
assign col_out_68 = {u_ca_out_68[5:0],u_ca_out_67[23:6], u_ca_out_66[41:24], u_ca_out_65[47:42]};
assign col_out_69 = {u_ca_out_69[5:0],u_ca_out_68[23:6], u_ca_out_67[41:24], u_ca_out_66[47:42]};
assign col_out_70 = {u_ca_out_70[5:0],u_ca_out_69[23:6], u_ca_out_68[41:24], u_ca_out_67[47:42]};
assign col_out_71 = {u_ca_out_71[5:0],u_ca_out_70[23:6], u_ca_out_69[41:24], u_ca_out_68[47:42]};
assign col_out_72 = {u_ca_out_72[5:0],u_ca_out_71[23:6], u_ca_out_70[41:24], u_ca_out_69[47:42]};
assign col_out_73 = {u_ca_out_73[5:0],u_ca_out_72[23:6], u_ca_out_71[41:24], u_ca_out_70[47:42]};
assign col_out_74 = {u_ca_out_74[5:0],u_ca_out_73[23:6], u_ca_out_72[41:24], u_ca_out_71[47:42]};
assign col_out_75 = {u_ca_out_75[5:0],u_ca_out_74[23:6], u_ca_out_73[41:24], u_ca_out_72[47:42]};
assign col_out_76 = {u_ca_out_76[5:0],u_ca_out_75[23:6], u_ca_out_74[41:24], u_ca_out_73[47:42]};
assign col_out_77 = {u_ca_out_77[5:0],u_ca_out_76[23:6], u_ca_out_75[41:24], u_ca_out_74[47:42]};
assign col_out_78 = {u_ca_out_78[5:0],u_ca_out_77[23:6], u_ca_out_76[41:24], u_ca_out_75[47:42]};
assign col_out_79 = {u_ca_out_79[5:0],u_ca_out_78[23:6], u_ca_out_77[41:24], u_ca_out_76[47:42]};
assign col_out_80 = {u_ca_out_80[5:0],u_ca_out_79[23:6], u_ca_out_78[41:24], u_ca_out_77[47:42]};
assign col_out_81 = {u_ca_out_81[5:0],u_ca_out_80[23:6], u_ca_out_79[41:24], u_ca_out_78[47:42]};
assign col_out_82 = {u_ca_out_82[5:0],u_ca_out_81[23:6], u_ca_out_80[41:24], u_ca_out_79[47:42]};
assign col_out_83 = {u_ca_out_83[5:0],u_ca_out_82[23:6], u_ca_out_81[41:24], u_ca_out_80[47:42]};
assign col_out_84 = {u_ca_out_84[5:0],u_ca_out_83[23:6], u_ca_out_82[41:24], u_ca_out_81[47:42]};
assign col_out_85 = {u_ca_out_85[5:0],u_ca_out_84[23:6], u_ca_out_83[41:24], u_ca_out_82[47:42]};
assign col_out_86 = {u_ca_out_86[5:0],u_ca_out_85[23:6], u_ca_out_84[41:24], u_ca_out_83[47:42]};
assign col_out_87 = {u_ca_out_87[5:0],u_ca_out_86[23:6], u_ca_out_85[41:24], u_ca_out_84[47:42]};
assign col_out_88 = {u_ca_out_88[5:0],u_ca_out_87[23:6], u_ca_out_86[41:24], u_ca_out_85[47:42]};
assign col_out_89 = {u_ca_out_89[5:0],u_ca_out_88[23:6], u_ca_out_87[41:24], u_ca_out_86[47:42]};
assign col_out_90 = {u_ca_out_90[5:0],u_ca_out_89[23:6], u_ca_out_88[41:24], u_ca_out_87[47:42]};
assign col_out_91 = {u_ca_out_91[5:0],u_ca_out_90[23:6], u_ca_out_89[41:24], u_ca_out_88[47:42]};
assign col_out_92 = {u_ca_out_92[5:0],u_ca_out_91[23:6], u_ca_out_90[41:24], u_ca_out_89[47:42]};
assign col_out_93 = {u_ca_out_93[5:0],u_ca_out_92[23:6], u_ca_out_91[41:24], u_ca_out_90[47:42]};
assign col_out_94 = {u_ca_out_94[5:0],u_ca_out_93[23:6], u_ca_out_92[41:24], u_ca_out_91[47:42]};
assign col_out_95 = {u_ca_out_95[5:0],u_ca_out_94[23:6], u_ca_out_93[41:24], u_ca_out_92[47:42]};
assign col_out_96 = {u_ca_out_96[5:0],u_ca_out_95[23:6], u_ca_out_94[41:24], u_ca_out_93[47:42]};
assign col_out_97 = {u_ca_out_97[5:0],u_ca_out_96[23:6], u_ca_out_95[41:24], u_ca_out_94[47:42]};
assign col_out_98 = {u_ca_out_98[5:0],u_ca_out_97[23:6], u_ca_out_96[41:24], u_ca_out_95[47:42]};
assign col_out_99 = {u_ca_out_99[5:0],u_ca_out_98[23:6], u_ca_out_97[41:24], u_ca_out_96[47:42]};
assign col_out_100 = {u_ca_out_100[5:0],u_ca_out_99[23:6], u_ca_out_98[41:24], u_ca_out_97[47:42]};
assign col_out_101 = {u_ca_out_101[5:0],u_ca_out_100[23:6], u_ca_out_99[41:24], u_ca_out_98[47:42]};
assign col_out_102 = {u_ca_out_102[5:0],u_ca_out_101[23:6], u_ca_out_100[41:24], u_ca_out_99[47:42]};
assign col_out_103 = {u_ca_out_103[5:0],u_ca_out_102[23:6], u_ca_out_101[41:24], u_ca_out_100[47:42]};
assign col_out_104 = {u_ca_out_104[5:0],u_ca_out_103[23:6], u_ca_out_102[41:24], u_ca_out_101[47:42]};
assign col_out_105 = {u_ca_out_105[5:0],u_ca_out_104[23:6], u_ca_out_103[41:24], u_ca_out_102[47:42]};
assign col_out_106 = {u_ca_out_106[5:0],u_ca_out_105[23:6], u_ca_out_104[41:24], u_ca_out_103[47:42]};
assign col_out_107 = {u_ca_out_107[5:0],u_ca_out_106[23:6], u_ca_out_105[41:24], u_ca_out_104[47:42]};
assign col_out_108 = {u_ca_out_108[5:0],u_ca_out_107[23:6], u_ca_out_106[41:24], u_ca_out_105[47:42]};
assign col_out_109 = {u_ca_out_109[5:0],u_ca_out_108[23:6], u_ca_out_107[41:24], u_ca_out_106[47:42]};
assign col_out_110 = {u_ca_out_110[5:0],u_ca_out_109[23:6], u_ca_out_108[41:24], u_ca_out_107[47:42]};
assign col_out_111 = {u_ca_out_111[5:0],u_ca_out_110[23:6], u_ca_out_109[41:24], u_ca_out_108[47:42]};
assign col_out_112 = {u_ca_out_112[5:0],u_ca_out_111[23:6], u_ca_out_110[41:24], u_ca_out_109[47:42]};
assign col_out_113 = {u_ca_out_113[5:0],u_ca_out_112[23:6], u_ca_out_111[41:24], u_ca_out_110[47:42]};
assign col_out_114 = {u_ca_out_114[5:0],u_ca_out_113[23:6], u_ca_out_112[41:24], u_ca_out_111[47:42]};
assign col_out_115 = {u_ca_out_115[5:0],u_ca_out_114[23:6], u_ca_out_113[41:24], u_ca_out_112[47:42]};
assign col_out_116 = {u_ca_out_116[5:0],u_ca_out_115[23:6], u_ca_out_114[41:24], u_ca_out_113[47:42]};
assign col_out_117 = {u_ca_out_117[5:0],u_ca_out_116[23:6], u_ca_out_115[41:24], u_ca_out_114[47:42]};
assign col_out_118 = {u_ca_out_118[5:0],u_ca_out_117[23:6], u_ca_out_116[41:24], u_ca_out_115[47:42]};
assign col_out_119 = {u_ca_out_119[5:0],u_ca_out_118[23:6], u_ca_out_117[41:24], u_ca_out_116[47:42]};
assign col_out_120 = {u_ca_out_120[5:0],u_ca_out_119[23:6], u_ca_out_118[41:24], u_ca_out_117[47:42]};
assign col_out_121 = {u_ca_out_121[5:0],u_ca_out_120[23:6], u_ca_out_119[41:24], u_ca_out_118[47:42]};
assign col_out_122 = {u_ca_out_122[5:0],u_ca_out_121[23:6], u_ca_out_120[41:24], u_ca_out_119[47:42]};
assign col_out_123 = {u_ca_out_123[5:0],u_ca_out_122[23:6], u_ca_out_121[41:24], u_ca_out_120[47:42]};
assign col_out_124 = {u_ca_out_124[5:0],u_ca_out_123[23:6], u_ca_out_122[41:24], u_ca_out_121[47:42]};
assign col_out_125 = {u_ca_out_125[5:0],u_ca_out_124[23:6], u_ca_out_123[41:24], u_ca_out_122[47:42]};
assign col_out_126 = {u_ca_out_126[5:0],u_ca_out_125[23:6], u_ca_out_124[41:24], u_ca_out_123[47:42]};
assign col_out_127 = {u_ca_out_127[5:0],u_ca_out_126[23:6], u_ca_out_125[41:24], u_ca_out_124[47:42]};
assign col_out_128 = {u_ca_out_128[5:0],u_ca_out_127[23:6], u_ca_out_126[41:24], u_ca_out_125[47:42]};
assign col_out_129 = {u_ca_out_129[5:0],u_ca_out_128[23:6], u_ca_out_127[41:24], u_ca_out_126[47:42]};
assign col_out_130 = {u_ca_out_130[5:0],u_ca_out_129[23:6], u_ca_out_128[41:24], u_ca_out_127[47:42]};
assign col_out_131 = {u_ca_out_131[5:0],u_ca_out_130[23:6], u_ca_out_129[41:24], u_ca_out_128[47:42]};
assign col_out_132 = {u_ca_out_132[5:0],u_ca_out_131[23:6], u_ca_out_130[41:24], u_ca_out_129[47:42]};
assign col_out_133 = {u_ca_out_133[5:0],u_ca_out_132[23:6], u_ca_out_131[41:24], u_ca_out_130[47:42]};
assign col_out_134 = {u_ca_out_134[5:0],u_ca_out_133[23:6], u_ca_out_132[41:24], u_ca_out_131[47:42]};
assign col_out_135 = {u_ca_out_135[5:0],u_ca_out_134[23:6], u_ca_out_133[41:24], u_ca_out_132[47:42]};
assign col_out_136 = {u_ca_out_136[5:0],u_ca_out_135[23:6], u_ca_out_134[41:24], u_ca_out_133[47:42]};
assign col_out_137 = {u_ca_out_137[5:0],u_ca_out_136[23:6], u_ca_out_135[41:24], u_ca_out_134[47:42]};
assign col_out_138 = {u_ca_out_138[5:0],u_ca_out_137[23:6], u_ca_out_136[41:24], u_ca_out_135[47:42]};
assign col_out_139 = {u_ca_out_139[5:0],u_ca_out_138[23:6], u_ca_out_137[41:24], u_ca_out_136[47:42]};
assign col_out_140 = {u_ca_out_140[5:0],u_ca_out_139[23:6], u_ca_out_138[41:24], u_ca_out_137[47:42]};
assign col_out_141 = {u_ca_out_141[5:0],u_ca_out_140[23:6], u_ca_out_139[41:24], u_ca_out_138[47:42]};
assign col_out_142 = {u_ca_out_142[5:0],u_ca_out_141[23:6], u_ca_out_140[41:24], u_ca_out_139[47:42]};
assign col_out_143 = {u_ca_out_143[5:0],u_ca_out_142[23:6], u_ca_out_141[41:24], u_ca_out_140[47:42]};
assign col_out_144 = {u_ca_out_144[5:0],u_ca_out_143[23:6], u_ca_out_142[41:24], u_ca_out_141[47:42]};
assign col_out_145 = {u_ca_out_145[5:0],u_ca_out_144[23:6], u_ca_out_143[41:24], u_ca_out_142[47:42]};
assign col_out_146 = {u_ca_out_146[5:0],u_ca_out_145[23:6], u_ca_out_144[41:24], u_ca_out_143[47:42]};
assign col_out_147 = {u_ca_out_147[5:0],u_ca_out_146[23:6], u_ca_out_145[41:24], u_ca_out_144[47:42]};
assign col_out_148 = {u_ca_out_148[5:0],u_ca_out_147[23:6], u_ca_out_146[41:24], u_ca_out_145[47:42]};
assign col_out_149 = {u_ca_out_149[5:0],u_ca_out_148[23:6], u_ca_out_147[41:24], u_ca_out_146[47:42]};
assign col_out_150 = {u_ca_out_150[5:0],u_ca_out_149[23:6], u_ca_out_148[41:24], u_ca_out_147[47:42]};
assign col_out_151 = {u_ca_out_151[5:0],u_ca_out_150[23:6], u_ca_out_149[41:24], u_ca_out_148[47:42]};
assign col_out_152 = {u_ca_out_152[5:0],u_ca_out_151[23:6], u_ca_out_150[41:24], u_ca_out_149[47:42]};
assign col_out_153 = {u_ca_out_153[5:0],u_ca_out_152[23:6], u_ca_out_151[41:24], u_ca_out_150[47:42]};
assign col_out_154 = {u_ca_out_154[5:0],u_ca_out_153[23:6], u_ca_out_152[41:24], u_ca_out_151[47:42]};
assign col_out_155 = {u_ca_out_155[5:0],u_ca_out_154[23:6], u_ca_out_153[41:24], u_ca_out_152[47:42]};
assign col_out_156 = {u_ca_out_156[5:0],u_ca_out_155[23:6], u_ca_out_154[41:24], u_ca_out_153[47:42]};
assign col_out_157 = {u_ca_out_157[5:0],u_ca_out_156[23:6], u_ca_out_155[41:24], u_ca_out_154[47:42]};
assign col_out_158 = {u_ca_out_158[5:0],u_ca_out_157[23:6], u_ca_out_156[41:24], u_ca_out_155[47:42]};
assign col_out_159 = {u_ca_out_159[5:0],u_ca_out_158[23:6], u_ca_out_157[41:24], u_ca_out_156[47:42]};
assign col_out_160 = {u_ca_out_160[5:0],u_ca_out_159[23:6], u_ca_out_158[41:24], u_ca_out_157[47:42]};
assign col_out_161 = {u_ca_out_161[5:0],u_ca_out_160[23:6], u_ca_out_159[41:24], u_ca_out_158[47:42]};
assign col_out_162 = {u_ca_out_162[5:0],u_ca_out_161[23:6], u_ca_out_160[41:24], u_ca_out_159[47:42]};
assign col_out_163 = {u_ca_out_163[5:0],u_ca_out_162[23:6], u_ca_out_161[41:24], u_ca_out_160[47:42]};
assign col_out_164 = {u_ca_out_164[5:0],u_ca_out_163[23:6], u_ca_out_162[41:24], u_ca_out_161[47:42]};
assign col_out_165 = {u_ca_out_165[5:0],u_ca_out_164[23:6], u_ca_out_163[41:24], u_ca_out_162[47:42]};
assign col_out_166 = {u_ca_out_166[5:0],u_ca_out_165[23:6], u_ca_out_164[41:24], u_ca_out_163[47:42]};
assign col_out_167 = {u_ca_out_167[5:0],u_ca_out_166[23:6], u_ca_out_165[41:24], u_ca_out_164[47:42]};
assign col_out_168 = {u_ca_out_168[5:0],u_ca_out_167[23:6], u_ca_out_166[41:24], u_ca_out_165[47:42]};
assign col_out_169 = {u_ca_out_169[5:0],u_ca_out_168[23:6], u_ca_out_167[41:24], u_ca_out_166[47:42]};
assign col_out_170 = {u_ca_out_170[5:0],u_ca_out_169[23:6], u_ca_out_168[41:24], u_ca_out_167[47:42]};
assign col_out_171 = {u_ca_out_171[5:0],u_ca_out_170[23:6], u_ca_out_169[41:24], u_ca_out_168[47:42]};
assign col_out_172 = {u_ca_out_172[5:0],u_ca_out_171[23:6], u_ca_out_170[41:24], u_ca_out_169[47:42]};
assign col_out_173 = {u_ca_out_173[5:0],u_ca_out_172[23:6], u_ca_out_171[41:24], u_ca_out_170[47:42]};
assign col_out_174 = {u_ca_out_174[5:0],u_ca_out_173[23:6], u_ca_out_172[41:24], u_ca_out_171[47:42]};
assign col_out_175 = {u_ca_out_175[5:0],u_ca_out_174[23:6], u_ca_out_173[41:24], u_ca_out_172[47:42]};
assign col_out_176 = {u_ca_out_176[5:0],u_ca_out_175[23:6], u_ca_out_174[41:24], u_ca_out_173[47:42]};
assign col_out_177 = {u_ca_out_177[5:0],u_ca_out_176[23:6], u_ca_out_175[41:24], u_ca_out_174[47:42]};
assign col_out_178 = {u_ca_out_178[5:0],u_ca_out_177[23:6], u_ca_out_176[41:24], u_ca_out_175[47:42]};
assign col_out_179 = {u_ca_out_179[5:0],u_ca_out_178[23:6], u_ca_out_177[41:24], u_ca_out_176[47:42]};
assign col_out_180 = {u_ca_out_180[5:0],u_ca_out_179[23:6], u_ca_out_178[41:24], u_ca_out_177[47:42]};
assign col_out_181 = {u_ca_out_181[5:0],u_ca_out_180[23:6], u_ca_out_179[41:24], u_ca_out_178[47:42]};
assign col_out_182 = {u_ca_out_182[5:0],u_ca_out_181[23:6], u_ca_out_180[41:24], u_ca_out_179[47:42]};
assign col_out_183 = {u_ca_out_183[5:0],u_ca_out_182[23:6], u_ca_out_181[41:24], u_ca_out_180[47:42]};
assign col_out_184 = {u_ca_out_184[5:0],u_ca_out_183[23:6], u_ca_out_182[41:24], u_ca_out_181[47:42]};
assign col_out_185 = {u_ca_out_185[5:0],u_ca_out_184[23:6], u_ca_out_183[41:24], u_ca_out_182[47:42]};
assign col_out_186 = {u_ca_out_186[5:0],u_ca_out_185[23:6], u_ca_out_184[41:24], u_ca_out_183[47:42]};
assign col_out_187 = {u_ca_out_187[5:0],u_ca_out_186[23:6], u_ca_out_185[41:24], u_ca_out_184[47:42]};
assign col_out_188 = {u_ca_out_188[5:0],u_ca_out_187[23:6], u_ca_out_186[41:24], u_ca_out_185[47:42]};
assign col_out_189 = {u_ca_out_189[5:0],u_ca_out_188[23:6], u_ca_out_187[41:24], u_ca_out_186[47:42]};
assign col_out_190 = {u_ca_out_190[5:0],u_ca_out_189[23:6], u_ca_out_188[41:24], u_ca_out_187[47:42]};
assign col_out_191 = {u_ca_out_191[5:0],u_ca_out_190[23:6], u_ca_out_189[41:24], u_ca_out_188[47:42]};
assign col_out_192 = {u_ca_out_192[5:0],u_ca_out_191[23:6], u_ca_out_190[41:24], u_ca_out_189[47:42]};
assign col_out_193 = {u_ca_out_193[5:0],u_ca_out_192[23:6], u_ca_out_191[41:24], u_ca_out_190[47:42]};
assign col_out_194 = {u_ca_out_194[5:0],u_ca_out_193[23:6], u_ca_out_192[41:24], u_ca_out_191[47:42]};
assign col_out_195 = {u_ca_out_195[5:0],u_ca_out_194[23:6], u_ca_out_193[41:24], u_ca_out_192[47:42]};
assign col_out_196 = {u_ca_out_196[5:0],u_ca_out_195[23:6], u_ca_out_194[41:24], u_ca_out_193[47:42]};
assign col_out_197 = {u_ca_out_197[5:0],u_ca_out_196[23:6], u_ca_out_195[41:24], u_ca_out_194[47:42]};
assign col_out_198 = {u_ca_out_198[5:0],u_ca_out_197[23:6], u_ca_out_196[41:24], u_ca_out_195[47:42]};
assign col_out_199 = {u_ca_out_199[5:0],u_ca_out_198[23:6], u_ca_out_197[41:24], u_ca_out_196[47:42]};
assign col_out_200 = {u_ca_out_200[5:0],u_ca_out_199[23:6], u_ca_out_198[41:24], u_ca_out_197[47:42]};
assign col_out_201 = {u_ca_out_201[5:0],u_ca_out_200[23:6], u_ca_out_199[41:24], u_ca_out_198[47:42]};
assign col_out_202 = {u_ca_out_202[5:0],u_ca_out_201[23:6], u_ca_out_200[41:24], u_ca_out_199[47:42]};
assign col_out_203 = {u_ca_out_203[5:0],u_ca_out_202[23:6], u_ca_out_201[41:24], u_ca_out_200[47:42]};
assign col_out_204 = {u_ca_out_204[5:0],u_ca_out_203[23:6], u_ca_out_202[41:24], u_ca_out_201[47:42]};
assign col_out_205 = {u_ca_out_205[5:0],u_ca_out_204[23:6], u_ca_out_203[41:24], u_ca_out_202[47:42]};
assign col_out_206 = {u_ca_out_206[5:0],u_ca_out_205[23:6], u_ca_out_204[41:24], u_ca_out_203[47:42]};
assign col_out_207 = {u_ca_out_207[5:0],u_ca_out_206[23:6], u_ca_out_205[41:24], u_ca_out_204[47:42]};
assign col_out_208 = {u_ca_out_208[5:0],u_ca_out_207[23:6], u_ca_out_206[41:24], u_ca_out_205[47:42]};
assign col_out_209 = {u_ca_out_209[5:0],u_ca_out_208[23:6], u_ca_out_207[41:24], u_ca_out_206[47:42]};
assign col_out_210 = {u_ca_out_210[5:0],u_ca_out_209[23:6], u_ca_out_208[41:24], u_ca_out_207[47:42]};
assign col_out_211 = {u_ca_out_211[5:0],u_ca_out_210[23:6], u_ca_out_209[41:24], u_ca_out_208[47:42]};
assign col_out_212 = {u_ca_out_212[5:0],u_ca_out_211[23:6], u_ca_out_210[41:24], u_ca_out_209[47:42]};
assign col_out_213 = {u_ca_out_213[5:0],u_ca_out_212[23:6], u_ca_out_211[41:24], u_ca_out_210[47:42]};
assign col_out_214 = {u_ca_out_214[5:0],u_ca_out_213[23:6], u_ca_out_212[41:24], u_ca_out_211[47:42]};
assign col_out_215 = {u_ca_out_215[5:0],u_ca_out_214[23:6], u_ca_out_213[41:24], u_ca_out_212[47:42]};
assign col_out_216 = {u_ca_out_216[5:0],u_ca_out_215[23:6], u_ca_out_214[41:24], u_ca_out_213[47:42]};
assign col_out_217 = {u_ca_out_217[5:0],u_ca_out_216[23:6], u_ca_out_215[41:24], u_ca_out_214[47:42]};
assign col_out_218 = {u_ca_out_218[5:0],u_ca_out_217[23:6], u_ca_out_216[41:24], u_ca_out_215[47:42]};
assign col_out_219 = {u_ca_out_219[5:0],u_ca_out_218[23:6], u_ca_out_217[41:24], u_ca_out_216[47:42]};
assign col_out_220 = {u_ca_out_220[5:0],u_ca_out_219[23:6], u_ca_out_218[41:24], u_ca_out_217[47:42]};
assign col_out_221 = {u_ca_out_221[5:0],u_ca_out_220[23:6], u_ca_out_219[41:24], u_ca_out_218[47:42]};
assign col_out_222 = {u_ca_out_222[5:0],u_ca_out_221[23:6], u_ca_out_220[41:24], u_ca_out_219[47:42]};
assign col_out_223 = {u_ca_out_223[5:0],u_ca_out_222[23:6], u_ca_out_221[41:24], u_ca_out_220[47:42]};
assign col_out_224 = {u_ca_out_224[5:0],u_ca_out_223[23:6], u_ca_out_222[41:24], u_ca_out_221[47:42]};
assign col_out_225 = {u_ca_out_225[5:0],u_ca_out_224[23:6], u_ca_out_223[41:24], u_ca_out_222[47:42]};
assign col_out_226 = {u_ca_out_226[5:0],u_ca_out_225[23:6], u_ca_out_224[41:24], u_ca_out_223[47:42]};
assign col_out_227 = {u_ca_out_227[5:0],u_ca_out_226[23:6], u_ca_out_225[41:24], u_ca_out_224[47:42]};
assign col_out_228 = {u_ca_out_228[5:0],u_ca_out_227[23:6], u_ca_out_226[41:24], u_ca_out_225[47:42]};
assign col_out_229 = {u_ca_out_229[5:0],u_ca_out_228[23:6], u_ca_out_227[41:24], u_ca_out_226[47:42]};
assign col_out_230 = {u_ca_out_230[5:0],u_ca_out_229[23:6], u_ca_out_228[41:24], u_ca_out_227[47:42]};
assign col_out_231 = {u_ca_out_231[5:0],u_ca_out_230[23:6], u_ca_out_229[41:24], u_ca_out_228[47:42]};
assign col_out_232 = {u_ca_out_232[5:0],u_ca_out_231[23:6], u_ca_out_230[41:24], u_ca_out_229[47:42]};
assign col_out_233 = {u_ca_out_233[5:0],u_ca_out_232[23:6], u_ca_out_231[41:24], u_ca_out_230[47:42]};
assign col_out_234 = {u_ca_out_234[5:0],u_ca_out_233[23:6], u_ca_out_232[41:24], u_ca_out_231[47:42]};
assign col_out_235 = {u_ca_out_235[5:0],u_ca_out_234[23:6], u_ca_out_233[41:24], u_ca_out_232[47:42]};
assign col_out_236 = {u_ca_out_236[5:0],u_ca_out_235[23:6], u_ca_out_234[41:24], u_ca_out_233[47:42]};
assign col_out_237 = {u_ca_out_237[5:0],u_ca_out_236[23:6], u_ca_out_235[41:24], u_ca_out_234[47:42]};
assign col_out_238 = {u_ca_out_238[5:0],u_ca_out_237[23:6], u_ca_out_236[41:24], u_ca_out_235[47:42]};
assign col_out_239 = {u_ca_out_239[5:0],u_ca_out_238[23:6], u_ca_out_237[41:24], u_ca_out_236[47:42]};
assign col_out_240 = {u_ca_out_240[5:0],u_ca_out_239[23:6], u_ca_out_238[41:24], u_ca_out_237[47:42]};
assign col_out_241 = {u_ca_out_241[5:0],u_ca_out_240[23:6], u_ca_out_239[41:24], u_ca_out_238[47:42]};
assign col_out_242 = {u_ca_out_242[5:0],u_ca_out_241[23:6], u_ca_out_240[41:24], u_ca_out_239[47:42]};
assign col_out_243 = {u_ca_out_243[5:0],u_ca_out_242[23:6], u_ca_out_241[41:24], u_ca_out_240[47:42]};
assign col_out_244 = {u_ca_out_244[5:0],u_ca_out_243[23:6], u_ca_out_242[41:24], u_ca_out_241[47:42]};
assign col_out_245 = {u_ca_out_245[5:0],u_ca_out_244[23:6], u_ca_out_243[41:24], u_ca_out_242[47:42]};
assign col_out_246 = {u_ca_out_246[5:0],u_ca_out_245[23:6], u_ca_out_244[41:24], u_ca_out_243[47:42]};
assign col_out_247 = {u_ca_out_247[5:0],u_ca_out_246[23:6], u_ca_out_245[41:24], u_ca_out_244[47:42]};
assign col_out_248 = {u_ca_out_248[5:0],u_ca_out_247[23:6], u_ca_out_246[41:24], u_ca_out_245[47:42]};
assign col_out_249 = {u_ca_out_249[5:0],u_ca_out_248[23:6], u_ca_out_247[41:24], u_ca_out_246[47:42]};
assign col_out_250 = {u_ca_out_250[5:0],u_ca_out_249[23:6], u_ca_out_248[41:24], u_ca_out_247[47:42]};
assign col_out_251 = {u_ca_out_251[5:0],u_ca_out_250[23:6], u_ca_out_249[41:24], u_ca_out_248[47:42]};
assign col_out_252 = {u_ca_out_252[5:0],u_ca_out_251[23:6], u_ca_out_250[41:24], u_ca_out_249[47:42]};
assign col_out_253 = {u_ca_out_253[5:0],u_ca_out_252[23:6], u_ca_out_251[41:24], u_ca_out_250[47:42]};
assign col_out_254 = {u_ca_out_254[5:0],u_ca_out_253[23:6], u_ca_out_252[41:24], u_ca_out_251[47:42]};
assign col_out_255 = {u_ca_out_255[5:0],u_ca_out_254[23:6], u_ca_out_253[41:24], u_ca_out_252[47:42]};
assign col_out_256 = {u_ca_out_256[5:0],u_ca_out_255[23:6], u_ca_out_254[41:24], u_ca_out_253[47:42]};
assign col_out_257 = {u_ca_out_257[5:0],u_ca_out_256[23:6], u_ca_out_255[41:24], u_ca_out_254[47:42]};
assign col_out_258 = {u_ca_out_258[5:0],u_ca_out_257[23:6], u_ca_out_256[41:24], u_ca_out_255[47:42]};
assign col_out_259 = {u_ca_out_259[5:0],u_ca_out_258[23:6], u_ca_out_257[41:24], u_ca_out_256[47:42]};
assign col_out_260 = {u_ca_out_260[5:0],u_ca_out_259[23:6], u_ca_out_258[41:24], u_ca_out_257[47:42]};
assign col_out_261 = {u_ca_out_261[5:0],u_ca_out_260[23:6], u_ca_out_259[41:24], u_ca_out_258[47:42]};
assign col_out_262 = {u_ca_out_262[5:0],u_ca_out_261[23:6], u_ca_out_260[41:24], u_ca_out_259[47:42]};
assign col_out_263 = {u_ca_out_263[5:0],u_ca_out_262[23:6], u_ca_out_261[41:24], u_ca_out_260[47:42]};
assign col_out_264 = {u_ca_out_264[5:0],u_ca_out_263[23:6], u_ca_out_262[41:24], u_ca_out_261[47:42]};
assign col_out_265 = {u_ca_out_265[5:0],u_ca_out_264[23:6], u_ca_out_263[41:24], u_ca_out_262[47:42]};
assign col_out_266 = {u_ca_out_266[5:0],u_ca_out_265[23:6], u_ca_out_264[41:24], u_ca_out_263[47:42]};
assign col_out_267 = {u_ca_out_267[5:0],u_ca_out_266[23:6], u_ca_out_265[41:24], u_ca_out_264[47:42]};
assign col_out_268 = {u_ca_out_268[5:0],u_ca_out_267[23:6], u_ca_out_266[41:24], u_ca_out_265[47:42]};
assign col_out_269 = {u_ca_out_269[5:0],u_ca_out_268[23:6], u_ca_out_267[41:24], u_ca_out_266[47:42]};
assign col_out_270 = {u_ca_out_270[5:0],u_ca_out_269[23:6], u_ca_out_268[41:24], u_ca_out_267[47:42]};
assign col_out_271 = {u_ca_out_271[5:0],u_ca_out_270[23:6], u_ca_out_269[41:24], u_ca_out_268[47:42]};
assign col_out_272 = {u_ca_out_272[5:0],u_ca_out_271[23:6], u_ca_out_270[41:24], u_ca_out_269[47:42]};
assign col_out_273 = {u_ca_out_273[5:0],u_ca_out_272[23:6], u_ca_out_271[41:24], u_ca_out_270[47:42]};
assign col_out_274 = {u_ca_out_274[5:0],u_ca_out_273[23:6], u_ca_out_272[41:24], u_ca_out_271[47:42]};
assign col_out_275 = {u_ca_out_275[5:0],u_ca_out_274[23:6], u_ca_out_273[41:24], u_ca_out_272[47:42]};
assign col_out_276 = {u_ca_out_276[5:0],u_ca_out_275[23:6], u_ca_out_274[41:24], u_ca_out_273[47:42]};
assign col_out_277 = {u_ca_out_277[5:0],u_ca_out_276[23:6], u_ca_out_275[41:24], u_ca_out_274[47:42]};
assign col_out_278 = {u_ca_out_278[5:0],u_ca_out_277[23:6], u_ca_out_276[41:24], u_ca_out_275[47:42]};
assign col_out_279 = {u_ca_out_279[5:0],u_ca_out_278[23:6], u_ca_out_277[41:24], u_ca_out_276[47:42]};
assign col_out_280 = {u_ca_out_280[5:0],u_ca_out_279[23:6], u_ca_out_278[41:24], u_ca_out_277[47:42]};
assign col_out_281 = {u_ca_out_281[5:0],u_ca_out_280[23:6], u_ca_out_279[41:24], u_ca_out_278[47:42]};
assign col_out_282 = {u_ca_out_282[5:0],u_ca_out_281[23:6], u_ca_out_280[41:24], u_ca_out_279[47:42]};
assign col_out_283 = {u_ca_out_283[5:0],u_ca_out_282[23:6], u_ca_out_281[41:24], u_ca_out_280[47:42]};
assign col_out_284 = {u_ca_out_284[5:0],u_ca_out_283[23:6], u_ca_out_282[41:24], u_ca_out_281[47:42]};
assign col_out_285 = {u_ca_out_285[5:0],u_ca_out_284[23:6], u_ca_out_283[41:24], u_ca_out_282[47:42]};
assign col_out_286 = {u_ca_out_286[5:0],u_ca_out_285[23:6], u_ca_out_284[41:24], u_ca_out_283[47:42]};
assign col_out_287 = {u_ca_out_287[5:0],u_ca_out_286[23:6], u_ca_out_285[41:24], u_ca_out_284[47:42]};
assign col_out_288 = {u_ca_out_288[5:0],u_ca_out_287[23:6], u_ca_out_286[41:24], u_ca_out_285[47:42]};
assign col_out_289 = {u_ca_out_289[5:0],u_ca_out_288[23:6], u_ca_out_287[41:24], u_ca_out_286[47:42]};
assign col_out_290 = {u_ca_out_290[5:0],u_ca_out_289[23:6], u_ca_out_288[41:24], u_ca_out_287[47:42]};
assign col_out_291 = {u_ca_out_291[5:0],u_ca_out_290[23:6], u_ca_out_289[41:24], u_ca_out_288[47:42]};
assign col_out_292 = {u_ca_out_292[5:0],u_ca_out_291[23:6], u_ca_out_290[41:24], u_ca_out_289[47:42]};
assign col_out_293 = {u_ca_out_293[5:0],u_ca_out_292[23:6], u_ca_out_291[41:24], u_ca_out_290[47:42]};
assign col_out_294 = {u_ca_out_294[5:0],u_ca_out_293[23:6], u_ca_out_292[41:24], u_ca_out_291[47:42]};
assign col_out_295 = {u_ca_out_295[5:0],u_ca_out_294[23:6], u_ca_out_293[41:24], u_ca_out_292[47:42]};
assign col_out_296 = {u_ca_out_296[5:0],u_ca_out_295[23:6], u_ca_out_294[41:24], u_ca_out_293[47:42]};
assign col_out_297 = {u_ca_out_297[5:0],u_ca_out_296[23:6], u_ca_out_295[41:24], u_ca_out_294[47:42]};
assign col_out_298 = {u_ca_out_298[5:0],u_ca_out_297[23:6], u_ca_out_296[41:24], u_ca_out_295[47:42]};
assign col_out_299 = {u_ca_out_299[5:0],u_ca_out_298[23:6], u_ca_out_297[41:24], u_ca_out_296[47:42]};
assign col_out_300 = {u_ca_out_300[5:0],u_ca_out_299[23:6], u_ca_out_298[41:24], u_ca_out_297[47:42]};
assign col_out_301 = {u_ca_out_301[5:0],u_ca_out_300[23:6], u_ca_out_299[41:24], u_ca_out_298[47:42]};
assign col_out_302 = {u_ca_out_302[5:0],u_ca_out_301[23:6], u_ca_out_300[41:24], u_ca_out_299[47:42]};
assign col_out_303 = {u_ca_out_303[5:0],u_ca_out_302[23:6], u_ca_out_301[41:24], u_ca_out_300[47:42]};
assign col_out_304 = {u_ca_out_304[5:0],u_ca_out_303[23:6], u_ca_out_302[41:24], u_ca_out_301[47:42]};
assign col_out_305 = {u_ca_out_305[5:0],u_ca_out_304[23:6], u_ca_out_303[41:24], u_ca_out_302[47:42]};
assign col_out_306 = {u_ca_out_306[5:0],u_ca_out_305[23:6], u_ca_out_304[41:24], u_ca_out_303[47:42]};
assign col_out_307 = {u_ca_out_307[5:0],u_ca_out_306[23:6], u_ca_out_305[41:24], u_ca_out_304[47:42]};
assign col_out_308 = {u_ca_out_308[5:0],u_ca_out_307[23:6], u_ca_out_306[41:24], u_ca_out_305[47:42]};
assign col_out_309 = {u_ca_out_309[5:0],u_ca_out_308[23:6], u_ca_out_307[41:24], u_ca_out_306[47:42]};
assign col_out_310 = {u_ca_out_310[5:0],u_ca_out_309[23:6], u_ca_out_308[41:24], u_ca_out_307[47:42]};
assign col_out_311 = {u_ca_out_311[5:0],u_ca_out_310[23:6], u_ca_out_309[41:24], u_ca_out_308[47:42]};
assign col_out_312 = {u_ca_out_312[5:0],u_ca_out_311[23:6], u_ca_out_310[41:24], u_ca_out_309[47:42]};
assign col_out_313 = {u_ca_out_313[5:0],u_ca_out_312[23:6], u_ca_out_311[41:24], u_ca_out_310[47:42]};
assign col_out_314 = {u_ca_out_314[5:0],u_ca_out_313[23:6], u_ca_out_312[41:24], u_ca_out_311[47:42]};
assign col_out_315 = {u_ca_out_315[5:0],u_ca_out_314[23:6], u_ca_out_313[41:24], u_ca_out_312[47:42]};
assign col_out_316 = {u_ca_out_316[5:0],u_ca_out_315[23:6], u_ca_out_314[41:24], u_ca_out_313[47:42]};
assign col_out_317 = {u_ca_out_317[5:0],u_ca_out_316[23:6], u_ca_out_315[41:24], u_ca_out_314[47:42]};
assign col_out_318 = {u_ca_out_318[5:0],u_ca_out_317[23:6], u_ca_out_316[41:24], u_ca_out_315[47:42]};
assign col_out_319 = {u_ca_out_319[5:0],u_ca_out_318[23:6], u_ca_out_317[41:24], u_ca_out_316[47:42]};
assign col_out_320 = {u_ca_out_320[5:0],u_ca_out_319[23:6], u_ca_out_318[41:24], u_ca_out_317[47:42]};
assign col_out_321 = {u_ca_out_321[5:0],u_ca_out_320[23:6], u_ca_out_319[41:24], u_ca_out_318[47:42]};
assign col_out_322 = {u_ca_out_322[5:0],u_ca_out_321[23:6], u_ca_out_320[41:24], u_ca_out_319[47:42]};
assign col_out_323 = {u_ca_out_323[5:0],u_ca_out_322[23:6], u_ca_out_321[41:24], u_ca_out_320[47:42]};
assign col_out_324 = {u_ca_out_324[5:0],u_ca_out_323[23:6], u_ca_out_322[41:24], u_ca_out_321[47:42]};
assign col_out_325 = {u_ca_out_325[5:0],u_ca_out_324[23:6], u_ca_out_323[41:24], u_ca_out_322[47:42]};
assign col_out_326 = {u_ca_out_326[5:0],u_ca_out_325[23:6], u_ca_out_324[41:24], u_ca_out_323[47:42]};
assign col_out_327 = {u_ca_out_327[5:0],u_ca_out_326[23:6], u_ca_out_325[41:24], u_ca_out_324[47:42]};
assign col_out_328 = {u_ca_out_328[5:0],u_ca_out_327[23:6], u_ca_out_326[41:24], u_ca_out_325[47:42]};
assign col_out_329 = {u_ca_out_329[5:0],u_ca_out_328[23:6], u_ca_out_327[41:24], u_ca_out_326[47:42]};
assign col_out_330 = {u_ca_out_330[5:0],u_ca_out_329[23:6], u_ca_out_328[41:24], u_ca_out_327[47:42]};
assign col_out_331 = {u_ca_out_331[5:0],u_ca_out_330[23:6], u_ca_out_329[41:24], u_ca_out_328[47:42]};
assign col_out_332 = {u_ca_out_332[5:0],u_ca_out_331[23:6], u_ca_out_330[41:24], u_ca_out_329[47:42]};
assign col_out_333 = {u_ca_out_333[5:0],u_ca_out_332[23:6], u_ca_out_331[41:24], u_ca_out_330[47:42]};
assign col_out_334 = {u_ca_out_334[5:0],u_ca_out_333[23:6], u_ca_out_332[41:24], u_ca_out_331[47:42]};
assign col_out_335 = {u_ca_out_335[5:0],u_ca_out_334[23:6], u_ca_out_333[41:24], u_ca_out_332[47:42]};
assign col_out_336 = {u_ca_out_336[5:0],u_ca_out_335[23:6], u_ca_out_334[41:24], u_ca_out_333[47:42]};
assign col_out_337 = {u_ca_out_337[5:0],u_ca_out_336[23:6], u_ca_out_335[41:24], u_ca_out_334[47:42]};
assign col_out_338 = {u_ca_out_338[5:0],u_ca_out_337[23:6], u_ca_out_336[41:24], u_ca_out_335[47:42]};
assign col_out_339 = {u_ca_out_339[5:0],u_ca_out_338[23:6], u_ca_out_337[41:24], u_ca_out_336[47:42]};
assign col_out_340 = {u_ca_out_340[5:0],u_ca_out_339[23:6], u_ca_out_338[41:24], u_ca_out_337[47:42]};
assign col_out_341 = {u_ca_out_341[5:0],u_ca_out_340[23:6], u_ca_out_339[41:24], u_ca_out_338[47:42]};
assign col_out_342 = {u_ca_out_342[5:0],u_ca_out_341[23:6], u_ca_out_340[41:24], u_ca_out_339[47:42]};
assign col_out_343 = {u_ca_out_343[5:0],u_ca_out_342[23:6], u_ca_out_341[41:24], u_ca_out_340[47:42]};
assign col_out_344 = {u_ca_out_344[5:0],u_ca_out_343[23:6], u_ca_out_342[41:24], u_ca_out_341[47:42]};
assign col_out_345 = {u_ca_out_345[5:0],u_ca_out_344[23:6], u_ca_out_343[41:24], u_ca_out_342[47:42]};
assign col_out_346 = {u_ca_out_346[5:0],u_ca_out_345[23:6], u_ca_out_344[41:24], u_ca_out_343[47:42]};
assign col_out_347 = {u_ca_out_347[5:0],u_ca_out_346[23:6], u_ca_out_345[41:24], u_ca_out_344[47:42]};
assign col_out_348 = {u_ca_out_348[5:0],u_ca_out_347[23:6], u_ca_out_346[41:24], u_ca_out_345[47:42]};
assign col_out_349 = {u_ca_out_349[5:0],u_ca_out_348[23:6], u_ca_out_347[41:24], u_ca_out_346[47:42]};
assign col_out_350 = {u_ca_out_350[5:0],u_ca_out_349[23:6], u_ca_out_348[41:24], u_ca_out_347[47:42]};
assign col_out_351 = {u_ca_out_351[5:0],u_ca_out_350[23:6], u_ca_out_349[41:24], u_ca_out_348[47:42]};
assign col_out_352 = {u_ca_out_352[5:0],u_ca_out_351[23:6], u_ca_out_350[41:24], u_ca_out_349[47:42]};
assign col_out_353 = {u_ca_out_353[5:0],u_ca_out_352[23:6], u_ca_out_351[41:24], u_ca_out_350[47:42]};
assign col_out_354 = {u_ca_out_354[5:0],u_ca_out_353[23:6], u_ca_out_352[41:24], u_ca_out_351[47:42]};
assign col_out_355 = {u_ca_out_355[5:0],u_ca_out_354[23:6], u_ca_out_353[41:24], u_ca_out_352[47:42]};
assign col_out_356 = {u_ca_out_356[5:0],u_ca_out_355[23:6], u_ca_out_354[41:24], u_ca_out_353[47:42]};
assign col_out_357 = {u_ca_out_357[5:0],u_ca_out_356[23:6], u_ca_out_355[41:24], u_ca_out_354[47:42]};
assign col_out_358 = {u_ca_out_358[5:0],u_ca_out_357[23:6], u_ca_out_356[41:24], u_ca_out_355[47:42]};
assign col_out_359 = {u_ca_out_359[5:0],u_ca_out_358[23:6], u_ca_out_357[41:24], u_ca_out_356[47:42]};
assign col_out_360 = {u_ca_out_360[5:0],u_ca_out_359[23:6], u_ca_out_358[41:24], u_ca_out_357[47:42]};
assign col_out_361 = {u_ca_out_361[5:0],u_ca_out_360[23:6], u_ca_out_359[41:24], u_ca_out_358[47:42]};
assign col_out_362 = {u_ca_out_362[5:0],u_ca_out_361[23:6], u_ca_out_360[41:24], u_ca_out_359[47:42]};
assign col_out_363 = {u_ca_out_363[5:0],u_ca_out_362[23:6], u_ca_out_361[41:24], u_ca_out_360[47:42]};
assign col_out_364 = {u_ca_out_364[5:0],u_ca_out_363[23:6], u_ca_out_362[41:24], u_ca_out_361[47:42]};
assign col_out_365 = {u_ca_out_365[5:0],u_ca_out_364[23:6], u_ca_out_363[41:24], u_ca_out_362[47:42]};
assign col_out_366 = {u_ca_out_366[5:0],u_ca_out_365[23:6], u_ca_out_364[41:24], u_ca_out_363[47:42]};
assign col_out_367 = {u_ca_out_367[5:0],u_ca_out_366[23:6], u_ca_out_365[41:24], u_ca_out_364[47:42]};
assign col_out_368 = {u_ca_out_368[5:0],u_ca_out_367[23:6], u_ca_out_366[41:24], u_ca_out_365[47:42]};
assign col_out_369 = {u_ca_out_369[5:0],u_ca_out_368[23:6], u_ca_out_367[41:24], u_ca_out_366[47:42]};
assign col_out_370 = {u_ca_out_370[5:0],u_ca_out_369[23:6], u_ca_out_368[41:24], u_ca_out_367[47:42]};
assign col_out_371 = {u_ca_out_371[5:0],u_ca_out_370[23:6], u_ca_out_369[41:24], u_ca_out_368[47:42]};
assign col_out_372 = {u_ca_out_372[5:0],u_ca_out_371[23:6], u_ca_out_370[41:24], u_ca_out_369[47:42]};
assign col_out_373 = {u_ca_out_373[5:0],u_ca_out_372[23:6], u_ca_out_371[41:24], u_ca_out_370[47:42]};
assign col_out_374 = {u_ca_out_374[5:0],u_ca_out_373[23:6], u_ca_out_372[41:24], u_ca_out_371[47:42]};
assign col_out_375 = {u_ca_out_375[5:0],u_ca_out_374[23:6], u_ca_out_373[41:24], u_ca_out_372[47:42]};
assign col_out_376 = {u_ca_out_376[5:0],u_ca_out_375[23:6], u_ca_out_374[41:24], u_ca_out_373[47:42]};
assign col_out_377 = {u_ca_out_377[5:0],u_ca_out_376[23:6], u_ca_out_375[41:24], u_ca_out_374[47:42]};
assign col_out_378 = {u_ca_out_378[5:0],u_ca_out_377[23:6], u_ca_out_376[41:24], u_ca_out_375[47:42]};
assign col_out_379 = {u_ca_out_379[5:0],u_ca_out_378[23:6], u_ca_out_377[41:24], u_ca_out_376[47:42]};
assign col_out_380 = {u_ca_out_380[5:0],u_ca_out_379[23:6], u_ca_out_378[41:24], u_ca_out_377[47:42]};
assign col_out_381 = {u_ca_out_381[5:0],u_ca_out_380[23:6], u_ca_out_379[41:24], u_ca_out_378[47:42]};
assign col_out_382 = {u_ca_out_382[5:0],u_ca_out_381[23:6], u_ca_out_380[41:24], u_ca_out_379[47:42]};
assign col_out_383 = {u_ca_out_383[5:0],u_ca_out_382[23:6], u_ca_out_381[41:24], u_ca_out_380[47:42]};
assign col_out_384 = {u_ca_out_384[5:0],u_ca_out_383[23:6], u_ca_out_382[41:24], u_ca_out_381[47:42]};
assign col_out_385 = {u_ca_out_385[5:0],u_ca_out_384[23:6], u_ca_out_383[41:24], u_ca_out_382[47:42]};
assign col_out_386 = {u_ca_out_386[5:0],u_ca_out_385[23:6], u_ca_out_384[41:24], u_ca_out_383[47:42]};
assign col_out_387 = {u_ca_out_387[5:0],u_ca_out_386[23:6], u_ca_out_385[41:24], u_ca_out_384[47:42]};
assign col_out_388 = {u_ca_out_388[5:0],u_ca_out_387[23:6], u_ca_out_386[41:24], u_ca_out_385[47:42]};
assign col_out_389 = {u_ca_out_389[5:0],u_ca_out_388[23:6], u_ca_out_387[41:24], u_ca_out_386[47:42]};
assign col_out_390 = {u_ca_out_390[5:0],u_ca_out_389[23:6], u_ca_out_388[41:24], u_ca_out_387[47:42]};
assign col_out_391 = {u_ca_out_391[5:0],u_ca_out_390[23:6], u_ca_out_389[41:24], u_ca_out_388[47:42]};
assign col_out_392 = {u_ca_out_392[5:0],u_ca_out_391[23:6], u_ca_out_390[41:24], u_ca_out_389[47:42]};
assign col_out_393 = {u_ca_out_393[5:0],u_ca_out_392[23:6], u_ca_out_391[41:24], u_ca_out_390[47:42]};
assign col_out_394 = {u_ca_out_394[5:0],u_ca_out_393[23:6], u_ca_out_392[41:24], u_ca_out_391[47:42]};
assign col_out_395 = {u_ca_out_395[5:0],u_ca_out_394[23:6], u_ca_out_393[41:24], u_ca_out_392[47:42]};
assign col_out_396 = {u_ca_out_396[5:0],u_ca_out_395[23:6], u_ca_out_394[41:24], u_ca_out_393[47:42]};
assign col_out_397 = {u_ca_out_397[5:0],u_ca_out_396[23:6], u_ca_out_395[41:24], u_ca_out_394[47:42]};
assign col_out_398 = {u_ca_out_398[5:0],u_ca_out_397[23:6], u_ca_out_396[41:24], u_ca_out_395[47:42]};
assign col_out_399 = {u_ca_out_399[5:0],u_ca_out_398[23:6], u_ca_out_397[41:24], u_ca_out_396[47:42]};
assign col_out_400 = {u_ca_out_400[5:0],u_ca_out_399[23:6], u_ca_out_398[41:24], u_ca_out_397[47:42]};
assign col_out_401 = {u_ca_out_401[5:0],u_ca_out_400[23:6], u_ca_out_399[41:24], u_ca_out_398[47:42]};
assign col_out_402 = {u_ca_out_402[5:0],u_ca_out_401[23:6], u_ca_out_400[41:24], u_ca_out_399[47:42]};
assign col_out_403 = {u_ca_out_403[5:0],u_ca_out_402[23:6], u_ca_out_401[41:24], u_ca_out_400[47:42]};
assign col_out_404 = {u_ca_out_404[5:0],u_ca_out_403[23:6], u_ca_out_402[41:24], u_ca_out_401[47:42]};
assign col_out_405 = {u_ca_out_405[5:0],u_ca_out_404[23:6], u_ca_out_403[41:24], u_ca_out_402[47:42]};
assign col_out_406 = {u_ca_out_406[5:0],u_ca_out_405[23:6], u_ca_out_404[41:24], u_ca_out_403[47:42]};
assign col_out_407 = {u_ca_out_407[5:0],u_ca_out_406[23:6], u_ca_out_405[41:24], u_ca_out_404[47:42]};
assign col_out_408 = {u_ca_out_408[5:0],u_ca_out_407[23:6], u_ca_out_406[41:24], u_ca_out_405[47:42]};
assign col_out_409 = {u_ca_out_409[5:0],u_ca_out_408[23:6], u_ca_out_407[41:24], u_ca_out_406[47:42]};
assign col_out_410 = {u_ca_out_410[5:0],u_ca_out_409[23:6], u_ca_out_408[41:24], u_ca_out_407[47:42]};
assign col_out_411 = {u_ca_out_411[5:0],u_ca_out_410[23:6], u_ca_out_409[41:24], u_ca_out_408[47:42]};
assign col_out_412 = {u_ca_out_412[5:0],u_ca_out_411[23:6], u_ca_out_410[41:24], u_ca_out_409[47:42]};
assign col_out_413 = {u_ca_out_413[5:0],u_ca_out_412[23:6], u_ca_out_411[41:24], u_ca_out_410[47:42]};
assign col_out_414 = {u_ca_out_414[5:0],u_ca_out_413[23:6], u_ca_out_412[41:24], u_ca_out_411[47:42]};
assign col_out_415 = {u_ca_out_415[5:0],u_ca_out_414[23:6], u_ca_out_413[41:24], u_ca_out_412[47:42]};
assign col_out_416 = {u_ca_out_416[5:0],u_ca_out_415[23:6], u_ca_out_414[41:24], u_ca_out_413[47:42]};
assign col_out_417 = {u_ca_out_417[5:0],u_ca_out_416[23:6], u_ca_out_415[41:24], u_ca_out_414[47:42]};
assign col_out_418 = {u_ca_out_418[5:0],u_ca_out_417[23:6], u_ca_out_416[41:24], u_ca_out_415[47:42]};
assign col_out_419 = {u_ca_out_419[5:0],u_ca_out_418[23:6], u_ca_out_417[41:24], u_ca_out_416[47:42]};
assign col_out_420 = {u_ca_out_420[5:0],u_ca_out_419[23:6], u_ca_out_418[41:24], u_ca_out_417[47:42]};
assign col_out_421 = {u_ca_out_421[5:0],u_ca_out_420[23:6], u_ca_out_419[41:24], u_ca_out_418[47:42]};
assign col_out_422 = {u_ca_out_422[5:0],u_ca_out_421[23:6], u_ca_out_420[41:24], u_ca_out_419[47:42]};
assign col_out_423 = {u_ca_out_423[5:0],u_ca_out_422[23:6], u_ca_out_421[41:24], u_ca_out_420[47:42]};
assign col_out_424 = {u_ca_out_424[5:0],u_ca_out_423[23:6], u_ca_out_422[41:24], u_ca_out_421[47:42]};
assign col_out_425 = {u_ca_out_425[5:0],u_ca_out_424[23:6], u_ca_out_423[41:24], u_ca_out_422[47:42]};
assign col_out_426 = {u_ca_out_426[5:0],u_ca_out_425[23:6], u_ca_out_424[41:24], u_ca_out_423[47:42]};
assign col_out_427 = {u_ca_out_427[5:0],u_ca_out_426[23:6], u_ca_out_425[41:24], u_ca_out_424[47:42]};
assign col_out_428 = {u_ca_out_428[5:0],u_ca_out_427[23:6], u_ca_out_426[41:24], u_ca_out_425[47:42]};
assign col_out_429 = {u_ca_out_429[5:0],u_ca_out_428[23:6], u_ca_out_427[41:24], u_ca_out_426[47:42]};
assign col_out_430 = {u_ca_out_430[5:0],u_ca_out_429[23:6], u_ca_out_428[41:24], u_ca_out_427[47:42]};
assign col_out_431 = {u_ca_out_431[5:0],u_ca_out_430[23:6], u_ca_out_429[41:24], u_ca_out_428[47:42]};
assign col_out_432 = {u_ca_out_432[5:0],u_ca_out_431[23:6], u_ca_out_430[41:24], u_ca_out_429[47:42]};
assign col_out_433 = {u_ca_out_433[5:0],u_ca_out_432[23:6], u_ca_out_431[41:24], u_ca_out_430[47:42]};
assign col_out_434 = {u_ca_out_434[5:0],u_ca_out_433[23:6], u_ca_out_432[41:24], u_ca_out_431[47:42]};
assign col_out_435 = {u_ca_out_435[5:0],u_ca_out_434[23:6], u_ca_out_433[41:24], u_ca_out_432[47:42]};
assign col_out_436 = {u_ca_out_436[5:0],u_ca_out_435[23:6], u_ca_out_434[41:24], u_ca_out_433[47:42]};
assign col_out_437 = {u_ca_out_437[5:0],u_ca_out_436[23:6], u_ca_out_435[41:24], u_ca_out_434[47:42]};
assign col_out_438 = {u_ca_out_438[5:0],u_ca_out_437[23:6], u_ca_out_436[41:24], u_ca_out_435[47:42]};
assign col_out_439 = {u_ca_out_439[5:0],u_ca_out_438[23:6], u_ca_out_437[41:24], u_ca_out_436[47:42]};
assign col_out_440 = {u_ca_out_440[5:0],u_ca_out_439[23:6], u_ca_out_438[41:24], u_ca_out_437[47:42]};
assign col_out_441 = {u_ca_out_441[5:0],u_ca_out_440[23:6], u_ca_out_439[41:24], u_ca_out_438[47:42]};
assign col_out_442 = {u_ca_out_442[5:0],u_ca_out_441[23:6], u_ca_out_440[41:24], u_ca_out_439[47:42]};
assign col_out_443 = {u_ca_out_443[5:0],u_ca_out_442[23:6], u_ca_out_441[41:24], u_ca_out_440[47:42]};
assign col_out_444 = {u_ca_out_444[5:0],u_ca_out_443[23:6], u_ca_out_442[41:24], u_ca_out_441[47:42]};
assign col_out_445 = {u_ca_out_445[5:0],u_ca_out_444[23:6], u_ca_out_443[41:24], u_ca_out_442[47:42]};
assign col_out_446 = {u_ca_out_446[5:0],u_ca_out_445[23:6], u_ca_out_444[41:24], u_ca_out_443[47:42]};
assign col_out_447 = {u_ca_out_447[5:0],u_ca_out_446[23:6], u_ca_out_445[41:24], u_ca_out_444[47:42]};
assign col_out_448 = {u_ca_out_448[5:0],u_ca_out_447[23:6], u_ca_out_446[41:24], u_ca_out_445[47:42]};
assign col_out_449 = {u_ca_out_449[5:0],u_ca_out_448[23:6], u_ca_out_447[41:24], u_ca_out_446[47:42]};
assign col_out_450 = {u_ca_out_450[5:0],u_ca_out_449[23:6], u_ca_out_448[41:24], u_ca_out_447[47:42]};
assign col_out_451 = {u_ca_out_451[5:0],u_ca_out_450[23:6], u_ca_out_449[41:24], u_ca_out_448[47:42]};
assign col_out_452 = {u_ca_out_452[5:0],u_ca_out_451[23:6], u_ca_out_450[41:24], u_ca_out_449[47:42]};
assign col_out_453 = {u_ca_out_453[5:0],u_ca_out_452[23:6], u_ca_out_451[41:24], u_ca_out_450[47:42]};
assign col_out_454 = {u_ca_out_454[5:0],u_ca_out_453[23:6], u_ca_out_452[41:24], u_ca_out_451[47:42]};
assign col_out_455 = {u_ca_out_455[5:0],u_ca_out_454[23:6], u_ca_out_453[41:24], u_ca_out_452[47:42]};
assign col_out_456 = {u_ca_out_456[5:0],u_ca_out_455[23:6], u_ca_out_454[41:24], u_ca_out_453[47:42]};
assign col_out_457 = {u_ca_out_457[5:0],u_ca_out_456[23:6], u_ca_out_455[41:24], u_ca_out_454[47:42]};
assign col_out_458 = {u_ca_out_458[5:0],u_ca_out_457[23:6], u_ca_out_456[41:24], u_ca_out_455[47:42]};
assign col_out_459 = {u_ca_out_459[5:0],u_ca_out_458[23:6], u_ca_out_457[41:24], u_ca_out_456[47:42]};
assign col_out_460 = {u_ca_out_460[5:0],u_ca_out_459[23:6], u_ca_out_458[41:24], u_ca_out_457[47:42]};
assign col_out_461 = {u_ca_out_461[5:0],u_ca_out_460[23:6], u_ca_out_459[41:24], u_ca_out_458[47:42]};
assign col_out_462 = {u_ca_out_462[5:0],u_ca_out_461[23:6], u_ca_out_460[41:24], u_ca_out_459[47:42]};
assign col_out_463 = {u_ca_out_463[5:0],u_ca_out_462[23:6], u_ca_out_461[41:24], u_ca_out_460[47:42]};
assign col_out_464 = {u_ca_out_464[5:0],u_ca_out_463[23:6], u_ca_out_462[41:24], u_ca_out_461[47:42]};
assign col_out_465 = {u_ca_out_465[5:0],u_ca_out_464[23:6], u_ca_out_463[41:24], u_ca_out_462[47:42]};
assign col_out_466 = {u_ca_out_466[5:0],u_ca_out_465[23:6], u_ca_out_464[41:24], u_ca_out_463[47:42]};
assign col_out_467 = {u_ca_out_467[5:0],u_ca_out_466[23:6], u_ca_out_465[41:24], u_ca_out_464[47:42]};
assign col_out_468 = {u_ca_out_468[5:0],u_ca_out_467[23:6], u_ca_out_466[41:24], u_ca_out_465[47:42]};
assign col_out_469 = {u_ca_out_469[5:0],u_ca_out_468[23:6], u_ca_out_467[41:24], u_ca_out_466[47:42]};
assign col_out_470 = {u_ca_out_470[5:0],u_ca_out_469[23:6], u_ca_out_468[41:24], u_ca_out_467[47:42]};
assign col_out_471 = {u_ca_out_471[5:0],u_ca_out_470[23:6], u_ca_out_469[41:24], u_ca_out_468[47:42]};
assign col_out_472 = {u_ca_out_472[5:0],u_ca_out_471[23:6], u_ca_out_470[41:24], u_ca_out_469[47:42]};
assign col_out_473 = {u_ca_out_473[5:0],u_ca_out_472[23:6], u_ca_out_471[41:24], u_ca_out_470[47:42]};
assign col_out_474 = {u_ca_out_474[5:0],u_ca_out_473[23:6], u_ca_out_472[41:24], u_ca_out_471[47:42]};
assign col_out_475 = {u_ca_out_475[5:0],u_ca_out_474[23:6], u_ca_out_473[41:24], u_ca_out_472[47:42]};
assign col_out_476 = {u_ca_out_476[5:0],u_ca_out_475[23:6], u_ca_out_474[41:24], u_ca_out_473[47:42]};
assign col_out_477 = {u_ca_out_477[5:0],u_ca_out_476[23:6], u_ca_out_475[41:24], u_ca_out_474[47:42]};
assign col_out_478 = {u_ca_out_478[5:0],u_ca_out_477[23:6], u_ca_out_476[41:24], u_ca_out_475[47:42]};
assign col_out_479 = {u_ca_out_479[5:0],u_ca_out_478[23:6], u_ca_out_477[41:24], u_ca_out_476[47:42]};
assign col_out_480 = {u_ca_out_480[5:0],u_ca_out_479[23:6], u_ca_out_478[41:24], u_ca_out_477[47:42]};
assign col_out_481 = {u_ca_out_481[5:0],u_ca_out_480[23:6], u_ca_out_479[41:24], u_ca_out_478[47:42]};
assign col_out_482 = {u_ca_out_482[5:0],u_ca_out_481[23:6], u_ca_out_480[41:24], u_ca_out_479[47:42]};
assign col_out_483 = {u_ca_out_483[5:0],u_ca_out_482[23:6], u_ca_out_481[41:24], u_ca_out_480[47:42]};
assign col_out_484 = {u_ca_out_484[5:0],u_ca_out_483[23:6], u_ca_out_482[41:24], u_ca_out_481[47:42]};
assign col_out_485 = {u_ca_out_485[5:0],u_ca_out_484[23:6], u_ca_out_483[41:24], u_ca_out_482[47:42]};
assign col_out_486 = {u_ca_out_486[5:0],u_ca_out_485[23:6], u_ca_out_484[41:24], u_ca_out_483[47:42]};
assign col_out_487 = {u_ca_out_487[5:0],u_ca_out_486[23:6], u_ca_out_485[41:24], u_ca_out_484[47:42]};
assign col_out_488 = {u_ca_out_488[5:0],u_ca_out_487[23:6], u_ca_out_486[41:24], u_ca_out_485[47:42]};
assign col_out_489 = {u_ca_out_489[5:0],u_ca_out_488[23:6], u_ca_out_487[41:24], u_ca_out_486[47:42]};
assign col_out_490 = {u_ca_out_490[5:0],u_ca_out_489[23:6], u_ca_out_488[41:24], u_ca_out_487[47:42]};
assign col_out_491 = {u_ca_out_491[5:0],u_ca_out_490[23:6], u_ca_out_489[41:24], u_ca_out_488[47:42]};
assign col_out_492 = {u_ca_out_492[5:0],u_ca_out_491[23:6], u_ca_out_490[41:24], u_ca_out_489[47:42]};
assign col_out_493 = {u_ca_out_493[5:0],u_ca_out_492[23:6], u_ca_out_491[41:24], u_ca_out_490[47:42]};
assign col_out_494 = {u_ca_out_494[5:0],u_ca_out_493[23:6], u_ca_out_492[41:24], u_ca_out_491[47:42]};
assign col_out_495 = {u_ca_out_495[5:0],u_ca_out_494[23:6], u_ca_out_493[41:24], u_ca_out_492[47:42]};
assign col_out_496 = {u_ca_out_496[5:0],u_ca_out_495[23:6], u_ca_out_494[41:24], u_ca_out_493[47:42]};
assign col_out_497 = {u_ca_out_497[5:0],u_ca_out_496[23:6], u_ca_out_495[41:24], u_ca_out_494[47:42]};
assign col_out_498 = {u_ca_out_498[5:0],u_ca_out_497[23:6], u_ca_out_496[41:24], u_ca_out_495[47:42]};
assign col_out_499 = {u_ca_out_499[5:0],u_ca_out_498[23:6], u_ca_out_497[41:24], u_ca_out_496[47:42]};
assign col_out_500 = {u_ca_out_500[5:0],u_ca_out_499[23:6], u_ca_out_498[41:24], u_ca_out_497[47:42]};
assign col_out_501 = {u_ca_out_501[5:0],u_ca_out_500[23:6], u_ca_out_499[41:24], u_ca_out_498[47:42]};
assign col_out_502 = {u_ca_out_502[5:0],u_ca_out_501[23:6], u_ca_out_500[41:24], u_ca_out_499[47:42]};
assign col_out_503 = {u_ca_out_503[5:0],u_ca_out_502[23:6], u_ca_out_501[41:24], u_ca_out_500[47:42]};
assign col_out_504 = {u_ca_out_504[5:0],u_ca_out_503[23:6], u_ca_out_502[41:24], u_ca_out_501[47:42]};
assign col_out_505 = {u_ca_out_505[5:0],u_ca_out_504[23:6], u_ca_out_503[41:24], u_ca_out_502[47:42]};
assign col_out_506 = {u_ca_out_506[5:0],u_ca_out_505[23:6], u_ca_out_504[41:24], u_ca_out_503[47:42]};
assign col_out_507 = {u_ca_out_507[5:0],u_ca_out_506[23:6], u_ca_out_505[41:24], u_ca_out_504[47:42]};
assign col_out_508 = {u_ca_out_508[5:0],u_ca_out_507[23:6], u_ca_out_506[41:24], u_ca_out_505[47:42]};
assign col_out_509 = {u_ca_out_509[5:0],u_ca_out_508[23:6], u_ca_out_507[41:24], u_ca_out_506[47:42]};
assign col_out_510 = {u_ca_out_510[5:0],u_ca_out_509[23:6], u_ca_out_508[41:24], u_ca_out_507[47:42]};
assign col_out_511 = {u_ca_out_511[5:0],u_ca_out_510[23:6], u_ca_out_509[41:24], u_ca_out_508[47:42]};
assign col_out_512 = {u_ca_out_512[5:0],u_ca_out_511[23:6], u_ca_out_510[41:24], u_ca_out_509[47:42]};
assign col_out_513 = {u_ca_out_513[5:0],u_ca_out_512[23:6], u_ca_out_511[41:24], u_ca_out_510[47:42]};
assign col_out_514 = {u_ca_out_514[5:0],u_ca_out_513[23:6], u_ca_out_512[41:24], u_ca_out_511[47:42]};
assign col_out_515 = {u_ca_out_515[5:0],u_ca_out_514[23:6], u_ca_out_513[41:24], u_ca_out_512[47:42]};
assign col_out_516 = {u_ca_out_516[5:0],u_ca_out_515[23:6], u_ca_out_514[41:24], u_ca_out_513[47:42]};
assign col_out_517 = {u_ca_out_517[5:0],u_ca_out_516[23:6], u_ca_out_515[41:24], u_ca_out_514[47:42]};
assign col_out_518 = {u_ca_out_518[5:0],u_ca_out_517[23:6], u_ca_out_516[41:24], u_ca_out_515[47:42]};
assign col_out_519 = {u_ca_out_519[5:0],u_ca_out_518[23:6], u_ca_out_517[41:24], u_ca_out_516[47:42]};
assign col_out_520 = {u_ca_out_520[5:0],u_ca_out_519[23:6], u_ca_out_518[41:24], u_ca_out_517[47:42]};
assign col_out_521 = {u_ca_out_521[5:0],u_ca_out_520[23:6], u_ca_out_519[41:24], u_ca_out_518[47:42]};
assign col_out_522 = {u_ca_out_522[5:0],u_ca_out_521[23:6], u_ca_out_520[41:24], u_ca_out_519[47:42]};
assign col_out_523 = {u_ca_out_523[5:0],u_ca_out_522[23:6], u_ca_out_521[41:24], u_ca_out_520[47:42]};
assign col_out_524 = {u_ca_out_524[5:0],u_ca_out_523[23:6], u_ca_out_522[41:24], u_ca_out_521[47:42]};
assign col_out_525 = {u_ca_out_525[5:0],u_ca_out_524[23:6], u_ca_out_523[41:24], u_ca_out_522[47:42]};
assign col_out_526 = {u_ca_out_526[5:0],u_ca_out_525[23:6], u_ca_out_524[41:24], u_ca_out_523[47:42]};
assign col_out_527 = {u_ca_out_527[5:0],u_ca_out_526[23:6], u_ca_out_525[41:24], u_ca_out_524[47:42]};
assign col_out_528 = {u_ca_out_528[5:0],u_ca_out_527[23:6], u_ca_out_526[41:24], u_ca_out_525[47:42]};
assign col_out_529 = {u_ca_out_529[5:0],u_ca_out_528[23:6], u_ca_out_527[41:24], u_ca_out_526[47:42]};
assign col_out_530 = {u_ca_out_530[5:0],u_ca_out_529[23:6], u_ca_out_528[41:24], u_ca_out_527[47:42]};
assign col_out_531 = {u_ca_out_531[5:0],u_ca_out_530[23:6], u_ca_out_529[41:24], u_ca_out_528[47:42]};
assign col_out_532 = {u_ca_out_532[5:0],u_ca_out_531[23:6], u_ca_out_530[41:24], u_ca_out_529[47:42]};
assign col_out_533 = {u_ca_out_533[5:0],u_ca_out_532[23:6], u_ca_out_531[41:24], u_ca_out_530[47:42]};
assign col_out_534 = {u_ca_out_534[5:0],u_ca_out_533[23:6], u_ca_out_532[41:24], u_ca_out_531[47:42]};
assign col_out_535 = {u_ca_out_535[5:0],u_ca_out_534[23:6], u_ca_out_533[41:24], u_ca_out_532[47:42]};
assign col_out_536 = {u_ca_out_536[5:0],u_ca_out_535[23:6], u_ca_out_534[41:24], u_ca_out_533[47:42]};
assign col_out_537 = {u_ca_out_537[5:0],u_ca_out_536[23:6], u_ca_out_535[41:24], u_ca_out_534[47:42]};
assign col_out_538 = {u_ca_out_538[5:0],u_ca_out_537[23:6], u_ca_out_536[41:24], u_ca_out_535[47:42]};
assign col_out_539 = {u_ca_out_539[5:0],u_ca_out_538[23:6], u_ca_out_537[41:24], u_ca_out_536[47:42]};
assign col_out_540 = {u_ca_out_540[5:0],u_ca_out_539[23:6], u_ca_out_538[41:24], u_ca_out_537[47:42]};
assign col_out_541 = {u_ca_out_541[5:0],u_ca_out_540[23:6], u_ca_out_539[41:24], u_ca_out_538[47:42]};
assign col_out_542 = {u_ca_out_542[5:0],u_ca_out_541[23:6], u_ca_out_540[41:24], u_ca_out_539[47:42]};
assign col_out_543 = {u_ca_out_543[5:0],u_ca_out_542[23:6], u_ca_out_541[41:24], u_ca_out_540[47:42]};
assign col_out_544 = {u_ca_out_544[5:0],u_ca_out_543[23:6], u_ca_out_542[41:24], u_ca_out_541[47:42]};
assign col_out_545 = {u_ca_out_545[5:0],u_ca_out_544[23:6], u_ca_out_543[41:24], u_ca_out_542[47:42]};
assign col_out_546 = {u_ca_out_546[5:0],u_ca_out_545[23:6], u_ca_out_544[41:24], u_ca_out_543[47:42]};
assign col_out_547 = {u_ca_out_547[5:0],u_ca_out_546[23:6], u_ca_out_545[41:24], u_ca_out_544[47:42]};
assign col_out_548 = {u_ca_out_548[5:0],u_ca_out_547[23:6], u_ca_out_546[41:24], u_ca_out_545[47:42]};
assign col_out_549 = {u_ca_out_549[5:0],u_ca_out_548[23:6], u_ca_out_547[41:24], u_ca_out_546[47:42]};
assign col_out_550 = {u_ca_out_550[5:0],u_ca_out_549[23:6], u_ca_out_548[41:24], u_ca_out_547[47:42]};
assign col_out_551 = {u_ca_out_551[5:0],u_ca_out_550[23:6], u_ca_out_549[41:24], u_ca_out_548[47:42]};
assign col_out_552 = {u_ca_out_552[5:0],u_ca_out_551[23:6], u_ca_out_550[41:24], u_ca_out_549[47:42]};
assign col_out_553 = {u_ca_out_553[5:0],u_ca_out_552[23:6], u_ca_out_551[41:24], u_ca_out_550[47:42]};
assign col_out_554 = {u_ca_out_554[5:0],u_ca_out_553[23:6], u_ca_out_552[41:24], u_ca_out_551[47:42]};
assign col_out_555 = {u_ca_out_555[5:0],u_ca_out_554[23:6], u_ca_out_553[41:24], u_ca_out_552[47:42]};
assign col_out_556 = {u_ca_out_556[5:0],u_ca_out_555[23:6], u_ca_out_554[41:24], u_ca_out_553[47:42]};
assign col_out_557 = {u_ca_out_557[5:0],u_ca_out_556[23:6], u_ca_out_555[41:24], u_ca_out_554[47:42]};
assign col_out_558 = {u_ca_out_558[5:0],u_ca_out_557[23:6], u_ca_out_556[41:24], u_ca_out_555[47:42]};
assign col_out_559 = {u_ca_out_559[5:0],u_ca_out_558[23:6], u_ca_out_557[41:24], u_ca_out_556[47:42]};
assign col_out_560 = {u_ca_out_560[5:0],u_ca_out_559[23:6], u_ca_out_558[41:24], u_ca_out_557[47:42]};
assign col_out_561 = {u_ca_out_561[5:0],u_ca_out_560[23:6], u_ca_out_559[41:24], u_ca_out_558[47:42]};
assign col_out_562 = {u_ca_out_562[5:0],u_ca_out_561[23:6], u_ca_out_560[41:24], u_ca_out_559[47:42]};
assign col_out_563 = {u_ca_out_563[5:0],u_ca_out_562[23:6], u_ca_out_561[41:24], u_ca_out_560[47:42]};
assign col_out_564 = {u_ca_out_564[5:0],u_ca_out_563[23:6], u_ca_out_562[41:24], u_ca_out_561[47:42]};
assign col_out_565 = {u_ca_out_565[5:0],u_ca_out_564[23:6], u_ca_out_563[41:24], u_ca_out_562[47:42]};
assign col_out_566 = {u_ca_out_566[5:0],u_ca_out_565[23:6], u_ca_out_564[41:24], u_ca_out_563[47:42]};
assign col_out_567 = {u_ca_out_567[5:0],u_ca_out_566[23:6], u_ca_out_565[41:24], u_ca_out_564[47:42]};
assign col_out_568 = {u_ca_out_568[5:0],u_ca_out_567[23:6], u_ca_out_566[41:24], u_ca_out_565[47:42]};
assign col_out_569 = {u_ca_out_569[5:0],u_ca_out_568[23:6], u_ca_out_567[41:24], u_ca_out_566[47:42]};
assign col_out_570 = {u_ca_out_570[5:0],u_ca_out_569[23:6], u_ca_out_568[41:24], u_ca_out_567[47:42]};
assign col_out_571 = {u_ca_out_571[5:0],u_ca_out_570[23:6], u_ca_out_569[41:24], u_ca_out_568[47:42]};
assign col_out_572 = {u_ca_out_572[5:0],u_ca_out_571[23:6], u_ca_out_570[41:24], u_ca_out_569[47:42]};
assign col_out_573 = {u_ca_out_573[5:0],u_ca_out_572[23:6], u_ca_out_571[41:24], u_ca_out_570[47:42]};
assign col_out_574 = {u_ca_out_574[5:0],u_ca_out_573[23:6], u_ca_out_572[41:24], u_ca_out_571[47:42]};
assign col_out_575 = {u_ca_out_575[5:0],u_ca_out_574[23:6], u_ca_out_573[41:24], u_ca_out_572[47:42]};
assign col_out_576 = {u_ca_out_576[5:0],u_ca_out_575[23:6], u_ca_out_574[41:24], u_ca_out_573[47:42]};
assign col_out_577 = {u_ca_out_577[5:0],u_ca_out_576[23:6], u_ca_out_575[41:24], u_ca_out_574[47:42]};
assign col_out_578 = {u_ca_out_578[5:0],u_ca_out_577[23:6], u_ca_out_576[41:24], u_ca_out_575[47:42]};
assign col_out_579 = {u_ca_out_579[5:0],u_ca_out_578[23:6], u_ca_out_577[41:24], u_ca_out_576[47:42]};
assign col_out_580 = {u_ca_out_580[5:0],u_ca_out_579[23:6], u_ca_out_578[41:24], u_ca_out_577[47:42]};
assign col_out_581 = {u_ca_out_581[5:0],u_ca_out_580[23:6], u_ca_out_579[41:24], u_ca_out_578[47:42]};
assign col_out_582 = {u_ca_out_582[5:0],u_ca_out_581[23:6], u_ca_out_580[41:24], u_ca_out_579[47:42]};
assign col_out_583 = {u_ca_out_583[5:0],u_ca_out_582[23:6], u_ca_out_581[41:24], u_ca_out_580[47:42]};
assign col_out_584 = {u_ca_out_584[5:0],u_ca_out_583[23:6], u_ca_out_582[41:24], u_ca_out_581[47:42]};
assign col_out_585 = {u_ca_out_585[5:0],u_ca_out_584[23:6], u_ca_out_583[41:24], u_ca_out_582[47:42]};
assign col_out_586 = {u_ca_out_586[5:0],u_ca_out_585[23:6], u_ca_out_584[41:24], u_ca_out_583[47:42]};
assign col_out_587 = {u_ca_out_587[5:0],u_ca_out_586[23:6], u_ca_out_585[41:24], u_ca_out_584[47:42]};
assign col_out_588 = {u_ca_out_588[5:0],u_ca_out_587[23:6], u_ca_out_586[41:24], u_ca_out_585[47:42]};
assign col_out_589 = {u_ca_out_589[5:0],u_ca_out_588[23:6], u_ca_out_587[41:24], u_ca_out_586[47:42]};
assign col_out_590 = {u_ca_out_590[5:0],u_ca_out_589[23:6], u_ca_out_588[41:24], u_ca_out_587[47:42]};
assign col_out_591 = {u_ca_out_591[5:0],u_ca_out_590[23:6], u_ca_out_589[41:24], u_ca_out_588[47:42]};
assign col_out_592 = {u_ca_out_592[5:0],u_ca_out_591[23:6], u_ca_out_590[41:24], u_ca_out_589[47:42]};
assign col_out_593 = {u_ca_out_593[5:0],u_ca_out_592[23:6], u_ca_out_591[41:24], u_ca_out_590[47:42]};
assign col_out_594 = {u_ca_out_594[5:0],u_ca_out_593[23:6], u_ca_out_592[41:24], u_ca_out_591[47:42]};
assign col_out_595 = {u_ca_out_595[5:0],u_ca_out_594[23:6], u_ca_out_593[41:24], u_ca_out_592[47:42]};
assign col_out_596 = {u_ca_out_596[5:0],u_ca_out_595[23:6], u_ca_out_594[41:24], u_ca_out_593[47:42]};
assign col_out_597 = {u_ca_out_597[5:0],u_ca_out_596[23:6], u_ca_out_595[41:24], u_ca_out_594[47:42]};
assign col_out_598 = {u_ca_out_598[5:0],u_ca_out_597[23:6], u_ca_out_596[41:24], u_ca_out_595[47:42]};
assign col_out_599 = {u_ca_out_599[5:0],u_ca_out_598[23:6], u_ca_out_597[41:24], u_ca_out_596[47:42]};
assign col_out_600 = {u_ca_out_600[5:0],u_ca_out_599[23:6], u_ca_out_598[41:24], u_ca_out_597[47:42]};
assign col_out_601 = {u_ca_out_601[5:0],u_ca_out_600[23:6], u_ca_out_599[41:24], u_ca_out_598[47:42]};
assign col_out_602 = {u_ca_out_602[5:0],u_ca_out_601[23:6], u_ca_out_600[41:24], u_ca_out_599[47:42]};
assign col_out_603 = {u_ca_out_603[5:0],u_ca_out_602[23:6], u_ca_out_601[41:24], u_ca_out_600[47:42]};
assign col_out_604 = {u_ca_out_604[5:0],u_ca_out_603[23:6], u_ca_out_602[41:24], u_ca_out_601[47:42]};
assign col_out_605 = {u_ca_out_605[5:0],u_ca_out_604[23:6], u_ca_out_603[41:24], u_ca_out_602[47:42]};
assign col_out_606 = {u_ca_out_606[5:0],u_ca_out_605[23:6], u_ca_out_604[41:24], u_ca_out_603[47:42]};
assign col_out_607 = {u_ca_out_607[5:0],u_ca_out_606[23:6], u_ca_out_605[41:24], u_ca_out_604[47:42]};
assign col_out_608 = {u_ca_out_608[5:0],u_ca_out_607[23:6], u_ca_out_606[41:24], u_ca_out_605[47:42]};
assign col_out_609 = {u_ca_out_609[5:0],u_ca_out_608[23:6], u_ca_out_607[41:24], u_ca_out_606[47:42]};
assign col_out_610 = {u_ca_out_610[5:0],u_ca_out_609[23:6], u_ca_out_608[41:24], u_ca_out_607[47:42]};
assign col_out_611 = {u_ca_out_611[5:0],u_ca_out_610[23:6], u_ca_out_609[41:24], u_ca_out_608[47:42]};
assign col_out_612 = {u_ca_out_612[5:0],u_ca_out_611[23:6], u_ca_out_610[41:24], u_ca_out_609[47:42]};
assign col_out_613 = {u_ca_out_613[5:0],u_ca_out_612[23:6], u_ca_out_611[41:24], u_ca_out_610[47:42]};
assign col_out_614 = {u_ca_out_614[5:0],u_ca_out_613[23:6], u_ca_out_612[41:24], u_ca_out_611[47:42]};
assign col_out_615 = {u_ca_out_615[5:0],u_ca_out_614[23:6], u_ca_out_613[41:24], u_ca_out_612[47:42]};
assign col_out_616 = {u_ca_out_616[5:0],u_ca_out_615[23:6], u_ca_out_614[41:24], u_ca_out_613[47:42]};
assign col_out_617 = {u_ca_out_617[5:0],u_ca_out_616[23:6], u_ca_out_615[41:24], u_ca_out_614[47:42]};
assign col_out_618 = {u_ca_out_618[5:0],u_ca_out_617[23:6], u_ca_out_616[41:24], u_ca_out_615[47:42]};
assign col_out_619 = {u_ca_out_619[5:0],u_ca_out_618[23:6], u_ca_out_617[41:24], u_ca_out_616[47:42]};
assign col_out_620 = {u_ca_out_620[5:0],u_ca_out_619[23:6], u_ca_out_618[41:24], u_ca_out_617[47:42]};
assign col_out_621 = {u_ca_out_621[5:0],u_ca_out_620[23:6], u_ca_out_619[41:24], u_ca_out_618[47:42]};
assign col_out_622 = {u_ca_out_622[5:0],u_ca_out_621[23:6], u_ca_out_620[41:24], u_ca_out_619[47:42]};
assign col_out_623 = {u_ca_out_623[5:0],u_ca_out_622[23:6], u_ca_out_621[41:24], u_ca_out_620[47:42]};
assign col_out_624 = {u_ca_out_624[5:0],u_ca_out_623[23:6], u_ca_out_622[41:24], u_ca_out_621[47:42]};
assign col_out_625 = {u_ca_out_625[5:0],u_ca_out_624[23:6], u_ca_out_623[41:24], u_ca_out_622[47:42]};
assign col_out_626 = {u_ca_out_626[5:0],u_ca_out_625[23:6], u_ca_out_624[41:24], u_ca_out_623[47:42]};
assign col_out_627 = {u_ca_out_627[5:0],u_ca_out_626[23:6], u_ca_out_625[41:24], u_ca_out_624[47:42]};
assign col_out_628 = {u_ca_out_628[5:0],u_ca_out_627[23:6], u_ca_out_626[41:24], u_ca_out_625[47:42]};
assign col_out_629 = {u_ca_out_629[5:0],u_ca_out_628[23:6], u_ca_out_627[41:24], u_ca_out_626[47:42]};
assign col_out_630 = {u_ca_out_630[5:0],u_ca_out_629[23:6], u_ca_out_628[41:24], u_ca_out_627[47:42]};
assign col_out_631 = {u_ca_out_631[5:0],u_ca_out_630[23:6], u_ca_out_629[41:24], u_ca_out_628[47:42]};
assign col_out_632 = {u_ca_out_632[5:0],u_ca_out_631[23:6], u_ca_out_630[41:24], u_ca_out_629[47:42]};
assign col_out_633 = {u_ca_out_633[5:0],u_ca_out_632[23:6], u_ca_out_631[41:24], u_ca_out_630[47:42]};
assign col_out_634 = {u_ca_out_634[5:0],u_ca_out_633[23:6], u_ca_out_632[41:24], u_ca_out_631[47:42]};
assign col_out_635 = {u_ca_out_635[5:0],u_ca_out_634[23:6], u_ca_out_633[41:24], u_ca_out_632[47:42]};
assign col_out_636 = {u_ca_out_636[5:0],u_ca_out_635[23:6], u_ca_out_634[41:24], u_ca_out_633[47:42]};
assign col_out_637 = {u_ca_out_637[5:0],u_ca_out_636[23:6], u_ca_out_635[41:24], u_ca_out_634[47:42]};
assign col_out_638 = {u_ca_out_638[5:0],u_ca_out_637[23:6], u_ca_out_636[41:24], u_ca_out_635[47:42]};
assign col_out_639 = {u_ca_out_639[5:0],u_ca_out_638[23:6], u_ca_out_637[41:24], u_ca_out_636[47:42]};
assign col_out_640 = {u_ca_out_640[5:0],u_ca_out_639[23:6], u_ca_out_638[41:24], u_ca_out_637[47:42]};
assign col_out_641 = {u_ca_out_641[5:0],u_ca_out_640[23:6], u_ca_out_639[41:24], u_ca_out_638[47:42]};
assign col_out_642 = {u_ca_out_642[5:0],u_ca_out_641[23:6], u_ca_out_640[41:24], u_ca_out_639[47:42]};
assign col_out_643 = {u_ca_out_643[5:0],u_ca_out_642[23:6], u_ca_out_641[41:24], u_ca_out_640[47:42]};
assign col_out_644 = {u_ca_out_644[5:0],u_ca_out_643[23:6], u_ca_out_642[41:24], u_ca_out_641[47:42]};
assign col_out_645 = {u_ca_out_645[5:0],u_ca_out_644[23:6], u_ca_out_643[41:24], u_ca_out_642[47:42]};
assign col_out_646 = {u_ca_out_646[5:0],u_ca_out_645[23:6], u_ca_out_644[41:24], u_ca_out_643[47:42]};
assign col_out_647 = {u_ca_out_647[5:0],u_ca_out_646[23:6], u_ca_out_645[41:24], u_ca_out_644[47:42]};
assign col_out_648 = {u_ca_out_648[5:0],u_ca_out_647[23:6], u_ca_out_646[41:24], u_ca_out_645[47:42]};
assign col_out_649 = {u_ca_out_649[5:0],u_ca_out_648[23:6], u_ca_out_647[41:24], u_ca_out_646[47:42]};
assign col_out_650 = {u_ca_out_650[5:0],u_ca_out_649[23:6], u_ca_out_648[41:24], u_ca_out_647[47:42]};
assign col_out_651 = {u_ca_out_651[5:0],u_ca_out_650[23:6], u_ca_out_649[41:24], u_ca_out_648[47:42]};
assign col_out_652 = {u_ca_out_652[5:0],u_ca_out_651[23:6], u_ca_out_650[41:24], u_ca_out_649[47:42]};
assign col_out_653 = {u_ca_out_653[5:0],u_ca_out_652[23:6], u_ca_out_651[41:24], u_ca_out_650[47:42]};
assign col_out_654 = {u_ca_out_654[5:0],u_ca_out_653[23:6], u_ca_out_652[41:24], u_ca_out_651[47:42]};
assign col_out_655 = {u_ca_out_655[5:0],u_ca_out_654[23:6], u_ca_out_653[41:24], u_ca_out_652[47:42]};
assign col_out_656 = {u_ca_out_656[5:0],u_ca_out_655[23:6], u_ca_out_654[41:24], u_ca_out_653[47:42]};
assign col_out_657 = {u_ca_out_657[5:0],u_ca_out_656[23:6], u_ca_out_655[41:24], u_ca_out_654[47:42]};
assign col_out_658 = {u_ca_out_658[5:0],u_ca_out_657[23:6], u_ca_out_656[41:24], u_ca_out_655[47:42]};
assign col_out_659 = {u_ca_out_659[5:0],u_ca_out_658[23:6], u_ca_out_657[41:24], u_ca_out_656[47:42]};
assign col_out_660 = {u_ca_out_660[5:0],u_ca_out_659[23:6], u_ca_out_658[41:24], u_ca_out_657[47:42]};
assign col_out_661 = {u_ca_out_661[5:0],u_ca_out_660[23:6], u_ca_out_659[41:24], u_ca_out_658[47:42]};
assign col_out_662 = {u_ca_out_662[5:0],u_ca_out_661[23:6], u_ca_out_660[41:24], u_ca_out_659[47:42]};
assign col_out_663 = {u_ca_out_663[5:0],u_ca_out_662[23:6], u_ca_out_661[41:24], u_ca_out_660[47:42]};
assign col_out_664 = {u_ca_out_664[5:0],u_ca_out_663[23:6], u_ca_out_662[41:24], u_ca_out_661[47:42]};
assign col_out_665 = {u_ca_out_665[5:0],u_ca_out_664[23:6], u_ca_out_663[41:24], u_ca_out_662[47:42]};
assign col_out_666 = {u_ca_out_666[5:0],u_ca_out_665[23:6], u_ca_out_664[41:24], u_ca_out_663[47:42]};
assign col_out_667 = {u_ca_out_667[5:0],u_ca_out_666[23:6], u_ca_out_665[41:24], u_ca_out_664[47:42]};
assign col_out_668 = {u_ca_out_668[5:0],u_ca_out_667[23:6], u_ca_out_666[41:24], u_ca_out_665[47:42]};
assign col_out_669 = {u_ca_out_669[5:0],u_ca_out_668[23:6], u_ca_out_667[41:24], u_ca_out_666[47:42]};
assign col_out_670 = {u_ca_out_670[5:0],u_ca_out_669[23:6], u_ca_out_668[41:24], u_ca_out_667[47:42]};
assign col_out_671 = {u_ca_out_671[5:0],u_ca_out_670[23:6], u_ca_out_669[41:24], u_ca_out_668[47:42]};
assign col_out_672 = {u_ca_out_672[5:0],u_ca_out_671[23:6], u_ca_out_670[41:24], u_ca_out_669[47:42]};
assign col_out_673 = {u_ca_out_673[5:0],u_ca_out_672[23:6], u_ca_out_671[41:24], u_ca_out_670[47:42]};
assign col_out_674 = {u_ca_out_674[5:0],u_ca_out_673[23:6], u_ca_out_672[41:24], u_ca_out_671[47:42]};
assign col_out_675 = {u_ca_out_675[5:0],u_ca_out_674[23:6], u_ca_out_673[41:24], u_ca_out_672[47:42]};
assign col_out_676 = {u_ca_out_676[5:0],u_ca_out_675[23:6], u_ca_out_674[41:24], u_ca_out_673[47:42]};
assign col_out_677 = {u_ca_out_677[5:0],u_ca_out_676[23:6], u_ca_out_675[41:24], u_ca_out_674[47:42]};
assign col_out_678 = {u_ca_out_678[5:0],u_ca_out_677[23:6], u_ca_out_676[41:24], u_ca_out_675[47:42]};
assign col_out_679 = {u_ca_out_679[5:0],u_ca_out_678[23:6], u_ca_out_677[41:24], u_ca_out_676[47:42]};
assign col_out_680 = {u_ca_out_680[5:0],u_ca_out_679[23:6], u_ca_out_678[41:24], u_ca_out_677[47:42]};
assign col_out_681 = {u_ca_out_681[5:0],u_ca_out_680[23:6], u_ca_out_679[41:24], u_ca_out_678[47:42]};
assign col_out_682 = {u_ca_out_682[5:0],u_ca_out_681[23:6], u_ca_out_680[41:24], u_ca_out_679[47:42]};
assign col_out_683 = {u_ca_out_683[5:0],u_ca_out_682[23:6], u_ca_out_681[41:24], u_ca_out_680[47:42]};
assign col_out_684 = {u_ca_out_684[5:0],u_ca_out_683[23:6], u_ca_out_682[41:24], u_ca_out_681[47:42]};
assign col_out_685 = {u_ca_out_685[5:0],u_ca_out_684[23:6], u_ca_out_683[41:24], u_ca_out_682[47:42]};
assign col_out_686 = {u_ca_out_686[5:0],u_ca_out_685[23:6], u_ca_out_684[41:24], u_ca_out_683[47:42]};
assign col_out_687 = {u_ca_out_687[5:0],u_ca_out_686[23:6], u_ca_out_685[41:24], u_ca_out_684[47:42]};
assign col_out_688 = {u_ca_out_688[5:0],u_ca_out_687[23:6], u_ca_out_686[41:24], u_ca_out_685[47:42]};
assign col_out_689 = {u_ca_out_689[5:0],u_ca_out_688[23:6], u_ca_out_687[41:24], u_ca_out_686[47:42]};
assign col_out_690 = {u_ca_out_690[5:0],u_ca_out_689[23:6], u_ca_out_688[41:24], u_ca_out_687[47:42]};
assign col_out_691 = {u_ca_out_691[5:0],u_ca_out_690[23:6], u_ca_out_689[41:24], u_ca_out_688[47:42]};
assign col_out_692 = {u_ca_out_692[5:0],u_ca_out_691[23:6], u_ca_out_690[41:24], u_ca_out_689[47:42]};
assign col_out_693 = {u_ca_out_693[5:0],u_ca_out_692[23:6], u_ca_out_691[41:24], u_ca_out_690[47:42]};
assign col_out_694 = {u_ca_out_694[5:0],u_ca_out_693[23:6], u_ca_out_692[41:24], u_ca_out_691[47:42]};
assign col_out_695 = {u_ca_out_695[5:0],u_ca_out_694[23:6], u_ca_out_693[41:24], u_ca_out_692[47:42]};
assign col_out_696 = {u_ca_out_696[5:0],u_ca_out_695[23:6], u_ca_out_694[41:24], u_ca_out_693[47:42]};
assign col_out_697 = {u_ca_out_697[5:0],u_ca_out_696[23:6], u_ca_out_695[41:24], u_ca_out_694[47:42]};
assign col_out_698 = {u_ca_out_698[5:0],u_ca_out_697[23:6], u_ca_out_696[41:24], u_ca_out_695[47:42]};
assign col_out_699 = {u_ca_out_699[5:0],u_ca_out_698[23:6], u_ca_out_697[41:24], u_ca_out_696[47:42]};
assign col_out_700 = {u_ca_out_700[5:0],u_ca_out_699[23:6], u_ca_out_698[41:24], u_ca_out_697[47:42]};
assign col_out_701 = {u_ca_out_701[5:0],u_ca_out_700[23:6], u_ca_out_699[41:24], u_ca_out_698[47:42]};
assign col_out_702 = {u_ca_out_702[5:0],u_ca_out_701[23:6], u_ca_out_700[41:24], u_ca_out_699[47:42]};
assign col_out_703 = {u_ca_out_703[5:0],u_ca_out_702[23:6], u_ca_out_701[41:24], u_ca_out_700[47:42]};
assign col_out_704 = {u_ca_out_704[5:0],u_ca_out_703[23:6], u_ca_out_702[41:24], u_ca_out_701[47:42]};
assign col_out_705 = {u_ca_out_705[5:0],u_ca_out_704[23:6], u_ca_out_703[41:24], u_ca_out_702[47:42]};
assign col_out_706 = {u_ca_out_706[5:0],u_ca_out_705[23:6], u_ca_out_704[41:24], u_ca_out_703[47:42]};
assign col_out_707 = {u_ca_out_707[5:0],u_ca_out_706[23:6], u_ca_out_705[41:24], u_ca_out_704[47:42]};
assign col_out_708 = {u_ca_out_708[5:0],u_ca_out_707[23:6], u_ca_out_706[41:24], u_ca_out_705[47:42]};
assign col_out_709 = {u_ca_out_709[5:0],u_ca_out_708[23:6], u_ca_out_707[41:24], u_ca_out_706[47:42]};
assign col_out_710 = {u_ca_out_710[5:0],u_ca_out_709[23:6], u_ca_out_708[41:24], u_ca_out_707[47:42]};
assign col_out_711 = {u_ca_out_711[5:0],u_ca_out_710[23:6], u_ca_out_709[41:24], u_ca_out_708[47:42]};
assign col_out_712 = {u_ca_out_712[5:0],u_ca_out_711[23:6], u_ca_out_710[41:24], u_ca_out_709[47:42]};
assign col_out_713 = {u_ca_out_713[5:0],u_ca_out_712[23:6], u_ca_out_711[41:24], u_ca_out_710[47:42]};
assign col_out_714 = {u_ca_out_714[5:0],u_ca_out_713[23:6], u_ca_out_712[41:24], u_ca_out_711[47:42]};
assign col_out_715 = {u_ca_out_715[5:0],u_ca_out_714[23:6], u_ca_out_713[41:24], u_ca_out_712[47:42]};
assign col_out_716 = {u_ca_out_716[5:0],u_ca_out_715[23:6], u_ca_out_714[41:24], u_ca_out_713[47:42]};
assign col_out_717 = {u_ca_out_717[5:0],u_ca_out_716[23:6], u_ca_out_715[41:24], u_ca_out_714[47:42]};
assign col_out_718 = {u_ca_out_718[5:0],u_ca_out_717[23:6], u_ca_out_716[41:24], u_ca_out_715[47:42]};
assign col_out_719 = {u_ca_out_719[5:0],u_ca_out_718[23:6], u_ca_out_717[41:24], u_ca_out_716[47:42]};
assign col_out_720 = {u_ca_out_720[5:0],u_ca_out_719[23:6], u_ca_out_718[41:24], u_ca_out_717[47:42]};
assign col_out_721 = {u_ca_out_721[5:0],u_ca_out_720[23:6], u_ca_out_719[41:24], u_ca_out_718[47:42]};
assign col_out_722 = {u_ca_out_722[5:0],u_ca_out_721[23:6], u_ca_out_720[41:24], u_ca_out_719[47:42]};
assign col_out_723 = {u_ca_out_723[5:0],u_ca_out_722[23:6], u_ca_out_721[41:24], u_ca_out_720[47:42]};
assign col_out_724 = {u_ca_out_724[5:0],u_ca_out_723[23:6], u_ca_out_722[41:24], u_ca_out_721[47:42]};
assign col_out_725 = {u_ca_out_725[5:0],u_ca_out_724[23:6], u_ca_out_723[41:24], u_ca_out_722[47:42]};
assign col_out_726 = {u_ca_out_726[5:0],u_ca_out_725[23:6], u_ca_out_724[41:24], u_ca_out_723[47:42]};
assign col_out_727 = {u_ca_out_727[5:0],u_ca_out_726[23:6], u_ca_out_725[41:24], u_ca_out_724[47:42]};
assign col_out_728 = {u_ca_out_728[5:0],u_ca_out_727[23:6], u_ca_out_726[41:24], u_ca_out_725[47:42]};
assign col_out_729 = {u_ca_out_729[5:0],u_ca_out_728[23:6], u_ca_out_727[41:24], u_ca_out_726[47:42]};
assign col_out_730 = {u_ca_out_730[5:0],u_ca_out_729[23:6], u_ca_out_728[41:24], u_ca_out_727[47:42]};
assign col_out_731 = {u_ca_out_731[5:0],u_ca_out_730[23:6], u_ca_out_729[41:24], u_ca_out_728[47:42]};
assign col_out_732 = {u_ca_out_732[5:0],u_ca_out_731[23:6], u_ca_out_730[41:24], u_ca_out_729[47:42]};
assign col_out_733 = {u_ca_out_733[5:0],u_ca_out_732[23:6], u_ca_out_731[41:24], u_ca_out_730[47:42]};
assign col_out_734 = {u_ca_out_734[5:0],u_ca_out_733[23:6], u_ca_out_732[41:24], u_ca_out_731[47:42]};
assign col_out_735 = {u_ca_out_735[5:0],u_ca_out_734[23:6], u_ca_out_733[41:24], u_ca_out_732[47:42]};
assign col_out_736 = {u_ca_out_736[5:0],u_ca_out_735[23:6], u_ca_out_734[41:24], u_ca_out_733[47:42]};
assign col_out_737 = {u_ca_out_737[5:0],u_ca_out_736[23:6], u_ca_out_735[41:24], u_ca_out_734[47:42]};
assign col_out_738 = {u_ca_out_738[5:0],u_ca_out_737[23:6], u_ca_out_736[41:24], u_ca_out_735[47:42]};
assign col_out_739 = {u_ca_out_739[5:0],u_ca_out_738[23:6], u_ca_out_737[41:24], u_ca_out_736[47:42]};
assign col_out_740 = {u_ca_out_740[5:0],u_ca_out_739[23:6], u_ca_out_738[41:24], u_ca_out_737[47:42]};
assign col_out_741 = {u_ca_out_741[5:0],u_ca_out_740[23:6], u_ca_out_739[41:24], u_ca_out_738[47:42]};
assign col_out_742 = {u_ca_out_742[5:0],u_ca_out_741[23:6], u_ca_out_740[41:24], u_ca_out_739[47:42]};
assign col_out_743 = {u_ca_out_743[5:0],u_ca_out_742[23:6], u_ca_out_741[41:24], u_ca_out_740[47:42]};
assign col_out_744 = {u_ca_out_744[5:0],u_ca_out_743[23:6], u_ca_out_742[41:24], u_ca_out_741[47:42]};
assign col_out_745 = {u_ca_out_745[5:0],u_ca_out_744[23:6], u_ca_out_743[41:24], u_ca_out_742[47:42]};
assign col_out_746 = {u_ca_out_746[5:0],u_ca_out_745[23:6], u_ca_out_744[41:24], u_ca_out_743[47:42]};
assign col_out_747 = {u_ca_out_747[5:0],u_ca_out_746[23:6], u_ca_out_745[41:24], u_ca_out_744[47:42]};
assign col_out_748 = {u_ca_out_748[5:0],u_ca_out_747[23:6], u_ca_out_746[41:24], u_ca_out_745[47:42]};
assign col_out_749 = {u_ca_out_749[5:0],u_ca_out_748[23:6], u_ca_out_747[41:24], u_ca_out_746[47:42]};
assign col_out_750 = {u_ca_out_750[5:0],u_ca_out_749[23:6], u_ca_out_748[41:24], u_ca_out_747[47:42]};
assign col_out_751 = {u_ca_out_751[5:0],u_ca_out_750[23:6], u_ca_out_749[41:24], u_ca_out_748[47:42]};
assign col_out_752 = {u_ca_out_752[5:0],u_ca_out_751[23:6], u_ca_out_750[41:24], u_ca_out_749[47:42]};
assign col_out_753 = {u_ca_out_753[5:0],u_ca_out_752[23:6], u_ca_out_751[41:24], u_ca_out_750[47:42]};
assign col_out_754 = {u_ca_out_754[5:0],u_ca_out_753[23:6], u_ca_out_752[41:24], u_ca_out_751[47:42]};
assign col_out_755 = {u_ca_out_755[5:0],u_ca_out_754[23:6], u_ca_out_753[41:24], u_ca_out_752[47:42]};
assign col_out_756 = {u_ca_out_756[5:0],u_ca_out_755[23:6], u_ca_out_754[41:24], u_ca_out_753[47:42]};
assign col_out_757 = {u_ca_out_757[5:0],u_ca_out_756[23:6], u_ca_out_755[41:24], u_ca_out_754[47:42]};
assign col_out_758 = {u_ca_out_758[5:0],u_ca_out_757[23:6], u_ca_out_756[41:24], u_ca_out_755[47:42]};
assign col_out_759 = {u_ca_out_759[5:0],u_ca_out_758[23:6], u_ca_out_757[41:24], u_ca_out_756[47:42]};
assign col_out_760 = {u_ca_out_760[5:0],u_ca_out_759[23:6], u_ca_out_758[41:24], u_ca_out_757[47:42]};
assign col_out_761 = {u_ca_out_761[5:0],u_ca_out_760[23:6], u_ca_out_759[41:24], u_ca_out_758[47:42]};
assign col_out_762 = {u_ca_out_762[5:0],u_ca_out_761[23:6], u_ca_out_760[41:24], u_ca_out_759[47:42]};
assign col_out_763 = {u_ca_out_763[5:0],u_ca_out_762[23:6], u_ca_out_761[41:24], u_ca_out_760[47:42]};
assign col_out_764 = {u_ca_out_764[5:0],u_ca_out_763[23:6], u_ca_out_762[41:24], u_ca_out_761[47:42]};
assign col_out_765 = {u_ca_out_765[5:0],u_ca_out_764[23:6], u_ca_out_763[41:24], u_ca_out_762[47:42]};
assign col_out_766 = {u_ca_out_766[5:0],u_ca_out_765[23:6], u_ca_out_764[41:24], u_ca_out_763[47:42]};
assign col_out_767 = {u_ca_out_767[5:0],u_ca_out_766[23:6], u_ca_out_765[41:24], u_ca_out_764[47:42]};
assign col_out_768 = {u_ca_out_768[5:0],u_ca_out_767[23:6], u_ca_out_766[41:24], u_ca_out_765[47:42]};
assign col_out_769 = {u_ca_out_769[5:0],u_ca_out_768[23:6], u_ca_out_767[41:24], u_ca_out_766[47:42]};
assign col_out_770 = {u_ca_out_770[5:0],u_ca_out_769[23:6], u_ca_out_768[41:24], u_ca_out_767[47:42]};
assign col_out_771 = {u_ca_out_771[5:0],u_ca_out_770[23:6], u_ca_out_769[41:24], u_ca_out_768[47:42]};
assign col_out_772 = {u_ca_out_772[5:0],u_ca_out_771[23:6], u_ca_out_770[41:24], u_ca_out_769[47:42]};
assign col_out_773 = {u_ca_out_773[5:0],u_ca_out_772[23:6], u_ca_out_771[41:24], u_ca_out_770[47:42]};
assign col_out_774 = {u_ca_out_774[5:0],u_ca_out_773[23:6], u_ca_out_772[41:24], u_ca_out_771[47:42]};
assign col_out_775 = {u_ca_out_775[5:0],u_ca_out_774[23:6], u_ca_out_773[41:24], u_ca_out_772[47:42]};
assign col_out_776 = {u_ca_out_776[5:0],u_ca_out_775[23:6], u_ca_out_774[41:24], u_ca_out_773[47:42]};
assign col_out_777 = {u_ca_out_777[5:0],u_ca_out_776[23:6], u_ca_out_775[41:24], u_ca_out_774[47:42]};
assign col_out_778 = {u_ca_out_778[5:0],u_ca_out_777[23:6], u_ca_out_776[41:24], u_ca_out_775[47:42]};
assign col_out_779 = {u_ca_out_779[5:0],u_ca_out_778[23:6], u_ca_out_777[41:24], u_ca_out_776[47:42]};
assign col_out_780 = {u_ca_out_780[5:0],u_ca_out_779[23:6], u_ca_out_778[41:24], u_ca_out_777[47:42]};
assign col_out_781 = {u_ca_out_781[5:0],u_ca_out_780[23:6], u_ca_out_779[41:24], u_ca_out_778[47:42]};
assign col_out_782 = {u_ca_out_782[5:0],u_ca_out_781[23:6], u_ca_out_780[41:24], u_ca_out_779[47:42]};
assign col_out_783 = {u_ca_out_783[5:0],u_ca_out_782[23:6], u_ca_out_781[41:24], u_ca_out_780[47:42]};
assign col_out_784 = {u_ca_out_784[5:0],u_ca_out_783[23:6], u_ca_out_782[41:24], u_ca_out_781[47:42]};
assign col_out_785 = {u_ca_out_785[5:0],u_ca_out_784[23:6], u_ca_out_783[41:24], u_ca_out_782[47:42]};
assign col_out_786 = {u_ca_out_786[5:0],u_ca_out_785[23:6], u_ca_out_784[41:24], u_ca_out_783[47:42]};
assign col_out_787 = {u_ca_out_787[5:0],u_ca_out_786[23:6], u_ca_out_785[41:24], u_ca_out_784[47:42]};
assign col_out_788 = {u_ca_out_788[5:0],u_ca_out_787[23:6], u_ca_out_786[41:24], u_ca_out_785[47:42]};
assign col_out_789 = {u_ca_out_789[5:0],u_ca_out_788[23:6], u_ca_out_787[41:24], u_ca_out_786[47:42]};
assign col_out_790 = {u_ca_out_790[5:0],u_ca_out_789[23:6], u_ca_out_788[41:24], u_ca_out_787[47:42]};
assign col_out_791 = {u_ca_out_791[5:0],u_ca_out_790[23:6], u_ca_out_789[41:24], u_ca_out_788[47:42]};
assign col_out_792 = {u_ca_out_792[5:0],u_ca_out_791[23:6], u_ca_out_790[41:24], u_ca_out_789[47:42]};
assign col_out_793 = {u_ca_out_793[5:0],u_ca_out_792[23:6], u_ca_out_791[41:24], u_ca_out_790[47:42]};
assign col_out_794 = {u_ca_out_794[5:0],u_ca_out_793[23:6], u_ca_out_792[41:24], u_ca_out_791[47:42]};
assign col_out_795 = {u_ca_out_795[5:0],u_ca_out_794[23:6], u_ca_out_793[41:24], u_ca_out_792[47:42]};
assign col_out_796 = {u_ca_out_796[5:0],u_ca_out_795[23:6], u_ca_out_794[41:24], u_ca_out_793[47:42]};
assign col_out_797 = {u_ca_out_797[5:0],u_ca_out_796[23:6], u_ca_out_795[41:24], u_ca_out_794[47:42]};
assign col_out_798 = {u_ca_out_798[5:0],u_ca_out_797[23:6], u_ca_out_796[41:24], u_ca_out_795[47:42]};
assign col_out_799 = {u_ca_out_799[5:0],u_ca_out_798[23:6], u_ca_out_797[41:24], u_ca_out_796[47:42]};
assign col_out_800 = {u_ca_out_800[5:0],u_ca_out_799[23:6], u_ca_out_798[41:24], u_ca_out_797[47:42]};
assign col_out_801 = {u_ca_out_801[5:0],u_ca_out_800[23:6], u_ca_out_799[41:24], u_ca_out_798[47:42]};
assign col_out_802 = {u_ca_out_802[5:0],u_ca_out_801[23:6], u_ca_out_800[41:24], u_ca_out_799[47:42]};
assign col_out_803 = {u_ca_out_803[5:0],u_ca_out_802[23:6], u_ca_out_801[41:24], u_ca_out_800[47:42]};
assign col_out_804 = {u_ca_out_804[5:0],u_ca_out_803[23:6], u_ca_out_802[41:24], u_ca_out_801[47:42]};
assign col_out_805 = {u_ca_out_805[5:0],u_ca_out_804[23:6], u_ca_out_803[41:24], u_ca_out_802[47:42]};
assign col_out_806 = {u_ca_out_806[5:0],u_ca_out_805[23:6], u_ca_out_804[41:24], u_ca_out_803[47:42]};
assign col_out_807 = {u_ca_out_807[5:0],u_ca_out_806[23:6], u_ca_out_805[41:24], u_ca_out_804[47:42]};
assign col_out_808 = {u_ca_out_808[5:0],u_ca_out_807[23:6], u_ca_out_806[41:24], u_ca_out_805[47:42]};
assign col_out_809 = {u_ca_out_809[5:0],u_ca_out_808[23:6], u_ca_out_807[41:24], u_ca_out_806[47:42]};
assign col_out_810 = {u_ca_out_810[5:0],u_ca_out_809[23:6], u_ca_out_808[41:24], u_ca_out_807[47:42]};
assign col_out_811 = {u_ca_out_811[5:0],u_ca_out_810[23:6], u_ca_out_809[41:24], u_ca_out_808[47:42]};
assign col_out_812 = {u_ca_out_812[5:0],u_ca_out_811[23:6], u_ca_out_810[41:24], u_ca_out_809[47:42]};
assign col_out_813 = {u_ca_out_813[5:0],u_ca_out_812[23:6], u_ca_out_811[41:24], u_ca_out_810[47:42]};
assign col_out_814 = {u_ca_out_814[5:0],u_ca_out_813[23:6], u_ca_out_812[41:24], u_ca_out_811[47:42]};
assign col_out_815 = {u_ca_out_815[5:0],u_ca_out_814[23:6], u_ca_out_813[41:24], u_ca_out_812[47:42]};
assign col_out_816 = {u_ca_out_816[5:0],u_ca_out_815[23:6], u_ca_out_814[41:24], u_ca_out_813[47:42]};
assign col_out_817 = {u_ca_out_817[5:0],u_ca_out_816[23:6], u_ca_out_815[41:24], u_ca_out_814[47:42]};
assign col_out_818 = {u_ca_out_818[5:0],u_ca_out_817[23:6], u_ca_out_816[41:24], u_ca_out_815[47:42]};
assign col_out_819 = {u_ca_out_819[5:0],u_ca_out_818[23:6], u_ca_out_817[41:24], u_ca_out_816[47:42]};
assign col_out_820 = {u_ca_out_820[5:0],u_ca_out_819[23:6], u_ca_out_818[41:24], u_ca_out_817[47:42]};
assign col_out_821 = {u_ca_out_821[5:0],u_ca_out_820[23:6], u_ca_out_819[41:24], u_ca_out_818[47:42]};
assign col_out_822 = {u_ca_out_822[5:0],u_ca_out_821[23:6], u_ca_out_820[41:24], u_ca_out_819[47:42]};
assign col_out_823 = {u_ca_out_823[5:0],u_ca_out_822[23:6], u_ca_out_821[41:24], u_ca_out_820[47:42]};
assign col_out_824 = {u_ca_out_824[5:0],u_ca_out_823[23:6], u_ca_out_822[41:24], u_ca_out_821[47:42]};
assign col_out_825 = {u_ca_out_825[5:0],u_ca_out_824[23:6], u_ca_out_823[41:24], u_ca_out_822[47:42]};
assign col_out_826 = {u_ca_out_826[5:0],u_ca_out_825[23:6], u_ca_out_824[41:24], u_ca_out_823[47:42]};
assign col_out_827 = {u_ca_out_827[5:0],u_ca_out_826[23:6], u_ca_out_825[41:24], u_ca_out_824[47:42]};
assign col_out_828 = {u_ca_out_828[5:0],u_ca_out_827[23:6], u_ca_out_826[41:24], u_ca_out_825[47:42]};
assign col_out_829 = {u_ca_out_829[5:0],u_ca_out_828[23:6], u_ca_out_827[41:24], u_ca_out_826[47:42]};
assign col_out_830 = {u_ca_out_830[5:0],u_ca_out_829[23:6], u_ca_out_828[41:24], u_ca_out_827[47:42]};
assign col_out_831 = {u_ca_out_831[5:0],u_ca_out_830[23:6], u_ca_out_829[41:24], u_ca_out_828[47:42]};
assign col_out_832 = {u_ca_out_832[5:0],u_ca_out_831[23:6], u_ca_out_830[41:24], u_ca_out_829[47:42]};
assign col_out_833 = {u_ca_out_833[5:0],u_ca_out_832[23:6], u_ca_out_831[41:24], u_ca_out_830[47:42]};
assign col_out_834 = {u_ca_out_834[5:0],u_ca_out_833[23:6], u_ca_out_832[41:24], u_ca_out_831[47:42]};
assign col_out_835 = {u_ca_out_835[5:0],u_ca_out_834[23:6], u_ca_out_833[41:24], u_ca_out_832[47:42]};
assign col_out_836 = {u_ca_out_836[5:0],u_ca_out_835[23:6], u_ca_out_834[41:24], u_ca_out_833[47:42]};
assign col_out_837 = {u_ca_out_837[5:0],u_ca_out_836[23:6], u_ca_out_835[41:24], u_ca_out_834[47:42]};
assign col_out_838 = {u_ca_out_838[5:0],u_ca_out_837[23:6], u_ca_out_836[41:24], u_ca_out_835[47:42]};
assign col_out_839 = {u_ca_out_839[5:0],u_ca_out_838[23:6], u_ca_out_837[41:24], u_ca_out_836[47:42]};
assign col_out_840 = {u_ca_out_840[5:0],u_ca_out_839[23:6], u_ca_out_838[41:24], u_ca_out_837[47:42]};
assign col_out_841 = {u_ca_out_841[5:0],u_ca_out_840[23:6], u_ca_out_839[41:24], u_ca_out_838[47:42]};
assign col_out_842 = {u_ca_out_842[5:0],u_ca_out_841[23:6], u_ca_out_840[41:24], u_ca_out_839[47:42]};
assign col_out_843 = {u_ca_out_843[5:0],u_ca_out_842[23:6], u_ca_out_841[41:24], u_ca_out_840[47:42]};
assign col_out_844 = {u_ca_out_844[5:0],u_ca_out_843[23:6], u_ca_out_842[41:24], u_ca_out_841[47:42]};
assign col_out_845 = {u_ca_out_845[5:0],u_ca_out_844[23:6], u_ca_out_843[41:24], u_ca_out_842[47:42]};
assign col_out_846 = {u_ca_out_846[5:0],u_ca_out_845[23:6], u_ca_out_844[41:24], u_ca_out_843[47:42]};
assign col_out_847 = {u_ca_out_847[5:0],u_ca_out_846[23:6], u_ca_out_845[41:24], u_ca_out_844[47:42]};
assign col_out_848 = {u_ca_out_848[5:0],u_ca_out_847[23:6], u_ca_out_846[41:24], u_ca_out_845[47:42]};
assign col_out_849 = {u_ca_out_849[5:0],u_ca_out_848[23:6], u_ca_out_847[41:24], u_ca_out_846[47:42]};
assign col_out_850 = {u_ca_out_850[5:0],u_ca_out_849[23:6], u_ca_out_848[41:24], u_ca_out_847[47:42]};
assign col_out_851 = {u_ca_out_851[5:0],u_ca_out_850[23:6], u_ca_out_849[41:24], u_ca_out_848[47:42]};
assign col_out_852 = {u_ca_out_852[5:0],u_ca_out_851[23:6], u_ca_out_850[41:24], u_ca_out_849[47:42]};
assign col_out_853 = {u_ca_out_853[5:0],u_ca_out_852[23:6], u_ca_out_851[41:24], u_ca_out_850[47:42]};
assign col_out_854 = {u_ca_out_854[5:0],u_ca_out_853[23:6], u_ca_out_852[41:24], u_ca_out_851[47:42]};
assign col_out_855 = {u_ca_out_855[5:0],u_ca_out_854[23:6], u_ca_out_853[41:24], u_ca_out_852[47:42]};
assign col_out_856 = {u_ca_out_856[5:0],u_ca_out_855[23:6], u_ca_out_854[41:24], u_ca_out_853[47:42]};
assign col_out_857 = {u_ca_out_857[5:0],u_ca_out_856[23:6], u_ca_out_855[41:24], u_ca_out_854[47:42]};
assign col_out_858 = {u_ca_out_858[5:0],u_ca_out_857[23:6], u_ca_out_856[41:24], u_ca_out_855[47:42]};
assign col_out_859 = {u_ca_out_859[5:0],u_ca_out_858[23:6], u_ca_out_857[41:24], u_ca_out_856[47:42]};
assign col_out_860 = {u_ca_out_860[5:0],u_ca_out_859[23:6], u_ca_out_858[41:24], u_ca_out_857[47:42]};
assign col_out_861 = {u_ca_out_861[5:0],u_ca_out_860[23:6], u_ca_out_859[41:24], u_ca_out_858[47:42]};
assign col_out_862 = {u_ca_out_862[5:0],u_ca_out_861[23:6], u_ca_out_860[41:24], u_ca_out_859[47:42]};
assign col_out_863 = {u_ca_out_863[5:0],u_ca_out_862[23:6], u_ca_out_861[41:24], u_ca_out_860[47:42]};
assign col_out_864 = {u_ca_out_864[5:0],u_ca_out_863[23:6], u_ca_out_862[41:24], u_ca_out_861[47:42]};
assign col_out_865 = {u_ca_out_865[5:0],u_ca_out_864[23:6], u_ca_out_863[41:24], u_ca_out_862[47:42]};
assign col_out_866 = {u_ca_out_866[5:0],u_ca_out_865[23:6], u_ca_out_864[41:24], u_ca_out_863[47:42]};
assign col_out_867 = {u_ca_out_867[5:0],u_ca_out_866[23:6], u_ca_out_865[41:24], u_ca_out_864[47:42]};
assign col_out_868 = {u_ca_out_868[5:0],u_ca_out_867[23:6], u_ca_out_866[41:24], u_ca_out_865[47:42]};
assign col_out_869 = {u_ca_out_869[5:0],u_ca_out_868[23:6], u_ca_out_867[41:24], u_ca_out_866[47:42]};
assign col_out_870 = {u_ca_out_870[5:0],u_ca_out_869[23:6], u_ca_out_868[41:24], u_ca_out_867[47:42]};
assign col_out_871 = {u_ca_out_871[5:0],u_ca_out_870[23:6], u_ca_out_869[41:24], u_ca_out_868[47:42]};
assign col_out_872 = {u_ca_out_872[5:0],u_ca_out_871[23:6], u_ca_out_870[41:24], u_ca_out_869[47:42]};
assign col_out_873 = {u_ca_out_873[5:0],u_ca_out_872[23:6], u_ca_out_871[41:24], u_ca_out_870[47:42]};
assign col_out_874 = {u_ca_out_874[5:0],u_ca_out_873[23:6], u_ca_out_872[41:24], u_ca_out_871[47:42]};
assign col_out_875 = {u_ca_out_875[5:0],u_ca_out_874[23:6], u_ca_out_873[41:24], u_ca_out_872[47:42]};
assign col_out_876 = {u_ca_out_876[5:0],u_ca_out_875[23:6], u_ca_out_874[41:24], u_ca_out_873[47:42]};
assign col_out_877 = {u_ca_out_877[5:0],u_ca_out_876[23:6], u_ca_out_875[41:24], u_ca_out_874[47:42]};
assign col_out_878 = {u_ca_out_878[5:0],u_ca_out_877[23:6], u_ca_out_876[41:24], u_ca_out_875[47:42]};
assign col_out_879 = {u_ca_out_879[5:0],u_ca_out_878[23:6], u_ca_out_877[41:24], u_ca_out_876[47:42]};
assign col_out_880 = {u_ca_out_880[5:0],u_ca_out_879[23:6], u_ca_out_878[41:24], u_ca_out_877[47:42]};
assign col_out_881 = {u_ca_out_881[5:0],u_ca_out_880[23:6], u_ca_out_879[41:24], u_ca_out_878[47:42]};
assign col_out_882 = {u_ca_out_882[5:0],u_ca_out_881[23:6], u_ca_out_880[41:24], u_ca_out_879[47:42]};
assign col_out_883 = {u_ca_out_883[5:0],u_ca_out_882[23:6], u_ca_out_881[41:24], u_ca_out_880[47:42]};
assign col_out_884 = {u_ca_out_884[5:0],u_ca_out_883[23:6], u_ca_out_882[41:24], u_ca_out_881[47:42]};
assign col_out_885 = {u_ca_out_885[5:0],u_ca_out_884[23:6], u_ca_out_883[41:24], u_ca_out_882[47:42]};
assign col_out_886 = {u_ca_out_886[5:0],u_ca_out_885[23:6], u_ca_out_884[41:24], u_ca_out_883[47:42]};
assign col_out_887 = {u_ca_out_887[5:0],u_ca_out_886[23:6], u_ca_out_885[41:24], u_ca_out_884[47:42]};
assign col_out_888 = {u_ca_out_888[5:0],u_ca_out_887[23:6], u_ca_out_886[41:24], u_ca_out_885[47:42]};
assign col_out_889 = {u_ca_out_889[5:0],u_ca_out_888[23:6], u_ca_out_887[41:24], u_ca_out_886[47:42]};
assign col_out_890 = {u_ca_out_890[5:0],u_ca_out_889[23:6], u_ca_out_888[41:24], u_ca_out_887[47:42]};
assign col_out_891 = {u_ca_out_891[5:0],u_ca_out_890[23:6], u_ca_out_889[41:24], u_ca_out_888[47:42]};
assign col_out_892 = {u_ca_out_892[5:0],u_ca_out_891[23:6], u_ca_out_890[41:24], u_ca_out_889[47:42]};
assign col_out_893 = {u_ca_out_893[5:0],u_ca_out_892[23:6], u_ca_out_891[41:24], u_ca_out_890[47:42]};
assign col_out_894 = {u_ca_out_894[5:0],u_ca_out_893[23:6], u_ca_out_892[41:24], u_ca_out_891[47:42]};
assign col_out_895 = {u_ca_out_895[5:0],u_ca_out_894[23:6], u_ca_out_893[41:24], u_ca_out_892[47:42]};
assign col_out_896 = {u_ca_out_896[5:0],u_ca_out_895[23:6], u_ca_out_894[41:24], u_ca_out_893[47:42]};
assign col_out_897 = {u_ca_out_897[5:0],u_ca_out_896[23:6], u_ca_out_895[41:24], u_ca_out_894[47:42]};
assign col_out_898 = {u_ca_out_898[5:0],u_ca_out_897[23:6], u_ca_out_896[41:24], u_ca_out_895[47:42]};
assign col_out_899 = {u_ca_out_899[5:0],u_ca_out_898[23:6], u_ca_out_897[41:24], u_ca_out_896[47:42]};
assign col_out_900 = {u_ca_out_900[5:0],u_ca_out_899[23:6], u_ca_out_898[41:24], u_ca_out_897[47:42]};
assign col_out_901 = {u_ca_out_901[5:0],u_ca_out_900[23:6], u_ca_out_899[41:24], u_ca_out_898[47:42]};
assign col_out_902 = {u_ca_out_902[5:0],u_ca_out_901[23:6], u_ca_out_900[41:24], u_ca_out_899[47:42]};
assign col_out_903 = {u_ca_out_903[5:0],u_ca_out_902[23:6], u_ca_out_901[41:24], u_ca_out_900[47:42]};
assign col_out_904 = {u_ca_out_904[5:0],u_ca_out_903[23:6], u_ca_out_902[41:24], u_ca_out_901[47:42]};
assign col_out_905 = {u_ca_out_905[5:0],u_ca_out_904[23:6], u_ca_out_903[41:24], u_ca_out_902[47:42]};
assign col_out_906 = {u_ca_out_906[5:0],u_ca_out_905[23:6], u_ca_out_904[41:24], u_ca_out_903[47:42]};
assign col_out_907 = {u_ca_out_907[5:0],u_ca_out_906[23:6], u_ca_out_905[41:24], u_ca_out_904[47:42]};
assign col_out_908 = {u_ca_out_908[5:0],u_ca_out_907[23:6], u_ca_out_906[41:24], u_ca_out_905[47:42]};
assign col_out_909 = {u_ca_out_909[5:0],u_ca_out_908[23:6], u_ca_out_907[41:24], u_ca_out_906[47:42]};
assign col_out_910 = {u_ca_out_910[5:0],u_ca_out_909[23:6], u_ca_out_908[41:24], u_ca_out_907[47:42]};
assign col_out_911 = {u_ca_out_911[5:0],u_ca_out_910[23:6], u_ca_out_909[41:24], u_ca_out_908[47:42]};
assign col_out_912 = {u_ca_out_912[5:0],u_ca_out_911[23:6], u_ca_out_910[41:24], u_ca_out_909[47:42]};
assign col_out_913 = {u_ca_out_913[5:0],u_ca_out_912[23:6], u_ca_out_911[41:24], u_ca_out_910[47:42]};
assign col_out_914 = {u_ca_out_914[5:0],u_ca_out_913[23:6], u_ca_out_912[41:24], u_ca_out_911[47:42]};
assign col_out_915 = {u_ca_out_915[5:0],u_ca_out_914[23:6], u_ca_out_913[41:24], u_ca_out_912[47:42]};
assign col_out_916 = {u_ca_out_916[5:0],u_ca_out_915[23:6], u_ca_out_914[41:24], u_ca_out_913[47:42]};
assign col_out_917 = {u_ca_out_917[5:0],u_ca_out_916[23:6], u_ca_out_915[41:24], u_ca_out_914[47:42]};
assign col_out_918 = {u_ca_out_918[5:0],u_ca_out_917[23:6], u_ca_out_916[41:24], u_ca_out_915[47:42]};
assign col_out_919 = {u_ca_out_919[5:0],u_ca_out_918[23:6], u_ca_out_917[41:24], u_ca_out_916[47:42]};
assign col_out_920 = {u_ca_out_920[5:0],u_ca_out_919[23:6], u_ca_out_918[41:24], u_ca_out_917[47:42]};
assign col_out_921 = {u_ca_out_921[5:0],u_ca_out_920[23:6], u_ca_out_919[41:24], u_ca_out_918[47:42]};
assign col_out_922 = {u_ca_out_922[5:0],u_ca_out_921[23:6], u_ca_out_920[41:24], u_ca_out_919[47:42]};
assign col_out_923 = {u_ca_out_923[5:0],u_ca_out_922[23:6], u_ca_out_921[41:24], u_ca_out_920[47:42]};
assign col_out_924 = {u_ca_out_924[5:0],u_ca_out_923[23:6], u_ca_out_922[41:24], u_ca_out_921[47:42]};
assign col_out_925 = {u_ca_out_925[5:0],u_ca_out_924[23:6], u_ca_out_923[41:24], u_ca_out_922[47:42]};
assign col_out_926 = {u_ca_out_926[5:0],u_ca_out_925[23:6], u_ca_out_924[41:24], u_ca_out_923[47:42]};
assign col_out_927 = {u_ca_out_927[5:0],u_ca_out_926[23:6], u_ca_out_925[41:24], u_ca_out_924[47:42]};
assign col_out_928 = {u_ca_out_928[5:0],u_ca_out_927[23:6], u_ca_out_926[41:24], u_ca_out_925[47:42]};
assign col_out_929 = {u_ca_out_929[5:0],u_ca_out_928[23:6], u_ca_out_927[41:24], u_ca_out_926[47:42]};
assign col_out_930 = {u_ca_out_930[5:0],u_ca_out_929[23:6], u_ca_out_928[41:24], u_ca_out_927[47:42]};
assign col_out_931 = {u_ca_out_931[5:0],u_ca_out_930[23:6], u_ca_out_929[41:24], u_ca_out_928[47:42]};
assign col_out_932 = {u_ca_out_932[5:0],u_ca_out_931[23:6], u_ca_out_930[41:24], u_ca_out_929[47:42]};
assign col_out_933 = {u_ca_out_933[5:0],u_ca_out_932[23:6], u_ca_out_931[41:24], u_ca_out_930[47:42]};
assign col_out_934 = {u_ca_out_934[5:0],u_ca_out_933[23:6], u_ca_out_932[41:24], u_ca_out_931[47:42]};
assign col_out_935 = {u_ca_out_935[5:0],u_ca_out_934[23:6], u_ca_out_933[41:24], u_ca_out_932[47:42]};
assign col_out_936 = {u_ca_out_936[5:0],u_ca_out_935[23:6], u_ca_out_934[41:24], u_ca_out_933[47:42]};
assign col_out_937 = {u_ca_out_937[5:0],u_ca_out_936[23:6], u_ca_out_935[41:24], u_ca_out_934[47:42]};
assign col_out_938 = {u_ca_out_938[5:0],u_ca_out_937[23:6], u_ca_out_936[41:24], u_ca_out_935[47:42]};
assign col_out_939 = {u_ca_out_939[5:0],u_ca_out_938[23:6], u_ca_out_937[41:24], u_ca_out_936[47:42]};
assign col_out_940 = {u_ca_out_940[5:0],u_ca_out_939[23:6], u_ca_out_938[41:24], u_ca_out_937[47:42]};
assign col_out_941 = {u_ca_out_941[5:0],u_ca_out_940[23:6], u_ca_out_939[41:24], u_ca_out_938[47:42]};
assign col_out_942 = {u_ca_out_942[5:0],u_ca_out_941[23:6], u_ca_out_940[41:24], u_ca_out_939[47:42]};
assign col_out_943 = {u_ca_out_943[5:0],u_ca_out_942[23:6], u_ca_out_941[41:24], u_ca_out_940[47:42]};
assign col_out_944 = {u_ca_out_944[5:0],u_ca_out_943[23:6], u_ca_out_942[41:24], u_ca_out_941[47:42]};
assign col_out_945 = {u_ca_out_945[5:0],u_ca_out_944[23:6], u_ca_out_943[41:24], u_ca_out_942[47:42]};
assign col_out_946 = {u_ca_out_946[5:0],u_ca_out_945[23:6], u_ca_out_944[41:24], u_ca_out_943[47:42]};
assign col_out_947 = {u_ca_out_947[5:0],u_ca_out_946[23:6], u_ca_out_945[41:24], u_ca_out_944[47:42]};
assign col_out_948 = {u_ca_out_948[5:0],u_ca_out_947[23:6], u_ca_out_946[41:24], u_ca_out_945[47:42]};
assign col_out_949 = {u_ca_out_949[5:0],u_ca_out_948[23:6], u_ca_out_947[41:24], u_ca_out_946[47:42]};
assign col_out_950 = {u_ca_out_950[5:0],u_ca_out_949[23:6], u_ca_out_948[41:24], u_ca_out_947[47:42]};
assign col_out_951 = {u_ca_out_951[5:0],u_ca_out_950[23:6], u_ca_out_949[41:24], u_ca_out_948[47:42]};
assign col_out_952 = {u_ca_out_952[5:0],u_ca_out_951[23:6], u_ca_out_950[41:24], u_ca_out_949[47:42]};
assign col_out_953 = {u_ca_out_953[5:0],u_ca_out_952[23:6], u_ca_out_951[41:24], u_ca_out_950[47:42]};
assign col_out_954 = {u_ca_out_954[5:0],u_ca_out_953[23:6], u_ca_out_952[41:24], u_ca_out_951[47:42]};
assign col_out_955 = {u_ca_out_955[5:0],u_ca_out_954[23:6], u_ca_out_953[41:24], u_ca_out_952[47:42]};
assign col_out_956 = {u_ca_out_956[5:0],u_ca_out_955[23:6], u_ca_out_954[41:24], u_ca_out_953[47:42]};
assign col_out_957 = {u_ca_out_957[5:0],u_ca_out_956[23:6], u_ca_out_955[41:24], u_ca_out_954[47:42]};
assign col_out_958 = {u_ca_out_958[5:0],u_ca_out_957[23:6], u_ca_out_956[41:24], u_ca_out_955[47:42]};
assign col_out_959 = {u_ca_out_959[5:0],u_ca_out_958[23:6], u_ca_out_957[41:24], u_ca_out_956[47:42]};
assign col_out_960 = {u_ca_out_960[5:0],u_ca_out_959[23:6], u_ca_out_958[41:24], u_ca_out_957[47:42]};
assign col_out_961 = {u_ca_out_961[5:0],u_ca_out_960[23:6], u_ca_out_959[41:24], u_ca_out_958[47:42]};
assign col_out_962 = {u_ca_out_962[5:0],u_ca_out_961[23:6], u_ca_out_960[41:24], u_ca_out_959[47:42]};
assign col_out_963 = {u_ca_out_963[5:0],u_ca_out_962[23:6], u_ca_out_961[41:24], u_ca_out_960[47:42]};
assign col_out_964 = {u_ca_out_964[5:0],u_ca_out_963[23:6], u_ca_out_962[41:24], u_ca_out_961[47:42]};
assign col_out_965 = {u_ca_out_965[5:0],u_ca_out_964[23:6], u_ca_out_963[41:24], u_ca_out_962[47:42]};
assign col_out_966 = {u_ca_out_966[5:0],u_ca_out_965[23:6], u_ca_out_964[41:24], u_ca_out_963[47:42]};
assign col_out_967 = {u_ca_out_967[5:0],u_ca_out_966[23:6], u_ca_out_965[41:24], u_ca_out_964[47:42]};
assign col_out_968 = {u_ca_out_968[5:0],u_ca_out_967[23:6], u_ca_out_966[41:24], u_ca_out_965[47:42]};
assign col_out_969 = {u_ca_out_969[5:0],u_ca_out_968[23:6], u_ca_out_967[41:24], u_ca_out_966[47:42]};
assign col_out_970 = {u_ca_out_970[5:0],u_ca_out_969[23:6], u_ca_out_968[41:24], u_ca_out_967[47:42]};
assign col_out_971 = {u_ca_out_971[5:0],u_ca_out_970[23:6], u_ca_out_969[41:24], u_ca_out_968[47:42]};
assign col_out_972 = {u_ca_out_972[5:0],u_ca_out_971[23:6], u_ca_out_970[41:24], u_ca_out_969[47:42]};
assign col_out_973 = {u_ca_out_973[5:0],u_ca_out_972[23:6], u_ca_out_971[41:24], u_ca_out_970[47:42]};
assign col_out_974 = {u_ca_out_974[5:0],u_ca_out_973[23:6], u_ca_out_972[41:24], u_ca_out_971[47:42]};
assign col_out_975 = {u_ca_out_975[5:0],u_ca_out_974[23:6], u_ca_out_973[41:24], u_ca_out_972[47:42]};
assign col_out_976 = {u_ca_out_976[5:0],u_ca_out_975[23:6], u_ca_out_974[41:24], u_ca_out_973[47:42]};
assign col_out_977 = {u_ca_out_977[5:0],u_ca_out_976[23:6], u_ca_out_975[41:24], u_ca_out_974[47:42]};
assign col_out_978 = {u_ca_out_978[5:0],u_ca_out_977[23:6], u_ca_out_976[41:24], u_ca_out_975[47:42]};
assign col_out_979 = {u_ca_out_979[5:0],u_ca_out_978[23:6], u_ca_out_977[41:24], u_ca_out_976[47:42]};
assign col_out_980 = {u_ca_out_980[5:0],u_ca_out_979[23:6], u_ca_out_978[41:24], u_ca_out_977[47:42]};
assign col_out_981 = {u_ca_out_981[5:0],u_ca_out_980[23:6], u_ca_out_979[41:24], u_ca_out_978[47:42]};
assign col_out_982 = {u_ca_out_982[5:0],u_ca_out_981[23:6], u_ca_out_980[41:24], u_ca_out_979[47:42]};
assign col_out_983 = {u_ca_out_983[5:0],u_ca_out_982[23:6], u_ca_out_981[41:24], u_ca_out_980[47:42]};
assign col_out_984 = {u_ca_out_984[5:0],u_ca_out_983[23:6], u_ca_out_982[41:24], u_ca_out_981[47:42]};
assign col_out_985 = {u_ca_out_985[5:0],u_ca_out_984[23:6], u_ca_out_983[41:24], u_ca_out_982[47:42]};
assign col_out_986 = {u_ca_out_986[5:0],u_ca_out_985[23:6], u_ca_out_984[41:24], u_ca_out_983[47:42]};
assign col_out_987 = {u_ca_out_987[5:0],u_ca_out_986[23:6], u_ca_out_985[41:24], u_ca_out_984[47:42]};
assign col_out_988 = {u_ca_out_988[5:0],u_ca_out_987[23:6], u_ca_out_986[41:24], u_ca_out_985[47:42]};
assign col_out_989 = {u_ca_out_989[5:0],u_ca_out_988[23:6], u_ca_out_987[41:24], u_ca_out_986[47:42]};
assign col_out_990 = {u_ca_out_990[5:0],u_ca_out_989[23:6], u_ca_out_988[41:24], u_ca_out_987[47:42]};
assign col_out_991 = {u_ca_out_991[5:0],u_ca_out_990[23:6], u_ca_out_989[41:24], u_ca_out_988[47:42]};
assign col_out_992 = {u_ca_out_992[5:0],u_ca_out_991[23:6], u_ca_out_990[41:24], u_ca_out_989[47:42]};
assign col_out_993 = {u_ca_out_993[5:0],u_ca_out_992[23:6], u_ca_out_991[41:24], u_ca_out_990[47:42]};
assign col_out_994 = {u_ca_out_994[5:0],u_ca_out_993[23:6], u_ca_out_992[41:24], u_ca_out_991[47:42]};
assign col_out_995 = {u_ca_out_995[5:0],u_ca_out_994[23:6], u_ca_out_993[41:24], u_ca_out_992[47:42]};
assign col_out_996 = {u_ca_out_996[5:0],u_ca_out_995[23:6], u_ca_out_994[41:24], u_ca_out_993[47:42]};
assign col_out_997 = {u_ca_out_997[5:0],u_ca_out_996[23:6], u_ca_out_995[41:24], u_ca_out_994[47:42]};
assign col_out_998 = {u_ca_out_998[5:0],u_ca_out_997[23:6], u_ca_out_996[41:24], u_ca_out_995[47:42]};
assign col_out_999 = {u_ca_out_999[5:0],u_ca_out_998[23:6], u_ca_out_997[41:24], u_ca_out_996[47:42]};
assign col_out_1000 = {u_ca_out_1000[5:0],u_ca_out_999[23:6], u_ca_out_998[41:24], u_ca_out_997[47:42]};
assign col_out_1001 = {u_ca_out_1001[5:0],u_ca_out_1000[23:6], u_ca_out_999[41:24], u_ca_out_998[47:42]};
assign col_out_1002 = {u_ca_out_1002[5:0],u_ca_out_1001[23:6], u_ca_out_1000[41:24], u_ca_out_999[47:42]};
assign col_out_1003 = {u_ca_out_1003[5:0],u_ca_out_1002[23:6], u_ca_out_1001[41:24], u_ca_out_1000[47:42]};
assign col_out_1004 = {u_ca_out_1004[5:0],u_ca_out_1003[23:6], u_ca_out_1002[41:24], u_ca_out_1001[47:42]};
assign col_out_1005 = {u_ca_out_1005[5:0],u_ca_out_1004[23:6], u_ca_out_1003[41:24], u_ca_out_1002[47:42]};
assign col_out_1006 = {u_ca_out_1006[5:0],u_ca_out_1005[23:6], u_ca_out_1004[41:24], u_ca_out_1003[47:42]};
assign col_out_1007 = {u_ca_out_1007[5:0],u_ca_out_1006[23:6], u_ca_out_1005[41:24], u_ca_out_1004[47:42]};
assign col_out_1008 = {u_ca_out_1008[5:0],u_ca_out_1007[23:6], u_ca_out_1006[41:24], u_ca_out_1005[47:42]};
assign col_out_1009 = {u_ca_out_1009[5:0],u_ca_out_1008[23:6], u_ca_out_1007[41:24], u_ca_out_1006[47:42]};
assign col_out_1010 = {u_ca_out_1010[5:0],u_ca_out_1009[23:6], u_ca_out_1008[41:24], u_ca_out_1007[47:42]};
assign col_out_1011 = {u_ca_out_1011[5:0],u_ca_out_1010[23:6], u_ca_out_1009[41:24], u_ca_out_1008[47:42]};
assign col_out_1012 = {u_ca_out_1012[5:0],u_ca_out_1011[23:6], u_ca_out_1010[41:24], u_ca_out_1009[47:42]};
assign col_out_1013 = {u_ca_out_1013[5:0],u_ca_out_1012[23:6], u_ca_out_1011[41:24], u_ca_out_1010[47:42]};
assign col_out_1014 = {u_ca_out_1014[5:0],u_ca_out_1013[23:6], u_ca_out_1012[41:24], u_ca_out_1011[47:42]};
assign col_out_1015 = {u_ca_out_1015[5:0],u_ca_out_1014[23:6], u_ca_out_1013[41:24], u_ca_out_1012[47:42]};
assign col_out_1016 = {u_ca_out_1016[5:0],u_ca_out_1015[23:6], u_ca_out_1014[41:24], u_ca_out_1013[47:42]};
assign col_out_1017 = {u_ca_out_1017[5:0],u_ca_out_1016[23:6], u_ca_out_1015[41:24], u_ca_out_1014[47:42]};
assign col_out_1018 = {u_ca_out_1018[5:0],u_ca_out_1017[23:6], u_ca_out_1016[41:24], u_ca_out_1015[47:42]};
assign col_out_1019 = {u_ca_out_1019[5:0],u_ca_out_1018[23:6], u_ca_out_1017[41:24], u_ca_out_1016[47:42]};
assign col_out_1020 = {u_ca_out_1020[5:0],u_ca_out_1019[23:6], u_ca_out_1018[41:24], u_ca_out_1017[47:42]};
assign col_out_1021 = {u_ca_out_1021[5:0],u_ca_out_1020[23:6], u_ca_out_1019[41:24], u_ca_out_1018[47:42]};
assign col_out_1022 = {u_ca_out_1022[5:0],u_ca_out_1021[23:6], u_ca_out_1020[41:24], u_ca_out_1019[47:42]};
assign col_out_1023 = {u_ca_out_1023[5:0],u_ca_out_1022[23:6], u_ca_out_1021[41:24], u_ca_out_1020[47:42]};
assign col_out_1024 = {u_ca_out_1024[5:0],u_ca_out_1023[23:6], u_ca_out_1022[41:24], u_ca_out_1021[47:42]};
assign col_out_1025 = {u_ca_out_1025[5:0],u_ca_out_1024[23:6], u_ca_out_1023[41:24], u_ca_out_1022[47:42]};
assign col_out_1026 = {u_ca_out_1026[5:0],u_ca_out_1025[23:6], u_ca_out_1024[41:24], u_ca_out_1023[47:42]};
assign col_out_1027 = {{6{1'b0}}, u_ca_out_1026[23:6], u_ca_out_1025[41:24], u_ca_out_1024[47:42]};
assign col_out_1028 = {{24{1'b0}}, u_ca_out_1026[41:24], u_ca_out_1025[47:42]};
assign col_out_1029 = {{42{1'b0}}, u_ca_out_1026[47:42]};

//---------------------------------------------------------


endmodule
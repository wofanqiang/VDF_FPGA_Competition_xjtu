module xpb_5_860
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h7fb489ba0dff27455772d26a2a52ec28a95e6a3029a715b75933911d2a47ae91bce3dac85fb282edcb9a55a88231f28589221999195e53cc21017952132be43cd27b23bcb62d9d072d8e5ef5afc6048de974f5352e99fde10e252a9d0ed16987458214a77c054b9852cf58529982e6ee29ef5d346f32df3ce5d2e44aedc065a2;
    5'b00010 : xpb = 1024'h4ebbce1e5a1019c1e3e02cfd444b90ffe146d12f7dd68af7348a68e4a18cb01b767f3817f53e874cf7d66c0a2105d440ae2a0b4c1009d74c9163b345eb8553c830a712cabcca3cc94882bb48c6b044eadee4f0d1d0adceb166bdc33f6378307c5bfc972547419ea31edec9c63b35a7b30504db868e1a614985364d91529e64d9;
    5'b00011 : xpb = 1024'h1dc31282a6210c3e704d87905e4435d7192f382ed20600370fe140ac18d1b1a5301a95678aca8bac2412826bbfd9b5fbd331fcff06b55acd01c5ed39c3dec3538ed301d8c366dc8b6377179bdd9a8547d454ec6e72c19f81bf565be1b81ef771727719a3127df1adeaee3b39dce86877e01a59d8ad01e3562499b6d7b77c6410;
    5'b00100 : xpb = 1024'h9d779c3cb4203383c7c059fa889721ffc28da25efbad15ee6914d1c943196036ecfe702fea7d0e99efacd814420ba8815c5416982013ae9922c7668bd70aa790614e259579947992910576918d6089d5bdc9e1a3a15b9d62cd7b867ec6f060f8b7f92e4a8e833d463dbd938c766b4f660a09b70d1c34c2930a6c9b22a53cc9b2;
    5'b00101 : xpb = 1024'h6c7ee0a100312600542db48da28fc6d6fa76095e4fdc8b2e446ba990ba5e61c0a699cd7f800912f91be8ee75e0df8a3c815c084b16bf32199329a07faf64171bbf7a14a380311954abf9d2e4a44aca32b339dd40436f6e3326141f211b9727edce73b0c859bf905109cd0500181e102ae51f355f3b1c449fa9d004690a1ac8e9;
    5'b00110 : xpb = 1024'h3b8625054c42187ce09b0f20bc886bae325e705da40c006e1fc2815831a3634a60352acf15951758482504d77fb36bf7a663f9fe0d6ab59a038bda7387bd86a71da603b186cdb916c6ee2f37bb350a8fa8a9d8dce5833f037eacb7c3703deee2e4ee334624fbe35bd5dc7673b9d0d0efc034b3b15a03c6ac49336daf6ef8c820;
    5'b00111 : xpb = 1024'ha8d696998530af96d0869b3d68110856a46d75cf83b75adfb19591fa8e864d419d0881eab211bb774611b391e874db2cb6bebb10416391a73ee14676016f6327bd1f2bf8d6a58d8e1e28b8ad21f4aec9e19d47987970fd3d7455065c4e4b5d7fb68b5c3f0383666a1ebe7e75b8391b49b4a320378eb48b8e896d6f5d3d6c757;
    5'b01000 : xpb = 1024'h8a41f323a652323ec47b3c1e00d3fcae13a5418d21e28b65544cea3cd3301365d6b462e70ad39ea53ffb70e1a0b94038548e054a1d748ce694ef8db97342da6f4e4d167c4397f5e00f70ea8081e54f7a878ec9aeb6310db4e56a7b02d3b61f5f40eaca6b6c3d81fef4bb4039f50678a2c5398f37e81e27f5ce69bb40c1972cf9;
    5'b01001 : xpb = 1024'h59493787f26324bb50e896b11acca1854b8da88c761200a52fa3c2044a7514ef904fc036a05fa3046c3787433f8d21f37995f6fd142010670551c7ad4b9c49faac79058a4a3495a22a6546d398cf8fd77cfec54b5844de853e0313a5285ce65457654ce93779d509c0cab1ad96b93967a04f0d8a0705aa026dcd248726752c30;
    5'b01010 : xpb = 1024'h28507bec3e741737dd55f14434c5465c83760f8bca4175e50afa99cbc1ba167949eb1d8635eba76398739da4de6103ae9e9de8b00acb93e775b401a123f5b9860aa4f49850d135644559a326afb9d034726ec0e7fa58af55969bac477d03ad496ddfcf6702b628148cda2321386bfa2c7b648bdc25ed2c0f0d308dcd8b532b67;
    5'b01011 : xpb = 1024'ha80505a64c733e7d34c8c3ae5f1832852cd479bbf3e88b9c642e2ae8ec01c50b06cef84e959e2a51640df34d6092f63427c002492429e7b396b57af337219dc2dd20185506fed26b72e8021c5f7fd4c25be3b61d28f2ad36a4c0d6e48bd516d0b361e40e7ebb73acdfa97b73d1eee11aa553e91095200b4bf303721879139109;
    5'b01100 : xpb = 1024'h770c4a0a988430f9c1361e417910d75c64bce0bb481800dc3f8502b06346c694c06a559e2b2a2eb0904a09aeff66d7ef4cc7f3fc1ad56b340717b4e70f7b0d4e3b4c07630d9b722d8ddc5e6f766a151f5153b1b9cb067e06fd596f86e07bddc5c9dc668c49f7c6b7abb8ece773a1a1df80696762b4078d589266db5eddf19040;
    5'b01101 : xpb = 1024'h46138e6ee49523764da378d493097c339ca547ba9c47761c1adbda77da8bc81e7a05b2edc0b6330fbc8620109e3ab9aa71cfe5af1180eeb47779eedae7d47cd99977f671143811efa8d0bac28d54557c46c3ad566d1a4ed755f208293522a4bae056e90a153419c277c85e5b155462a45b7ee5b4d2ef0f6531ca44a542cf8f77;
    5'b01110 : xpb = 1024'h151ad2d330a615f2da10d367ad02210ad48daeb9f076eb5bf632b23f51d0c9a833a1103d5642376ee8c236723d0e9b6596d7d762082c7234e7dc28cec02dec64f7a3e57f1ad4b1b1c3c51715a43e95d93c33a8f30f2e1fa7ae8aa0cb89c96baff6d16b87e0706ccd43d7cfceb707236936946406f1d69171d12dadeba7ad8eae;
    5'b01111 : xpb = 1024'h94cf5c8d3ea53d383183a5d1d7550d337dec18ea1a1e01134f66435c7c187839f084eb05b5f4ba5cb45c8c1abf408deb1ff9f0fb218ac60108dda220d359d0a1ca1f093bd1024eb8f153760b54049a6725a89e283dc81d88bcafcb68989ad5373c53802f5c75b86596a72821508a0a576083c13b610970aeb7009236956df450;
    5'b10000 : xpb = 1024'h63d6a0f18ab62fb4bdf10064f14db20ab5d47fe96e4d76532abd1b23f35d79c3aa2048554b80bebbe098a27c5e146fa64501e2ae18364981793fdc14abb3402d284af849d79eee7b0c47d25e6aeedac41b1899c4dfdbee591548640aed419c2c52ce02ad27b20b7062b69994f23ccb1c3b993f8d7ff0f2bb5663fb7cfa4bf387;
    5'b10001 : xpb = 1024'h32dde555d6c722314a5e5af80b4656e1edbce6e8c27ceb930613f2eb6aa27b4d63bba5a4e10cc31b0cd4b8ddfce851616a09d4610ee1cd01e9a21608840cafb88676e757de3b8e3d273c2eb181d91b211088956181efbf296de0fcad41e863216948852af2ee5e7b2ec60b0893ef8be116aebddf9ed874c7f5c764c35f29f2be;
    5'b10010 : xpb = 1024'h1e529ba22d814add6cbb58b253efbb925a54de816ac60d2e16acab2e1e77cd71d5702f47698c77a3910cf3f9bbc331c8f11c614058d50825a044ffc5c661f43e4a2d665e4d82dff42308b0498c35b7e05f890fe24038ff9c679954f968f2a167fc307a8be2ab185fad57c7c35a24ca5f1c43c31bdbff6d4952ace09c407f1f5;
    5'b10011 : xpb = 1024'h8199b37430d73bf32e3e87f54f91e7e1cf03b8184053768a3a9e5bd00c2f2b68da3addbcd64b4a6804ab24e81dee25a21833dfad1eeba44e7b05c94e6f920380b71dfa229b05cb066fbee9fa4889600bef6d8633529d8ddad49ebfeca560939dc5451c503a2ffd1e4da4d4cecf2533941bb399662cf2d6117afdb254b1c85797;
    5'b10100 : xpb = 1024'h50a0f7d87ce82e6fbaabe288698a8cb906ec1f179482ebca15f5339783742cf293d63b0c6bd74ec730e73b49bcc2075d3d3bd160159727ceeb68034247eb730c1549e930a1a26ac88ab3464d5f73a068e4dd81cff4b15eab2d37588efa075a92dbbf9ece056c502919b4464270d7f458f6c917b84bda581e1a611b9b16a656ce;
    5'b10101 : xpb = 1024'h1fa83c3cc8f920ec47193d1b838331903ed48616e8b26109f14c0b5efab92e7c4d71985c016353265d2351ab5b95e9186243c3130c42ab4f5bca3d362044e2977375d83ea83f0a8aa5a7a2a0765de0c5da4d7d6c96c52f7b85cff1314eae2187f23a214bd0a8a333e5c3b7b6128ab51dd1de960a6ac1da2ab9c484e17b845605;
    5'b10110 : xpb = 1024'h9f5cc5f6d6f848319e8c0f85add61db8e832f047125976c14a7f9c7c2500dd0e0a5573246115d61428bda753ddc7db9deb65dcac25a0ff1b7ccbb6883370c6d445f0fbfb5e6ca791d33601962623e553c3c272a1c55f2d5c93f51bce5d7f8b0f37bc35f34cadeecc38931008ac0d9c0bfbcdf33ed9f4b9679f97692c6944bba7;
    5'b10111 : xpb = 1024'h6e640a5b23093aae2af96a18c7cec290201b57466688ec0125d674439c45de97c3f0d073f6a1da7354f9bdb57c9bbd59106dce5f1c4c829bed2df07c0bca365fa41ceb0965094753ee2a5de93d0e25b0b9326e3e6772fe2cec8db470b22652044e36b87117ea41d704a2817c4dc05cd0d6e37190f8dc3b743efad272ce22bade;
    5'b11000 : xpb = 1024'h3d6b4ebf6f1a2d2ab766c4abe1c767675803be45bab86141012d4c0b138ae0217d8c2dc38c2dded28135d4171b6f9f143575c01212f8061c5d902a6fe423a5eb0248da176ba5e716091eba3c53f8660daea269db0986cefd45264d1306cd18f964b13aeee32694e1d0b1f2efef731d95b1f8efe317c3bd80de5e3bb93300ba15;
    5'b11001 : xpb = 1024'hc729323bb2b1fa743d41f3efbc00c3e8fec25450ee7d680dc8423d28acfe1ab37278b1321b9e331ad71ea78ba4380cf5a7db1c509a3899ccdf26463bc7d15766074c925724286d82413168f6ae2a66aa4126577ab9a9fcd9dbee5b55b73dfee7b2bbd6cae62e7ec9cc164639125de5a8d0e6e3536ab3f8d7dc1a4ff97deb94c;
    5'b11010 : xpb = 1024'h8c271cddc92a46ec9b46f1a92612f867394a8f75388eec3835b7b4efb517903cf40b65db816c661f790c40213c757354e39fcb5e2301dd68eef3ddb5cfa8f9b332efece2287023df51a175851aa8aaf88d875aacda349daeabe410526a454975c0add2142a683384ef90bcb62aa8c548b6fdcb69a5de1eca6394894a859f1eee;
    5'b11011 : xpb = 1024'h5b2e6142153b396927b44c3c400b9d3e7132f6748cbe6178110e8cb72c5c91c6ada6c32b16f86a7ea5485682db49551008a7bd1119ad60e95f5617a9a802693e911bdbf02f0cc3a16c95d1d83192eb5582f756497c486e7f047ca8f4beec106ad7285491f5a4868fbba02e29cc5b860d921349bbc4c5a0d702f7f290ea7d1e25;
    5'b11100 : xpb = 1024'h2a35a5a6614c2be5b421a6cf5a044215a91b5d73e0edd6b7ec65647ea3a193506742207aac846eddd1846ce47a1d36cb2dafaec41058e469cfb8519d805bd8c9ef47cafe35a96363878a2e2b487d2bb2786751e61e5c3f4f5d1541971392d75feda2d70fc0e0d99a87af9f9d6e0e46d26d28c80de3ad22e3a25b5bd74f5b1d5c;
    5'b11101 : xpb = 1024'ha9ea2f606f4b532b0b94793984572e3e5279c7a40a94ec6f4598f59bcde941e22425fb430c36f1cb9d1ec28cfc4f2950b6d1c85d29b73835f0b9caef9387bd06c1c2eebaebd7006ab5188d20f843304061dc471b4cf63d306b3a6c34226440e73324ebb73ce62532da7ef7f007912dc09718254252e00220882e40223d1b82fe;
    5'b11110 : xpb = 1024'h78f173c4bb5c45a79801d3cc9e4fd3158a622ea35ec461af20efcd63452e436bddc15892a1c2f62ac95ad8ee9b230b0bdbd9ba102062bbb6611c04e36be12c921feeddc8f273a02cd00ce9740f2d709d574c42b7ef0a0e00c3d304d6770b07dc499f6e350822783da68e6963a943ee85722da39471c7842d2791a968a1f98235;
    5'b11111 : xpb = 1024'h47f8b829076d3824246f2e5fb84877ecc24a95a2b2f3d6eefc46a52abc7344f5975cb5e2374efa89f596ef5039f6ecc700e1abc3170e3f36d17e3ed7443a9c1d7e1accd6f9103feeeb0145c72617b0fa4cbc3e54911dded11c6b9d78cbb1ced16019f0b2d35ecb48729ddad74af6af4a4d4321e690af0639c6f512af06d7816c;
    endcase
end

endmodule

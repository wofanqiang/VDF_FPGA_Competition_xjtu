module xpb_5_375
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h541319b3268d9a0bfe6b719fe04b305996f19388bc59bbe770046dda4bcf88dfdff6fdbdfc9a8d5d10c4352a1729d3e46dc1826ccb0aa67475523520c9ded23ceaa901888937f2d37fdc48176c5899a59453214fcd28ac636858e5464c452be74e9e3d1124d3952111b59e958bb3c71c4788016d7eda4b7d424dcb3e04b45039;
    5'b00010 : xpb = 1024'ha82633664d1b3417fcd6e33fc09660b32de3271178b377cee008dbb4979f11bfbfedfb7bf9351aba21886a542e53a7c8db8304d996154ce8eaa46a4193bda479d5520311126fe5a6ffb8902ed8b1334b28a6429f9a5158c6d0b1ca8c988a57ce9d3c7a2249a72a42236b3d2b17678e388f1002dafdb496fa849b967c0968a072;
    5'b00011 : xpb = 1024'h4b8c07c3b1ba995b303cdd08908749bb535eb7695f95933ed2309039306bed979c9c7bc12ba9298892ee6037621f6ae2e52a5f603e6d2311af57600422ca02054babcfeaec16db356cfad5a3ac2e08bfc8f46a56daf3d819837e1dd82aa4e123bcd32509bdb1c6d5ae60f4e1ab4b2f2b87be25662c4385478079e6b5853a8a40;
    5'b00100 : xpb = 1024'h9f9f2176d84833672ea84ea870d27a14ea504af21bef4f264234fe137c3b76777c93797f2843b6e5a3b2956179493ec752ebe1cd0977c98624a99524eca8d4423654d173754ece08ecd71dbb1886a2655d478ba6a81c847cebd7031e76ea0d0b0b71621ae2855bf6c016937736fef647cf4626d3ab1dd0c4c2c7b1f389eeda79;
    5'b00101 : xpb = 1024'h4304f5d43ce798aa620e487140c3631d0fcbdb4a02d16a96345cb2981508524f5941f9c45ab7c5b415188b44ad1501e15c933c53b1cf9faee95c8ae77bb531cdacae9e4d4ef5c3975a19632fec0377d9fd95b35de8bf03cf9ea3566a090496602b080d02568ff88a4b0c4b2dcae2973ac7f4495ed9acbf11bea6022d05c0c447;
    5'b00110 : xpb = 1024'h97180f87637532b66079ba11210e9376a6bd6ed2bf2b267da461207260d7db2f3938f7825752531125dcc06ec43ed5c5ca54bec07cda46235eaec0084594040a97579fd5d82db66ad9f5ab47585c117f91e8d4adb5e7b03306fc3bb05549c24779a64a137b638dab5cc1e9c356965e570f7c4acc58870a8f00f3cd6b0a751480;
    5'b00111 : xpb = 1024'h3a7de3e4c81497f993dfb3d9f0ff7c7ecc38ff2aa60d41ed9688d4f6f9a4b70715e777c789c661df9742b651f80a98dfd3fc194725321c4c2361b5cad4a061960db16cafb1d4abf94737f0bc2bd8e6f43236fc64f68a2f85b9c88efbe7644b9c993cf4faef6e2a3ee7b7a179ea79ff4a082a6d578715f8dbfcd21da48646fe4e;
    5'b01000 : xpb = 1024'h8e90fd97eea23205924b2579d14aacd8632a92b36266fdd5068d42d145743fe6f5de75858660ef3ca806eb7c0f346cc441bd9bb3f03cc2c098b3eaeb9e7f33d2f85a6e383b0c9eccc71438d398318099c68a1db4c3b2dbe92221744233a97783e7db320c1441bf5ff96d400f762dc6664fb26ec505f044593f1fe8e28afb4e87;
    5'b01001 : xpb = 1024'h31f6d1f553419748c5b11f42a13b95e088a6230b49491944f8b4f755de411bbed28cf5cab8d4fe0b196ce15f43002fde4b64f63a989498e95d66e0ae2d8b915e6eb43b1214b3945b34567e486bae560e66d8456c04555b3bd4edc78dc5c400d90771dcf3884c5bf38462f7c60a11675948609150347f32a63afe391c06cd3855;
    5'b01010 : xpb = 1024'h8609eba879cf3154c41c90e28186c63a1f97b69405a2d52c68b965302a10a49eb283f388b56f8b682a3116895a2a03c2b92678a7639f3f5dd2b915cef76a639b595d3c9a9deb872eb432c65fd806efb3fb2b66bbd17e079f3d46acd412092cc056101a04ad1ff1149618965b95c52e758fe892bdb3597e237d4c045a0b81888e;
    5'b01011 : xpb = 1024'h296fc005de6e9697f7828aab5177af42451346ebec84f09c5ae119b4c2dd80768f3273cde7e39a369b970c6c8df5c6dcc2cdd32e0bf71586976c0b918676c126cfb7097477927cbd21750bd4ab83c5289b798e73122086f1f013001fa423b61575a6c4ec212a8da8210e4e1229a8cf688896b548e1e86c70792a54938753725c;
    5'b01100 : xpb = 1024'h7d82d9b904fc30a3f5edfc4b31c2df9bdc04da74a8deac83cae5878f0ead09566f29718be47e2793ac5b4196a51f9ac1308f559ad701bbfb0cbe40b250559363ba600afd00ca6f90a15153ec17dc5ece2fccafc2df493355586be565f068e1fcc44501fd45fe22c932c3eca7b55c9684d01eb6b660c2b7edbb781fd18c07c295;
    5'b01101 : xpb = 1024'h20e8ae16699b95e72953f61401b3c8a401806acc8fc0c7f3bd0d3c13a779e52e4bd7f1d116f236621dc13779d8eb5ddb3a36b0217f599223d1713674df61f0ef30b9d7d6da71651f0e939960eb593442d01ad77a1febb2a80b3838b182836b51e3dbace4ba08bf5cbdb9a45e49403777c8ccd9418f51a63ab756700b07d9ac63;
    5'b01110 : xpb = 1024'h74fbc7c990292ff327bf67b3e1fef8fd9871fe554c1a83db2d11a9edf3496e0e2bceef8f138cc3bf2e856ca3f01531bfa7f8328e4a64389846c36b95a940c32c1b62d95f63a957f28e6fe17857b1cde8646df8c9ed145f0b73911df7cec897393279e9f5dedc547dcf6f42f3d4f3fe941054daaf0e2bf1b7f9a43b490c8dfc9c;
    5'b01111 : xpb = 1024'h18619c26f4c895365b25617cb1efe205bded8ead32fc9f4b1f395e728c1649e6087d6fd44600d28d9feb628723e0f4d9b19f8d14f2bc0ec10b766158384d20b791bca6393d504d80fbb226ed2b2ea35d04bc20812db6de5e265d714360e3208e521094dd52e6f1115a64faaa68d79f870902fd3a3cbae004f5828b82885fe66a;
    5'b10000 : xpb = 1024'h6c74b5da1b562f425990d31c923b125f54df2235ef565b328f3dcc4cd7e5d2c5e8746d92429b5feab0af97b13b0ac8be1f610f81bdc6b53580c89679022bf2f47c65a7c1c68840547b8e6f0497873d02990f41d0fadf8ac18eb65689ad284c75a0aed1ee77ba86326c1a993ff48b66a3508afea7bb952b8237d056c08d1436a3;
    5'b10001 : xpb = 1024'hfda8a377ff594858cf6cce5622bfb677a5ab28dd63876a2816580d170b2ae9dc522edd7750f6eb922158d946ed68bd829086a08661e8b5e457b8c3b9138507ff2bf749ba02f35e2e8d0b4796b041277395d69883b820a144182a9d53f42d5cac0457cd5ebc522c5f71050f6886f079649392132ea2419cf33aea6fa08e62071;
    5'b10010 : xpb = 1024'h63eda3eaa6832e918b623e8542772bc1114c461692923289f169eeabbc82377da519eb9571a9fc1632d9c2be86005fbc96c9ec75312931d2bacdc15c5b1722bcdd687624296728b668acfc90d75cac1ccdb08ad808aab677a9db8f1b8b8801b20ee3b9e71098b7e708c5ef8c1422ceb290c122a068fe654c75fc72380d9a70aa;
    5'b10011 : xpb = 1024'h75378480b2293d4bec8384e126814c936c7d66e79744df9e391a330554f135581c86bdaa41e0ae4a43fb8a1b9cc22d6a07146fbd98107fb7f80b71eea23804853c242fe030e1e44d5ef4205aad981916dfeb28f494d35ca5ca7e2671da28b072e7a64ce84a3547a93bba742a8066fa5896f452b978d539971dac271896c5a78;
    5'b10100 : xpb = 1024'h5b6691fb31b02de0bd33a9edf2b34522cdb969f735ce09e15396110aa11e9c3561bf6998a0b89841b503edcbd0f5f6bb0e32c968a48bae6ff4d2ec3fb40252853e6b44868c46111855cb8a1d17321b370251d3df1675e22dc500c7ad69e7b6ee7d18a1dfa976e99ba57145d833ba36c1d0f7469916679f16b4288daf8e20aab1;
    5'b10101 : xpb = 1024'haf79abae583dc7ecbb9f1b8dd2fe757c64aafd7ff227c5c8c39a7ee4ecee251541b667569d53259ec5c822f5e81fca9f7bf44bd56f9654e46a2521607de124c22914460f157e03ebd5a7d234838ab4dc96a4f52ee39e8e912d59acf3b62ce2d5cbb6def0ce4a7ebcb726e46dbf6dfdde187f48069541ea93f67658ed92d4faea;
    5'b10110 : xpb = 1024'h52df800bbcdd2d2fef051556a2ef5e848a268dd7d909e138b5c2336985bb00ed1e64e79bcfc7346d372e18d91beb8db9859ba65c17ee2b0d2ed817230ced824d9f6e12e8ef24f97a42ea17a957078a5136f31ce624410de3e026003f48476c2aeb4d89d842551b50421c9c2453519ed1112d6a91c3d0d8e0f254a9270ea6e4b8;
    5'b10111 : xpb = 1024'ha6f299bee36ac73bed7086f6833a8ede2118216095639d2025c6a143d18a89ccfe5be559cc61c1ca47f24e033315619df35d28c8e2f8d181a42a4c43d6cc548a8a171471785cec4dc2c65fc0c36023f6cb463e35f169ba47487ee585948c981239ebc6e96728b07153d23ab9df0565ed58b56bff42ab245e34a27465135b34f1;
    5'b11000 : xpb = 1024'h4a586e1c480a2c7f20d680bf532b77e64693b1b87c45b89017ee55c86a5765a4db0a659efed5d098b95843e666e124b7fd04834f8b50a7aa68dd420665d8b2160070e14b5203e1dc3008a53596dcf96b6b9465ed320c3999fb4b38d126a72167598271d0db334d04dec7f27072e906e051638e8a713a12ab3080c49e8f2d1ebf;
    5'b11001 : xpb = 1024'h9e6b87cf6e97c68b1f41f25f3376a83fdd854541389f747787f2c3a2b626ee84bb01635cfb705df5ca1c79107e0af89c6ac605bc565b4e1ede2f77272fb78452eb19e2d3db3bd4afafe4ed4d03359310ffe7873cff34e5fd63a41e1772ec4d4ea820aee20006e225f07d9105fe9ccdfc98eb8ff7f0145e2872ce8fdc93e16ef8;
    5'b11010 : xpb = 1024'h41d15c2cd3372bce52a7ec28036791480300d5991f818fe77a1a78274ef3ca5c97afe3a22de46cc43b826ef3b1d6bbb6746d6042feb32447a2e26ce9bec3e1de6173afadb4e2ca3e1d2732c1d6b26885a035aef43fd76550167071630506d6a3c7b759c974117eb97b7348bc92806eef9199b2831ea34c756eace0160fb358c6;
    5'b11011 : xpb = 1024'h95e475dff9c4c5da51135dc7e3b2c1a199f26921dbdb4bceea1ee6019ac3533c77a6e1602a7efa214c46a41dc9008f9ae22ee2afc9bdcabc1834a20a88a2b41b4c1cb1363e1abd119d037ad9430b022b3488d0440d0011b37ec956a9514c028b165596da98e513da8d28e7521e34360bd921b3f09d7d97f2b0faab541467a8ff;
    5'b11100 : xpb = 1024'h394a4a3d5e642b1d84795790b3a3aaa9bf6df979c2bd673edc469a8633902f14545561a55cf308efbdac9a00fccc52b4ebd63d367215a0e4dce797cd17af11a6c2767e1017c1b2a00a45c04e1687d79fd4d6f7fb4da291063195a9f4e3668be035ec41c20cefb06e181e9f08b217d6fed1cfd67bcc0c863facd8fb8d903992cd;
    5'b11101 : xpb = 1024'h8d5d63f084f1c52982e4c93093eedb03565f8d027f1723264c4b08607f5fb7f4344c5f63598d964cce70cf2b13f626995997bfa33d2047595239ccede18de3e3ad1f7f98a0f9a5738a22086582e07145692a194b1acb3d6999ee8f3b2fabb7c7848a7ed331c3458f29d43d9e3dcb9e1b1957d7e94ae6d1bcef26c6cb94ede306;
    5'b11110 : xpb = 1024'h30c3384de9912a6cb64ac2f963dfc40b7bdb1d5a65f93e963e72bce5182c93cc10fadfa88c01a51b3fd6c50e47c1e9b3633f1a29e5781d8216ecc2b0709a416f23794c727aa09b01f7644dda565d46ba097841025b6dbcbc4cbae286c1c6411ca42129baa5cde222b4c9f554d1af3f0e1205fa747975c009eb05170510bfccd4;
    5'b11111 : xpb = 1024'h84d65201101ec478b4b63499442af46512ccb0e32252fa7dae772abf63fc1cabf0f1dd66889c3278509afa385eebbd97d1009c96b082c3f68c3ef7d13a7913ac0e224dfb03d88dd5774095f1c2b5e05f9dcb62522896691fb513c7cd0e0b6d03f2bf66cbcaa17743c67f93ea5d63062a598dfbe1f8500b872d52e24315741d0d;
    endcase
end

endmodule

module xpb_5_75
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h1689caec76c5c4178a1778f2ffb895fdac5536157bcbc4b651f64365d3a640dabecf25ecb59291531a89e021cc8a3588438f32f1b8dcc16619228cd4f1b9f86613dbfc6f08d842bc1ed929e636aacf45d8422d04308d1a2d55c04a52fe53631cdbd161e565ba9094413139035405a8dcb74a8778d60f23bc6d06fc379666f46b;
    5'b00010 : xpb = 1024'h2d1395d8ed8b882f142ef1e5ff712bfb58aa6c2af797896ca3ec86cba74c81b57d9e4bd96b2522a63513c04399146b10871e65e371b982cc324519a9e373f0cc27b7f8de11b085783db253cc6d559e8bb0845a08611a345aab8094a5fca6c639b7a2c3cacb75212882627206a80b51b96e950ef1ac1e4778da0df86f2ccde8d6;
    5'b00011 : xpb = 1024'h439d60c564514c469e466ad8ff29c1f904ffa24073634e22f5e2ca317af2c2903c6d71c620b7b3f94f9da065659ea098caad98d52a9644324b67a67ed52de9323b93f54d1a88c8345c8b7db2a4006dd188c6870c91a74e880140def8fafa2956937425b0312fb1bcc393ab09fc10fa9625df966a822d6b354714f4a6c334dd41;
    5'b00100 : xpb = 1024'h5a272bb1db17105e285de3cbfee257f6b154d855ef2f12d947d90d974e99036afb3c97b2d64a454c6a2780873228d6210e3ccbc6e3730598648a3353c6e7e1984f6ff1bc23610af07b64a798daab3d176108b410c23468b55701294bf94d8c736f45879596ea425104c4e40d5016a372dd2a1de3583c8ef1b41bf0de599bd1ac;
    5'b00101 : xpb = 1024'h70b0f69e51dcd475b2755cbefe9aedf45daa0e6b6afad78f99cf50fd223f4445ba0bbd9f8bdcd69f84b160a8feb30ba951cbfeb89c4fc6fe7dacc028b8a1d9fe634bee2b2c394dac9a3dd17f11560c5d394ae114f2c182e2acc1739ef7a0ef904b16e97afca4d2e545f61d10a41c4c4f9474a55c2e4bb2ae2122ed15f002c617;
    5'b00110 : xpb = 1024'h873ac18ac8a2988d3c8cd5b1fe5383f209ff4480e6c69c45ebc59462f5e5852078dae38c416f67f29f3b40cacb3d4131955b31aa552c886496cf4cfdaa5bd2647727ea9a35119068b916fb654800dba3118d0e19234e9d100281bdf1f5f452ad26e84b60625f637987275613f821f52c4bbf2cd5045ad66a8e29e94d8669ba82;
    5'b00111 : xpb = 1024'h9dc48c773f685ca4c6a44ea4fe0c19efb6547a96629260fc3dbbd7c8c98bc5fb37aa0978f701f945b9c520ec97c776b9d8ea649c0e0949caaff1d9d29c15caca8b03e7093de9d324d7f0254b7eabaae8e9cf3b1d53dbb73d58420844f447b5ca02b9ad45c819f40dc8588f174c279e090309b44dda69fa26fb30e5851cd0aeed;
    5'b01000 : xpb = 1024'h3a1120df43febf385b64fc0ed6a689bf133ad7b08e6853b11d561d8ea2f59cdf330b1ece26e0c0a34f0c1c780f39b77b85f6fa7a4333ae51875274952fd4e7f2a90aec99731189be42f4c8f1c7ab5fdce0c6e88f7e2a459f875c09d38707654af837d017d0b8c1482c9e13ba85d20bc6b7a5ce4602dc0b321c866b82a553ced;
    5'b01001 : xpb = 1024'h1a2adcfa6b05b00b0fcdc8b3ed22fe999d88e39084b249f163cba53ebdd59aa8b1ffd7d998009d5d4f7aa1e94d7dd0fffbeea2995d0ffc4b3197b41e44b746e53e6cab38a0095b580308767553258543a64e9b8d286fbe874e360af036c3d9718b54dee6e2c61ca8c3fb1a3efc62c99922c4e45d363ce46f8ecf62efc0bc3158;
    5'b01010 : xpb = 1024'h30b4a7e6e1cb742299e541a6ecdb949749de19a6007e0ea7b5c1e8a4917bdb8370cefdc64d932eb06a04820b1a0806883f7dd58b15ecbdb14aba40f336713f4b5248a7a7a8e19e1421e1a05b89d054897e90c89158fcd8b4a3f6554335173c8e672640cc4880ad3d052c534250687275da0f6bd60c4c082bfbd65f27572325c3;
    5'b01011 : xpb = 1024'h473e72d35891383a23fcba99ec942a94f6334fbb7c49d35e07b82c0a65221c5e2f9e23b30325c003848e622ce6923c10830d087ccec97f1763dccdc8282b37b16624a416b1b9e0d040baca41c07b23cf56d2f5958989f2e1f9b69f96336a9fab42f7a2b1ae3b3dd1465d8c45a46e1b529159f34ee25b2be868dd5b5eed8a1a2e;
    5'b01100 : xpb = 1024'h5dc83dbfcf56fc51ae14338cec4cc092a28885d0f815981459ae6f7038c85d38ee6d499fb8b851569f18424eb31c7198c69c3b6e87a6407d7cff5a9d19e530177a00a085ba92238c5f93f427f725f3152f152299ba170d0f4f76e9e931be02c81ec9049713f5ce65878ec548f873c42f48a47ac7b86a4fa4d5e4579683f10e99;
    5'b01101 : xpb = 1024'h745208ac461cc069382bac7fec0556904eddbbe673e15ccaaba4b2d60c6e9e13ad3c6f8c6e4ae2a9b9a222707fa6a7210a2b6e60408301e39621e7720b9f287d8ddc9cf4c36a66487e6d1e0e2dd0c25b07574f9deaa4273ca537343c301165e4fa9a667c79b05ef9c8bffe4c4c796d0bffef02408e79736142eb53ce1a580304;
    5'b01110 : xpb = 1024'h8adbd398bce28480c2432572ebbdec8dfb32f1fbefad2180fd9af63be014deee6c0b957923dd73fcd42c02924c30dca94dbaa151f95fc349af447446fd5920e3a1b89963cc42a9049d4647f4647b91a0df997ca21b314169faf77e8f2e64c901d66bc861df6aef8e09f1374fa07f15e8b73989b96488971daff25005b0bef76f;
    5'b01111 : xpb = 1024'ha1659e8533a848984c5a9e65eb76828ba78828116b78e6374f9139a1b3bb1fc92adabb65d970054feeb5e2b418bb12319149d443b23c84afc867011bef131949b59495d2d51aebc0bc1f71da9b2660e6b7dba9a64bbe5b9750b7c8e22cb82c1eb23d2a47452580224b227052f484bec56e8411323a97bada1cf94c3d4725ebda;
    5'b10000 : xpb = 1024'h742241be87fd7e70b6c9f81dad4d137e2675af611cd0a7623aac3b1d45eb39be66163d9c4dc181469e1838f01e736ef70bedf4f486675ca30ea4e92a5fa9cfe55215d932e623137c85e991e38f56bfb9c18dd11efc548b3f0eb813a70e0eca95f06fa02fa1718290593c27750ba4178d6f4b9c8c05b81664390cd7054aa79da;
    5'b10001 : xpb = 1024'h1dcbef085f459bfe95841874da8d67358ebc910b8d98cf2c75a10717a804f476a53089c67a6ea967846b63b0ce716c77b44e1241014337304a0cdb6797b4956468fd5a02373a73f3e737c3046fa03b41745b0a16205262e146abcb8d6f344fc63ad85be85fd1a8bd46c4fb7aa4bfea558e3f4141966aa522b097c9a7eb116e45;
    5'b10010 : xpb = 1024'h3455b9f4d60b60161f9b9167da45fd333b11c721096493e2c7974a7d7bab355163ffafb330013aba9ef543d29afba1fff7dd4532ba1ff896632f683c896e8dca7cd956714012b6b00610eceaa64b0a874c9d371a50df7d0e9c6c15e06d87b2e316a9bdcdc58c395187f6347df8c593324589c8ba6c79c8df1d9ec5df817862b0;
    5'b10011 : xpb = 1024'h4adf84e14cd1242da9b30a5ad9fe9330e766fd3685305899198d8de34f51762c22ced59fe593cc0db97f23f46785d7883b6c782472fcb9fc7c51f5117b28863090b552e048eaf96c24ea16d0dcf5d9cd24df641e816c973bf22c60336bdb15fff27b1fb32b46c9e5c9276d814ccb3c0efcd450334288ec9b8aa5c21717df571b;
    5'b10100 : xpb = 1024'h61694fcdc396e84533ca834dd9b7292e93bc334c00fc1d4f6b83d14922f7b706e19dfb8c9b265d60d409041634100d107efbab162bd97b62957481e66ce27e96a4914f4f51c33c2843c340b713a0a912fd219122b1f9b16947ecaa866a2e791cce4c819891015a7a0a58a684a0d0e4ebb41ed7ac18981057f7acbe4eae464b86;
    5'b10101 : xpb = 1024'h77f31aba3a5cac5cbde1fc40d96fbf2c401169617cc7e205bd7a14aef69df7e1a06d217950b8eeb3ee92e438009a4298c28ade07e4b63cc8ae970ebb5e9c76fcb86d4bbe5a9b7ee4629c6a9d4a4b7858d563be26e286cb969dacf4d96881dc39aa1de37df6bbeb0e4b89df87f4d68dc86b695f24eea7341464b3ba8644ad3ff1;
    5'b10110 : xpb = 1024'h8e7ce5a6b122707447f97533d9285529ec669f76f893a6bc0f705814ca4438bc5f3c4766064b8007091cc459cd247821061a10f99d92fe2ec7b99b9050566f62cc49482d6373c1a08175948380f6479eada5eb2b1313e5c3f36d3f2c66d53f5685ef45635c767ba28cbb188b48dc36a522b3e69dc4b657d0d1bab6bddb14345c;
    5'b10111 : xpb = 1024'ha506b09327e8348bd210ee26d8e0eb2798bbd58c745f6b7261669b7a9dea79971e0b6d52bbde115a23a6a47b99aeada949a943eb566fbf94e0dc2865421067c8e025449c6c4c045ca04ebe69b7a116e485e8182f43a0fff1492d897f6528a27361c0a748c2310c36cdec518e9ce1df81d9fe6e169ac57b8d3ec1b2f5717b28c7;
    5'b11000 : xpb = 1024'hae33629dcbfc3da9122ef42c83f39d3d39b08711ab38fb13580258abe8e0d69d99215c6a74a241e9ed2455682dad267291e4ef6ec99b0af495f75dbf8f7eb7d7fb20c5cc59349d3ac8de5ad557021f96a254b9ae7a7ed0de96141d7a95162fe0e8a77047722a43d885da3b2f9176235426f16ad20894219655934287effb6c7;
    5'b11001 : xpb = 1024'h216d0116538587f21b3a6835c7f7cfd17ff03e86967f5467877668f092344e4498613bb35cdcb571b95c25784f6507ef6cad81e8a5767215628202b0eab1e3e3938e08cbce6b8c8fcb670f938c1af13f4267789f1835073b3f218c2aa7a4c61aea5bd8e9dcdd34d1c98edcb64d1d0b11f9b99e25f69865d5d26030601566ab32;
    5'b11010 : xpb = 1024'h37f6cc02ca4b4c09a551e128c7b065cf2c45749c124b191dd96cac5665da8f1f573061a0126f46c4d3e6059a1bef3d77b03cb4da5e53337b7ba48f85dc6bdc49a76a053ad743cf4bea403979c2c5c0851aa9a5a348c2216894e1d67da5f82937c62d3acf4297c5660ac015b9a122b3eeb104259ecca789923f672c97abcd9f9d;
    5'b11011 : xpb = 1024'h4e8096ef411110212f695a1bc768fbccd89aaab18e16ddd42b62efbc3980cffa15ff878cc801d817ee6fe5bbe87972fff3cbe7cc172ff4e194c71c5ace25d4afbb4601a9e01c12080919635ff9708fcaf2ebd2a7794f3b95eaa220d0a44b8c54a1fe9cb4a85255fa4bf14ebcf5285ccb684ead17a2b6ad4eac6e28cf42349408;
    5'b11100 : xpb = 1024'h650a61dbb7d6d438b980d30ec72191ca84efe0c709e2a28a7d5933220d2710d4d4cead797d94696b08f9c5ddb503a888375b1abdd00cb647ade9a92fbfdfcd15cf21fe18e8f454c427f28d46301b5f10cb2dffaba9dc55c340626b23a29eef717dcffe9a0e0ce68e8d2287c0492e05a81f99349078c5d10b19752506d89b8873;
    5'b11101 : xpb = 1024'h7b942cc82e9c985043984c01c6da27c8314516dc85ae6740cf4f7687e0cd51af939dd3663326fabe2383a5ff818dde107aea4daf88e977adc70c3604b199c57be2fdfa87f1cc978046cbb72c66c62e56a3702cafda696ff09622b576a0f2528e59a1607f73c77722ce53c0c39d33ae84d6e3bc094ed4f4c7867c213e6f027cde;
    5'b11110 : xpb = 1024'h921df7b4a5625c67cdafc4f4c692bdc5dd9a4cf2017a2bf72145b9edb473928a526cf952e8b98c113e0d86214e181398be7980a141c63913e02ec2d9a353bde1f6d9f6f6faa4da3c65a4e1129d70fd9c7bb259b40af68a1debe2ffc99f45b5ab3572c264d98207b70f84f9c6f13957618e2e438224e41883f3831d7605697149;
    5'b11111 : xpb = 1024'ha8a7c2a11c28207f57c73de7c64b53c389ef83077d45f0ad733bfd538819d365113c1f3f9e4c1d64589766431aa249210208b392faa2fa79f9514fae950db6480ab5f366037d1cf8847e0af8d41bcce253f486b83b83a44b41a34a1c9d9918c81144244a3f3c984b50b632ca453f003e4578cafafaf33c40608a19ad9bd065b4;
    endcase
end

endmodule

module xpb_5_275
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h6c00899b5a852da8200eda1677a8eb5368444be39d65b88991fa86a140db8a59512ecda5871a4505627d381d587090065f0d94d6d8f0f3180d12ea2d048067f59336c5e44dad8b8d1b15e8619788fab407b120fdab02b1774b799442225e81bac8c16bb8d4b9d085675c9819b5c1db2b3d525912090d6110bbafb89cc07ed8ec;
    5'b00010 : xpb = 1024'h2753cde0f31c268775183c55def78f555f1294966553d09ba61853ecceb467aa9f151dd2440e0b7c259c30f3cd830f425a0101c78f2f15e4698694fbce2e5b39b21e5719ebca19d52391ce20963631371b5d4862c97f35dde16696898a9260e3627b4547f8aaa87d47f9495473b3902d2bcad341c1cf64f130eff634f81b4b6d;
    5'b00011 : xpb = 1024'h9354577c4da1542f9527166c56a07aa8c756e07a02b989253812da8e0f8ff203f043eb77cb2850818819691125f39f48b90e969e682008fc76997f28d2aec32f45551cfe3977a5623ea7b6822dbf2beb230e69607481e7552ce02acbacf0e29e2b3cb100cd647902af55e16e29756b58691d2c53cadcc601ec9faed1b89a2459;
    5'b00100 : xpb = 1024'h4ea79bc1e6384d0eea3078abbdef1eaabe25292ccaa7a1374c30a7d99d68cf553e2a3ba4881c16f84b3861e79b061e84b402038f1e5e2bc8d30d29f79c5cb673643cae33d79433aa47239c412c6c626e36ba90c592fe6bbbc2cd2d131524c1c6c4f68a8ff15550fa8ff292a8e767205a5795a683839ec9e261dfec69f03696da;
    5'b00101 : xpb = 1024'h9fae0077ecf45ee3f39daeb253dc2acb4f371df9295b949604e75252b41aca68c108bd1450fdd6f0e575abe10189dc0aef5707fd49c4e952f80d4c6660aa9b783243f6975b0c1f24f9f82002b1998f14a66b82ab17af02258ba2f5a7d58a0ef5eb0641f154628f2708f43e3a558d55c460e20b33c60cdc2d7202a0227d3095b;
    5'b00110 : xpb = 1024'h75fb69a2d95473965f48b5019ce6ae001d37bdc32ffb71d2f248fbc66c1d36ffdd3f5976cc2a227470d492db68892dc70e030556ad8d41ad3c93bef36a8b11ad165b054dc35e4d7f6ab56a61c2a293a55217d9285c7da199a433c39c9fb722aa2771cfd7e9fff977d7ebdbfd5b1ab087836079c5456e2ed392cfe29ee851e247;
    5'b00111 : xpb = 1024'h314eade871eb6c75b45217410435520214060675f7e989e50666c911f9f614512b25a9a3891de8eb33f38bb1dd9bad0308f6724763cb6479990769c2343904f135429683617adbc773315020c14fca2865c4008d7afa26003a20c5e407eb01d2c12ba9670df0d16fb8888d38190c658971d8f3f4fe3032b4081020371fee54c8;
    5'b01000 : xpb = 1024'h9d4f3783cc709a1dd460f1577bde3d557c4a5259954f426e98614fb33ad19eaa7c54774910382df09670c3cf360c3d096804071e3cbc5791a61a53ef38b96ce6c8795c67af2867548e47388258d8c4dc6d75218b25fcd777859a5a262a49838d89ed151fe2aaa1f51fe52551cece40b4af2b4d07073d93c4c3bfd8d3e06d2db4;
    5'b01001 : xpb = 1024'h58a27bc9650792fd296a5396e32ce15773189b0c5d3d5a80ac7f1cfec8aa7bfbca3ac775cd2bf467598fbca5ab1ebc4562f7740ef2fa7a5e028dfebe0267602ae760ed9d4d44f59c96c31e415785fb5f812148f044795bde1b875c6d927d62b623a6eeaf069b79ed0081d68c8cbff5b69da3c736bfff97a53900166c1809a035;
    5'b01010 : xpb = 1024'h13f5c00efd9e8bdc7e73b5d64a7b855969e6e3bf252b7292c09cea4a5683594d182117a28a1fbade1caeb57c20313b815deae0ffa9389d2a5f01a98ccc15536f06487ed2eb6183e49f3f0400563331e294cd705562f5e044b1745eb4fab141debd60c83e2a8c51e4e11e87c74ab1aab88c1c416678c19b85ae4054044fa612b6;
    5'b01011 : xpb = 1024'h7ff649aa5823b9849e828fecc22470acd22b2fa2c2912b1c529770eb975ee3a6694fe5481139ffe37f2bed9978a1cb87bcf875d6822990426c1493b9d095bb64997f44b7390f0f71ba54ec61edbc2c969c7e91530df891bbfcedf2f71d0fc399862233f6ff46226a487b1fe1007385e3c96e9a7881cefc9669f00ca11024eba2;
    5'b01100 : xpb = 1024'h3b498deff0bab263f38bf22c297314aec8f978558a7f432e66b53e372537c0f7b7363574ce2dc65a424ae66fedb44ac3b7ebe2c73867b30ec8883e889a43aea8b866d5ecd72b9db9c2d0d220ec696319b02ab8b82c75162292daf53e8543a2c21fdc0d862336fa622917d11bbe653ae5b7e714a83a910076df304a3947c15e23;
    5'b01101 : xpb = 1024'ha74a178b4b3fe00c139acc42a11c0002313dc43927e4fbb7f8afc4d866134b510865031a55480b5fa4c81e8d4624daca16f9779e1158a626d59b28b59ec4169e4b9d9bd124d92946dde6ba8283f25dcdb7dbd9b5d777c799de548980a7a2247ce89d793ef7f0cae79074693574271610f5396dba439e61879ae002d60840370f;
    5'b01110 : xpb = 1024'h629d5bd0e3d6d8eb68a42e82086aa404280c0cebefd313ca0ccd9223f3ec28a2564b5347123bd1d667e71763bb375a0611ece48ec796c8f3320ed384687209e26a852d06c2f5b78ee662a041829f9450cb88011af5f44c0074418bc80fd603a5825752ce1be1a2df71111a703218cb12e3b1e7e9fc6065681020406e3fdca990;
    5'b01111 : xpb = 1024'h1df0a0167c6dd1cabdad90c16fb948061eda559eb7c12bdc20eb5f6f81c505f3a431a373cf2f984d2b06103a3049d9420ce0517f7dd4ebbf8e827e53321ffd26896cbe3c611245d6eede8600814ccad3df3428801470d0670a2e8e0f7809e2ce1c112c5d3fd27ad751adcbaaf00a8014d22a6219b522694885607e0677791c11;
    5'b10000 : xpb = 1024'h89f129b1d6f2ff72ddbc6ad7e7623359871ea1825526e465b2e5e610c2a0904cf56071195649dd528d83485788ba69486bede65656c5ded79b95688036a0651c1ca38420aebfd16409f46e6218d5c587e6e5497dbf7381de55a822519a686488e4d29816148c4b5cb90a63c4a5cc5b400f7cbb2bbe2fca59411036a337f7f4fd;
    5'b10001 : xpb = 1024'h45446df76f89f85232c5cd174eb0d75b7decea351d14fc77c703b35c50796d9e4346c146133da3c950a2412dfdcce88466e153470d0401a3f809134f004e58603b8b15564cdc5fac127054211782fc0afa9170e2ddf00644eb952499029c43b17e8c71a5387d235499a714ff63be1041fdf5355b76f1ce39b650743b6f94677e;
    5'b10010 : xpb = 1024'h97b23d0820f13187cf2f56b5ff7b5d74bb32e7e5031489db2180a7de524aef912d1172d0316a4013c13a0472df67c061d4c037c3422470547cbe1dc9fc4ba45a72a68beaf8edf41aec39e01630328e0e3d9847fc6c8aab818226e06ad022da18464b345c6dfb4c7a43c63a21afc543ec6daf8b2fb3d21a2b90b1d3a730d9ff;
    5'b10011 : xpb = 1024'h6c983bd862a61ed9a7de096d2da866b0dcff7ecb8268cd136d1c07491f2dd548e25bdf18574baf45763e7221cb4ff7c6c0e2550e9c331788618fa84ace7cb399eda96c7038a6798136022241adb92d4215eeb945a76f3c22ccfbbb228d2ea494e107b6ed3127cbd1e1a05e53d771a06f29c0089d38c1332ae7406a7067afb2eb;
    5'b10100 : xpb = 1024'h27eb801dfb3d17b8fce76bac94f70ab2d3cdc77e4a56e5258139d494ad06b29a30422f45143f75bc395d6af840627702bbd5c1ff52713a54be035319982aa6de0c90fda5d6c307c93e7e0800ac6663c5299ae0aac5ebc08962e8bd69f56283bd7ac1907c5518a3c9c23d0f8e95635571183882ccf183370b5c80a8089f4c256c;
    5'b10101 : xpb = 1024'h93ec09b955c245611cf645c30c9ff6063c121361e7bc9daf13345b35ede23cf38170fcea9b59bac19bdaa31598d307091ae356d62b622d6ccb163d469cab0ed39fc7c38a247093565993f06243ef5e79314c01a870ee7200ae6251ac17c105784382fc3529d2744f2999a7a84b25309c558adbdefa90981c183060a55fcafe58;
    5'b10110 : xpb = 1024'h4f3f4dfeee593e4071ffa80273ee9a0832e05c14afaab5c1275228817bbb1a44cf574d17584d81385ef99bec0de5864515d6c3c6e1a050392789e81566590217beaf54bfc28d219e620fd621429c94fc44f8290d8f6af667444f53f37ff4e4a0dd3cd5c44dc34c470a3658e30916e59e4403560eb3529bfc8d709e3d976770d9;
    5'b10111 : xpb = 1024'ha92924486f0371fc7090a41db3d3e0a29aea4c77798cdd33b6ff5cd0993f7961d3d9d44154147af221894c282f8058110ca30b797de730583fd92e43006f55bdd96e5f560a9afe66a8bbbe04149cb7f58a45072ade77acdda3c563ae828c3c976f6af5371b4243eead30a1dc7089aa0327bd03e6c149fdd02b0dbd5cf03e35a;
    5'b11000 : xpb = 1024'h76931bdfe17564c7e717e45852e6295d91f2f0ab14fe865ccd6a7c6e4a6f81ef6e6c6ae99c5b8cb48495ccdfdb6895876fd7c58e70cf661d91107d1134875d5170cdabd9ae573b7385a1a441d8d2c6336055717058ea2c4525b5ea7d0a8745843fb81b0c466df4c4522fa2377cca75cb6fce2950752200edbe6094728f82bc46;
    5'b11001 : xpb = 1024'h31e660257a0c5da73c214697ba34cd5f88c1395ddcec9e6ee18849b9d8485f40bc52bb16594f532b47b4c5b6507b14c36acb327f270d88e9ed8427dffe3550958fb53d0f4c73c9bb8e1d8a00d77ffcb6740198d57766b0abbba2ecc472bb24acd971f49b6a5eccbc32cc53723abc2acd5e46a3802de404ce33a0d20ac71f2ec7;
    5'b11010 : xpb = 1024'h9de6e9c0d4918b4f5c3020ae31ddb8b2f10585417a5256f87382d05b1923e99a0d8188bbe0699830aa31fdd3a8eba4c9c9d8c755fffe7c01fa97120d02b5b88b22ec02f39a215548a93372626f08f76a7bb2b9d322696223071c81069519a667a23360543f189d419a28eb8bf07e05f89b98fc9236f165deef508aa7879e07b3;
    5'b11011 : xpb = 1024'h593a2e066d28842eb13982ed992c5cb4e7d3cdf442406f0a87a09da6a6fcc6eb5b67d8e89d5d5ea76d50f6aa1dfe2405c4cc3446b63c9ece570abcdbcc63abcf41d39429383de390b1af58216db62ded8f5ee13840e5e6899d09834dfd4d85903bed39e3630975397ac59cc6ae6fbafa8a1176c1efb369bf6490c83fbf3a7a34;
    5'b11100 : xpb = 1024'h148d724c05bf7d0e0642e52d007b00b6dea216a70a2e871c9bbe6af234d5a43ca94e29155a51251e306fef809310a341bfbfa1376c7ac19ab37e67aa96119f1360bb255ed65a71d8ba2b3de06c636470a30b089d5f626af032f68595658164b8d5a7137286fa4d315b624e016c616ffc7889f0f1a8756d9fd9d105d7f6d6ecb5;
    5'b11101 : xpb = 1024'h808dfbe76044aab62651bf437823ec0a46e6628aa7943fa62db8f19375b12e95fa7cf6bae16b6a2392ed279deb8133481ecd360e456bb4b2c09151d79a920708f3f1eb432407fd65d541264203ec5f24aabc299b0a651c677e7019d787dfe6739e687f2b5bb41db6c2bee61b22234b27b5dc4a03b182ceb09580be74b755c5a1;
    5'b11110 : xpb = 1024'h3be1402cf8dba3957b5b2182df72900c3db4ab3d6f8257b841d6bedf038a0be7486346e79e5f309a560c20746093b28419c0a2fefba9d77f1d04fca6643ffa4d12d97c78c2248badddbd0c01029995a7be68510028e1a0ce145d1c1ef013c59c382258ba7fa4f5aea35b9755e0150029a454c4336a44d2910ac0fc0ceef23822;
    5'b11111 : xpb = 1024'ha7e1c9c85360d13d9b69fb99571b7b5fa5f8f7210ce81041d3d14580446596409992148d2579759fb8895891b904428a78ce37d5d49aca972a17e6d368c06242a610425d0fd2173af8d2f4629a22905bc61971fdd3e452455fd6b0611272475700e3c473545ec6340ab82f6f95d6db54e1a71d45735233a1c670b4a9af71110e;
    endcase
end

endmodule

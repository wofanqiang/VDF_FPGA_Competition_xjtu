module xpb_5_995
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h1fa4044cf463e42fbb91056d24f0ad9b2656b4eee0cfc626857fb123da69c1fb4beeaee1b0db47a51aa516722b09ade2fb5e0dc24e3b7a92e082ae365e55624f3bc1e5d87f42cebd579e4b18993ab77ed1d34157ae1deae48ce078d7cfa20965b6c64fa82d5c0202a54949993831e1ed092f304770df058b2aa1585b187de81;
    5'b00010 : xpb = 1024'h3f480899e8c7c85f77220ada49e15b364cad69ddc19f8c4d0aff6247b4d383f697dd5dc361b68f4a354a2ce456135bc5f6bc1b849c76f525c1055c6cbcaac49e7783cbb0fe859d7aaf3c963132756efda3a682af5c3bd5c919c0f1af9f4412cb6d8c9f505ab804054a9293327063c3da125e608ee1be0b165542b0b630fbd02;
    5'b00011 : xpb = 1024'h5eec0ce6dd2bac8f32b310476ed208d173041ecca26f5273907f136b8f3d45f1e3cc0ca51291d6ef4fef4356811d09a8f21a2946eab26fb8a1880aa31b0026edb345b1897dc86c3806dae149cbb0267c7579c4070a59c0ada6a16a876ee61c312452eef888140607efdbdccba895a5c71b8d90d6529d10a17fe409114979b83;
    5'b00100 : xpb = 1024'h7e901133d18f90beee4415b493c2b66c995ad3bb833f189a15fec48f69a707ed2fbabb86c36d1e946a9459c8ac26b78bed78370938edea4b820ab8d97955893cef079761fd0b3af55e792c6264eaddfb474d055eb877ab923381e35f3e882596db193ea0b570080a95252664e0c787b424bcc11dc37c162caa85616c61f7a04;
    5'b00101 : xpb = 1024'h9e341580c5f374eea9d51b21b8b36407bfb188aa640edec09b7e75b34410c9e87ba96a68744866398539703ad730656ee8d644cb872964de628d670fd7aaeb8c2ac97d3a7c4e09b2b617777afe25957a192046b666959676c0625c370e2a2efc91df8e48e2cc0a0d3a6e6ffe18f969a12debf165345b1bb7d526b9c77a75885;
    5'b00110 : xpb = 1024'hbdd819cdba57591e6566208edda411a2e6083d9944dea4e720fe26d71e7a8be3c798194a2523adde9fde86ad023a1351e434528dd564df714310154636004ddb668b6312fb90d8700db5c29397604cf8eaf3880e14b3815b4d42d50eddcc386248a5ddf110280c0fdfb7b997512b4b8e371b21aca53a2142ffc8122292f3706;
    5'b00111 : xpb = 1024'hdd7c1e1aaebb3d4e20f725fc0294bf3e0c5ef28825ae6b0da67dd7faf8e44ddf1386c82bd5fef583ba839d1f2d43c134df92605023a05a042392c37c9455b02aa24d48eb7ad3a72d65540dac309b0477bcc6c965c2d16c3fda234de6ad6e41c7ff6c2d993d840e1285010330895d2d7b404a51f4161926ce2a696a7dab71587;
    5'b01000 : xpb = 1024'hfd202267a31f217ddc882b6927856cd932b5a777067e31342bfd891ed34e0fda5f75770d86da3d28d528b391584d6f17daf06e1271dbd497041571b2f2ab1279de0f2ec3fa1675eabcf258c4c9d5bbf68e9a0abd70ef57246703c6be7d104b2db6327d416ae010152a4a4cc9c18f0f684979823b86f82c59550ac2d8c3ef408;
    5'b01001 : xpb = 1024'h11cc426b4978305ad981930d64c761a74590c5c65e74df75ab17d3a42adb7d1d5ab6425ef37b584cdefcdca0383571cfad64e7bd4c0174f29e4981fe9510074c919d1149c795944a81490a3dd63107375606d4c151f0d4208f3e43f964cb254936cf8cce9983c1217cf939662f9c0f15552a8b282f7d731e47fac1b33dc6d289;
    5'b01010 : xpb = 1024'h13c682b018be6e9dd53aa36437166c80f7f631154c81dbd8136fceb66882193d0f752d4d0e890cc730a72e075ae60caddd1ac89970e52c9bcc51ace1faf55d7185592fa74f89c13656c2eeef5fc4b2af432408d6ccd2b2ced80c4b86e1c545df923bf1c91c598141a74dcdffc31f2d3425bd7e2ca68b6376faa4d738ef4eb10a;
    5'b01011 : xpb = 1024'h15c0c2f4e804ace0d0f3b3bb0965775aaa5b9c643a8ed83a7bc7c9c8a628b55cc434183b2996c14182517f6e7d96a78c0cd0a97595c8e444fa59d7c560dab39679154e04d77dee222c3cd3a0e9585e2730413cec47b4917d20da53145ebf6675eda856c39f2f4161d1a2629956a24b52f65071311d9953cfad4eecbea0d68f8b;
    5'b01100 : xpb = 1024'h17bb0339b74aeb23ccacc411dbb482345cc107b3289bd49ce41fc4dae3cf517c78f3032944a475bbd3fbd0d5a047426a3c868a51baac9bee286202a8c6c009bb6cd16c625f721b0e01b6b85272ec099f1d5e7101c296702b69a85aa1dbb9870c4914bbbe22050181fbf6f732ea256971c6e3643594a744285ff90244525e6e0c;
    5'b01101 : xpb = 1024'h19b5437e86912966c865d468ae038d0e0f26730216a8d0ff4c77bfed2175ed9c2db1ee175fb22a3625a6223cc2f7dd486c3c6b2ddf905397566a2d8c2ca55fe0608d8abfe76647f9d7309d03fc7fb5170a7ba5173d784ed9b276622f58b3a7a2a48120b8a4dac1a2264b8bcc7da887909776573a0bb5348112a317ca03e64c8d;
    5'b01110 : xpb = 1024'h1baf83c355d767a9c41ee4bf805297e7c18bde5104b5cd61b4cfbaff5f1c89bbe270d9057abfdeb0775073a3e5a878269bf24c0a04740b408472586f928ab6055449a91d6f5a74e5acaa81b58613608ef798d92cb85a2d87fb4469bcd5adc838ffed85b327b081c250a02066112ba5af68094a3e82c324d9c54d2d4fb56e2b0e;
    5'b01111 : xpb = 1024'h1da9c408251da5ecbfd7f51652a1a2c173f1499ff2c2c9c41d27b6119cc325db972fc3f395cd932ac8fac50b08591304cba82ce62957c2e9b27a8352f8700c2a4805c77af74ea1d1822466670fa70c06e4b60d42333c0c364412714a52a7e8cf5b59eaadaa8641e27af4b4ffa4aec3ce389c3d42f9d1153277f742d566f6098f;
    5'b10000 : xpb = 1024'h1fa4044cf463e42fbb91056d24f0ad9b2656b4eee0cfc626857fb123da69c1fb4beeaee1b0db47a51aa516722b09ade2fb5e0dc24e3b7a92e082ae365e55624f3bc1e5d87f42cebd579e4b18993ab77ed1d34157ae1deae48ce078d7cfa20965b6c64fa82d5c0202a54949993831e1ed092f304770df058b2aa1585b187de810;
    5'b10001 : xpb = 1024'h219e4491c3aa2272b74a15c3f73fb874d8bc203dcedcc288edd7ac3618105e1b00ad99cfcbe8fc1f6c4f67d94dba48c12b13ee9e731f323c0e8ad919c43ab8742f7e04360736fba92d182fca22ce62f6bef0756d28ffc992d5ae80654c9c29fc1232b4a2b031c222cf9dde32cbb5000bd9c2234be7ecf5e3dd4b6de0ca05c691;
    5'b10010 : xpb = 1024'h239884d692f060b5b303261ac98ec34e8b218b8cbce9beeb562fa74855b6fa3ab56c84bde6f6b099bdf9b940706ae39f5ac9cf7a9802e9e53c9303fd2a200e99233a22938f2b28950292147bac620e6eac0da982a3e1a8411e7c87f2c9964a926d9f199d33078242f9f272cc5f381e2aaa5516505efae63c8ff583667b8da512;
    5'b10011 : xpb = 1024'h2592c51b62369ef8aebc36719bddce283d86f6dbaaf6bb4dbe87a25a935d965a6a2b6fac020465140fa40aa7931b7e7d8a7fb056bce6a18e6a9b2ee0900564be16f640f1171f5580d80bf92d35f5b9e6992add981ec386ef674a8f8046906b28c90b7e97b5dd426324470765f2bb3c497ae80954d608d695429f98ec2d158393;
    5'b10100 : xpb = 1024'h278d0560317cdd3baa7546c86e2cd901efec622a9903b7b026df9d6cd104327a1eea5a9a1d12198e614e5c0eb5cc195bba359132e1ca593798a359c3f5eabae30ab25f4e9f13826cad85dddebf89655e864811ad99a5659db018970dc38a8bbf2477e39238b302834e9b9bff863e5a684b7afc594d16c6edf549ae71de9d6214;
    5'b10101 : xpb = 1024'h298745a500c31b7ea62e571f407be3dba251cd798710b4128f37987f0eaace99d3a94588381fce08b2f8ad75d87cb439e9eb720f06ae10e0c6ab84a75bd01107fe6e7dac2707af5882ffc290491d10d6736545c31487444bf8e69e9b4084ac557fe4488cbb88c2a378f0309919c178871c0def5dc424b746a7f3c3f790254095;
    5'b10110 : xpb = 1024'h2b8185e9d00959c1a1e7677612caeeb554b738c8751db074f78f93914c516ab988683076532d828304a2fedcfb2d4f1819a152eb2b91c889f4b3af8ac1b5672cf22a9c09aefbdc445879a741d2b0bc4e608279d88f6922fa41b4a628bd7eccebdb50ad873e5e82c3a344c532ad4496a5eca0e2623b32a79f5a9dd97d41ad1f16;
    5'b10111 : xpb = 1024'h2d7bc62e9f4f98049da077cce519f98f071ca417632aacd75fe78ea389f806d93d271b646e3b36fd564d50441ddde9f6495733c75075803322bbda6e279abd51e5e6ba6736f009302df38bf35c4467c64d9fadee0a4b01a88a82adb63a78ed8236bd1281c13442e3cd9959cc40c7b4c4bd33d566b24097f80d47ef02f334fd97;
    5'b11000 : xpb = 1024'h2f7606736e95d64799598823b7690468b9820f665137a939c83f89b5c79ea2f8f1e606528948eb77a7f7a1ab408e84d4790d14a3755937dc50c405518d801376d9a2d8c4bee4361c036d70a4e5d8133e3abce203852ce056d350b543b7730e189229777c440a0303f7edee65d44ad2e38dc6c86b294e8850bff20488a4bcdc18;
    5'b11001 : xpb = 1024'h317046b83ddc148a9512987a89b80f426be77ab53f44a59c309784c805453f18a6a4f140a4569ff1f9a1f312633f1fb2a8c2f57f9a3cef857ecc3034f365699bcd5ef72246d86307d8e755566f6bbeb627da1619000ebf051c1ebcd1346d2eaeed95dc76c6dfc324224282ff67cdf1025e59bb6fa05c78a9729c1a0e5644ba99;
    5'b11010 : xpb = 1024'h336a86fd0d2252cd90cba8d15c071a1c1e4ce6042d51a1fe98ef7fda42ebdb385b63dc2ebf64546c4b4c447985efba90d878d65bbf20a72eacd45b18594abfc0c11b157fcecc8ff3ae613a07f8ff6a2e14f74a2e7af09db364ecc45eb1674f454902417149b583444c971798fb510f212eecae74176a690225462f9407cc991a;
    5'b11011 : xpb = 1024'h3564c741dc6891108c84b9282e5624f5d0b251531b5e9e6101477aec809277581022c71cda7208e69cf695e0a8a0556f082eb737e4045ed7dadc85fbbf3015e5b4d733dd56c0bcdf83db1eb9829315a602147e43f5d27c61adbacbec2e616fdba46ea66bcc8b436476ebac328ed42d3fff7fa1788e78595ad7f04519b954779b;
    5'b11100 : xpb = 1024'h375f0786abaecf53883dc97f00a52fcf8317bca2096b9ac3699f75febe391377c4e1b20af57fbd60eea0e747cb50f04d37e4981408e8168108e4b0df25156c0aa893523adeb4e9cb5955036b0c26c11def31b25970b45b0ff688d379ab5b9071ffdb0b664f610384a14040cc22574b5ed012947d058649b38a9a5a9f6adc561c;
    5'b11101 : xpb = 1024'h395947cb7af50d9683f6d9d5d2f43aa9357d27f0f7789725d1f77110fbdfaf9779a09cf9108d71db404b38aeee018b2b679a78f02dcbce2a36ecdbc28afac22f9c4f709866a916b72ecee81c95ba6c95dc4ee66eeb9639be3f56db072855b1085b477060d236c3a4cb94d565b5da697da0a587817c943a0c3d4470251c64349d;
    5'b11110 : xpb = 1024'h3b5388104a3b4bd97fafea2ca5434582e7e2933fe58593883a4f6c2339864bb72e5f87e72b9b265591f58a1610b22609975059cc52af85d364f506a5f0e01854900b8ef5ee9d43a30448ccce1f4e180dc96c1a846678186c8824e294a54fd19eb6b3d55b550c83c4f5e969ff495d879c71387a85f3a22a64efee85aacdec131e;
    5'b11111 : xpb = 1024'h3d4dc85519818a1c7b68fa837792505c9a47fe8ed3928feaa2a76735772ce7d6e31e72d546a8dacfe39fdb7d3362c0e7c7063aa877933d7c92fd318956c56e7983c7ad537691708ed9c2b17fa8e1c385b6894e99e159f71ad0f2ea222249f23512203a55d7e243e5203dfe98dce0a5bb41cb6d8a6ab01abda2989b307f73f19f;
    endcase
end

endmodule

module compressor_array_72_24_1283
(
    input  [71:0] col_in_0,
    input  [71:0] col_in_1,
    input  [71:0] col_in_2,
    input  [71:0] col_in_3,
    input  [71:0] col_in_4,
    input  [71:0] col_in_5,
    input  [71:0] col_in_6,
    input  [71:0] col_in_7,
    input  [71:0] col_in_8,
    input  [71:0] col_in_9,
    input  [71:0] col_in_10,
    input  [71:0] col_in_11,
    input  [71:0] col_in_12,
    input  [71:0] col_in_13,
    input  [71:0] col_in_14,
    input  [71:0] col_in_15,
    input  [71:0] col_in_16,
    input  [71:0] col_in_17,
    input  [71:0] col_in_18,
    input  [71:0] col_in_19,
    input  [71:0] col_in_20,
    input  [71:0] col_in_21,
    input  [71:0] col_in_22,
    input  [71:0] col_in_23,
    input  [71:0] col_in_24,
    input  [71:0] col_in_25,
    input  [71:0] col_in_26,
    input  [71:0] col_in_27,
    input  [71:0] col_in_28,
    input  [71:0] col_in_29,
    input  [71:0] col_in_30,
    input  [71:0] col_in_31,
    input  [71:0] col_in_32,
    input  [71:0] col_in_33,
    input  [71:0] col_in_34,
    input  [71:0] col_in_35,
    input  [71:0] col_in_36,
    input  [71:0] col_in_37,
    input  [71:0] col_in_38,
    input  [71:0] col_in_39,
    input  [71:0] col_in_40,
    input  [71:0] col_in_41,
    input  [71:0] col_in_42,
    input  [71:0] col_in_43,
    input  [71:0] col_in_44,
    input  [71:0] col_in_45,
    input  [71:0] col_in_46,
    input  [71:0] col_in_47,
    input  [71:0] col_in_48,
    input  [71:0] col_in_49,
    input  [71:0] col_in_50,
    input  [71:0] col_in_51,
    input  [71:0] col_in_52,
    input  [71:0] col_in_53,
    input  [71:0] col_in_54,
    input  [71:0] col_in_55,
    input  [71:0] col_in_56,
    input  [71:0] col_in_57,
    input  [71:0] col_in_58,
    input  [71:0] col_in_59,
    input  [71:0] col_in_60,
    input  [71:0] col_in_61,
    input  [71:0] col_in_62,
    input  [71:0] col_in_63,
    input  [71:0] col_in_64,
    input  [71:0] col_in_65,
    input  [71:0] col_in_66,
    input  [71:0] col_in_67,
    input  [71:0] col_in_68,
    input  [71:0] col_in_69,
    input  [71:0] col_in_70,
    input  [71:0] col_in_71,
    input  [71:0] col_in_72,
    input  [71:0] col_in_73,
    input  [71:0] col_in_74,
    input  [71:0] col_in_75,
    input  [71:0] col_in_76,
    input  [71:0] col_in_77,
    input  [71:0] col_in_78,
    input  [71:0] col_in_79,
    input  [71:0] col_in_80,
    input  [71:0] col_in_81,
    input  [71:0] col_in_82,
    input  [71:0] col_in_83,
    input  [71:0] col_in_84,
    input  [71:0] col_in_85,
    input  [71:0] col_in_86,
    input  [71:0] col_in_87,
    input  [71:0] col_in_88,
    input  [71:0] col_in_89,
    input  [71:0] col_in_90,
    input  [71:0] col_in_91,
    input  [71:0] col_in_92,
    input  [71:0] col_in_93,
    input  [71:0] col_in_94,
    input  [71:0] col_in_95,
    input  [71:0] col_in_96,
    input  [71:0] col_in_97,
    input  [71:0] col_in_98,
    input  [71:0] col_in_99,
    input  [71:0] col_in_100,
    input  [71:0] col_in_101,
    input  [71:0] col_in_102,
    input  [71:0] col_in_103,
    input  [71:0] col_in_104,
    input  [71:0] col_in_105,
    input  [71:0] col_in_106,
    input  [71:0] col_in_107,
    input  [71:0] col_in_108,
    input  [71:0] col_in_109,
    input  [71:0] col_in_110,
    input  [71:0] col_in_111,
    input  [71:0] col_in_112,
    input  [71:0] col_in_113,
    input  [71:0] col_in_114,
    input  [71:0] col_in_115,
    input  [71:0] col_in_116,
    input  [71:0] col_in_117,
    input  [71:0] col_in_118,
    input  [71:0] col_in_119,
    input  [71:0] col_in_120,
    input  [71:0] col_in_121,
    input  [71:0] col_in_122,
    input  [71:0] col_in_123,
    input  [71:0] col_in_124,
    input  [71:0] col_in_125,
    input  [71:0] col_in_126,
    input  [71:0] col_in_127,
    input  [71:0] col_in_128,
    input  [71:0] col_in_129,
    input  [71:0] col_in_130,
    input  [71:0] col_in_131,
    input  [71:0] col_in_132,
    input  [71:0] col_in_133,
    input  [71:0] col_in_134,
    input  [71:0] col_in_135,
    input  [71:0] col_in_136,
    input  [71:0] col_in_137,
    input  [71:0] col_in_138,
    input  [71:0] col_in_139,
    input  [71:0] col_in_140,
    input  [71:0] col_in_141,
    input  [71:0] col_in_142,
    input  [71:0] col_in_143,
    input  [71:0] col_in_144,
    input  [71:0] col_in_145,
    input  [71:0] col_in_146,
    input  [71:0] col_in_147,
    input  [71:0] col_in_148,
    input  [71:0] col_in_149,
    input  [71:0] col_in_150,
    input  [71:0] col_in_151,
    input  [71:0] col_in_152,
    input  [71:0] col_in_153,
    input  [71:0] col_in_154,
    input  [71:0] col_in_155,
    input  [71:0] col_in_156,
    input  [71:0] col_in_157,
    input  [71:0] col_in_158,
    input  [71:0] col_in_159,
    input  [71:0] col_in_160,
    input  [71:0] col_in_161,
    input  [71:0] col_in_162,
    input  [71:0] col_in_163,
    input  [71:0] col_in_164,
    input  [71:0] col_in_165,
    input  [71:0] col_in_166,
    input  [71:0] col_in_167,
    input  [71:0] col_in_168,
    input  [71:0] col_in_169,
    input  [71:0] col_in_170,
    input  [71:0] col_in_171,
    input  [71:0] col_in_172,
    input  [71:0] col_in_173,
    input  [71:0] col_in_174,
    input  [71:0] col_in_175,
    input  [71:0] col_in_176,
    input  [71:0] col_in_177,
    input  [71:0] col_in_178,
    input  [71:0] col_in_179,
    input  [71:0] col_in_180,
    input  [71:0] col_in_181,
    input  [71:0] col_in_182,
    input  [71:0] col_in_183,
    input  [71:0] col_in_184,
    input  [71:0] col_in_185,
    input  [71:0] col_in_186,
    input  [71:0] col_in_187,
    input  [71:0] col_in_188,
    input  [71:0] col_in_189,
    input  [71:0] col_in_190,
    input  [71:0] col_in_191,
    input  [71:0] col_in_192,
    input  [71:0] col_in_193,
    input  [71:0] col_in_194,
    input  [71:0] col_in_195,
    input  [71:0] col_in_196,
    input  [71:0] col_in_197,
    input  [71:0] col_in_198,
    input  [71:0] col_in_199,
    input  [71:0] col_in_200,
    input  [71:0] col_in_201,
    input  [71:0] col_in_202,
    input  [71:0] col_in_203,
    input  [71:0] col_in_204,
    input  [71:0] col_in_205,
    input  [71:0] col_in_206,
    input  [71:0] col_in_207,
    input  [71:0] col_in_208,
    input  [71:0] col_in_209,
    input  [71:0] col_in_210,
    input  [71:0] col_in_211,
    input  [71:0] col_in_212,
    input  [71:0] col_in_213,
    input  [71:0] col_in_214,
    input  [71:0] col_in_215,
    input  [71:0] col_in_216,
    input  [71:0] col_in_217,
    input  [71:0] col_in_218,
    input  [71:0] col_in_219,
    input  [71:0] col_in_220,
    input  [71:0] col_in_221,
    input  [71:0] col_in_222,
    input  [71:0] col_in_223,
    input  [71:0] col_in_224,
    input  [71:0] col_in_225,
    input  [71:0] col_in_226,
    input  [71:0] col_in_227,
    input  [71:0] col_in_228,
    input  [71:0] col_in_229,
    input  [71:0] col_in_230,
    input  [71:0] col_in_231,
    input  [71:0] col_in_232,
    input  [71:0] col_in_233,
    input  [71:0] col_in_234,
    input  [71:0] col_in_235,
    input  [71:0] col_in_236,
    input  [71:0] col_in_237,
    input  [71:0] col_in_238,
    input  [71:0] col_in_239,
    input  [71:0] col_in_240,
    input  [71:0] col_in_241,
    input  [71:0] col_in_242,
    input  [71:0] col_in_243,
    input  [71:0] col_in_244,
    input  [71:0] col_in_245,
    input  [71:0] col_in_246,
    input  [71:0] col_in_247,
    input  [71:0] col_in_248,
    input  [71:0] col_in_249,
    input  [71:0] col_in_250,
    input  [71:0] col_in_251,
    input  [71:0] col_in_252,
    input  [71:0] col_in_253,
    input  [71:0] col_in_254,
    input  [71:0] col_in_255,
    input  [71:0] col_in_256,
    input  [71:0] col_in_257,
    input  [71:0] col_in_258,
    input  [71:0] col_in_259,
    input  [71:0] col_in_260,
    input  [71:0] col_in_261,
    input  [71:0] col_in_262,
    input  [71:0] col_in_263,
    input  [71:0] col_in_264,
    input  [71:0] col_in_265,
    input  [71:0] col_in_266,
    input  [71:0] col_in_267,
    input  [71:0] col_in_268,
    input  [71:0] col_in_269,
    input  [71:0] col_in_270,
    input  [71:0] col_in_271,
    input  [71:0] col_in_272,
    input  [71:0] col_in_273,
    input  [71:0] col_in_274,
    input  [71:0] col_in_275,
    input  [71:0] col_in_276,
    input  [71:0] col_in_277,
    input  [71:0] col_in_278,
    input  [71:0] col_in_279,
    input  [71:0] col_in_280,
    input  [71:0] col_in_281,
    input  [71:0] col_in_282,
    input  [71:0] col_in_283,
    input  [71:0] col_in_284,
    input  [71:0] col_in_285,
    input  [71:0] col_in_286,
    input  [71:0] col_in_287,
    input  [71:0] col_in_288,
    input  [71:0] col_in_289,
    input  [71:0] col_in_290,
    input  [71:0] col_in_291,
    input  [71:0] col_in_292,
    input  [71:0] col_in_293,
    input  [71:0] col_in_294,
    input  [71:0] col_in_295,
    input  [71:0] col_in_296,
    input  [71:0] col_in_297,
    input  [71:0] col_in_298,
    input  [71:0] col_in_299,
    input  [71:0] col_in_300,
    input  [71:0] col_in_301,
    input  [71:0] col_in_302,
    input  [71:0] col_in_303,
    input  [71:0] col_in_304,
    input  [71:0] col_in_305,
    input  [71:0] col_in_306,
    input  [71:0] col_in_307,
    input  [71:0] col_in_308,
    input  [71:0] col_in_309,
    input  [71:0] col_in_310,
    input  [71:0] col_in_311,
    input  [71:0] col_in_312,
    input  [71:0] col_in_313,
    input  [71:0] col_in_314,
    input  [71:0] col_in_315,
    input  [71:0] col_in_316,
    input  [71:0] col_in_317,
    input  [71:0] col_in_318,
    input  [71:0] col_in_319,
    input  [71:0] col_in_320,
    input  [71:0] col_in_321,
    input  [71:0] col_in_322,
    input  [71:0] col_in_323,
    input  [71:0] col_in_324,
    input  [71:0] col_in_325,
    input  [71:0] col_in_326,
    input  [71:0] col_in_327,
    input  [71:0] col_in_328,
    input  [71:0] col_in_329,
    input  [71:0] col_in_330,
    input  [71:0] col_in_331,
    input  [71:0] col_in_332,
    input  [71:0] col_in_333,
    input  [71:0] col_in_334,
    input  [71:0] col_in_335,
    input  [71:0] col_in_336,
    input  [71:0] col_in_337,
    input  [71:0] col_in_338,
    input  [71:0] col_in_339,
    input  [71:0] col_in_340,
    input  [71:0] col_in_341,
    input  [71:0] col_in_342,
    input  [71:0] col_in_343,
    input  [71:0] col_in_344,
    input  [71:0] col_in_345,
    input  [71:0] col_in_346,
    input  [71:0] col_in_347,
    input  [71:0] col_in_348,
    input  [71:0] col_in_349,
    input  [71:0] col_in_350,
    input  [71:0] col_in_351,
    input  [71:0] col_in_352,
    input  [71:0] col_in_353,
    input  [71:0] col_in_354,
    input  [71:0] col_in_355,
    input  [71:0] col_in_356,
    input  [71:0] col_in_357,
    input  [71:0] col_in_358,
    input  [71:0] col_in_359,
    input  [71:0] col_in_360,
    input  [71:0] col_in_361,
    input  [71:0] col_in_362,
    input  [71:0] col_in_363,
    input  [71:0] col_in_364,
    input  [71:0] col_in_365,
    input  [71:0] col_in_366,
    input  [71:0] col_in_367,
    input  [71:0] col_in_368,
    input  [71:0] col_in_369,
    input  [71:0] col_in_370,
    input  [71:0] col_in_371,
    input  [71:0] col_in_372,
    input  [71:0] col_in_373,
    input  [71:0] col_in_374,
    input  [71:0] col_in_375,
    input  [71:0] col_in_376,
    input  [71:0] col_in_377,
    input  [71:0] col_in_378,
    input  [71:0] col_in_379,
    input  [71:0] col_in_380,
    input  [71:0] col_in_381,
    input  [71:0] col_in_382,
    input  [71:0] col_in_383,
    input  [71:0] col_in_384,
    input  [71:0] col_in_385,
    input  [71:0] col_in_386,
    input  [71:0] col_in_387,
    input  [71:0] col_in_388,
    input  [71:0] col_in_389,
    input  [71:0] col_in_390,
    input  [71:0] col_in_391,
    input  [71:0] col_in_392,
    input  [71:0] col_in_393,
    input  [71:0] col_in_394,
    input  [71:0] col_in_395,
    input  [71:0] col_in_396,
    input  [71:0] col_in_397,
    input  [71:0] col_in_398,
    input  [71:0] col_in_399,
    input  [71:0] col_in_400,
    input  [71:0] col_in_401,
    input  [71:0] col_in_402,
    input  [71:0] col_in_403,
    input  [71:0] col_in_404,
    input  [71:0] col_in_405,
    input  [71:0] col_in_406,
    input  [71:0] col_in_407,
    input  [71:0] col_in_408,
    input  [71:0] col_in_409,
    input  [71:0] col_in_410,
    input  [71:0] col_in_411,
    input  [71:0] col_in_412,
    input  [71:0] col_in_413,
    input  [71:0] col_in_414,
    input  [71:0] col_in_415,
    input  [71:0] col_in_416,
    input  [71:0] col_in_417,
    input  [71:0] col_in_418,
    input  [71:0] col_in_419,
    input  [71:0] col_in_420,
    input  [71:0] col_in_421,
    input  [71:0] col_in_422,
    input  [71:0] col_in_423,
    input  [71:0] col_in_424,
    input  [71:0] col_in_425,
    input  [71:0] col_in_426,
    input  [71:0] col_in_427,
    input  [71:0] col_in_428,
    input  [71:0] col_in_429,
    input  [71:0] col_in_430,
    input  [71:0] col_in_431,
    input  [71:0] col_in_432,
    input  [71:0] col_in_433,
    input  [71:0] col_in_434,
    input  [71:0] col_in_435,
    input  [71:0] col_in_436,
    input  [71:0] col_in_437,
    input  [71:0] col_in_438,
    input  [71:0] col_in_439,
    input  [71:0] col_in_440,
    input  [71:0] col_in_441,
    input  [71:0] col_in_442,
    input  [71:0] col_in_443,
    input  [71:0] col_in_444,
    input  [71:0] col_in_445,
    input  [71:0] col_in_446,
    input  [71:0] col_in_447,
    input  [71:0] col_in_448,
    input  [71:0] col_in_449,
    input  [71:0] col_in_450,
    input  [71:0] col_in_451,
    input  [71:0] col_in_452,
    input  [71:0] col_in_453,
    input  [71:0] col_in_454,
    input  [71:0] col_in_455,
    input  [71:0] col_in_456,
    input  [71:0] col_in_457,
    input  [71:0] col_in_458,
    input  [71:0] col_in_459,
    input  [71:0] col_in_460,
    input  [71:0] col_in_461,
    input  [71:0] col_in_462,
    input  [71:0] col_in_463,
    input  [71:0] col_in_464,
    input  [71:0] col_in_465,
    input  [71:0] col_in_466,
    input  [71:0] col_in_467,
    input  [71:0] col_in_468,
    input  [71:0] col_in_469,
    input  [71:0] col_in_470,
    input  [71:0] col_in_471,
    input  [71:0] col_in_472,
    input  [71:0] col_in_473,
    input  [71:0] col_in_474,
    input  [71:0] col_in_475,
    input  [71:0] col_in_476,
    input  [71:0] col_in_477,
    input  [71:0] col_in_478,
    input  [71:0] col_in_479,
    input  [71:0] col_in_480,
    input  [71:0] col_in_481,
    input  [71:0] col_in_482,
    input  [71:0] col_in_483,
    input  [71:0] col_in_484,
    input  [71:0] col_in_485,
    input  [71:0] col_in_486,
    input  [71:0] col_in_487,
    input  [71:0] col_in_488,
    input  [71:0] col_in_489,
    input  [71:0] col_in_490,
    input  [71:0] col_in_491,
    input  [71:0] col_in_492,
    input  [71:0] col_in_493,
    input  [71:0] col_in_494,
    input  [71:0] col_in_495,
    input  [71:0] col_in_496,
    input  [71:0] col_in_497,
    input  [71:0] col_in_498,
    input  [71:0] col_in_499,
    input  [71:0] col_in_500,
    input  [71:0] col_in_501,
    input  [71:0] col_in_502,
    input  [71:0] col_in_503,
    input  [71:0] col_in_504,
    input  [71:0] col_in_505,
    input  [71:0] col_in_506,
    input  [71:0] col_in_507,
    input  [71:0] col_in_508,
    input  [71:0] col_in_509,
    input  [71:0] col_in_510,
    input  [71:0] col_in_511,
    input  [71:0] col_in_512,
    input  [71:0] col_in_513,
    input  [71:0] col_in_514,
    input  [71:0] col_in_515,
    input  [71:0] col_in_516,
    input  [71:0] col_in_517,
    input  [71:0] col_in_518,
    input  [71:0] col_in_519,
    input  [71:0] col_in_520,
    input  [71:0] col_in_521,
    input  [71:0] col_in_522,
    input  [71:0] col_in_523,
    input  [71:0] col_in_524,
    input  [71:0] col_in_525,
    input  [71:0] col_in_526,
    input  [71:0] col_in_527,
    input  [71:0] col_in_528,
    input  [71:0] col_in_529,
    input  [71:0] col_in_530,
    input  [71:0] col_in_531,
    input  [71:0] col_in_532,
    input  [71:0] col_in_533,
    input  [71:0] col_in_534,
    input  [71:0] col_in_535,
    input  [71:0] col_in_536,
    input  [71:0] col_in_537,
    input  [71:0] col_in_538,
    input  [71:0] col_in_539,
    input  [71:0] col_in_540,
    input  [71:0] col_in_541,
    input  [71:0] col_in_542,
    input  [71:0] col_in_543,
    input  [71:0] col_in_544,
    input  [71:0] col_in_545,
    input  [71:0] col_in_546,
    input  [71:0] col_in_547,
    input  [71:0] col_in_548,
    input  [71:0] col_in_549,
    input  [71:0] col_in_550,
    input  [71:0] col_in_551,
    input  [71:0] col_in_552,
    input  [71:0] col_in_553,
    input  [71:0] col_in_554,
    input  [71:0] col_in_555,
    input  [71:0] col_in_556,
    input  [71:0] col_in_557,
    input  [71:0] col_in_558,
    input  [71:0] col_in_559,
    input  [71:0] col_in_560,
    input  [71:0] col_in_561,
    input  [71:0] col_in_562,
    input  [71:0] col_in_563,
    input  [71:0] col_in_564,
    input  [71:0] col_in_565,
    input  [71:0] col_in_566,
    input  [71:0] col_in_567,
    input  [71:0] col_in_568,
    input  [71:0] col_in_569,
    input  [71:0] col_in_570,
    input  [71:0] col_in_571,
    input  [71:0] col_in_572,
    input  [71:0] col_in_573,
    input  [71:0] col_in_574,
    input  [71:0] col_in_575,
    input  [71:0] col_in_576,
    input  [71:0] col_in_577,
    input  [71:0] col_in_578,
    input  [71:0] col_in_579,
    input  [71:0] col_in_580,
    input  [71:0] col_in_581,
    input  [71:0] col_in_582,
    input  [71:0] col_in_583,
    input  [71:0] col_in_584,
    input  [71:0] col_in_585,
    input  [71:0] col_in_586,
    input  [71:0] col_in_587,
    input  [71:0] col_in_588,
    input  [71:0] col_in_589,
    input  [71:0] col_in_590,
    input  [71:0] col_in_591,
    input  [71:0] col_in_592,
    input  [71:0] col_in_593,
    input  [71:0] col_in_594,
    input  [71:0] col_in_595,
    input  [71:0] col_in_596,
    input  [71:0] col_in_597,
    input  [71:0] col_in_598,
    input  [71:0] col_in_599,
    input  [71:0] col_in_600,
    input  [71:0] col_in_601,
    input  [71:0] col_in_602,
    input  [71:0] col_in_603,
    input  [71:0] col_in_604,
    input  [71:0] col_in_605,
    input  [71:0] col_in_606,
    input  [71:0] col_in_607,
    input  [71:0] col_in_608,
    input  [71:0] col_in_609,
    input  [71:0] col_in_610,
    input  [71:0] col_in_611,
    input  [71:0] col_in_612,
    input  [71:0] col_in_613,
    input  [71:0] col_in_614,
    input  [71:0] col_in_615,
    input  [71:0] col_in_616,
    input  [71:0] col_in_617,
    input  [71:0] col_in_618,
    input  [71:0] col_in_619,
    input  [71:0] col_in_620,
    input  [71:0] col_in_621,
    input  [71:0] col_in_622,
    input  [71:0] col_in_623,
    input  [71:0] col_in_624,
    input  [71:0] col_in_625,
    input  [71:0] col_in_626,
    input  [71:0] col_in_627,
    input  [71:0] col_in_628,
    input  [71:0] col_in_629,
    input  [71:0] col_in_630,
    input  [71:0] col_in_631,
    input  [71:0] col_in_632,
    input  [71:0] col_in_633,
    input  [71:0] col_in_634,
    input  [71:0] col_in_635,
    input  [71:0] col_in_636,
    input  [71:0] col_in_637,
    input  [71:0] col_in_638,
    input  [71:0] col_in_639,
    input  [71:0] col_in_640,
    input  [71:0] col_in_641,
    input  [71:0] col_in_642,
    input  [71:0] col_in_643,
    input  [71:0] col_in_644,
    input  [71:0] col_in_645,
    input  [71:0] col_in_646,
    input  [71:0] col_in_647,
    input  [71:0] col_in_648,
    input  [71:0] col_in_649,
    input  [71:0] col_in_650,
    input  [71:0] col_in_651,
    input  [71:0] col_in_652,
    input  [71:0] col_in_653,
    input  [71:0] col_in_654,
    input  [71:0] col_in_655,
    input  [71:0] col_in_656,
    input  [71:0] col_in_657,
    input  [71:0] col_in_658,
    input  [71:0] col_in_659,
    input  [71:0] col_in_660,
    input  [71:0] col_in_661,
    input  [71:0] col_in_662,
    input  [71:0] col_in_663,
    input  [71:0] col_in_664,
    input  [71:0] col_in_665,
    input  [71:0] col_in_666,
    input  [71:0] col_in_667,
    input  [71:0] col_in_668,
    input  [71:0] col_in_669,
    input  [71:0] col_in_670,
    input  [71:0] col_in_671,
    input  [71:0] col_in_672,
    input  [71:0] col_in_673,
    input  [71:0] col_in_674,
    input  [71:0] col_in_675,
    input  [71:0] col_in_676,
    input  [71:0] col_in_677,
    input  [71:0] col_in_678,
    input  [71:0] col_in_679,
    input  [71:0] col_in_680,
    input  [71:0] col_in_681,
    input  [71:0] col_in_682,
    input  [71:0] col_in_683,
    input  [71:0] col_in_684,
    input  [71:0] col_in_685,
    input  [71:0] col_in_686,
    input  [71:0] col_in_687,
    input  [71:0] col_in_688,
    input  [71:0] col_in_689,
    input  [71:0] col_in_690,
    input  [71:0] col_in_691,
    input  [71:0] col_in_692,
    input  [71:0] col_in_693,
    input  [71:0] col_in_694,
    input  [71:0] col_in_695,
    input  [71:0] col_in_696,
    input  [71:0] col_in_697,
    input  [71:0] col_in_698,
    input  [71:0] col_in_699,
    input  [71:0] col_in_700,
    input  [71:0] col_in_701,
    input  [71:0] col_in_702,
    input  [71:0] col_in_703,
    input  [71:0] col_in_704,
    input  [71:0] col_in_705,
    input  [71:0] col_in_706,
    input  [71:0] col_in_707,
    input  [71:0] col_in_708,
    input  [71:0] col_in_709,
    input  [71:0] col_in_710,
    input  [71:0] col_in_711,
    input  [71:0] col_in_712,
    input  [71:0] col_in_713,
    input  [71:0] col_in_714,
    input  [71:0] col_in_715,
    input  [71:0] col_in_716,
    input  [71:0] col_in_717,
    input  [71:0] col_in_718,
    input  [71:0] col_in_719,
    input  [71:0] col_in_720,
    input  [71:0] col_in_721,
    input  [71:0] col_in_722,
    input  [71:0] col_in_723,
    input  [71:0] col_in_724,
    input  [71:0] col_in_725,
    input  [71:0] col_in_726,
    input  [71:0] col_in_727,
    input  [71:0] col_in_728,
    input  [71:0] col_in_729,
    input  [71:0] col_in_730,
    input  [71:0] col_in_731,
    input  [71:0] col_in_732,
    input  [71:0] col_in_733,
    input  [71:0] col_in_734,
    input  [71:0] col_in_735,
    input  [71:0] col_in_736,
    input  [71:0] col_in_737,
    input  [71:0] col_in_738,
    input  [71:0] col_in_739,
    input  [71:0] col_in_740,
    input  [71:0] col_in_741,
    input  [71:0] col_in_742,
    input  [71:0] col_in_743,
    input  [71:0] col_in_744,
    input  [71:0] col_in_745,
    input  [71:0] col_in_746,
    input  [71:0] col_in_747,
    input  [71:0] col_in_748,
    input  [71:0] col_in_749,
    input  [71:0] col_in_750,
    input  [71:0] col_in_751,
    input  [71:0] col_in_752,
    input  [71:0] col_in_753,
    input  [71:0] col_in_754,
    input  [71:0] col_in_755,
    input  [71:0] col_in_756,
    input  [71:0] col_in_757,
    input  [71:0] col_in_758,
    input  [71:0] col_in_759,
    input  [71:0] col_in_760,
    input  [71:0] col_in_761,
    input  [71:0] col_in_762,
    input  [71:0] col_in_763,
    input  [71:0] col_in_764,
    input  [71:0] col_in_765,
    input  [71:0] col_in_766,
    input  [71:0] col_in_767,
    input  [71:0] col_in_768,
    input  [71:0] col_in_769,
    input  [71:0] col_in_770,
    input  [71:0] col_in_771,
    input  [71:0] col_in_772,
    input  [71:0] col_in_773,
    input  [71:0] col_in_774,
    input  [71:0] col_in_775,
    input  [71:0] col_in_776,
    input  [71:0] col_in_777,
    input  [71:0] col_in_778,
    input  [71:0] col_in_779,
    input  [71:0] col_in_780,
    input  [71:0] col_in_781,
    input  [71:0] col_in_782,
    input  [71:0] col_in_783,
    input  [71:0] col_in_784,
    input  [71:0] col_in_785,
    input  [71:0] col_in_786,
    input  [71:0] col_in_787,
    input  [71:0] col_in_788,
    input  [71:0] col_in_789,
    input  [71:0] col_in_790,
    input  [71:0] col_in_791,
    input  [71:0] col_in_792,
    input  [71:0] col_in_793,
    input  [71:0] col_in_794,
    input  [71:0] col_in_795,
    input  [71:0] col_in_796,
    input  [71:0] col_in_797,
    input  [71:0] col_in_798,
    input  [71:0] col_in_799,
    input  [71:0] col_in_800,
    input  [71:0] col_in_801,
    input  [71:0] col_in_802,
    input  [71:0] col_in_803,
    input  [71:0] col_in_804,
    input  [71:0] col_in_805,
    input  [71:0] col_in_806,
    input  [71:0] col_in_807,
    input  [71:0] col_in_808,
    input  [71:0] col_in_809,
    input  [71:0] col_in_810,
    input  [71:0] col_in_811,
    input  [71:0] col_in_812,
    input  [71:0] col_in_813,
    input  [71:0] col_in_814,
    input  [71:0] col_in_815,
    input  [71:0] col_in_816,
    input  [71:0] col_in_817,
    input  [71:0] col_in_818,
    input  [71:0] col_in_819,
    input  [71:0] col_in_820,
    input  [71:0] col_in_821,
    input  [71:0] col_in_822,
    input  [71:0] col_in_823,
    input  [71:0] col_in_824,
    input  [71:0] col_in_825,
    input  [71:0] col_in_826,
    input  [71:0] col_in_827,
    input  [71:0] col_in_828,
    input  [71:0] col_in_829,
    input  [71:0] col_in_830,
    input  [71:0] col_in_831,
    input  [71:0] col_in_832,
    input  [71:0] col_in_833,
    input  [71:0] col_in_834,
    input  [71:0] col_in_835,
    input  [71:0] col_in_836,
    input  [71:0] col_in_837,
    input  [71:0] col_in_838,
    input  [71:0] col_in_839,
    input  [71:0] col_in_840,
    input  [71:0] col_in_841,
    input  [71:0] col_in_842,
    input  [71:0] col_in_843,
    input  [71:0] col_in_844,
    input  [71:0] col_in_845,
    input  [71:0] col_in_846,
    input  [71:0] col_in_847,
    input  [71:0] col_in_848,
    input  [71:0] col_in_849,
    input  [71:0] col_in_850,
    input  [71:0] col_in_851,
    input  [71:0] col_in_852,
    input  [71:0] col_in_853,
    input  [71:0] col_in_854,
    input  [71:0] col_in_855,
    input  [71:0] col_in_856,
    input  [71:0] col_in_857,
    input  [71:0] col_in_858,
    input  [71:0] col_in_859,
    input  [71:0] col_in_860,
    input  [71:0] col_in_861,
    input  [71:0] col_in_862,
    input  [71:0] col_in_863,
    input  [71:0] col_in_864,
    input  [71:0] col_in_865,
    input  [71:0] col_in_866,
    input  [71:0] col_in_867,
    input  [71:0] col_in_868,
    input  [71:0] col_in_869,
    input  [71:0] col_in_870,
    input  [71:0] col_in_871,
    input  [71:0] col_in_872,
    input  [71:0] col_in_873,
    input  [71:0] col_in_874,
    input  [71:0] col_in_875,
    input  [71:0] col_in_876,
    input  [71:0] col_in_877,
    input  [71:0] col_in_878,
    input  [71:0] col_in_879,
    input  [71:0] col_in_880,
    input  [71:0] col_in_881,
    input  [71:0] col_in_882,
    input  [71:0] col_in_883,
    input  [71:0] col_in_884,
    input  [71:0] col_in_885,
    input  [71:0] col_in_886,
    input  [71:0] col_in_887,
    input  [71:0] col_in_888,
    input  [71:0] col_in_889,
    input  [71:0] col_in_890,
    input  [71:0] col_in_891,
    input  [71:0] col_in_892,
    input  [71:0] col_in_893,
    input  [71:0] col_in_894,
    input  [71:0] col_in_895,
    input  [71:0] col_in_896,
    input  [71:0] col_in_897,
    input  [71:0] col_in_898,
    input  [71:0] col_in_899,
    input  [71:0] col_in_900,
    input  [71:0] col_in_901,
    input  [71:0] col_in_902,
    input  [71:0] col_in_903,
    input  [71:0] col_in_904,
    input  [71:0] col_in_905,
    input  [71:0] col_in_906,
    input  [71:0] col_in_907,
    input  [71:0] col_in_908,
    input  [71:0] col_in_909,
    input  [71:0] col_in_910,
    input  [71:0] col_in_911,
    input  [71:0] col_in_912,
    input  [71:0] col_in_913,
    input  [71:0] col_in_914,
    input  [71:0] col_in_915,
    input  [71:0] col_in_916,
    input  [71:0] col_in_917,
    input  [71:0] col_in_918,
    input  [71:0] col_in_919,
    input  [71:0] col_in_920,
    input  [71:0] col_in_921,
    input  [71:0] col_in_922,
    input  [71:0] col_in_923,
    input  [71:0] col_in_924,
    input  [71:0] col_in_925,
    input  [71:0] col_in_926,
    input  [71:0] col_in_927,
    input  [71:0] col_in_928,
    input  [71:0] col_in_929,
    input  [71:0] col_in_930,
    input  [71:0] col_in_931,
    input  [71:0] col_in_932,
    input  [71:0] col_in_933,
    input  [71:0] col_in_934,
    input  [71:0] col_in_935,
    input  [71:0] col_in_936,
    input  [71:0] col_in_937,
    input  [71:0] col_in_938,
    input  [71:0] col_in_939,
    input  [71:0] col_in_940,
    input  [71:0] col_in_941,
    input  [71:0] col_in_942,
    input  [71:0] col_in_943,
    input  [71:0] col_in_944,
    input  [71:0] col_in_945,
    input  [71:0] col_in_946,
    input  [71:0] col_in_947,
    input  [71:0] col_in_948,
    input  [71:0] col_in_949,
    input  [71:0] col_in_950,
    input  [71:0] col_in_951,
    input  [71:0] col_in_952,
    input  [71:0] col_in_953,
    input  [71:0] col_in_954,
    input  [71:0] col_in_955,
    input  [71:0] col_in_956,
    input  [71:0] col_in_957,
    input  [71:0] col_in_958,
    input  [71:0] col_in_959,
    input  [71:0] col_in_960,
    input  [71:0] col_in_961,
    input  [71:0] col_in_962,
    input  [71:0] col_in_963,
    input  [71:0] col_in_964,
    input  [71:0] col_in_965,
    input  [71:0] col_in_966,
    input  [71:0] col_in_967,
    input  [71:0] col_in_968,
    input  [71:0] col_in_969,
    input  [71:0] col_in_970,
    input  [71:0] col_in_971,
    input  [71:0] col_in_972,
    input  [71:0] col_in_973,
    input  [71:0] col_in_974,
    input  [71:0] col_in_975,
    input  [71:0] col_in_976,
    input  [71:0] col_in_977,
    input  [71:0] col_in_978,
    input  [71:0] col_in_979,
    input  [71:0] col_in_980,
    input  [71:0] col_in_981,
    input  [71:0] col_in_982,
    input  [71:0] col_in_983,
    input  [71:0] col_in_984,
    input  [71:0] col_in_985,
    input  [71:0] col_in_986,
    input  [71:0] col_in_987,
    input  [71:0] col_in_988,
    input  [71:0] col_in_989,
    input  [71:0] col_in_990,
    input  [71:0] col_in_991,
    input  [71:0] col_in_992,
    input  [71:0] col_in_993,
    input  [71:0] col_in_994,
    input  [71:0] col_in_995,
    input  [71:0] col_in_996,
    input  [71:0] col_in_997,
    input  [71:0] col_in_998,
    input  [71:0] col_in_999,
    input  [71:0] col_in_1000,
    input  [71:0] col_in_1001,
    input  [71:0] col_in_1002,
    input  [71:0] col_in_1003,
    input  [71:0] col_in_1004,
    input  [71:0] col_in_1005,
    input  [71:0] col_in_1006,
    input  [71:0] col_in_1007,
    input  [71:0] col_in_1008,
    input  [71:0] col_in_1009,
    input  [71:0] col_in_1010,
    input  [71:0] col_in_1011,
    input  [71:0] col_in_1012,
    input  [71:0] col_in_1013,
    input  [71:0] col_in_1014,
    input  [71:0] col_in_1015,
    input  [71:0] col_in_1016,
    input  [71:0] col_in_1017,
    input  [71:0] col_in_1018,
    input  [71:0] col_in_1019,
    input  [71:0] col_in_1020,
    input  [71:0] col_in_1021,
    input  [71:0] col_in_1022,
    input  [71:0] col_in_1023,
    input  [71:0] col_in_1024,
    input  [71:0] col_in_1025,
    input  [71:0] col_in_1026,
    input  [71:0] col_in_1027,
    input  [71:0] col_in_1028,
    input  [71:0] col_in_1029,
    input  [71:0] col_in_1030,
    input  [71:0] col_in_1031,
    input  [71:0] col_in_1032,
    input  [71:0] col_in_1033,
    input  [71:0] col_in_1034,
    input  [71:0] col_in_1035,
    input  [71:0] col_in_1036,
    input  [71:0] col_in_1037,
    input  [71:0] col_in_1038,
    input  [71:0] col_in_1039,
    input  [71:0] col_in_1040,
    input  [71:0] col_in_1041,
    input  [71:0] col_in_1042,
    input  [71:0] col_in_1043,
    input  [71:0] col_in_1044,
    input  [71:0] col_in_1045,
    input  [71:0] col_in_1046,
    input  [71:0] col_in_1047,
    input  [71:0] col_in_1048,
    input  [71:0] col_in_1049,
    input  [71:0] col_in_1050,
    input  [71:0] col_in_1051,
    input  [71:0] col_in_1052,
    input  [71:0] col_in_1053,
    input  [71:0] col_in_1054,
    input  [71:0] col_in_1055,
    input  [71:0] col_in_1056,
    input  [71:0] col_in_1057,
    input  [71:0] col_in_1058,
    input  [71:0] col_in_1059,
    input  [71:0] col_in_1060,
    input  [71:0] col_in_1061,
    input  [71:0] col_in_1062,
    input  [71:0] col_in_1063,
    input  [71:0] col_in_1064,
    input  [71:0] col_in_1065,
    input  [71:0] col_in_1066,
    input  [71:0] col_in_1067,
    input  [71:0] col_in_1068,
    input  [71:0] col_in_1069,
    input  [71:0] col_in_1070,
    input  [71:0] col_in_1071,
    input  [71:0] col_in_1072,
    input  [71:0] col_in_1073,
    input  [71:0] col_in_1074,
    input  [71:0] col_in_1075,
    input  [71:0] col_in_1076,
    input  [71:0] col_in_1077,
    input  [71:0] col_in_1078,
    input  [71:0] col_in_1079,
    input  [71:0] col_in_1080,
    input  [71:0] col_in_1081,
    input  [71:0] col_in_1082,
    input  [71:0] col_in_1083,
    input  [71:0] col_in_1084,
    input  [71:0] col_in_1085,
    input  [71:0] col_in_1086,
    input  [71:0] col_in_1087,
    input  [71:0] col_in_1088,
    input  [71:0] col_in_1089,
    input  [71:0] col_in_1090,
    input  [71:0] col_in_1091,
    input  [71:0] col_in_1092,
    input  [71:0] col_in_1093,
    input  [71:0] col_in_1094,
    input  [71:0] col_in_1095,
    input  [71:0] col_in_1096,
    input  [71:0] col_in_1097,
    input  [71:0] col_in_1098,
    input  [71:0] col_in_1099,
    input  [71:0] col_in_1100,
    input  [71:0] col_in_1101,
    input  [71:0] col_in_1102,
    input  [71:0] col_in_1103,
    input  [71:0] col_in_1104,
    input  [71:0] col_in_1105,
    input  [71:0] col_in_1106,
    input  [71:0] col_in_1107,
    input  [71:0] col_in_1108,
    input  [71:0] col_in_1109,
    input  [71:0] col_in_1110,
    input  [71:0] col_in_1111,
    input  [71:0] col_in_1112,
    input  [71:0] col_in_1113,
    input  [71:0] col_in_1114,
    input  [71:0] col_in_1115,
    input  [71:0] col_in_1116,
    input  [71:0] col_in_1117,
    input  [71:0] col_in_1118,
    input  [71:0] col_in_1119,
    input  [71:0] col_in_1120,
    input  [71:0] col_in_1121,
    input  [71:0] col_in_1122,
    input  [71:0] col_in_1123,
    input  [71:0] col_in_1124,
    input  [71:0] col_in_1125,
    input  [71:0] col_in_1126,
    input  [71:0] col_in_1127,
    input  [71:0] col_in_1128,
    input  [71:0] col_in_1129,
    input  [71:0] col_in_1130,
    input  [71:0] col_in_1131,
    input  [71:0] col_in_1132,
    input  [71:0] col_in_1133,
    input  [71:0] col_in_1134,
    input  [71:0] col_in_1135,
    input  [71:0] col_in_1136,
    input  [71:0] col_in_1137,
    input  [71:0] col_in_1138,
    input  [71:0] col_in_1139,
    input  [71:0] col_in_1140,
    input  [71:0] col_in_1141,
    input  [71:0] col_in_1142,
    input  [71:0] col_in_1143,
    input  [71:0] col_in_1144,
    input  [71:0] col_in_1145,
    input  [71:0] col_in_1146,
    input  [71:0] col_in_1147,
    input  [71:0] col_in_1148,
    input  [71:0] col_in_1149,
    input  [71:0] col_in_1150,
    input  [71:0] col_in_1151,
    input  [71:0] col_in_1152,
    input  [71:0] col_in_1153,
    input  [71:0] col_in_1154,
    input  [71:0] col_in_1155,
    input  [71:0] col_in_1156,
    input  [71:0] col_in_1157,
    input  [71:0] col_in_1158,
    input  [71:0] col_in_1159,
    input  [71:0] col_in_1160,
    input  [71:0] col_in_1161,
    input  [71:0] col_in_1162,
    input  [71:0] col_in_1163,
    input  [71:0] col_in_1164,
    input  [71:0] col_in_1165,
    input  [71:0] col_in_1166,
    input  [71:0] col_in_1167,
    input  [71:0] col_in_1168,
    input  [71:0] col_in_1169,
    input  [71:0] col_in_1170,
    input  [71:0] col_in_1171,
    input  [71:0] col_in_1172,
    input  [71:0] col_in_1173,
    input  [71:0] col_in_1174,
    input  [71:0] col_in_1175,
    input  [71:0] col_in_1176,
    input  [71:0] col_in_1177,
    input  [71:0] col_in_1178,
    input  [71:0] col_in_1179,
    input  [71:0] col_in_1180,
    input  [71:0] col_in_1181,
    input  [71:0] col_in_1182,
    input  [71:0] col_in_1183,
    input  [71:0] col_in_1184,
    input  [71:0] col_in_1185,
    input  [71:0] col_in_1186,
    input  [71:0] col_in_1187,
    input  [71:0] col_in_1188,
    input  [71:0] col_in_1189,
    input  [71:0] col_in_1190,
    input  [71:0] col_in_1191,
    input  [71:0] col_in_1192,
    input  [71:0] col_in_1193,
    input  [71:0] col_in_1194,
    input  [71:0] col_in_1195,
    input  [71:0] col_in_1196,
    input  [71:0] col_in_1197,
    input  [71:0] col_in_1198,
    input  [71:0] col_in_1199,
    input  [71:0] col_in_1200,
    input  [71:0] col_in_1201,
    input  [71:0] col_in_1202,
    input  [71:0] col_in_1203,
    input  [71:0] col_in_1204,
    input  [71:0] col_in_1205,
    input  [71:0] col_in_1206,
    input  [71:0] col_in_1207,
    input  [71:0] col_in_1208,
    input  [71:0] col_in_1209,
    input  [71:0] col_in_1210,
    input  [71:0] col_in_1211,
    input  [71:0] col_in_1212,
    input  [71:0] col_in_1213,
    input  [71:0] col_in_1214,
    input  [71:0] col_in_1215,
    input  [71:0] col_in_1216,
    input  [71:0] col_in_1217,
    input  [71:0] col_in_1218,
    input  [71:0] col_in_1219,
    input  [71:0] col_in_1220,
    input  [71:0] col_in_1221,
    input  [71:0] col_in_1222,
    input  [71:0] col_in_1223,
    input  [71:0] col_in_1224,
    input  [71:0] col_in_1225,
    input  [71:0] col_in_1226,
    input  [71:0] col_in_1227,
    input  [71:0] col_in_1228,
    input  [71:0] col_in_1229,
    input  [71:0] col_in_1230,
    input  [71:0] col_in_1231,
    input  [71:0] col_in_1232,
    input  [71:0] col_in_1233,
    input  [71:0] col_in_1234,
    input  [71:0] col_in_1235,
    input  [71:0] col_in_1236,
    input  [71:0] col_in_1237,
    input  [71:0] col_in_1238,
    input  [71:0] col_in_1239,
    input  [71:0] col_in_1240,
    input  [71:0] col_in_1241,
    input  [71:0] col_in_1242,
    input  [71:0] col_in_1243,
    input  [71:0] col_in_1244,
    input  [71:0] col_in_1245,
    input  [71:0] col_in_1246,
    input  [71:0] col_in_1247,
    input  [71:0] col_in_1248,
    input  [71:0] col_in_1249,
    input  [71:0] col_in_1250,
    input  [71:0] col_in_1251,
    input  [71:0] col_in_1252,
    input  [71:0] col_in_1253,
    input  [71:0] col_in_1254,
    input  [71:0] col_in_1255,
    input  [71:0] col_in_1256,
    input  [71:0] col_in_1257,
    input  [71:0] col_in_1258,
    input  [71:0] col_in_1259,
    input  [71:0] col_in_1260,
    input  [71:0] col_in_1261,
    input  [71:0] col_in_1262,
    input  [71:0] col_in_1263,
    input  [71:0] col_in_1264,
    input  [71:0] col_in_1265,
    input  [71:0] col_in_1266,
    input  [71:0] col_in_1267,
    input  [71:0] col_in_1268,
    input  [71:0] col_in_1269,
    input  [71:0] col_in_1270,
    input  [71:0] col_in_1271,
    input  [71:0] col_in_1272,
    input  [71:0] col_in_1273,
    input  [71:0] col_in_1274,
    input  [71:0] col_in_1275,
    input  [71:0] col_in_1276,
    input  [71:0] col_in_1277,
    input  [71:0] col_in_1278,
    input  [71:0] col_in_1279,
    input  [71:0] col_in_1280,
    input  [71:0] col_in_1281,
    input  [71:0] col_in_1282,

    output [23:0] col_out_0,
    output [23:0] col_out_1,
    output [23:0] col_out_2,
    output [23:0] col_out_3,
    output [23:0] col_out_4,
    output [23:0] col_out_5,
    output [23:0] col_out_6,
    output [23:0] col_out_7,
    output [23:0] col_out_8,
    output [23:0] col_out_9,
    output [23:0] col_out_10,
    output [23:0] col_out_11,
    output [23:0] col_out_12,
    output [23:0] col_out_13,
    output [23:0] col_out_14,
    output [23:0] col_out_15,
    output [23:0] col_out_16,
    output [23:0] col_out_17,
    output [23:0] col_out_18,
    output [23:0] col_out_19,
    output [23:0] col_out_20,
    output [23:0] col_out_21,
    output [23:0] col_out_22,
    output [23:0] col_out_23,
    output [23:0] col_out_24,
    output [23:0] col_out_25,
    output [23:0] col_out_26,
    output [23:0] col_out_27,
    output [23:0] col_out_28,
    output [23:0] col_out_29,
    output [23:0] col_out_30,
    output [23:0] col_out_31,
    output [23:0] col_out_32,
    output [23:0] col_out_33,
    output [23:0] col_out_34,
    output [23:0] col_out_35,
    output [23:0] col_out_36,
    output [23:0] col_out_37,
    output [23:0] col_out_38,
    output [23:0] col_out_39,
    output [23:0] col_out_40,
    output [23:0] col_out_41,
    output [23:0] col_out_42,
    output [23:0] col_out_43,
    output [23:0] col_out_44,
    output [23:0] col_out_45,
    output [23:0] col_out_46,
    output [23:0] col_out_47,
    output [23:0] col_out_48,
    output [23:0] col_out_49,
    output [23:0] col_out_50,
    output [23:0] col_out_51,
    output [23:0] col_out_52,
    output [23:0] col_out_53,
    output [23:0] col_out_54,
    output [23:0] col_out_55,
    output [23:0] col_out_56,
    output [23:0] col_out_57,
    output [23:0] col_out_58,
    output [23:0] col_out_59,
    output [23:0] col_out_60,
    output [23:0] col_out_61,
    output [23:0] col_out_62,
    output [23:0] col_out_63,
    output [23:0] col_out_64,
    output [23:0] col_out_65,
    output [23:0] col_out_66,
    output [23:0] col_out_67,
    output [23:0] col_out_68,
    output [23:0] col_out_69,
    output [23:0] col_out_70,
    output [23:0] col_out_71,
    output [23:0] col_out_72,
    output [23:0] col_out_73,
    output [23:0] col_out_74,
    output [23:0] col_out_75,
    output [23:0] col_out_76,
    output [23:0] col_out_77,
    output [23:0] col_out_78,
    output [23:0] col_out_79,
    output [23:0] col_out_80,
    output [23:0] col_out_81,
    output [23:0] col_out_82,
    output [23:0] col_out_83,
    output [23:0] col_out_84,
    output [23:0] col_out_85,
    output [23:0] col_out_86,
    output [23:0] col_out_87,
    output [23:0] col_out_88,
    output [23:0] col_out_89,
    output [23:0] col_out_90,
    output [23:0] col_out_91,
    output [23:0] col_out_92,
    output [23:0] col_out_93,
    output [23:0] col_out_94,
    output [23:0] col_out_95,
    output [23:0] col_out_96,
    output [23:0] col_out_97,
    output [23:0] col_out_98,
    output [23:0] col_out_99,
    output [23:0] col_out_100,
    output [23:0] col_out_101,
    output [23:0] col_out_102,
    output [23:0] col_out_103,
    output [23:0] col_out_104,
    output [23:0] col_out_105,
    output [23:0] col_out_106,
    output [23:0] col_out_107,
    output [23:0] col_out_108,
    output [23:0] col_out_109,
    output [23:0] col_out_110,
    output [23:0] col_out_111,
    output [23:0] col_out_112,
    output [23:0] col_out_113,
    output [23:0] col_out_114,
    output [23:0] col_out_115,
    output [23:0] col_out_116,
    output [23:0] col_out_117,
    output [23:0] col_out_118,
    output [23:0] col_out_119,
    output [23:0] col_out_120,
    output [23:0] col_out_121,
    output [23:0] col_out_122,
    output [23:0] col_out_123,
    output [23:0] col_out_124,
    output [23:0] col_out_125,
    output [23:0] col_out_126,
    output [23:0] col_out_127,
    output [23:0] col_out_128,
    output [23:0] col_out_129,
    output [23:0] col_out_130,
    output [23:0] col_out_131,
    output [23:0] col_out_132,
    output [23:0] col_out_133,
    output [23:0] col_out_134,
    output [23:0] col_out_135,
    output [23:0] col_out_136,
    output [23:0] col_out_137,
    output [23:0] col_out_138,
    output [23:0] col_out_139,
    output [23:0] col_out_140,
    output [23:0] col_out_141,
    output [23:0] col_out_142,
    output [23:0] col_out_143,
    output [23:0] col_out_144,
    output [23:0] col_out_145,
    output [23:0] col_out_146,
    output [23:0] col_out_147,
    output [23:0] col_out_148,
    output [23:0] col_out_149,
    output [23:0] col_out_150,
    output [23:0] col_out_151,
    output [23:0] col_out_152,
    output [23:0] col_out_153,
    output [23:0] col_out_154,
    output [23:0] col_out_155,
    output [23:0] col_out_156,
    output [23:0] col_out_157,
    output [23:0] col_out_158,
    output [23:0] col_out_159,
    output [23:0] col_out_160,
    output [23:0] col_out_161,
    output [23:0] col_out_162,
    output [23:0] col_out_163,
    output [23:0] col_out_164,
    output [23:0] col_out_165,
    output [23:0] col_out_166,
    output [23:0] col_out_167,
    output [23:0] col_out_168,
    output [23:0] col_out_169,
    output [23:0] col_out_170,
    output [23:0] col_out_171,
    output [23:0] col_out_172,
    output [23:0] col_out_173,
    output [23:0] col_out_174,
    output [23:0] col_out_175,
    output [23:0] col_out_176,
    output [23:0] col_out_177,
    output [23:0] col_out_178,
    output [23:0] col_out_179,
    output [23:0] col_out_180,
    output [23:0] col_out_181,
    output [23:0] col_out_182,
    output [23:0] col_out_183,
    output [23:0] col_out_184,
    output [23:0] col_out_185,
    output [23:0] col_out_186,
    output [23:0] col_out_187,
    output [23:0] col_out_188,
    output [23:0] col_out_189,
    output [23:0] col_out_190,
    output [23:0] col_out_191,
    output [23:0] col_out_192,
    output [23:0] col_out_193,
    output [23:0] col_out_194,
    output [23:0] col_out_195,
    output [23:0] col_out_196,
    output [23:0] col_out_197,
    output [23:0] col_out_198,
    output [23:0] col_out_199,
    output [23:0] col_out_200,
    output [23:0] col_out_201,
    output [23:0] col_out_202,
    output [23:0] col_out_203,
    output [23:0] col_out_204,
    output [23:0] col_out_205,
    output [23:0] col_out_206,
    output [23:0] col_out_207,
    output [23:0] col_out_208,
    output [23:0] col_out_209,
    output [23:0] col_out_210,
    output [23:0] col_out_211,
    output [23:0] col_out_212,
    output [23:0] col_out_213,
    output [23:0] col_out_214,
    output [23:0] col_out_215,
    output [23:0] col_out_216,
    output [23:0] col_out_217,
    output [23:0] col_out_218,
    output [23:0] col_out_219,
    output [23:0] col_out_220,
    output [23:0] col_out_221,
    output [23:0] col_out_222,
    output [23:0] col_out_223,
    output [23:0] col_out_224,
    output [23:0] col_out_225,
    output [23:0] col_out_226,
    output [23:0] col_out_227,
    output [23:0] col_out_228,
    output [23:0] col_out_229,
    output [23:0] col_out_230,
    output [23:0] col_out_231,
    output [23:0] col_out_232,
    output [23:0] col_out_233,
    output [23:0] col_out_234,
    output [23:0] col_out_235,
    output [23:0] col_out_236,
    output [23:0] col_out_237,
    output [23:0] col_out_238,
    output [23:0] col_out_239,
    output [23:0] col_out_240,
    output [23:0] col_out_241,
    output [23:0] col_out_242,
    output [23:0] col_out_243,
    output [23:0] col_out_244,
    output [23:0] col_out_245,
    output [23:0] col_out_246,
    output [23:0] col_out_247,
    output [23:0] col_out_248,
    output [23:0] col_out_249,
    output [23:0] col_out_250,
    output [23:0] col_out_251,
    output [23:0] col_out_252,
    output [23:0] col_out_253,
    output [23:0] col_out_254,
    output [23:0] col_out_255,
    output [23:0] col_out_256,
    output [23:0] col_out_257,
    output [23:0] col_out_258,
    output [23:0] col_out_259,
    output [23:0] col_out_260,
    output [23:0] col_out_261,
    output [23:0] col_out_262,
    output [23:0] col_out_263,
    output [23:0] col_out_264,
    output [23:0] col_out_265,
    output [23:0] col_out_266,
    output [23:0] col_out_267,
    output [23:0] col_out_268,
    output [23:0] col_out_269,
    output [23:0] col_out_270,
    output [23:0] col_out_271,
    output [23:0] col_out_272,
    output [23:0] col_out_273,
    output [23:0] col_out_274,
    output [23:0] col_out_275,
    output [23:0] col_out_276,
    output [23:0] col_out_277,
    output [23:0] col_out_278,
    output [23:0] col_out_279,
    output [23:0] col_out_280,
    output [23:0] col_out_281,
    output [23:0] col_out_282,
    output [23:0] col_out_283,
    output [23:0] col_out_284,
    output [23:0] col_out_285,
    output [23:0] col_out_286,
    output [23:0] col_out_287,
    output [23:0] col_out_288,
    output [23:0] col_out_289,
    output [23:0] col_out_290,
    output [23:0] col_out_291,
    output [23:0] col_out_292,
    output [23:0] col_out_293,
    output [23:0] col_out_294,
    output [23:0] col_out_295,
    output [23:0] col_out_296,
    output [23:0] col_out_297,
    output [23:0] col_out_298,
    output [23:0] col_out_299,
    output [23:0] col_out_300,
    output [23:0] col_out_301,
    output [23:0] col_out_302,
    output [23:0] col_out_303,
    output [23:0] col_out_304,
    output [23:0] col_out_305,
    output [23:0] col_out_306,
    output [23:0] col_out_307,
    output [23:0] col_out_308,
    output [23:0] col_out_309,
    output [23:0] col_out_310,
    output [23:0] col_out_311,
    output [23:0] col_out_312,
    output [23:0] col_out_313,
    output [23:0] col_out_314,
    output [23:0] col_out_315,
    output [23:0] col_out_316,
    output [23:0] col_out_317,
    output [23:0] col_out_318,
    output [23:0] col_out_319,
    output [23:0] col_out_320,
    output [23:0] col_out_321,
    output [23:0] col_out_322,
    output [23:0] col_out_323,
    output [23:0] col_out_324,
    output [23:0] col_out_325,
    output [23:0] col_out_326,
    output [23:0] col_out_327,
    output [23:0] col_out_328,
    output [23:0] col_out_329,
    output [23:0] col_out_330,
    output [23:0] col_out_331,
    output [23:0] col_out_332,
    output [23:0] col_out_333,
    output [23:0] col_out_334,
    output [23:0] col_out_335,
    output [23:0] col_out_336,
    output [23:0] col_out_337,
    output [23:0] col_out_338,
    output [23:0] col_out_339,
    output [23:0] col_out_340,
    output [23:0] col_out_341,
    output [23:0] col_out_342,
    output [23:0] col_out_343,
    output [23:0] col_out_344,
    output [23:0] col_out_345,
    output [23:0] col_out_346,
    output [23:0] col_out_347,
    output [23:0] col_out_348,
    output [23:0] col_out_349,
    output [23:0] col_out_350,
    output [23:0] col_out_351,
    output [23:0] col_out_352,
    output [23:0] col_out_353,
    output [23:0] col_out_354,
    output [23:0] col_out_355,
    output [23:0] col_out_356,
    output [23:0] col_out_357,
    output [23:0] col_out_358,
    output [23:0] col_out_359,
    output [23:0] col_out_360,
    output [23:0] col_out_361,
    output [23:0] col_out_362,
    output [23:0] col_out_363,
    output [23:0] col_out_364,
    output [23:0] col_out_365,
    output [23:0] col_out_366,
    output [23:0] col_out_367,
    output [23:0] col_out_368,
    output [23:0] col_out_369,
    output [23:0] col_out_370,
    output [23:0] col_out_371,
    output [23:0] col_out_372,
    output [23:0] col_out_373,
    output [23:0] col_out_374,
    output [23:0] col_out_375,
    output [23:0] col_out_376,
    output [23:0] col_out_377,
    output [23:0] col_out_378,
    output [23:0] col_out_379,
    output [23:0] col_out_380,
    output [23:0] col_out_381,
    output [23:0] col_out_382,
    output [23:0] col_out_383,
    output [23:0] col_out_384,
    output [23:0] col_out_385,
    output [23:0] col_out_386,
    output [23:0] col_out_387,
    output [23:0] col_out_388,
    output [23:0] col_out_389,
    output [23:0] col_out_390,
    output [23:0] col_out_391,
    output [23:0] col_out_392,
    output [23:0] col_out_393,
    output [23:0] col_out_394,
    output [23:0] col_out_395,
    output [23:0] col_out_396,
    output [23:0] col_out_397,
    output [23:0] col_out_398,
    output [23:0] col_out_399,
    output [23:0] col_out_400,
    output [23:0] col_out_401,
    output [23:0] col_out_402,
    output [23:0] col_out_403,
    output [23:0] col_out_404,
    output [23:0] col_out_405,
    output [23:0] col_out_406,
    output [23:0] col_out_407,
    output [23:0] col_out_408,
    output [23:0] col_out_409,
    output [23:0] col_out_410,
    output [23:0] col_out_411,
    output [23:0] col_out_412,
    output [23:0] col_out_413,
    output [23:0] col_out_414,
    output [23:0] col_out_415,
    output [23:0] col_out_416,
    output [23:0] col_out_417,
    output [23:0] col_out_418,
    output [23:0] col_out_419,
    output [23:0] col_out_420,
    output [23:0] col_out_421,
    output [23:0] col_out_422,
    output [23:0] col_out_423,
    output [23:0] col_out_424,
    output [23:0] col_out_425,
    output [23:0] col_out_426,
    output [23:0] col_out_427,
    output [23:0] col_out_428,
    output [23:0] col_out_429,
    output [23:0] col_out_430,
    output [23:0] col_out_431,
    output [23:0] col_out_432,
    output [23:0] col_out_433,
    output [23:0] col_out_434,
    output [23:0] col_out_435,
    output [23:0] col_out_436,
    output [23:0] col_out_437,
    output [23:0] col_out_438,
    output [23:0] col_out_439,
    output [23:0] col_out_440,
    output [23:0] col_out_441,
    output [23:0] col_out_442,
    output [23:0] col_out_443,
    output [23:0] col_out_444,
    output [23:0] col_out_445,
    output [23:0] col_out_446,
    output [23:0] col_out_447,
    output [23:0] col_out_448,
    output [23:0] col_out_449,
    output [23:0] col_out_450,
    output [23:0] col_out_451,
    output [23:0] col_out_452,
    output [23:0] col_out_453,
    output [23:0] col_out_454,
    output [23:0] col_out_455,
    output [23:0] col_out_456,
    output [23:0] col_out_457,
    output [23:0] col_out_458,
    output [23:0] col_out_459,
    output [23:0] col_out_460,
    output [23:0] col_out_461,
    output [23:0] col_out_462,
    output [23:0] col_out_463,
    output [23:0] col_out_464,
    output [23:0] col_out_465,
    output [23:0] col_out_466,
    output [23:0] col_out_467,
    output [23:0] col_out_468,
    output [23:0] col_out_469,
    output [23:0] col_out_470,
    output [23:0] col_out_471,
    output [23:0] col_out_472,
    output [23:0] col_out_473,
    output [23:0] col_out_474,
    output [23:0] col_out_475,
    output [23:0] col_out_476,
    output [23:0] col_out_477,
    output [23:0] col_out_478,
    output [23:0] col_out_479,
    output [23:0] col_out_480,
    output [23:0] col_out_481,
    output [23:0] col_out_482,
    output [23:0] col_out_483,
    output [23:0] col_out_484,
    output [23:0] col_out_485,
    output [23:0] col_out_486,
    output [23:0] col_out_487,
    output [23:0] col_out_488,
    output [23:0] col_out_489,
    output [23:0] col_out_490,
    output [23:0] col_out_491,
    output [23:0] col_out_492,
    output [23:0] col_out_493,
    output [23:0] col_out_494,
    output [23:0] col_out_495,
    output [23:0] col_out_496,
    output [23:0] col_out_497,
    output [23:0] col_out_498,
    output [23:0] col_out_499,
    output [23:0] col_out_500,
    output [23:0] col_out_501,
    output [23:0] col_out_502,
    output [23:0] col_out_503,
    output [23:0] col_out_504,
    output [23:0] col_out_505,
    output [23:0] col_out_506,
    output [23:0] col_out_507,
    output [23:0] col_out_508,
    output [23:0] col_out_509,
    output [23:0] col_out_510,
    output [23:0] col_out_511,
    output [23:0] col_out_512,
    output [23:0] col_out_513,
    output [23:0] col_out_514,
    output [23:0] col_out_515,
    output [23:0] col_out_516,
    output [23:0] col_out_517,
    output [23:0] col_out_518,
    output [23:0] col_out_519,
    output [23:0] col_out_520,
    output [23:0] col_out_521,
    output [23:0] col_out_522,
    output [23:0] col_out_523,
    output [23:0] col_out_524,
    output [23:0] col_out_525,
    output [23:0] col_out_526,
    output [23:0] col_out_527,
    output [23:0] col_out_528,
    output [23:0] col_out_529,
    output [23:0] col_out_530,
    output [23:0] col_out_531,
    output [23:0] col_out_532,
    output [23:0] col_out_533,
    output [23:0] col_out_534,
    output [23:0] col_out_535,
    output [23:0] col_out_536,
    output [23:0] col_out_537,
    output [23:0] col_out_538,
    output [23:0] col_out_539,
    output [23:0] col_out_540,
    output [23:0] col_out_541,
    output [23:0] col_out_542,
    output [23:0] col_out_543,
    output [23:0] col_out_544,
    output [23:0] col_out_545,
    output [23:0] col_out_546,
    output [23:0] col_out_547,
    output [23:0] col_out_548,
    output [23:0] col_out_549,
    output [23:0] col_out_550,
    output [23:0] col_out_551,
    output [23:0] col_out_552,
    output [23:0] col_out_553,
    output [23:0] col_out_554,
    output [23:0] col_out_555,
    output [23:0] col_out_556,
    output [23:0] col_out_557,
    output [23:0] col_out_558,
    output [23:0] col_out_559,
    output [23:0] col_out_560,
    output [23:0] col_out_561,
    output [23:0] col_out_562,
    output [23:0] col_out_563,
    output [23:0] col_out_564,
    output [23:0] col_out_565,
    output [23:0] col_out_566,
    output [23:0] col_out_567,
    output [23:0] col_out_568,
    output [23:0] col_out_569,
    output [23:0] col_out_570,
    output [23:0] col_out_571,
    output [23:0] col_out_572,
    output [23:0] col_out_573,
    output [23:0] col_out_574,
    output [23:0] col_out_575,
    output [23:0] col_out_576,
    output [23:0] col_out_577,
    output [23:0] col_out_578,
    output [23:0] col_out_579,
    output [23:0] col_out_580,
    output [23:0] col_out_581,
    output [23:0] col_out_582,
    output [23:0] col_out_583,
    output [23:0] col_out_584,
    output [23:0] col_out_585,
    output [23:0] col_out_586,
    output [23:0] col_out_587,
    output [23:0] col_out_588,
    output [23:0] col_out_589,
    output [23:0] col_out_590,
    output [23:0] col_out_591,
    output [23:0] col_out_592,
    output [23:0] col_out_593,
    output [23:0] col_out_594,
    output [23:0] col_out_595,
    output [23:0] col_out_596,
    output [23:0] col_out_597,
    output [23:0] col_out_598,
    output [23:0] col_out_599,
    output [23:0] col_out_600,
    output [23:0] col_out_601,
    output [23:0] col_out_602,
    output [23:0] col_out_603,
    output [23:0] col_out_604,
    output [23:0] col_out_605,
    output [23:0] col_out_606,
    output [23:0] col_out_607,
    output [23:0] col_out_608,
    output [23:0] col_out_609,
    output [23:0] col_out_610,
    output [23:0] col_out_611,
    output [23:0] col_out_612,
    output [23:0] col_out_613,
    output [23:0] col_out_614,
    output [23:0] col_out_615,
    output [23:0] col_out_616,
    output [23:0] col_out_617,
    output [23:0] col_out_618,
    output [23:0] col_out_619,
    output [23:0] col_out_620,
    output [23:0] col_out_621,
    output [23:0] col_out_622,
    output [23:0] col_out_623,
    output [23:0] col_out_624,
    output [23:0] col_out_625,
    output [23:0] col_out_626,
    output [23:0] col_out_627,
    output [23:0] col_out_628,
    output [23:0] col_out_629,
    output [23:0] col_out_630,
    output [23:0] col_out_631,
    output [23:0] col_out_632,
    output [23:0] col_out_633,
    output [23:0] col_out_634,
    output [23:0] col_out_635,
    output [23:0] col_out_636,
    output [23:0] col_out_637,
    output [23:0] col_out_638,
    output [23:0] col_out_639,
    output [23:0] col_out_640,
    output [23:0] col_out_641,
    output [23:0] col_out_642,
    output [23:0] col_out_643,
    output [23:0] col_out_644,
    output [23:0] col_out_645,
    output [23:0] col_out_646,
    output [23:0] col_out_647,
    output [23:0] col_out_648,
    output [23:0] col_out_649,
    output [23:0] col_out_650,
    output [23:0] col_out_651,
    output [23:0] col_out_652,
    output [23:0] col_out_653,
    output [23:0] col_out_654,
    output [23:0] col_out_655,
    output [23:0] col_out_656,
    output [23:0] col_out_657,
    output [23:0] col_out_658,
    output [23:0] col_out_659,
    output [23:0] col_out_660,
    output [23:0] col_out_661,
    output [23:0] col_out_662,
    output [23:0] col_out_663,
    output [23:0] col_out_664,
    output [23:0] col_out_665,
    output [23:0] col_out_666,
    output [23:0] col_out_667,
    output [23:0] col_out_668,
    output [23:0] col_out_669,
    output [23:0] col_out_670,
    output [23:0] col_out_671,
    output [23:0] col_out_672,
    output [23:0] col_out_673,
    output [23:0] col_out_674,
    output [23:0] col_out_675,
    output [23:0] col_out_676,
    output [23:0] col_out_677,
    output [23:0] col_out_678,
    output [23:0] col_out_679,
    output [23:0] col_out_680,
    output [23:0] col_out_681,
    output [23:0] col_out_682,
    output [23:0] col_out_683,
    output [23:0] col_out_684,
    output [23:0] col_out_685,
    output [23:0] col_out_686,
    output [23:0] col_out_687,
    output [23:0] col_out_688,
    output [23:0] col_out_689,
    output [23:0] col_out_690,
    output [23:0] col_out_691,
    output [23:0] col_out_692,
    output [23:0] col_out_693,
    output [23:0] col_out_694,
    output [23:0] col_out_695,
    output [23:0] col_out_696,
    output [23:0] col_out_697,
    output [23:0] col_out_698,
    output [23:0] col_out_699,
    output [23:0] col_out_700,
    output [23:0] col_out_701,
    output [23:0] col_out_702,
    output [23:0] col_out_703,
    output [23:0] col_out_704,
    output [23:0] col_out_705,
    output [23:0] col_out_706,
    output [23:0] col_out_707,
    output [23:0] col_out_708,
    output [23:0] col_out_709,
    output [23:0] col_out_710,
    output [23:0] col_out_711,
    output [23:0] col_out_712,
    output [23:0] col_out_713,
    output [23:0] col_out_714,
    output [23:0] col_out_715,
    output [23:0] col_out_716,
    output [23:0] col_out_717,
    output [23:0] col_out_718,
    output [23:0] col_out_719,
    output [23:0] col_out_720,
    output [23:0] col_out_721,
    output [23:0] col_out_722,
    output [23:0] col_out_723,
    output [23:0] col_out_724,
    output [23:0] col_out_725,
    output [23:0] col_out_726,
    output [23:0] col_out_727,
    output [23:0] col_out_728,
    output [23:0] col_out_729,
    output [23:0] col_out_730,
    output [23:0] col_out_731,
    output [23:0] col_out_732,
    output [23:0] col_out_733,
    output [23:0] col_out_734,
    output [23:0] col_out_735,
    output [23:0] col_out_736,
    output [23:0] col_out_737,
    output [23:0] col_out_738,
    output [23:0] col_out_739,
    output [23:0] col_out_740,
    output [23:0] col_out_741,
    output [23:0] col_out_742,
    output [23:0] col_out_743,
    output [23:0] col_out_744,
    output [23:0] col_out_745,
    output [23:0] col_out_746,
    output [23:0] col_out_747,
    output [23:0] col_out_748,
    output [23:0] col_out_749,
    output [23:0] col_out_750,
    output [23:0] col_out_751,
    output [23:0] col_out_752,
    output [23:0] col_out_753,
    output [23:0] col_out_754,
    output [23:0] col_out_755,
    output [23:0] col_out_756,
    output [23:0] col_out_757,
    output [23:0] col_out_758,
    output [23:0] col_out_759,
    output [23:0] col_out_760,
    output [23:0] col_out_761,
    output [23:0] col_out_762,
    output [23:0] col_out_763,
    output [23:0] col_out_764,
    output [23:0] col_out_765,
    output [23:0] col_out_766,
    output [23:0] col_out_767,
    output [23:0] col_out_768,
    output [23:0] col_out_769,
    output [23:0] col_out_770,
    output [23:0] col_out_771,
    output [23:0] col_out_772,
    output [23:0] col_out_773,
    output [23:0] col_out_774,
    output [23:0] col_out_775,
    output [23:0] col_out_776,
    output [23:0] col_out_777,
    output [23:0] col_out_778,
    output [23:0] col_out_779,
    output [23:0] col_out_780,
    output [23:0] col_out_781,
    output [23:0] col_out_782,
    output [23:0] col_out_783,
    output [23:0] col_out_784,
    output [23:0] col_out_785,
    output [23:0] col_out_786,
    output [23:0] col_out_787,
    output [23:0] col_out_788,
    output [23:0] col_out_789,
    output [23:0] col_out_790,
    output [23:0] col_out_791,
    output [23:0] col_out_792,
    output [23:0] col_out_793,
    output [23:0] col_out_794,
    output [23:0] col_out_795,
    output [23:0] col_out_796,
    output [23:0] col_out_797,
    output [23:0] col_out_798,
    output [23:0] col_out_799,
    output [23:0] col_out_800,
    output [23:0] col_out_801,
    output [23:0] col_out_802,
    output [23:0] col_out_803,
    output [23:0] col_out_804,
    output [23:0] col_out_805,
    output [23:0] col_out_806,
    output [23:0] col_out_807,
    output [23:0] col_out_808,
    output [23:0] col_out_809,
    output [23:0] col_out_810,
    output [23:0] col_out_811,
    output [23:0] col_out_812,
    output [23:0] col_out_813,
    output [23:0] col_out_814,
    output [23:0] col_out_815,
    output [23:0] col_out_816,
    output [23:0] col_out_817,
    output [23:0] col_out_818,
    output [23:0] col_out_819,
    output [23:0] col_out_820,
    output [23:0] col_out_821,
    output [23:0] col_out_822,
    output [23:0] col_out_823,
    output [23:0] col_out_824,
    output [23:0] col_out_825,
    output [23:0] col_out_826,
    output [23:0] col_out_827,
    output [23:0] col_out_828,
    output [23:0] col_out_829,
    output [23:0] col_out_830,
    output [23:0] col_out_831,
    output [23:0] col_out_832,
    output [23:0] col_out_833,
    output [23:0] col_out_834,
    output [23:0] col_out_835,
    output [23:0] col_out_836,
    output [23:0] col_out_837,
    output [23:0] col_out_838,
    output [23:0] col_out_839,
    output [23:0] col_out_840,
    output [23:0] col_out_841,
    output [23:0] col_out_842,
    output [23:0] col_out_843,
    output [23:0] col_out_844,
    output [23:0] col_out_845,
    output [23:0] col_out_846,
    output [23:0] col_out_847,
    output [23:0] col_out_848,
    output [23:0] col_out_849,
    output [23:0] col_out_850,
    output [23:0] col_out_851,
    output [23:0] col_out_852,
    output [23:0] col_out_853,
    output [23:0] col_out_854,
    output [23:0] col_out_855,
    output [23:0] col_out_856,
    output [23:0] col_out_857,
    output [23:0] col_out_858,
    output [23:0] col_out_859,
    output [23:0] col_out_860,
    output [23:0] col_out_861,
    output [23:0] col_out_862,
    output [23:0] col_out_863,
    output [23:0] col_out_864,
    output [23:0] col_out_865,
    output [23:0] col_out_866,
    output [23:0] col_out_867,
    output [23:0] col_out_868,
    output [23:0] col_out_869,
    output [23:0] col_out_870,
    output [23:0] col_out_871,
    output [23:0] col_out_872,
    output [23:0] col_out_873,
    output [23:0] col_out_874,
    output [23:0] col_out_875,
    output [23:0] col_out_876,
    output [23:0] col_out_877,
    output [23:0] col_out_878,
    output [23:0] col_out_879,
    output [23:0] col_out_880,
    output [23:0] col_out_881,
    output [23:0] col_out_882,
    output [23:0] col_out_883,
    output [23:0] col_out_884,
    output [23:0] col_out_885,
    output [23:0] col_out_886,
    output [23:0] col_out_887,
    output [23:0] col_out_888,
    output [23:0] col_out_889,
    output [23:0] col_out_890,
    output [23:0] col_out_891,
    output [23:0] col_out_892,
    output [23:0] col_out_893,
    output [23:0] col_out_894,
    output [23:0] col_out_895,
    output [23:0] col_out_896,
    output [23:0] col_out_897,
    output [23:0] col_out_898,
    output [23:0] col_out_899,
    output [23:0] col_out_900,
    output [23:0] col_out_901,
    output [23:0] col_out_902,
    output [23:0] col_out_903,
    output [23:0] col_out_904,
    output [23:0] col_out_905,
    output [23:0] col_out_906,
    output [23:0] col_out_907,
    output [23:0] col_out_908,
    output [23:0] col_out_909,
    output [23:0] col_out_910,
    output [23:0] col_out_911,
    output [23:0] col_out_912,
    output [23:0] col_out_913,
    output [23:0] col_out_914,
    output [23:0] col_out_915,
    output [23:0] col_out_916,
    output [23:0] col_out_917,
    output [23:0] col_out_918,
    output [23:0] col_out_919,
    output [23:0] col_out_920,
    output [23:0] col_out_921,
    output [23:0] col_out_922,
    output [23:0] col_out_923,
    output [23:0] col_out_924,
    output [23:0] col_out_925,
    output [23:0] col_out_926,
    output [23:0] col_out_927,
    output [23:0] col_out_928,
    output [23:0] col_out_929,
    output [23:0] col_out_930,
    output [23:0] col_out_931,
    output [23:0] col_out_932,
    output [23:0] col_out_933,
    output [23:0] col_out_934,
    output [23:0] col_out_935,
    output [23:0] col_out_936,
    output [23:0] col_out_937,
    output [23:0] col_out_938,
    output [23:0] col_out_939,
    output [23:0] col_out_940,
    output [23:0] col_out_941,
    output [23:0] col_out_942,
    output [23:0] col_out_943,
    output [23:0] col_out_944,
    output [23:0] col_out_945,
    output [23:0] col_out_946,
    output [23:0] col_out_947,
    output [23:0] col_out_948,
    output [23:0] col_out_949,
    output [23:0] col_out_950,
    output [23:0] col_out_951,
    output [23:0] col_out_952,
    output [23:0] col_out_953,
    output [23:0] col_out_954,
    output [23:0] col_out_955,
    output [23:0] col_out_956,
    output [23:0] col_out_957,
    output [23:0] col_out_958,
    output [23:0] col_out_959,
    output [23:0] col_out_960,
    output [23:0] col_out_961,
    output [23:0] col_out_962,
    output [23:0] col_out_963,
    output [23:0] col_out_964,
    output [23:0] col_out_965,
    output [23:0] col_out_966,
    output [23:0] col_out_967,
    output [23:0] col_out_968,
    output [23:0] col_out_969,
    output [23:0] col_out_970,
    output [23:0] col_out_971,
    output [23:0] col_out_972,
    output [23:0] col_out_973,
    output [23:0] col_out_974,
    output [23:0] col_out_975,
    output [23:0] col_out_976,
    output [23:0] col_out_977,
    output [23:0] col_out_978,
    output [23:0] col_out_979,
    output [23:0] col_out_980,
    output [23:0] col_out_981,
    output [23:0] col_out_982,
    output [23:0] col_out_983,
    output [23:0] col_out_984,
    output [23:0] col_out_985,
    output [23:0] col_out_986,
    output [23:0] col_out_987,
    output [23:0] col_out_988,
    output [23:0] col_out_989,
    output [23:0] col_out_990,
    output [23:0] col_out_991,
    output [23:0] col_out_992,
    output [23:0] col_out_993,
    output [23:0] col_out_994,
    output [23:0] col_out_995,
    output [23:0] col_out_996,
    output [23:0] col_out_997,
    output [23:0] col_out_998,
    output [23:0] col_out_999,
    output [23:0] col_out_1000,
    output [23:0] col_out_1001,
    output [23:0] col_out_1002,
    output [23:0] col_out_1003,
    output [23:0] col_out_1004,
    output [23:0] col_out_1005,
    output [23:0] col_out_1006,
    output [23:0] col_out_1007,
    output [23:0] col_out_1008,
    output [23:0] col_out_1009,
    output [23:0] col_out_1010,
    output [23:0] col_out_1011,
    output [23:0] col_out_1012,
    output [23:0] col_out_1013,
    output [23:0] col_out_1014,
    output [23:0] col_out_1015,
    output [23:0] col_out_1016,
    output [23:0] col_out_1017,
    output [23:0] col_out_1018,
    output [23:0] col_out_1019,
    output [23:0] col_out_1020,
    output [23:0] col_out_1021,
    output [23:0] col_out_1022,
    output [23:0] col_out_1023,
    output [23:0] col_out_1024,
    output [23:0] col_out_1025,
    output [23:0] col_out_1026,
    output [23:0] col_out_1027,
    output [23:0] col_out_1028,
    output [23:0] col_out_1029,
    output [23:0] col_out_1030,
    output [23:0] col_out_1031,
    output [23:0] col_out_1032,
    output [23:0] col_out_1033,
    output [23:0] col_out_1034,
    output [23:0] col_out_1035,
    output [23:0] col_out_1036,
    output [23:0] col_out_1037,
    output [23:0] col_out_1038,
    output [23:0] col_out_1039,
    output [23:0] col_out_1040,
    output [23:0] col_out_1041,
    output [23:0] col_out_1042,
    output [23:0] col_out_1043,
    output [23:0] col_out_1044,
    output [23:0] col_out_1045,
    output [23:0] col_out_1046,
    output [23:0] col_out_1047,
    output [23:0] col_out_1048,
    output [23:0] col_out_1049,
    output [23:0] col_out_1050,
    output [23:0] col_out_1051,
    output [23:0] col_out_1052,
    output [23:0] col_out_1053,
    output [23:0] col_out_1054,
    output [23:0] col_out_1055,
    output [23:0] col_out_1056,
    output [23:0] col_out_1057,
    output [23:0] col_out_1058,
    output [23:0] col_out_1059,
    output [23:0] col_out_1060,
    output [23:0] col_out_1061,
    output [23:0] col_out_1062,
    output [23:0] col_out_1063,
    output [23:0] col_out_1064,
    output [23:0] col_out_1065,
    output [23:0] col_out_1066,
    output [23:0] col_out_1067,
    output [23:0] col_out_1068,
    output [23:0] col_out_1069,
    output [23:0] col_out_1070,
    output [23:0] col_out_1071,
    output [23:0] col_out_1072,
    output [23:0] col_out_1073,
    output [23:0] col_out_1074,
    output [23:0] col_out_1075,
    output [23:0] col_out_1076,
    output [23:0] col_out_1077,
    output [23:0] col_out_1078,
    output [23:0] col_out_1079,
    output [23:0] col_out_1080,
    output [23:0] col_out_1081,
    output [23:0] col_out_1082,
    output [23:0] col_out_1083,
    output [23:0] col_out_1084,
    output [23:0] col_out_1085,
    output [23:0] col_out_1086,
    output [23:0] col_out_1087,
    output [23:0] col_out_1088,
    output [23:0] col_out_1089,
    output [23:0] col_out_1090,
    output [23:0] col_out_1091,
    output [23:0] col_out_1092,
    output [23:0] col_out_1093,
    output [23:0] col_out_1094,
    output [23:0] col_out_1095,
    output [23:0] col_out_1096,
    output [23:0] col_out_1097,
    output [23:0] col_out_1098,
    output [23:0] col_out_1099,
    output [23:0] col_out_1100,
    output [23:0] col_out_1101,
    output [23:0] col_out_1102,
    output [23:0] col_out_1103,
    output [23:0] col_out_1104,
    output [23:0] col_out_1105,
    output [23:0] col_out_1106,
    output [23:0] col_out_1107,
    output [23:0] col_out_1108,
    output [23:0] col_out_1109,
    output [23:0] col_out_1110,
    output [23:0] col_out_1111,
    output [23:0] col_out_1112,
    output [23:0] col_out_1113,
    output [23:0] col_out_1114,
    output [23:0] col_out_1115,
    output [23:0] col_out_1116,
    output [23:0] col_out_1117,
    output [23:0] col_out_1118,
    output [23:0] col_out_1119,
    output [23:0] col_out_1120,
    output [23:0] col_out_1121,
    output [23:0] col_out_1122,
    output [23:0] col_out_1123,
    output [23:0] col_out_1124,
    output [23:0] col_out_1125,
    output [23:0] col_out_1126,
    output [23:0] col_out_1127,
    output [23:0] col_out_1128,
    output [23:0] col_out_1129,
    output [23:0] col_out_1130,
    output [23:0] col_out_1131,
    output [23:0] col_out_1132,
    output [23:0] col_out_1133,
    output [23:0] col_out_1134,
    output [23:0] col_out_1135,
    output [23:0] col_out_1136,
    output [23:0] col_out_1137,
    output [23:0] col_out_1138,
    output [23:0] col_out_1139,
    output [23:0] col_out_1140,
    output [23:0] col_out_1141,
    output [23:0] col_out_1142,
    output [23:0] col_out_1143,
    output [23:0] col_out_1144,
    output [23:0] col_out_1145,
    output [23:0] col_out_1146,
    output [23:0] col_out_1147,
    output [23:0] col_out_1148,
    output [23:0] col_out_1149,
    output [23:0] col_out_1150,
    output [23:0] col_out_1151,
    output [23:0] col_out_1152,
    output [23:0] col_out_1153,
    output [23:0] col_out_1154,
    output [23:0] col_out_1155,
    output [23:0] col_out_1156,
    output [23:0] col_out_1157,
    output [23:0] col_out_1158,
    output [23:0] col_out_1159,
    output [23:0] col_out_1160,
    output [23:0] col_out_1161,
    output [23:0] col_out_1162,
    output [23:0] col_out_1163,
    output [23:0] col_out_1164,
    output [23:0] col_out_1165,
    output [23:0] col_out_1166,
    output [23:0] col_out_1167,
    output [23:0] col_out_1168,
    output [23:0] col_out_1169,
    output [23:0] col_out_1170,
    output [23:0] col_out_1171,
    output [23:0] col_out_1172,
    output [23:0] col_out_1173,
    output [23:0] col_out_1174,
    output [23:0] col_out_1175,
    output [23:0] col_out_1176,
    output [23:0] col_out_1177,
    output [23:0] col_out_1178,
    output [23:0] col_out_1179,
    output [23:0] col_out_1180,
    output [23:0] col_out_1181,
    output [23:0] col_out_1182,
    output [23:0] col_out_1183,
    output [23:0] col_out_1184,
    output [23:0] col_out_1185,
    output [23:0] col_out_1186,
    output [23:0] col_out_1187,
    output [23:0] col_out_1188,
    output [23:0] col_out_1189,
    output [23:0] col_out_1190,
    output [23:0] col_out_1191,
    output [23:0] col_out_1192,
    output [23:0] col_out_1193,
    output [23:0] col_out_1194,
    output [23:0] col_out_1195,
    output [23:0] col_out_1196,
    output [23:0] col_out_1197,
    output [23:0] col_out_1198,
    output [23:0] col_out_1199,
    output [23:0] col_out_1200,
    output [23:0] col_out_1201,
    output [23:0] col_out_1202,
    output [23:0] col_out_1203,
    output [23:0] col_out_1204,
    output [23:0] col_out_1205,
    output [23:0] col_out_1206,
    output [23:0] col_out_1207,
    output [23:0] col_out_1208,
    output [23:0] col_out_1209,
    output [23:0] col_out_1210,
    output [23:0] col_out_1211,
    output [23:0] col_out_1212,
    output [23:0] col_out_1213,
    output [23:0] col_out_1214,
    output [23:0] col_out_1215,
    output [23:0] col_out_1216,
    output [23:0] col_out_1217,
    output [23:0] col_out_1218,
    output [23:0] col_out_1219,
    output [23:0] col_out_1220,
    output [23:0] col_out_1221,
    output [23:0] col_out_1222,
    output [23:0] col_out_1223,
    output [23:0] col_out_1224,
    output [23:0] col_out_1225,
    output [23:0] col_out_1226,
    output [23:0] col_out_1227,
    output [23:0] col_out_1228,
    output [23:0] col_out_1229,
    output [23:0] col_out_1230,
    output [23:0] col_out_1231,
    output [23:0] col_out_1232,
    output [23:0] col_out_1233,
    output [23:0] col_out_1234,
    output [23:0] col_out_1235,
    output [23:0] col_out_1236,
    output [23:0] col_out_1237,
    output [23:0] col_out_1238,
    output [23:0] col_out_1239,
    output [23:0] col_out_1240,
    output [23:0] col_out_1241,
    output [23:0] col_out_1242,
    output [23:0] col_out_1243,
    output [23:0] col_out_1244,
    output [23:0] col_out_1245,
    output [23:0] col_out_1246,
    output [23:0] col_out_1247,
    output [23:0] col_out_1248,
    output [23:0] col_out_1249,
    output [23:0] col_out_1250,
    output [23:0] col_out_1251,
    output [23:0] col_out_1252,
    output [23:0] col_out_1253,
    output [23:0] col_out_1254,
    output [23:0] col_out_1255,
    output [23:0] col_out_1256,
    output [23:0] col_out_1257,
    output [23:0] col_out_1258,
    output [23:0] col_out_1259,
    output [23:0] col_out_1260,
    output [23:0] col_out_1261,
    output [23:0] col_out_1262,
    output [23:0] col_out_1263,
    output [23:0] col_out_1264,
    output [23:0] col_out_1265,
    output [23:0] col_out_1266,
    output [23:0] col_out_1267,
    output [23:0] col_out_1268,
    output [23:0] col_out_1269,
    output [23:0] col_out_1270,
    output [23:0] col_out_1271,
    output [23:0] col_out_1272,
    output [23:0] col_out_1273,
    output [23:0] col_out_1274,
    output [23:0] col_out_1275,
    output [23:0] col_out_1276,
    output [23:0] col_out_1277,
    output [23:0] col_out_1278,
    output [23:0] col_out_1279,
    output [23:0] col_out_1280,
    output [23:0] col_out_1281,
    output [23:0] col_out_1282,
    output [23:0] col_out_1283,
    output [23:0] col_out_1284,
    output [23:0] col_out_1285
);



//--compressor_array input and output----------------------

wire [80:0] u_ca_in_0;
wire [80:0] u_ca_in_1;
wire [80:0] u_ca_in_2;
wire [80:0] u_ca_in_3;
wire [80:0] u_ca_in_4;
wire [80:0] u_ca_in_5;
wire [80:0] u_ca_in_6;
wire [80:0] u_ca_in_7;
wire [80:0] u_ca_in_8;
wire [80:0] u_ca_in_9;
wire [80:0] u_ca_in_10;
wire [80:0] u_ca_in_11;
wire [80:0] u_ca_in_12;
wire [80:0] u_ca_in_13;
wire [80:0] u_ca_in_14;
wire [80:0] u_ca_in_15;
wire [80:0] u_ca_in_16;
wire [80:0] u_ca_in_17;
wire [80:0] u_ca_in_18;
wire [80:0] u_ca_in_19;
wire [80:0] u_ca_in_20;
wire [80:0] u_ca_in_21;
wire [80:0] u_ca_in_22;
wire [80:0] u_ca_in_23;
wire [80:0] u_ca_in_24;
wire [80:0] u_ca_in_25;
wire [80:0] u_ca_in_26;
wire [80:0] u_ca_in_27;
wire [80:0] u_ca_in_28;
wire [80:0] u_ca_in_29;
wire [80:0] u_ca_in_30;
wire [80:0] u_ca_in_31;
wire [80:0] u_ca_in_32;
wire [80:0] u_ca_in_33;
wire [80:0] u_ca_in_34;
wire [80:0] u_ca_in_35;
wire [80:0] u_ca_in_36;
wire [80:0] u_ca_in_37;
wire [80:0] u_ca_in_38;
wire [80:0] u_ca_in_39;
wire [80:0] u_ca_in_40;
wire [80:0] u_ca_in_41;
wire [80:0] u_ca_in_42;
wire [80:0] u_ca_in_43;
wire [80:0] u_ca_in_44;
wire [80:0] u_ca_in_45;
wire [80:0] u_ca_in_46;
wire [80:0] u_ca_in_47;
wire [80:0] u_ca_in_48;
wire [80:0] u_ca_in_49;
wire [80:0] u_ca_in_50;
wire [80:0] u_ca_in_51;
wire [80:0] u_ca_in_52;
wire [80:0] u_ca_in_53;
wire [80:0] u_ca_in_54;
wire [80:0] u_ca_in_55;
wire [80:0] u_ca_in_56;
wire [80:0] u_ca_in_57;
wire [80:0] u_ca_in_58;
wire [80:0] u_ca_in_59;
wire [80:0] u_ca_in_60;
wire [80:0] u_ca_in_61;
wire [80:0] u_ca_in_62;
wire [80:0] u_ca_in_63;
wire [80:0] u_ca_in_64;
wire [80:0] u_ca_in_65;
wire [80:0] u_ca_in_66;
wire [80:0] u_ca_in_67;
wire [80:0] u_ca_in_68;
wire [80:0] u_ca_in_69;
wire [80:0] u_ca_in_70;
wire [80:0] u_ca_in_71;
wire [80:0] u_ca_in_72;
wire [80:0] u_ca_in_73;
wire [80:0] u_ca_in_74;
wire [80:0] u_ca_in_75;
wire [80:0] u_ca_in_76;
wire [80:0] u_ca_in_77;
wire [80:0] u_ca_in_78;
wire [80:0] u_ca_in_79;
wire [80:0] u_ca_in_80;
wire [80:0] u_ca_in_81;
wire [80:0] u_ca_in_82;
wire [80:0] u_ca_in_83;
wire [80:0] u_ca_in_84;
wire [80:0] u_ca_in_85;
wire [80:0] u_ca_in_86;
wire [80:0] u_ca_in_87;
wire [80:0] u_ca_in_88;
wire [80:0] u_ca_in_89;
wire [80:0] u_ca_in_90;
wire [80:0] u_ca_in_91;
wire [80:0] u_ca_in_92;
wire [80:0] u_ca_in_93;
wire [80:0] u_ca_in_94;
wire [80:0] u_ca_in_95;
wire [80:0] u_ca_in_96;
wire [80:0] u_ca_in_97;
wire [80:0] u_ca_in_98;
wire [80:0] u_ca_in_99;
wire [80:0] u_ca_in_100;
wire [80:0] u_ca_in_101;
wire [80:0] u_ca_in_102;
wire [80:0] u_ca_in_103;
wire [80:0] u_ca_in_104;
wire [80:0] u_ca_in_105;
wire [80:0] u_ca_in_106;
wire [80:0] u_ca_in_107;
wire [80:0] u_ca_in_108;
wire [80:0] u_ca_in_109;
wire [80:0] u_ca_in_110;
wire [80:0] u_ca_in_111;
wire [80:0] u_ca_in_112;
wire [80:0] u_ca_in_113;
wire [80:0] u_ca_in_114;
wire [80:0] u_ca_in_115;
wire [80:0] u_ca_in_116;
wire [80:0] u_ca_in_117;
wire [80:0] u_ca_in_118;
wire [80:0] u_ca_in_119;
wire [80:0] u_ca_in_120;
wire [80:0] u_ca_in_121;
wire [80:0] u_ca_in_122;
wire [80:0] u_ca_in_123;
wire [80:0] u_ca_in_124;
wire [80:0] u_ca_in_125;
wire [80:0] u_ca_in_126;
wire [80:0] u_ca_in_127;
wire [80:0] u_ca_in_128;
wire [80:0] u_ca_in_129;
wire [80:0] u_ca_in_130;
wire [80:0] u_ca_in_131;
wire [80:0] u_ca_in_132;
wire [80:0] u_ca_in_133;
wire [80:0] u_ca_in_134;
wire [80:0] u_ca_in_135;
wire [80:0] u_ca_in_136;
wire [80:0] u_ca_in_137;
wire [80:0] u_ca_in_138;
wire [80:0] u_ca_in_139;
wire [80:0] u_ca_in_140;
wire [80:0] u_ca_in_141;
wire [80:0] u_ca_in_142;
wire [80:0] u_ca_in_143;
wire [80:0] u_ca_in_144;
wire [80:0] u_ca_in_145;
wire [80:0] u_ca_in_146;
wire [80:0] u_ca_in_147;
wire [80:0] u_ca_in_148;
wire [80:0] u_ca_in_149;
wire [80:0] u_ca_in_150;
wire [80:0] u_ca_in_151;
wire [80:0] u_ca_in_152;
wire [80:0] u_ca_in_153;
wire [80:0] u_ca_in_154;
wire [80:0] u_ca_in_155;
wire [80:0] u_ca_in_156;
wire [80:0] u_ca_in_157;
wire [80:0] u_ca_in_158;
wire [80:0] u_ca_in_159;
wire [80:0] u_ca_in_160;
wire [80:0] u_ca_in_161;
wire [80:0] u_ca_in_162;
wire [80:0] u_ca_in_163;
wire [80:0] u_ca_in_164;
wire [80:0] u_ca_in_165;
wire [80:0] u_ca_in_166;
wire [80:0] u_ca_in_167;
wire [80:0] u_ca_in_168;
wire [80:0] u_ca_in_169;
wire [80:0] u_ca_in_170;
wire [80:0] u_ca_in_171;
wire [80:0] u_ca_in_172;
wire [80:0] u_ca_in_173;
wire [80:0] u_ca_in_174;
wire [80:0] u_ca_in_175;
wire [80:0] u_ca_in_176;
wire [80:0] u_ca_in_177;
wire [80:0] u_ca_in_178;
wire [80:0] u_ca_in_179;
wire [80:0] u_ca_in_180;
wire [80:0] u_ca_in_181;
wire [80:0] u_ca_in_182;
wire [80:0] u_ca_in_183;
wire [80:0] u_ca_in_184;
wire [80:0] u_ca_in_185;
wire [80:0] u_ca_in_186;
wire [80:0] u_ca_in_187;
wire [80:0] u_ca_in_188;
wire [80:0] u_ca_in_189;
wire [80:0] u_ca_in_190;
wire [80:0] u_ca_in_191;
wire [80:0] u_ca_in_192;
wire [80:0] u_ca_in_193;
wire [80:0] u_ca_in_194;
wire [80:0] u_ca_in_195;
wire [80:0] u_ca_in_196;
wire [80:0] u_ca_in_197;
wire [80:0] u_ca_in_198;
wire [80:0] u_ca_in_199;
wire [80:0] u_ca_in_200;
wire [80:0] u_ca_in_201;
wire [80:0] u_ca_in_202;
wire [80:0] u_ca_in_203;
wire [80:0] u_ca_in_204;
wire [80:0] u_ca_in_205;
wire [80:0] u_ca_in_206;
wire [80:0] u_ca_in_207;
wire [80:0] u_ca_in_208;
wire [80:0] u_ca_in_209;
wire [80:0] u_ca_in_210;
wire [80:0] u_ca_in_211;
wire [80:0] u_ca_in_212;
wire [80:0] u_ca_in_213;
wire [80:0] u_ca_in_214;
wire [80:0] u_ca_in_215;
wire [80:0] u_ca_in_216;
wire [80:0] u_ca_in_217;
wire [80:0] u_ca_in_218;
wire [80:0] u_ca_in_219;
wire [80:0] u_ca_in_220;
wire [80:0] u_ca_in_221;
wire [80:0] u_ca_in_222;
wire [80:0] u_ca_in_223;
wire [80:0] u_ca_in_224;
wire [80:0] u_ca_in_225;
wire [80:0] u_ca_in_226;
wire [80:0] u_ca_in_227;
wire [80:0] u_ca_in_228;
wire [80:0] u_ca_in_229;
wire [80:0] u_ca_in_230;
wire [80:0] u_ca_in_231;
wire [80:0] u_ca_in_232;
wire [80:0] u_ca_in_233;
wire [80:0] u_ca_in_234;
wire [80:0] u_ca_in_235;
wire [80:0] u_ca_in_236;
wire [80:0] u_ca_in_237;
wire [80:0] u_ca_in_238;
wire [80:0] u_ca_in_239;
wire [80:0] u_ca_in_240;
wire [80:0] u_ca_in_241;
wire [80:0] u_ca_in_242;
wire [80:0] u_ca_in_243;
wire [80:0] u_ca_in_244;
wire [80:0] u_ca_in_245;
wire [80:0] u_ca_in_246;
wire [80:0] u_ca_in_247;
wire [80:0] u_ca_in_248;
wire [80:0] u_ca_in_249;
wire [80:0] u_ca_in_250;
wire [80:0] u_ca_in_251;
wire [80:0] u_ca_in_252;
wire [80:0] u_ca_in_253;
wire [80:0] u_ca_in_254;
wire [80:0] u_ca_in_255;
wire [80:0] u_ca_in_256;
wire [80:0] u_ca_in_257;
wire [80:0] u_ca_in_258;
wire [80:0] u_ca_in_259;
wire [80:0] u_ca_in_260;
wire [80:0] u_ca_in_261;
wire [80:0] u_ca_in_262;
wire [80:0] u_ca_in_263;
wire [80:0] u_ca_in_264;
wire [80:0] u_ca_in_265;
wire [80:0] u_ca_in_266;
wire [80:0] u_ca_in_267;
wire [80:0] u_ca_in_268;
wire [80:0] u_ca_in_269;
wire [80:0] u_ca_in_270;
wire [80:0] u_ca_in_271;
wire [80:0] u_ca_in_272;
wire [80:0] u_ca_in_273;
wire [80:0] u_ca_in_274;
wire [80:0] u_ca_in_275;
wire [80:0] u_ca_in_276;
wire [80:0] u_ca_in_277;
wire [80:0] u_ca_in_278;
wire [80:0] u_ca_in_279;
wire [80:0] u_ca_in_280;
wire [80:0] u_ca_in_281;
wire [80:0] u_ca_in_282;
wire [80:0] u_ca_in_283;
wire [80:0] u_ca_in_284;
wire [80:0] u_ca_in_285;
wire [80:0] u_ca_in_286;
wire [80:0] u_ca_in_287;
wire [80:0] u_ca_in_288;
wire [80:0] u_ca_in_289;
wire [80:0] u_ca_in_290;
wire [80:0] u_ca_in_291;
wire [80:0] u_ca_in_292;
wire [80:0] u_ca_in_293;
wire [80:0] u_ca_in_294;
wire [80:0] u_ca_in_295;
wire [80:0] u_ca_in_296;
wire [80:0] u_ca_in_297;
wire [80:0] u_ca_in_298;
wire [80:0] u_ca_in_299;
wire [80:0] u_ca_in_300;
wire [80:0] u_ca_in_301;
wire [80:0] u_ca_in_302;
wire [80:0] u_ca_in_303;
wire [80:0] u_ca_in_304;
wire [80:0] u_ca_in_305;
wire [80:0] u_ca_in_306;
wire [80:0] u_ca_in_307;
wire [80:0] u_ca_in_308;
wire [80:0] u_ca_in_309;
wire [80:0] u_ca_in_310;
wire [80:0] u_ca_in_311;
wire [80:0] u_ca_in_312;
wire [80:0] u_ca_in_313;
wire [80:0] u_ca_in_314;
wire [80:0] u_ca_in_315;
wire [80:0] u_ca_in_316;
wire [80:0] u_ca_in_317;
wire [80:0] u_ca_in_318;
wire [80:0] u_ca_in_319;
wire [80:0] u_ca_in_320;
wire [80:0] u_ca_in_321;
wire [80:0] u_ca_in_322;
wire [80:0] u_ca_in_323;
wire [80:0] u_ca_in_324;
wire [80:0] u_ca_in_325;
wire [80:0] u_ca_in_326;
wire [80:0] u_ca_in_327;
wire [80:0] u_ca_in_328;
wire [80:0] u_ca_in_329;
wire [80:0] u_ca_in_330;
wire [80:0] u_ca_in_331;
wire [80:0] u_ca_in_332;
wire [80:0] u_ca_in_333;
wire [80:0] u_ca_in_334;
wire [80:0] u_ca_in_335;
wire [80:0] u_ca_in_336;
wire [80:0] u_ca_in_337;
wire [80:0] u_ca_in_338;
wire [80:0] u_ca_in_339;
wire [80:0] u_ca_in_340;
wire [80:0] u_ca_in_341;
wire [80:0] u_ca_in_342;
wire [80:0] u_ca_in_343;
wire [80:0] u_ca_in_344;
wire [80:0] u_ca_in_345;
wire [80:0] u_ca_in_346;
wire [80:0] u_ca_in_347;
wire [80:0] u_ca_in_348;
wire [80:0] u_ca_in_349;
wire [80:0] u_ca_in_350;
wire [80:0] u_ca_in_351;
wire [80:0] u_ca_in_352;
wire [80:0] u_ca_in_353;
wire [80:0] u_ca_in_354;
wire [80:0] u_ca_in_355;
wire [80:0] u_ca_in_356;
wire [80:0] u_ca_in_357;
wire [80:0] u_ca_in_358;
wire [80:0] u_ca_in_359;
wire [80:0] u_ca_in_360;
wire [80:0] u_ca_in_361;
wire [80:0] u_ca_in_362;
wire [80:0] u_ca_in_363;
wire [80:0] u_ca_in_364;
wire [80:0] u_ca_in_365;
wire [80:0] u_ca_in_366;
wire [80:0] u_ca_in_367;
wire [80:0] u_ca_in_368;
wire [80:0] u_ca_in_369;
wire [80:0] u_ca_in_370;
wire [80:0] u_ca_in_371;
wire [80:0] u_ca_in_372;
wire [80:0] u_ca_in_373;
wire [80:0] u_ca_in_374;
wire [80:0] u_ca_in_375;
wire [80:0] u_ca_in_376;
wire [80:0] u_ca_in_377;
wire [80:0] u_ca_in_378;
wire [80:0] u_ca_in_379;
wire [80:0] u_ca_in_380;
wire [80:0] u_ca_in_381;
wire [80:0] u_ca_in_382;
wire [80:0] u_ca_in_383;
wire [80:0] u_ca_in_384;
wire [80:0] u_ca_in_385;
wire [80:0] u_ca_in_386;
wire [80:0] u_ca_in_387;
wire [80:0] u_ca_in_388;
wire [80:0] u_ca_in_389;
wire [80:0] u_ca_in_390;
wire [80:0] u_ca_in_391;
wire [80:0] u_ca_in_392;
wire [80:0] u_ca_in_393;
wire [80:0] u_ca_in_394;
wire [80:0] u_ca_in_395;
wire [80:0] u_ca_in_396;
wire [80:0] u_ca_in_397;
wire [80:0] u_ca_in_398;
wire [80:0] u_ca_in_399;
wire [80:0] u_ca_in_400;
wire [80:0] u_ca_in_401;
wire [80:0] u_ca_in_402;
wire [80:0] u_ca_in_403;
wire [80:0] u_ca_in_404;
wire [80:0] u_ca_in_405;
wire [80:0] u_ca_in_406;
wire [80:0] u_ca_in_407;
wire [80:0] u_ca_in_408;
wire [80:0] u_ca_in_409;
wire [80:0] u_ca_in_410;
wire [80:0] u_ca_in_411;
wire [80:0] u_ca_in_412;
wire [80:0] u_ca_in_413;
wire [80:0] u_ca_in_414;
wire [80:0] u_ca_in_415;
wire [80:0] u_ca_in_416;
wire [80:0] u_ca_in_417;
wire [80:0] u_ca_in_418;
wire [80:0] u_ca_in_419;
wire [80:0] u_ca_in_420;
wire [80:0] u_ca_in_421;
wire [80:0] u_ca_in_422;
wire [80:0] u_ca_in_423;
wire [80:0] u_ca_in_424;
wire [80:0] u_ca_in_425;
wire [80:0] u_ca_in_426;
wire [80:0] u_ca_in_427;
wire [80:0] u_ca_in_428;
wire [80:0] u_ca_in_429;
wire [80:0] u_ca_in_430;
wire [80:0] u_ca_in_431;
wire [80:0] u_ca_in_432;
wire [80:0] u_ca_in_433;
wire [80:0] u_ca_in_434;
wire [80:0] u_ca_in_435;
wire [80:0] u_ca_in_436;
wire [80:0] u_ca_in_437;
wire [80:0] u_ca_in_438;
wire [80:0] u_ca_in_439;
wire [80:0] u_ca_in_440;
wire [80:0] u_ca_in_441;
wire [80:0] u_ca_in_442;
wire [80:0] u_ca_in_443;
wire [80:0] u_ca_in_444;
wire [80:0] u_ca_in_445;
wire [80:0] u_ca_in_446;
wire [80:0] u_ca_in_447;
wire [80:0] u_ca_in_448;
wire [80:0] u_ca_in_449;
wire [80:0] u_ca_in_450;
wire [80:0] u_ca_in_451;
wire [80:0] u_ca_in_452;
wire [80:0] u_ca_in_453;
wire [80:0] u_ca_in_454;
wire [80:0] u_ca_in_455;
wire [80:0] u_ca_in_456;
wire [80:0] u_ca_in_457;
wire [80:0] u_ca_in_458;
wire [80:0] u_ca_in_459;
wire [80:0] u_ca_in_460;
wire [80:0] u_ca_in_461;
wire [80:0] u_ca_in_462;
wire [80:0] u_ca_in_463;
wire [80:0] u_ca_in_464;
wire [80:0] u_ca_in_465;
wire [80:0] u_ca_in_466;
wire [80:0] u_ca_in_467;
wire [80:0] u_ca_in_468;
wire [80:0] u_ca_in_469;
wire [80:0] u_ca_in_470;
wire [80:0] u_ca_in_471;
wire [80:0] u_ca_in_472;
wire [80:0] u_ca_in_473;
wire [80:0] u_ca_in_474;
wire [80:0] u_ca_in_475;
wire [80:0] u_ca_in_476;
wire [80:0] u_ca_in_477;
wire [80:0] u_ca_in_478;
wire [80:0] u_ca_in_479;
wire [80:0] u_ca_in_480;
wire [80:0] u_ca_in_481;
wire [80:0] u_ca_in_482;
wire [80:0] u_ca_in_483;
wire [80:0] u_ca_in_484;
wire [80:0] u_ca_in_485;
wire [80:0] u_ca_in_486;
wire [80:0] u_ca_in_487;
wire [80:0] u_ca_in_488;
wire [80:0] u_ca_in_489;
wire [80:0] u_ca_in_490;
wire [80:0] u_ca_in_491;
wire [80:0] u_ca_in_492;
wire [80:0] u_ca_in_493;
wire [80:0] u_ca_in_494;
wire [80:0] u_ca_in_495;
wire [80:0] u_ca_in_496;
wire [80:0] u_ca_in_497;
wire [80:0] u_ca_in_498;
wire [80:0] u_ca_in_499;
wire [80:0] u_ca_in_500;
wire [80:0] u_ca_in_501;
wire [80:0] u_ca_in_502;
wire [80:0] u_ca_in_503;
wire [80:0] u_ca_in_504;
wire [80:0] u_ca_in_505;
wire [80:0] u_ca_in_506;
wire [80:0] u_ca_in_507;
wire [80:0] u_ca_in_508;
wire [80:0] u_ca_in_509;
wire [80:0] u_ca_in_510;
wire [80:0] u_ca_in_511;
wire [80:0] u_ca_in_512;
wire [80:0] u_ca_in_513;
wire [80:0] u_ca_in_514;
wire [80:0] u_ca_in_515;
wire [80:0] u_ca_in_516;
wire [80:0] u_ca_in_517;
wire [80:0] u_ca_in_518;
wire [80:0] u_ca_in_519;
wire [80:0] u_ca_in_520;
wire [80:0] u_ca_in_521;
wire [80:0] u_ca_in_522;
wire [80:0] u_ca_in_523;
wire [80:0] u_ca_in_524;
wire [80:0] u_ca_in_525;
wire [80:0] u_ca_in_526;
wire [80:0] u_ca_in_527;
wire [80:0] u_ca_in_528;
wire [80:0] u_ca_in_529;
wire [80:0] u_ca_in_530;
wire [80:0] u_ca_in_531;
wire [80:0] u_ca_in_532;
wire [80:0] u_ca_in_533;
wire [80:0] u_ca_in_534;
wire [80:0] u_ca_in_535;
wire [80:0] u_ca_in_536;
wire [80:0] u_ca_in_537;
wire [80:0] u_ca_in_538;
wire [80:0] u_ca_in_539;
wire [80:0] u_ca_in_540;
wire [80:0] u_ca_in_541;
wire [80:0] u_ca_in_542;
wire [80:0] u_ca_in_543;
wire [80:0] u_ca_in_544;
wire [80:0] u_ca_in_545;
wire [80:0] u_ca_in_546;
wire [80:0] u_ca_in_547;
wire [80:0] u_ca_in_548;
wire [80:0] u_ca_in_549;
wire [80:0] u_ca_in_550;
wire [80:0] u_ca_in_551;
wire [80:0] u_ca_in_552;
wire [80:0] u_ca_in_553;
wire [80:0] u_ca_in_554;
wire [80:0] u_ca_in_555;
wire [80:0] u_ca_in_556;
wire [80:0] u_ca_in_557;
wire [80:0] u_ca_in_558;
wire [80:0] u_ca_in_559;
wire [80:0] u_ca_in_560;
wire [80:0] u_ca_in_561;
wire [80:0] u_ca_in_562;
wire [80:0] u_ca_in_563;
wire [80:0] u_ca_in_564;
wire [80:0] u_ca_in_565;
wire [80:0] u_ca_in_566;
wire [80:0] u_ca_in_567;
wire [80:0] u_ca_in_568;
wire [80:0] u_ca_in_569;
wire [80:0] u_ca_in_570;
wire [80:0] u_ca_in_571;
wire [80:0] u_ca_in_572;
wire [80:0] u_ca_in_573;
wire [80:0] u_ca_in_574;
wire [80:0] u_ca_in_575;
wire [80:0] u_ca_in_576;
wire [80:0] u_ca_in_577;
wire [80:0] u_ca_in_578;
wire [80:0] u_ca_in_579;
wire [80:0] u_ca_in_580;
wire [80:0] u_ca_in_581;
wire [80:0] u_ca_in_582;
wire [80:0] u_ca_in_583;
wire [80:0] u_ca_in_584;
wire [80:0] u_ca_in_585;
wire [80:0] u_ca_in_586;
wire [80:0] u_ca_in_587;
wire [80:0] u_ca_in_588;
wire [80:0] u_ca_in_589;
wire [80:0] u_ca_in_590;
wire [80:0] u_ca_in_591;
wire [80:0] u_ca_in_592;
wire [80:0] u_ca_in_593;
wire [80:0] u_ca_in_594;
wire [80:0] u_ca_in_595;
wire [80:0] u_ca_in_596;
wire [80:0] u_ca_in_597;
wire [80:0] u_ca_in_598;
wire [80:0] u_ca_in_599;
wire [80:0] u_ca_in_600;
wire [80:0] u_ca_in_601;
wire [80:0] u_ca_in_602;
wire [80:0] u_ca_in_603;
wire [80:0] u_ca_in_604;
wire [80:0] u_ca_in_605;
wire [80:0] u_ca_in_606;
wire [80:0] u_ca_in_607;
wire [80:0] u_ca_in_608;
wire [80:0] u_ca_in_609;
wire [80:0] u_ca_in_610;
wire [80:0] u_ca_in_611;
wire [80:0] u_ca_in_612;
wire [80:0] u_ca_in_613;
wire [80:0] u_ca_in_614;
wire [80:0] u_ca_in_615;
wire [80:0] u_ca_in_616;
wire [80:0] u_ca_in_617;
wire [80:0] u_ca_in_618;
wire [80:0] u_ca_in_619;
wire [80:0] u_ca_in_620;
wire [80:0] u_ca_in_621;
wire [80:0] u_ca_in_622;
wire [80:0] u_ca_in_623;
wire [80:0] u_ca_in_624;
wire [80:0] u_ca_in_625;
wire [80:0] u_ca_in_626;
wire [80:0] u_ca_in_627;
wire [80:0] u_ca_in_628;
wire [80:0] u_ca_in_629;
wire [80:0] u_ca_in_630;
wire [80:0] u_ca_in_631;
wire [80:0] u_ca_in_632;
wire [80:0] u_ca_in_633;
wire [80:0] u_ca_in_634;
wire [80:0] u_ca_in_635;
wire [80:0] u_ca_in_636;
wire [80:0] u_ca_in_637;
wire [80:0] u_ca_in_638;
wire [80:0] u_ca_in_639;
wire [80:0] u_ca_in_640;
wire [80:0] u_ca_in_641;
wire [80:0] u_ca_in_642;
wire [80:0] u_ca_in_643;
wire [80:0] u_ca_in_644;
wire [80:0] u_ca_in_645;
wire [80:0] u_ca_in_646;
wire [80:0] u_ca_in_647;
wire [80:0] u_ca_in_648;
wire [80:0] u_ca_in_649;
wire [80:0] u_ca_in_650;
wire [80:0] u_ca_in_651;
wire [80:0] u_ca_in_652;
wire [80:0] u_ca_in_653;
wire [80:0] u_ca_in_654;
wire [80:0] u_ca_in_655;
wire [80:0] u_ca_in_656;
wire [80:0] u_ca_in_657;
wire [80:0] u_ca_in_658;
wire [80:0] u_ca_in_659;
wire [80:0] u_ca_in_660;
wire [80:0] u_ca_in_661;
wire [80:0] u_ca_in_662;
wire [80:0] u_ca_in_663;
wire [80:0] u_ca_in_664;
wire [80:0] u_ca_in_665;
wire [80:0] u_ca_in_666;
wire [80:0] u_ca_in_667;
wire [80:0] u_ca_in_668;
wire [80:0] u_ca_in_669;
wire [80:0] u_ca_in_670;
wire [80:0] u_ca_in_671;
wire [80:0] u_ca_in_672;
wire [80:0] u_ca_in_673;
wire [80:0] u_ca_in_674;
wire [80:0] u_ca_in_675;
wire [80:0] u_ca_in_676;
wire [80:0] u_ca_in_677;
wire [80:0] u_ca_in_678;
wire [80:0] u_ca_in_679;
wire [80:0] u_ca_in_680;
wire [80:0] u_ca_in_681;
wire [80:0] u_ca_in_682;
wire [80:0] u_ca_in_683;
wire [80:0] u_ca_in_684;
wire [80:0] u_ca_in_685;
wire [80:0] u_ca_in_686;
wire [80:0] u_ca_in_687;
wire [80:0] u_ca_in_688;
wire [80:0] u_ca_in_689;
wire [80:0] u_ca_in_690;
wire [80:0] u_ca_in_691;
wire [80:0] u_ca_in_692;
wire [80:0] u_ca_in_693;
wire [80:0] u_ca_in_694;
wire [80:0] u_ca_in_695;
wire [80:0] u_ca_in_696;
wire [80:0] u_ca_in_697;
wire [80:0] u_ca_in_698;
wire [80:0] u_ca_in_699;
wire [80:0] u_ca_in_700;
wire [80:0] u_ca_in_701;
wire [80:0] u_ca_in_702;
wire [80:0] u_ca_in_703;
wire [80:0] u_ca_in_704;
wire [80:0] u_ca_in_705;
wire [80:0] u_ca_in_706;
wire [80:0] u_ca_in_707;
wire [80:0] u_ca_in_708;
wire [80:0] u_ca_in_709;
wire [80:0] u_ca_in_710;
wire [80:0] u_ca_in_711;
wire [80:0] u_ca_in_712;
wire [80:0] u_ca_in_713;
wire [80:0] u_ca_in_714;
wire [80:0] u_ca_in_715;
wire [80:0] u_ca_in_716;
wire [80:0] u_ca_in_717;
wire [80:0] u_ca_in_718;
wire [80:0] u_ca_in_719;
wire [80:0] u_ca_in_720;
wire [80:0] u_ca_in_721;
wire [80:0] u_ca_in_722;
wire [80:0] u_ca_in_723;
wire [80:0] u_ca_in_724;
wire [80:0] u_ca_in_725;
wire [80:0] u_ca_in_726;
wire [80:0] u_ca_in_727;
wire [80:0] u_ca_in_728;
wire [80:0] u_ca_in_729;
wire [80:0] u_ca_in_730;
wire [80:0] u_ca_in_731;
wire [80:0] u_ca_in_732;
wire [80:0] u_ca_in_733;
wire [80:0] u_ca_in_734;
wire [80:0] u_ca_in_735;
wire [80:0] u_ca_in_736;
wire [80:0] u_ca_in_737;
wire [80:0] u_ca_in_738;
wire [80:0] u_ca_in_739;
wire [80:0] u_ca_in_740;
wire [80:0] u_ca_in_741;
wire [80:0] u_ca_in_742;
wire [80:0] u_ca_in_743;
wire [80:0] u_ca_in_744;
wire [80:0] u_ca_in_745;
wire [80:0] u_ca_in_746;
wire [80:0] u_ca_in_747;
wire [80:0] u_ca_in_748;
wire [80:0] u_ca_in_749;
wire [80:0] u_ca_in_750;
wire [80:0] u_ca_in_751;
wire [80:0] u_ca_in_752;
wire [80:0] u_ca_in_753;
wire [80:0] u_ca_in_754;
wire [80:0] u_ca_in_755;
wire [80:0] u_ca_in_756;
wire [80:0] u_ca_in_757;
wire [80:0] u_ca_in_758;
wire [80:0] u_ca_in_759;
wire [80:0] u_ca_in_760;
wire [80:0] u_ca_in_761;
wire [80:0] u_ca_in_762;
wire [80:0] u_ca_in_763;
wire [80:0] u_ca_in_764;
wire [80:0] u_ca_in_765;
wire [80:0] u_ca_in_766;
wire [80:0] u_ca_in_767;
wire [80:0] u_ca_in_768;
wire [80:0] u_ca_in_769;
wire [80:0] u_ca_in_770;
wire [80:0] u_ca_in_771;
wire [80:0] u_ca_in_772;
wire [80:0] u_ca_in_773;
wire [80:0] u_ca_in_774;
wire [80:0] u_ca_in_775;
wire [80:0] u_ca_in_776;
wire [80:0] u_ca_in_777;
wire [80:0] u_ca_in_778;
wire [80:0] u_ca_in_779;
wire [80:0] u_ca_in_780;
wire [80:0] u_ca_in_781;
wire [80:0] u_ca_in_782;
wire [80:0] u_ca_in_783;
wire [80:0] u_ca_in_784;
wire [80:0] u_ca_in_785;
wire [80:0] u_ca_in_786;
wire [80:0] u_ca_in_787;
wire [80:0] u_ca_in_788;
wire [80:0] u_ca_in_789;
wire [80:0] u_ca_in_790;
wire [80:0] u_ca_in_791;
wire [80:0] u_ca_in_792;
wire [80:0] u_ca_in_793;
wire [80:0] u_ca_in_794;
wire [80:0] u_ca_in_795;
wire [80:0] u_ca_in_796;
wire [80:0] u_ca_in_797;
wire [80:0] u_ca_in_798;
wire [80:0] u_ca_in_799;
wire [80:0] u_ca_in_800;
wire [80:0] u_ca_in_801;
wire [80:0] u_ca_in_802;
wire [80:0] u_ca_in_803;
wire [80:0] u_ca_in_804;
wire [80:0] u_ca_in_805;
wire [80:0] u_ca_in_806;
wire [80:0] u_ca_in_807;
wire [80:0] u_ca_in_808;
wire [80:0] u_ca_in_809;
wire [80:0] u_ca_in_810;
wire [80:0] u_ca_in_811;
wire [80:0] u_ca_in_812;
wire [80:0] u_ca_in_813;
wire [80:0] u_ca_in_814;
wire [80:0] u_ca_in_815;
wire [80:0] u_ca_in_816;
wire [80:0] u_ca_in_817;
wire [80:0] u_ca_in_818;
wire [80:0] u_ca_in_819;
wire [80:0] u_ca_in_820;
wire [80:0] u_ca_in_821;
wire [80:0] u_ca_in_822;
wire [80:0] u_ca_in_823;
wire [80:0] u_ca_in_824;
wire [80:0] u_ca_in_825;
wire [80:0] u_ca_in_826;
wire [80:0] u_ca_in_827;
wire [80:0] u_ca_in_828;
wire [80:0] u_ca_in_829;
wire [80:0] u_ca_in_830;
wire [80:0] u_ca_in_831;
wire [80:0] u_ca_in_832;
wire [80:0] u_ca_in_833;
wire [80:0] u_ca_in_834;
wire [80:0] u_ca_in_835;
wire [80:0] u_ca_in_836;
wire [80:0] u_ca_in_837;
wire [80:0] u_ca_in_838;
wire [80:0] u_ca_in_839;
wire [80:0] u_ca_in_840;
wire [80:0] u_ca_in_841;
wire [80:0] u_ca_in_842;
wire [80:0] u_ca_in_843;
wire [80:0] u_ca_in_844;
wire [80:0] u_ca_in_845;
wire [80:0] u_ca_in_846;
wire [80:0] u_ca_in_847;
wire [80:0] u_ca_in_848;
wire [80:0] u_ca_in_849;
wire [80:0] u_ca_in_850;
wire [80:0] u_ca_in_851;
wire [80:0] u_ca_in_852;
wire [80:0] u_ca_in_853;
wire [80:0] u_ca_in_854;
wire [80:0] u_ca_in_855;
wire [80:0] u_ca_in_856;
wire [80:0] u_ca_in_857;
wire [80:0] u_ca_in_858;
wire [80:0] u_ca_in_859;
wire [80:0] u_ca_in_860;
wire [80:0] u_ca_in_861;
wire [80:0] u_ca_in_862;
wire [80:0] u_ca_in_863;
wire [80:0] u_ca_in_864;
wire [80:0] u_ca_in_865;
wire [80:0] u_ca_in_866;
wire [80:0] u_ca_in_867;
wire [80:0] u_ca_in_868;
wire [80:0] u_ca_in_869;
wire [80:0] u_ca_in_870;
wire [80:0] u_ca_in_871;
wire [80:0] u_ca_in_872;
wire [80:0] u_ca_in_873;
wire [80:0] u_ca_in_874;
wire [80:0] u_ca_in_875;
wire [80:0] u_ca_in_876;
wire [80:0] u_ca_in_877;
wire [80:0] u_ca_in_878;
wire [80:0] u_ca_in_879;
wire [80:0] u_ca_in_880;
wire [80:0] u_ca_in_881;
wire [80:0] u_ca_in_882;
wire [80:0] u_ca_in_883;
wire [80:0] u_ca_in_884;
wire [80:0] u_ca_in_885;
wire [80:0] u_ca_in_886;
wire [80:0] u_ca_in_887;
wire [80:0] u_ca_in_888;
wire [80:0] u_ca_in_889;
wire [80:0] u_ca_in_890;
wire [80:0] u_ca_in_891;
wire [80:0] u_ca_in_892;
wire [80:0] u_ca_in_893;
wire [80:0] u_ca_in_894;
wire [80:0] u_ca_in_895;
wire [80:0] u_ca_in_896;
wire [80:0] u_ca_in_897;
wire [80:0] u_ca_in_898;
wire [80:0] u_ca_in_899;
wire [80:0] u_ca_in_900;
wire [80:0] u_ca_in_901;
wire [80:0] u_ca_in_902;
wire [80:0] u_ca_in_903;
wire [80:0] u_ca_in_904;
wire [80:0] u_ca_in_905;
wire [80:0] u_ca_in_906;
wire [80:0] u_ca_in_907;
wire [80:0] u_ca_in_908;
wire [80:0] u_ca_in_909;
wire [80:0] u_ca_in_910;
wire [80:0] u_ca_in_911;
wire [80:0] u_ca_in_912;
wire [80:0] u_ca_in_913;
wire [80:0] u_ca_in_914;
wire [80:0] u_ca_in_915;
wire [80:0] u_ca_in_916;
wire [80:0] u_ca_in_917;
wire [80:0] u_ca_in_918;
wire [80:0] u_ca_in_919;
wire [80:0] u_ca_in_920;
wire [80:0] u_ca_in_921;
wire [80:0] u_ca_in_922;
wire [80:0] u_ca_in_923;
wire [80:0] u_ca_in_924;
wire [80:0] u_ca_in_925;
wire [80:0] u_ca_in_926;
wire [80:0] u_ca_in_927;
wire [80:0] u_ca_in_928;
wire [80:0] u_ca_in_929;
wire [80:0] u_ca_in_930;
wire [80:0] u_ca_in_931;
wire [80:0] u_ca_in_932;
wire [80:0] u_ca_in_933;
wire [80:0] u_ca_in_934;
wire [80:0] u_ca_in_935;
wire [80:0] u_ca_in_936;
wire [80:0] u_ca_in_937;
wire [80:0] u_ca_in_938;
wire [80:0] u_ca_in_939;
wire [80:0] u_ca_in_940;
wire [80:0] u_ca_in_941;
wire [80:0] u_ca_in_942;
wire [80:0] u_ca_in_943;
wire [80:0] u_ca_in_944;
wire [80:0] u_ca_in_945;
wire [80:0] u_ca_in_946;
wire [80:0] u_ca_in_947;
wire [80:0] u_ca_in_948;
wire [80:0] u_ca_in_949;
wire [80:0] u_ca_in_950;
wire [80:0] u_ca_in_951;
wire [80:0] u_ca_in_952;
wire [80:0] u_ca_in_953;
wire [80:0] u_ca_in_954;
wire [80:0] u_ca_in_955;
wire [80:0] u_ca_in_956;
wire [80:0] u_ca_in_957;
wire [80:0] u_ca_in_958;
wire [80:0] u_ca_in_959;
wire [80:0] u_ca_in_960;
wire [80:0] u_ca_in_961;
wire [80:0] u_ca_in_962;
wire [80:0] u_ca_in_963;
wire [80:0] u_ca_in_964;
wire [80:0] u_ca_in_965;
wire [80:0] u_ca_in_966;
wire [80:0] u_ca_in_967;
wire [80:0] u_ca_in_968;
wire [80:0] u_ca_in_969;
wire [80:0] u_ca_in_970;
wire [80:0] u_ca_in_971;
wire [80:0] u_ca_in_972;
wire [80:0] u_ca_in_973;
wire [80:0] u_ca_in_974;
wire [80:0] u_ca_in_975;
wire [80:0] u_ca_in_976;
wire [80:0] u_ca_in_977;
wire [80:0] u_ca_in_978;
wire [80:0] u_ca_in_979;
wire [80:0] u_ca_in_980;
wire [80:0] u_ca_in_981;
wire [80:0] u_ca_in_982;
wire [80:0] u_ca_in_983;
wire [80:0] u_ca_in_984;
wire [80:0] u_ca_in_985;
wire [80:0] u_ca_in_986;
wire [80:0] u_ca_in_987;
wire [80:0] u_ca_in_988;
wire [80:0] u_ca_in_989;
wire [80:0] u_ca_in_990;
wire [80:0] u_ca_in_991;
wire [80:0] u_ca_in_992;
wire [80:0] u_ca_in_993;
wire [80:0] u_ca_in_994;
wire [80:0] u_ca_in_995;
wire [80:0] u_ca_in_996;
wire [80:0] u_ca_in_997;
wire [80:0] u_ca_in_998;
wire [80:0] u_ca_in_999;
wire [80:0] u_ca_in_1000;
wire [80:0] u_ca_in_1001;
wire [80:0] u_ca_in_1002;
wire [80:0] u_ca_in_1003;
wire [80:0] u_ca_in_1004;
wire [80:0] u_ca_in_1005;
wire [80:0] u_ca_in_1006;
wire [80:0] u_ca_in_1007;
wire [80:0] u_ca_in_1008;
wire [80:0] u_ca_in_1009;
wire [80:0] u_ca_in_1010;
wire [80:0] u_ca_in_1011;
wire [80:0] u_ca_in_1012;
wire [80:0] u_ca_in_1013;
wire [80:0] u_ca_in_1014;
wire [80:0] u_ca_in_1015;
wire [80:0] u_ca_in_1016;
wire [80:0] u_ca_in_1017;
wire [80:0] u_ca_in_1018;
wire [80:0] u_ca_in_1019;
wire [80:0] u_ca_in_1020;
wire [80:0] u_ca_in_1021;
wire [80:0] u_ca_in_1022;
wire [80:0] u_ca_in_1023;
wire [80:0] u_ca_in_1024;
wire [80:0] u_ca_in_1025;
wire [80:0] u_ca_in_1026;
wire [80:0] u_ca_in_1027;
wire [80:0] u_ca_in_1028;
wire [80:0] u_ca_in_1029;
wire [80:0] u_ca_in_1030;
wire [80:0] u_ca_in_1031;
wire [80:0] u_ca_in_1032;
wire [80:0] u_ca_in_1033;
wire [80:0] u_ca_in_1034;
wire [80:0] u_ca_in_1035;
wire [80:0] u_ca_in_1036;
wire [80:0] u_ca_in_1037;
wire [80:0] u_ca_in_1038;
wire [80:0] u_ca_in_1039;
wire [80:0] u_ca_in_1040;
wire [80:0] u_ca_in_1041;
wire [80:0] u_ca_in_1042;
wire [80:0] u_ca_in_1043;
wire [80:0] u_ca_in_1044;
wire [80:0] u_ca_in_1045;
wire [80:0] u_ca_in_1046;
wire [80:0] u_ca_in_1047;
wire [80:0] u_ca_in_1048;
wire [80:0] u_ca_in_1049;
wire [80:0] u_ca_in_1050;
wire [80:0] u_ca_in_1051;
wire [80:0] u_ca_in_1052;
wire [80:0] u_ca_in_1053;
wire [80:0] u_ca_in_1054;
wire [80:0] u_ca_in_1055;
wire [80:0] u_ca_in_1056;
wire [80:0] u_ca_in_1057;
wire [80:0] u_ca_in_1058;
wire [80:0] u_ca_in_1059;
wire [80:0] u_ca_in_1060;
wire [80:0] u_ca_in_1061;
wire [80:0] u_ca_in_1062;
wire [80:0] u_ca_in_1063;
wire [80:0] u_ca_in_1064;
wire [80:0] u_ca_in_1065;
wire [80:0] u_ca_in_1066;
wire [80:0] u_ca_in_1067;
wire [80:0] u_ca_in_1068;
wire [80:0] u_ca_in_1069;
wire [80:0] u_ca_in_1070;
wire [80:0] u_ca_in_1071;
wire [80:0] u_ca_in_1072;
wire [80:0] u_ca_in_1073;
wire [80:0] u_ca_in_1074;
wire [80:0] u_ca_in_1075;
wire [80:0] u_ca_in_1076;
wire [80:0] u_ca_in_1077;
wire [80:0] u_ca_in_1078;
wire [80:0] u_ca_in_1079;
wire [80:0] u_ca_in_1080;
wire [80:0] u_ca_in_1081;
wire [80:0] u_ca_in_1082;
wire [80:0] u_ca_in_1083;
wire [80:0] u_ca_in_1084;
wire [80:0] u_ca_in_1085;
wire [80:0] u_ca_in_1086;
wire [80:0] u_ca_in_1087;
wire [80:0] u_ca_in_1088;
wire [80:0] u_ca_in_1089;
wire [80:0] u_ca_in_1090;
wire [80:0] u_ca_in_1091;
wire [80:0] u_ca_in_1092;
wire [80:0] u_ca_in_1093;
wire [80:0] u_ca_in_1094;
wire [80:0] u_ca_in_1095;
wire [80:0] u_ca_in_1096;
wire [80:0] u_ca_in_1097;
wire [80:0] u_ca_in_1098;
wire [80:0] u_ca_in_1099;
wire [80:0] u_ca_in_1100;
wire [80:0] u_ca_in_1101;
wire [80:0] u_ca_in_1102;
wire [80:0] u_ca_in_1103;
wire [80:0] u_ca_in_1104;
wire [80:0] u_ca_in_1105;
wire [80:0] u_ca_in_1106;
wire [80:0] u_ca_in_1107;
wire [80:0] u_ca_in_1108;
wire [80:0] u_ca_in_1109;
wire [80:0] u_ca_in_1110;
wire [80:0] u_ca_in_1111;
wire [80:0] u_ca_in_1112;
wire [80:0] u_ca_in_1113;
wire [80:0] u_ca_in_1114;
wire [80:0] u_ca_in_1115;
wire [80:0] u_ca_in_1116;
wire [80:0] u_ca_in_1117;
wire [80:0] u_ca_in_1118;
wire [80:0] u_ca_in_1119;
wire [80:0] u_ca_in_1120;
wire [80:0] u_ca_in_1121;
wire [80:0] u_ca_in_1122;
wire [80:0] u_ca_in_1123;
wire [80:0] u_ca_in_1124;
wire [80:0] u_ca_in_1125;
wire [80:0] u_ca_in_1126;
wire [80:0] u_ca_in_1127;
wire [80:0] u_ca_in_1128;
wire [80:0] u_ca_in_1129;
wire [80:0] u_ca_in_1130;
wire [80:0] u_ca_in_1131;
wire [80:0] u_ca_in_1132;
wire [80:0] u_ca_in_1133;
wire [80:0] u_ca_in_1134;
wire [80:0] u_ca_in_1135;
wire [80:0] u_ca_in_1136;
wire [80:0] u_ca_in_1137;
wire [80:0] u_ca_in_1138;
wire [80:0] u_ca_in_1139;
wire [80:0] u_ca_in_1140;
wire [80:0] u_ca_in_1141;
wire [80:0] u_ca_in_1142;
wire [80:0] u_ca_in_1143;
wire [80:0] u_ca_in_1144;
wire [80:0] u_ca_in_1145;
wire [80:0] u_ca_in_1146;
wire [80:0] u_ca_in_1147;
wire [80:0] u_ca_in_1148;
wire [80:0] u_ca_in_1149;
wire [80:0] u_ca_in_1150;
wire [80:0] u_ca_in_1151;
wire [80:0] u_ca_in_1152;
wire [80:0] u_ca_in_1153;
wire [80:0] u_ca_in_1154;
wire [80:0] u_ca_in_1155;
wire [80:0] u_ca_in_1156;
wire [80:0] u_ca_in_1157;
wire [80:0] u_ca_in_1158;
wire [80:0] u_ca_in_1159;
wire [80:0] u_ca_in_1160;
wire [80:0] u_ca_in_1161;
wire [80:0] u_ca_in_1162;
wire [80:0] u_ca_in_1163;
wire [80:0] u_ca_in_1164;
wire [80:0] u_ca_in_1165;
wire [80:0] u_ca_in_1166;
wire [80:0] u_ca_in_1167;
wire [80:0] u_ca_in_1168;
wire [80:0] u_ca_in_1169;
wire [80:0] u_ca_in_1170;
wire [80:0] u_ca_in_1171;
wire [80:0] u_ca_in_1172;
wire [80:0] u_ca_in_1173;
wire [80:0] u_ca_in_1174;
wire [80:0] u_ca_in_1175;
wire [80:0] u_ca_in_1176;
wire [80:0] u_ca_in_1177;
wire [80:0] u_ca_in_1178;
wire [80:0] u_ca_in_1179;
wire [80:0] u_ca_in_1180;
wire [80:0] u_ca_in_1181;
wire [80:0] u_ca_in_1182;
wire [80:0] u_ca_in_1183;
wire [80:0] u_ca_in_1184;
wire [80:0] u_ca_in_1185;
wire [80:0] u_ca_in_1186;
wire [80:0] u_ca_in_1187;
wire [80:0] u_ca_in_1188;
wire [80:0] u_ca_in_1189;
wire [80:0] u_ca_in_1190;
wire [80:0] u_ca_in_1191;
wire [80:0] u_ca_in_1192;
wire [80:0] u_ca_in_1193;
wire [80:0] u_ca_in_1194;
wire [80:0] u_ca_in_1195;
wire [80:0] u_ca_in_1196;
wire [80:0] u_ca_in_1197;
wire [80:0] u_ca_in_1198;
wire [80:0] u_ca_in_1199;
wire [80:0] u_ca_in_1200;
wire [80:0] u_ca_in_1201;
wire [80:0] u_ca_in_1202;
wire [80:0] u_ca_in_1203;
wire [80:0] u_ca_in_1204;
wire [80:0] u_ca_in_1205;
wire [80:0] u_ca_in_1206;
wire [80:0] u_ca_in_1207;
wire [80:0] u_ca_in_1208;
wire [80:0] u_ca_in_1209;
wire [80:0] u_ca_in_1210;
wire [80:0] u_ca_in_1211;
wire [80:0] u_ca_in_1212;
wire [80:0] u_ca_in_1213;
wire [80:0] u_ca_in_1214;
wire [80:0] u_ca_in_1215;
wire [80:0] u_ca_in_1216;
wire [80:0] u_ca_in_1217;
wire [80:0] u_ca_in_1218;
wire [80:0] u_ca_in_1219;
wire [80:0] u_ca_in_1220;
wire [80:0] u_ca_in_1221;
wire [80:0] u_ca_in_1222;
wire [80:0] u_ca_in_1223;
wire [80:0] u_ca_in_1224;
wire [80:0] u_ca_in_1225;
wire [80:0] u_ca_in_1226;
wire [80:0] u_ca_in_1227;
wire [80:0] u_ca_in_1228;
wire [80:0] u_ca_in_1229;
wire [80:0] u_ca_in_1230;
wire [80:0] u_ca_in_1231;
wire [80:0] u_ca_in_1232;
wire [80:0] u_ca_in_1233;
wire [80:0] u_ca_in_1234;
wire [80:0] u_ca_in_1235;
wire [80:0] u_ca_in_1236;
wire [80:0] u_ca_in_1237;
wire [80:0] u_ca_in_1238;
wire [80:0] u_ca_in_1239;
wire [80:0] u_ca_in_1240;
wire [80:0] u_ca_in_1241;
wire [80:0] u_ca_in_1242;
wire [80:0] u_ca_in_1243;
wire [80:0] u_ca_in_1244;
wire [80:0] u_ca_in_1245;
wire [80:0] u_ca_in_1246;
wire [80:0] u_ca_in_1247;
wire [80:0] u_ca_in_1248;
wire [80:0] u_ca_in_1249;
wire [80:0] u_ca_in_1250;
wire [80:0] u_ca_in_1251;
wire [80:0] u_ca_in_1252;
wire [80:0] u_ca_in_1253;
wire [80:0] u_ca_in_1254;
wire [80:0] u_ca_in_1255;
wire [80:0] u_ca_in_1256;
wire [80:0] u_ca_in_1257;
wire [80:0] u_ca_in_1258;
wire [80:0] u_ca_in_1259;
wire [80:0] u_ca_in_1260;
wire [80:0] u_ca_in_1261;
wire [80:0] u_ca_in_1262;
wire [80:0] u_ca_in_1263;
wire [80:0] u_ca_in_1264;
wire [80:0] u_ca_in_1265;
wire [80:0] u_ca_in_1266;
wire [80:0] u_ca_in_1267;
wire [80:0] u_ca_in_1268;
wire [80:0] u_ca_in_1269;
wire [80:0] u_ca_in_1270;
wire [80:0] u_ca_in_1271;
wire [80:0] u_ca_in_1272;
wire [80:0] u_ca_in_1273;
wire [80:0] u_ca_in_1274;
wire [80:0] u_ca_in_1275;
wire [80:0] u_ca_in_1276;
wire [80:0] u_ca_in_1277;
wire [80:0] u_ca_in_1278;
wire [80:0] u_ca_in_1279;
wire [80:0] u_ca_in_1280;
wire [80:0] u_ca_in_1281;
wire [80:0] u_ca_in_1282;


wire [23:0] u_ca_out_0;
wire [23:0] u_ca_out_1;
wire [23:0] u_ca_out_2;
wire [23:0] u_ca_out_3;
wire [23:0] u_ca_out_4;
wire [23:0] u_ca_out_5;
wire [23:0] u_ca_out_6;
wire [23:0] u_ca_out_7;
wire [23:0] u_ca_out_8;
wire [23:0] u_ca_out_9;
wire [23:0] u_ca_out_10;
wire [23:0] u_ca_out_11;
wire [23:0] u_ca_out_12;
wire [23:0] u_ca_out_13;
wire [23:0] u_ca_out_14;
wire [23:0] u_ca_out_15;
wire [23:0] u_ca_out_16;
wire [23:0] u_ca_out_17;
wire [23:0] u_ca_out_18;
wire [23:0] u_ca_out_19;
wire [23:0] u_ca_out_20;
wire [23:0] u_ca_out_21;
wire [23:0] u_ca_out_22;
wire [23:0] u_ca_out_23;
wire [23:0] u_ca_out_24;
wire [23:0] u_ca_out_25;
wire [23:0] u_ca_out_26;
wire [23:0] u_ca_out_27;
wire [23:0] u_ca_out_28;
wire [23:0] u_ca_out_29;
wire [23:0] u_ca_out_30;
wire [23:0] u_ca_out_31;
wire [23:0] u_ca_out_32;
wire [23:0] u_ca_out_33;
wire [23:0] u_ca_out_34;
wire [23:0] u_ca_out_35;
wire [23:0] u_ca_out_36;
wire [23:0] u_ca_out_37;
wire [23:0] u_ca_out_38;
wire [23:0] u_ca_out_39;
wire [23:0] u_ca_out_40;
wire [23:0] u_ca_out_41;
wire [23:0] u_ca_out_42;
wire [23:0] u_ca_out_43;
wire [23:0] u_ca_out_44;
wire [23:0] u_ca_out_45;
wire [23:0] u_ca_out_46;
wire [23:0] u_ca_out_47;
wire [23:0] u_ca_out_48;
wire [23:0] u_ca_out_49;
wire [23:0] u_ca_out_50;
wire [23:0] u_ca_out_51;
wire [23:0] u_ca_out_52;
wire [23:0] u_ca_out_53;
wire [23:0] u_ca_out_54;
wire [23:0] u_ca_out_55;
wire [23:0] u_ca_out_56;
wire [23:0] u_ca_out_57;
wire [23:0] u_ca_out_58;
wire [23:0] u_ca_out_59;
wire [23:0] u_ca_out_60;
wire [23:0] u_ca_out_61;
wire [23:0] u_ca_out_62;
wire [23:0] u_ca_out_63;
wire [23:0] u_ca_out_64;
wire [23:0] u_ca_out_65;
wire [23:0] u_ca_out_66;
wire [23:0] u_ca_out_67;
wire [23:0] u_ca_out_68;
wire [23:0] u_ca_out_69;
wire [23:0] u_ca_out_70;
wire [23:0] u_ca_out_71;
wire [23:0] u_ca_out_72;
wire [23:0] u_ca_out_73;
wire [23:0] u_ca_out_74;
wire [23:0] u_ca_out_75;
wire [23:0] u_ca_out_76;
wire [23:0] u_ca_out_77;
wire [23:0] u_ca_out_78;
wire [23:0] u_ca_out_79;
wire [23:0] u_ca_out_80;
wire [23:0] u_ca_out_81;
wire [23:0] u_ca_out_82;
wire [23:0] u_ca_out_83;
wire [23:0] u_ca_out_84;
wire [23:0] u_ca_out_85;
wire [23:0] u_ca_out_86;
wire [23:0] u_ca_out_87;
wire [23:0] u_ca_out_88;
wire [23:0] u_ca_out_89;
wire [23:0] u_ca_out_90;
wire [23:0] u_ca_out_91;
wire [23:0] u_ca_out_92;
wire [23:0] u_ca_out_93;
wire [23:0] u_ca_out_94;
wire [23:0] u_ca_out_95;
wire [23:0] u_ca_out_96;
wire [23:0] u_ca_out_97;
wire [23:0] u_ca_out_98;
wire [23:0] u_ca_out_99;
wire [23:0] u_ca_out_100;
wire [23:0] u_ca_out_101;
wire [23:0] u_ca_out_102;
wire [23:0] u_ca_out_103;
wire [23:0] u_ca_out_104;
wire [23:0] u_ca_out_105;
wire [23:0] u_ca_out_106;
wire [23:0] u_ca_out_107;
wire [23:0] u_ca_out_108;
wire [23:0] u_ca_out_109;
wire [23:0] u_ca_out_110;
wire [23:0] u_ca_out_111;
wire [23:0] u_ca_out_112;
wire [23:0] u_ca_out_113;
wire [23:0] u_ca_out_114;
wire [23:0] u_ca_out_115;
wire [23:0] u_ca_out_116;
wire [23:0] u_ca_out_117;
wire [23:0] u_ca_out_118;
wire [23:0] u_ca_out_119;
wire [23:0] u_ca_out_120;
wire [23:0] u_ca_out_121;
wire [23:0] u_ca_out_122;
wire [23:0] u_ca_out_123;
wire [23:0] u_ca_out_124;
wire [23:0] u_ca_out_125;
wire [23:0] u_ca_out_126;
wire [23:0] u_ca_out_127;
wire [23:0] u_ca_out_128;
wire [23:0] u_ca_out_129;
wire [23:0] u_ca_out_130;
wire [23:0] u_ca_out_131;
wire [23:0] u_ca_out_132;
wire [23:0] u_ca_out_133;
wire [23:0] u_ca_out_134;
wire [23:0] u_ca_out_135;
wire [23:0] u_ca_out_136;
wire [23:0] u_ca_out_137;
wire [23:0] u_ca_out_138;
wire [23:0] u_ca_out_139;
wire [23:0] u_ca_out_140;
wire [23:0] u_ca_out_141;
wire [23:0] u_ca_out_142;
wire [23:0] u_ca_out_143;
wire [23:0] u_ca_out_144;
wire [23:0] u_ca_out_145;
wire [23:0] u_ca_out_146;
wire [23:0] u_ca_out_147;
wire [23:0] u_ca_out_148;
wire [23:0] u_ca_out_149;
wire [23:0] u_ca_out_150;
wire [23:0] u_ca_out_151;
wire [23:0] u_ca_out_152;
wire [23:0] u_ca_out_153;
wire [23:0] u_ca_out_154;
wire [23:0] u_ca_out_155;
wire [23:0] u_ca_out_156;
wire [23:0] u_ca_out_157;
wire [23:0] u_ca_out_158;
wire [23:0] u_ca_out_159;
wire [23:0] u_ca_out_160;
wire [23:0] u_ca_out_161;
wire [23:0] u_ca_out_162;
wire [23:0] u_ca_out_163;
wire [23:0] u_ca_out_164;
wire [23:0] u_ca_out_165;
wire [23:0] u_ca_out_166;
wire [23:0] u_ca_out_167;
wire [23:0] u_ca_out_168;
wire [23:0] u_ca_out_169;
wire [23:0] u_ca_out_170;
wire [23:0] u_ca_out_171;
wire [23:0] u_ca_out_172;
wire [23:0] u_ca_out_173;
wire [23:0] u_ca_out_174;
wire [23:0] u_ca_out_175;
wire [23:0] u_ca_out_176;
wire [23:0] u_ca_out_177;
wire [23:0] u_ca_out_178;
wire [23:0] u_ca_out_179;
wire [23:0] u_ca_out_180;
wire [23:0] u_ca_out_181;
wire [23:0] u_ca_out_182;
wire [23:0] u_ca_out_183;
wire [23:0] u_ca_out_184;
wire [23:0] u_ca_out_185;
wire [23:0] u_ca_out_186;
wire [23:0] u_ca_out_187;
wire [23:0] u_ca_out_188;
wire [23:0] u_ca_out_189;
wire [23:0] u_ca_out_190;
wire [23:0] u_ca_out_191;
wire [23:0] u_ca_out_192;
wire [23:0] u_ca_out_193;
wire [23:0] u_ca_out_194;
wire [23:0] u_ca_out_195;
wire [23:0] u_ca_out_196;
wire [23:0] u_ca_out_197;
wire [23:0] u_ca_out_198;
wire [23:0] u_ca_out_199;
wire [23:0] u_ca_out_200;
wire [23:0] u_ca_out_201;
wire [23:0] u_ca_out_202;
wire [23:0] u_ca_out_203;
wire [23:0] u_ca_out_204;
wire [23:0] u_ca_out_205;
wire [23:0] u_ca_out_206;
wire [23:0] u_ca_out_207;
wire [23:0] u_ca_out_208;
wire [23:0] u_ca_out_209;
wire [23:0] u_ca_out_210;
wire [23:0] u_ca_out_211;
wire [23:0] u_ca_out_212;
wire [23:0] u_ca_out_213;
wire [23:0] u_ca_out_214;
wire [23:0] u_ca_out_215;
wire [23:0] u_ca_out_216;
wire [23:0] u_ca_out_217;
wire [23:0] u_ca_out_218;
wire [23:0] u_ca_out_219;
wire [23:0] u_ca_out_220;
wire [23:0] u_ca_out_221;
wire [23:0] u_ca_out_222;
wire [23:0] u_ca_out_223;
wire [23:0] u_ca_out_224;
wire [23:0] u_ca_out_225;
wire [23:0] u_ca_out_226;
wire [23:0] u_ca_out_227;
wire [23:0] u_ca_out_228;
wire [23:0] u_ca_out_229;
wire [23:0] u_ca_out_230;
wire [23:0] u_ca_out_231;
wire [23:0] u_ca_out_232;
wire [23:0] u_ca_out_233;
wire [23:0] u_ca_out_234;
wire [23:0] u_ca_out_235;
wire [23:0] u_ca_out_236;
wire [23:0] u_ca_out_237;
wire [23:0] u_ca_out_238;
wire [23:0] u_ca_out_239;
wire [23:0] u_ca_out_240;
wire [23:0] u_ca_out_241;
wire [23:0] u_ca_out_242;
wire [23:0] u_ca_out_243;
wire [23:0] u_ca_out_244;
wire [23:0] u_ca_out_245;
wire [23:0] u_ca_out_246;
wire [23:0] u_ca_out_247;
wire [23:0] u_ca_out_248;
wire [23:0] u_ca_out_249;
wire [23:0] u_ca_out_250;
wire [23:0] u_ca_out_251;
wire [23:0] u_ca_out_252;
wire [23:0] u_ca_out_253;
wire [23:0] u_ca_out_254;
wire [23:0] u_ca_out_255;
wire [23:0] u_ca_out_256;
wire [23:0] u_ca_out_257;
wire [23:0] u_ca_out_258;
wire [23:0] u_ca_out_259;
wire [23:0] u_ca_out_260;
wire [23:0] u_ca_out_261;
wire [23:0] u_ca_out_262;
wire [23:0] u_ca_out_263;
wire [23:0] u_ca_out_264;
wire [23:0] u_ca_out_265;
wire [23:0] u_ca_out_266;
wire [23:0] u_ca_out_267;
wire [23:0] u_ca_out_268;
wire [23:0] u_ca_out_269;
wire [23:0] u_ca_out_270;
wire [23:0] u_ca_out_271;
wire [23:0] u_ca_out_272;
wire [23:0] u_ca_out_273;
wire [23:0] u_ca_out_274;
wire [23:0] u_ca_out_275;
wire [23:0] u_ca_out_276;
wire [23:0] u_ca_out_277;
wire [23:0] u_ca_out_278;
wire [23:0] u_ca_out_279;
wire [23:0] u_ca_out_280;
wire [23:0] u_ca_out_281;
wire [23:0] u_ca_out_282;
wire [23:0] u_ca_out_283;
wire [23:0] u_ca_out_284;
wire [23:0] u_ca_out_285;
wire [23:0] u_ca_out_286;
wire [23:0] u_ca_out_287;
wire [23:0] u_ca_out_288;
wire [23:0] u_ca_out_289;
wire [23:0] u_ca_out_290;
wire [23:0] u_ca_out_291;
wire [23:0] u_ca_out_292;
wire [23:0] u_ca_out_293;
wire [23:0] u_ca_out_294;
wire [23:0] u_ca_out_295;
wire [23:0] u_ca_out_296;
wire [23:0] u_ca_out_297;
wire [23:0] u_ca_out_298;
wire [23:0] u_ca_out_299;
wire [23:0] u_ca_out_300;
wire [23:0] u_ca_out_301;
wire [23:0] u_ca_out_302;
wire [23:0] u_ca_out_303;
wire [23:0] u_ca_out_304;
wire [23:0] u_ca_out_305;
wire [23:0] u_ca_out_306;
wire [23:0] u_ca_out_307;
wire [23:0] u_ca_out_308;
wire [23:0] u_ca_out_309;
wire [23:0] u_ca_out_310;
wire [23:0] u_ca_out_311;
wire [23:0] u_ca_out_312;
wire [23:0] u_ca_out_313;
wire [23:0] u_ca_out_314;
wire [23:0] u_ca_out_315;
wire [23:0] u_ca_out_316;
wire [23:0] u_ca_out_317;
wire [23:0] u_ca_out_318;
wire [23:0] u_ca_out_319;
wire [23:0] u_ca_out_320;
wire [23:0] u_ca_out_321;
wire [23:0] u_ca_out_322;
wire [23:0] u_ca_out_323;
wire [23:0] u_ca_out_324;
wire [23:0] u_ca_out_325;
wire [23:0] u_ca_out_326;
wire [23:0] u_ca_out_327;
wire [23:0] u_ca_out_328;
wire [23:0] u_ca_out_329;
wire [23:0] u_ca_out_330;
wire [23:0] u_ca_out_331;
wire [23:0] u_ca_out_332;
wire [23:0] u_ca_out_333;
wire [23:0] u_ca_out_334;
wire [23:0] u_ca_out_335;
wire [23:0] u_ca_out_336;
wire [23:0] u_ca_out_337;
wire [23:0] u_ca_out_338;
wire [23:0] u_ca_out_339;
wire [23:0] u_ca_out_340;
wire [23:0] u_ca_out_341;
wire [23:0] u_ca_out_342;
wire [23:0] u_ca_out_343;
wire [23:0] u_ca_out_344;
wire [23:0] u_ca_out_345;
wire [23:0] u_ca_out_346;
wire [23:0] u_ca_out_347;
wire [23:0] u_ca_out_348;
wire [23:0] u_ca_out_349;
wire [23:0] u_ca_out_350;
wire [23:0] u_ca_out_351;
wire [23:0] u_ca_out_352;
wire [23:0] u_ca_out_353;
wire [23:0] u_ca_out_354;
wire [23:0] u_ca_out_355;
wire [23:0] u_ca_out_356;
wire [23:0] u_ca_out_357;
wire [23:0] u_ca_out_358;
wire [23:0] u_ca_out_359;
wire [23:0] u_ca_out_360;
wire [23:0] u_ca_out_361;
wire [23:0] u_ca_out_362;
wire [23:0] u_ca_out_363;
wire [23:0] u_ca_out_364;
wire [23:0] u_ca_out_365;
wire [23:0] u_ca_out_366;
wire [23:0] u_ca_out_367;
wire [23:0] u_ca_out_368;
wire [23:0] u_ca_out_369;
wire [23:0] u_ca_out_370;
wire [23:0] u_ca_out_371;
wire [23:0] u_ca_out_372;
wire [23:0] u_ca_out_373;
wire [23:0] u_ca_out_374;
wire [23:0] u_ca_out_375;
wire [23:0] u_ca_out_376;
wire [23:0] u_ca_out_377;
wire [23:0] u_ca_out_378;
wire [23:0] u_ca_out_379;
wire [23:0] u_ca_out_380;
wire [23:0] u_ca_out_381;
wire [23:0] u_ca_out_382;
wire [23:0] u_ca_out_383;
wire [23:0] u_ca_out_384;
wire [23:0] u_ca_out_385;
wire [23:0] u_ca_out_386;
wire [23:0] u_ca_out_387;
wire [23:0] u_ca_out_388;
wire [23:0] u_ca_out_389;
wire [23:0] u_ca_out_390;
wire [23:0] u_ca_out_391;
wire [23:0] u_ca_out_392;
wire [23:0] u_ca_out_393;
wire [23:0] u_ca_out_394;
wire [23:0] u_ca_out_395;
wire [23:0] u_ca_out_396;
wire [23:0] u_ca_out_397;
wire [23:0] u_ca_out_398;
wire [23:0] u_ca_out_399;
wire [23:0] u_ca_out_400;
wire [23:0] u_ca_out_401;
wire [23:0] u_ca_out_402;
wire [23:0] u_ca_out_403;
wire [23:0] u_ca_out_404;
wire [23:0] u_ca_out_405;
wire [23:0] u_ca_out_406;
wire [23:0] u_ca_out_407;
wire [23:0] u_ca_out_408;
wire [23:0] u_ca_out_409;
wire [23:0] u_ca_out_410;
wire [23:0] u_ca_out_411;
wire [23:0] u_ca_out_412;
wire [23:0] u_ca_out_413;
wire [23:0] u_ca_out_414;
wire [23:0] u_ca_out_415;
wire [23:0] u_ca_out_416;
wire [23:0] u_ca_out_417;
wire [23:0] u_ca_out_418;
wire [23:0] u_ca_out_419;
wire [23:0] u_ca_out_420;
wire [23:0] u_ca_out_421;
wire [23:0] u_ca_out_422;
wire [23:0] u_ca_out_423;
wire [23:0] u_ca_out_424;
wire [23:0] u_ca_out_425;
wire [23:0] u_ca_out_426;
wire [23:0] u_ca_out_427;
wire [23:0] u_ca_out_428;
wire [23:0] u_ca_out_429;
wire [23:0] u_ca_out_430;
wire [23:0] u_ca_out_431;
wire [23:0] u_ca_out_432;
wire [23:0] u_ca_out_433;
wire [23:0] u_ca_out_434;
wire [23:0] u_ca_out_435;
wire [23:0] u_ca_out_436;
wire [23:0] u_ca_out_437;
wire [23:0] u_ca_out_438;
wire [23:0] u_ca_out_439;
wire [23:0] u_ca_out_440;
wire [23:0] u_ca_out_441;
wire [23:0] u_ca_out_442;
wire [23:0] u_ca_out_443;
wire [23:0] u_ca_out_444;
wire [23:0] u_ca_out_445;
wire [23:0] u_ca_out_446;
wire [23:0] u_ca_out_447;
wire [23:0] u_ca_out_448;
wire [23:0] u_ca_out_449;
wire [23:0] u_ca_out_450;
wire [23:0] u_ca_out_451;
wire [23:0] u_ca_out_452;
wire [23:0] u_ca_out_453;
wire [23:0] u_ca_out_454;
wire [23:0] u_ca_out_455;
wire [23:0] u_ca_out_456;
wire [23:0] u_ca_out_457;
wire [23:0] u_ca_out_458;
wire [23:0] u_ca_out_459;
wire [23:0] u_ca_out_460;
wire [23:0] u_ca_out_461;
wire [23:0] u_ca_out_462;
wire [23:0] u_ca_out_463;
wire [23:0] u_ca_out_464;
wire [23:0] u_ca_out_465;
wire [23:0] u_ca_out_466;
wire [23:0] u_ca_out_467;
wire [23:0] u_ca_out_468;
wire [23:0] u_ca_out_469;
wire [23:0] u_ca_out_470;
wire [23:0] u_ca_out_471;
wire [23:0] u_ca_out_472;
wire [23:0] u_ca_out_473;
wire [23:0] u_ca_out_474;
wire [23:0] u_ca_out_475;
wire [23:0] u_ca_out_476;
wire [23:0] u_ca_out_477;
wire [23:0] u_ca_out_478;
wire [23:0] u_ca_out_479;
wire [23:0] u_ca_out_480;
wire [23:0] u_ca_out_481;
wire [23:0] u_ca_out_482;
wire [23:0] u_ca_out_483;
wire [23:0] u_ca_out_484;
wire [23:0] u_ca_out_485;
wire [23:0] u_ca_out_486;
wire [23:0] u_ca_out_487;
wire [23:0] u_ca_out_488;
wire [23:0] u_ca_out_489;
wire [23:0] u_ca_out_490;
wire [23:0] u_ca_out_491;
wire [23:0] u_ca_out_492;
wire [23:0] u_ca_out_493;
wire [23:0] u_ca_out_494;
wire [23:0] u_ca_out_495;
wire [23:0] u_ca_out_496;
wire [23:0] u_ca_out_497;
wire [23:0] u_ca_out_498;
wire [23:0] u_ca_out_499;
wire [23:0] u_ca_out_500;
wire [23:0] u_ca_out_501;
wire [23:0] u_ca_out_502;
wire [23:0] u_ca_out_503;
wire [23:0] u_ca_out_504;
wire [23:0] u_ca_out_505;
wire [23:0] u_ca_out_506;
wire [23:0] u_ca_out_507;
wire [23:0] u_ca_out_508;
wire [23:0] u_ca_out_509;
wire [23:0] u_ca_out_510;
wire [23:0] u_ca_out_511;
wire [23:0] u_ca_out_512;
wire [23:0] u_ca_out_513;
wire [23:0] u_ca_out_514;
wire [23:0] u_ca_out_515;
wire [23:0] u_ca_out_516;
wire [23:0] u_ca_out_517;
wire [23:0] u_ca_out_518;
wire [23:0] u_ca_out_519;
wire [23:0] u_ca_out_520;
wire [23:0] u_ca_out_521;
wire [23:0] u_ca_out_522;
wire [23:0] u_ca_out_523;
wire [23:0] u_ca_out_524;
wire [23:0] u_ca_out_525;
wire [23:0] u_ca_out_526;
wire [23:0] u_ca_out_527;
wire [23:0] u_ca_out_528;
wire [23:0] u_ca_out_529;
wire [23:0] u_ca_out_530;
wire [23:0] u_ca_out_531;
wire [23:0] u_ca_out_532;
wire [23:0] u_ca_out_533;
wire [23:0] u_ca_out_534;
wire [23:0] u_ca_out_535;
wire [23:0] u_ca_out_536;
wire [23:0] u_ca_out_537;
wire [23:0] u_ca_out_538;
wire [23:0] u_ca_out_539;
wire [23:0] u_ca_out_540;
wire [23:0] u_ca_out_541;
wire [23:0] u_ca_out_542;
wire [23:0] u_ca_out_543;
wire [23:0] u_ca_out_544;
wire [23:0] u_ca_out_545;
wire [23:0] u_ca_out_546;
wire [23:0] u_ca_out_547;
wire [23:0] u_ca_out_548;
wire [23:0] u_ca_out_549;
wire [23:0] u_ca_out_550;
wire [23:0] u_ca_out_551;
wire [23:0] u_ca_out_552;
wire [23:0] u_ca_out_553;
wire [23:0] u_ca_out_554;
wire [23:0] u_ca_out_555;
wire [23:0] u_ca_out_556;
wire [23:0] u_ca_out_557;
wire [23:0] u_ca_out_558;
wire [23:0] u_ca_out_559;
wire [23:0] u_ca_out_560;
wire [23:0] u_ca_out_561;
wire [23:0] u_ca_out_562;
wire [23:0] u_ca_out_563;
wire [23:0] u_ca_out_564;
wire [23:0] u_ca_out_565;
wire [23:0] u_ca_out_566;
wire [23:0] u_ca_out_567;
wire [23:0] u_ca_out_568;
wire [23:0] u_ca_out_569;
wire [23:0] u_ca_out_570;
wire [23:0] u_ca_out_571;
wire [23:0] u_ca_out_572;
wire [23:0] u_ca_out_573;
wire [23:0] u_ca_out_574;
wire [23:0] u_ca_out_575;
wire [23:0] u_ca_out_576;
wire [23:0] u_ca_out_577;
wire [23:0] u_ca_out_578;
wire [23:0] u_ca_out_579;
wire [23:0] u_ca_out_580;
wire [23:0] u_ca_out_581;
wire [23:0] u_ca_out_582;
wire [23:0] u_ca_out_583;
wire [23:0] u_ca_out_584;
wire [23:0] u_ca_out_585;
wire [23:0] u_ca_out_586;
wire [23:0] u_ca_out_587;
wire [23:0] u_ca_out_588;
wire [23:0] u_ca_out_589;
wire [23:0] u_ca_out_590;
wire [23:0] u_ca_out_591;
wire [23:0] u_ca_out_592;
wire [23:0] u_ca_out_593;
wire [23:0] u_ca_out_594;
wire [23:0] u_ca_out_595;
wire [23:0] u_ca_out_596;
wire [23:0] u_ca_out_597;
wire [23:0] u_ca_out_598;
wire [23:0] u_ca_out_599;
wire [23:0] u_ca_out_600;
wire [23:0] u_ca_out_601;
wire [23:0] u_ca_out_602;
wire [23:0] u_ca_out_603;
wire [23:0] u_ca_out_604;
wire [23:0] u_ca_out_605;
wire [23:0] u_ca_out_606;
wire [23:0] u_ca_out_607;
wire [23:0] u_ca_out_608;
wire [23:0] u_ca_out_609;
wire [23:0] u_ca_out_610;
wire [23:0] u_ca_out_611;
wire [23:0] u_ca_out_612;
wire [23:0] u_ca_out_613;
wire [23:0] u_ca_out_614;
wire [23:0] u_ca_out_615;
wire [23:0] u_ca_out_616;
wire [23:0] u_ca_out_617;
wire [23:0] u_ca_out_618;
wire [23:0] u_ca_out_619;
wire [23:0] u_ca_out_620;
wire [23:0] u_ca_out_621;
wire [23:0] u_ca_out_622;
wire [23:0] u_ca_out_623;
wire [23:0] u_ca_out_624;
wire [23:0] u_ca_out_625;
wire [23:0] u_ca_out_626;
wire [23:0] u_ca_out_627;
wire [23:0] u_ca_out_628;
wire [23:0] u_ca_out_629;
wire [23:0] u_ca_out_630;
wire [23:0] u_ca_out_631;
wire [23:0] u_ca_out_632;
wire [23:0] u_ca_out_633;
wire [23:0] u_ca_out_634;
wire [23:0] u_ca_out_635;
wire [23:0] u_ca_out_636;
wire [23:0] u_ca_out_637;
wire [23:0] u_ca_out_638;
wire [23:0] u_ca_out_639;
wire [23:0] u_ca_out_640;
wire [23:0] u_ca_out_641;
wire [23:0] u_ca_out_642;
wire [23:0] u_ca_out_643;
wire [23:0] u_ca_out_644;
wire [23:0] u_ca_out_645;
wire [23:0] u_ca_out_646;
wire [23:0] u_ca_out_647;
wire [23:0] u_ca_out_648;
wire [23:0] u_ca_out_649;
wire [23:0] u_ca_out_650;
wire [23:0] u_ca_out_651;
wire [23:0] u_ca_out_652;
wire [23:0] u_ca_out_653;
wire [23:0] u_ca_out_654;
wire [23:0] u_ca_out_655;
wire [23:0] u_ca_out_656;
wire [23:0] u_ca_out_657;
wire [23:0] u_ca_out_658;
wire [23:0] u_ca_out_659;
wire [23:0] u_ca_out_660;
wire [23:0] u_ca_out_661;
wire [23:0] u_ca_out_662;
wire [23:0] u_ca_out_663;
wire [23:0] u_ca_out_664;
wire [23:0] u_ca_out_665;
wire [23:0] u_ca_out_666;
wire [23:0] u_ca_out_667;
wire [23:0] u_ca_out_668;
wire [23:0] u_ca_out_669;
wire [23:0] u_ca_out_670;
wire [23:0] u_ca_out_671;
wire [23:0] u_ca_out_672;
wire [23:0] u_ca_out_673;
wire [23:0] u_ca_out_674;
wire [23:0] u_ca_out_675;
wire [23:0] u_ca_out_676;
wire [23:0] u_ca_out_677;
wire [23:0] u_ca_out_678;
wire [23:0] u_ca_out_679;
wire [23:0] u_ca_out_680;
wire [23:0] u_ca_out_681;
wire [23:0] u_ca_out_682;
wire [23:0] u_ca_out_683;
wire [23:0] u_ca_out_684;
wire [23:0] u_ca_out_685;
wire [23:0] u_ca_out_686;
wire [23:0] u_ca_out_687;
wire [23:0] u_ca_out_688;
wire [23:0] u_ca_out_689;
wire [23:0] u_ca_out_690;
wire [23:0] u_ca_out_691;
wire [23:0] u_ca_out_692;
wire [23:0] u_ca_out_693;
wire [23:0] u_ca_out_694;
wire [23:0] u_ca_out_695;
wire [23:0] u_ca_out_696;
wire [23:0] u_ca_out_697;
wire [23:0] u_ca_out_698;
wire [23:0] u_ca_out_699;
wire [23:0] u_ca_out_700;
wire [23:0] u_ca_out_701;
wire [23:0] u_ca_out_702;
wire [23:0] u_ca_out_703;
wire [23:0] u_ca_out_704;
wire [23:0] u_ca_out_705;
wire [23:0] u_ca_out_706;
wire [23:0] u_ca_out_707;
wire [23:0] u_ca_out_708;
wire [23:0] u_ca_out_709;
wire [23:0] u_ca_out_710;
wire [23:0] u_ca_out_711;
wire [23:0] u_ca_out_712;
wire [23:0] u_ca_out_713;
wire [23:0] u_ca_out_714;
wire [23:0] u_ca_out_715;
wire [23:0] u_ca_out_716;
wire [23:0] u_ca_out_717;
wire [23:0] u_ca_out_718;
wire [23:0] u_ca_out_719;
wire [23:0] u_ca_out_720;
wire [23:0] u_ca_out_721;
wire [23:0] u_ca_out_722;
wire [23:0] u_ca_out_723;
wire [23:0] u_ca_out_724;
wire [23:0] u_ca_out_725;
wire [23:0] u_ca_out_726;
wire [23:0] u_ca_out_727;
wire [23:0] u_ca_out_728;
wire [23:0] u_ca_out_729;
wire [23:0] u_ca_out_730;
wire [23:0] u_ca_out_731;
wire [23:0] u_ca_out_732;
wire [23:0] u_ca_out_733;
wire [23:0] u_ca_out_734;
wire [23:0] u_ca_out_735;
wire [23:0] u_ca_out_736;
wire [23:0] u_ca_out_737;
wire [23:0] u_ca_out_738;
wire [23:0] u_ca_out_739;
wire [23:0] u_ca_out_740;
wire [23:0] u_ca_out_741;
wire [23:0] u_ca_out_742;
wire [23:0] u_ca_out_743;
wire [23:0] u_ca_out_744;
wire [23:0] u_ca_out_745;
wire [23:0] u_ca_out_746;
wire [23:0] u_ca_out_747;
wire [23:0] u_ca_out_748;
wire [23:0] u_ca_out_749;
wire [23:0] u_ca_out_750;
wire [23:0] u_ca_out_751;
wire [23:0] u_ca_out_752;
wire [23:0] u_ca_out_753;
wire [23:0] u_ca_out_754;
wire [23:0] u_ca_out_755;
wire [23:0] u_ca_out_756;
wire [23:0] u_ca_out_757;
wire [23:0] u_ca_out_758;
wire [23:0] u_ca_out_759;
wire [23:0] u_ca_out_760;
wire [23:0] u_ca_out_761;
wire [23:0] u_ca_out_762;
wire [23:0] u_ca_out_763;
wire [23:0] u_ca_out_764;
wire [23:0] u_ca_out_765;
wire [23:0] u_ca_out_766;
wire [23:0] u_ca_out_767;
wire [23:0] u_ca_out_768;
wire [23:0] u_ca_out_769;
wire [23:0] u_ca_out_770;
wire [23:0] u_ca_out_771;
wire [23:0] u_ca_out_772;
wire [23:0] u_ca_out_773;
wire [23:0] u_ca_out_774;
wire [23:0] u_ca_out_775;
wire [23:0] u_ca_out_776;
wire [23:0] u_ca_out_777;
wire [23:0] u_ca_out_778;
wire [23:0] u_ca_out_779;
wire [23:0] u_ca_out_780;
wire [23:0] u_ca_out_781;
wire [23:0] u_ca_out_782;
wire [23:0] u_ca_out_783;
wire [23:0] u_ca_out_784;
wire [23:0] u_ca_out_785;
wire [23:0] u_ca_out_786;
wire [23:0] u_ca_out_787;
wire [23:0] u_ca_out_788;
wire [23:0] u_ca_out_789;
wire [23:0] u_ca_out_790;
wire [23:0] u_ca_out_791;
wire [23:0] u_ca_out_792;
wire [23:0] u_ca_out_793;
wire [23:0] u_ca_out_794;
wire [23:0] u_ca_out_795;
wire [23:0] u_ca_out_796;
wire [23:0] u_ca_out_797;
wire [23:0] u_ca_out_798;
wire [23:0] u_ca_out_799;
wire [23:0] u_ca_out_800;
wire [23:0] u_ca_out_801;
wire [23:0] u_ca_out_802;
wire [23:0] u_ca_out_803;
wire [23:0] u_ca_out_804;
wire [23:0] u_ca_out_805;
wire [23:0] u_ca_out_806;
wire [23:0] u_ca_out_807;
wire [23:0] u_ca_out_808;
wire [23:0] u_ca_out_809;
wire [23:0] u_ca_out_810;
wire [23:0] u_ca_out_811;
wire [23:0] u_ca_out_812;
wire [23:0] u_ca_out_813;
wire [23:0] u_ca_out_814;
wire [23:0] u_ca_out_815;
wire [23:0] u_ca_out_816;
wire [23:0] u_ca_out_817;
wire [23:0] u_ca_out_818;
wire [23:0] u_ca_out_819;
wire [23:0] u_ca_out_820;
wire [23:0] u_ca_out_821;
wire [23:0] u_ca_out_822;
wire [23:0] u_ca_out_823;
wire [23:0] u_ca_out_824;
wire [23:0] u_ca_out_825;
wire [23:0] u_ca_out_826;
wire [23:0] u_ca_out_827;
wire [23:0] u_ca_out_828;
wire [23:0] u_ca_out_829;
wire [23:0] u_ca_out_830;
wire [23:0] u_ca_out_831;
wire [23:0] u_ca_out_832;
wire [23:0] u_ca_out_833;
wire [23:0] u_ca_out_834;
wire [23:0] u_ca_out_835;
wire [23:0] u_ca_out_836;
wire [23:0] u_ca_out_837;
wire [23:0] u_ca_out_838;
wire [23:0] u_ca_out_839;
wire [23:0] u_ca_out_840;
wire [23:0] u_ca_out_841;
wire [23:0] u_ca_out_842;
wire [23:0] u_ca_out_843;
wire [23:0] u_ca_out_844;
wire [23:0] u_ca_out_845;
wire [23:0] u_ca_out_846;
wire [23:0] u_ca_out_847;
wire [23:0] u_ca_out_848;
wire [23:0] u_ca_out_849;
wire [23:0] u_ca_out_850;
wire [23:0] u_ca_out_851;
wire [23:0] u_ca_out_852;
wire [23:0] u_ca_out_853;
wire [23:0] u_ca_out_854;
wire [23:0] u_ca_out_855;
wire [23:0] u_ca_out_856;
wire [23:0] u_ca_out_857;
wire [23:0] u_ca_out_858;
wire [23:0] u_ca_out_859;
wire [23:0] u_ca_out_860;
wire [23:0] u_ca_out_861;
wire [23:0] u_ca_out_862;
wire [23:0] u_ca_out_863;
wire [23:0] u_ca_out_864;
wire [23:0] u_ca_out_865;
wire [23:0] u_ca_out_866;
wire [23:0] u_ca_out_867;
wire [23:0] u_ca_out_868;
wire [23:0] u_ca_out_869;
wire [23:0] u_ca_out_870;
wire [23:0] u_ca_out_871;
wire [23:0] u_ca_out_872;
wire [23:0] u_ca_out_873;
wire [23:0] u_ca_out_874;
wire [23:0] u_ca_out_875;
wire [23:0] u_ca_out_876;
wire [23:0] u_ca_out_877;
wire [23:0] u_ca_out_878;
wire [23:0] u_ca_out_879;
wire [23:0] u_ca_out_880;
wire [23:0] u_ca_out_881;
wire [23:0] u_ca_out_882;
wire [23:0] u_ca_out_883;
wire [23:0] u_ca_out_884;
wire [23:0] u_ca_out_885;
wire [23:0] u_ca_out_886;
wire [23:0] u_ca_out_887;
wire [23:0] u_ca_out_888;
wire [23:0] u_ca_out_889;
wire [23:0] u_ca_out_890;
wire [23:0] u_ca_out_891;
wire [23:0] u_ca_out_892;
wire [23:0] u_ca_out_893;
wire [23:0] u_ca_out_894;
wire [23:0] u_ca_out_895;
wire [23:0] u_ca_out_896;
wire [23:0] u_ca_out_897;
wire [23:0] u_ca_out_898;
wire [23:0] u_ca_out_899;
wire [23:0] u_ca_out_900;
wire [23:0] u_ca_out_901;
wire [23:0] u_ca_out_902;
wire [23:0] u_ca_out_903;
wire [23:0] u_ca_out_904;
wire [23:0] u_ca_out_905;
wire [23:0] u_ca_out_906;
wire [23:0] u_ca_out_907;
wire [23:0] u_ca_out_908;
wire [23:0] u_ca_out_909;
wire [23:0] u_ca_out_910;
wire [23:0] u_ca_out_911;
wire [23:0] u_ca_out_912;
wire [23:0] u_ca_out_913;
wire [23:0] u_ca_out_914;
wire [23:0] u_ca_out_915;
wire [23:0] u_ca_out_916;
wire [23:0] u_ca_out_917;
wire [23:0] u_ca_out_918;
wire [23:0] u_ca_out_919;
wire [23:0] u_ca_out_920;
wire [23:0] u_ca_out_921;
wire [23:0] u_ca_out_922;
wire [23:0] u_ca_out_923;
wire [23:0] u_ca_out_924;
wire [23:0] u_ca_out_925;
wire [23:0] u_ca_out_926;
wire [23:0] u_ca_out_927;
wire [23:0] u_ca_out_928;
wire [23:0] u_ca_out_929;
wire [23:0] u_ca_out_930;
wire [23:0] u_ca_out_931;
wire [23:0] u_ca_out_932;
wire [23:0] u_ca_out_933;
wire [23:0] u_ca_out_934;
wire [23:0] u_ca_out_935;
wire [23:0] u_ca_out_936;
wire [23:0] u_ca_out_937;
wire [23:0] u_ca_out_938;
wire [23:0] u_ca_out_939;
wire [23:0] u_ca_out_940;
wire [23:0] u_ca_out_941;
wire [23:0] u_ca_out_942;
wire [23:0] u_ca_out_943;
wire [23:0] u_ca_out_944;
wire [23:0] u_ca_out_945;
wire [23:0] u_ca_out_946;
wire [23:0] u_ca_out_947;
wire [23:0] u_ca_out_948;
wire [23:0] u_ca_out_949;
wire [23:0] u_ca_out_950;
wire [23:0] u_ca_out_951;
wire [23:0] u_ca_out_952;
wire [23:0] u_ca_out_953;
wire [23:0] u_ca_out_954;
wire [23:0] u_ca_out_955;
wire [23:0] u_ca_out_956;
wire [23:0] u_ca_out_957;
wire [23:0] u_ca_out_958;
wire [23:0] u_ca_out_959;
wire [23:0] u_ca_out_960;
wire [23:0] u_ca_out_961;
wire [23:0] u_ca_out_962;
wire [23:0] u_ca_out_963;
wire [23:0] u_ca_out_964;
wire [23:0] u_ca_out_965;
wire [23:0] u_ca_out_966;
wire [23:0] u_ca_out_967;
wire [23:0] u_ca_out_968;
wire [23:0] u_ca_out_969;
wire [23:0] u_ca_out_970;
wire [23:0] u_ca_out_971;
wire [23:0] u_ca_out_972;
wire [23:0] u_ca_out_973;
wire [23:0] u_ca_out_974;
wire [23:0] u_ca_out_975;
wire [23:0] u_ca_out_976;
wire [23:0] u_ca_out_977;
wire [23:0] u_ca_out_978;
wire [23:0] u_ca_out_979;
wire [23:0] u_ca_out_980;
wire [23:0] u_ca_out_981;
wire [23:0] u_ca_out_982;
wire [23:0] u_ca_out_983;
wire [23:0] u_ca_out_984;
wire [23:0] u_ca_out_985;
wire [23:0] u_ca_out_986;
wire [23:0] u_ca_out_987;
wire [23:0] u_ca_out_988;
wire [23:0] u_ca_out_989;
wire [23:0] u_ca_out_990;
wire [23:0] u_ca_out_991;
wire [23:0] u_ca_out_992;
wire [23:0] u_ca_out_993;
wire [23:0] u_ca_out_994;
wire [23:0] u_ca_out_995;
wire [23:0] u_ca_out_996;
wire [23:0] u_ca_out_997;
wire [23:0] u_ca_out_998;
wire [23:0] u_ca_out_999;
wire [23:0] u_ca_out_1000;
wire [23:0] u_ca_out_1001;
wire [23:0] u_ca_out_1002;
wire [23:0] u_ca_out_1003;
wire [23:0] u_ca_out_1004;
wire [23:0] u_ca_out_1005;
wire [23:0] u_ca_out_1006;
wire [23:0] u_ca_out_1007;
wire [23:0] u_ca_out_1008;
wire [23:0] u_ca_out_1009;
wire [23:0] u_ca_out_1010;
wire [23:0] u_ca_out_1011;
wire [23:0] u_ca_out_1012;
wire [23:0] u_ca_out_1013;
wire [23:0] u_ca_out_1014;
wire [23:0] u_ca_out_1015;
wire [23:0] u_ca_out_1016;
wire [23:0] u_ca_out_1017;
wire [23:0] u_ca_out_1018;
wire [23:0] u_ca_out_1019;
wire [23:0] u_ca_out_1020;
wire [23:0] u_ca_out_1021;
wire [23:0] u_ca_out_1022;
wire [23:0] u_ca_out_1023;
wire [23:0] u_ca_out_1024;
wire [23:0] u_ca_out_1025;
wire [23:0] u_ca_out_1026;
wire [23:0] u_ca_out_1027;
wire [23:0] u_ca_out_1028;
wire [23:0] u_ca_out_1029;
wire [23:0] u_ca_out_1030;
wire [23:0] u_ca_out_1031;
wire [23:0] u_ca_out_1032;
wire [23:0] u_ca_out_1033;
wire [23:0] u_ca_out_1034;
wire [23:0] u_ca_out_1035;
wire [23:0] u_ca_out_1036;
wire [23:0] u_ca_out_1037;
wire [23:0] u_ca_out_1038;
wire [23:0] u_ca_out_1039;
wire [23:0] u_ca_out_1040;
wire [23:0] u_ca_out_1041;
wire [23:0] u_ca_out_1042;
wire [23:0] u_ca_out_1043;
wire [23:0] u_ca_out_1044;
wire [23:0] u_ca_out_1045;
wire [23:0] u_ca_out_1046;
wire [23:0] u_ca_out_1047;
wire [23:0] u_ca_out_1048;
wire [23:0] u_ca_out_1049;
wire [23:0] u_ca_out_1050;
wire [23:0] u_ca_out_1051;
wire [23:0] u_ca_out_1052;
wire [23:0] u_ca_out_1053;
wire [23:0] u_ca_out_1054;
wire [23:0] u_ca_out_1055;
wire [23:0] u_ca_out_1056;
wire [23:0] u_ca_out_1057;
wire [23:0] u_ca_out_1058;
wire [23:0] u_ca_out_1059;
wire [23:0] u_ca_out_1060;
wire [23:0] u_ca_out_1061;
wire [23:0] u_ca_out_1062;
wire [23:0] u_ca_out_1063;
wire [23:0] u_ca_out_1064;
wire [23:0] u_ca_out_1065;
wire [23:0] u_ca_out_1066;
wire [23:0] u_ca_out_1067;
wire [23:0] u_ca_out_1068;
wire [23:0] u_ca_out_1069;
wire [23:0] u_ca_out_1070;
wire [23:0] u_ca_out_1071;
wire [23:0] u_ca_out_1072;
wire [23:0] u_ca_out_1073;
wire [23:0] u_ca_out_1074;
wire [23:0] u_ca_out_1075;
wire [23:0] u_ca_out_1076;
wire [23:0] u_ca_out_1077;
wire [23:0] u_ca_out_1078;
wire [23:0] u_ca_out_1079;
wire [23:0] u_ca_out_1080;
wire [23:0] u_ca_out_1081;
wire [23:0] u_ca_out_1082;
wire [23:0] u_ca_out_1083;
wire [23:0] u_ca_out_1084;
wire [23:0] u_ca_out_1085;
wire [23:0] u_ca_out_1086;
wire [23:0] u_ca_out_1087;
wire [23:0] u_ca_out_1088;
wire [23:0] u_ca_out_1089;
wire [23:0] u_ca_out_1090;
wire [23:0] u_ca_out_1091;
wire [23:0] u_ca_out_1092;
wire [23:0] u_ca_out_1093;
wire [23:0] u_ca_out_1094;
wire [23:0] u_ca_out_1095;
wire [23:0] u_ca_out_1096;
wire [23:0] u_ca_out_1097;
wire [23:0] u_ca_out_1098;
wire [23:0] u_ca_out_1099;
wire [23:0] u_ca_out_1100;
wire [23:0] u_ca_out_1101;
wire [23:0] u_ca_out_1102;
wire [23:0] u_ca_out_1103;
wire [23:0] u_ca_out_1104;
wire [23:0] u_ca_out_1105;
wire [23:0] u_ca_out_1106;
wire [23:0] u_ca_out_1107;
wire [23:0] u_ca_out_1108;
wire [23:0] u_ca_out_1109;
wire [23:0] u_ca_out_1110;
wire [23:0] u_ca_out_1111;
wire [23:0] u_ca_out_1112;
wire [23:0] u_ca_out_1113;
wire [23:0] u_ca_out_1114;
wire [23:0] u_ca_out_1115;
wire [23:0] u_ca_out_1116;
wire [23:0] u_ca_out_1117;
wire [23:0] u_ca_out_1118;
wire [23:0] u_ca_out_1119;
wire [23:0] u_ca_out_1120;
wire [23:0] u_ca_out_1121;
wire [23:0] u_ca_out_1122;
wire [23:0] u_ca_out_1123;
wire [23:0] u_ca_out_1124;
wire [23:0] u_ca_out_1125;
wire [23:0] u_ca_out_1126;
wire [23:0] u_ca_out_1127;
wire [23:0] u_ca_out_1128;
wire [23:0] u_ca_out_1129;
wire [23:0] u_ca_out_1130;
wire [23:0] u_ca_out_1131;
wire [23:0] u_ca_out_1132;
wire [23:0] u_ca_out_1133;
wire [23:0] u_ca_out_1134;
wire [23:0] u_ca_out_1135;
wire [23:0] u_ca_out_1136;
wire [23:0] u_ca_out_1137;
wire [23:0] u_ca_out_1138;
wire [23:0] u_ca_out_1139;
wire [23:0] u_ca_out_1140;
wire [23:0] u_ca_out_1141;
wire [23:0] u_ca_out_1142;
wire [23:0] u_ca_out_1143;
wire [23:0] u_ca_out_1144;
wire [23:0] u_ca_out_1145;
wire [23:0] u_ca_out_1146;
wire [23:0] u_ca_out_1147;
wire [23:0] u_ca_out_1148;
wire [23:0] u_ca_out_1149;
wire [23:0] u_ca_out_1150;
wire [23:0] u_ca_out_1151;
wire [23:0] u_ca_out_1152;
wire [23:0] u_ca_out_1153;
wire [23:0] u_ca_out_1154;
wire [23:0] u_ca_out_1155;
wire [23:0] u_ca_out_1156;
wire [23:0] u_ca_out_1157;
wire [23:0] u_ca_out_1158;
wire [23:0] u_ca_out_1159;
wire [23:0] u_ca_out_1160;
wire [23:0] u_ca_out_1161;
wire [23:0] u_ca_out_1162;
wire [23:0] u_ca_out_1163;
wire [23:0] u_ca_out_1164;
wire [23:0] u_ca_out_1165;
wire [23:0] u_ca_out_1166;
wire [23:0] u_ca_out_1167;
wire [23:0] u_ca_out_1168;
wire [23:0] u_ca_out_1169;
wire [23:0] u_ca_out_1170;
wire [23:0] u_ca_out_1171;
wire [23:0] u_ca_out_1172;
wire [23:0] u_ca_out_1173;
wire [23:0] u_ca_out_1174;
wire [23:0] u_ca_out_1175;
wire [23:0] u_ca_out_1176;
wire [23:0] u_ca_out_1177;
wire [23:0] u_ca_out_1178;
wire [23:0] u_ca_out_1179;
wire [23:0] u_ca_out_1180;
wire [23:0] u_ca_out_1181;
wire [23:0] u_ca_out_1182;
wire [23:0] u_ca_out_1183;
wire [23:0] u_ca_out_1184;
wire [23:0] u_ca_out_1185;
wire [23:0] u_ca_out_1186;
wire [23:0] u_ca_out_1187;
wire [23:0] u_ca_out_1188;
wire [23:0] u_ca_out_1189;
wire [23:0] u_ca_out_1190;
wire [23:0] u_ca_out_1191;
wire [23:0] u_ca_out_1192;
wire [23:0] u_ca_out_1193;
wire [23:0] u_ca_out_1194;
wire [23:0] u_ca_out_1195;
wire [23:0] u_ca_out_1196;
wire [23:0] u_ca_out_1197;
wire [23:0] u_ca_out_1198;
wire [23:0] u_ca_out_1199;
wire [23:0] u_ca_out_1200;
wire [23:0] u_ca_out_1201;
wire [23:0] u_ca_out_1202;
wire [23:0] u_ca_out_1203;
wire [23:0] u_ca_out_1204;
wire [23:0] u_ca_out_1205;
wire [23:0] u_ca_out_1206;
wire [23:0] u_ca_out_1207;
wire [23:0] u_ca_out_1208;
wire [23:0] u_ca_out_1209;
wire [23:0] u_ca_out_1210;
wire [23:0] u_ca_out_1211;
wire [23:0] u_ca_out_1212;
wire [23:0] u_ca_out_1213;
wire [23:0] u_ca_out_1214;
wire [23:0] u_ca_out_1215;
wire [23:0] u_ca_out_1216;
wire [23:0] u_ca_out_1217;
wire [23:0] u_ca_out_1218;
wire [23:0] u_ca_out_1219;
wire [23:0] u_ca_out_1220;
wire [23:0] u_ca_out_1221;
wire [23:0] u_ca_out_1222;
wire [23:0] u_ca_out_1223;
wire [23:0] u_ca_out_1224;
wire [23:0] u_ca_out_1225;
wire [23:0] u_ca_out_1226;
wire [23:0] u_ca_out_1227;
wire [23:0] u_ca_out_1228;
wire [23:0] u_ca_out_1229;
wire [23:0] u_ca_out_1230;
wire [23:0] u_ca_out_1231;
wire [23:0] u_ca_out_1232;
wire [23:0] u_ca_out_1233;
wire [23:0] u_ca_out_1234;
wire [23:0] u_ca_out_1235;
wire [23:0] u_ca_out_1236;
wire [23:0] u_ca_out_1237;
wire [23:0] u_ca_out_1238;
wire [23:0] u_ca_out_1239;
wire [23:0] u_ca_out_1240;
wire [23:0] u_ca_out_1241;
wire [23:0] u_ca_out_1242;
wire [23:0] u_ca_out_1243;
wire [23:0] u_ca_out_1244;
wire [23:0] u_ca_out_1245;
wire [23:0] u_ca_out_1246;
wire [23:0] u_ca_out_1247;
wire [23:0] u_ca_out_1248;
wire [23:0] u_ca_out_1249;
wire [23:0] u_ca_out_1250;
wire [23:0] u_ca_out_1251;
wire [23:0] u_ca_out_1252;
wire [23:0] u_ca_out_1253;
wire [23:0] u_ca_out_1254;
wire [23:0] u_ca_out_1255;
wire [23:0] u_ca_out_1256;
wire [23:0] u_ca_out_1257;
wire [23:0] u_ca_out_1258;
wire [23:0] u_ca_out_1259;
wire [23:0] u_ca_out_1260;
wire [23:0] u_ca_out_1261;
wire [23:0] u_ca_out_1262;
wire [23:0] u_ca_out_1263;
wire [23:0] u_ca_out_1264;
wire [23:0] u_ca_out_1265;
wire [23:0] u_ca_out_1266;
wire [23:0] u_ca_out_1267;
wire [23:0] u_ca_out_1268;
wire [23:0] u_ca_out_1269;
wire [23:0] u_ca_out_1270;
wire [23:0] u_ca_out_1271;
wire [23:0] u_ca_out_1272;
wire [23:0] u_ca_out_1273;
wire [23:0] u_ca_out_1274;
wire [23:0] u_ca_out_1275;
wire [23:0] u_ca_out_1276;
wire [23:0] u_ca_out_1277;
wire [23:0] u_ca_out_1278;
wire [23:0] u_ca_out_1279;
wire [23:0] u_ca_out_1280;
wire [23:0] u_ca_out_1281;
wire [23:0] u_ca_out_1282;

assign u_ca_in_0 = {{9{1'b0}}, col_in_0};
assign u_ca_in_1 = {{9{1'b0}}, col_in_1};
assign u_ca_in_2 = {{9{1'b0}}, col_in_2};
assign u_ca_in_3 = {{9{1'b0}}, col_in_3};
assign u_ca_in_4 = {{9{1'b0}}, col_in_4};
assign u_ca_in_5 = {{9{1'b0}}, col_in_5};
assign u_ca_in_6 = {{9{1'b0}}, col_in_6};
assign u_ca_in_7 = {{9{1'b0}}, col_in_7};
assign u_ca_in_8 = {{9{1'b0}}, col_in_8};
assign u_ca_in_9 = {{9{1'b0}}, col_in_9};
assign u_ca_in_10 = {{9{1'b0}}, col_in_10};
assign u_ca_in_11 = {{9{1'b0}}, col_in_11};
assign u_ca_in_12 = {{9{1'b0}}, col_in_12};
assign u_ca_in_13 = {{9{1'b0}}, col_in_13};
assign u_ca_in_14 = {{9{1'b0}}, col_in_14};
assign u_ca_in_15 = {{9{1'b0}}, col_in_15};
assign u_ca_in_16 = {{9{1'b0}}, col_in_16};
assign u_ca_in_17 = {{9{1'b0}}, col_in_17};
assign u_ca_in_18 = {{9{1'b0}}, col_in_18};
assign u_ca_in_19 = {{9{1'b0}}, col_in_19};
assign u_ca_in_20 = {{9{1'b0}}, col_in_20};
assign u_ca_in_21 = {{9{1'b0}}, col_in_21};
assign u_ca_in_22 = {{9{1'b0}}, col_in_22};
assign u_ca_in_23 = {{9{1'b0}}, col_in_23};
assign u_ca_in_24 = {{9{1'b0}}, col_in_24};
assign u_ca_in_25 = {{9{1'b0}}, col_in_25};
assign u_ca_in_26 = {{9{1'b0}}, col_in_26};
assign u_ca_in_27 = {{9{1'b0}}, col_in_27};
assign u_ca_in_28 = {{9{1'b0}}, col_in_28};
assign u_ca_in_29 = {{9{1'b0}}, col_in_29};
assign u_ca_in_30 = {{9{1'b0}}, col_in_30};
assign u_ca_in_31 = {{9{1'b0}}, col_in_31};
assign u_ca_in_32 = {{9{1'b0}}, col_in_32};
assign u_ca_in_33 = {{9{1'b0}}, col_in_33};
assign u_ca_in_34 = {{9{1'b0}}, col_in_34};
assign u_ca_in_35 = {{9{1'b0}}, col_in_35};
assign u_ca_in_36 = {{9{1'b0}}, col_in_36};
assign u_ca_in_37 = {{9{1'b0}}, col_in_37};
assign u_ca_in_38 = {{9{1'b0}}, col_in_38};
assign u_ca_in_39 = {{9{1'b0}}, col_in_39};
assign u_ca_in_40 = {{9{1'b0}}, col_in_40};
assign u_ca_in_41 = {{9{1'b0}}, col_in_41};
assign u_ca_in_42 = {{9{1'b0}}, col_in_42};
assign u_ca_in_43 = {{9{1'b0}}, col_in_43};
assign u_ca_in_44 = {{9{1'b0}}, col_in_44};
assign u_ca_in_45 = {{9{1'b0}}, col_in_45};
assign u_ca_in_46 = {{9{1'b0}}, col_in_46};
assign u_ca_in_47 = {{9{1'b0}}, col_in_47};
assign u_ca_in_48 = {{9{1'b0}}, col_in_48};
assign u_ca_in_49 = {{9{1'b0}}, col_in_49};
assign u_ca_in_50 = {{9{1'b0}}, col_in_50};
assign u_ca_in_51 = {{9{1'b0}}, col_in_51};
assign u_ca_in_52 = {{9{1'b0}}, col_in_52};
assign u_ca_in_53 = {{9{1'b0}}, col_in_53};
assign u_ca_in_54 = {{9{1'b0}}, col_in_54};
assign u_ca_in_55 = {{9{1'b0}}, col_in_55};
assign u_ca_in_56 = {{9{1'b0}}, col_in_56};
assign u_ca_in_57 = {{9{1'b0}}, col_in_57};
assign u_ca_in_58 = {{9{1'b0}}, col_in_58};
assign u_ca_in_59 = {{9{1'b0}}, col_in_59};
assign u_ca_in_60 = {{9{1'b0}}, col_in_60};
assign u_ca_in_61 = {{9{1'b0}}, col_in_61};
assign u_ca_in_62 = {{9{1'b0}}, col_in_62};
assign u_ca_in_63 = {{9{1'b0}}, col_in_63};
assign u_ca_in_64 = {{9{1'b0}}, col_in_64};
assign u_ca_in_65 = {{9{1'b0}}, col_in_65};
assign u_ca_in_66 = {{9{1'b0}}, col_in_66};
assign u_ca_in_67 = {{9{1'b0}}, col_in_67};
assign u_ca_in_68 = {{9{1'b0}}, col_in_68};
assign u_ca_in_69 = {{9{1'b0}}, col_in_69};
assign u_ca_in_70 = {{9{1'b0}}, col_in_70};
assign u_ca_in_71 = {{9{1'b0}}, col_in_71};
assign u_ca_in_72 = {{9{1'b0}}, col_in_72};
assign u_ca_in_73 = {{9{1'b0}}, col_in_73};
assign u_ca_in_74 = {{9{1'b0}}, col_in_74};
assign u_ca_in_75 = {{9{1'b0}}, col_in_75};
assign u_ca_in_76 = {{9{1'b0}}, col_in_76};
assign u_ca_in_77 = {{9{1'b0}}, col_in_77};
assign u_ca_in_78 = {{9{1'b0}}, col_in_78};
assign u_ca_in_79 = {{9{1'b0}}, col_in_79};
assign u_ca_in_80 = {{9{1'b0}}, col_in_80};
assign u_ca_in_81 = {{9{1'b0}}, col_in_81};
assign u_ca_in_82 = {{9{1'b0}}, col_in_82};
assign u_ca_in_83 = {{9{1'b0}}, col_in_83};
assign u_ca_in_84 = {{9{1'b0}}, col_in_84};
assign u_ca_in_85 = {{9{1'b0}}, col_in_85};
assign u_ca_in_86 = {{9{1'b0}}, col_in_86};
assign u_ca_in_87 = {{9{1'b0}}, col_in_87};
assign u_ca_in_88 = {{9{1'b0}}, col_in_88};
assign u_ca_in_89 = {{9{1'b0}}, col_in_89};
assign u_ca_in_90 = {{9{1'b0}}, col_in_90};
assign u_ca_in_91 = {{9{1'b0}}, col_in_91};
assign u_ca_in_92 = {{9{1'b0}}, col_in_92};
assign u_ca_in_93 = {{9{1'b0}}, col_in_93};
assign u_ca_in_94 = {{9{1'b0}}, col_in_94};
assign u_ca_in_95 = {{9{1'b0}}, col_in_95};
assign u_ca_in_96 = {{9{1'b0}}, col_in_96};
assign u_ca_in_97 = {{9{1'b0}}, col_in_97};
assign u_ca_in_98 = {{9{1'b0}}, col_in_98};
assign u_ca_in_99 = {{9{1'b0}}, col_in_99};
assign u_ca_in_100 = {{9{1'b0}}, col_in_100};
assign u_ca_in_101 = {{9{1'b0}}, col_in_101};
assign u_ca_in_102 = {{9{1'b0}}, col_in_102};
assign u_ca_in_103 = {{9{1'b0}}, col_in_103};
assign u_ca_in_104 = {{9{1'b0}}, col_in_104};
assign u_ca_in_105 = {{9{1'b0}}, col_in_105};
assign u_ca_in_106 = {{9{1'b0}}, col_in_106};
assign u_ca_in_107 = {{9{1'b0}}, col_in_107};
assign u_ca_in_108 = {{9{1'b0}}, col_in_108};
assign u_ca_in_109 = {{9{1'b0}}, col_in_109};
assign u_ca_in_110 = {{9{1'b0}}, col_in_110};
assign u_ca_in_111 = {{9{1'b0}}, col_in_111};
assign u_ca_in_112 = {{9{1'b0}}, col_in_112};
assign u_ca_in_113 = {{9{1'b0}}, col_in_113};
assign u_ca_in_114 = {{9{1'b0}}, col_in_114};
assign u_ca_in_115 = {{9{1'b0}}, col_in_115};
assign u_ca_in_116 = {{9{1'b0}}, col_in_116};
assign u_ca_in_117 = {{9{1'b0}}, col_in_117};
assign u_ca_in_118 = {{9{1'b0}}, col_in_118};
assign u_ca_in_119 = {{9{1'b0}}, col_in_119};
assign u_ca_in_120 = {{9{1'b0}}, col_in_120};
assign u_ca_in_121 = {{9{1'b0}}, col_in_121};
assign u_ca_in_122 = {{9{1'b0}}, col_in_122};
assign u_ca_in_123 = {{9{1'b0}}, col_in_123};
assign u_ca_in_124 = {{9{1'b0}}, col_in_124};
assign u_ca_in_125 = {{9{1'b0}}, col_in_125};
assign u_ca_in_126 = {{9{1'b0}}, col_in_126};
assign u_ca_in_127 = {{9{1'b0}}, col_in_127};
assign u_ca_in_128 = {{9{1'b0}}, col_in_128};
assign u_ca_in_129 = {{9{1'b0}}, col_in_129};
assign u_ca_in_130 = {{9{1'b0}}, col_in_130};
assign u_ca_in_131 = {{9{1'b0}}, col_in_131};
assign u_ca_in_132 = {{9{1'b0}}, col_in_132};
assign u_ca_in_133 = {{9{1'b0}}, col_in_133};
assign u_ca_in_134 = {{9{1'b0}}, col_in_134};
assign u_ca_in_135 = {{9{1'b0}}, col_in_135};
assign u_ca_in_136 = {{9{1'b0}}, col_in_136};
assign u_ca_in_137 = {{9{1'b0}}, col_in_137};
assign u_ca_in_138 = {{9{1'b0}}, col_in_138};
assign u_ca_in_139 = {{9{1'b0}}, col_in_139};
assign u_ca_in_140 = {{9{1'b0}}, col_in_140};
assign u_ca_in_141 = {{9{1'b0}}, col_in_141};
assign u_ca_in_142 = {{9{1'b0}}, col_in_142};
assign u_ca_in_143 = {{9{1'b0}}, col_in_143};
assign u_ca_in_144 = {{9{1'b0}}, col_in_144};
assign u_ca_in_145 = {{9{1'b0}}, col_in_145};
assign u_ca_in_146 = {{9{1'b0}}, col_in_146};
assign u_ca_in_147 = {{9{1'b0}}, col_in_147};
assign u_ca_in_148 = {{9{1'b0}}, col_in_148};
assign u_ca_in_149 = {{9{1'b0}}, col_in_149};
assign u_ca_in_150 = {{9{1'b0}}, col_in_150};
assign u_ca_in_151 = {{9{1'b0}}, col_in_151};
assign u_ca_in_152 = {{9{1'b0}}, col_in_152};
assign u_ca_in_153 = {{9{1'b0}}, col_in_153};
assign u_ca_in_154 = {{9{1'b0}}, col_in_154};
assign u_ca_in_155 = {{9{1'b0}}, col_in_155};
assign u_ca_in_156 = {{9{1'b0}}, col_in_156};
assign u_ca_in_157 = {{9{1'b0}}, col_in_157};
assign u_ca_in_158 = {{9{1'b0}}, col_in_158};
assign u_ca_in_159 = {{9{1'b0}}, col_in_159};
assign u_ca_in_160 = {{9{1'b0}}, col_in_160};
assign u_ca_in_161 = {{9{1'b0}}, col_in_161};
assign u_ca_in_162 = {{9{1'b0}}, col_in_162};
assign u_ca_in_163 = {{9{1'b0}}, col_in_163};
assign u_ca_in_164 = {{9{1'b0}}, col_in_164};
assign u_ca_in_165 = {{9{1'b0}}, col_in_165};
assign u_ca_in_166 = {{9{1'b0}}, col_in_166};
assign u_ca_in_167 = {{9{1'b0}}, col_in_167};
assign u_ca_in_168 = {{9{1'b0}}, col_in_168};
assign u_ca_in_169 = {{9{1'b0}}, col_in_169};
assign u_ca_in_170 = {{9{1'b0}}, col_in_170};
assign u_ca_in_171 = {{9{1'b0}}, col_in_171};
assign u_ca_in_172 = {{9{1'b0}}, col_in_172};
assign u_ca_in_173 = {{9{1'b0}}, col_in_173};
assign u_ca_in_174 = {{9{1'b0}}, col_in_174};
assign u_ca_in_175 = {{9{1'b0}}, col_in_175};
assign u_ca_in_176 = {{9{1'b0}}, col_in_176};
assign u_ca_in_177 = {{9{1'b0}}, col_in_177};
assign u_ca_in_178 = {{9{1'b0}}, col_in_178};
assign u_ca_in_179 = {{9{1'b0}}, col_in_179};
assign u_ca_in_180 = {{9{1'b0}}, col_in_180};
assign u_ca_in_181 = {{9{1'b0}}, col_in_181};
assign u_ca_in_182 = {{9{1'b0}}, col_in_182};
assign u_ca_in_183 = {{9{1'b0}}, col_in_183};
assign u_ca_in_184 = {{9{1'b0}}, col_in_184};
assign u_ca_in_185 = {{9{1'b0}}, col_in_185};
assign u_ca_in_186 = {{9{1'b0}}, col_in_186};
assign u_ca_in_187 = {{9{1'b0}}, col_in_187};
assign u_ca_in_188 = {{9{1'b0}}, col_in_188};
assign u_ca_in_189 = {{9{1'b0}}, col_in_189};
assign u_ca_in_190 = {{9{1'b0}}, col_in_190};
assign u_ca_in_191 = {{9{1'b0}}, col_in_191};
assign u_ca_in_192 = {{9{1'b0}}, col_in_192};
assign u_ca_in_193 = {{9{1'b0}}, col_in_193};
assign u_ca_in_194 = {{9{1'b0}}, col_in_194};
assign u_ca_in_195 = {{9{1'b0}}, col_in_195};
assign u_ca_in_196 = {{9{1'b0}}, col_in_196};
assign u_ca_in_197 = {{9{1'b0}}, col_in_197};
assign u_ca_in_198 = {{9{1'b0}}, col_in_198};
assign u_ca_in_199 = {{9{1'b0}}, col_in_199};
assign u_ca_in_200 = {{9{1'b0}}, col_in_200};
assign u_ca_in_201 = {{9{1'b0}}, col_in_201};
assign u_ca_in_202 = {{9{1'b0}}, col_in_202};
assign u_ca_in_203 = {{9{1'b0}}, col_in_203};
assign u_ca_in_204 = {{9{1'b0}}, col_in_204};
assign u_ca_in_205 = {{9{1'b0}}, col_in_205};
assign u_ca_in_206 = {{9{1'b0}}, col_in_206};
assign u_ca_in_207 = {{9{1'b0}}, col_in_207};
assign u_ca_in_208 = {{9{1'b0}}, col_in_208};
assign u_ca_in_209 = {{9{1'b0}}, col_in_209};
assign u_ca_in_210 = {{9{1'b0}}, col_in_210};
assign u_ca_in_211 = {{9{1'b0}}, col_in_211};
assign u_ca_in_212 = {{9{1'b0}}, col_in_212};
assign u_ca_in_213 = {{9{1'b0}}, col_in_213};
assign u_ca_in_214 = {{9{1'b0}}, col_in_214};
assign u_ca_in_215 = {{9{1'b0}}, col_in_215};
assign u_ca_in_216 = {{9{1'b0}}, col_in_216};
assign u_ca_in_217 = {{9{1'b0}}, col_in_217};
assign u_ca_in_218 = {{9{1'b0}}, col_in_218};
assign u_ca_in_219 = {{9{1'b0}}, col_in_219};
assign u_ca_in_220 = {{9{1'b0}}, col_in_220};
assign u_ca_in_221 = {{9{1'b0}}, col_in_221};
assign u_ca_in_222 = {{9{1'b0}}, col_in_222};
assign u_ca_in_223 = {{9{1'b0}}, col_in_223};
assign u_ca_in_224 = {{9{1'b0}}, col_in_224};
assign u_ca_in_225 = {{9{1'b0}}, col_in_225};
assign u_ca_in_226 = {{9{1'b0}}, col_in_226};
assign u_ca_in_227 = {{9{1'b0}}, col_in_227};
assign u_ca_in_228 = {{9{1'b0}}, col_in_228};
assign u_ca_in_229 = {{9{1'b0}}, col_in_229};
assign u_ca_in_230 = {{9{1'b0}}, col_in_230};
assign u_ca_in_231 = {{9{1'b0}}, col_in_231};
assign u_ca_in_232 = {{9{1'b0}}, col_in_232};
assign u_ca_in_233 = {{9{1'b0}}, col_in_233};
assign u_ca_in_234 = {{9{1'b0}}, col_in_234};
assign u_ca_in_235 = {{9{1'b0}}, col_in_235};
assign u_ca_in_236 = {{9{1'b0}}, col_in_236};
assign u_ca_in_237 = {{9{1'b0}}, col_in_237};
assign u_ca_in_238 = {{9{1'b0}}, col_in_238};
assign u_ca_in_239 = {{9{1'b0}}, col_in_239};
assign u_ca_in_240 = {{9{1'b0}}, col_in_240};
assign u_ca_in_241 = {{9{1'b0}}, col_in_241};
assign u_ca_in_242 = {{9{1'b0}}, col_in_242};
assign u_ca_in_243 = {{9{1'b0}}, col_in_243};
assign u_ca_in_244 = {{9{1'b0}}, col_in_244};
assign u_ca_in_245 = {{9{1'b0}}, col_in_245};
assign u_ca_in_246 = {{9{1'b0}}, col_in_246};
assign u_ca_in_247 = {{9{1'b0}}, col_in_247};
assign u_ca_in_248 = {{9{1'b0}}, col_in_248};
assign u_ca_in_249 = {{9{1'b0}}, col_in_249};
assign u_ca_in_250 = {{9{1'b0}}, col_in_250};
assign u_ca_in_251 = {{9{1'b0}}, col_in_251};
assign u_ca_in_252 = {{9{1'b0}}, col_in_252};
assign u_ca_in_253 = {{9{1'b0}}, col_in_253};
assign u_ca_in_254 = {{9{1'b0}}, col_in_254};
assign u_ca_in_255 = {{9{1'b0}}, col_in_255};
assign u_ca_in_256 = {{9{1'b0}}, col_in_256};
assign u_ca_in_257 = {{9{1'b0}}, col_in_257};
assign u_ca_in_258 = {{9{1'b0}}, col_in_258};
assign u_ca_in_259 = {{9{1'b0}}, col_in_259};
assign u_ca_in_260 = {{9{1'b0}}, col_in_260};
assign u_ca_in_261 = {{9{1'b0}}, col_in_261};
assign u_ca_in_262 = {{9{1'b0}}, col_in_262};
assign u_ca_in_263 = {{9{1'b0}}, col_in_263};
assign u_ca_in_264 = {{9{1'b0}}, col_in_264};
assign u_ca_in_265 = {{9{1'b0}}, col_in_265};
assign u_ca_in_266 = {{9{1'b0}}, col_in_266};
assign u_ca_in_267 = {{9{1'b0}}, col_in_267};
assign u_ca_in_268 = {{9{1'b0}}, col_in_268};
assign u_ca_in_269 = {{9{1'b0}}, col_in_269};
assign u_ca_in_270 = {{9{1'b0}}, col_in_270};
assign u_ca_in_271 = {{9{1'b0}}, col_in_271};
assign u_ca_in_272 = {{9{1'b0}}, col_in_272};
assign u_ca_in_273 = {{9{1'b0}}, col_in_273};
assign u_ca_in_274 = {{9{1'b0}}, col_in_274};
assign u_ca_in_275 = {{9{1'b0}}, col_in_275};
assign u_ca_in_276 = {{9{1'b0}}, col_in_276};
assign u_ca_in_277 = {{9{1'b0}}, col_in_277};
assign u_ca_in_278 = {{9{1'b0}}, col_in_278};
assign u_ca_in_279 = {{9{1'b0}}, col_in_279};
assign u_ca_in_280 = {{9{1'b0}}, col_in_280};
assign u_ca_in_281 = {{9{1'b0}}, col_in_281};
assign u_ca_in_282 = {{9{1'b0}}, col_in_282};
assign u_ca_in_283 = {{9{1'b0}}, col_in_283};
assign u_ca_in_284 = {{9{1'b0}}, col_in_284};
assign u_ca_in_285 = {{9{1'b0}}, col_in_285};
assign u_ca_in_286 = {{9{1'b0}}, col_in_286};
assign u_ca_in_287 = {{9{1'b0}}, col_in_287};
assign u_ca_in_288 = {{9{1'b0}}, col_in_288};
assign u_ca_in_289 = {{9{1'b0}}, col_in_289};
assign u_ca_in_290 = {{9{1'b0}}, col_in_290};
assign u_ca_in_291 = {{9{1'b0}}, col_in_291};
assign u_ca_in_292 = {{9{1'b0}}, col_in_292};
assign u_ca_in_293 = {{9{1'b0}}, col_in_293};
assign u_ca_in_294 = {{9{1'b0}}, col_in_294};
assign u_ca_in_295 = {{9{1'b0}}, col_in_295};
assign u_ca_in_296 = {{9{1'b0}}, col_in_296};
assign u_ca_in_297 = {{9{1'b0}}, col_in_297};
assign u_ca_in_298 = {{9{1'b0}}, col_in_298};
assign u_ca_in_299 = {{9{1'b0}}, col_in_299};
assign u_ca_in_300 = {{9{1'b0}}, col_in_300};
assign u_ca_in_301 = {{9{1'b0}}, col_in_301};
assign u_ca_in_302 = {{9{1'b0}}, col_in_302};
assign u_ca_in_303 = {{9{1'b0}}, col_in_303};
assign u_ca_in_304 = {{9{1'b0}}, col_in_304};
assign u_ca_in_305 = {{9{1'b0}}, col_in_305};
assign u_ca_in_306 = {{9{1'b0}}, col_in_306};
assign u_ca_in_307 = {{9{1'b0}}, col_in_307};
assign u_ca_in_308 = {{9{1'b0}}, col_in_308};
assign u_ca_in_309 = {{9{1'b0}}, col_in_309};
assign u_ca_in_310 = {{9{1'b0}}, col_in_310};
assign u_ca_in_311 = {{9{1'b0}}, col_in_311};
assign u_ca_in_312 = {{9{1'b0}}, col_in_312};
assign u_ca_in_313 = {{9{1'b0}}, col_in_313};
assign u_ca_in_314 = {{9{1'b0}}, col_in_314};
assign u_ca_in_315 = {{9{1'b0}}, col_in_315};
assign u_ca_in_316 = {{9{1'b0}}, col_in_316};
assign u_ca_in_317 = {{9{1'b0}}, col_in_317};
assign u_ca_in_318 = {{9{1'b0}}, col_in_318};
assign u_ca_in_319 = {{9{1'b0}}, col_in_319};
assign u_ca_in_320 = {{9{1'b0}}, col_in_320};
assign u_ca_in_321 = {{9{1'b0}}, col_in_321};
assign u_ca_in_322 = {{9{1'b0}}, col_in_322};
assign u_ca_in_323 = {{9{1'b0}}, col_in_323};
assign u_ca_in_324 = {{9{1'b0}}, col_in_324};
assign u_ca_in_325 = {{9{1'b0}}, col_in_325};
assign u_ca_in_326 = {{9{1'b0}}, col_in_326};
assign u_ca_in_327 = {{9{1'b0}}, col_in_327};
assign u_ca_in_328 = {{9{1'b0}}, col_in_328};
assign u_ca_in_329 = {{9{1'b0}}, col_in_329};
assign u_ca_in_330 = {{9{1'b0}}, col_in_330};
assign u_ca_in_331 = {{9{1'b0}}, col_in_331};
assign u_ca_in_332 = {{9{1'b0}}, col_in_332};
assign u_ca_in_333 = {{9{1'b0}}, col_in_333};
assign u_ca_in_334 = {{9{1'b0}}, col_in_334};
assign u_ca_in_335 = {{9{1'b0}}, col_in_335};
assign u_ca_in_336 = {{9{1'b0}}, col_in_336};
assign u_ca_in_337 = {{9{1'b0}}, col_in_337};
assign u_ca_in_338 = {{9{1'b0}}, col_in_338};
assign u_ca_in_339 = {{9{1'b0}}, col_in_339};
assign u_ca_in_340 = {{9{1'b0}}, col_in_340};
assign u_ca_in_341 = {{9{1'b0}}, col_in_341};
assign u_ca_in_342 = {{9{1'b0}}, col_in_342};
assign u_ca_in_343 = {{9{1'b0}}, col_in_343};
assign u_ca_in_344 = {{9{1'b0}}, col_in_344};
assign u_ca_in_345 = {{9{1'b0}}, col_in_345};
assign u_ca_in_346 = {{9{1'b0}}, col_in_346};
assign u_ca_in_347 = {{9{1'b0}}, col_in_347};
assign u_ca_in_348 = {{9{1'b0}}, col_in_348};
assign u_ca_in_349 = {{9{1'b0}}, col_in_349};
assign u_ca_in_350 = {{9{1'b0}}, col_in_350};
assign u_ca_in_351 = {{9{1'b0}}, col_in_351};
assign u_ca_in_352 = {{9{1'b0}}, col_in_352};
assign u_ca_in_353 = {{9{1'b0}}, col_in_353};
assign u_ca_in_354 = {{9{1'b0}}, col_in_354};
assign u_ca_in_355 = {{9{1'b0}}, col_in_355};
assign u_ca_in_356 = {{9{1'b0}}, col_in_356};
assign u_ca_in_357 = {{9{1'b0}}, col_in_357};
assign u_ca_in_358 = {{9{1'b0}}, col_in_358};
assign u_ca_in_359 = {{9{1'b0}}, col_in_359};
assign u_ca_in_360 = {{9{1'b0}}, col_in_360};
assign u_ca_in_361 = {{9{1'b0}}, col_in_361};
assign u_ca_in_362 = {{9{1'b0}}, col_in_362};
assign u_ca_in_363 = {{9{1'b0}}, col_in_363};
assign u_ca_in_364 = {{9{1'b0}}, col_in_364};
assign u_ca_in_365 = {{9{1'b0}}, col_in_365};
assign u_ca_in_366 = {{9{1'b0}}, col_in_366};
assign u_ca_in_367 = {{9{1'b0}}, col_in_367};
assign u_ca_in_368 = {{9{1'b0}}, col_in_368};
assign u_ca_in_369 = {{9{1'b0}}, col_in_369};
assign u_ca_in_370 = {{9{1'b0}}, col_in_370};
assign u_ca_in_371 = {{9{1'b0}}, col_in_371};
assign u_ca_in_372 = {{9{1'b0}}, col_in_372};
assign u_ca_in_373 = {{9{1'b0}}, col_in_373};
assign u_ca_in_374 = {{9{1'b0}}, col_in_374};
assign u_ca_in_375 = {{9{1'b0}}, col_in_375};
assign u_ca_in_376 = {{9{1'b0}}, col_in_376};
assign u_ca_in_377 = {{9{1'b0}}, col_in_377};
assign u_ca_in_378 = {{9{1'b0}}, col_in_378};
assign u_ca_in_379 = {{9{1'b0}}, col_in_379};
assign u_ca_in_380 = {{9{1'b0}}, col_in_380};
assign u_ca_in_381 = {{9{1'b0}}, col_in_381};
assign u_ca_in_382 = {{9{1'b0}}, col_in_382};
assign u_ca_in_383 = {{9{1'b0}}, col_in_383};
assign u_ca_in_384 = {{9{1'b0}}, col_in_384};
assign u_ca_in_385 = {{9{1'b0}}, col_in_385};
assign u_ca_in_386 = {{9{1'b0}}, col_in_386};
assign u_ca_in_387 = {{9{1'b0}}, col_in_387};
assign u_ca_in_388 = {{9{1'b0}}, col_in_388};
assign u_ca_in_389 = {{9{1'b0}}, col_in_389};
assign u_ca_in_390 = {{9{1'b0}}, col_in_390};
assign u_ca_in_391 = {{9{1'b0}}, col_in_391};
assign u_ca_in_392 = {{9{1'b0}}, col_in_392};
assign u_ca_in_393 = {{9{1'b0}}, col_in_393};
assign u_ca_in_394 = {{9{1'b0}}, col_in_394};
assign u_ca_in_395 = {{9{1'b0}}, col_in_395};
assign u_ca_in_396 = {{9{1'b0}}, col_in_396};
assign u_ca_in_397 = {{9{1'b0}}, col_in_397};
assign u_ca_in_398 = {{9{1'b0}}, col_in_398};
assign u_ca_in_399 = {{9{1'b0}}, col_in_399};
assign u_ca_in_400 = {{9{1'b0}}, col_in_400};
assign u_ca_in_401 = {{9{1'b0}}, col_in_401};
assign u_ca_in_402 = {{9{1'b0}}, col_in_402};
assign u_ca_in_403 = {{9{1'b0}}, col_in_403};
assign u_ca_in_404 = {{9{1'b0}}, col_in_404};
assign u_ca_in_405 = {{9{1'b0}}, col_in_405};
assign u_ca_in_406 = {{9{1'b0}}, col_in_406};
assign u_ca_in_407 = {{9{1'b0}}, col_in_407};
assign u_ca_in_408 = {{9{1'b0}}, col_in_408};
assign u_ca_in_409 = {{9{1'b0}}, col_in_409};
assign u_ca_in_410 = {{9{1'b0}}, col_in_410};
assign u_ca_in_411 = {{9{1'b0}}, col_in_411};
assign u_ca_in_412 = {{9{1'b0}}, col_in_412};
assign u_ca_in_413 = {{9{1'b0}}, col_in_413};
assign u_ca_in_414 = {{9{1'b0}}, col_in_414};
assign u_ca_in_415 = {{9{1'b0}}, col_in_415};
assign u_ca_in_416 = {{9{1'b0}}, col_in_416};
assign u_ca_in_417 = {{9{1'b0}}, col_in_417};
assign u_ca_in_418 = {{9{1'b0}}, col_in_418};
assign u_ca_in_419 = {{9{1'b0}}, col_in_419};
assign u_ca_in_420 = {{9{1'b0}}, col_in_420};
assign u_ca_in_421 = {{9{1'b0}}, col_in_421};
assign u_ca_in_422 = {{9{1'b0}}, col_in_422};
assign u_ca_in_423 = {{9{1'b0}}, col_in_423};
assign u_ca_in_424 = {{9{1'b0}}, col_in_424};
assign u_ca_in_425 = {{9{1'b0}}, col_in_425};
assign u_ca_in_426 = {{9{1'b0}}, col_in_426};
assign u_ca_in_427 = {{9{1'b0}}, col_in_427};
assign u_ca_in_428 = {{9{1'b0}}, col_in_428};
assign u_ca_in_429 = {{9{1'b0}}, col_in_429};
assign u_ca_in_430 = {{9{1'b0}}, col_in_430};
assign u_ca_in_431 = {{9{1'b0}}, col_in_431};
assign u_ca_in_432 = {{9{1'b0}}, col_in_432};
assign u_ca_in_433 = {{9{1'b0}}, col_in_433};
assign u_ca_in_434 = {{9{1'b0}}, col_in_434};
assign u_ca_in_435 = {{9{1'b0}}, col_in_435};
assign u_ca_in_436 = {{9{1'b0}}, col_in_436};
assign u_ca_in_437 = {{9{1'b0}}, col_in_437};
assign u_ca_in_438 = {{9{1'b0}}, col_in_438};
assign u_ca_in_439 = {{9{1'b0}}, col_in_439};
assign u_ca_in_440 = {{9{1'b0}}, col_in_440};
assign u_ca_in_441 = {{9{1'b0}}, col_in_441};
assign u_ca_in_442 = {{9{1'b0}}, col_in_442};
assign u_ca_in_443 = {{9{1'b0}}, col_in_443};
assign u_ca_in_444 = {{9{1'b0}}, col_in_444};
assign u_ca_in_445 = {{9{1'b0}}, col_in_445};
assign u_ca_in_446 = {{9{1'b0}}, col_in_446};
assign u_ca_in_447 = {{9{1'b0}}, col_in_447};
assign u_ca_in_448 = {{9{1'b0}}, col_in_448};
assign u_ca_in_449 = {{9{1'b0}}, col_in_449};
assign u_ca_in_450 = {{9{1'b0}}, col_in_450};
assign u_ca_in_451 = {{9{1'b0}}, col_in_451};
assign u_ca_in_452 = {{9{1'b0}}, col_in_452};
assign u_ca_in_453 = {{9{1'b0}}, col_in_453};
assign u_ca_in_454 = {{9{1'b0}}, col_in_454};
assign u_ca_in_455 = {{9{1'b0}}, col_in_455};
assign u_ca_in_456 = {{9{1'b0}}, col_in_456};
assign u_ca_in_457 = {{9{1'b0}}, col_in_457};
assign u_ca_in_458 = {{9{1'b0}}, col_in_458};
assign u_ca_in_459 = {{9{1'b0}}, col_in_459};
assign u_ca_in_460 = {{9{1'b0}}, col_in_460};
assign u_ca_in_461 = {{9{1'b0}}, col_in_461};
assign u_ca_in_462 = {{9{1'b0}}, col_in_462};
assign u_ca_in_463 = {{9{1'b0}}, col_in_463};
assign u_ca_in_464 = {{9{1'b0}}, col_in_464};
assign u_ca_in_465 = {{9{1'b0}}, col_in_465};
assign u_ca_in_466 = {{9{1'b0}}, col_in_466};
assign u_ca_in_467 = {{9{1'b0}}, col_in_467};
assign u_ca_in_468 = {{9{1'b0}}, col_in_468};
assign u_ca_in_469 = {{9{1'b0}}, col_in_469};
assign u_ca_in_470 = {{9{1'b0}}, col_in_470};
assign u_ca_in_471 = {{9{1'b0}}, col_in_471};
assign u_ca_in_472 = {{9{1'b0}}, col_in_472};
assign u_ca_in_473 = {{9{1'b0}}, col_in_473};
assign u_ca_in_474 = {{9{1'b0}}, col_in_474};
assign u_ca_in_475 = {{9{1'b0}}, col_in_475};
assign u_ca_in_476 = {{9{1'b0}}, col_in_476};
assign u_ca_in_477 = {{9{1'b0}}, col_in_477};
assign u_ca_in_478 = {{9{1'b0}}, col_in_478};
assign u_ca_in_479 = {{9{1'b0}}, col_in_479};
assign u_ca_in_480 = {{9{1'b0}}, col_in_480};
assign u_ca_in_481 = {{9{1'b0}}, col_in_481};
assign u_ca_in_482 = {{9{1'b0}}, col_in_482};
assign u_ca_in_483 = {{9{1'b0}}, col_in_483};
assign u_ca_in_484 = {{9{1'b0}}, col_in_484};
assign u_ca_in_485 = {{9{1'b0}}, col_in_485};
assign u_ca_in_486 = {{9{1'b0}}, col_in_486};
assign u_ca_in_487 = {{9{1'b0}}, col_in_487};
assign u_ca_in_488 = {{9{1'b0}}, col_in_488};
assign u_ca_in_489 = {{9{1'b0}}, col_in_489};
assign u_ca_in_490 = {{9{1'b0}}, col_in_490};
assign u_ca_in_491 = {{9{1'b0}}, col_in_491};
assign u_ca_in_492 = {{9{1'b0}}, col_in_492};
assign u_ca_in_493 = {{9{1'b0}}, col_in_493};
assign u_ca_in_494 = {{9{1'b0}}, col_in_494};
assign u_ca_in_495 = {{9{1'b0}}, col_in_495};
assign u_ca_in_496 = {{9{1'b0}}, col_in_496};
assign u_ca_in_497 = {{9{1'b0}}, col_in_497};
assign u_ca_in_498 = {{9{1'b0}}, col_in_498};
assign u_ca_in_499 = {{9{1'b0}}, col_in_499};
assign u_ca_in_500 = {{9{1'b0}}, col_in_500};
assign u_ca_in_501 = {{9{1'b0}}, col_in_501};
assign u_ca_in_502 = {{9{1'b0}}, col_in_502};
assign u_ca_in_503 = {{9{1'b0}}, col_in_503};
assign u_ca_in_504 = {{9{1'b0}}, col_in_504};
assign u_ca_in_505 = {{9{1'b0}}, col_in_505};
assign u_ca_in_506 = {{9{1'b0}}, col_in_506};
assign u_ca_in_507 = {{9{1'b0}}, col_in_507};
assign u_ca_in_508 = {{9{1'b0}}, col_in_508};
assign u_ca_in_509 = {{9{1'b0}}, col_in_509};
assign u_ca_in_510 = {{9{1'b0}}, col_in_510};
assign u_ca_in_511 = {{9{1'b0}}, col_in_511};
assign u_ca_in_512 = {{9{1'b0}}, col_in_512};
assign u_ca_in_513 = {{9{1'b0}}, col_in_513};
assign u_ca_in_514 = {{9{1'b0}}, col_in_514};
assign u_ca_in_515 = {{9{1'b0}}, col_in_515};
assign u_ca_in_516 = {{9{1'b0}}, col_in_516};
assign u_ca_in_517 = {{9{1'b0}}, col_in_517};
assign u_ca_in_518 = {{9{1'b0}}, col_in_518};
assign u_ca_in_519 = {{9{1'b0}}, col_in_519};
assign u_ca_in_520 = {{9{1'b0}}, col_in_520};
assign u_ca_in_521 = {{9{1'b0}}, col_in_521};
assign u_ca_in_522 = {{9{1'b0}}, col_in_522};
assign u_ca_in_523 = {{9{1'b0}}, col_in_523};
assign u_ca_in_524 = {{9{1'b0}}, col_in_524};
assign u_ca_in_525 = {{9{1'b0}}, col_in_525};
assign u_ca_in_526 = {{9{1'b0}}, col_in_526};
assign u_ca_in_527 = {{9{1'b0}}, col_in_527};
assign u_ca_in_528 = {{9{1'b0}}, col_in_528};
assign u_ca_in_529 = {{9{1'b0}}, col_in_529};
assign u_ca_in_530 = {{9{1'b0}}, col_in_530};
assign u_ca_in_531 = {{9{1'b0}}, col_in_531};
assign u_ca_in_532 = {{9{1'b0}}, col_in_532};
assign u_ca_in_533 = {{9{1'b0}}, col_in_533};
assign u_ca_in_534 = {{9{1'b0}}, col_in_534};
assign u_ca_in_535 = {{9{1'b0}}, col_in_535};
assign u_ca_in_536 = {{9{1'b0}}, col_in_536};
assign u_ca_in_537 = {{9{1'b0}}, col_in_537};
assign u_ca_in_538 = {{9{1'b0}}, col_in_538};
assign u_ca_in_539 = {{9{1'b0}}, col_in_539};
assign u_ca_in_540 = {{9{1'b0}}, col_in_540};
assign u_ca_in_541 = {{9{1'b0}}, col_in_541};
assign u_ca_in_542 = {{9{1'b0}}, col_in_542};
assign u_ca_in_543 = {{9{1'b0}}, col_in_543};
assign u_ca_in_544 = {{9{1'b0}}, col_in_544};
assign u_ca_in_545 = {{9{1'b0}}, col_in_545};
assign u_ca_in_546 = {{9{1'b0}}, col_in_546};
assign u_ca_in_547 = {{9{1'b0}}, col_in_547};
assign u_ca_in_548 = {{9{1'b0}}, col_in_548};
assign u_ca_in_549 = {{9{1'b0}}, col_in_549};
assign u_ca_in_550 = {{9{1'b0}}, col_in_550};
assign u_ca_in_551 = {{9{1'b0}}, col_in_551};
assign u_ca_in_552 = {{9{1'b0}}, col_in_552};
assign u_ca_in_553 = {{9{1'b0}}, col_in_553};
assign u_ca_in_554 = {{9{1'b0}}, col_in_554};
assign u_ca_in_555 = {{9{1'b0}}, col_in_555};
assign u_ca_in_556 = {{9{1'b0}}, col_in_556};
assign u_ca_in_557 = {{9{1'b0}}, col_in_557};
assign u_ca_in_558 = {{9{1'b0}}, col_in_558};
assign u_ca_in_559 = {{9{1'b0}}, col_in_559};
assign u_ca_in_560 = {{9{1'b0}}, col_in_560};
assign u_ca_in_561 = {{9{1'b0}}, col_in_561};
assign u_ca_in_562 = {{9{1'b0}}, col_in_562};
assign u_ca_in_563 = {{9{1'b0}}, col_in_563};
assign u_ca_in_564 = {{9{1'b0}}, col_in_564};
assign u_ca_in_565 = {{9{1'b0}}, col_in_565};
assign u_ca_in_566 = {{9{1'b0}}, col_in_566};
assign u_ca_in_567 = {{9{1'b0}}, col_in_567};
assign u_ca_in_568 = {{9{1'b0}}, col_in_568};
assign u_ca_in_569 = {{9{1'b0}}, col_in_569};
assign u_ca_in_570 = {{9{1'b0}}, col_in_570};
assign u_ca_in_571 = {{9{1'b0}}, col_in_571};
assign u_ca_in_572 = {{9{1'b0}}, col_in_572};
assign u_ca_in_573 = {{9{1'b0}}, col_in_573};
assign u_ca_in_574 = {{9{1'b0}}, col_in_574};
assign u_ca_in_575 = {{9{1'b0}}, col_in_575};
assign u_ca_in_576 = {{9{1'b0}}, col_in_576};
assign u_ca_in_577 = {{9{1'b0}}, col_in_577};
assign u_ca_in_578 = {{9{1'b0}}, col_in_578};
assign u_ca_in_579 = {{9{1'b0}}, col_in_579};
assign u_ca_in_580 = {{9{1'b0}}, col_in_580};
assign u_ca_in_581 = {{9{1'b0}}, col_in_581};
assign u_ca_in_582 = {{9{1'b0}}, col_in_582};
assign u_ca_in_583 = {{9{1'b0}}, col_in_583};
assign u_ca_in_584 = {{9{1'b0}}, col_in_584};
assign u_ca_in_585 = {{9{1'b0}}, col_in_585};
assign u_ca_in_586 = {{9{1'b0}}, col_in_586};
assign u_ca_in_587 = {{9{1'b0}}, col_in_587};
assign u_ca_in_588 = {{9{1'b0}}, col_in_588};
assign u_ca_in_589 = {{9{1'b0}}, col_in_589};
assign u_ca_in_590 = {{9{1'b0}}, col_in_590};
assign u_ca_in_591 = {{9{1'b0}}, col_in_591};
assign u_ca_in_592 = {{9{1'b0}}, col_in_592};
assign u_ca_in_593 = {{9{1'b0}}, col_in_593};
assign u_ca_in_594 = {{9{1'b0}}, col_in_594};
assign u_ca_in_595 = {{9{1'b0}}, col_in_595};
assign u_ca_in_596 = {{9{1'b0}}, col_in_596};
assign u_ca_in_597 = {{9{1'b0}}, col_in_597};
assign u_ca_in_598 = {{9{1'b0}}, col_in_598};
assign u_ca_in_599 = {{9{1'b0}}, col_in_599};
assign u_ca_in_600 = {{9{1'b0}}, col_in_600};
assign u_ca_in_601 = {{9{1'b0}}, col_in_601};
assign u_ca_in_602 = {{9{1'b0}}, col_in_602};
assign u_ca_in_603 = {{9{1'b0}}, col_in_603};
assign u_ca_in_604 = {{9{1'b0}}, col_in_604};
assign u_ca_in_605 = {{9{1'b0}}, col_in_605};
assign u_ca_in_606 = {{9{1'b0}}, col_in_606};
assign u_ca_in_607 = {{9{1'b0}}, col_in_607};
assign u_ca_in_608 = {{9{1'b0}}, col_in_608};
assign u_ca_in_609 = {{9{1'b0}}, col_in_609};
assign u_ca_in_610 = {{9{1'b0}}, col_in_610};
assign u_ca_in_611 = {{9{1'b0}}, col_in_611};
assign u_ca_in_612 = {{9{1'b0}}, col_in_612};
assign u_ca_in_613 = {{9{1'b0}}, col_in_613};
assign u_ca_in_614 = {{9{1'b0}}, col_in_614};
assign u_ca_in_615 = {{9{1'b0}}, col_in_615};
assign u_ca_in_616 = {{9{1'b0}}, col_in_616};
assign u_ca_in_617 = {{9{1'b0}}, col_in_617};
assign u_ca_in_618 = {{9{1'b0}}, col_in_618};
assign u_ca_in_619 = {{9{1'b0}}, col_in_619};
assign u_ca_in_620 = {{9{1'b0}}, col_in_620};
assign u_ca_in_621 = {{9{1'b0}}, col_in_621};
assign u_ca_in_622 = {{9{1'b0}}, col_in_622};
assign u_ca_in_623 = {{9{1'b0}}, col_in_623};
assign u_ca_in_624 = {{9{1'b0}}, col_in_624};
assign u_ca_in_625 = {{9{1'b0}}, col_in_625};
assign u_ca_in_626 = {{9{1'b0}}, col_in_626};
assign u_ca_in_627 = {{9{1'b0}}, col_in_627};
assign u_ca_in_628 = {{9{1'b0}}, col_in_628};
assign u_ca_in_629 = {{9{1'b0}}, col_in_629};
assign u_ca_in_630 = {{9{1'b0}}, col_in_630};
assign u_ca_in_631 = {{9{1'b0}}, col_in_631};
assign u_ca_in_632 = {{9{1'b0}}, col_in_632};
assign u_ca_in_633 = {{9{1'b0}}, col_in_633};
assign u_ca_in_634 = {{9{1'b0}}, col_in_634};
assign u_ca_in_635 = {{9{1'b0}}, col_in_635};
assign u_ca_in_636 = {{9{1'b0}}, col_in_636};
assign u_ca_in_637 = {{9{1'b0}}, col_in_637};
assign u_ca_in_638 = {{9{1'b0}}, col_in_638};
assign u_ca_in_639 = {{9{1'b0}}, col_in_639};
assign u_ca_in_640 = {{9{1'b0}}, col_in_640};
assign u_ca_in_641 = {{9{1'b0}}, col_in_641};
assign u_ca_in_642 = {{9{1'b0}}, col_in_642};
assign u_ca_in_643 = {{9{1'b0}}, col_in_643};
assign u_ca_in_644 = {{9{1'b0}}, col_in_644};
assign u_ca_in_645 = {{9{1'b0}}, col_in_645};
assign u_ca_in_646 = {{9{1'b0}}, col_in_646};
assign u_ca_in_647 = {{9{1'b0}}, col_in_647};
assign u_ca_in_648 = {{9{1'b0}}, col_in_648};
assign u_ca_in_649 = {{9{1'b0}}, col_in_649};
assign u_ca_in_650 = {{9{1'b0}}, col_in_650};
assign u_ca_in_651 = {{9{1'b0}}, col_in_651};
assign u_ca_in_652 = {{9{1'b0}}, col_in_652};
assign u_ca_in_653 = {{9{1'b0}}, col_in_653};
assign u_ca_in_654 = {{9{1'b0}}, col_in_654};
assign u_ca_in_655 = {{9{1'b0}}, col_in_655};
assign u_ca_in_656 = {{9{1'b0}}, col_in_656};
assign u_ca_in_657 = {{9{1'b0}}, col_in_657};
assign u_ca_in_658 = {{9{1'b0}}, col_in_658};
assign u_ca_in_659 = {{9{1'b0}}, col_in_659};
assign u_ca_in_660 = {{9{1'b0}}, col_in_660};
assign u_ca_in_661 = {{9{1'b0}}, col_in_661};
assign u_ca_in_662 = {{9{1'b0}}, col_in_662};
assign u_ca_in_663 = {{9{1'b0}}, col_in_663};
assign u_ca_in_664 = {{9{1'b0}}, col_in_664};
assign u_ca_in_665 = {{9{1'b0}}, col_in_665};
assign u_ca_in_666 = {{9{1'b0}}, col_in_666};
assign u_ca_in_667 = {{9{1'b0}}, col_in_667};
assign u_ca_in_668 = {{9{1'b0}}, col_in_668};
assign u_ca_in_669 = {{9{1'b0}}, col_in_669};
assign u_ca_in_670 = {{9{1'b0}}, col_in_670};
assign u_ca_in_671 = {{9{1'b0}}, col_in_671};
assign u_ca_in_672 = {{9{1'b0}}, col_in_672};
assign u_ca_in_673 = {{9{1'b0}}, col_in_673};
assign u_ca_in_674 = {{9{1'b0}}, col_in_674};
assign u_ca_in_675 = {{9{1'b0}}, col_in_675};
assign u_ca_in_676 = {{9{1'b0}}, col_in_676};
assign u_ca_in_677 = {{9{1'b0}}, col_in_677};
assign u_ca_in_678 = {{9{1'b0}}, col_in_678};
assign u_ca_in_679 = {{9{1'b0}}, col_in_679};
assign u_ca_in_680 = {{9{1'b0}}, col_in_680};
assign u_ca_in_681 = {{9{1'b0}}, col_in_681};
assign u_ca_in_682 = {{9{1'b0}}, col_in_682};
assign u_ca_in_683 = {{9{1'b0}}, col_in_683};
assign u_ca_in_684 = {{9{1'b0}}, col_in_684};
assign u_ca_in_685 = {{9{1'b0}}, col_in_685};
assign u_ca_in_686 = {{9{1'b0}}, col_in_686};
assign u_ca_in_687 = {{9{1'b0}}, col_in_687};
assign u_ca_in_688 = {{9{1'b0}}, col_in_688};
assign u_ca_in_689 = {{9{1'b0}}, col_in_689};
assign u_ca_in_690 = {{9{1'b0}}, col_in_690};
assign u_ca_in_691 = {{9{1'b0}}, col_in_691};
assign u_ca_in_692 = {{9{1'b0}}, col_in_692};
assign u_ca_in_693 = {{9{1'b0}}, col_in_693};
assign u_ca_in_694 = {{9{1'b0}}, col_in_694};
assign u_ca_in_695 = {{9{1'b0}}, col_in_695};
assign u_ca_in_696 = {{9{1'b0}}, col_in_696};
assign u_ca_in_697 = {{9{1'b0}}, col_in_697};
assign u_ca_in_698 = {{9{1'b0}}, col_in_698};
assign u_ca_in_699 = {{9{1'b0}}, col_in_699};
assign u_ca_in_700 = {{9{1'b0}}, col_in_700};
assign u_ca_in_701 = {{9{1'b0}}, col_in_701};
assign u_ca_in_702 = {{9{1'b0}}, col_in_702};
assign u_ca_in_703 = {{9{1'b0}}, col_in_703};
assign u_ca_in_704 = {{9{1'b0}}, col_in_704};
assign u_ca_in_705 = {{9{1'b0}}, col_in_705};
assign u_ca_in_706 = {{9{1'b0}}, col_in_706};
assign u_ca_in_707 = {{9{1'b0}}, col_in_707};
assign u_ca_in_708 = {{9{1'b0}}, col_in_708};
assign u_ca_in_709 = {{9{1'b0}}, col_in_709};
assign u_ca_in_710 = {{9{1'b0}}, col_in_710};
assign u_ca_in_711 = {{9{1'b0}}, col_in_711};
assign u_ca_in_712 = {{9{1'b0}}, col_in_712};
assign u_ca_in_713 = {{9{1'b0}}, col_in_713};
assign u_ca_in_714 = {{9{1'b0}}, col_in_714};
assign u_ca_in_715 = {{9{1'b0}}, col_in_715};
assign u_ca_in_716 = {{9{1'b0}}, col_in_716};
assign u_ca_in_717 = {{9{1'b0}}, col_in_717};
assign u_ca_in_718 = {{9{1'b0}}, col_in_718};
assign u_ca_in_719 = {{9{1'b0}}, col_in_719};
assign u_ca_in_720 = {{9{1'b0}}, col_in_720};
assign u_ca_in_721 = {{9{1'b0}}, col_in_721};
assign u_ca_in_722 = {{9{1'b0}}, col_in_722};
assign u_ca_in_723 = {{9{1'b0}}, col_in_723};
assign u_ca_in_724 = {{9{1'b0}}, col_in_724};
assign u_ca_in_725 = {{9{1'b0}}, col_in_725};
assign u_ca_in_726 = {{9{1'b0}}, col_in_726};
assign u_ca_in_727 = {{9{1'b0}}, col_in_727};
assign u_ca_in_728 = {{9{1'b0}}, col_in_728};
assign u_ca_in_729 = {{9{1'b0}}, col_in_729};
assign u_ca_in_730 = {{9{1'b0}}, col_in_730};
assign u_ca_in_731 = {{9{1'b0}}, col_in_731};
assign u_ca_in_732 = {{9{1'b0}}, col_in_732};
assign u_ca_in_733 = {{9{1'b0}}, col_in_733};
assign u_ca_in_734 = {{9{1'b0}}, col_in_734};
assign u_ca_in_735 = {{9{1'b0}}, col_in_735};
assign u_ca_in_736 = {{9{1'b0}}, col_in_736};
assign u_ca_in_737 = {{9{1'b0}}, col_in_737};
assign u_ca_in_738 = {{9{1'b0}}, col_in_738};
assign u_ca_in_739 = {{9{1'b0}}, col_in_739};
assign u_ca_in_740 = {{9{1'b0}}, col_in_740};
assign u_ca_in_741 = {{9{1'b0}}, col_in_741};
assign u_ca_in_742 = {{9{1'b0}}, col_in_742};
assign u_ca_in_743 = {{9{1'b0}}, col_in_743};
assign u_ca_in_744 = {{9{1'b0}}, col_in_744};
assign u_ca_in_745 = {{9{1'b0}}, col_in_745};
assign u_ca_in_746 = {{9{1'b0}}, col_in_746};
assign u_ca_in_747 = {{9{1'b0}}, col_in_747};
assign u_ca_in_748 = {{9{1'b0}}, col_in_748};
assign u_ca_in_749 = {{9{1'b0}}, col_in_749};
assign u_ca_in_750 = {{9{1'b0}}, col_in_750};
assign u_ca_in_751 = {{9{1'b0}}, col_in_751};
assign u_ca_in_752 = {{9{1'b0}}, col_in_752};
assign u_ca_in_753 = {{9{1'b0}}, col_in_753};
assign u_ca_in_754 = {{9{1'b0}}, col_in_754};
assign u_ca_in_755 = {{9{1'b0}}, col_in_755};
assign u_ca_in_756 = {{9{1'b0}}, col_in_756};
assign u_ca_in_757 = {{9{1'b0}}, col_in_757};
assign u_ca_in_758 = {{9{1'b0}}, col_in_758};
assign u_ca_in_759 = {{9{1'b0}}, col_in_759};
assign u_ca_in_760 = {{9{1'b0}}, col_in_760};
assign u_ca_in_761 = {{9{1'b0}}, col_in_761};
assign u_ca_in_762 = {{9{1'b0}}, col_in_762};
assign u_ca_in_763 = {{9{1'b0}}, col_in_763};
assign u_ca_in_764 = {{9{1'b0}}, col_in_764};
assign u_ca_in_765 = {{9{1'b0}}, col_in_765};
assign u_ca_in_766 = {{9{1'b0}}, col_in_766};
assign u_ca_in_767 = {{9{1'b0}}, col_in_767};
assign u_ca_in_768 = {{9{1'b0}}, col_in_768};
assign u_ca_in_769 = {{9{1'b0}}, col_in_769};
assign u_ca_in_770 = {{9{1'b0}}, col_in_770};
assign u_ca_in_771 = {{9{1'b0}}, col_in_771};
assign u_ca_in_772 = {{9{1'b0}}, col_in_772};
assign u_ca_in_773 = {{9{1'b0}}, col_in_773};
assign u_ca_in_774 = {{9{1'b0}}, col_in_774};
assign u_ca_in_775 = {{9{1'b0}}, col_in_775};
assign u_ca_in_776 = {{9{1'b0}}, col_in_776};
assign u_ca_in_777 = {{9{1'b0}}, col_in_777};
assign u_ca_in_778 = {{9{1'b0}}, col_in_778};
assign u_ca_in_779 = {{9{1'b0}}, col_in_779};
assign u_ca_in_780 = {{9{1'b0}}, col_in_780};
assign u_ca_in_781 = {{9{1'b0}}, col_in_781};
assign u_ca_in_782 = {{9{1'b0}}, col_in_782};
assign u_ca_in_783 = {{9{1'b0}}, col_in_783};
assign u_ca_in_784 = {{9{1'b0}}, col_in_784};
assign u_ca_in_785 = {{9{1'b0}}, col_in_785};
assign u_ca_in_786 = {{9{1'b0}}, col_in_786};
assign u_ca_in_787 = {{9{1'b0}}, col_in_787};
assign u_ca_in_788 = {{9{1'b0}}, col_in_788};
assign u_ca_in_789 = {{9{1'b0}}, col_in_789};
assign u_ca_in_790 = {{9{1'b0}}, col_in_790};
assign u_ca_in_791 = {{9{1'b0}}, col_in_791};
assign u_ca_in_792 = {{9{1'b0}}, col_in_792};
assign u_ca_in_793 = {{9{1'b0}}, col_in_793};
assign u_ca_in_794 = {{9{1'b0}}, col_in_794};
assign u_ca_in_795 = {{9{1'b0}}, col_in_795};
assign u_ca_in_796 = {{9{1'b0}}, col_in_796};
assign u_ca_in_797 = {{9{1'b0}}, col_in_797};
assign u_ca_in_798 = {{9{1'b0}}, col_in_798};
assign u_ca_in_799 = {{9{1'b0}}, col_in_799};
assign u_ca_in_800 = {{9{1'b0}}, col_in_800};
assign u_ca_in_801 = {{9{1'b0}}, col_in_801};
assign u_ca_in_802 = {{9{1'b0}}, col_in_802};
assign u_ca_in_803 = {{9{1'b0}}, col_in_803};
assign u_ca_in_804 = {{9{1'b0}}, col_in_804};
assign u_ca_in_805 = {{9{1'b0}}, col_in_805};
assign u_ca_in_806 = {{9{1'b0}}, col_in_806};
assign u_ca_in_807 = {{9{1'b0}}, col_in_807};
assign u_ca_in_808 = {{9{1'b0}}, col_in_808};
assign u_ca_in_809 = {{9{1'b0}}, col_in_809};
assign u_ca_in_810 = {{9{1'b0}}, col_in_810};
assign u_ca_in_811 = {{9{1'b0}}, col_in_811};
assign u_ca_in_812 = {{9{1'b0}}, col_in_812};
assign u_ca_in_813 = {{9{1'b0}}, col_in_813};
assign u_ca_in_814 = {{9{1'b0}}, col_in_814};
assign u_ca_in_815 = {{9{1'b0}}, col_in_815};
assign u_ca_in_816 = {{9{1'b0}}, col_in_816};
assign u_ca_in_817 = {{9{1'b0}}, col_in_817};
assign u_ca_in_818 = {{9{1'b0}}, col_in_818};
assign u_ca_in_819 = {{9{1'b0}}, col_in_819};
assign u_ca_in_820 = {{9{1'b0}}, col_in_820};
assign u_ca_in_821 = {{9{1'b0}}, col_in_821};
assign u_ca_in_822 = {{9{1'b0}}, col_in_822};
assign u_ca_in_823 = {{9{1'b0}}, col_in_823};
assign u_ca_in_824 = {{9{1'b0}}, col_in_824};
assign u_ca_in_825 = {{9{1'b0}}, col_in_825};
assign u_ca_in_826 = {{9{1'b0}}, col_in_826};
assign u_ca_in_827 = {{9{1'b0}}, col_in_827};
assign u_ca_in_828 = {{9{1'b0}}, col_in_828};
assign u_ca_in_829 = {{9{1'b0}}, col_in_829};
assign u_ca_in_830 = {{9{1'b0}}, col_in_830};
assign u_ca_in_831 = {{9{1'b0}}, col_in_831};
assign u_ca_in_832 = {{9{1'b0}}, col_in_832};
assign u_ca_in_833 = {{9{1'b0}}, col_in_833};
assign u_ca_in_834 = {{9{1'b0}}, col_in_834};
assign u_ca_in_835 = {{9{1'b0}}, col_in_835};
assign u_ca_in_836 = {{9{1'b0}}, col_in_836};
assign u_ca_in_837 = {{9{1'b0}}, col_in_837};
assign u_ca_in_838 = {{9{1'b0}}, col_in_838};
assign u_ca_in_839 = {{9{1'b0}}, col_in_839};
assign u_ca_in_840 = {{9{1'b0}}, col_in_840};
assign u_ca_in_841 = {{9{1'b0}}, col_in_841};
assign u_ca_in_842 = {{9{1'b0}}, col_in_842};
assign u_ca_in_843 = {{9{1'b0}}, col_in_843};
assign u_ca_in_844 = {{9{1'b0}}, col_in_844};
assign u_ca_in_845 = {{9{1'b0}}, col_in_845};
assign u_ca_in_846 = {{9{1'b0}}, col_in_846};
assign u_ca_in_847 = {{9{1'b0}}, col_in_847};
assign u_ca_in_848 = {{9{1'b0}}, col_in_848};
assign u_ca_in_849 = {{9{1'b0}}, col_in_849};
assign u_ca_in_850 = {{9{1'b0}}, col_in_850};
assign u_ca_in_851 = {{9{1'b0}}, col_in_851};
assign u_ca_in_852 = {{9{1'b0}}, col_in_852};
assign u_ca_in_853 = {{9{1'b0}}, col_in_853};
assign u_ca_in_854 = {{9{1'b0}}, col_in_854};
assign u_ca_in_855 = {{9{1'b0}}, col_in_855};
assign u_ca_in_856 = {{9{1'b0}}, col_in_856};
assign u_ca_in_857 = {{9{1'b0}}, col_in_857};
assign u_ca_in_858 = {{9{1'b0}}, col_in_858};
assign u_ca_in_859 = {{9{1'b0}}, col_in_859};
assign u_ca_in_860 = {{9{1'b0}}, col_in_860};
assign u_ca_in_861 = {{9{1'b0}}, col_in_861};
assign u_ca_in_862 = {{9{1'b0}}, col_in_862};
assign u_ca_in_863 = {{9{1'b0}}, col_in_863};
assign u_ca_in_864 = {{9{1'b0}}, col_in_864};
assign u_ca_in_865 = {{9{1'b0}}, col_in_865};
assign u_ca_in_866 = {{9{1'b0}}, col_in_866};
assign u_ca_in_867 = {{9{1'b0}}, col_in_867};
assign u_ca_in_868 = {{9{1'b0}}, col_in_868};
assign u_ca_in_869 = {{9{1'b0}}, col_in_869};
assign u_ca_in_870 = {{9{1'b0}}, col_in_870};
assign u_ca_in_871 = {{9{1'b0}}, col_in_871};
assign u_ca_in_872 = {{9{1'b0}}, col_in_872};
assign u_ca_in_873 = {{9{1'b0}}, col_in_873};
assign u_ca_in_874 = {{9{1'b0}}, col_in_874};
assign u_ca_in_875 = {{9{1'b0}}, col_in_875};
assign u_ca_in_876 = {{9{1'b0}}, col_in_876};
assign u_ca_in_877 = {{9{1'b0}}, col_in_877};
assign u_ca_in_878 = {{9{1'b0}}, col_in_878};
assign u_ca_in_879 = {{9{1'b0}}, col_in_879};
assign u_ca_in_880 = {{9{1'b0}}, col_in_880};
assign u_ca_in_881 = {{9{1'b0}}, col_in_881};
assign u_ca_in_882 = {{9{1'b0}}, col_in_882};
assign u_ca_in_883 = {{9{1'b0}}, col_in_883};
assign u_ca_in_884 = {{9{1'b0}}, col_in_884};
assign u_ca_in_885 = {{9{1'b0}}, col_in_885};
assign u_ca_in_886 = {{9{1'b0}}, col_in_886};
assign u_ca_in_887 = {{9{1'b0}}, col_in_887};
assign u_ca_in_888 = {{9{1'b0}}, col_in_888};
assign u_ca_in_889 = {{9{1'b0}}, col_in_889};
assign u_ca_in_890 = {{9{1'b0}}, col_in_890};
assign u_ca_in_891 = {{9{1'b0}}, col_in_891};
assign u_ca_in_892 = {{9{1'b0}}, col_in_892};
assign u_ca_in_893 = {{9{1'b0}}, col_in_893};
assign u_ca_in_894 = {{9{1'b0}}, col_in_894};
assign u_ca_in_895 = {{9{1'b0}}, col_in_895};
assign u_ca_in_896 = {{9{1'b0}}, col_in_896};
assign u_ca_in_897 = {{9{1'b0}}, col_in_897};
assign u_ca_in_898 = {{9{1'b0}}, col_in_898};
assign u_ca_in_899 = {{9{1'b0}}, col_in_899};
assign u_ca_in_900 = {{9{1'b0}}, col_in_900};
assign u_ca_in_901 = {{9{1'b0}}, col_in_901};
assign u_ca_in_902 = {{9{1'b0}}, col_in_902};
assign u_ca_in_903 = {{9{1'b0}}, col_in_903};
assign u_ca_in_904 = {{9{1'b0}}, col_in_904};
assign u_ca_in_905 = {{9{1'b0}}, col_in_905};
assign u_ca_in_906 = {{9{1'b0}}, col_in_906};
assign u_ca_in_907 = {{9{1'b0}}, col_in_907};
assign u_ca_in_908 = {{9{1'b0}}, col_in_908};
assign u_ca_in_909 = {{9{1'b0}}, col_in_909};
assign u_ca_in_910 = {{9{1'b0}}, col_in_910};
assign u_ca_in_911 = {{9{1'b0}}, col_in_911};
assign u_ca_in_912 = {{9{1'b0}}, col_in_912};
assign u_ca_in_913 = {{9{1'b0}}, col_in_913};
assign u_ca_in_914 = {{9{1'b0}}, col_in_914};
assign u_ca_in_915 = {{9{1'b0}}, col_in_915};
assign u_ca_in_916 = {{9{1'b0}}, col_in_916};
assign u_ca_in_917 = {{9{1'b0}}, col_in_917};
assign u_ca_in_918 = {{9{1'b0}}, col_in_918};
assign u_ca_in_919 = {{9{1'b0}}, col_in_919};
assign u_ca_in_920 = {{9{1'b0}}, col_in_920};
assign u_ca_in_921 = {{9{1'b0}}, col_in_921};
assign u_ca_in_922 = {{9{1'b0}}, col_in_922};
assign u_ca_in_923 = {{9{1'b0}}, col_in_923};
assign u_ca_in_924 = {{9{1'b0}}, col_in_924};
assign u_ca_in_925 = {{9{1'b0}}, col_in_925};
assign u_ca_in_926 = {{9{1'b0}}, col_in_926};
assign u_ca_in_927 = {{9{1'b0}}, col_in_927};
assign u_ca_in_928 = {{9{1'b0}}, col_in_928};
assign u_ca_in_929 = {{9{1'b0}}, col_in_929};
assign u_ca_in_930 = {{9{1'b0}}, col_in_930};
assign u_ca_in_931 = {{9{1'b0}}, col_in_931};
assign u_ca_in_932 = {{9{1'b0}}, col_in_932};
assign u_ca_in_933 = {{9{1'b0}}, col_in_933};
assign u_ca_in_934 = {{9{1'b0}}, col_in_934};
assign u_ca_in_935 = {{9{1'b0}}, col_in_935};
assign u_ca_in_936 = {{9{1'b0}}, col_in_936};
assign u_ca_in_937 = {{9{1'b0}}, col_in_937};
assign u_ca_in_938 = {{9{1'b0}}, col_in_938};
assign u_ca_in_939 = {{9{1'b0}}, col_in_939};
assign u_ca_in_940 = {{9{1'b0}}, col_in_940};
assign u_ca_in_941 = {{9{1'b0}}, col_in_941};
assign u_ca_in_942 = {{9{1'b0}}, col_in_942};
assign u_ca_in_943 = {{9{1'b0}}, col_in_943};
assign u_ca_in_944 = {{9{1'b0}}, col_in_944};
assign u_ca_in_945 = {{9{1'b0}}, col_in_945};
assign u_ca_in_946 = {{9{1'b0}}, col_in_946};
assign u_ca_in_947 = {{9{1'b0}}, col_in_947};
assign u_ca_in_948 = {{9{1'b0}}, col_in_948};
assign u_ca_in_949 = {{9{1'b0}}, col_in_949};
assign u_ca_in_950 = {{9{1'b0}}, col_in_950};
assign u_ca_in_951 = {{9{1'b0}}, col_in_951};
assign u_ca_in_952 = {{9{1'b0}}, col_in_952};
assign u_ca_in_953 = {{9{1'b0}}, col_in_953};
assign u_ca_in_954 = {{9{1'b0}}, col_in_954};
assign u_ca_in_955 = {{9{1'b0}}, col_in_955};
assign u_ca_in_956 = {{9{1'b0}}, col_in_956};
assign u_ca_in_957 = {{9{1'b0}}, col_in_957};
assign u_ca_in_958 = {{9{1'b0}}, col_in_958};
assign u_ca_in_959 = {{9{1'b0}}, col_in_959};
assign u_ca_in_960 = {{9{1'b0}}, col_in_960};
assign u_ca_in_961 = {{9{1'b0}}, col_in_961};
assign u_ca_in_962 = {{9{1'b0}}, col_in_962};
assign u_ca_in_963 = {{9{1'b0}}, col_in_963};
assign u_ca_in_964 = {{9{1'b0}}, col_in_964};
assign u_ca_in_965 = {{9{1'b0}}, col_in_965};
assign u_ca_in_966 = {{9{1'b0}}, col_in_966};
assign u_ca_in_967 = {{9{1'b0}}, col_in_967};
assign u_ca_in_968 = {{9{1'b0}}, col_in_968};
assign u_ca_in_969 = {{9{1'b0}}, col_in_969};
assign u_ca_in_970 = {{9{1'b0}}, col_in_970};
assign u_ca_in_971 = {{9{1'b0}}, col_in_971};
assign u_ca_in_972 = {{9{1'b0}}, col_in_972};
assign u_ca_in_973 = {{9{1'b0}}, col_in_973};
assign u_ca_in_974 = {{9{1'b0}}, col_in_974};
assign u_ca_in_975 = {{9{1'b0}}, col_in_975};
assign u_ca_in_976 = {{9{1'b0}}, col_in_976};
assign u_ca_in_977 = {{9{1'b0}}, col_in_977};
assign u_ca_in_978 = {{9{1'b0}}, col_in_978};
assign u_ca_in_979 = {{9{1'b0}}, col_in_979};
assign u_ca_in_980 = {{9{1'b0}}, col_in_980};
assign u_ca_in_981 = {{9{1'b0}}, col_in_981};
assign u_ca_in_982 = {{9{1'b0}}, col_in_982};
assign u_ca_in_983 = {{9{1'b0}}, col_in_983};
assign u_ca_in_984 = {{9{1'b0}}, col_in_984};
assign u_ca_in_985 = {{9{1'b0}}, col_in_985};
assign u_ca_in_986 = {{9{1'b0}}, col_in_986};
assign u_ca_in_987 = {{9{1'b0}}, col_in_987};
assign u_ca_in_988 = {{9{1'b0}}, col_in_988};
assign u_ca_in_989 = {{9{1'b0}}, col_in_989};
assign u_ca_in_990 = {{9{1'b0}}, col_in_990};
assign u_ca_in_991 = {{9{1'b0}}, col_in_991};
assign u_ca_in_992 = {{9{1'b0}}, col_in_992};
assign u_ca_in_993 = {{9{1'b0}}, col_in_993};
assign u_ca_in_994 = {{9{1'b0}}, col_in_994};
assign u_ca_in_995 = {{9{1'b0}}, col_in_995};
assign u_ca_in_996 = {{9{1'b0}}, col_in_996};
assign u_ca_in_997 = {{9{1'b0}}, col_in_997};
assign u_ca_in_998 = {{9{1'b0}}, col_in_998};
assign u_ca_in_999 = {{9{1'b0}}, col_in_999};
assign u_ca_in_1000 = {{9{1'b0}}, col_in_1000};
assign u_ca_in_1001 = {{9{1'b0}}, col_in_1001};
assign u_ca_in_1002 = {{9{1'b0}}, col_in_1002};
assign u_ca_in_1003 = {{9{1'b0}}, col_in_1003};
assign u_ca_in_1004 = {{9{1'b0}}, col_in_1004};
assign u_ca_in_1005 = {{9{1'b0}}, col_in_1005};
assign u_ca_in_1006 = {{9{1'b0}}, col_in_1006};
assign u_ca_in_1007 = {{9{1'b0}}, col_in_1007};
assign u_ca_in_1008 = {{9{1'b0}}, col_in_1008};
assign u_ca_in_1009 = {{9{1'b0}}, col_in_1009};
assign u_ca_in_1010 = {{9{1'b0}}, col_in_1010};
assign u_ca_in_1011 = {{9{1'b0}}, col_in_1011};
assign u_ca_in_1012 = {{9{1'b0}}, col_in_1012};
assign u_ca_in_1013 = {{9{1'b0}}, col_in_1013};
assign u_ca_in_1014 = {{9{1'b0}}, col_in_1014};
assign u_ca_in_1015 = {{9{1'b0}}, col_in_1015};
assign u_ca_in_1016 = {{9{1'b0}}, col_in_1016};
assign u_ca_in_1017 = {{9{1'b0}}, col_in_1017};
assign u_ca_in_1018 = {{9{1'b0}}, col_in_1018};
assign u_ca_in_1019 = {{9{1'b0}}, col_in_1019};
assign u_ca_in_1020 = {{9{1'b0}}, col_in_1020};
assign u_ca_in_1021 = {{9{1'b0}}, col_in_1021};
assign u_ca_in_1022 = {{9{1'b0}}, col_in_1022};
assign u_ca_in_1023 = {{9{1'b0}}, col_in_1023};
assign u_ca_in_1024 = {{9{1'b0}}, col_in_1024};
assign u_ca_in_1025 = {{9{1'b0}}, col_in_1025};
assign u_ca_in_1026 = {{9{1'b0}}, col_in_1026};
assign u_ca_in_1027 = {{9{1'b0}}, col_in_1027};
assign u_ca_in_1028 = {{9{1'b0}}, col_in_1028};
assign u_ca_in_1029 = {{9{1'b0}}, col_in_1029};
assign u_ca_in_1030 = {{9{1'b0}}, col_in_1030};
assign u_ca_in_1031 = {{9{1'b0}}, col_in_1031};
assign u_ca_in_1032 = {{9{1'b0}}, col_in_1032};
assign u_ca_in_1033 = {{9{1'b0}}, col_in_1033};
assign u_ca_in_1034 = {{9{1'b0}}, col_in_1034};
assign u_ca_in_1035 = {{9{1'b0}}, col_in_1035};
assign u_ca_in_1036 = {{9{1'b0}}, col_in_1036};
assign u_ca_in_1037 = {{9{1'b0}}, col_in_1037};
assign u_ca_in_1038 = {{9{1'b0}}, col_in_1038};
assign u_ca_in_1039 = {{9{1'b0}}, col_in_1039};
assign u_ca_in_1040 = {{9{1'b0}}, col_in_1040};
assign u_ca_in_1041 = {{9{1'b0}}, col_in_1041};
assign u_ca_in_1042 = {{9{1'b0}}, col_in_1042};
assign u_ca_in_1043 = {{9{1'b0}}, col_in_1043};
assign u_ca_in_1044 = {{9{1'b0}}, col_in_1044};
assign u_ca_in_1045 = {{9{1'b0}}, col_in_1045};
assign u_ca_in_1046 = {{9{1'b0}}, col_in_1046};
assign u_ca_in_1047 = {{9{1'b0}}, col_in_1047};
assign u_ca_in_1048 = {{9{1'b0}}, col_in_1048};
assign u_ca_in_1049 = {{9{1'b0}}, col_in_1049};
assign u_ca_in_1050 = {{9{1'b0}}, col_in_1050};
assign u_ca_in_1051 = {{9{1'b0}}, col_in_1051};
assign u_ca_in_1052 = {{9{1'b0}}, col_in_1052};
assign u_ca_in_1053 = {{9{1'b0}}, col_in_1053};
assign u_ca_in_1054 = {{9{1'b0}}, col_in_1054};
assign u_ca_in_1055 = {{9{1'b0}}, col_in_1055};
assign u_ca_in_1056 = {{9{1'b0}}, col_in_1056};
assign u_ca_in_1057 = {{9{1'b0}}, col_in_1057};
assign u_ca_in_1058 = {{9{1'b0}}, col_in_1058};
assign u_ca_in_1059 = {{9{1'b0}}, col_in_1059};
assign u_ca_in_1060 = {{9{1'b0}}, col_in_1060};
assign u_ca_in_1061 = {{9{1'b0}}, col_in_1061};
assign u_ca_in_1062 = {{9{1'b0}}, col_in_1062};
assign u_ca_in_1063 = {{9{1'b0}}, col_in_1063};
assign u_ca_in_1064 = {{9{1'b0}}, col_in_1064};
assign u_ca_in_1065 = {{9{1'b0}}, col_in_1065};
assign u_ca_in_1066 = {{9{1'b0}}, col_in_1066};
assign u_ca_in_1067 = {{9{1'b0}}, col_in_1067};
assign u_ca_in_1068 = {{9{1'b0}}, col_in_1068};
assign u_ca_in_1069 = {{9{1'b0}}, col_in_1069};
assign u_ca_in_1070 = {{9{1'b0}}, col_in_1070};
assign u_ca_in_1071 = {{9{1'b0}}, col_in_1071};
assign u_ca_in_1072 = {{9{1'b0}}, col_in_1072};
assign u_ca_in_1073 = {{9{1'b0}}, col_in_1073};
assign u_ca_in_1074 = {{9{1'b0}}, col_in_1074};
assign u_ca_in_1075 = {{9{1'b0}}, col_in_1075};
assign u_ca_in_1076 = {{9{1'b0}}, col_in_1076};
assign u_ca_in_1077 = {{9{1'b0}}, col_in_1077};
assign u_ca_in_1078 = {{9{1'b0}}, col_in_1078};
assign u_ca_in_1079 = {{9{1'b0}}, col_in_1079};
assign u_ca_in_1080 = {{9{1'b0}}, col_in_1080};
assign u_ca_in_1081 = {{9{1'b0}}, col_in_1081};
assign u_ca_in_1082 = {{9{1'b0}}, col_in_1082};
assign u_ca_in_1083 = {{9{1'b0}}, col_in_1083};
assign u_ca_in_1084 = {{9{1'b0}}, col_in_1084};
assign u_ca_in_1085 = {{9{1'b0}}, col_in_1085};
assign u_ca_in_1086 = {{9{1'b0}}, col_in_1086};
assign u_ca_in_1087 = {{9{1'b0}}, col_in_1087};
assign u_ca_in_1088 = {{9{1'b0}}, col_in_1088};
assign u_ca_in_1089 = {{9{1'b0}}, col_in_1089};
assign u_ca_in_1090 = {{9{1'b0}}, col_in_1090};
assign u_ca_in_1091 = {{9{1'b0}}, col_in_1091};
assign u_ca_in_1092 = {{9{1'b0}}, col_in_1092};
assign u_ca_in_1093 = {{9{1'b0}}, col_in_1093};
assign u_ca_in_1094 = {{9{1'b0}}, col_in_1094};
assign u_ca_in_1095 = {{9{1'b0}}, col_in_1095};
assign u_ca_in_1096 = {{9{1'b0}}, col_in_1096};
assign u_ca_in_1097 = {{9{1'b0}}, col_in_1097};
assign u_ca_in_1098 = {{9{1'b0}}, col_in_1098};
assign u_ca_in_1099 = {{9{1'b0}}, col_in_1099};
assign u_ca_in_1100 = {{9{1'b0}}, col_in_1100};
assign u_ca_in_1101 = {{9{1'b0}}, col_in_1101};
assign u_ca_in_1102 = {{9{1'b0}}, col_in_1102};
assign u_ca_in_1103 = {{9{1'b0}}, col_in_1103};
assign u_ca_in_1104 = {{9{1'b0}}, col_in_1104};
assign u_ca_in_1105 = {{9{1'b0}}, col_in_1105};
assign u_ca_in_1106 = {{9{1'b0}}, col_in_1106};
assign u_ca_in_1107 = {{9{1'b0}}, col_in_1107};
assign u_ca_in_1108 = {{9{1'b0}}, col_in_1108};
assign u_ca_in_1109 = {{9{1'b0}}, col_in_1109};
assign u_ca_in_1110 = {{9{1'b0}}, col_in_1110};
assign u_ca_in_1111 = {{9{1'b0}}, col_in_1111};
assign u_ca_in_1112 = {{9{1'b0}}, col_in_1112};
assign u_ca_in_1113 = {{9{1'b0}}, col_in_1113};
assign u_ca_in_1114 = {{9{1'b0}}, col_in_1114};
assign u_ca_in_1115 = {{9{1'b0}}, col_in_1115};
assign u_ca_in_1116 = {{9{1'b0}}, col_in_1116};
assign u_ca_in_1117 = {{9{1'b0}}, col_in_1117};
assign u_ca_in_1118 = {{9{1'b0}}, col_in_1118};
assign u_ca_in_1119 = {{9{1'b0}}, col_in_1119};
assign u_ca_in_1120 = {{9{1'b0}}, col_in_1120};
assign u_ca_in_1121 = {{9{1'b0}}, col_in_1121};
assign u_ca_in_1122 = {{9{1'b0}}, col_in_1122};
assign u_ca_in_1123 = {{9{1'b0}}, col_in_1123};
assign u_ca_in_1124 = {{9{1'b0}}, col_in_1124};
assign u_ca_in_1125 = {{9{1'b0}}, col_in_1125};
assign u_ca_in_1126 = {{9{1'b0}}, col_in_1126};
assign u_ca_in_1127 = {{9{1'b0}}, col_in_1127};
assign u_ca_in_1128 = {{9{1'b0}}, col_in_1128};
assign u_ca_in_1129 = {{9{1'b0}}, col_in_1129};
assign u_ca_in_1130 = {{9{1'b0}}, col_in_1130};
assign u_ca_in_1131 = {{9{1'b0}}, col_in_1131};
assign u_ca_in_1132 = {{9{1'b0}}, col_in_1132};
assign u_ca_in_1133 = {{9{1'b0}}, col_in_1133};
assign u_ca_in_1134 = {{9{1'b0}}, col_in_1134};
assign u_ca_in_1135 = {{9{1'b0}}, col_in_1135};
assign u_ca_in_1136 = {{9{1'b0}}, col_in_1136};
assign u_ca_in_1137 = {{9{1'b0}}, col_in_1137};
assign u_ca_in_1138 = {{9{1'b0}}, col_in_1138};
assign u_ca_in_1139 = {{9{1'b0}}, col_in_1139};
assign u_ca_in_1140 = {{9{1'b0}}, col_in_1140};
assign u_ca_in_1141 = {{9{1'b0}}, col_in_1141};
assign u_ca_in_1142 = {{9{1'b0}}, col_in_1142};
assign u_ca_in_1143 = {{9{1'b0}}, col_in_1143};
assign u_ca_in_1144 = {{9{1'b0}}, col_in_1144};
assign u_ca_in_1145 = {{9{1'b0}}, col_in_1145};
assign u_ca_in_1146 = {{9{1'b0}}, col_in_1146};
assign u_ca_in_1147 = {{9{1'b0}}, col_in_1147};
assign u_ca_in_1148 = {{9{1'b0}}, col_in_1148};
assign u_ca_in_1149 = {{9{1'b0}}, col_in_1149};
assign u_ca_in_1150 = {{9{1'b0}}, col_in_1150};
assign u_ca_in_1151 = {{9{1'b0}}, col_in_1151};
assign u_ca_in_1152 = {{9{1'b0}}, col_in_1152};
assign u_ca_in_1153 = {{9{1'b0}}, col_in_1153};
assign u_ca_in_1154 = {{9{1'b0}}, col_in_1154};
assign u_ca_in_1155 = {{9{1'b0}}, col_in_1155};
assign u_ca_in_1156 = {{9{1'b0}}, col_in_1156};
assign u_ca_in_1157 = {{9{1'b0}}, col_in_1157};
assign u_ca_in_1158 = {{9{1'b0}}, col_in_1158};
assign u_ca_in_1159 = {{9{1'b0}}, col_in_1159};
assign u_ca_in_1160 = {{9{1'b0}}, col_in_1160};
assign u_ca_in_1161 = {{9{1'b0}}, col_in_1161};
assign u_ca_in_1162 = {{9{1'b0}}, col_in_1162};
assign u_ca_in_1163 = {{9{1'b0}}, col_in_1163};
assign u_ca_in_1164 = {{9{1'b0}}, col_in_1164};
assign u_ca_in_1165 = {{9{1'b0}}, col_in_1165};
assign u_ca_in_1166 = {{9{1'b0}}, col_in_1166};
assign u_ca_in_1167 = {{9{1'b0}}, col_in_1167};
assign u_ca_in_1168 = {{9{1'b0}}, col_in_1168};
assign u_ca_in_1169 = {{9{1'b0}}, col_in_1169};
assign u_ca_in_1170 = {{9{1'b0}}, col_in_1170};
assign u_ca_in_1171 = {{9{1'b0}}, col_in_1171};
assign u_ca_in_1172 = {{9{1'b0}}, col_in_1172};
assign u_ca_in_1173 = {{9{1'b0}}, col_in_1173};
assign u_ca_in_1174 = {{9{1'b0}}, col_in_1174};
assign u_ca_in_1175 = {{9{1'b0}}, col_in_1175};
assign u_ca_in_1176 = {{9{1'b0}}, col_in_1176};
assign u_ca_in_1177 = {{9{1'b0}}, col_in_1177};
assign u_ca_in_1178 = {{9{1'b0}}, col_in_1178};
assign u_ca_in_1179 = {{9{1'b0}}, col_in_1179};
assign u_ca_in_1180 = {{9{1'b0}}, col_in_1180};
assign u_ca_in_1181 = {{9{1'b0}}, col_in_1181};
assign u_ca_in_1182 = {{9{1'b0}}, col_in_1182};
assign u_ca_in_1183 = {{9{1'b0}}, col_in_1183};
assign u_ca_in_1184 = {{9{1'b0}}, col_in_1184};
assign u_ca_in_1185 = {{9{1'b0}}, col_in_1185};
assign u_ca_in_1186 = {{9{1'b0}}, col_in_1186};
assign u_ca_in_1187 = {{9{1'b0}}, col_in_1187};
assign u_ca_in_1188 = {{9{1'b0}}, col_in_1188};
assign u_ca_in_1189 = {{9{1'b0}}, col_in_1189};
assign u_ca_in_1190 = {{9{1'b0}}, col_in_1190};
assign u_ca_in_1191 = {{9{1'b0}}, col_in_1191};
assign u_ca_in_1192 = {{9{1'b0}}, col_in_1192};
assign u_ca_in_1193 = {{9{1'b0}}, col_in_1193};
assign u_ca_in_1194 = {{9{1'b0}}, col_in_1194};
assign u_ca_in_1195 = {{9{1'b0}}, col_in_1195};
assign u_ca_in_1196 = {{9{1'b0}}, col_in_1196};
assign u_ca_in_1197 = {{9{1'b0}}, col_in_1197};
assign u_ca_in_1198 = {{9{1'b0}}, col_in_1198};
assign u_ca_in_1199 = {{9{1'b0}}, col_in_1199};
assign u_ca_in_1200 = {{9{1'b0}}, col_in_1200};
assign u_ca_in_1201 = {{9{1'b0}}, col_in_1201};
assign u_ca_in_1202 = {{9{1'b0}}, col_in_1202};
assign u_ca_in_1203 = {{9{1'b0}}, col_in_1203};
assign u_ca_in_1204 = {{9{1'b0}}, col_in_1204};
assign u_ca_in_1205 = {{9{1'b0}}, col_in_1205};
assign u_ca_in_1206 = {{9{1'b0}}, col_in_1206};
assign u_ca_in_1207 = {{9{1'b0}}, col_in_1207};
assign u_ca_in_1208 = {{9{1'b0}}, col_in_1208};
assign u_ca_in_1209 = {{9{1'b0}}, col_in_1209};
assign u_ca_in_1210 = {{9{1'b0}}, col_in_1210};
assign u_ca_in_1211 = {{9{1'b0}}, col_in_1211};
assign u_ca_in_1212 = {{9{1'b0}}, col_in_1212};
assign u_ca_in_1213 = {{9{1'b0}}, col_in_1213};
assign u_ca_in_1214 = {{9{1'b0}}, col_in_1214};
assign u_ca_in_1215 = {{9{1'b0}}, col_in_1215};
assign u_ca_in_1216 = {{9{1'b0}}, col_in_1216};
assign u_ca_in_1217 = {{9{1'b0}}, col_in_1217};
assign u_ca_in_1218 = {{9{1'b0}}, col_in_1218};
assign u_ca_in_1219 = {{9{1'b0}}, col_in_1219};
assign u_ca_in_1220 = {{9{1'b0}}, col_in_1220};
assign u_ca_in_1221 = {{9{1'b0}}, col_in_1221};
assign u_ca_in_1222 = {{9{1'b0}}, col_in_1222};
assign u_ca_in_1223 = {{9{1'b0}}, col_in_1223};
assign u_ca_in_1224 = {{9{1'b0}}, col_in_1224};
assign u_ca_in_1225 = {{9{1'b0}}, col_in_1225};
assign u_ca_in_1226 = {{9{1'b0}}, col_in_1226};
assign u_ca_in_1227 = {{9{1'b0}}, col_in_1227};
assign u_ca_in_1228 = {{9{1'b0}}, col_in_1228};
assign u_ca_in_1229 = {{9{1'b0}}, col_in_1229};
assign u_ca_in_1230 = {{9{1'b0}}, col_in_1230};
assign u_ca_in_1231 = {{9{1'b0}}, col_in_1231};
assign u_ca_in_1232 = {{9{1'b0}}, col_in_1232};
assign u_ca_in_1233 = {{9{1'b0}}, col_in_1233};
assign u_ca_in_1234 = {{9{1'b0}}, col_in_1234};
assign u_ca_in_1235 = {{9{1'b0}}, col_in_1235};
assign u_ca_in_1236 = {{9{1'b0}}, col_in_1236};
assign u_ca_in_1237 = {{9{1'b0}}, col_in_1237};
assign u_ca_in_1238 = {{9{1'b0}}, col_in_1238};
assign u_ca_in_1239 = {{9{1'b0}}, col_in_1239};
assign u_ca_in_1240 = {{9{1'b0}}, col_in_1240};
assign u_ca_in_1241 = {{9{1'b0}}, col_in_1241};
assign u_ca_in_1242 = {{9{1'b0}}, col_in_1242};
assign u_ca_in_1243 = {{9{1'b0}}, col_in_1243};
assign u_ca_in_1244 = {{9{1'b0}}, col_in_1244};
assign u_ca_in_1245 = {{9{1'b0}}, col_in_1245};
assign u_ca_in_1246 = {{9{1'b0}}, col_in_1246};
assign u_ca_in_1247 = {{9{1'b0}}, col_in_1247};
assign u_ca_in_1248 = {{9{1'b0}}, col_in_1248};
assign u_ca_in_1249 = {{9{1'b0}}, col_in_1249};
assign u_ca_in_1250 = {{9{1'b0}}, col_in_1250};
assign u_ca_in_1251 = {{9{1'b0}}, col_in_1251};
assign u_ca_in_1252 = {{9{1'b0}}, col_in_1252};
assign u_ca_in_1253 = {{9{1'b0}}, col_in_1253};
assign u_ca_in_1254 = {{9{1'b0}}, col_in_1254};
assign u_ca_in_1255 = {{9{1'b0}}, col_in_1255};
assign u_ca_in_1256 = {{9{1'b0}}, col_in_1256};
assign u_ca_in_1257 = {{9{1'b0}}, col_in_1257};
assign u_ca_in_1258 = {{9{1'b0}}, col_in_1258};
assign u_ca_in_1259 = {{9{1'b0}}, col_in_1259};
assign u_ca_in_1260 = {{9{1'b0}}, col_in_1260};
assign u_ca_in_1261 = {{9{1'b0}}, col_in_1261};
assign u_ca_in_1262 = {{9{1'b0}}, col_in_1262};
assign u_ca_in_1263 = {{9{1'b0}}, col_in_1263};
assign u_ca_in_1264 = {{9{1'b0}}, col_in_1264};
assign u_ca_in_1265 = {{9{1'b0}}, col_in_1265};
assign u_ca_in_1266 = {{9{1'b0}}, col_in_1266};
assign u_ca_in_1267 = {{9{1'b0}}, col_in_1267};
assign u_ca_in_1268 = {{9{1'b0}}, col_in_1268};
assign u_ca_in_1269 = {{9{1'b0}}, col_in_1269};
assign u_ca_in_1270 = {{9{1'b0}}, col_in_1270};
assign u_ca_in_1271 = {{9{1'b0}}, col_in_1271};
assign u_ca_in_1272 = {{9{1'b0}}, col_in_1272};
assign u_ca_in_1273 = {{9{1'b0}}, col_in_1273};
assign u_ca_in_1274 = {{9{1'b0}}, col_in_1274};
assign u_ca_in_1275 = {{9{1'b0}}, col_in_1275};
assign u_ca_in_1276 = {{9{1'b0}}, col_in_1276};
assign u_ca_in_1277 = {{9{1'b0}}, col_in_1277};
assign u_ca_in_1278 = {{9{1'b0}}, col_in_1278};
assign u_ca_in_1279 = {{9{1'b0}}, col_in_1279};
assign u_ca_in_1280 = {{9{1'b0}}, col_in_1280};
assign u_ca_in_1281 = {{9{1'b0}}, col_in_1281};
assign u_ca_in_1282 = {{9{1'b0}}, col_in_1282};

//---------------------------------------------------------


compressor_81_24 u_ca_81_24_0(.d_in(u_ca_in_0), .d_out(u_ca_out_0));
compressor_81_24 u_ca_81_24_1(.d_in(u_ca_in_1), .d_out(u_ca_out_1));
compressor_81_24 u_ca_81_24_2(.d_in(u_ca_in_2), .d_out(u_ca_out_2));
compressor_81_24 u_ca_81_24_3(.d_in(u_ca_in_3), .d_out(u_ca_out_3));
compressor_81_24 u_ca_81_24_4(.d_in(u_ca_in_4), .d_out(u_ca_out_4));
compressor_81_24 u_ca_81_24_5(.d_in(u_ca_in_5), .d_out(u_ca_out_5));
compressor_81_24 u_ca_81_24_6(.d_in(u_ca_in_6), .d_out(u_ca_out_6));
compressor_81_24 u_ca_81_24_7(.d_in(u_ca_in_7), .d_out(u_ca_out_7));
compressor_81_24 u_ca_81_24_8(.d_in(u_ca_in_8), .d_out(u_ca_out_8));
compressor_81_24 u_ca_81_24_9(.d_in(u_ca_in_9), .d_out(u_ca_out_9));
compressor_81_24 u_ca_81_24_10(.d_in(u_ca_in_10), .d_out(u_ca_out_10));
compressor_81_24 u_ca_81_24_11(.d_in(u_ca_in_11), .d_out(u_ca_out_11));
compressor_81_24 u_ca_81_24_12(.d_in(u_ca_in_12), .d_out(u_ca_out_12));
compressor_81_24 u_ca_81_24_13(.d_in(u_ca_in_13), .d_out(u_ca_out_13));
compressor_81_24 u_ca_81_24_14(.d_in(u_ca_in_14), .d_out(u_ca_out_14));
compressor_81_24 u_ca_81_24_15(.d_in(u_ca_in_15), .d_out(u_ca_out_15));
compressor_81_24 u_ca_81_24_16(.d_in(u_ca_in_16), .d_out(u_ca_out_16));
compressor_81_24 u_ca_81_24_17(.d_in(u_ca_in_17), .d_out(u_ca_out_17));
compressor_81_24 u_ca_81_24_18(.d_in(u_ca_in_18), .d_out(u_ca_out_18));
compressor_81_24 u_ca_81_24_19(.d_in(u_ca_in_19), .d_out(u_ca_out_19));
compressor_81_24 u_ca_81_24_20(.d_in(u_ca_in_20), .d_out(u_ca_out_20));
compressor_81_24 u_ca_81_24_21(.d_in(u_ca_in_21), .d_out(u_ca_out_21));
compressor_81_24 u_ca_81_24_22(.d_in(u_ca_in_22), .d_out(u_ca_out_22));
compressor_81_24 u_ca_81_24_23(.d_in(u_ca_in_23), .d_out(u_ca_out_23));
compressor_81_24 u_ca_81_24_24(.d_in(u_ca_in_24), .d_out(u_ca_out_24));
compressor_81_24 u_ca_81_24_25(.d_in(u_ca_in_25), .d_out(u_ca_out_25));
compressor_81_24 u_ca_81_24_26(.d_in(u_ca_in_26), .d_out(u_ca_out_26));
compressor_81_24 u_ca_81_24_27(.d_in(u_ca_in_27), .d_out(u_ca_out_27));
compressor_81_24 u_ca_81_24_28(.d_in(u_ca_in_28), .d_out(u_ca_out_28));
compressor_81_24 u_ca_81_24_29(.d_in(u_ca_in_29), .d_out(u_ca_out_29));
compressor_81_24 u_ca_81_24_30(.d_in(u_ca_in_30), .d_out(u_ca_out_30));
compressor_81_24 u_ca_81_24_31(.d_in(u_ca_in_31), .d_out(u_ca_out_31));
compressor_81_24 u_ca_81_24_32(.d_in(u_ca_in_32), .d_out(u_ca_out_32));
compressor_81_24 u_ca_81_24_33(.d_in(u_ca_in_33), .d_out(u_ca_out_33));
compressor_81_24 u_ca_81_24_34(.d_in(u_ca_in_34), .d_out(u_ca_out_34));
compressor_81_24 u_ca_81_24_35(.d_in(u_ca_in_35), .d_out(u_ca_out_35));
compressor_81_24 u_ca_81_24_36(.d_in(u_ca_in_36), .d_out(u_ca_out_36));
compressor_81_24 u_ca_81_24_37(.d_in(u_ca_in_37), .d_out(u_ca_out_37));
compressor_81_24 u_ca_81_24_38(.d_in(u_ca_in_38), .d_out(u_ca_out_38));
compressor_81_24 u_ca_81_24_39(.d_in(u_ca_in_39), .d_out(u_ca_out_39));
compressor_81_24 u_ca_81_24_40(.d_in(u_ca_in_40), .d_out(u_ca_out_40));
compressor_81_24 u_ca_81_24_41(.d_in(u_ca_in_41), .d_out(u_ca_out_41));
compressor_81_24 u_ca_81_24_42(.d_in(u_ca_in_42), .d_out(u_ca_out_42));
compressor_81_24 u_ca_81_24_43(.d_in(u_ca_in_43), .d_out(u_ca_out_43));
compressor_81_24 u_ca_81_24_44(.d_in(u_ca_in_44), .d_out(u_ca_out_44));
compressor_81_24 u_ca_81_24_45(.d_in(u_ca_in_45), .d_out(u_ca_out_45));
compressor_81_24 u_ca_81_24_46(.d_in(u_ca_in_46), .d_out(u_ca_out_46));
compressor_81_24 u_ca_81_24_47(.d_in(u_ca_in_47), .d_out(u_ca_out_47));
compressor_81_24 u_ca_81_24_48(.d_in(u_ca_in_48), .d_out(u_ca_out_48));
compressor_81_24 u_ca_81_24_49(.d_in(u_ca_in_49), .d_out(u_ca_out_49));
compressor_81_24 u_ca_81_24_50(.d_in(u_ca_in_50), .d_out(u_ca_out_50));
compressor_81_24 u_ca_81_24_51(.d_in(u_ca_in_51), .d_out(u_ca_out_51));
compressor_81_24 u_ca_81_24_52(.d_in(u_ca_in_52), .d_out(u_ca_out_52));
compressor_81_24 u_ca_81_24_53(.d_in(u_ca_in_53), .d_out(u_ca_out_53));
compressor_81_24 u_ca_81_24_54(.d_in(u_ca_in_54), .d_out(u_ca_out_54));
compressor_81_24 u_ca_81_24_55(.d_in(u_ca_in_55), .d_out(u_ca_out_55));
compressor_81_24 u_ca_81_24_56(.d_in(u_ca_in_56), .d_out(u_ca_out_56));
compressor_81_24 u_ca_81_24_57(.d_in(u_ca_in_57), .d_out(u_ca_out_57));
compressor_81_24 u_ca_81_24_58(.d_in(u_ca_in_58), .d_out(u_ca_out_58));
compressor_81_24 u_ca_81_24_59(.d_in(u_ca_in_59), .d_out(u_ca_out_59));
compressor_81_24 u_ca_81_24_60(.d_in(u_ca_in_60), .d_out(u_ca_out_60));
compressor_81_24 u_ca_81_24_61(.d_in(u_ca_in_61), .d_out(u_ca_out_61));
compressor_81_24 u_ca_81_24_62(.d_in(u_ca_in_62), .d_out(u_ca_out_62));
compressor_81_24 u_ca_81_24_63(.d_in(u_ca_in_63), .d_out(u_ca_out_63));
compressor_81_24 u_ca_81_24_64(.d_in(u_ca_in_64), .d_out(u_ca_out_64));
compressor_81_24 u_ca_81_24_65(.d_in(u_ca_in_65), .d_out(u_ca_out_65));
compressor_81_24 u_ca_81_24_66(.d_in(u_ca_in_66), .d_out(u_ca_out_66));
compressor_81_24 u_ca_81_24_67(.d_in(u_ca_in_67), .d_out(u_ca_out_67));
compressor_81_24 u_ca_81_24_68(.d_in(u_ca_in_68), .d_out(u_ca_out_68));
compressor_81_24 u_ca_81_24_69(.d_in(u_ca_in_69), .d_out(u_ca_out_69));
compressor_81_24 u_ca_81_24_70(.d_in(u_ca_in_70), .d_out(u_ca_out_70));
compressor_81_24 u_ca_81_24_71(.d_in(u_ca_in_71), .d_out(u_ca_out_71));
compressor_81_24 u_ca_81_24_72(.d_in(u_ca_in_72), .d_out(u_ca_out_72));
compressor_81_24 u_ca_81_24_73(.d_in(u_ca_in_73), .d_out(u_ca_out_73));
compressor_81_24 u_ca_81_24_74(.d_in(u_ca_in_74), .d_out(u_ca_out_74));
compressor_81_24 u_ca_81_24_75(.d_in(u_ca_in_75), .d_out(u_ca_out_75));
compressor_81_24 u_ca_81_24_76(.d_in(u_ca_in_76), .d_out(u_ca_out_76));
compressor_81_24 u_ca_81_24_77(.d_in(u_ca_in_77), .d_out(u_ca_out_77));
compressor_81_24 u_ca_81_24_78(.d_in(u_ca_in_78), .d_out(u_ca_out_78));
compressor_81_24 u_ca_81_24_79(.d_in(u_ca_in_79), .d_out(u_ca_out_79));
compressor_81_24 u_ca_81_24_80(.d_in(u_ca_in_80), .d_out(u_ca_out_80));
compressor_81_24 u_ca_81_24_81(.d_in(u_ca_in_81), .d_out(u_ca_out_81));
compressor_81_24 u_ca_81_24_82(.d_in(u_ca_in_82), .d_out(u_ca_out_82));
compressor_81_24 u_ca_81_24_83(.d_in(u_ca_in_83), .d_out(u_ca_out_83));
compressor_81_24 u_ca_81_24_84(.d_in(u_ca_in_84), .d_out(u_ca_out_84));
compressor_81_24 u_ca_81_24_85(.d_in(u_ca_in_85), .d_out(u_ca_out_85));
compressor_81_24 u_ca_81_24_86(.d_in(u_ca_in_86), .d_out(u_ca_out_86));
compressor_81_24 u_ca_81_24_87(.d_in(u_ca_in_87), .d_out(u_ca_out_87));
compressor_81_24 u_ca_81_24_88(.d_in(u_ca_in_88), .d_out(u_ca_out_88));
compressor_81_24 u_ca_81_24_89(.d_in(u_ca_in_89), .d_out(u_ca_out_89));
compressor_81_24 u_ca_81_24_90(.d_in(u_ca_in_90), .d_out(u_ca_out_90));
compressor_81_24 u_ca_81_24_91(.d_in(u_ca_in_91), .d_out(u_ca_out_91));
compressor_81_24 u_ca_81_24_92(.d_in(u_ca_in_92), .d_out(u_ca_out_92));
compressor_81_24 u_ca_81_24_93(.d_in(u_ca_in_93), .d_out(u_ca_out_93));
compressor_81_24 u_ca_81_24_94(.d_in(u_ca_in_94), .d_out(u_ca_out_94));
compressor_81_24 u_ca_81_24_95(.d_in(u_ca_in_95), .d_out(u_ca_out_95));
compressor_81_24 u_ca_81_24_96(.d_in(u_ca_in_96), .d_out(u_ca_out_96));
compressor_81_24 u_ca_81_24_97(.d_in(u_ca_in_97), .d_out(u_ca_out_97));
compressor_81_24 u_ca_81_24_98(.d_in(u_ca_in_98), .d_out(u_ca_out_98));
compressor_81_24 u_ca_81_24_99(.d_in(u_ca_in_99), .d_out(u_ca_out_99));
compressor_81_24 u_ca_81_24_100(.d_in(u_ca_in_100), .d_out(u_ca_out_100));
compressor_81_24 u_ca_81_24_101(.d_in(u_ca_in_101), .d_out(u_ca_out_101));
compressor_81_24 u_ca_81_24_102(.d_in(u_ca_in_102), .d_out(u_ca_out_102));
compressor_81_24 u_ca_81_24_103(.d_in(u_ca_in_103), .d_out(u_ca_out_103));
compressor_81_24 u_ca_81_24_104(.d_in(u_ca_in_104), .d_out(u_ca_out_104));
compressor_81_24 u_ca_81_24_105(.d_in(u_ca_in_105), .d_out(u_ca_out_105));
compressor_81_24 u_ca_81_24_106(.d_in(u_ca_in_106), .d_out(u_ca_out_106));
compressor_81_24 u_ca_81_24_107(.d_in(u_ca_in_107), .d_out(u_ca_out_107));
compressor_81_24 u_ca_81_24_108(.d_in(u_ca_in_108), .d_out(u_ca_out_108));
compressor_81_24 u_ca_81_24_109(.d_in(u_ca_in_109), .d_out(u_ca_out_109));
compressor_81_24 u_ca_81_24_110(.d_in(u_ca_in_110), .d_out(u_ca_out_110));
compressor_81_24 u_ca_81_24_111(.d_in(u_ca_in_111), .d_out(u_ca_out_111));
compressor_81_24 u_ca_81_24_112(.d_in(u_ca_in_112), .d_out(u_ca_out_112));
compressor_81_24 u_ca_81_24_113(.d_in(u_ca_in_113), .d_out(u_ca_out_113));
compressor_81_24 u_ca_81_24_114(.d_in(u_ca_in_114), .d_out(u_ca_out_114));
compressor_81_24 u_ca_81_24_115(.d_in(u_ca_in_115), .d_out(u_ca_out_115));
compressor_81_24 u_ca_81_24_116(.d_in(u_ca_in_116), .d_out(u_ca_out_116));
compressor_81_24 u_ca_81_24_117(.d_in(u_ca_in_117), .d_out(u_ca_out_117));
compressor_81_24 u_ca_81_24_118(.d_in(u_ca_in_118), .d_out(u_ca_out_118));
compressor_81_24 u_ca_81_24_119(.d_in(u_ca_in_119), .d_out(u_ca_out_119));
compressor_81_24 u_ca_81_24_120(.d_in(u_ca_in_120), .d_out(u_ca_out_120));
compressor_81_24 u_ca_81_24_121(.d_in(u_ca_in_121), .d_out(u_ca_out_121));
compressor_81_24 u_ca_81_24_122(.d_in(u_ca_in_122), .d_out(u_ca_out_122));
compressor_81_24 u_ca_81_24_123(.d_in(u_ca_in_123), .d_out(u_ca_out_123));
compressor_81_24 u_ca_81_24_124(.d_in(u_ca_in_124), .d_out(u_ca_out_124));
compressor_81_24 u_ca_81_24_125(.d_in(u_ca_in_125), .d_out(u_ca_out_125));
compressor_81_24 u_ca_81_24_126(.d_in(u_ca_in_126), .d_out(u_ca_out_126));
compressor_81_24 u_ca_81_24_127(.d_in(u_ca_in_127), .d_out(u_ca_out_127));
compressor_81_24 u_ca_81_24_128(.d_in(u_ca_in_128), .d_out(u_ca_out_128));
compressor_81_24 u_ca_81_24_129(.d_in(u_ca_in_129), .d_out(u_ca_out_129));
compressor_81_24 u_ca_81_24_130(.d_in(u_ca_in_130), .d_out(u_ca_out_130));
compressor_81_24 u_ca_81_24_131(.d_in(u_ca_in_131), .d_out(u_ca_out_131));
compressor_81_24 u_ca_81_24_132(.d_in(u_ca_in_132), .d_out(u_ca_out_132));
compressor_81_24 u_ca_81_24_133(.d_in(u_ca_in_133), .d_out(u_ca_out_133));
compressor_81_24 u_ca_81_24_134(.d_in(u_ca_in_134), .d_out(u_ca_out_134));
compressor_81_24 u_ca_81_24_135(.d_in(u_ca_in_135), .d_out(u_ca_out_135));
compressor_81_24 u_ca_81_24_136(.d_in(u_ca_in_136), .d_out(u_ca_out_136));
compressor_81_24 u_ca_81_24_137(.d_in(u_ca_in_137), .d_out(u_ca_out_137));
compressor_81_24 u_ca_81_24_138(.d_in(u_ca_in_138), .d_out(u_ca_out_138));
compressor_81_24 u_ca_81_24_139(.d_in(u_ca_in_139), .d_out(u_ca_out_139));
compressor_81_24 u_ca_81_24_140(.d_in(u_ca_in_140), .d_out(u_ca_out_140));
compressor_81_24 u_ca_81_24_141(.d_in(u_ca_in_141), .d_out(u_ca_out_141));
compressor_81_24 u_ca_81_24_142(.d_in(u_ca_in_142), .d_out(u_ca_out_142));
compressor_81_24 u_ca_81_24_143(.d_in(u_ca_in_143), .d_out(u_ca_out_143));
compressor_81_24 u_ca_81_24_144(.d_in(u_ca_in_144), .d_out(u_ca_out_144));
compressor_81_24 u_ca_81_24_145(.d_in(u_ca_in_145), .d_out(u_ca_out_145));
compressor_81_24 u_ca_81_24_146(.d_in(u_ca_in_146), .d_out(u_ca_out_146));
compressor_81_24 u_ca_81_24_147(.d_in(u_ca_in_147), .d_out(u_ca_out_147));
compressor_81_24 u_ca_81_24_148(.d_in(u_ca_in_148), .d_out(u_ca_out_148));
compressor_81_24 u_ca_81_24_149(.d_in(u_ca_in_149), .d_out(u_ca_out_149));
compressor_81_24 u_ca_81_24_150(.d_in(u_ca_in_150), .d_out(u_ca_out_150));
compressor_81_24 u_ca_81_24_151(.d_in(u_ca_in_151), .d_out(u_ca_out_151));
compressor_81_24 u_ca_81_24_152(.d_in(u_ca_in_152), .d_out(u_ca_out_152));
compressor_81_24 u_ca_81_24_153(.d_in(u_ca_in_153), .d_out(u_ca_out_153));
compressor_81_24 u_ca_81_24_154(.d_in(u_ca_in_154), .d_out(u_ca_out_154));
compressor_81_24 u_ca_81_24_155(.d_in(u_ca_in_155), .d_out(u_ca_out_155));
compressor_81_24 u_ca_81_24_156(.d_in(u_ca_in_156), .d_out(u_ca_out_156));
compressor_81_24 u_ca_81_24_157(.d_in(u_ca_in_157), .d_out(u_ca_out_157));
compressor_81_24 u_ca_81_24_158(.d_in(u_ca_in_158), .d_out(u_ca_out_158));
compressor_81_24 u_ca_81_24_159(.d_in(u_ca_in_159), .d_out(u_ca_out_159));
compressor_81_24 u_ca_81_24_160(.d_in(u_ca_in_160), .d_out(u_ca_out_160));
compressor_81_24 u_ca_81_24_161(.d_in(u_ca_in_161), .d_out(u_ca_out_161));
compressor_81_24 u_ca_81_24_162(.d_in(u_ca_in_162), .d_out(u_ca_out_162));
compressor_81_24 u_ca_81_24_163(.d_in(u_ca_in_163), .d_out(u_ca_out_163));
compressor_81_24 u_ca_81_24_164(.d_in(u_ca_in_164), .d_out(u_ca_out_164));
compressor_81_24 u_ca_81_24_165(.d_in(u_ca_in_165), .d_out(u_ca_out_165));
compressor_81_24 u_ca_81_24_166(.d_in(u_ca_in_166), .d_out(u_ca_out_166));
compressor_81_24 u_ca_81_24_167(.d_in(u_ca_in_167), .d_out(u_ca_out_167));
compressor_81_24 u_ca_81_24_168(.d_in(u_ca_in_168), .d_out(u_ca_out_168));
compressor_81_24 u_ca_81_24_169(.d_in(u_ca_in_169), .d_out(u_ca_out_169));
compressor_81_24 u_ca_81_24_170(.d_in(u_ca_in_170), .d_out(u_ca_out_170));
compressor_81_24 u_ca_81_24_171(.d_in(u_ca_in_171), .d_out(u_ca_out_171));
compressor_81_24 u_ca_81_24_172(.d_in(u_ca_in_172), .d_out(u_ca_out_172));
compressor_81_24 u_ca_81_24_173(.d_in(u_ca_in_173), .d_out(u_ca_out_173));
compressor_81_24 u_ca_81_24_174(.d_in(u_ca_in_174), .d_out(u_ca_out_174));
compressor_81_24 u_ca_81_24_175(.d_in(u_ca_in_175), .d_out(u_ca_out_175));
compressor_81_24 u_ca_81_24_176(.d_in(u_ca_in_176), .d_out(u_ca_out_176));
compressor_81_24 u_ca_81_24_177(.d_in(u_ca_in_177), .d_out(u_ca_out_177));
compressor_81_24 u_ca_81_24_178(.d_in(u_ca_in_178), .d_out(u_ca_out_178));
compressor_81_24 u_ca_81_24_179(.d_in(u_ca_in_179), .d_out(u_ca_out_179));
compressor_81_24 u_ca_81_24_180(.d_in(u_ca_in_180), .d_out(u_ca_out_180));
compressor_81_24 u_ca_81_24_181(.d_in(u_ca_in_181), .d_out(u_ca_out_181));
compressor_81_24 u_ca_81_24_182(.d_in(u_ca_in_182), .d_out(u_ca_out_182));
compressor_81_24 u_ca_81_24_183(.d_in(u_ca_in_183), .d_out(u_ca_out_183));
compressor_81_24 u_ca_81_24_184(.d_in(u_ca_in_184), .d_out(u_ca_out_184));
compressor_81_24 u_ca_81_24_185(.d_in(u_ca_in_185), .d_out(u_ca_out_185));
compressor_81_24 u_ca_81_24_186(.d_in(u_ca_in_186), .d_out(u_ca_out_186));
compressor_81_24 u_ca_81_24_187(.d_in(u_ca_in_187), .d_out(u_ca_out_187));
compressor_81_24 u_ca_81_24_188(.d_in(u_ca_in_188), .d_out(u_ca_out_188));
compressor_81_24 u_ca_81_24_189(.d_in(u_ca_in_189), .d_out(u_ca_out_189));
compressor_81_24 u_ca_81_24_190(.d_in(u_ca_in_190), .d_out(u_ca_out_190));
compressor_81_24 u_ca_81_24_191(.d_in(u_ca_in_191), .d_out(u_ca_out_191));
compressor_81_24 u_ca_81_24_192(.d_in(u_ca_in_192), .d_out(u_ca_out_192));
compressor_81_24 u_ca_81_24_193(.d_in(u_ca_in_193), .d_out(u_ca_out_193));
compressor_81_24 u_ca_81_24_194(.d_in(u_ca_in_194), .d_out(u_ca_out_194));
compressor_81_24 u_ca_81_24_195(.d_in(u_ca_in_195), .d_out(u_ca_out_195));
compressor_81_24 u_ca_81_24_196(.d_in(u_ca_in_196), .d_out(u_ca_out_196));
compressor_81_24 u_ca_81_24_197(.d_in(u_ca_in_197), .d_out(u_ca_out_197));
compressor_81_24 u_ca_81_24_198(.d_in(u_ca_in_198), .d_out(u_ca_out_198));
compressor_81_24 u_ca_81_24_199(.d_in(u_ca_in_199), .d_out(u_ca_out_199));
compressor_81_24 u_ca_81_24_200(.d_in(u_ca_in_200), .d_out(u_ca_out_200));
compressor_81_24 u_ca_81_24_201(.d_in(u_ca_in_201), .d_out(u_ca_out_201));
compressor_81_24 u_ca_81_24_202(.d_in(u_ca_in_202), .d_out(u_ca_out_202));
compressor_81_24 u_ca_81_24_203(.d_in(u_ca_in_203), .d_out(u_ca_out_203));
compressor_81_24 u_ca_81_24_204(.d_in(u_ca_in_204), .d_out(u_ca_out_204));
compressor_81_24 u_ca_81_24_205(.d_in(u_ca_in_205), .d_out(u_ca_out_205));
compressor_81_24 u_ca_81_24_206(.d_in(u_ca_in_206), .d_out(u_ca_out_206));
compressor_81_24 u_ca_81_24_207(.d_in(u_ca_in_207), .d_out(u_ca_out_207));
compressor_81_24 u_ca_81_24_208(.d_in(u_ca_in_208), .d_out(u_ca_out_208));
compressor_81_24 u_ca_81_24_209(.d_in(u_ca_in_209), .d_out(u_ca_out_209));
compressor_81_24 u_ca_81_24_210(.d_in(u_ca_in_210), .d_out(u_ca_out_210));
compressor_81_24 u_ca_81_24_211(.d_in(u_ca_in_211), .d_out(u_ca_out_211));
compressor_81_24 u_ca_81_24_212(.d_in(u_ca_in_212), .d_out(u_ca_out_212));
compressor_81_24 u_ca_81_24_213(.d_in(u_ca_in_213), .d_out(u_ca_out_213));
compressor_81_24 u_ca_81_24_214(.d_in(u_ca_in_214), .d_out(u_ca_out_214));
compressor_81_24 u_ca_81_24_215(.d_in(u_ca_in_215), .d_out(u_ca_out_215));
compressor_81_24 u_ca_81_24_216(.d_in(u_ca_in_216), .d_out(u_ca_out_216));
compressor_81_24 u_ca_81_24_217(.d_in(u_ca_in_217), .d_out(u_ca_out_217));
compressor_81_24 u_ca_81_24_218(.d_in(u_ca_in_218), .d_out(u_ca_out_218));
compressor_81_24 u_ca_81_24_219(.d_in(u_ca_in_219), .d_out(u_ca_out_219));
compressor_81_24 u_ca_81_24_220(.d_in(u_ca_in_220), .d_out(u_ca_out_220));
compressor_81_24 u_ca_81_24_221(.d_in(u_ca_in_221), .d_out(u_ca_out_221));
compressor_81_24 u_ca_81_24_222(.d_in(u_ca_in_222), .d_out(u_ca_out_222));
compressor_81_24 u_ca_81_24_223(.d_in(u_ca_in_223), .d_out(u_ca_out_223));
compressor_81_24 u_ca_81_24_224(.d_in(u_ca_in_224), .d_out(u_ca_out_224));
compressor_81_24 u_ca_81_24_225(.d_in(u_ca_in_225), .d_out(u_ca_out_225));
compressor_81_24 u_ca_81_24_226(.d_in(u_ca_in_226), .d_out(u_ca_out_226));
compressor_81_24 u_ca_81_24_227(.d_in(u_ca_in_227), .d_out(u_ca_out_227));
compressor_81_24 u_ca_81_24_228(.d_in(u_ca_in_228), .d_out(u_ca_out_228));
compressor_81_24 u_ca_81_24_229(.d_in(u_ca_in_229), .d_out(u_ca_out_229));
compressor_81_24 u_ca_81_24_230(.d_in(u_ca_in_230), .d_out(u_ca_out_230));
compressor_81_24 u_ca_81_24_231(.d_in(u_ca_in_231), .d_out(u_ca_out_231));
compressor_81_24 u_ca_81_24_232(.d_in(u_ca_in_232), .d_out(u_ca_out_232));
compressor_81_24 u_ca_81_24_233(.d_in(u_ca_in_233), .d_out(u_ca_out_233));
compressor_81_24 u_ca_81_24_234(.d_in(u_ca_in_234), .d_out(u_ca_out_234));
compressor_81_24 u_ca_81_24_235(.d_in(u_ca_in_235), .d_out(u_ca_out_235));
compressor_81_24 u_ca_81_24_236(.d_in(u_ca_in_236), .d_out(u_ca_out_236));
compressor_81_24 u_ca_81_24_237(.d_in(u_ca_in_237), .d_out(u_ca_out_237));
compressor_81_24 u_ca_81_24_238(.d_in(u_ca_in_238), .d_out(u_ca_out_238));
compressor_81_24 u_ca_81_24_239(.d_in(u_ca_in_239), .d_out(u_ca_out_239));
compressor_81_24 u_ca_81_24_240(.d_in(u_ca_in_240), .d_out(u_ca_out_240));
compressor_81_24 u_ca_81_24_241(.d_in(u_ca_in_241), .d_out(u_ca_out_241));
compressor_81_24 u_ca_81_24_242(.d_in(u_ca_in_242), .d_out(u_ca_out_242));
compressor_81_24 u_ca_81_24_243(.d_in(u_ca_in_243), .d_out(u_ca_out_243));
compressor_81_24 u_ca_81_24_244(.d_in(u_ca_in_244), .d_out(u_ca_out_244));
compressor_81_24 u_ca_81_24_245(.d_in(u_ca_in_245), .d_out(u_ca_out_245));
compressor_81_24 u_ca_81_24_246(.d_in(u_ca_in_246), .d_out(u_ca_out_246));
compressor_81_24 u_ca_81_24_247(.d_in(u_ca_in_247), .d_out(u_ca_out_247));
compressor_81_24 u_ca_81_24_248(.d_in(u_ca_in_248), .d_out(u_ca_out_248));
compressor_81_24 u_ca_81_24_249(.d_in(u_ca_in_249), .d_out(u_ca_out_249));
compressor_81_24 u_ca_81_24_250(.d_in(u_ca_in_250), .d_out(u_ca_out_250));
compressor_81_24 u_ca_81_24_251(.d_in(u_ca_in_251), .d_out(u_ca_out_251));
compressor_81_24 u_ca_81_24_252(.d_in(u_ca_in_252), .d_out(u_ca_out_252));
compressor_81_24 u_ca_81_24_253(.d_in(u_ca_in_253), .d_out(u_ca_out_253));
compressor_81_24 u_ca_81_24_254(.d_in(u_ca_in_254), .d_out(u_ca_out_254));
compressor_81_24 u_ca_81_24_255(.d_in(u_ca_in_255), .d_out(u_ca_out_255));
compressor_81_24 u_ca_81_24_256(.d_in(u_ca_in_256), .d_out(u_ca_out_256));
compressor_81_24 u_ca_81_24_257(.d_in(u_ca_in_257), .d_out(u_ca_out_257));
compressor_81_24 u_ca_81_24_258(.d_in(u_ca_in_258), .d_out(u_ca_out_258));
compressor_81_24 u_ca_81_24_259(.d_in(u_ca_in_259), .d_out(u_ca_out_259));
compressor_81_24 u_ca_81_24_260(.d_in(u_ca_in_260), .d_out(u_ca_out_260));
compressor_81_24 u_ca_81_24_261(.d_in(u_ca_in_261), .d_out(u_ca_out_261));
compressor_81_24 u_ca_81_24_262(.d_in(u_ca_in_262), .d_out(u_ca_out_262));
compressor_81_24 u_ca_81_24_263(.d_in(u_ca_in_263), .d_out(u_ca_out_263));
compressor_81_24 u_ca_81_24_264(.d_in(u_ca_in_264), .d_out(u_ca_out_264));
compressor_81_24 u_ca_81_24_265(.d_in(u_ca_in_265), .d_out(u_ca_out_265));
compressor_81_24 u_ca_81_24_266(.d_in(u_ca_in_266), .d_out(u_ca_out_266));
compressor_81_24 u_ca_81_24_267(.d_in(u_ca_in_267), .d_out(u_ca_out_267));
compressor_81_24 u_ca_81_24_268(.d_in(u_ca_in_268), .d_out(u_ca_out_268));
compressor_81_24 u_ca_81_24_269(.d_in(u_ca_in_269), .d_out(u_ca_out_269));
compressor_81_24 u_ca_81_24_270(.d_in(u_ca_in_270), .d_out(u_ca_out_270));
compressor_81_24 u_ca_81_24_271(.d_in(u_ca_in_271), .d_out(u_ca_out_271));
compressor_81_24 u_ca_81_24_272(.d_in(u_ca_in_272), .d_out(u_ca_out_272));
compressor_81_24 u_ca_81_24_273(.d_in(u_ca_in_273), .d_out(u_ca_out_273));
compressor_81_24 u_ca_81_24_274(.d_in(u_ca_in_274), .d_out(u_ca_out_274));
compressor_81_24 u_ca_81_24_275(.d_in(u_ca_in_275), .d_out(u_ca_out_275));
compressor_81_24 u_ca_81_24_276(.d_in(u_ca_in_276), .d_out(u_ca_out_276));
compressor_81_24 u_ca_81_24_277(.d_in(u_ca_in_277), .d_out(u_ca_out_277));
compressor_81_24 u_ca_81_24_278(.d_in(u_ca_in_278), .d_out(u_ca_out_278));
compressor_81_24 u_ca_81_24_279(.d_in(u_ca_in_279), .d_out(u_ca_out_279));
compressor_81_24 u_ca_81_24_280(.d_in(u_ca_in_280), .d_out(u_ca_out_280));
compressor_81_24 u_ca_81_24_281(.d_in(u_ca_in_281), .d_out(u_ca_out_281));
compressor_81_24 u_ca_81_24_282(.d_in(u_ca_in_282), .d_out(u_ca_out_282));
compressor_81_24 u_ca_81_24_283(.d_in(u_ca_in_283), .d_out(u_ca_out_283));
compressor_81_24 u_ca_81_24_284(.d_in(u_ca_in_284), .d_out(u_ca_out_284));
compressor_81_24 u_ca_81_24_285(.d_in(u_ca_in_285), .d_out(u_ca_out_285));
compressor_81_24 u_ca_81_24_286(.d_in(u_ca_in_286), .d_out(u_ca_out_286));
compressor_81_24 u_ca_81_24_287(.d_in(u_ca_in_287), .d_out(u_ca_out_287));
compressor_81_24 u_ca_81_24_288(.d_in(u_ca_in_288), .d_out(u_ca_out_288));
compressor_81_24 u_ca_81_24_289(.d_in(u_ca_in_289), .d_out(u_ca_out_289));
compressor_81_24 u_ca_81_24_290(.d_in(u_ca_in_290), .d_out(u_ca_out_290));
compressor_81_24 u_ca_81_24_291(.d_in(u_ca_in_291), .d_out(u_ca_out_291));
compressor_81_24 u_ca_81_24_292(.d_in(u_ca_in_292), .d_out(u_ca_out_292));
compressor_81_24 u_ca_81_24_293(.d_in(u_ca_in_293), .d_out(u_ca_out_293));
compressor_81_24 u_ca_81_24_294(.d_in(u_ca_in_294), .d_out(u_ca_out_294));
compressor_81_24 u_ca_81_24_295(.d_in(u_ca_in_295), .d_out(u_ca_out_295));
compressor_81_24 u_ca_81_24_296(.d_in(u_ca_in_296), .d_out(u_ca_out_296));
compressor_81_24 u_ca_81_24_297(.d_in(u_ca_in_297), .d_out(u_ca_out_297));
compressor_81_24 u_ca_81_24_298(.d_in(u_ca_in_298), .d_out(u_ca_out_298));
compressor_81_24 u_ca_81_24_299(.d_in(u_ca_in_299), .d_out(u_ca_out_299));
compressor_81_24 u_ca_81_24_300(.d_in(u_ca_in_300), .d_out(u_ca_out_300));
compressor_81_24 u_ca_81_24_301(.d_in(u_ca_in_301), .d_out(u_ca_out_301));
compressor_81_24 u_ca_81_24_302(.d_in(u_ca_in_302), .d_out(u_ca_out_302));
compressor_81_24 u_ca_81_24_303(.d_in(u_ca_in_303), .d_out(u_ca_out_303));
compressor_81_24 u_ca_81_24_304(.d_in(u_ca_in_304), .d_out(u_ca_out_304));
compressor_81_24 u_ca_81_24_305(.d_in(u_ca_in_305), .d_out(u_ca_out_305));
compressor_81_24 u_ca_81_24_306(.d_in(u_ca_in_306), .d_out(u_ca_out_306));
compressor_81_24 u_ca_81_24_307(.d_in(u_ca_in_307), .d_out(u_ca_out_307));
compressor_81_24 u_ca_81_24_308(.d_in(u_ca_in_308), .d_out(u_ca_out_308));
compressor_81_24 u_ca_81_24_309(.d_in(u_ca_in_309), .d_out(u_ca_out_309));
compressor_81_24 u_ca_81_24_310(.d_in(u_ca_in_310), .d_out(u_ca_out_310));
compressor_81_24 u_ca_81_24_311(.d_in(u_ca_in_311), .d_out(u_ca_out_311));
compressor_81_24 u_ca_81_24_312(.d_in(u_ca_in_312), .d_out(u_ca_out_312));
compressor_81_24 u_ca_81_24_313(.d_in(u_ca_in_313), .d_out(u_ca_out_313));
compressor_81_24 u_ca_81_24_314(.d_in(u_ca_in_314), .d_out(u_ca_out_314));
compressor_81_24 u_ca_81_24_315(.d_in(u_ca_in_315), .d_out(u_ca_out_315));
compressor_81_24 u_ca_81_24_316(.d_in(u_ca_in_316), .d_out(u_ca_out_316));
compressor_81_24 u_ca_81_24_317(.d_in(u_ca_in_317), .d_out(u_ca_out_317));
compressor_81_24 u_ca_81_24_318(.d_in(u_ca_in_318), .d_out(u_ca_out_318));
compressor_81_24 u_ca_81_24_319(.d_in(u_ca_in_319), .d_out(u_ca_out_319));
compressor_81_24 u_ca_81_24_320(.d_in(u_ca_in_320), .d_out(u_ca_out_320));
compressor_81_24 u_ca_81_24_321(.d_in(u_ca_in_321), .d_out(u_ca_out_321));
compressor_81_24 u_ca_81_24_322(.d_in(u_ca_in_322), .d_out(u_ca_out_322));
compressor_81_24 u_ca_81_24_323(.d_in(u_ca_in_323), .d_out(u_ca_out_323));
compressor_81_24 u_ca_81_24_324(.d_in(u_ca_in_324), .d_out(u_ca_out_324));
compressor_81_24 u_ca_81_24_325(.d_in(u_ca_in_325), .d_out(u_ca_out_325));
compressor_81_24 u_ca_81_24_326(.d_in(u_ca_in_326), .d_out(u_ca_out_326));
compressor_81_24 u_ca_81_24_327(.d_in(u_ca_in_327), .d_out(u_ca_out_327));
compressor_81_24 u_ca_81_24_328(.d_in(u_ca_in_328), .d_out(u_ca_out_328));
compressor_81_24 u_ca_81_24_329(.d_in(u_ca_in_329), .d_out(u_ca_out_329));
compressor_81_24 u_ca_81_24_330(.d_in(u_ca_in_330), .d_out(u_ca_out_330));
compressor_81_24 u_ca_81_24_331(.d_in(u_ca_in_331), .d_out(u_ca_out_331));
compressor_81_24 u_ca_81_24_332(.d_in(u_ca_in_332), .d_out(u_ca_out_332));
compressor_81_24 u_ca_81_24_333(.d_in(u_ca_in_333), .d_out(u_ca_out_333));
compressor_81_24 u_ca_81_24_334(.d_in(u_ca_in_334), .d_out(u_ca_out_334));
compressor_81_24 u_ca_81_24_335(.d_in(u_ca_in_335), .d_out(u_ca_out_335));
compressor_81_24 u_ca_81_24_336(.d_in(u_ca_in_336), .d_out(u_ca_out_336));
compressor_81_24 u_ca_81_24_337(.d_in(u_ca_in_337), .d_out(u_ca_out_337));
compressor_81_24 u_ca_81_24_338(.d_in(u_ca_in_338), .d_out(u_ca_out_338));
compressor_81_24 u_ca_81_24_339(.d_in(u_ca_in_339), .d_out(u_ca_out_339));
compressor_81_24 u_ca_81_24_340(.d_in(u_ca_in_340), .d_out(u_ca_out_340));
compressor_81_24 u_ca_81_24_341(.d_in(u_ca_in_341), .d_out(u_ca_out_341));
compressor_81_24 u_ca_81_24_342(.d_in(u_ca_in_342), .d_out(u_ca_out_342));
compressor_81_24 u_ca_81_24_343(.d_in(u_ca_in_343), .d_out(u_ca_out_343));
compressor_81_24 u_ca_81_24_344(.d_in(u_ca_in_344), .d_out(u_ca_out_344));
compressor_81_24 u_ca_81_24_345(.d_in(u_ca_in_345), .d_out(u_ca_out_345));
compressor_81_24 u_ca_81_24_346(.d_in(u_ca_in_346), .d_out(u_ca_out_346));
compressor_81_24 u_ca_81_24_347(.d_in(u_ca_in_347), .d_out(u_ca_out_347));
compressor_81_24 u_ca_81_24_348(.d_in(u_ca_in_348), .d_out(u_ca_out_348));
compressor_81_24 u_ca_81_24_349(.d_in(u_ca_in_349), .d_out(u_ca_out_349));
compressor_81_24 u_ca_81_24_350(.d_in(u_ca_in_350), .d_out(u_ca_out_350));
compressor_81_24 u_ca_81_24_351(.d_in(u_ca_in_351), .d_out(u_ca_out_351));
compressor_81_24 u_ca_81_24_352(.d_in(u_ca_in_352), .d_out(u_ca_out_352));
compressor_81_24 u_ca_81_24_353(.d_in(u_ca_in_353), .d_out(u_ca_out_353));
compressor_81_24 u_ca_81_24_354(.d_in(u_ca_in_354), .d_out(u_ca_out_354));
compressor_81_24 u_ca_81_24_355(.d_in(u_ca_in_355), .d_out(u_ca_out_355));
compressor_81_24 u_ca_81_24_356(.d_in(u_ca_in_356), .d_out(u_ca_out_356));
compressor_81_24 u_ca_81_24_357(.d_in(u_ca_in_357), .d_out(u_ca_out_357));
compressor_81_24 u_ca_81_24_358(.d_in(u_ca_in_358), .d_out(u_ca_out_358));
compressor_81_24 u_ca_81_24_359(.d_in(u_ca_in_359), .d_out(u_ca_out_359));
compressor_81_24 u_ca_81_24_360(.d_in(u_ca_in_360), .d_out(u_ca_out_360));
compressor_81_24 u_ca_81_24_361(.d_in(u_ca_in_361), .d_out(u_ca_out_361));
compressor_81_24 u_ca_81_24_362(.d_in(u_ca_in_362), .d_out(u_ca_out_362));
compressor_81_24 u_ca_81_24_363(.d_in(u_ca_in_363), .d_out(u_ca_out_363));
compressor_81_24 u_ca_81_24_364(.d_in(u_ca_in_364), .d_out(u_ca_out_364));
compressor_81_24 u_ca_81_24_365(.d_in(u_ca_in_365), .d_out(u_ca_out_365));
compressor_81_24 u_ca_81_24_366(.d_in(u_ca_in_366), .d_out(u_ca_out_366));
compressor_81_24 u_ca_81_24_367(.d_in(u_ca_in_367), .d_out(u_ca_out_367));
compressor_81_24 u_ca_81_24_368(.d_in(u_ca_in_368), .d_out(u_ca_out_368));
compressor_81_24 u_ca_81_24_369(.d_in(u_ca_in_369), .d_out(u_ca_out_369));
compressor_81_24 u_ca_81_24_370(.d_in(u_ca_in_370), .d_out(u_ca_out_370));
compressor_81_24 u_ca_81_24_371(.d_in(u_ca_in_371), .d_out(u_ca_out_371));
compressor_81_24 u_ca_81_24_372(.d_in(u_ca_in_372), .d_out(u_ca_out_372));
compressor_81_24 u_ca_81_24_373(.d_in(u_ca_in_373), .d_out(u_ca_out_373));
compressor_81_24 u_ca_81_24_374(.d_in(u_ca_in_374), .d_out(u_ca_out_374));
compressor_81_24 u_ca_81_24_375(.d_in(u_ca_in_375), .d_out(u_ca_out_375));
compressor_81_24 u_ca_81_24_376(.d_in(u_ca_in_376), .d_out(u_ca_out_376));
compressor_81_24 u_ca_81_24_377(.d_in(u_ca_in_377), .d_out(u_ca_out_377));
compressor_81_24 u_ca_81_24_378(.d_in(u_ca_in_378), .d_out(u_ca_out_378));
compressor_81_24 u_ca_81_24_379(.d_in(u_ca_in_379), .d_out(u_ca_out_379));
compressor_81_24 u_ca_81_24_380(.d_in(u_ca_in_380), .d_out(u_ca_out_380));
compressor_81_24 u_ca_81_24_381(.d_in(u_ca_in_381), .d_out(u_ca_out_381));
compressor_81_24 u_ca_81_24_382(.d_in(u_ca_in_382), .d_out(u_ca_out_382));
compressor_81_24 u_ca_81_24_383(.d_in(u_ca_in_383), .d_out(u_ca_out_383));
compressor_81_24 u_ca_81_24_384(.d_in(u_ca_in_384), .d_out(u_ca_out_384));
compressor_81_24 u_ca_81_24_385(.d_in(u_ca_in_385), .d_out(u_ca_out_385));
compressor_81_24 u_ca_81_24_386(.d_in(u_ca_in_386), .d_out(u_ca_out_386));
compressor_81_24 u_ca_81_24_387(.d_in(u_ca_in_387), .d_out(u_ca_out_387));
compressor_81_24 u_ca_81_24_388(.d_in(u_ca_in_388), .d_out(u_ca_out_388));
compressor_81_24 u_ca_81_24_389(.d_in(u_ca_in_389), .d_out(u_ca_out_389));
compressor_81_24 u_ca_81_24_390(.d_in(u_ca_in_390), .d_out(u_ca_out_390));
compressor_81_24 u_ca_81_24_391(.d_in(u_ca_in_391), .d_out(u_ca_out_391));
compressor_81_24 u_ca_81_24_392(.d_in(u_ca_in_392), .d_out(u_ca_out_392));
compressor_81_24 u_ca_81_24_393(.d_in(u_ca_in_393), .d_out(u_ca_out_393));
compressor_81_24 u_ca_81_24_394(.d_in(u_ca_in_394), .d_out(u_ca_out_394));
compressor_81_24 u_ca_81_24_395(.d_in(u_ca_in_395), .d_out(u_ca_out_395));
compressor_81_24 u_ca_81_24_396(.d_in(u_ca_in_396), .d_out(u_ca_out_396));
compressor_81_24 u_ca_81_24_397(.d_in(u_ca_in_397), .d_out(u_ca_out_397));
compressor_81_24 u_ca_81_24_398(.d_in(u_ca_in_398), .d_out(u_ca_out_398));
compressor_81_24 u_ca_81_24_399(.d_in(u_ca_in_399), .d_out(u_ca_out_399));
compressor_81_24 u_ca_81_24_400(.d_in(u_ca_in_400), .d_out(u_ca_out_400));
compressor_81_24 u_ca_81_24_401(.d_in(u_ca_in_401), .d_out(u_ca_out_401));
compressor_81_24 u_ca_81_24_402(.d_in(u_ca_in_402), .d_out(u_ca_out_402));
compressor_81_24 u_ca_81_24_403(.d_in(u_ca_in_403), .d_out(u_ca_out_403));
compressor_81_24 u_ca_81_24_404(.d_in(u_ca_in_404), .d_out(u_ca_out_404));
compressor_81_24 u_ca_81_24_405(.d_in(u_ca_in_405), .d_out(u_ca_out_405));
compressor_81_24 u_ca_81_24_406(.d_in(u_ca_in_406), .d_out(u_ca_out_406));
compressor_81_24 u_ca_81_24_407(.d_in(u_ca_in_407), .d_out(u_ca_out_407));
compressor_81_24 u_ca_81_24_408(.d_in(u_ca_in_408), .d_out(u_ca_out_408));
compressor_81_24 u_ca_81_24_409(.d_in(u_ca_in_409), .d_out(u_ca_out_409));
compressor_81_24 u_ca_81_24_410(.d_in(u_ca_in_410), .d_out(u_ca_out_410));
compressor_81_24 u_ca_81_24_411(.d_in(u_ca_in_411), .d_out(u_ca_out_411));
compressor_81_24 u_ca_81_24_412(.d_in(u_ca_in_412), .d_out(u_ca_out_412));
compressor_81_24 u_ca_81_24_413(.d_in(u_ca_in_413), .d_out(u_ca_out_413));
compressor_81_24 u_ca_81_24_414(.d_in(u_ca_in_414), .d_out(u_ca_out_414));
compressor_81_24 u_ca_81_24_415(.d_in(u_ca_in_415), .d_out(u_ca_out_415));
compressor_81_24 u_ca_81_24_416(.d_in(u_ca_in_416), .d_out(u_ca_out_416));
compressor_81_24 u_ca_81_24_417(.d_in(u_ca_in_417), .d_out(u_ca_out_417));
compressor_81_24 u_ca_81_24_418(.d_in(u_ca_in_418), .d_out(u_ca_out_418));
compressor_81_24 u_ca_81_24_419(.d_in(u_ca_in_419), .d_out(u_ca_out_419));
compressor_81_24 u_ca_81_24_420(.d_in(u_ca_in_420), .d_out(u_ca_out_420));
compressor_81_24 u_ca_81_24_421(.d_in(u_ca_in_421), .d_out(u_ca_out_421));
compressor_81_24 u_ca_81_24_422(.d_in(u_ca_in_422), .d_out(u_ca_out_422));
compressor_81_24 u_ca_81_24_423(.d_in(u_ca_in_423), .d_out(u_ca_out_423));
compressor_81_24 u_ca_81_24_424(.d_in(u_ca_in_424), .d_out(u_ca_out_424));
compressor_81_24 u_ca_81_24_425(.d_in(u_ca_in_425), .d_out(u_ca_out_425));
compressor_81_24 u_ca_81_24_426(.d_in(u_ca_in_426), .d_out(u_ca_out_426));
compressor_81_24 u_ca_81_24_427(.d_in(u_ca_in_427), .d_out(u_ca_out_427));
compressor_81_24 u_ca_81_24_428(.d_in(u_ca_in_428), .d_out(u_ca_out_428));
compressor_81_24 u_ca_81_24_429(.d_in(u_ca_in_429), .d_out(u_ca_out_429));
compressor_81_24 u_ca_81_24_430(.d_in(u_ca_in_430), .d_out(u_ca_out_430));
compressor_81_24 u_ca_81_24_431(.d_in(u_ca_in_431), .d_out(u_ca_out_431));
compressor_81_24 u_ca_81_24_432(.d_in(u_ca_in_432), .d_out(u_ca_out_432));
compressor_81_24 u_ca_81_24_433(.d_in(u_ca_in_433), .d_out(u_ca_out_433));
compressor_81_24 u_ca_81_24_434(.d_in(u_ca_in_434), .d_out(u_ca_out_434));
compressor_81_24 u_ca_81_24_435(.d_in(u_ca_in_435), .d_out(u_ca_out_435));
compressor_81_24 u_ca_81_24_436(.d_in(u_ca_in_436), .d_out(u_ca_out_436));
compressor_81_24 u_ca_81_24_437(.d_in(u_ca_in_437), .d_out(u_ca_out_437));
compressor_81_24 u_ca_81_24_438(.d_in(u_ca_in_438), .d_out(u_ca_out_438));
compressor_81_24 u_ca_81_24_439(.d_in(u_ca_in_439), .d_out(u_ca_out_439));
compressor_81_24 u_ca_81_24_440(.d_in(u_ca_in_440), .d_out(u_ca_out_440));
compressor_81_24 u_ca_81_24_441(.d_in(u_ca_in_441), .d_out(u_ca_out_441));
compressor_81_24 u_ca_81_24_442(.d_in(u_ca_in_442), .d_out(u_ca_out_442));
compressor_81_24 u_ca_81_24_443(.d_in(u_ca_in_443), .d_out(u_ca_out_443));
compressor_81_24 u_ca_81_24_444(.d_in(u_ca_in_444), .d_out(u_ca_out_444));
compressor_81_24 u_ca_81_24_445(.d_in(u_ca_in_445), .d_out(u_ca_out_445));
compressor_81_24 u_ca_81_24_446(.d_in(u_ca_in_446), .d_out(u_ca_out_446));
compressor_81_24 u_ca_81_24_447(.d_in(u_ca_in_447), .d_out(u_ca_out_447));
compressor_81_24 u_ca_81_24_448(.d_in(u_ca_in_448), .d_out(u_ca_out_448));
compressor_81_24 u_ca_81_24_449(.d_in(u_ca_in_449), .d_out(u_ca_out_449));
compressor_81_24 u_ca_81_24_450(.d_in(u_ca_in_450), .d_out(u_ca_out_450));
compressor_81_24 u_ca_81_24_451(.d_in(u_ca_in_451), .d_out(u_ca_out_451));
compressor_81_24 u_ca_81_24_452(.d_in(u_ca_in_452), .d_out(u_ca_out_452));
compressor_81_24 u_ca_81_24_453(.d_in(u_ca_in_453), .d_out(u_ca_out_453));
compressor_81_24 u_ca_81_24_454(.d_in(u_ca_in_454), .d_out(u_ca_out_454));
compressor_81_24 u_ca_81_24_455(.d_in(u_ca_in_455), .d_out(u_ca_out_455));
compressor_81_24 u_ca_81_24_456(.d_in(u_ca_in_456), .d_out(u_ca_out_456));
compressor_81_24 u_ca_81_24_457(.d_in(u_ca_in_457), .d_out(u_ca_out_457));
compressor_81_24 u_ca_81_24_458(.d_in(u_ca_in_458), .d_out(u_ca_out_458));
compressor_81_24 u_ca_81_24_459(.d_in(u_ca_in_459), .d_out(u_ca_out_459));
compressor_81_24 u_ca_81_24_460(.d_in(u_ca_in_460), .d_out(u_ca_out_460));
compressor_81_24 u_ca_81_24_461(.d_in(u_ca_in_461), .d_out(u_ca_out_461));
compressor_81_24 u_ca_81_24_462(.d_in(u_ca_in_462), .d_out(u_ca_out_462));
compressor_81_24 u_ca_81_24_463(.d_in(u_ca_in_463), .d_out(u_ca_out_463));
compressor_81_24 u_ca_81_24_464(.d_in(u_ca_in_464), .d_out(u_ca_out_464));
compressor_81_24 u_ca_81_24_465(.d_in(u_ca_in_465), .d_out(u_ca_out_465));
compressor_81_24 u_ca_81_24_466(.d_in(u_ca_in_466), .d_out(u_ca_out_466));
compressor_81_24 u_ca_81_24_467(.d_in(u_ca_in_467), .d_out(u_ca_out_467));
compressor_81_24 u_ca_81_24_468(.d_in(u_ca_in_468), .d_out(u_ca_out_468));
compressor_81_24 u_ca_81_24_469(.d_in(u_ca_in_469), .d_out(u_ca_out_469));
compressor_81_24 u_ca_81_24_470(.d_in(u_ca_in_470), .d_out(u_ca_out_470));
compressor_81_24 u_ca_81_24_471(.d_in(u_ca_in_471), .d_out(u_ca_out_471));
compressor_81_24 u_ca_81_24_472(.d_in(u_ca_in_472), .d_out(u_ca_out_472));
compressor_81_24 u_ca_81_24_473(.d_in(u_ca_in_473), .d_out(u_ca_out_473));
compressor_81_24 u_ca_81_24_474(.d_in(u_ca_in_474), .d_out(u_ca_out_474));
compressor_81_24 u_ca_81_24_475(.d_in(u_ca_in_475), .d_out(u_ca_out_475));
compressor_81_24 u_ca_81_24_476(.d_in(u_ca_in_476), .d_out(u_ca_out_476));
compressor_81_24 u_ca_81_24_477(.d_in(u_ca_in_477), .d_out(u_ca_out_477));
compressor_81_24 u_ca_81_24_478(.d_in(u_ca_in_478), .d_out(u_ca_out_478));
compressor_81_24 u_ca_81_24_479(.d_in(u_ca_in_479), .d_out(u_ca_out_479));
compressor_81_24 u_ca_81_24_480(.d_in(u_ca_in_480), .d_out(u_ca_out_480));
compressor_81_24 u_ca_81_24_481(.d_in(u_ca_in_481), .d_out(u_ca_out_481));
compressor_81_24 u_ca_81_24_482(.d_in(u_ca_in_482), .d_out(u_ca_out_482));
compressor_81_24 u_ca_81_24_483(.d_in(u_ca_in_483), .d_out(u_ca_out_483));
compressor_81_24 u_ca_81_24_484(.d_in(u_ca_in_484), .d_out(u_ca_out_484));
compressor_81_24 u_ca_81_24_485(.d_in(u_ca_in_485), .d_out(u_ca_out_485));
compressor_81_24 u_ca_81_24_486(.d_in(u_ca_in_486), .d_out(u_ca_out_486));
compressor_81_24 u_ca_81_24_487(.d_in(u_ca_in_487), .d_out(u_ca_out_487));
compressor_81_24 u_ca_81_24_488(.d_in(u_ca_in_488), .d_out(u_ca_out_488));
compressor_81_24 u_ca_81_24_489(.d_in(u_ca_in_489), .d_out(u_ca_out_489));
compressor_81_24 u_ca_81_24_490(.d_in(u_ca_in_490), .d_out(u_ca_out_490));
compressor_81_24 u_ca_81_24_491(.d_in(u_ca_in_491), .d_out(u_ca_out_491));
compressor_81_24 u_ca_81_24_492(.d_in(u_ca_in_492), .d_out(u_ca_out_492));
compressor_81_24 u_ca_81_24_493(.d_in(u_ca_in_493), .d_out(u_ca_out_493));
compressor_81_24 u_ca_81_24_494(.d_in(u_ca_in_494), .d_out(u_ca_out_494));
compressor_81_24 u_ca_81_24_495(.d_in(u_ca_in_495), .d_out(u_ca_out_495));
compressor_81_24 u_ca_81_24_496(.d_in(u_ca_in_496), .d_out(u_ca_out_496));
compressor_81_24 u_ca_81_24_497(.d_in(u_ca_in_497), .d_out(u_ca_out_497));
compressor_81_24 u_ca_81_24_498(.d_in(u_ca_in_498), .d_out(u_ca_out_498));
compressor_81_24 u_ca_81_24_499(.d_in(u_ca_in_499), .d_out(u_ca_out_499));
compressor_81_24 u_ca_81_24_500(.d_in(u_ca_in_500), .d_out(u_ca_out_500));
compressor_81_24 u_ca_81_24_501(.d_in(u_ca_in_501), .d_out(u_ca_out_501));
compressor_81_24 u_ca_81_24_502(.d_in(u_ca_in_502), .d_out(u_ca_out_502));
compressor_81_24 u_ca_81_24_503(.d_in(u_ca_in_503), .d_out(u_ca_out_503));
compressor_81_24 u_ca_81_24_504(.d_in(u_ca_in_504), .d_out(u_ca_out_504));
compressor_81_24 u_ca_81_24_505(.d_in(u_ca_in_505), .d_out(u_ca_out_505));
compressor_81_24 u_ca_81_24_506(.d_in(u_ca_in_506), .d_out(u_ca_out_506));
compressor_81_24 u_ca_81_24_507(.d_in(u_ca_in_507), .d_out(u_ca_out_507));
compressor_81_24 u_ca_81_24_508(.d_in(u_ca_in_508), .d_out(u_ca_out_508));
compressor_81_24 u_ca_81_24_509(.d_in(u_ca_in_509), .d_out(u_ca_out_509));
compressor_81_24 u_ca_81_24_510(.d_in(u_ca_in_510), .d_out(u_ca_out_510));
compressor_81_24 u_ca_81_24_511(.d_in(u_ca_in_511), .d_out(u_ca_out_511));
compressor_81_24 u_ca_81_24_512(.d_in(u_ca_in_512), .d_out(u_ca_out_512));
compressor_81_24 u_ca_81_24_513(.d_in(u_ca_in_513), .d_out(u_ca_out_513));
compressor_81_24 u_ca_81_24_514(.d_in(u_ca_in_514), .d_out(u_ca_out_514));
compressor_81_24 u_ca_81_24_515(.d_in(u_ca_in_515), .d_out(u_ca_out_515));
compressor_81_24 u_ca_81_24_516(.d_in(u_ca_in_516), .d_out(u_ca_out_516));
compressor_81_24 u_ca_81_24_517(.d_in(u_ca_in_517), .d_out(u_ca_out_517));
compressor_81_24 u_ca_81_24_518(.d_in(u_ca_in_518), .d_out(u_ca_out_518));
compressor_81_24 u_ca_81_24_519(.d_in(u_ca_in_519), .d_out(u_ca_out_519));
compressor_81_24 u_ca_81_24_520(.d_in(u_ca_in_520), .d_out(u_ca_out_520));
compressor_81_24 u_ca_81_24_521(.d_in(u_ca_in_521), .d_out(u_ca_out_521));
compressor_81_24 u_ca_81_24_522(.d_in(u_ca_in_522), .d_out(u_ca_out_522));
compressor_81_24 u_ca_81_24_523(.d_in(u_ca_in_523), .d_out(u_ca_out_523));
compressor_81_24 u_ca_81_24_524(.d_in(u_ca_in_524), .d_out(u_ca_out_524));
compressor_81_24 u_ca_81_24_525(.d_in(u_ca_in_525), .d_out(u_ca_out_525));
compressor_81_24 u_ca_81_24_526(.d_in(u_ca_in_526), .d_out(u_ca_out_526));
compressor_81_24 u_ca_81_24_527(.d_in(u_ca_in_527), .d_out(u_ca_out_527));
compressor_81_24 u_ca_81_24_528(.d_in(u_ca_in_528), .d_out(u_ca_out_528));
compressor_81_24 u_ca_81_24_529(.d_in(u_ca_in_529), .d_out(u_ca_out_529));
compressor_81_24 u_ca_81_24_530(.d_in(u_ca_in_530), .d_out(u_ca_out_530));
compressor_81_24 u_ca_81_24_531(.d_in(u_ca_in_531), .d_out(u_ca_out_531));
compressor_81_24 u_ca_81_24_532(.d_in(u_ca_in_532), .d_out(u_ca_out_532));
compressor_81_24 u_ca_81_24_533(.d_in(u_ca_in_533), .d_out(u_ca_out_533));
compressor_81_24 u_ca_81_24_534(.d_in(u_ca_in_534), .d_out(u_ca_out_534));
compressor_81_24 u_ca_81_24_535(.d_in(u_ca_in_535), .d_out(u_ca_out_535));
compressor_81_24 u_ca_81_24_536(.d_in(u_ca_in_536), .d_out(u_ca_out_536));
compressor_81_24 u_ca_81_24_537(.d_in(u_ca_in_537), .d_out(u_ca_out_537));
compressor_81_24 u_ca_81_24_538(.d_in(u_ca_in_538), .d_out(u_ca_out_538));
compressor_81_24 u_ca_81_24_539(.d_in(u_ca_in_539), .d_out(u_ca_out_539));
compressor_81_24 u_ca_81_24_540(.d_in(u_ca_in_540), .d_out(u_ca_out_540));
compressor_81_24 u_ca_81_24_541(.d_in(u_ca_in_541), .d_out(u_ca_out_541));
compressor_81_24 u_ca_81_24_542(.d_in(u_ca_in_542), .d_out(u_ca_out_542));
compressor_81_24 u_ca_81_24_543(.d_in(u_ca_in_543), .d_out(u_ca_out_543));
compressor_81_24 u_ca_81_24_544(.d_in(u_ca_in_544), .d_out(u_ca_out_544));
compressor_81_24 u_ca_81_24_545(.d_in(u_ca_in_545), .d_out(u_ca_out_545));
compressor_81_24 u_ca_81_24_546(.d_in(u_ca_in_546), .d_out(u_ca_out_546));
compressor_81_24 u_ca_81_24_547(.d_in(u_ca_in_547), .d_out(u_ca_out_547));
compressor_81_24 u_ca_81_24_548(.d_in(u_ca_in_548), .d_out(u_ca_out_548));
compressor_81_24 u_ca_81_24_549(.d_in(u_ca_in_549), .d_out(u_ca_out_549));
compressor_81_24 u_ca_81_24_550(.d_in(u_ca_in_550), .d_out(u_ca_out_550));
compressor_81_24 u_ca_81_24_551(.d_in(u_ca_in_551), .d_out(u_ca_out_551));
compressor_81_24 u_ca_81_24_552(.d_in(u_ca_in_552), .d_out(u_ca_out_552));
compressor_81_24 u_ca_81_24_553(.d_in(u_ca_in_553), .d_out(u_ca_out_553));
compressor_81_24 u_ca_81_24_554(.d_in(u_ca_in_554), .d_out(u_ca_out_554));
compressor_81_24 u_ca_81_24_555(.d_in(u_ca_in_555), .d_out(u_ca_out_555));
compressor_81_24 u_ca_81_24_556(.d_in(u_ca_in_556), .d_out(u_ca_out_556));
compressor_81_24 u_ca_81_24_557(.d_in(u_ca_in_557), .d_out(u_ca_out_557));
compressor_81_24 u_ca_81_24_558(.d_in(u_ca_in_558), .d_out(u_ca_out_558));
compressor_81_24 u_ca_81_24_559(.d_in(u_ca_in_559), .d_out(u_ca_out_559));
compressor_81_24 u_ca_81_24_560(.d_in(u_ca_in_560), .d_out(u_ca_out_560));
compressor_81_24 u_ca_81_24_561(.d_in(u_ca_in_561), .d_out(u_ca_out_561));
compressor_81_24 u_ca_81_24_562(.d_in(u_ca_in_562), .d_out(u_ca_out_562));
compressor_81_24 u_ca_81_24_563(.d_in(u_ca_in_563), .d_out(u_ca_out_563));
compressor_81_24 u_ca_81_24_564(.d_in(u_ca_in_564), .d_out(u_ca_out_564));
compressor_81_24 u_ca_81_24_565(.d_in(u_ca_in_565), .d_out(u_ca_out_565));
compressor_81_24 u_ca_81_24_566(.d_in(u_ca_in_566), .d_out(u_ca_out_566));
compressor_81_24 u_ca_81_24_567(.d_in(u_ca_in_567), .d_out(u_ca_out_567));
compressor_81_24 u_ca_81_24_568(.d_in(u_ca_in_568), .d_out(u_ca_out_568));
compressor_81_24 u_ca_81_24_569(.d_in(u_ca_in_569), .d_out(u_ca_out_569));
compressor_81_24 u_ca_81_24_570(.d_in(u_ca_in_570), .d_out(u_ca_out_570));
compressor_81_24 u_ca_81_24_571(.d_in(u_ca_in_571), .d_out(u_ca_out_571));
compressor_81_24 u_ca_81_24_572(.d_in(u_ca_in_572), .d_out(u_ca_out_572));
compressor_81_24 u_ca_81_24_573(.d_in(u_ca_in_573), .d_out(u_ca_out_573));
compressor_81_24 u_ca_81_24_574(.d_in(u_ca_in_574), .d_out(u_ca_out_574));
compressor_81_24 u_ca_81_24_575(.d_in(u_ca_in_575), .d_out(u_ca_out_575));
compressor_81_24 u_ca_81_24_576(.d_in(u_ca_in_576), .d_out(u_ca_out_576));
compressor_81_24 u_ca_81_24_577(.d_in(u_ca_in_577), .d_out(u_ca_out_577));
compressor_81_24 u_ca_81_24_578(.d_in(u_ca_in_578), .d_out(u_ca_out_578));
compressor_81_24 u_ca_81_24_579(.d_in(u_ca_in_579), .d_out(u_ca_out_579));
compressor_81_24 u_ca_81_24_580(.d_in(u_ca_in_580), .d_out(u_ca_out_580));
compressor_81_24 u_ca_81_24_581(.d_in(u_ca_in_581), .d_out(u_ca_out_581));
compressor_81_24 u_ca_81_24_582(.d_in(u_ca_in_582), .d_out(u_ca_out_582));
compressor_81_24 u_ca_81_24_583(.d_in(u_ca_in_583), .d_out(u_ca_out_583));
compressor_81_24 u_ca_81_24_584(.d_in(u_ca_in_584), .d_out(u_ca_out_584));
compressor_81_24 u_ca_81_24_585(.d_in(u_ca_in_585), .d_out(u_ca_out_585));
compressor_81_24 u_ca_81_24_586(.d_in(u_ca_in_586), .d_out(u_ca_out_586));
compressor_81_24 u_ca_81_24_587(.d_in(u_ca_in_587), .d_out(u_ca_out_587));
compressor_81_24 u_ca_81_24_588(.d_in(u_ca_in_588), .d_out(u_ca_out_588));
compressor_81_24 u_ca_81_24_589(.d_in(u_ca_in_589), .d_out(u_ca_out_589));
compressor_81_24 u_ca_81_24_590(.d_in(u_ca_in_590), .d_out(u_ca_out_590));
compressor_81_24 u_ca_81_24_591(.d_in(u_ca_in_591), .d_out(u_ca_out_591));
compressor_81_24 u_ca_81_24_592(.d_in(u_ca_in_592), .d_out(u_ca_out_592));
compressor_81_24 u_ca_81_24_593(.d_in(u_ca_in_593), .d_out(u_ca_out_593));
compressor_81_24 u_ca_81_24_594(.d_in(u_ca_in_594), .d_out(u_ca_out_594));
compressor_81_24 u_ca_81_24_595(.d_in(u_ca_in_595), .d_out(u_ca_out_595));
compressor_81_24 u_ca_81_24_596(.d_in(u_ca_in_596), .d_out(u_ca_out_596));
compressor_81_24 u_ca_81_24_597(.d_in(u_ca_in_597), .d_out(u_ca_out_597));
compressor_81_24 u_ca_81_24_598(.d_in(u_ca_in_598), .d_out(u_ca_out_598));
compressor_81_24 u_ca_81_24_599(.d_in(u_ca_in_599), .d_out(u_ca_out_599));
compressor_81_24 u_ca_81_24_600(.d_in(u_ca_in_600), .d_out(u_ca_out_600));
compressor_81_24 u_ca_81_24_601(.d_in(u_ca_in_601), .d_out(u_ca_out_601));
compressor_81_24 u_ca_81_24_602(.d_in(u_ca_in_602), .d_out(u_ca_out_602));
compressor_81_24 u_ca_81_24_603(.d_in(u_ca_in_603), .d_out(u_ca_out_603));
compressor_81_24 u_ca_81_24_604(.d_in(u_ca_in_604), .d_out(u_ca_out_604));
compressor_81_24 u_ca_81_24_605(.d_in(u_ca_in_605), .d_out(u_ca_out_605));
compressor_81_24 u_ca_81_24_606(.d_in(u_ca_in_606), .d_out(u_ca_out_606));
compressor_81_24 u_ca_81_24_607(.d_in(u_ca_in_607), .d_out(u_ca_out_607));
compressor_81_24 u_ca_81_24_608(.d_in(u_ca_in_608), .d_out(u_ca_out_608));
compressor_81_24 u_ca_81_24_609(.d_in(u_ca_in_609), .d_out(u_ca_out_609));
compressor_81_24 u_ca_81_24_610(.d_in(u_ca_in_610), .d_out(u_ca_out_610));
compressor_81_24 u_ca_81_24_611(.d_in(u_ca_in_611), .d_out(u_ca_out_611));
compressor_81_24 u_ca_81_24_612(.d_in(u_ca_in_612), .d_out(u_ca_out_612));
compressor_81_24 u_ca_81_24_613(.d_in(u_ca_in_613), .d_out(u_ca_out_613));
compressor_81_24 u_ca_81_24_614(.d_in(u_ca_in_614), .d_out(u_ca_out_614));
compressor_81_24 u_ca_81_24_615(.d_in(u_ca_in_615), .d_out(u_ca_out_615));
compressor_81_24 u_ca_81_24_616(.d_in(u_ca_in_616), .d_out(u_ca_out_616));
compressor_81_24 u_ca_81_24_617(.d_in(u_ca_in_617), .d_out(u_ca_out_617));
compressor_81_24 u_ca_81_24_618(.d_in(u_ca_in_618), .d_out(u_ca_out_618));
compressor_81_24 u_ca_81_24_619(.d_in(u_ca_in_619), .d_out(u_ca_out_619));
compressor_81_24 u_ca_81_24_620(.d_in(u_ca_in_620), .d_out(u_ca_out_620));
compressor_81_24 u_ca_81_24_621(.d_in(u_ca_in_621), .d_out(u_ca_out_621));
compressor_81_24 u_ca_81_24_622(.d_in(u_ca_in_622), .d_out(u_ca_out_622));
compressor_81_24 u_ca_81_24_623(.d_in(u_ca_in_623), .d_out(u_ca_out_623));
compressor_81_24 u_ca_81_24_624(.d_in(u_ca_in_624), .d_out(u_ca_out_624));
compressor_81_24 u_ca_81_24_625(.d_in(u_ca_in_625), .d_out(u_ca_out_625));
compressor_81_24 u_ca_81_24_626(.d_in(u_ca_in_626), .d_out(u_ca_out_626));
compressor_81_24 u_ca_81_24_627(.d_in(u_ca_in_627), .d_out(u_ca_out_627));
compressor_81_24 u_ca_81_24_628(.d_in(u_ca_in_628), .d_out(u_ca_out_628));
compressor_81_24 u_ca_81_24_629(.d_in(u_ca_in_629), .d_out(u_ca_out_629));
compressor_81_24 u_ca_81_24_630(.d_in(u_ca_in_630), .d_out(u_ca_out_630));
compressor_81_24 u_ca_81_24_631(.d_in(u_ca_in_631), .d_out(u_ca_out_631));
compressor_81_24 u_ca_81_24_632(.d_in(u_ca_in_632), .d_out(u_ca_out_632));
compressor_81_24 u_ca_81_24_633(.d_in(u_ca_in_633), .d_out(u_ca_out_633));
compressor_81_24 u_ca_81_24_634(.d_in(u_ca_in_634), .d_out(u_ca_out_634));
compressor_81_24 u_ca_81_24_635(.d_in(u_ca_in_635), .d_out(u_ca_out_635));
compressor_81_24 u_ca_81_24_636(.d_in(u_ca_in_636), .d_out(u_ca_out_636));
compressor_81_24 u_ca_81_24_637(.d_in(u_ca_in_637), .d_out(u_ca_out_637));
compressor_81_24 u_ca_81_24_638(.d_in(u_ca_in_638), .d_out(u_ca_out_638));
compressor_81_24 u_ca_81_24_639(.d_in(u_ca_in_639), .d_out(u_ca_out_639));
compressor_81_24 u_ca_81_24_640(.d_in(u_ca_in_640), .d_out(u_ca_out_640));
compressor_81_24 u_ca_81_24_641(.d_in(u_ca_in_641), .d_out(u_ca_out_641));
compressor_81_24 u_ca_81_24_642(.d_in(u_ca_in_642), .d_out(u_ca_out_642));
compressor_81_24 u_ca_81_24_643(.d_in(u_ca_in_643), .d_out(u_ca_out_643));
compressor_81_24 u_ca_81_24_644(.d_in(u_ca_in_644), .d_out(u_ca_out_644));
compressor_81_24 u_ca_81_24_645(.d_in(u_ca_in_645), .d_out(u_ca_out_645));
compressor_81_24 u_ca_81_24_646(.d_in(u_ca_in_646), .d_out(u_ca_out_646));
compressor_81_24 u_ca_81_24_647(.d_in(u_ca_in_647), .d_out(u_ca_out_647));
compressor_81_24 u_ca_81_24_648(.d_in(u_ca_in_648), .d_out(u_ca_out_648));
compressor_81_24 u_ca_81_24_649(.d_in(u_ca_in_649), .d_out(u_ca_out_649));
compressor_81_24 u_ca_81_24_650(.d_in(u_ca_in_650), .d_out(u_ca_out_650));
compressor_81_24 u_ca_81_24_651(.d_in(u_ca_in_651), .d_out(u_ca_out_651));
compressor_81_24 u_ca_81_24_652(.d_in(u_ca_in_652), .d_out(u_ca_out_652));
compressor_81_24 u_ca_81_24_653(.d_in(u_ca_in_653), .d_out(u_ca_out_653));
compressor_81_24 u_ca_81_24_654(.d_in(u_ca_in_654), .d_out(u_ca_out_654));
compressor_81_24 u_ca_81_24_655(.d_in(u_ca_in_655), .d_out(u_ca_out_655));
compressor_81_24 u_ca_81_24_656(.d_in(u_ca_in_656), .d_out(u_ca_out_656));
compressor_81_24 u_ca_81_24_657(.d_in(u_ca_in_657), .d_out(u_ca_out_657));
compressor_81_24 u_ca_81_24_658(.d_in(u_ca_in_658), .d_out(u_ca_out_658));
compressor_81_24 u_ca_81_24_659(.d_in(u_ca_in_659), .d_out(u_ca_out_659));
compressor_81_24 u_ca_81_24_660(.d_in(u_ca_in_660), .d_out(u_ca_out_660));
compressor_81_24 u_ca_81_24_661(.d_in(u_ca_in_661), .d_out(u_ca_out_661));
compressor_81_24 u_ca_81_24_662(.d_in(u_ca_in_662), .d_out(u_ca_out_662));
compressor_81_24 u_ca_81_24_663(.d_in(u_ca_in_663), .d_out(u_ca_out_663));
compressor_81_24 u_ca_81_24_664(.d_in(u_ca_in_664), .d_out(u_ca_out_664));
compressor_81_24 u_ca_81_24_665(.d_in(u_ca_in_665), .d_out(u_ca_out_665));
compressor_81_24 u_ca_81_24_666(.d_in(u_ca_in_666), .d_out(u_ca_out_666));
compressor_81_24 u_ca_81_24_667(.d_in(u_ca_in_667), .d_out(u_ca_out_667));
compressor_81_24 u_ca_81_24_668(.d_in(u_ca_in_668), .d_out(u_ca_out_668));
compressor_81_24 u_ca_81_24_669(.d_in(u_ca_in_669), .d_out(u_ca_out_669));
compressor_81_24 u_ca_81_24_670(.d_in(u_ca_in_670), .d_out(u_ca_out_670));
compressor_81_24 u_ca_81_24_671(.d_in(u_ca_in_671), .d_out(u_ca_out_671));
compressor_81_24 u_ca_81_24_672(.d_in(u_ca_in_672), .d_out(u_ca_out_672));
compressor_81_24 u_ca_81_24_673(.d_in(u_ca_in_673), .d_out(u_ca_out_673));
compressor_81_24 u_ca_81_24_674(.d_in(u_ca_in_674), .d_out(u_ca_out_674));
compressor_81_24 u_ca_81_24_675(.d_in(u_ca_in_675), .d_out(u_ca_out_675));
compressor_81_24 u_ca_81_24_676(.d_in(u_ca_in_676), .d_out(u_ca_out_676));
compressor_81_24 u_ca_81_24_677(.d_in(u_ca_in_677), .d_out(u_ca_out_677));
compressor_81_24 u_ca_81_24_678(.d_in(u_ca_in_678), .d_out(u_ca_out_678));
compressor_81_24 u_ca_81_24_679(.d_in(u_ca_in_679), .d_out(u_ca_out_679));
compressor_81_24 u_ca_81_24_680(.d_in(u_ca_in_680), .d_out(u_ca_out_680));
compressor_81_24 u_ca_81_24_681(.d_in(u_ca_in_681), .d_out(u_ca_out_681));
compressor_81_24 u_ca_81_24_682(.d_in(u_ca_in_682), .d_out(u_ca_out_682));
compressor_81_24 u_ca_81_24_683(.d_in(u_ca_in_683), .d_out(u_ca_out_683));
compressor_81_24 u_ca_81_24_684(.d_in(u_ca_in_684), .d_out(u_ca_out_684));
compressor_81_24 u_ca_81_24_685(.d_in(u_ca_in_685), .d_out(u_ca_out_685));
compressor_81_24 u_ca_81_24_686(.d_in(u_ca_in_686), .d_out(u_ca_out_686));
compressor_81_24 u_ca_81_24_687(.d_in(u_ca_in_687), .d_out(u_ca_out_687));
compressor_81_24 u_ca_81_24_688(.d_in(u_ca_in_688), .d_out(u_ca_out_688));
compressor_81_24 u_ca_81_24_689(.d_in(u_ca_in_689), .d_out(u_ca_out_689));
compressor_81_24 u_ca_81_24_690(.d_in(u_ca_in_690), .d_out(u_ca_out_690));
compressor_81_24 u_ca_81_24_691(.d_in(u_ca_in_691), .d_out(u_ca_out_691));
compressor_81_24 u_ca_81_24_692(.d_in(u_ca_in_692), .d_out(u_ca_out_692));
compressor_81_24 u_ca_81_24_693(.d_in(u_ca_in_693), .d_out(u_ca_out_693));
compressor_81_24 u_ca_81_24_694(.d_in(u_ca_in_694), .d_out(u_ca_out_694));
compressor_81_24 u_ca_81_24_695(.d_in(u_ca_in_695), .d_out(u_ca_out_695));
compressor_81_24 u_ca_81_24_696(.d_in(u_ca_in_696), .d_out(u_ca_out_696));
compressor_81_24 u_ca_81_24_697(.d_in(u_ca_in_697), .d_out(u_ca_out_697));
compressor_81_24 u_ca_81_24_698(.d_in(u_ca_in_698), .d_out(u_ca_out_698));
compressor_81_24 u_ca_81_24_699(.d_in(u_ca_in_699), .d_out(u_ca_out_699));
compressor_81_24 u_ca_81_24_700(.d_in(u_ca_in_700), .d_out(u_ca_out_700));
compressor_81_24 u_ca_81_24_701(.d_in(u_ca_in_701), .d_out(u_ca_out_701));
compressor_81_24 u_ca_81_24_702(.d_in(u_ca_in_702), .d_out(u_ca_out_702));
compressor_81_24 u_ca_81_24_703(.d_in(u_ca_in_703), .d_out(u_ca_out_703));
compressor_81_24 u_ca_81_24_704(.d_in(u_ca_in_704), .d_out(u_ca_out_704));
compressor_81_24 u_ca_81_24_705(.d_in(u_ca_in_705), .d_out(u_ca_out_705));
compressor_81_24 u_ca_81_24_706(.d_in(u_ca_in_706), .d_out(u_ca_out_706));
compressor_81_24 u_ca_81_24_707(.d_in(u_ca_in_707), .d_out(u_ca_out_707));
compressor_81_24 u_ca_81_24_708(.d_in(u_ca_in_708), .d_out(u_ca_out_708));
compressor_81_24 u_ca_81_24_709(.d_in(u_ca_in_709), .d_out(u_ca_out_709));
compressor_81_24 u_ca_81_24_710(.d_in(u_ca_in_710), .d_out(u_ca_out_710));
compressor_81_24 u_ca_81_24_711(.d_in(u_ca_in_711), .d_out(u_ca_out_711));
compressor_81_24 u_ca_81_24_712(.d_in(u_ca_in_712), .d_out(u_ca_out_712));
compressor_81_24 u_ca_81_24_713(.d_in(u_ca_in_713), .d_out(u_ca_out_713));
compressor_81_24 u_ca_81_24_714(.d_in(u_ca_in_714), .d_out(u_ca_out_714));
compressor_81_24 u_ca_81_24_715(.d_in(u_ca_in_715), .d_out(u_ca_out_715));
compressor_81_24 u_ca_81_24_716(.d_in(u_ca_in_716), .d_out(u_ca_out_716));
compressor_81_24 u_ca_81_24_717(.d_in(u_ca_in_717), .d_out(u_ca_out_717));
compressor_81_24 u_ca_81_24_718(.d_in(u_ca_in_718), .d_out(u_ca_out_718));
compressor_81_24 u_ca_81_24_719(.d_in(u_ca_in_719), .d_out(u_ca_out_719));
compressor_81_24 u_ca_81_24_720(.d_in(u_ca_in_720), .d_out(u_ca_out_720));
compressor_81_24 u_ca_81_24_721(.d_in(u_ca_in_721), .d_out(u_ca_out_721));
compressor_81_24 u_ca_81_24_722(.d_in(u_ca_in_722), .d_out(u_ca_out_722));
compressor_81_24 u_ca_81_24_723(.d_in(u_ca_in_723), .d_out(u_ca_out_723));
compressor_81_24 u_ca_81_24_724(.d_in(u_ca_in_724), .d_out(u_ca_out_724));
compressor_81_24 u_ca_81_24_725(.d_in(u_ca_in_725), .d_out(u_ca_out_725));
compressor_81_24 u_ca_81_24_726(.d_in(u_ca_in_726), .d_out(u_ca_out_726));
compressor_81_24 u_ca_81_24_727(.d_in(u_ca_in_727), .d_out(u_ca_out_727));
compressor_81_24 u_ca_81_24_728(.d_in(u_ca_in_728), .d_out(u_ca_out_728));
compressor_81_24 u_ca_81_24_729(.d_in(u_ca_in_729), .d_out(u_ca_out_729));
compressor_81_24 u_ca_81_24_730(.d_in(u_ca_in_730), .d_out(u_ca_out_730));
compressor_81_24 u_ca_81_24_731(.d_in(u_ca_in_731), .d_out(u_ca_out_731));
compressor_81_24 u_ca_81_24_732(.d_in(u_ca_in_732), .d_out(u_ca_out_732));
compressor_81_24 u_ca_81_24_733(.d_in(u_ca_in_733), .d_out(u_ca_out_733));
compressor_81_24 u_ca_81_24_734(.d_in(u_ca_in_734), .d_out(u_ca_out_734));
compressor_81_24 u_ca_81_24_735(.d_in(u_ca_in_735), .d_out(u_ca_out_735));
compressor_81_24 u_ca_81_24_736(.d_in(u_ca_in_736), .d_out(u_ca_out_736));
compressor_81_24 u_ca_81_24_737(.d_in(u_ca_in_737), .d_out(u_ca_out_737));
compressor_81_24 u_ca_81_24_738(.d_in(u_ca_in_738), .d_out(u_ca_out_738));
compressor_81_24 u_ca_81_24_739(.d_in(u_ca_in_739), .d_out(u_ca_out_739));
compressor_81_24 u_ca_81_24_740(.d_in(u_ca_in_740), .d_out(u_ca_out_740));
compressor_81_24 u_ca_81_24_741(.d_in(u_ca_in_741), .d_out(u_ca_out_741));
compressor_81_24 u_ca_81_24_742(.d_in(u_ca_in_742), .d_out(u_ca_out_742));
compressor_81_24 u_ca_81_24_743(.d_in(u_ca_in_743), .d_out(u_ca_out_743));
compressor_81_24 u_ca_81_24_744(.d_in(u_ca_in_744), .d_out(u_ca_out_744));
compressor_81_24 u_ca_81_24_745(.d_in(u_ca_in_745), .d_out(u_ca_out_745));
compressor_81_24 u_ca_81_24_746(.d_in(u_ca_in_746), .d_out(u_ca_out_746));
compressor_81_24 u_ca_81_24_747(.d_in(u_ca_in_747), .d_out(u_ca_out_747));
compressor_81_24 u_ca_81_24_748(.d_in(u_ca_in_748), .d_out(u_ca_out_748));
compressor_81_24 u_ca_81_24_749(.d_in(u_ca_in_749), .d_out(u_ca_out_749));
compressor_81_24 u_ca_81_24_750(.d_in(u_ca_in_750), .d_out(u_ca_out_750));
compressor_81_24 u_ca_81_24_751(.d_in(u_ca_in_751), .d_out(u_ca_out_751));
compressor_81_24 u_ca_81_24_752(.d_in(u_ca_in_752), .d_out(u_ca_out_752));
compressor_81_24 u_ca_81_24_753(.d_in(u_ca_in_753), .d_out(u_ca_out_753));
compressor_81_24 u_ca_81_24_754(.d_in(u_ca_in_754), .d_out(u_ca_out_754));
compressor_81_24 u_ca_81_24_755(.d_in(u_ca_in_755), .d_out(u_ca_out_755));
compressor_81_24 u_ca_81_24_756(.d_in(u_ca_in_756), .d_out(u_ca_out_756));
compressor_81_24 u_ca_81_24_757(.d_in(u_ca_in_757), .d_out(u_ca_out_757));
compressor_81_24 u_ca_81_24_758(.d_in(u_ca_in_758), .d_out(u_ca_out_758));
compressor_81_24 u_ca_81_24_759(.d_in(u_ca_in_759), .d_out(u_ca_out_759));
compressor_81_24 u_ca_81_24_760(.d_in(u_ca_in_760), .d_out(u_ca_out_760));
compressor_81_24 u_ca_81_24_761(.d_in(u_ca_in_761), .d_out(u_ca_out_761));
compressor_81_24 u_ca_81_24_762(.d_in(u_ca_in_762), .d_out(u_ca_out_762));
compressor_81_24 u_ca_81_24_763(.d_in(u_ca_in_763), .d_out(u_ca_out_763));
compressor_81_24 u_ca_81_24_764(.d_in(u_ca_in_764), .d_out(u_ca_out_764));
compressor_81_24 u_ca_81_24_765(.d_in(u_ca_in_765), .d_out(u_ca_out_765));
compressor_81_24 u_ca_81_24_766(.d_in(u_ca_in_766), .d_out(u_ca_out_766));
compressor_81_24 u_ca_81_24_767(.d_in(u_ca_in_767), .d_out(u_ca_out_767));
compressor_81_24 u_ca_81_24_768(.d_in(u_ca_in_768), .d_out(u_ca_out_768));
compressor_81_24 u_ca_81_24_769(.d_in(u_ca_in_769), .d_out(u_ca_out_769));
compressor_81_24 u_ca_81_24_770(.d_in(u_ca_in_770), .d_out(u_ca_out_770));
compressor_81_24 u_ca_81_24_771(.d_in(u_ca_in_771), .d_out(u_ca_out_771));
compressor_81_24 u_ca_81_24_772(.d_in(u_ca_in_772), .d_out(u_ca_out_772));
compressor_81_24 u_ca_81_24_773(.d_in(u_ca_in_773), .d_out(u_ca_out_773));
compressor_81_24 u_ca_81_24_774(.d_in(u_ca_in_774), .d_out(u_ca_out_774));
compressor_81_24 u_ca_81_24_775(.d_in(u_ca_in_775), .d_out(u_ca_out_775));
compressor_81_24 u_ca_81_24_776(.d_in(u_ca_in_776), .d_out(u_ca_out_776));
compressor_81_24 u_ca_81_24_777(.d_in(u_ca_in_777), .d_out(u_ca_out_777));
compressor_81_24 u_ca_81_24_778(.d_in(u_ca_in_778), .d_out(u_ca_out_778));
compressor_81_24 u_ca_81_24_779(.d_in(u_ca_in_779), .d_out(u_ca_out_779));
compressor_81_24 u_ca_81_24_780(.d_in(u_ca_in_780), .d_out(u_ca_out_780));
compressor_81_24 u_ca_81_24_781(.d_in(u_ca_in_781), .d_out(u_ca_out_781));
compressor_81_24 u_ca_81_24_782(.d_in(u_ca_in_782), .d_out(u_ca_out_782));
compressor_81_24 u_ca_81_24_783(.d_in(u_ca_in_783), .d_out(u_ca_out_783));
compressor_81_24 u_ca_81_24_784(.d_in(u_ca_in_784), .d_out(u_ca_out_784));
compressor_81_24 u_ca_81_24_785(.d_in(u_ca_in_785), .d_out(u_ca_out_785));
compressor_81_24 u_ca_81_24_786(.d_in(u_ca_in_786), .d_out(u_ca_out_786));
compressor_81_24 u_ca_81_24_787(.d_in(u_ca_in_787), .d_out(u_ca_out_787));
compressor_81_24 u_ca_81_24_788(.d_in(u_ca_in_788), .d_out(u_ca_out_788));
compressor_81_24 u_ca_81_24_789(.d_in(u_ca_in_789), .d_out(u_ca_out_789));
compressor_81_24 u_ca_81_24_790(.d_in(u_ca_in_790), .d_out(u_ca_out_790));
compressor_81_24 u_ca_81_24_791(.d_in(u_ca_in_791), .d_out(u_ca_out_791));
compressor_81_24 u_ca_81_24_792(.d_in(u_ca_in_792), .d_out(u_ca_out_792));
compressor_81_24 u_ca_81_24_793(.d_in(u_ca_in_793), .d_out(u_ca_out_793));
compressor_81_24 u_ca_81_24_794(.d_in(u_ca_in_794), .d_out(u_ca_out_794));
compressor_81_24 u_ca_81_24_795(.d_in(u_ca_in_795), .d_out(u_ca_out_795));
compressor_81_24 u_ca_81_24_796(.d_in(u_ca_in_796), .d_out(u_ca_out_796));
compressor_81_24 u_ca_81_24_797(.d_in(u_ca_in_797), .d_out(u_ca_out_797));
compressor_81_24 u_ca_81_24_798(.d_in(u_ca_in_798), .d_out(u_ca_out_798));
compressor_81_24 u_ca_81_24_799(.d_in(u_ca_in_799), .d_out(u_ca_out_799));
compressor_81_24 u_ca_81_24_800(.d_in(u_ca_in_800), .d_out(u_ca_out_800));
compressor_81_24 u_ca_81_24_801(.d_in(u_ca_in_801), .d_out(u_ca_out_801));
compressor_81_24 u_ca_81_24_802(.d_in(u_ca_in_802), .d_out(u_ca_out_802));
compressor_81_24 u_ca_81_24_803(.d_in(u_ca_in_803), .d_out(u_ca_out_803));
compressor_81_24 u_ca_81_24_804(.d_in(u_ca_in_804), .d_out(u_ca_out_804));
compressor_81_24 u_ca_81_24_805(.d_in(u_ca_in_805), .d_out(u_ca_out_805));
compressor_81_24 u_ca_81_24_806(.d_in(u_ca_in_806), .d_out(u_ca_out_806));
compressor_81_24 u_ca_81_24_807(.d_in(u_ca_in_807), .d_out(u_ca_out_807));
compressor_81_24 u_ca_81_24_808(.d_in(u_ca_in_808), .d_out(u_ca_out_808));
compressor_81_24 u_ca_81_24_809(.d_in(u_ca_in_809), .d_out(u_ca_out_809));
compressor_81_24 u_ca_81_24_810(.d_in(u_ca_in_810), .d_out(u_ca_out_810));
compressor_81_24 u_ca_81_24_811(.d_in(u_ca_in_811), .d_out(u_ca_out_811));
compressor_81_24 u_ca_81_24_812(.d_in(u_ca_in_812), .d_out(u_ca_out_812));
compressor_81_24 u_ca_81_24_813(.d_in(u_ca_in_813), .d_out(u_ca_out_813));
compressor_81_24 u_ca_81_24_814(.d_in(u_ca_in_814), .d_out(u_ca_out_814));
compressor_81_24 u_ca_81_24_815(.d_in(u_ca_in_815), .d_out(u_ca_out_815));
compressor_81_24 u_ca_81_24_816(.d_in(u_ca_in_816), .d_out(u_ca_out_816));
compressor_81_24 u_ca_81_24_817(.d_in(u_ca_in_817), .d_out(u_ca_out_817));
compressor_81_24 u_ca_81_24_818(.d_in(u_ca_in_818), .d_out(u_ca_out_818));
compressor_81_24 u_ca_81_24_819(.d_in(u_ca_in_819), .d_out(u_ca_out_819));
compressor_81_24 u_ca_81_24_820(.d_in(u_ca_in_820), .d_out(u_ca_out_820));
compressor_81_24 u_ca_81_24_821(.d_in(u_ca_in_821), .d_out(u_ca_out_821));
compressor_81_24 u_ca_81_24_822(.d_in(u_ca_in_822), .d_out(u_ca_out_822));
compressor_81_24 u_ca_81_24_823(.d_in(u_ca_in_823), .d_out(u_ca_out_823));
compressor_81_24 u_ca_81_24_824(.d_in(u_ca_in_824), .d_out(u_ca_out_824));
compressor_81_24 u_ca_81_24_825(.d_in(u_ca_in_825), .d_out(u_ca_out_825));
compressor_81_24 u_ca_81_24_826(.d_in(u_ca_in_826), .d_out(u_ca_out_826));
compressor_81_24 u_ca_81_24_827(.d_in(u_ca_in_827), .d_out(u_ca_out_827));
compressor_81_24 u_ca_81_24_828(.d_in(u_ca_in_828), .d_out(u_ca_out_828));
compressor_81_24 u_ca_81_24_829(.d_in(u_ca_in_829), .d_out(u_ca_out_829));
compressor_81_24 u_ca_81_24_830(.d_in(u_ca_in_830), .d_out(u_ca_out_830));
compressor_81_24 u_ca_81_24_831(.d_in(u_ca_in_831), .d_out(u_ca_out_831));
compressor_81_24 u_ca_81_24_832(.d_in(u_ca_in_832), .d_out(u_ca_out_832));
compressor_81_24 u_ca_81_24_833(.d_in(u_ca_in_833), .d_out(u_ca_out_833));
compressor_81_24 u_ca_81_24_834(.d_in(u_ca_in_834), .d_out(u_ca_out_834));
compressor_81_24 u_ca_81_24_835(.d_in(u_ca_in_835), .d_out(u_ca_out_835));
compressor_81_24 u_ca_81_24_836(.d_in(u_ca_in_836), .d_out(u_ca_out_836));
compressor_81_24 u_ca_81_24_837(.d_in(u_ca_in_837), .d_out(u_ca_out_837));
compressor_81_24 u_ca_81_24_838(.d_in(u_ca_in_838), .d_out(u_ca_out_838));
compressor_81_24 u_ca_81_24_839(.d_in(u_ca_in_839), .d_out(u_ca_out_839));
compressor_81_24 u_ca_81_24_840(.d_in(u_ca_in_840), .d_out(u_ca_out_840));
compressor_81_24 u_ca_81_24_841(.d_in(u_ca_in_841), .d_out(u_ca_out_841));
compressor_81_24 u_ca_81_24_842(.d_in(u_ca_in_842), .d_out(u_ca_out_842));
compressor_81_24 u_ca_81_24_843(.d_in(u_ca_in_843), .d_out(u_ca_out_843));
compressor_81_24 u_ca_81_24_844(.d_in(u_ca_in_844), .d_out(u_ca_out_844));
compressor_81_24 u_ca_81_24_845(.d_in(u_ca_in_845), .d_out(u_ca_out_845));
compressor_81_24 u_ca_81_24_846(.d_in(u_ca_in_846), .d_out(u_ca_out_846));
compressor_81_24 u_ca_81_24_847(.d_in(u_ca_in_847), .d_out(u_ca_out_847));
compressor_81_24 u_ca_81_24_848(.d_in(u_ca_in_848), .d_out(u_ca_out_848));
compressor_81_24 u_ca_81_24_849(.d_in(u_ca_in_849), .d_out(u_ca_out_849));
compressor_81_24 u_ca_81_24_850(.d_in(u_ca_in_850), .d_out(u_ca_out_850));
compressor_81_24 u_ca_81_24_851(.d_in(u_ca_in_851), .d_out(u_ca_out_851));
compressor_81_24 u_ca_81_24_852(.d_in(u_ca_in_852), .d_out(u_ca_out_852));
compressor_81_24 u_ca_81_24_853(.d_in(u_ca_in_853), .d_out(u_ca_out_853));
compressor_81_24 u_ca_81_24_854(.d_in(u_ca_in_854), .d_out(u_ca_out_854));
compressor_81_24 u_ca_81_24_855(.d_in(u_ca_in_855), .d_out(u_ca_out_855));
compressor_81_24 u_ca_81_24_856(.d_in(u_ca_in_856), .d_out(u_ca_out_856));
compressor_81_24 u_ca_81_24_857(.d_in(u_ca_in_857), .d_out(u_ca_out_857));
compressor_81_24 u_ca_81_24_858(.d_in(u_ca_in_858), .d_out(u_ca_out_858));
compressor_81_24 u_ca_81_24_859(.d_in(u_ca_in_859), .d_out(u_ca_out_859));
compressor_81_24 u_ca_81_24_860(.d_in(u_ca_in_860), .d_out(u_ca_out_860));
compressor_81_24 u_ca_81_24_861(.d_in(u_ca_in_861), .d_out(u_ca_out_861));
compressor_81_24 u_ca_81_24_862(.d_in(u_ca_in_862), .d_out(u_ca_out_862));
compressor_81_24 u_ca_81_24_863(.d_in(u_ca_in_863), .d_out(u_ca_out_863));
compressor_81_24 u_ca_81_24_864(.d_in(u_ca_in_864), .d_out(u_ca_out_864));
compressor_81_24 u_ca_81_24_865(.d_in(u_ca_in_865), .d_out(u_ca_out_865));
compressor_81_24 u_ca_81_24_866(.d_in(u_ca_in_866), .d_out(u_ca_out_866));
compressor_81_24 u_ca_81_24_867(.d_in(u_ca_in_867), .d_out(u_ca_out_867));
compressor_81_24 u_ca_81_24_868(.d_in(u_ca_in_868), .d_out(u_ca_out_868));
compressor_81_24 u_ca_81_24_869(.d_in(u_ca_in_869), .d_out(u_ca_out_869));
compressor_81_24 u_ca_81_24_870(.d_in(u_ca_in_870), .d_out(u_ca_out_870));
compressor_81_24 u_ca_81_24_871(.d_in(u_ca_in_871), .d_out(u_ca_out_871));
compressor_81_24 u_ca_81_24_872(.d_in(u_ca_in_872), .d_out(u_ca_out_872));
compressor_81_24 u_ca_81_24_873(.d_in(u_ca_in_873), .d_out(u_ca_out_873));
compressor_81_24 u_ca_81_24_874(.d_in(u_ca_in_874), .d_out(u_ca_out_874));
compressor_81_24 u_ca_81_24_875(.d_in(u_ca_in_875), .d_out(u_ca_out_875));
compressor_81_24 u_ca_81_24_876(.d_in(u_ca_in_876), .d_out(u_ca_out_876));
compressor_81_24 u_ca_81_24_877(.d_in(u_ca_in_877), .d_out(u_ca_out_877));
compressor_81_24 u_ca_81_24_878(.d_in(u_ca_in_878), .d_out(u_ca_out_878));
compressor_81_24 u_ca_81_24_879(.d_in(u_ca_in_879), .d_out(u_ca_out_879));
compressor_81_24 u_ca_81_24_880(.d_in(u_ca_in_880), .d_out(u_ca_out_880));
compressor_81_24 u_ca_81_24_881(.d_in(u_ca_in_881), .d_out(u_ca_out_881));
compressor_81_24 u_ca_81_24_882(.d_in(u_ca_in_882), .d_out(u_ca_out_882));
compressor_81_24 u_ca_81_24_883(.d_in(u_ca_in_883), .d_out(u_ca_out_883));
compressor_81_24 u_ca_81_24_884(.d_in(u_ca_in_884), .d_out(u_ca_out_884));
compressor_81_24 u_ca_81_24_885(.d_in(u_ca_in_885), .d_out(u_ca_out_885));
compressor_81_24 u_ca_81_24_886(.d_in(u_ca_in_886), .d_out(u_ca_out_886));
compressor_81_24 u_ca_81_24_887(.d_in(u_ca_in_887), .d_out(u_ca_out_887));
compressor_81_24 u_ca_81_24_888(.d_in(u_ca_in_888), .d_out(u_ca_out_888));
compressor_81_24 u_ca_81_24_889(.d_in(u_ca_in_889), .d_out(u_ca_out_889));
compressor_81_24 u_ca_81_24_890(.d_in(u_ca_in_890), .d_out(u_ca_out_890));
compressor_81_24 u_ca_81_24_891(.d_in(u_ca_in_891), .d_out(u_ca_out_891));
compressor_81_24 u_ca_81_24_892(.d_in(u_ca_in_892), .d_out(u_ca_out_892));
compressor_81_24 u_ca_81_24_893(.d_in(u_ca_in_893), .d_out(u_ca_out_893));
compressor_81_24 u_ca_81_24_894(.d_in(u_ca_in_894), .d_out(u_ca_out_894));
compressor_81_24 u_ca_81_24_895(.d_in(u_ca_in_895), .d_out(u_ca_out_895));
compressor_81_24 u_ca_81_24_896(.d_in(u_ca_in_896), .d_out(u_ca_out_896));
compressor_81_24 u_ca_81_24_897(.d_in(u_ca_in_897), .d_out(u_ca_out_897));
compressor_81_24 u_ca_81_24_898(.d_in(u_ca_in_898), .d_out(u_ca_out_898));
compressor_81_24 u_ca_81_24_899(.d_in(u_ca_in_899), .d_out(u_ca_out_899));
compressor_81_24 u_ca_81_24_900(.d_in(u_ca_in_900), .d_out(u_ca_out_900));
compressor_81_24 u_ca_81_24_901(.d_in(u_ca_in_901), .d_out(u_ca_out_901));
compressor_81_24 u_ca_81_24_902(.d_in(u_ca_in_902), .d_out(u_ca_out_902));
compressor_81_24 u_ca_81_24_903(.d_in(u_ca_in_903), .d_out(u_ca_out_903));
compressor_81_24 u_ca_81_24_904(.d_in(u_ca_in_904), .d_out(u_ca_out_904));
compressor_81_24 u_ca_81_24_905(.d_in(u_ca_in_905), .d_out(u_ca_out_905));
compressor_81_24 u_ca_81_24_906(.d_in(u_ca_in_906), .d_out(u_ca_out_906));
compressor_81_24 u_ca_81_24_907(.d_in(u_ca_in_907), .d_out(u_ca_out_907));
compressor_81_24 u_ca_81_24_908(.d_in(u_ca_in_908), .d_out(u_ca_out_908));
compressor_81_24 u_ca_81_24_909(.d_in(u_ca_in_909), .d_out(u_ca_out_909));
compressor_81_24 u_ca_81_24_910(.d_in(u_ca_in_910), .d_out(u_ca_out_910));
compressor_81_24 u_ca_81_24_911(.d_in(u_ca_in_911), .d_out(u_ca_out_911));
compressor_81_24 u_ca_81_24_912(.d_in(u_ca_in_912), .d_out(u_ca_out_912));
compressor_81_24 u_ca_81_24_913(.d_in(u_ca_in_913), .d_out(u_ca_out_913));
compressor_81_24 u_ca_81_24_914(.d_in(u_ca_in_914), .d_out(u_ca_out_914));
compressor_81_24 u_ca_81_24_915(.d_in(u_ca_in_915), .d_out(u_ca_out_915));
compressor_81_24 u_ca_81_24_916(.d_in(u_ca_in_916), .d_out(u_ca_out_916));
compressor_81_24 u_ca_81_24_917(.d_in(u_ca_in_917), .d_out(u_ca_out_917));
compressor_81_24 u_ca_81_24_918(.d_in(u_ca_in_918), .d_out(u_ca_out_918));
compressor_81_24 u_ca_81_24_919(.d_in(u_ca_in_919), .d_out(u_ca_out_919));
compressor_81_24 u_ca_81_24_920(.d_in(u_ca_in_920), .d_out(u_ca_out_920));
compressor_81_24 u_ca_81_24_921(.d_in(u_ca_in_921), .d_out(u_ca_out_921));
compressor_81_24 u_ca_81_24_922(.d_in(u_ca_in_922), .d_out(u_ca_out_922));
compressor_81_24 u_ca_81_24_923(.d_in(u_ca_in_923), .d_out(u_ca_out_923));
compressor_81_24 u_ca_81_24_924(.d_in(u_ca_in_924), .d_out(u_ca_out_924));
compressor_81_24 u_ca_81_24_925(.d_in(u_ca_in_925), .d_out(u_ca_out_925));
compressor_81_24 u_ca_81_24_926(.d_in(u_ca_in_926), .d_out(u_ca_out_926));
compressor_81_24 u_ca_81_24_927(.d_in(u_ca_in_927), .d_out(u_ca_out_927));
compressor_81_24 u_ca_81_24_928(.d_in(u_ca_in_928), .d_out(u_ca_out_928));
compressor_81_24 u_ca_81_24_929(.d_in(u_ca_in_929), .d_out(u_ca_out_929));
compressor_81_24 u_ca_81_24_930(.d_in(u_ca_in_930), .d_out(u_ca_out_930));
compressor_81_24 u_ca_81_24_931(.d_in(u_ca_in_931), .d_out(u_ca_out_931));
compressor_81_24 u_ca_81_24_932(.d_in(u_ca_in_932), .d_out(u_ca_out_932));
compressor_81_24 u_ca_81_24_933(.d_in(u_ca_in_933), .d_out(u_ca_out_933));
compressor_81_24 u_ca_81_24_934(.d_in(u_ca_in_934), .d_out(u_ca_out_934));
compressor_81_24 u_ca_81_24_935(.d_in(u_ca_in_935), .d_out(u_ca_out_935));
compressor_81_24 u_ca_81_24_936(.d_in(u_ca_in_936), .d_out(u_ca_out_936));
compressor_81_24 u_ca_81_24_937(.d_in(u_ca_in_937), .d_out(u_ca_out_937));
compressor_81_24 u_ca_81_24_938(.d_in(u_ca_in_938), .d_out(u_ca_out_938));
compressor_81_24 u_ca_81_24_939(.d_in(u_ca_in_939), .d_out(u_ca_out_939));
compressor_81_24 u_ca_81_24_940(.d_in(u_ca_in_940), .d_out(u_ca_out_940));
compressor_81_24 u_ca_81_24_941(.d_in(u_ca_in_941), .d_out(u_ca_out_941));
compressor_81_24 u_ca_81_24_942(.d_in(u_ca_in_942), .d_out(u_ca_out_942));
compressor_81_24 u_ca_81_24_943(.d_in(u_ca_in_943), .d_out(u_ca_out_943));
compressor_81_24 u_ca_81_24_944(.d_in(u_ca_in_944), .d_out(u_ca_out_944));
compressor_81_24 u_ca_81_24_945(.d_in(u_ca_in_945), .d_out(u_ca_out_945));
compressor_81_24 u_ca_81_24_946(.d_in(u_ca_in_946), .d_out(u_ca_out_946));
compressor_81_24 u_ca_81_24_947(.d_in(u_ca_in_947), .d_out(u_ca_out_947));
compressor_81_24 u_ca_81_24_948(.d_in(u_ca_in_948), .d_out(u_ca_out_948));
compressor_81_24 u_ca_81_24_949(.d_in(u_ca_in_949), .d_out(u_ca_out_949));
compressor_81_24 u_ca_81_24_950(.d_in(u_ca_in_950), .d_out(u_ca_out_950));
compressor_81_24 u_ca_81_24_951(.d_in(u_ca_in_951), .d_out(u_ca_out_951));
compressor_81_24 u_ca_81_24_952(.d_in(u_ca_in_952), .d_out(u_ca_out_952));
compressor_81_24 u_ca_81_24_953(.d_in(u_ca_in_953), .d_out(u_ca_out_953));
compressor_81_24 u_ca_81_24_954(.d_in(u_ca_in_954), .d_out(u_ca_out_954));
compressor_81_24 u_ca_81_24_955(.d_in(u_ca_in_955), .d_out(u_ca_out_955));
compressor_81_24 u_ca_81_24_956(.d_in(u_ca_in_956), .d_out(u_ca_out_956));
compressor_81_24 u_ca_81_24_957(.d_in(u_ca_in_957), .d_out(u_ca_out_957));
compressor_81_24 u_ca_81_24_958(.d_in(u_ca_in_958), .d_out(u_ca_out_958));
compressor_81_24 u_ca_81_24_959(.d_in(u_ca_in_959), .d_out(u_ca_out_959));
compressor_81_24 u_ca_81_24_960(.d_in(u_ca_in_960), .d_out(u_ca_out_960));
compressor_81_24 u_ca_81_24_961(.d_in(u_ca_in_961), .d_out(u_ca_out_961));
compressor_81_24 u_ca_81_24_962(.d_in(u_ca_in_962), .d_out(u_ca_out_962));
compressor_81_24 u_ca_81_24_963(.d_in(u_ca_in_963), .d_out(u_ca_out_963));
compressor_81_24 u_ca_81_24_964(.d_in(u_ca_in_964), .d_out(u_ca_out_964));
compressor_81_24 u_ca_81_24_965(.d_in(u_ca_in_965), .d_out(u_ca_out_965));
compressor_81_24 u_ca_81_24_966(.d_in(u_ca_in_966), .d_out(u_ca_out_966));
compressor_81_24 u_ca_81_24_967(.d_in(u_ca_in_967), .d_out(u_ca_out_967));
compressor_81_24 u_ca_81_24_968(.d_in(u_ca_in_968), .d_out(u_ca_out_968));
compressor_81_24 u_ca_81_24_969(.d_in(u_ca_in_969), .d_out(u_ca_out_969));
compressor_81_24 u_ca_81_24_970(.d_in(u_ca_in_970), .d_out(u_ca_out_970));
compressor_81_24 u_ca_81_24_971(.d_in(u_ca_in_971), .d_out(u_ca_out_971));
compressor_81_24 u_ca_81_24_972(.d_in(u_ca_in_972), .d_out(u_ca_out_972));
compressor_81_24 u_ca_81_24_973(.d_in(u_ca_in_973), .d_out(u_ca_out_973));
compressor_81_24 u_ca_81_24_974(.d_in(u_ca_in_974), .d_out(u_ca_out_974));
compressor_81_24 u_ca_81_24_975(.d_in(u_ca_in_975), .d_out(u_ca_out_975));
compressor_81_24 u_ca_81_24_976(.d_in(u_ca_in_976), .d_out(u_ca_out_976));
compressor_81_24 u_ca_81_24_977(.d_in(u_ca_in_977), .d_out(u_ca_out_977));
compressor_81_24 u_ca_81_24_978(.d_in(u_ca_in_978), .d_out(u_ca_out_978));
compressor_81_24 u_ca_81_24_979(.d_in(u_ca_in_979), .d_out(u_ca_out_979));
compressor_81_24 u_ca_81_24_980(.d_in(u_ca_in_980), .d_out(u_ca_out_980));
compressor_81_24 u_ca_81_24_981(.d_in(u_ca_in_981), .d_out(u_ca_out_981));
compressor_81_24 u_ca_81_24_982(.d_in(u_ca_in_982), .d_out(u_ca_out_982));
compressor_81_24 u_ca_81_24_983(.d_in(u_ca_in_983), .d_out(u_ca_out_983));
compressor_81_24 u_ca_81_24_984(.d_in(u_ca_in_984), .d_out(u_ca_out_984));
compressor_81_24 u_ca_81_24_985(.d_in(u_ca_in_985), .d_out(u_ca_out_985));
compressor_81_24 u_ca_81_24_986(.d_in(u_ca_in_986), .d_out(u_ca_out_986));
compressor_81_24 u_ca_81_24_987(.d_in(u_ca_in_987), .d_out(u_ca_out_987));
compressor_81_24 u_ca_81_24_988(.d_in(u_ca_in_988), .d_out(u_ca_out_988));
compressor_81_24 u_ca_81_24_989(.d_in(u_ca_in_989), .d_out(u_ca_out_989));
compressor_81_24 u_ca_81_24_990(.d_in(u_ca_in_990), .d_out(u_ca_out_990));
compressor_81_24 u_ca_81_24_991(.d_in(u_ca_in_991), .d_out(u_ca_out_991));
compressor_81_24 u_ca_81_24_992(.d_in(u_ca_in_992), .d_out(u_ca_out_992));
compressor_81_24 u_ca_81_24_993(.d_in(u_ca_in_993), .d_out(u_ca_out_993));
compressor_81_24 u_ca_81_24_994(.d_in(u_ca_in_994), .d_out(u_ca_out_994));
compressor_81_24 u_ca_81_24_995(.d_in(u_ca_in_995), .d_out(u_ca_out_995));
compressor_81_24 u_ca_81_24_996(.d_in(u_ca_in_996), .d_out(u_ca_out_996));
compressor_81_24 u_ca_81_24_997(.d_in(u_ca_in_997), .d_out(u_ca_out_997));
compressor_81_24 u_ca_81_24_998(.d_in(u_ca_in_998), .d_out(u_ca_out_998));
compressor_81_24 u_ca_81_24_999(.d_in(u_ca_in_999), .d_out(u_ca_out_999));
compressor_81_24 u_ca_81_24_1000(.d_in(u_ca_in_1000), .d_out(u_ca_out_1000));
compressor_81_24 u_ca_81_24_1001(.d_in(u_ca_in_1001), .d_out(u_ca_out_1001));
compressor_81_24 u_ca_81_24_1002(.d_in(u_ca_in_1002), .d_out(u_ca_out_1002));
compressor_81_24 u_ca_81_24_1003(.d_in(u_ca_in_1003), .d_out(u_ca_out_1003));
compressor_81_24 u_ca_81_24_1004(.d_in(u_ca_in_1004), .d_out(u_ca_out_1004));
compressor_81_24 u_ca_81_24_1005(.d_in(u_ca_in_1005), .d_out(u_ca_out_1005));
compressor_81_24 u_ca_81_24_1006(.d_in(u_ca_in_1006), .d_out(u_ca_out_1006));
compressor_81_24 u_ca_81_24_1007(.d_in(u_ca_in_1007), .d_out(u_ca_out_1007));
compressor_81_24 u_ca_81_24_1008(.d_in(u_ca_in_1008), .d_out(u_ca_out_1008));
compressor_81_24 u_ca_81_24_1009(.d_in(u_ca_in_1009), .d_out(u_ca_out_1009));
compressor_81_24 u_ca_81_24_1010(.d_in(u_ca_in_1010), .d_out(u_ca_out_1010));
compressor_81_24 u_ca_81_24_1011(.d_in(u_ca_in_1011), .d_out(u_ca_out_1011));
compressor_81_24 u_ca_81_24_1012(.d_in(u_ca_in_1012), .d_out(u_ca_out_1012));
compressor_81_24 u_ca_81_24_1013(.d_in(u_ca_in_1013), .d_out(u_ca_out_1013));
compressor_81_24 u_ca_81_24_1014(.d_in(u_ca_in_1014), .d_out(u_ca_out_1014));
compressor_81_24 u_ca_81_24_1015(.d_in(u_ca_in_1015), .d_out(u_ca_out_1015));
compressor_81_24 u_ca_81_24_1016(.d_in(u_ca_in_1016), .d_out(u_ca_out_1016));
compressor_81_24 u_ca_81_24_1017(.d_in(u_ca_in_1017), .d_out(u_ca_out_1017));
compressor_81_24 u_ca_81_24_1018(.d_in(u_ca_in_1018), .d_out(u_ca_out_1018));
compressor_81_24 u_ca_81_24_1019(.d_in(u_ca_in_1019), .d_out(u_ca_out_1019));
compressor_81_24 u_ca_81_24_1020(.d_in(u_ca_in_1020), .d_out(u_ca_out_1020));
compressor_81_24 u_ca_81_24_1021(.d_in(u_ca_in_1021), .d_out(u_ca_out_1021));
compressor_81_24 u_ca_81_24_1022(.d_in(u_ca_in_1022), .d_out(u_ca_out_1022));
compressor_81_24 u_ca_81_24_1023(.d_in(u_ca_in_1023), .d_out(u_ca_out_1023));
compressor_81_24 u_ca_81_24_1024(.d_in(u_ca_in_1024), .d_out(u_ca_out_1024));
compressor_81_24 u_ca_81_24_1025(.d_in(u_ca_in_1025), .d_out(u_ca_out_1025));
compressor_81_24 u_ca_81_24_1026(.d_in(u_ca_in_1026), .d_out(u_ca_out_1026));
compressor_81_24 u_ca_81_24_1027(.d_in(u_ca_in_1027), .d_out(u_ca_out_1027));
compressor_81_24 u_ca_81_24_1028(.d_in(u_ca_in_1028), .d_out(u_ca_out_1028));
compressor_81_24 u_ca_81_24_1029(.d_in(u_ca_in_1029), .d_out(u_ca_out_1029));
compressor_81_24 u_ca_81_24_1030(.d_in(u_ca_in_1030), .d_out(u_ca_out_1030));
compressor_81_24 u_ca_81_24_1031(.d_in(u_ca_in_1031), .d_out(u_ca_out_1031));
compressor_81_24 u_ca_81_24_1032(.d_in(u_ca_in_1032), .d_out(u_ca_out_1032));
compressor_81_24 u_ca_81_24_1033(.d_in(u_ca_in_1033), .d_out(u_ca_out_1033));
compressor_81_24 u_ca_81_24_1034(.d_in(u_ca_in_1034), .d_out(u_ca_out_1034));
compressor_81_24 u_ca_81_24_1035(.d_in(u_ca_in_1035), .d_out(u_ca_out_1035));
compressor_81_24 u_ca_81_24_1036(.d_in(u_ca_in_1036), .d_out(u_ca_out_1036));
compressor_81_24 u_ca_81_24_1037(.d_in(u_ca_in_1037), .d_out(u_ca_out_1037));
compressor_81_24 u_ca_81_24_1038(.d_in(u_ca_in_1038), .d_out(u_ca_out_1038));
compressor_81_24 u_ca_81_24_1039(.d_in(u_ca_in_1039), .d_out(u_ca_out_1039));
compressor_81_24 u_ca_81_24_1040(.d_in(u_ca_in_1040), .d_out(u_ca_out_1040));
compressor_81_24 u_ca_81_24_1041(.d_in(u_ca_in_1041), .d_out(u_ca_out_1041));
compressor_81_24 u_ca_81_24_1042(.d_in(u_ca_in_1042), .d_out(u_ca_out_1042));
compressor_81_24 u_ca_81_24_1043(.d_in(u_ca_in_1043), .d_out(u_ca_out_1043));
compressor_81_24 u_ca_81_24_1044(.d_in(u_ca_in_1044), .d_out(u_ca_out_1044));
compressor_81_24 u_ca_81_24_1045(.d_in(u_ca_in_1045), .d_out(u_ca_out_1045));
compressor_81_24 u_ca_81_24_1046(.d_in(u_ca_in_1046), .d_out(u_ca_out_1046));
compressor_81_24 u_ca_81_24_1047(.d_in(u_ca_in_1047), .d_out(u_ca_out_1047));
compressor_81_24 u_ca_81_24_1048(.d_in(u_ca_in_1048), .d_out(u_ca_out_1048));
compressor_81_24 u_ca_81_24_1049(.d_in(u_ca_in_1049), .d_out(u_ca_out_1049));
compressor_81_24 u_ca_81_24_1050(.d_in(u_ca_in_1050), .d_out(u_ca_out_1050));
compressor_81_24 u_ca_81_24_1051(.d_in(u_ca_in_1051), .d_out(u_ca_out_1051));
compressor_81_24 u_ca_81_24_1052(.d_in(u_ca_in_1052), .d_out(u_ca_out_1052));
compressor_81_24 u_ca_81_24_1053(.d_in(u_ca_in_1053), .d_out(u_ca_out_1053));
compressor_81_24 u_ca_81_24_1054(.d_in(u_ca_in_1054), .d_out(u_ca_out_1054));
compressor_81_24 u_ca_81_24_1055(.d_in(u_ca_in_1055), .d_out(u_ca_out_1055));
compressor_81_24 u_ca_81_24_1056(.d_in(u_ca_in_1056), .d_out(u_ca_out_1056));
compressor_81_24 u_ca_81_24_1057(.d_in(u_ca_in_1057), .d_out(u_ca_out_1057));
compressor_81_24 u_ca_81_24_1058(.d_in(u_ca_in_1058), .d_out(u_ca_out_1058));
compressor_81_24 u_ca_81_24_1059(.d_in(u_ca_in_1059), .d_out(u_ca_out_1059));
compressor_81_24 u_ca_81_24_1060(.d_in(u_ca_in_1060), .d_out(u_ca_out_1060));
compressor_81_24 u_ca_81_24_1061(.d_in(u_ca_in_1061), .d_out(u_ca_out_1061));
compressor_81_24 u_ca_81_24_1062(.d_in(u_ca_in_1062), .d_out(u_ca_out_1062));
compressor_81_24 u_ca_81_24_1063(.d_in(u_ca_in_1063), .d_out(u_ca_out_1063));
compressor_81_24 u_ca_81_24_1064(.d_in(u_ca_in_1064), .d_out(u_ca_out_1064));
compressor_81_24 u_ca_81_24_1065(.d_in(u_ca_in_1065), .d_out(u_ca_out_1065));
compressor_81_24 u_ca_81_24_1066(.d_in(u_ca_in_1066), .d_out(u_ca_out_1066));
compressor_81_24 u_ca_81_24_1067(.d_in(u_ca_in_1067), .d_out(u_ca_out_1067));
compressor_81_24 u_ca_81_24_1068(.d_in(u_ca_in_1068), .d_out(u_ca_out_1068));
compressor_81_24 u_ca_81_24_1069(.d_in(u_ca_in_1069), .d_out(u_ca_out_1069));
compressor_81_24 u_ca_81_24_1070(.d_in(u_ca_in_1070), .d_out(u_ca_out_1070));
compressor_81_24 u_ca_81_24_1071(.d_in(u_ca_in_1071), .d_out(u_ca_out_1071));
compressor_81_24 u_ca_81_24_1072(.d_in(u_ca_in_1072), .d_out(u_ca_out_1072));
compressor_81_24 u_ca_81_24_1073(.d_in(u_ca_in_1073), .d_out(u_ca_out_1073));
compressor_81_24 u_ca_81_24_1074(.d_in(u_ca_in_1074), .d_out(u_ca_out_1074));
compressor_81_24 u_ca_81_24_1075(.d_in(u_ca_in_1075), .d_out(u_ca_out_1075));
compressor_81_24 u_ca_81_24_1076(.d_in(u_ca_in_1076), .d_out(u_ca_out_1076));
compressor_81_24 u_ca_81_24_1077(.d_in(u_ca_in_1077), .d_out(u_ca_out_1077));
compressor_81_24 u_ca_81_24_1078(.d_in(u_ca_in_1078), .d_out(u_ca_out_1078));
compressor_81_24 u_ca_81_24_1079(.d_in(u_ca_in_1079), .d_out(u_ca_out_1079));
compressor_81_24 u_ca_81_24_1080(.d_in(u_ca_in_1080), .d_out(u_ca_out_1080));
compressor_81_24 u_ca_81_24_1081(.d_in(u_ca_in_1081), .d_out(u_ca_out_1081));
compressor_81_24 u_ca_81_24_1082(.d_in(u_ca_in_1082), .d_out(u_ca_out_1082));
compressor_81_24 u_ca_81_24_1083(.d_in(u_ca_in_1083), .d_out(u_ca_out_1083));
compressor_81_24 u_ca_81_24_1084(.d_in(u_ca_in_1084), .d_out(u_ca_out_1084));
compressor_81_24 u_ca_81_24_1085(.d_in(u_ca_in_1085), .d_out(u_ca_out_1085));
compressor_81_24 u_ca_81_24_1086(.d_in(u_ca_in_1086), .d_out(u_ca_out_1086));
compressor_81_24 u_ca_81_24_1087(.d_in(u_ca_in_1087), .d_out(u_ca_out_1087));
compressor_81_24 u_ca_81_24_1088(.d_in(u_ca_in_1088), .d_out(u_ca_out_1088));
compressor_81_24 u_ca_81_24_1089(.d_in(u_ca_in_1089), .d_out(u_ca_out_1089));
compressor_81_24 u_ca_81_24_1090(.d_in(u_ca_in_1090), .d_out(u_ca_out_1090));
compressor_81_24 u_ca_81_24_1091(.d_in(u_ca_in_1091), .d_out(u_ca_out_1091));
compressor_81_24 u_ca_81_24_1092(.d_in(u_ca_in_1092), .d_out(u_ca_out_1092));
compressor_81_24 u_ca_81_24_1093(.d_in(u_ca_in_1093), .d_out(u_ca_out_1093));
compressor_81_24 u_ca_81_24_1094(.d_in(u_ca_in_1094), .d_out(u_ca_out_1094));
compressor_81_24 u_ca_81_24_1095(.d_in(u_ca_in_1095), .d_out(u_ca_out_1095));
compressor_81_24 u_ca_81_24_1096(.d_in(u_ca_in_1096), .d_out(u_ca_out_1096));
compressor_81_24 u_ca_81_24_1097(.d_in(u_ca_in_1097), .d_out(u_ca_out_1097));
compressor_81_24 u_ca_81_24_1098(.d_in(u_ca_in_1098), .d_out(u_ca_out_1098));
compressor_81_24 u_ca_81_24_1099(.d_in(u_ca_in_1099), .d_out(u_ca_out_1099));
compressor_81_24 u_ca_81_24_1100(.d_in(u_ca_in_1100), .d_out(u_ca_out_1100));
compressor_81_24 u_ca_81_24_1101(.d_in(u_ca_in_1101), .d_out(u_ca_out_1101));
compressor_81_24 u_ca_81_24_1102(.d_in(u_ca_in_1102), .d_out(u_ca_out_1102));
compressor_81_24 u_ca_81_24_1103(.d_in(u_ca_in_1103), .d_out(u_ca_out_1103));
compressor_81_24 u_ca_81_24_1104(.d_in(u_ca_in_1104), .d_out(u_ca_out_1104));
compressor_81_24 u_ca_81_24_1105(.d_in(u_ca_in_1105), .d_out(u_ca_out_1105));
compressor_81_24 u_ca_81_24_1106(.d_in(u_ca_in_1106), .d_out(u_ca_out_1106));
compressor_81_24 u_ca_81_24_1107(.d_in(u_ca_in_1107), .d_out(u_ca_out_1107));
compressor_81_24 u_ca_81_24_1108(.d_in(u_ca_in_1108), .d_out(u_ca_out_1108));
compressor_81_24 u_ca_81_24_1109(.d_in(u_ca_in_1109), .d_out(u_ca_out_1109));
compressor_81_24 u_ca_81_24_1110(.d_in(u_ca_in_1110), .d_out(u_ca_out_1110));
compressor_81_24 u_ca_81_24_1111(.d_in(u_ca_in_1111), .d_out(u_ca_out_1111));
compressor_81_24 u_ca_81_24_1112(.d_in(u_ca_in_1112), .d_out(u_ca_out_1112));
compressor_81_24 u_ca_81_24_1113(.d_in(u_ca_in_1113), .d_out(u_ca_out_1113));
compressor_81_24 u_ca_81_24_1114(.d_in(u_ca_in_1114), .d_out(u_ca_out_1114));
compressor_81_24 u_ca_81_24_1115(.d_in(u_ca_in_1115), .d_out(u_ca_out_1115));
compressor_81_24 u_ca_81_24_1116(.d_in(u_ca_in_1116), .d_out(u_ca_out_1116));
compressor_81_24 u_ca_81_24_1117(.d_in(u_ca_in_1117), .d_out(u_ca_out_1117));
compressor_81_24 u_ca_81_24_1118(.d_in(u_ca_in_1118), .d_out(u_ca_out_1118));
compressor_81_24 u_ca_81_24_1119(.d_in(u_ca_in_1119), .d_out(u_ca_out_1119));
compressor_81_24 u_ca_81_24_1120(.d_in(u_ca_in_1120), .d_out(u_ca_out_1120));
compressor_81_24 u_ca_81_24_1121(.d_in(u_ca_in_1121), .d_out(u_ca_out_1121));
compressor_81_24 u_ca_81_24_1122(.d_in(u_ca_in_1122), .d_out(u_ca_out_1122));
compressor_81_24 u_ca_81_24_1123(.d_in(u_ca_in_1123), .d_out(u_ca_out_1123));
compressor_81_24 u_ca_81_24_1124(.d_in(u_ca_in_1124), .d_out(u_ca_out_1124));
compressor_81_24 u_ca_81_24_1125(.d_in(u_ca_in_1125), .d_out(u_ca_out_1125));
compressor_81_24 u_ca_81_24_1126(.d_in(u_ca_in_1126), .d_out(u_ca_out_1126));
compressor_81_24 u_ca_81_24_1127(.d_in(u_ca_in_1127), .d_out(u_ca_out_1127));
compressor_81_24 u_ca_81_24_1128(.d_in(u_ca_in_1128), .d_out(u_ca_out_1128));
compressor_81_24 u_ca_81_24_1129(.d_in(u_ca_in_1129), .d_out(u_ca_out_1129));
compressor_81_24 u_ca_81_24_1130(.d_in(u_ca_in_1130), .d_out(u_ca_out_1130));
compressor_81_24 u_ca_81_24_1131(.d_in(u_ca_in_1131), .d_out(u_ca_out_1131));
compressor_81_24 u_ca_81_24_1132(.d_in(u_ca_in_1132), .d_out(u_ca_out_1132));
compressor_81_24 u_ca_81_24_1133(.d_in(u_ca_in_1133), .d_out(u_ca_out_1133));
compressor_81_24 u_ca_81_24_1134(.d_in(u_ca_in_1134), .d_out(u_ca_out_1134));
compressor_81_24 u_ca_81_24_1135(.d_in(u_ca_in_1135), .d_out(u_ca_out_1135));
compressor_81_24 u_ca_81_24_1136(.d_in(u_ca_in_1136), .d_out(u_ca_out_1136));
compressor_81_24 u_ca_81_24_1137(.d_in(u_ca_in_1137), .d_out(u_ca_out_1137));
compressor_81_24 u_ca_81_24_1138(.d_in(u_ca_in_1138), .d_out(u_ca_out_1138));
compressor_81_24 u_ca_81_24_1139(.d_in(u_ca_in_1139), .d_out(u_ca_out_1139));
compressor_81_24 u_ca_81_24_1140(.d_in(u_ca_in_1140), .d_out(u_ca_out_1140));
compressor_81_24 u_ca_81_24_1141(.d_in(u_ca_in_1141), .d_out(u_ca_out_1141));
compressor_81_24 u_ca_81_24_1142(.d_in(u_ca_in_1142), .d_out(u_ca_out_1142));
compressor_81_24 u_ca_81_24_1143(.d_in(u_ca_in_1143), .d_out(u_ca_out_1143));
compressor_81_24 u_ca_81_24_1144(.d_in(u_ca_in_1144), .d_out(u_ca_out_1144));
compressor_81_24 u_ca_81_24_1145(.d_in(u_ca_in_1145), .d_out(u_ca_out_1145));
compressor_81_24 u_ca_81_24_1146(.d_in(u_ca_in_1146), .d_out(u_ca_out_1146));
compressor_81_24 u_ca_81_24_1147(.d_in(u_ca_in_1147), .d_out(u_ca_out_1147));
compressor_81_24 u_ca_81_24_1148(.d_in(u_ca_in_1148), .d_out(u_ca_out_1148));
compressor_81_24 u_ca_81_24_1149(.d_in(u_ca_in_1149), .d_out(u_ca_out_1149));
compressor_81_24 u_ca_81_24_1150(.d_in(u_ca_in_1150), .d_out(u_ca_out_1150));
compressor_81_24 u_ca_81_24_1151(.d_in(u_ca_in_1151), .d_out(u_ca_out_1151));
compressor_81_24 u_ca_81_24_1152(.d_in(u_ca_in_1152), .d_out(u_ca_out_1152));
compressor_81_24 u_ca_81_24_1153(.d_in(u_ca_in_1153), .d_out(u_ca_out_1153));
compressor_81_24 u_ca_81_24_1154(.d_in(u_ca_in_1154), .d_out(u_ca_out_1154));
compressor_81_24 u_ca_81_24_1155(.d_in(u_ca_in_1155), .d_out(u_ca_out_1155));
compressor_81_24 u_ca_81_24_1156(.d_in(u_ca_in_1156), .d_out(u_ca_out_1156));
compressor_81_24 u_ca_81_24_1157(.d_in(u_ca_in_1157), .d_out(u_ca_out_1157));
compressor_81_24 u_ca_81_24_1158(.d_in(u_ca_in_1158), .d_out(u_ca_out_1158));
compressor_81_24 u_ca_81_24_1159(.d_in(u_ca_in_1159), .d_out(u_ca_out_1159));
compressor_81_24 u_ca_81_24_1160(.d_in(u_ca_in_1160), .d_out(u_ca_out_1160));
compressor_81_24 u_ca_81_24_1161(.d_in(u_ca_in_1161), .d_out(u_ca_out_1161));
compressor_81_24 u_ca_81_24_1162(.d_in(u_ca_in_1162), .d_out(u_ca_out_1162));
compressor_81_24 u_ca_81_24_1163(.d_in(u_ca_in_1163), .d_out(u_ca_out_1163));
compressor_81_24 u_ca_81_24_1164(.d_in(u_ca_in_1164), .d_out(u_ca_out_1164));
compressor_81_24 u_ca_81_24_1165(.d_in(u_ca_in_1165), .d_out(u_ca_out_1165));
compressor_81_24 u_ca_81_24_1166(.d_in(u_ca_in_1166), .d_out(u_ca_out_1166));
compressor_81_24 u_ca_81_24_1167(.d_in(u_ca_in_1167), .d_out(u_ca_out_1167));
compressor_81_24 u_ca_81_24_1168(.d_in(u_ca_in_1168), .d_out(u_ca_out_1168));
compressor_81_24 u_ca_81_24_1169(.d_in(u_ca_in_1169), .d_out(u_ca_out_1169));
compressor_81_24 u_ca_81_24_1170(.d_in(u_ca_in_1170), .d_out(u_ca_out_1170));
compressor_81_24 u_ca_81_24_1171(.d_in(u_ca_in_1171), .d_out(u_ca_out_1171));
compressor_81_24 u_ca_81_24_1172(.d_in(u_ca_in_1172), .d_out(u_ca_out_1172));
compressor_81_24 u_ca_81_24_1173(.d_in(u_ca_in_1173), .d_out(u_ca_out_1173));
compressor_81_24 u_ca_81_24_1174(.d_in(u_ca_in_1174), .d_out(u_ca_out_1174));
compressor_81_24 u_ca_81_24_1175(.d_in(u_ca_in_1175), .d_out(u_ca_out_1175));
compressor_81_24 u_ca_81_24_1176(.d_in(u_ca_in_1176), .d_out(u_ca_out_1176));
compressor_81_24 u_ca_81_24_1177(.d_in(u_ca_in_1177), .d_out(u_ca_out_1177));
compressor_81_24 u_ca_81_24_1178(.d_in(u_ca_in_1178), .d_out(u_ca_out_1178));
compressor_81_24 u_ca_81_24_1179(.d_in(u_ca_in_1179), .d_out(u_ca_out_1179));
compressor_81_24 u_ca_81_24_1180(.d_in(u_ca_in_1180), .d_out(u_ca_out_1180));
compressor_81_24 u_ca_81_24_1181(.d_in(u_ca_in_1181), .d_out(u_ca_out_1181));
compressor_81_24 u_ca_81_24_1182(.d_in(u_ca_in_1182), .d_out(u_ca_out_1182));
compressor_81_24 u_ca_81_24_1183(.d_in(u_ca_in_1183), .d_out(u_ca_out_1183));
compressor_81_24 u_ca_81_24_1184(.d_in(u_ca_in_1184), .d_out(u_ca_out_1184));
compressor_81_24 u_ca_81_24_1185(.d_in(u_ca_in_1185), .d_out(u_ca_out_1185));
compressor_81_24 u_ca_81_24_1186(.d_in(u_ca_in_1186), .d_out(u_ca_out_1186));
compressor_81_24 u_ca_81_24_1187(.d_in(u_ca_in_1187), .d_out(u_ca_out_1187));
compressor_81_24 u_ca_81_24_1188(.d_in(u_ca_in_1188), .d_out(u_ca_out_1188));
compressor_81_24 u_ca_81_24_1189(.d_in(u_ca_in_1189), .d_out(u_ca_out_1189));
compressor_81_24 u_ca_81_24_1190(.d_in(u_ca_in_1190), .d_out(u_ca_out_1190));
compressor_81_24 u_ca_81_24_1191(.d_in(u_ca_in_1191), .d_out(u_ca_out_1191));
compressor_81_24 u_ca_81_24_1192(.d_in(u_ca_in_1192), .d_out(u_ca_out_1192));
compressor_81_24 u_ca_81_24_1193(.d_in(u_ca_in_1193), .d_out(u_ca_out_1193));
compressor_81_24 u_ca_81_24_1194(.d_in(u_ca_in_1194), .d_out(u_ca_out_1194));
compressor_81_24 u_ca_81_24_1195(.d_in(u_ca_in_1195), .d_out(u_ca_out_1195));
compressor_81_24 u_ca_81_24_1196(.d_in(u_ca_in_1196), .d_out(u_ca_out_1196));
compressor_81_24 u_ca_81_24_1197(.d_in(u_ca_in_1197), .d_out(u_ca_out_1197));
compressor_81_24 u_ca_81_24_1198(.d_in(u_ca_in_1198), .d_out(u_ca_out_1198));
compressor_81_24 u_ca_81_24_1199(.d_in(u_ca_in_1199), .d_out(u_ca_out_1199));
compressor_81_24 u_ca_81_24_1200(.d_in(u_ca_in_1200), .d_out(u_ca_out_1200));
compressor_81_24 u_ca_81_24_1201(.d_in(u_ca_in_1201), .d_out(u_ca_out_1201));
compressor_81_24 u_ca_81_24_1202(.d_in(u_ca_in_1202), .d_out(u_ca_out_1202));
compressor_81_24 u_ca_81_24_1203(.d_in(u_ca_in_1203), .d_out(u_ca_out_1203));
compressor_81_24 u_ca_81_24_1204(.d_in(u_ca_in_1204), .d_out(u_ca_out_1204));
compressor_81_24 u_ca_81_24_1205(.d_in(u_ca_in_1205), .d_out(u_ca_out_1205));
compressor_81_24 u_ca_81_24_1206(.d_in(u_ca_in_1206), .d_out(u_ca_out_1206));
compressor_81_24 u_ca_81_24_1207(.d_in(u_ca_in_1207), .d_out(u_ca_out_1207));
compressor_81_24 u_ca_81_24_1208(.d_in(u_ca_in_1208), .d_out(u_ca_out_1208));
compressor_81_24 u_ca_81_24_1209(.d_in(u_ca_in_1209), .d_out(u_ca_out_1209));
compressor_81_24 u_ca_81_24_1210(.d_in(u_ca_in_1210), .d_out(u_ca_out_1210));
compressor_81_24 u_ca_81_24_1211(.d_in(u_ca_in_1211), .d_out(u_ca_out_1211));
compressor_81_24 u_ca_81_24_1212(.d_in(u_ca_in_1212), .d_out(u_ca_out_1212));
compressor_81_24 u_ca_81_24_1213(.d_in(u_ca_in_1213), .d_out(u_ca_out_1213));
compressor_81_24 u_ca_81_24_1214(.d_in(u_ca_in_1214), .d_out(u_ca_out_1214));
compressor_81_24 u_ca_81_24_1215(.d_in(u_ca_in_1215), .d_out(u_ca_out_1215));
compressor_81_24 u_ca_81_24_1216(.d_in(u_ca_in_1216), .d_out(u_ca_out_1216));
compressor_81_24 u_ca_81_24_1217(.d_in(u_ca_in_1217), .d_out(u_ca_out_1217));
compressor_81_24 u_ca_81_24_1218(.d_in(u_ca_in_1218), .d_out(u_ca_out_1218));
compressor_81_24 u_ca_81_24_1219(.d_in(u_ca_in_1219), .d_out(u_ca_out_1219));
compressor_81_24 u_ca_81_24_1220(.d_in(u_ca_in_1220), .d_out(u_ca_out_1220));
compressor_81_24 u_ca_81_24_1221(.d_in(u_ca_in_1221), .d_out(u_ca_out_1221));
compressor_81_24 u_ca_81_24_1222(.d_in(u_ca_in_1222), .d_out(u_ca_out_1222));
compressor_81_24 u_ca_81_24_1223(.d_in(u_ca_in_1223), .d_out(u_ca_out_1223));
compressor_81_24 u_ca_81_24_1224(.d_in(u_ca_in_1224), .d_out(u_ca_out_1224));
compressor_81_24 u_ca_81_24_1225(.d_in(u_ca_in_1225), .d_out(u_ca_out_1225));
compressor_81_24 u_ca_81_24_1226(.d_in(u_ca_in_1226), .d_out(u_ca_out_1226));
compressor_81_24 u_ca_81_24_1227(.d_in(u_ca_in_1227), .d_out(u_ca_out_1227));
compressor_81_24 u_ca_81_24_1228(.d_in(u_ca_in_1228), .d_out(u_ca_out_1228));
compressor_81_24 u_ca_81_24_1229(.d_in(u_ca_in_1229), .d_out(u_ca_out_1229));
compressor_81_24 u_ca_81_24_1230(.d_in(u_ca_in_1230), .d_out(u_ca_out_1230));
compressor_81_24 u_ca_81_24_1231(.d_in(u_ca_in_1231), .d_out(u_ca_out_1231));
compressor_81_24 u_ca_81_24_1232(.d_in(u_ca_in_1232), .d_out(u_ca_out_1232));
compressor_81_24 u_ca_81_24_1233(.d_in(u_ca_in_1233), .d_out(u_ca_out_1233));
compressor_81_24 u_ca_81_24_1234(.d_in(u_ca_in_1234), .d_out(u_ca_out_1234));
compressor_81_24 u_ca_81_24_1235(.d_in(u_ca_in_1235), .d_out(u_ca_out_1235));
compressor_81_24 u_ca_81_24_1236(.d_in(u_ca_in_1236), .d_out(u_ca_out_1236));
compressor_81_24 u_ca_81_24_1237(.d_in(u_ca_in_1237), .d_out(u_ca_out_1237));
compressor_81_24 u_ca_81_24_1238(.d_in(u_ca_in_1238), .d_out(u_ca_out_1238));
compressor_81_24 u_ca_81_24_1239(.d_in(u_ca_in_1239), .d_out(u_ca_out_1239));
compressor_81_24 u_ca_81_24_1240(.d_in(u_ca_in_1240), .d_out(u_ca_out_1240));
compressor_81_24 u_ca_81_24_1241(.d_in(u_ca_in_1241), .d_out(u_ca_out_1241));
compressor_81_24 u_ca_81_24_1242(.d_in(u_ca_in_1242), .d_out(u_ca_out_1242));
compressor_81_24 u_ca_81_24_1243(.d_in(u_ca_in_1243), .d_out(u_ca_out_1243));
compressor_81_24 u_ca_81_24_1244(.d_in(u_ca_in_1244), .d_out(u_ca_out_1244));
compressor_81_24 u_ca_81_24_1245(.d_in(u_ca_in_1245), .d_out(u_ca_out_1245));
compressor_81_24 u_ca_81_24_1246(.d_in(u_ca_in_1246), .d_out(u_ca_out_1246));
compressor_81_24 u_ca_81_24_1247(.d_in(u_ca_in_1247), .d_out(u_ca_out_1247));
compressor_81_24 u_ca_81_24_1248(.d_in(u_ca_in_1248), .d_out(u_ca_out_1248));
compressor_81_24 u_ca_81_24_1249(.d_in(u_ca_in_1249), .d_out(u_ca_out_1249));
compressor_81_24 u_ca_81_24_1250(.d_in(u_ca_in_1250), .d_out(u_ca_out_1250));
compressor_81_24 u_ca_81_24_1251(.d_in(u_ca_in_1251), .d_out(u_ca_out_1251));
compressor_81_24 u_ca_81_24_1252(.d_in(u_ca_in_1252), .d_out(u_ca_out_1252));
compressor_81_24 u_ca_81_24_1253(.d_in(u_ca_in_1253), .d_out(u_ca_out_1253));
compressor_81_24 u_ca_81_24_1254(.d_in(u_ca_in_1254), .d_out(u_ca_out_1254));
compressor_81_24 u_ca_81_24_1255(.d_in(u_ca_in_1255), .d_out(u_ca_out_1255));
compressor_81_24 u_ca_81_24_1256(.d_in(u_ca_in_1256), .d_out(u_ca_out_1256));
compressor_81_24 u_ca_81_24_1257(.d_in(u_ca_in_1257), .d_out(u_ca_out_1257));
compressor_81_24 u_ca_81_24_1258(.d_in(u_ca_in_1258), .d_out(u_ca_out_1258));
compressor_81_24 u_ca_81_24_1259(.d_in(u_ca_in_1259), .d_out(u_ca_out_1259));
compressor_81_24 u_ca_81_24_1260(.d_in(u_ca_in_1260), .d_out(u_ca_out_1260));
compressor_81_24 u_ca_81_24_1261(.d_in(u_ca_in_1261), .d_out(u_ca_out_1261));
compressor_81_24 u_ca_81_24_1262(.d_in(u_ca_in_1262), .d_out(u_ca_out_1262));
compressor_81_24 u_ca_81_24_1263(.d_in(u_ca_in_1263), .d_out(u_ca_out_1263));
compressor_81_24 u_ca_81_24_1264(.d_in(u_ca_in_1264), .d_out(u_ca_out_1264));
compressor_81_24 u_ca_81_24_1265(.d_in(u_ca_in_1265), .d_out(u_ca_out_1265));
compressor_81_24 u_ca_81_24_1266(.d_in(u_ca_in_1266), .d_out(u_ca_out_1266));
compressor_81_24 u_ca_81_24_1267(.d_in(u_ca_in_1267), .d_out(u_ca_out_1267));
compressor_81_24 u_ca_81_24_1268(.d_in(u_ca_in_1268), .d_out(u_ca_out_1268));
compressor_81_24 u_ca_81_24_1269(.d_in(u_ca_in_1269), .d_out(u_ca_out_1269));
compressor_81_24 u_ca_81_24_1270(.d_in(u_ca_in_1270), .d_out(u_ca_out_1270));
compressor_81_24 u_ca_81_24_1271(.d_in(u_ca_in_1271), .d_out(u_ca_out_1271));
compressor_81_24 u_ca_81_24_1272(.d_in(u_ca_in_1272), .d_out(u_ca_out_1272));
compressor_81_24 u_ca_81_24_1273(.d_in(u_ca_in_1273), .d_out(u_ca_out_1273));
compressor_81_24 u_ca_81_24_1274(.d_in(u_ca_in_1274), .d_out(u_ca_out_1274));
compressor_81_24 u_ca_81_24_1275(.d_in(u_ca_in_1275), .d_out(u_ca_out_1275));
compressor_81_24 u_ca_81_24_1276(.d_in(u_ca_in_1276), .d_out(u_ca_out_1276));
compressor_81_24 u_ca_81_24_1277(.d_in(u_ca_in_1277), .d_out(u_ca_out_1277));
compressor_81_24 u_ca_81_24_1278(.d_in(u_ca_in_1278), .d_out(u_ca_out_1278));
compressor_81_24 u_ca_81_24_1279(.d_in(u_ca_in_1279), .d_out(u_ca_out_1279));
compressor_81_24 u_ca_81_24_1280(.d_in(u_ca_in_1280), .d_out(u_ca_out_1280));
compressor_81_24 u_ca_81_24_1281(.d_in(u_ca_in_1281), .d_out(u_ca_out_1281));
compressor_81_24 u_ca_81_24_1282(.d_in(u_ca_in_1282), .d_out(u_ca_out_1282));

//---------------------------------------------------------



//--output-------------------------------------------------

assign col_out_0 = {{21{1'b0}}, u_ca_out_0[2:0]};
assign col_out_1 = {{12{1'b0}}, u_ca_out_1[2:0], u_ca_out_0[11:3]};
assign col_out_2 = {{3{1'b0}}, u_ca_out_2[2:0], u_ca_out_1[11:3], u_ca_out_0[20:12]};
assign col_out_3 = {u_ca_out_3[2:0],u_ca_out_2[11:3], u_ca_out_1[20:12], u_ca_out_0[23:21]};
assign col_out_4 = {u_ca_out_4[2:0],u_ca_out_3[11:3], u_ca_out_2[20:12], u_ca_out_1[23:21]};
assign col_out_5 = {u_ca_out_5[2:0],u_ca_out_4[11:3], u_ca_out_3[20:12], u_ca_out_2[23:21]};
assign col_out_6 = {u_ca_out_6[2:0],u_ca_out_5[11:3], u_ca_out_4[20:12], u_ca_out_3[23:21]};
assign col_out_7 = {u_ca_out_7[2:0],u_ca_out_6[11:3], u_ca_out_5[20:12], u_ca_out_4[23:21]};
assign col_out_8 = {u_ca_out_8[2:0],u_ca_out_7[11:3], u_ca_out_6[20:12], u_ca_out_5[23:21]};
assign col_out_9 = {u_ca_out_9[2:0],u_ca_out_8[11:3], u_ca_out_7[20:12], u_ca_out_6[23:21]};
assign col_out_10 = {u_ca_out_10[2:0],u_ca_out_9[11:3], u_ca_out_8[20:12], u_ca_out_7[23:21]};
assign col_out_11 = {u_ca_out_11[2:0],u_ca_out_10[11:3], u_ca_out_9[20:12], u_ca_out_8[23:21]};
assign col_out_12 = {u_ca_out_12[2:0],u_ca_out_11[11:3], u_ca_out_10[20:12], u_ca_out_9[23:21]};
assign col_out_13 = {u_ca_out_13[2:0],u_ca_out_12[11:3], u_ca_out_11[20:12], u_ca_out_10[23:21]};
assign col_out_14 = {u_ca_out_14[2:0],u_ca_out_13[11:3], u_ca_out_12[20:12], u_ca_out_11[23:21]};
assign col_out_15 = {u_ca_out_15[2:0],u_ca_out_14[11:3], u_ca_out_13[20:12], u_ca_out_12[23:21]};
assign col_out_16 = {u_ca_out_16[2:0],u_ca_out_15[11:3], u_ca_out_14[20:12], u_ca_out_13[23:21]};
assign col_out_17 = {u_ca_out_17[2:0],u_ca_out_16[11:3], u_ca_out_15[20:12], u_ca_out_14[23:21]};
assign col_out_18 = {u_ca_out_18[2:0],u_ca_out_17[11:3], u_ca_out_16[20:12], u_ca_out_15[23:21]};
assign col_out_19 = {u_ca_out_19[2:0],u_ca_out_18[11:3], u_ca_out_17[20:12], u_ca_out_16[23:21]};
assign col_out_20 = {u_ca_out_20[2:0],u_ca_out_19[11:3], u_ca_out_18[20:12], u_ca_out_17[23:21]};
assign col_out_21 = {u_ca_out_21[2:0],u_ca_out_20[11:3], u_ca_out_19[20:12], u_ca_out_18[23:21]};
assign col_out_22 = {u_ca_out_22[2:0],u_ca_out_21[11:3], u_ca_out_20[20:12], u_ca_out_19[23:21]};
assign col_out_23 = {u_ca_out_23[2:0],u_ca_out_22[11:3], u_ca_out_21[20:12], u_ca_out_20[23:21]};
assign col_out_24 = {u_ca_out_24[2:0],u_ca_out_23[11:3], u_ca_out_22[20:12], u_ca_out_21[23:21]};
assign col_out_25 = {u_ca_out_25[2:0],u_ca_out_24[11:3], u_ca_out_23[20:12], u_ca_out_22[23:21]};
assign col_out_26 = {u_ca_out_26[2:0],u_ca_out_25[11:3], u_ca_out_24[20:12], u_ca_out_23[23:21]};
assign col_out_27 = {u_ca_out_27[2:0],u_ca_out_26[11:3], u_ca_out_25[20:12], u_ca_out_24[23:21]};
assign col_out_28 = {u_ca_out_28[2:0],u_ca_out_27[11:3], u_ca_out_26[20:12], u_ca_out_25[23:21]};
assign col_out_29 = {u_ca_out_29[2:0],u_ca_out_28[11:3], u_ca_out_27[20:12], u_ca_out_26[23:21]};
assign col_out_30 = {u_ca_out_30[2:0],u_ca_out_29[11:3], u_ca_out_28[20:12], u_ca_out_27[23:21]};
assign col_out_31 = {u_ca_out_31[2:0],u_ca_out_30[11:3], u_ca_out_29[20:12], u_ca_out_28[23:21]};
assign col_out_32 = {u_ca_out_32[2:0],u_ca_out_31[11:3], u_ca_out_30[20:12], u_ca_out_29[23:21]};
assign col_out_33 = {u_ca_out_33[2:0],u_ca_out_32[11:3], u_ca_out_31[20:12], u_ca_out_30[23:21]};
assign col_out_34 = {u_ca_out_34[2:0],u_ca_out_33[11:3], u_ca_out_32[20:12], u_ca_out_31[23:21]};
assign col_out_35 = {u_ca_out_35[2:0],u_ca_out_34[11:3], u_ca_out_33[20:12], u_ca_out_32[23:21]};
assign col_out_36 = {u_ca_out_36[2:0],u_ca_out_35[11:3], u_ca_out_34[20:12], u_ca_out_33[23:21]};
assign col_out_37 = {u_ca_out_37[2:0],u_ca_out_36[11:3], u_ca_out_35[20:12], u_ca_out_34[23:21]};
assign col_out_38 = {u_ca_out_38[2:0],u_ca_out_37[11:3], u_ca_out_36[20:12], u_ca_out_35[23:21]};
assign col_out_39 = {u_ca_out_39[2:0],u_ca_out_38[11:3], u_ca_out_37[20:12], u_ca_out_36[23:21]};
assign col_out_40 = {u_ca_out_40[2:0],u_ca_out_39[11:3], u_ca_out_38[20:12], u_ca_out_37[23:21]};
assign col_out_41 = {u_ca_out_41[2:0],u_ca_out_40[11:3], u_ca_out_39[20:12], u_ca_out_38[23:21]};
assign col_out_42 = {u_ca_out_42[2:0],u_ca_out_41[11:3], u_ca_out_40[20:12], u_ca_out_39[23:21]};
assign col_out_43 = {u_ca_out_43[2:0],u_ca_out_42[11:3], u_ca_out_41[20:12], u_ca_out_40[23:21]};
assign col_out_44 = {u_ca_out_44[2:0],u_ca_out_43[11:3], u_ca_out_42[20:12], u_ca_out_41[23:21]};
assign col_out_45 = {u_ca_out_45[2:0],u_ca_out_44[11:3], u_ca_out_43[20:12], u_ca_out_42[23:21]};
assign col_out_46 = {u_ca_out_46[2:0],u_ca_out_45[11:3], u_ca_out_44[20:12], u_ca_out_43[23:21]};
assign col_out_47 = {u_ca_out_47[2:0],u_ca_out_46[11:3], u_ca_out_45[20:12], u_ca_out_44[23:21]};
assign col_out_48 = {u_ca_out_48[2:0],u_ca_out_47[11:3], u_ca_out_46[20:12], u_ca_out_45[23:21]};
assign col_out_49 = {u_ca_out_49[2:0],u_ca_out_48[11:3], u_ca_out_47[20:12], u_ca_out_46[23:21]};
assign col_out_50 = {u_ca_out_50[2:0],u_ca_out_49[11:3], u_ca_out_48[20:12], u_ca_out_47[23:21]};
assign col_out_51 = {u_ca_out_51[2:0],u_ca_out_50[11:3], u_ca_out_49[20:12], u_ca_out_48[23:21]};
assign col_out_52 = {u_ca_out_52[2:0],u_ca_out_51[11:3], u_ca_out_50[20:12], u_ca_out_49[23:21]};
assign col_out_53 = {u_ca_out_53[2:0],u_ca_out_52[11:3], u_ca_out_51[20:12], u_ca_out_50[23:21]};
assign col_out_54 = {u_ca_out_54[2:0],u_ca_out_53[11:3], u_ca_out_52[20:12], u_ca_out_51[23:21]};
assign col_out_55 = {u_ca_out_55[2:0],u_ca_out_54[11:3], u_ca_out_53[20:12], u_ca_out_52[23:21]};
assign col_out_56 = {u_ca_out_56[2:0],u_ca_out_55[11:3], u_ca_out_54[20:12], u_ca_out_53[23:21]};
assign col_out_57 = {u_ca_out_57[2:0],u_ca_out_56[11:3], u_ca_out_55[20:12], u_ca_out_54[23:21]};
assign col_out_58 = {u_ca_out_58[2:0],u_ca_out_57[11:3], u_ca_out_56[20:12], u_ca_out_55[23:21]};
assign col_out_59 = {u_ca_out_59[2:0],u_ca_out_58[11:3], u_ca_out_57[20:12], u_ca_out_56[23:21]};
assign col_out_60 = {u_ca_out_60[2:0],u_ca_out_59[11:3], u_ca_out_58[20:12], u_ca_out_57[23:21]};
assign col_out_61 = {u_ca_out_61[2:0],u_ca_out_60[11:3], u_ca_out_59[20:12], u_ca_out_58[23:21]};
assign col_out_62 = {u_ca_out_62[2:0],u_ca_out_61[11:3], u_ca_out_60[20:12], u_ca_out_59[23:21]};
assign col_out_63 = {u_ca_out_63[2:0],u_ca_out_62[11:3], u_ca_out_61[20:12], u_ca_out_60[23:21]};
assign col_out_64 = {u_ca_out_64[2:0],u_ca_out_63[11:3], u_ca_out_62[20:12], u_ca_out_61[23:21]};
assign col_out_65 = {u_ca_out_65[2:0],u_ca_out_64[11:3], u_ca_out_63[20:12], u_ca_out_62[23:21]};
assign col_out_66 = {u_ca_out_66[2:0],u_ca_out_65[11:3], u_ca_out_64[20:12], u_ca_out_63[23:21]};
assign col_out_67 = {u_ca_out_67[2:0],u_ca_out_66[11:3], u_ca_out_65[20:12], u_ca_out_64[23:21]};
assign col_out_68 = {u_ca_out_68[2:0],u_ca_out_67[11:3], u_ca_out_66[20:12], u_ca_out_65[23:21]};
assign col_out_69 = {u_ca_out_69[2:0],u_ca_out_68[11:3], u_ca_out_67[20:12], u_ca_out_66[23:21]};
assign col_out_70 = {u_ca_out_70[2:0],u_ca_out_69[11:3], u_ca_out_68[20:12], u_ca_out_67[23:21]};
assign col_out_71 = {u_ca_out_71[2:0],u_ca_out_70[11:3], u_ca_out_69[20:12], u_ca_out_68[23:21]};
assign col_out_72 = {u_ca_out_72[2:0],u_ca_out_71[11:3], u_ca_out_70[20:12], u_ca_out_69[23:21]};
assign col_out_73 = {u_ca_out_73[2:0],u_ca_out_72[11:3], u_ca_out_71[20:12], u_ca_out_70[23:21]};
assign col_out_74 = {u_ca_out_74[2:0],u_ca_out_73[11:3], u_ca_out_72[20:12], u_ca_out_71[23:21]};
assign col_out_75 = {u_ca_out_75[2:0],u_ca_out_74[11:3], u_ca_out_73[20:12], u_ca_out_72[23:21]};
assign col_out_76 = {u_ca_out_76[2:0],u_ca_out_75[11:3], u_ca_out_74[20:12], u_ca_out_73[23:21]};
assign col_out_77 = {u_ca_out_77[2:0],u_ca_out_76[11:3], u_ca_out_75[20:12], u_ca_out_74[23:21]};
assign col_out_78 = {u_ca_out_78[2:0],u_ca_out_77[11:3], u_ca_out_76[20:12], u_ca_out_75[23:21]};
assign col_out_79 = {u_ca_out_79[2:0],u_ca_out_78[11:3], u_ca_out_77[20:12], u_ca_out_76[23:21]};
assign col_out_80 = {u_ca_out_80[2:0],u_ca_out_79[11:3], u_ca_out_78[20:12], u_ca_out_77[23:21]};
assign col_out_81 = {u_ca_out_81[2:0],u_ca_out_80[11:3], u_ca_out_79[20:12], u_ca_out_78[23:21]};
assign col_out_82 = {u_ca_out_82[2:0],u_ca_out_81[11:3], u_ca_out_80[20:12], u_ca_out_79[23:21]};
assign col_out_83 = {u_ca_out_83[2:0],u_ca_out_82[11:3], u_ca_out_81[20:12], u_ca_out_80[23:21]};
assign col_out_84 = {u_ca_out_84[2:0],u_ca_out_83[11:3], u_ca_out_82[20:12], u_ca_out_81[23:21]};
assign col_out_85 = {u_ca_out_85[2:0],u_ca_out_84[11:3], u_ca_out_83[20:12], u_ca_out_82[23:21]};
assign col_out_86 = {u_ca_out_86[2:0],u_ca_out_85[11:3], u_ca_out_84[20:12], u_ca_out_83[23:21]};
assign col_out_87 = {u_ca_out_87[2:0],u_ca_out_86[11:3], u_ca_out_85[20:12], u_ca_out_84[23:21]};
assign col_out_88 = {u_ca_out_88[2:0],u_ca_out_87[11:3], u_ca_out_86[20:12], u_ca_out_85[23:21]};
assign col_out_89 = {u_ca_out_89[2:0],u_ca_out_88[11:3], u_ca_out_87[20:12], u_ca_out_86[23:21]};
assign col_out_90 = {u_ca_out_90[2:0],u_ca_out_89[11:3], u_ca_out_88[20:12], u_ca_out_87[23:21]};
assign col_out_91 = {u_ca_out_91[2:0],u_ca_out_90[11:3], u_ca_out_89[20:12], u_ca_out_88[23:21]};
assign col_out_92 = {u_ca_out_92[2:0],u_ca_out_91[11:3], u_ca_out_90[20:12], u_ca_out_89[23:21]};
assign col_out_93 = {u_ca_out_93[2:0],u_ca_out_92[11:3], u_ca_out_91[20:12], u_ca_out_90[23:21]};
assign col_out_94 = {u_ca_out_94[2:0],u_ca_out_93[11:3], u_ca_out_92[20:12], u_ca_out_91[23:21]};
assign col_out_95 = {u_ca_out_95[2:0],u_ca_out_94[11:3], u_ca_out_93[20:12], u_ca_out_92[23:21]};
assign col_out_96 = {u_ca_out_96[2:0],u_ca_out_95[11:3], u_ca_out_94[20:12], u_ca_out_93[23:21]};
assign col_out_97 = {u_ca_out_97[2:0],u_ca_out_96[11:3], u_ca_out_95[20:12], u_ca_out_94[23:21]};
assign col_out_98 = {u_ca_out_98[2:0],u_ca_out_97[11:3], u_ca_out_96[20:12], u_ca_out_95[23:21]};
assign col_out_99 = {u_ca_out_99[2:0],u_ca_out_98[11:3], u_ca_out_97[20:12], u_ca_out_96[23:21]};
assign col_out_100 = {u_ca_out_100[2:0],u_ca_out_99[11:3], u_ca_out_98[20:12], u_ca_out_97[23:21]};
assign col_out_101 = {u_ca_out_101[2:0],u_ca_out_100[11:3], u_ca_out_99[20:12], u_ca_out_98[23:21]};
assign col_out_102 = {u_ca_out_102[2:0],u_ca_out_101[11:3], u_ca_out_100[20:12], u_ca_out_99[23:21]};
assign col_out_103 = {u_ca_out_103[2:0],u_ca_out_102[11:3], u_ca_out_101[20:12], u_ca_out_100[23:21]};
assign col_out_104 = {u_ca_out_104[2:0],u_ca_out_103[11:3], u_ca_out_102[20:12], u_ca_out_101[23:21]};
assign col_out_105 = {u_ca_out_105[2:0],u_ca_out_104[11:3], u_ca_out_103[20:12], u_ca_out_102[23:21]};
assign col_out_106 = {u_ca_out_106[2:0],u_ca_out_105[11:3], u_ca_out_104[20:12], u_ca_out_103[23:21]};
assign col_out_107 = {u_ca_out_107[2:0],u_ca_out_106[11:3], u_ca_out_105[20:12], u_ca_out_104[23:21]};
assign col_out_108 = {u_ca_out_108[2:0],u_ca_out_107[11:3], u_ca_out_106[20:12], u_ca_out_105[23:21]};
assign col_out_109 = {u_ca_out_109[2:0],u_ca_out_108[11:3], u_ca_out_107[20:12], u_ca_out_106[23:21]};
assign col_out_110 = {u_ca_out_110[2:0],u_ca_out_109[11:3], u_ca_out_108[20:12], u_ca_out_107[23:21]};
assign col_out_111 = {u_ca_out_111[2:0],u_ca_out_110[11:3], u_ca_out_109[20:12], u_ca_out_108[23:21]};
assign col_out_112 = {u_ca_out_112[2:0],u_ca_out_111[11:3], u_ca_out_110[20:12], u_ca_out_109[23:21]};
assign col_out_113 = {u_ca_out_113[2:0],u_ca_out_112[11:3], u_ca_out_111[20:12], u_ca_out_110[23:21]};
assign col_out_114 = {u_ca_out_114[2:0],u_ca_out_113[11:3], u_ca_out_112[20:12], u_ca_out_111[23:21]};
assign col_out_115 = {u_ca_out_115[2:0],u_ca_out_114[11:3], u_ca_out_113[20:12], u_ca_out_112[23:21]};
assign col_out_116 = {u_ca_out_116[2:0],u_ca_out_115[11:3], u_ca_out_114[20:12], u_ca_out_113[23:21]};
assign col_out_117 = {u_ca_out_117[2:0],u_ca_out_116[11:3], u_ca_out_115[20:12], u_ca_out_114[23:21]};
assign col_out_118 = {u_ca_out_118[2:0],u_ca_out_117[11:3], u_ca_out_116[20:12], u_ca_out_115[23:21]};
assign col_out_119 = {u_ca_out_119[2:0],u_ca_out_118[11:3], u_ca_out_117[20:12], u_ca_out_116[23:21]};
assign col_out_120 = {u_ca_out_120[2:0],u_ca_out_119[11:3], u_ca_out_118[20:12], u_ca_out_117[23:21]};
assign col_out_121 = {u_ca_out_121[2:0],u_ca_out_120[11:3], u_ca_out_119[20:12], u_ca_out_118[23:21]};
assign col_out_122 = {u_ca_out_122[2:0],u_ca_out_121[11:3], u_ca_out_120[20:12], u_ca_out_119[23:21]};
assign col_out_123 = {u_ca_out_123[2:0],u_ca_out_122[11:3], u_ca_out_121[20:12], u_ca_out_120[23:21]};
assign col_out_124 = {u_ca_out_124[2:0],u_ca_out_123[11:3], u_ca_out_122[20:12], u_ca_out_121[23:21]};
assign col_out_125 = {u_ca_out_125[2:0],u_ca_out_124[11:3], u_ca_out_123[20:12], u_ca_out_122[23:21]};
assign col_out_126 = {u_ca_out_126[2:0],u_ca_out_125[11:3], u_ca_out_124[20:12], u_ca_out_123[23:21]};
assign col_out_127 = {u_ca_out_127[2:0],u_ca_out_126[11:3], u_ca_out_125[20:12], u_ca_out_124[23:21]};
assign col_out_128 = {u_ca_out_128[2:0],u_ca_out_127[11:3], u_ca_out_126[20:12], u_ca_out_125[23:21]};
assign col_out_129 = {u_ca_out_129[2:0],u_ca_out_128[11:3], u_ca_out_127[20:12], u_ca_out_126[23:21]};
assign col_out_130 = {u_ca_out_130[2:0],u_ca_out_129[11:3], u_ca_out_128[20:12], u_ca_out_127[23:21]};
assign col_out_131 = {u_ca_out_131[2:0],u_ca_out_130[11:3], u_ca_out_129[20:12], u_ca_out_128[23:21]};
assign col_out_132 = {u_ca_out_132[2:0],u_ca_out_131[11:3], u_ca_out_130[20:12], u_ca_out_129[23:21]};
assign col_out_133 = {u_ca_out_133[2:0],u_ca_out_132[11:3], u_ca_out_131[20:12], u_ca_out_130[23:21]};
assign col_out_134 = {u_ca_out_134[2:0],u_ca_out_133[11:3], u_ca_out_132[20:12], u_ca_out_131[23:21]};
assign col_out_135 = {u_ca_out_135[2:0],u_ca_out_134[11:3], u_ca_out_133[20:12], u_ca_out_132[23:21]};
assign col_out_136 = {u_ca_out_136[2:0],u_ca_out_135[11:3], u_ca_out_134[20:12], u_ca_out_133[23:21]};
assign col_out_137 = {u_ca_out_137[2:0],u_ca_out_136[11:3], u_ca_out_135[20:12], u_ca_out_134[23:21]};
assign col_out_138 = {u_ca_out_138[2:0],u_ca_out_137[11:3], u_ca_out_136[20:12], u_ca_out_135[23:21]};
assign col_out_139 = {u_ca_out_139[2:0],u_ca_out_138[11:3], u_ca_out_137[20:12], u_ca_out_136[23:21]};
assign col_out_140 = {u_ca_out_140[2:0],u_ca_out_139[11:3], u_ca_out_138[20:12], u_ca_out_137[23:21]};
assign col_out_141 = {u_ca_out_141[2:0],u_ca_out_140[11:3], u_ca_out_139[20:12], u_ca_out_138[23:21]};
assign col_out_142 = {u_ca_out_142[2:0],u_ca_out_141[11:3], u_ca_out_140[20:12], u_ca_out_139[23:21]};
assign col_out_143 = {u_ca_out_143[2:0],u_ca_out_142[11:3], u_ca_out_141[20:12], u_ca_out_140[23:21]};
assign col_out_144 = {u_ca_out_144[2:0],u_ca_out_143[11:3], u_ca_out_142[20:12], u_ca_out_141[23:21]};
assign col_out_145 = {u_ca_out_145[2:0],u_ca_out_144[11:3], u_ca_out_143[20:12], u_ca_out_142[23:21]};
assign col_out_146 = {u_ca_out_146[2:0],u_ca_out_145[11:3], u_ca_out_144[20:12], u_ca_out_143[23:21]};
assign col_out_147 = {u_ca_out_147[2:0],u_ca_out_146[11:3], u_ca_out_145[20:12], u_ca_out_144[23:21]};
assign col_out_148 = {u_ca_out_148[2:0],u_ca_out_147[11:3], u_ca_out_146[20:12], u_ca_out_145[23:21]};
assign col_out_149 = {u_ca_out_149[2:0],u_ca_out_148[11:3], u_ca_out_147[20:12], u_ca_out_146[23:21]};
assign col_out_150 = {u_ca_out_150[2:0],u_ca_out_149[11:3], u_ca_out_148[20:12], u_ca_out_147[23:21]};
assign col_out_151 = {u_ca_out_151[2:0],u_ca_out_150[11:3], u_ca_out_149[20:12], u_ca_out_148[23:21]};
assign col_out_152 = {u_ca_out_152[2:0],u_ca_out_151[11:3], u_ca_out_150[20:12], u_ca_out_149[23:21]};
assign col_out_153 = {u_ca_out_153[2:0],u_ca_out_152[11:3], u_ca_out_151[20:12], u_ca_out_150[23:21]};
assign col_out_154 = {u_ca_out_154[2:0],u_ca_out_153[11:3], u_ca_out_152[20:12], u_ca_out_151[23:21]};
assign col_out_155 = {u_ca_out_155[2:0],u_ca_out_154[11:3], u_ca_out_153[20:12], u_ca_out_152[23:21]};
assign col_out_156 = {u_ca_out_156[2:0],u_ca_out_155[11:3], u_ca_out_154[20:12], u_ca_out_153[23:21]};
assign col_out_157 = {u_ca_out_157[2:0],u_ca_out_156[11:3], u_ca_out_155[20:12], u_ca_out_154[23:21]};
assign col_out_158 = {u_ca_out_158[2:0],u_ca_out_157[11:3], u_ca_out_156[20:12], u_ca_out_155[23:21]};
assign col_out_159 = {u_ca_out_159[2:0],u_ca_out_158[11:3], u_ca_out_157[20:12], u_ca_out_156[23:21]};
assign col_out_160 = {u_ca_out_160[2:0],u_ca_out_159[11:3], u_ca_out_158[20:12], u_ca_out_157[23:21]};
assign col_out_161 = {u_ca_out_161[2:0],u_ca_out_160[11:3], u_ca_out_159[20:12], u_ca_out_158[23:21]};
assign col_out_162 = {u_ca_out_162[2:0],u_ca_out_161[11:3], u_ca_out_160[20:12], u_ca_out_159[23:21]};
assign col_out_163 = {u_ca_out_163[2:0],u_ca_out_162[11:3], u_ca_out_161[20:12], u_ca_out_160[23:21]};
assign col_out_164 = {u_ca_out_164[2:0],u_ca_out_163[11:3], u_ca_out_162[20:12], u_ca_out_161[23:21]};
assign col_out_165 = {u_ca_out_165[2:0],u_ca_out_164[11:3], u_ca_out_163[20:12], u_ca_out_162[23:21]};
assign col_out_166 = {u_ca_out_166[2:0],u_ca_out_165[11:3], u_ca_out_164[20:12], u_ca_out_163[23:21]};
assign col_out_167 = {u_ca_out_167[2:0],u_ca_out_166[11:3], u_ca_out_165[20:12], u_ca_out_164[23:21]};
assign col_out_168 = {u_ca_out_168[2:0],u_ca_out_167[11:3], u_ca_out_166[20:12], u_ca_out_165[23:21]};
assign col_out_169 = {u_ca_out_169[2:0],u_ca_out_168[11:3], u_ca_out_167[20:12], u_ca_out_166[23:21]};
assign col_out_170 = {u_ca_out_170[2:0],u_ca_out_169[11:3], u_ca_out_168[20:12], u_ca_out_167[23:21]};
assign col_out_171 = {u_ca_out_171[2:0],u_ca_out_170[11:3], u_ca_out_169[20:12], u_ca_out_168[23:21]};
assign col_out_172 = {u_ca_out_172[2:0],u_ca_out_171[11:3], u_ca_out_170[20:12], u_ca_out_169[23:21]};
assign col_out_173 = {u_ca_out_173[2:0],u_ca_out_172[11:3], u_ca_out_171[20:12], u_ca_out_170[23:21]};
assign col_out_174 = {u_ca_out_174[2:0],u_ca_out_173[11:3], u_ca_out_172[20:12], u_ca_out_171[23:21]};
assign col_out_175 = {u_ca_out_175[2:0],u_ca_out_174[11:3], u_ca_out_173[20:12], u_ca_out_172[23:21]};
assign col_out_176 = {u_ca_out_176[2:0],u_ca_out_175[11:3], u_ca_out_174[20:12], u_ca_out_173[23:21]};
assign col_out_177 = {u_ca_out_177[2:0],u_ca_out_176[11:3], u_ca_out_175[20:12], u_ca_out_174[23:21]};
assign col_out_178 = {u_ca_out_178[2:0],u_ca_out_177[11:3], u_ca_out_176[20:12], u_ca_out_175[23:21]};
assign col_out_179 = {u_ca_out_179[2:0],u_ca_out_178[11:3], u_ca_out_177[20:12], u_ca_out_176[23:21]};
assign col_out_180 = {u_ca_out_180[2:0],u_ca_out_179[11:3], u_ca_out_178[20:12], u_ca_out_177[23:21]};
assign col_out_181 = {u_ca_out_181[2:0],u_ca_out_180[11:3], u_ca_out_179[20:12], u_ca_out_178[23:21]};
assign col_out_182 = {u_ca_out_182[2:0],u_ca_out_181[11:3], u_ca_out_180[20:12], u_ca_out_179[23:21]};
assign col_out_183 = {u_ca_out_183[2:0],u_ca_out_182[11:3], u_ca_out_181[20:12], u_ca_out_180[23:21]};
assign col_out_184 = {u_ca_out_184[2:0],u_ca_out_183[11:3], u_ca_out_182[20:12], u_ca_out_181[23:21]};
assign col_out_185 = {u_ca_out_185[2:0],u_ca_out_184[11:3], u_ca_out_183[20:12], u_ca_out_182[23:21]};
assign col_out_186 = {u_ca_out_186[2:0],u_ca_out_185[11:3], u_ca_out_184[20:12], u_ca_out_183[23:21]};
assign col_out_187 = {u_ca_out_187[2:0],u_ca_out_186[11:3], u_ca_out_185[20:12], u_ca_out_184[23:21]};
assign col_out_188 = {u_ca_out_188[2:0],u_ca_out_187[11:3], u_ca_out_186[20:12], u_ca_out_185[23:21]};
assign col_out_189 = {u_ca_out_189[2:0],u_ca_out_188[11:3], u_ca_out_187[20:12], u_ca_out_186[23:21]};
assign col_out_190 = {u_ca_out_190[2:0],u_ca_out_189[11:3], u_ca_out_188[20:12], u_ca_out_187[23:21]};
assign col_out_191 = {u_ca_out_191[2:0],u_ca_out_190[11:3], u_ca_out_189[20:12], u_ca_out_188[23:21]};
assign col_out_192 = {u_ca_out_192[2:0],u_ca_out_191[11:3], u_ca_out_190[20:12], u_ca_out_189[23:21]};
assign col_out_193 = {u_ca_out_193[2:0],u_ca_out_192[11:3], u_ca_out_191[20:12], u_ca_out_190[23:21]};
assign col_out_194 = {u_ca_out_194[2:0],u_ca_out_193[11:3], u_ca_out_192[20:12], u_ca_out_191[23:21]};
assign col_out_195 = {u_ca_out_195[2:0],u_ca_out_194[11:3], u_ca_out_193[20:12], u_ca_out_192[23:21]};
assign col_out_196 = {u_ca_out_196[2:0],u_ca_out_195[11:3], u_ca_out_194[20:12], u_ca_out_193[23:21]};
assign col_out_197 = {u_ca_out_197[2:0],u_ca_out_196[11:3], u_ca_out_195[20:12], u_ca_out_194[23:21]};
assign col_out_198 = {u_ca_out_198[2:0],u_ca_out_197[11:3], u_ca_out_196[20:12], u_ca_out_195[23:21]};
assign col_out_199 = {u_ca_out_199[2:0],u_ca_out_198[11:3], u_ca_out_197[20:12], u_ca_out_196[23:21]};
assign col_out_200 = {u_ca_out_200[2:0],u_ca_out_199[11:3], u_ca_out_198[20:12], u_ca_out_197[23:21]};
assign col_out_201 = {u_ca_out_201[2:0],u_ca_out_200[11:3], u_ca_out_199[20:12], u_ca_out_198[23:21]};
assign col_out_202 = {u_ca_out_202[2:0],u_ca_out_201[11:3], u_ca_out_200[20:12], u_ca_out_199[23:21]};
assign col_out_203 = {u_ca_out_203[2:0],u_ca_out_202[11:3], u_ca_out_201[20:12], u_ca_out_200[23:21]};
assign col_out_204 = {u_ca_out_204[2:0],u_ca_out_203[11:3], u_ca_out_202[20:12], u_ca_out_201[23:21]};
assign col_out_205 = {u_ca_out_205[2:0],u_ca_out_204[11:3], u_ca_out_203[20:12], u_ca_out_202[23:21]};
assign col_out_206 = {u_ca_out_206[2:0],u_ca_out_205[11:3], u_ca_out_204[20:12], u_ca_out_203[23:21]};
assign col_out_207 = {u_ca_out_207[2:0],u_ca_out_206[11:3], u_ca_out_205[20:12], u_ca_out_204[23:21]};
assign col_out_208 = {u_ca_out_208[2:0],u_ca_out_207[11:3], u_ca_out_206[20:12], u_ca_out_205[23:21]};
assign col_out_209 = {u_ca_out_209[2:0],u_ca_out_208[11:3], u_ca_out_207[20:12], u_ca_out_206[23:21]};
assign col_out_210 = {u_ca_out_210[2:0],u_ca_out_209[11:3], u_ca_out_208[20:12], u_ca_out_207[23:21]};
assign col_out_211 = {u_ca_out_211[2:0],u_ca_out_210[11:3], u_ca_out_209[20:12], u_ca_out_208[23:21]};
assign col_out_212 = {u_ca_out_212[2:0],u_ca_out_211[11:3], u_ca_out_210[20:12], u_ca_out_209[23:21]};
assign col_out_213 = {u_ca_out_213[2:0],u_ca_out_212[11:3], u_ca_out_211[20:12], u_ca_out_210[23:21]};
assign col_out_214 = {u_ca_out_214[2:0],u_ca_out_213[11:3], u_ca_out_212[20:12], u_ca_out_211[23:21]};
assign col_out_215 = {u_ca_out_215[2:0],u_ca_out_214[11:3], u_ca_out_213[20:12], u_ca_out_212[23:21]};
assign col_out_216 = {u_ca_out_216[2:0],u_ca_out_215[11:3], u_ca_out_214[20:12], u_ca_out_213[23:21]};
assign col_out_217 = {u_ca_out_217[2:0],u_ca_out_216[11:3], u_ca_out_215[20:12], u_ca_out_214[23:21]};
assign col_out_218 = {u_ca_out_218[2:0],u_ca_out_217[11:3], u_ca_out_216[20:12], u_ca_out_215[23:21]};
assign col_out_219 = {u_ca_out_219[2:0],u_ca_out_218[11:3], u_ca_out_217[20:12], u_ca_out_216[23:21]};
assign col_out_220 = {u_ca_out_220[2:0],u_ca_out_219[11:3], u_ca_out_218[20:12], u_ca_out_217[23:21]};
assign col_out_221 = {u_ca_out_221[2:0],u_ca_out_220[11:3], u_ca_out_219[20:12], u_ca_out_218[23:21]};
assign col_out_222 = {u_ca_out_222[2:0],u_ca_out_221[11:3], u_ca_out_220[20:12], u_ca_out_219[23:21]};
assign col_out_223 = {u_ca_out_223[2:0],u_ca_out_222[11:3], u_ca_out_221[20:12], u_ca_out_220[23:21]};
assign col_out_224 = {u_ca_out_224[2:0],u_ca_out_223[11:3], u_ca_out_222[20:12], u_ca_out_221[23:21]};
assign col_out_225 = {u_ca_out_225[2:0],u_ca_out_224[11:3], u_ca_out_223[20:12], u_ca_out_222[23:21]};
assign col_out_226 = {u_ca_out_226[2:0],u_ca_out_225[11:3], u_ca_out_224[20:12], u_ca_out_223[23:21]};
assign col_out_227 = {u_ca_out_227[2:0],u_ca_out_226[11:3], u_ca_out_225[20:12], u_ca_out_224[23:21]};
assign col_out_228 = {u_ca_out_228[2:0],u_ca_out_227[11:3], u_ca_out_226[20:12], u_ca_out_225[23:21]};
assign col_out_229 = {u_ca_out_229[2:0],u_ca_out_228[11:3], u_ca_out_227[20:12], u_ca_out_226[23:21]};
assign col_out_230 = {u_ca_out_230[2:0],u_ca_out_229[11:3], u_ca_out_228[20:12], u_ca_out_227[23:21]};
assign col_out_231 = {u_ca_out_231[2:0],u_ca_out_230[11:3], u_ca_out_229[20:12], u_ca_out_228[23:21]};
assign col_out_232 = {u_ca_out_232[2:0],u_ca_out_231[11:3], u_ca_out_230[20:12], u_ca_out_229[23:21]};
assign col_out_233 = {u_ca_out_233[2:0],u_ca_out_232[11:3], u_ca_out_231[20:12], u_ca_out_230[23:21]};
assign col_out_234 = {u_ca_out_234[2:0],u_ca_out_233[11:3], u_ca_out_232[20:12], u_ca_out_231[23:21]};
assign col_out_235 = {u_ca_out_235[2:0],u_ca_out_234[11:3], u_ca_out_233[20:12], u_ca_out_232[23:21]};
assign col_out_236 = {u_ca_out_236[2:0],u_ca_out_235[11:3], u_ca_out_234[20:12], u_ca_out_233[23:21]};
assign col_out_237 = {u_ca_out_237[2:0],u_ca_out_236[11:3], u_ca_out_235[20:12], u_ca_out_234[23:21]};
assign col_out_238 = {u_ca_out_238[2:0],u_ca_out_237[11:3], u_ca_out_236[20:12], u_ca_out_235[23:21]};
assign col_out_239 = {u_ca_out_239[2:0],u_ca_out_238[11:3], u_ca_out_237[20:12], u_ca_out_236[23:21]};
assign col_out_240 = {u_ca_out_240[2:0],u_ca_out_239[11:3], u_ca_out_238[20:12], u_ca_out_237[23:21]};
assign col_out_241 = {u_ca_out_241[2:0],u_ca_out_240[11:3], u_ca_out_239[20:12], u_ca_out_238[23:21]};
assign col_out_242 = {u_ca_out_242[2:0],u_ca_out_241[11:3], u_ca_out_240[20:12], u_ca_out_239[23:21]};
assign col_out_243 = {u_ca_out_243[2:0],u_ca_out_242[11:3], u_ca_out_241[20:12], u_ca_out_240[23:21]};
assign col_out_244 = {u_ca_out_244[2:0],u_ca_out_243[11:3], u_ca_out_242[20:12], u_ca_out_241[23:21]};
assign col_out_245 = {u_ca_out_245[2:0],u_ca_out_244[11:3], u_ca_out_243[20:12], u_ca_out_242[23:21]};
assign col_out_246 = {u_ca_out_246[2:0],u_ca_out_245[11:3], u_ca_out_244[20:12], u_ca_out_243[23:21]};
assign col_out_247 = {u_ca_out_247[2:0],u_ca_out_246[11:3], u_ca_out_245[20:12], u_ca_out_244[23:21]};
assign col_out_248 = {u_ca_out_248[2:0],u_ca_out_247[11:3], u_ca_out_246[20:12], u_ca_out_245[23:21]};
assign col_out_249 = {u_ca_out_249[2:0],u_ca_out_248[11:3], u_ca_out_247[20:12], u_ca_out_246[23:21]};
assign col_out_250 = {u_ca_out_250[2:0],u_ca_out_249[11:3], u_ca_out_248[20:12], u_ca_out_247[23:21]};
assign col_out_251 = {u_ca_out_251[2:0],u_ca_out_250[11:3], u_ca_out_249[20:12], u_ca_out_248[23:21]};
assign col_out_252 = {u_ca_out_252[2:0],u_ca_out_251[11:3], u_ca_out_250[20:12], u_ca_out_249[23:21]};
assign col_out_253 = {u_ca_out_253[2:0],u_ca_out_252[11:3], u_ca_out_251[20:12], u_ca_out_250[23:21]};
assign col_out_254 = {u_ca_out_254[2:0],u_ca_out_253[11:3], u_ca_out_252[20:12], u_ca_out_251[23:21]};
assign col_out_255 = {u_ca_out_255[2:0],u_ca_out_254[11:3], u_ca_out_253[20:12], u_ca_out_252[23:21]};
assign col_out_256 = {u_ca_out_256[2:0],u_ca_out_255[11:3], u_ca_out_254[20:12], u_ca_out_253[23:21]};
assign col_out_257 = {u_ca_out_257[2:0],u_ca_out_256[11:3], u_ca_out_255[20:12], u_ca_out_254[23:21]};
assign col_out_258 = {u_ca_out_258[2:0],u_ca_out_257[11:3], u_ca_out_256[20:12], u_ca_out_255[23:21]};
assign col_out_259 = {u_ca_out_259[2:0],u_ca_out_258[11:3], u_ca_out_257[20:12], u_ca_out_256[23:21]};
assign col_out_260 = {u_ca_out_260[2:0],u_ca_out_259[11:3], u_ca_out_258[20:12], u_ca_out_257[23:21]};
assign col_out_261 = {u_ca_out_261[2:0],u_ca_out_260[11:3], u_ca_out_259[20:12], u_ca_out_258[23:21]};
assign col_out_262 = {u_ca_out_262[2:0],u_ca_out_261[11:3], u_ca_out_260[20:12], u_ca_out_259[23:21]};
assign col_out_263 = {u_ca_out_263[2:0],u_ca_out_262[11:3], u_ca_out_261[20:12], u_ca_out_260[23:21]};
assign col_out_264 = {u_ca_out_264[2:0],u_ca_out_263[11:3], u_ca_out_262[20:12], u_ca_out_261[23:21]};
assign col_out_265 = {u_ca_out_265[2:0],u_ca_out_264[11:3], u_ca_out_263[20:12], u_ca_out_262[23:21]};
assign col_out_266 = {u_ca_out_266[2:0],u_ca_out_265[11:3], u_ca_out_264[20:12], u_ca_out_263[23:21]};
assign col_out_267 = {u_ca_out_267[2:0],u_ca_out_266[11:3], u_ca_out_265[20:12], u_ca_out_264[23:21]};
assign col_out_268 = {u_ca_out_268[2:0],u_ca_out_267[11:3], u_ca_out_266[20:12], u_ca_out_265[23:21]};
assign col_out_269 = {u_ca_out_269[2:0],u_ca_out_268[11:3], u_ca_out_267[20:12], u_ca_out_266[23:21]};
assign col_out_270 = {u_ca_out_270[2:0],u_ca_out_269[11:3], u_ca_out_268[20:12], u_ca_out_267[23:21]};
assign col_out_271 = {u_ca_out_271[2:0],u_ca_out_270[11:3], u_ca_out_269[20:12], u_ca_out_268[23:21]};
assign col_out_272 = {u_ca_out_272[2:0],u_ca_out_271[11:3], u_ca_out_270[20:12], u_ca_out_269[23:21]};
assign col_out_273 = {u_ca_out_273[2:0],u_ca_out_272[11:3], u_ca_out_271[20:12], u_ca_out_270[23:21]};
assign col_out_274 = {u_ca_out_274[2:0],u_ca_out_273[11:3], u_ca_out_272[20:12], u_ca_out_271[23:21]};
assign col_out_275 = {u_ca_out_275[2:0],u_ca_out_274[11:3], u_ca_out_273[20:12], u_ca_out_272[23:21]};
assign col_out_276 = {u_ca_out_276[2:0],u_ca_out_275[11:3], u_ca_out_274[20:12], u_ca_out_273[23:21]};
assign col_out_277 = {u_ca_out_277[2:0],u_ca_out_276[11:3], u_ca_out_275[20:12], u_ca_out_274[23:21]};
assign col_out_278 = {u_ca_out_278[2:0],u_ca_out_277[11:3], u_ca_out_276[20:12], u_ca_out_275[23:21]};
assign col_out_279 = {u_ca_out_279[2:0],u_ca_out_278[11:3], u_ca_out_277[20:12], u_ca_out_276[23:21]};
assign col_out_280 = {u_ca_out_280[2:0],u_ca_out_279[11:3], u_ca_out_278[20:12], u_ca_out_277[23:21]};
assign col_out_281 = {u_ca_out_281[2:0],u_ca_out_280[11:3], u_ca_out_279[20:12], u_ca_out_278[23:21]};
assign col_out_282 = {u_ca_out_282[2:0],u_ca_out_281[11:3], u_ca_out_280[20:12], u_ca_out_279[23:21]};
assign col_out_283 = {u_ca_out_283[2:0],u_ca_out_282[11:3], u_ca_out_281[20:12], u_ca_out_280[23:21]};
assign col_out_284 = {u_ca_out_284[2:0],u_ca_out_283[11:3], u_ca_out_282[20:12], u_ca_out_281[23:21]};
assign col_out_285 = {u_ca_out_285[2:0],u_ca_out_284[11:3], u_ca_out_283[20:12], u_ca_out_282[23:21]};
assign col_out_286 = {u_ca_out_286[2:0],u_ca_out_285[11:3], u_ca_out_284[20:12], u_ca_out_283[23:21]};
assign col_out_287 = {u_ca_out_287[2:0],u_ca_out_286[11:3], u_ca_out_285[20:12], u_ca_out_284[23:21]};
assign col_out_288 = {u_ca_out_288[2:0],u_ca_out_287[11:3], u_ca_out_286[20:12], u_ca_out_285[23:21]};
assign col_out_289 = {u_ca_out_289[2:0],u_ca_out_288[11:3], u_ca_out_287[20:12], u_ca_out_286[23:21]};
assign col_out_290 = {u_ca_out_290[2:0],u_ca_out_289[11:3], u_ca_out_288[20:12], u_ca_out_287[23:21]};
assign col_out_291 = {u_ca_out_291[2:0],u_ca_out_290[11:3], u_ca_out_289[20:12], u_ca_out_288[23:21]};
assign col_out_292 = {u_ca_out_292[2:0],u_ca_out_291[11:3], u_ca_out_290[20:12], u_ca_out_289[23:21]};
assign col_out_293 = {u_ca_out_293[2:0],u_ca_out_292[11:3], u_ca_out_291[20:12], u_ca_out_290[23:21]};
assign col_out_294 = {u_ca_out_294[2:0],u_ca_out_293[11:3], u_ca_out_292[20:12], u_ca_out_291[23:21]};
assign col_out_295 = {u_ca_out_295[2:0],u_ca_out_294[11:3], u_ca_out_293[20:12], u_ca_out_292[23:21]};
assign col_out_296 = {u_ca_out_296[2:0],u_ca_out_295[11:3], u_ca_out_294[20:12], u_ca_out_293[23:21]};
assign col_out_297 = {u_ca_out_297[2:0],u_ca_out_296[11:3], u_ca_out_295[20:12], u_ca_out_294[23:21]};
assign col_out_298 = {u_ca_out_298[2:0],u_ca_out_297[11:3], u_ca_out_296[20:12], u_ca_out_295[23:21]};
assign col_out_299 = {u_ca_out_299[2:0],u_ca_out_298[11:3], u_ca_out_297[20:12], u_ca_out_296[23:21]};
assign col_out_300 = {u_ca_out_300[2:0],u_ca_out_299[11:3], u_ca_out_298[20:12], u_ca_out_297[23:21]};
assign col_out_301 = {u_ca_out_301[2:0],u_ca_out_300[11:3], u_ca_out_299[20:12], u_ca_out_298[23:21]};
assign col_out_302 = {u_ca_out_302[2:0],u_ca_out_301[11:3], u_ca_out_300[20:12], u_ca_out_299[23:21]};
assign col_out_303 = {u_ca_out_303[2:0],u_ca_out_302[11:3], u_ca_out_301[20:12], u_ca_out_300[23:21]};
assign col_out_304 = {u_ca_out_304[2:0],u_ca_out_303[11:3], u_ca_out_302[20:12], u_ca_out_301[23:21]};
assign col_out_305 = {u_ca_out_305[2:0],u_ca_out_304[11:3], u_ca_out_303[20:12], u_ca_out_302[23:21]};
assign col_out_306 = {u_ca_out_306[2:0],u_ca_out_305[11:3], u_ca_out_304[20:12], u_ca_out_303[23:21]};
assign col_out_307 = {u_ca_out_307[2:0],u_ca_out_306[11:3], u_ca_out_305[20:12], u_ca_out_304[23:21]};
assign col_out_308 = {u_ca_out_308[2:0],u_ca_out_307[11:3], u_ca_out_306[20:12], u_ca_out_305[23:21]};
assign col_out_309 = {u_ca_out_309[2:0],u_ca_out_308[11:3], u_ca_out_307[20:12], u_ca_out_306[23:21]};
assign col_out_310 = {u_ca_out_310[2:0],u_ca_out_309[11:3], u_ca_out_308[20:12], u_ca_out_307[23:21]};
assign col_out_311 = {u_ca_out_311[2:0],u_ca_out_310[11:3], u_ca_out_309[20:12], u_ca_out_308[23:21]};
assign col_out_312 = {u_ca_out_312[2:0],u_ca_out_311[11:3], u_ca_out_310[20:12], u_ca_out_309[23:21]};
assign col_out_313 = {u_ca_out_313[2:0],u_ca_out_312[11:3], u_ca_out_311[20:12], u_ca_out_310[23:21]};
assign col_out_314 = {u_ca_out_314[2:0],u_ca_out_313[11:3], u_ca_out_312[20:12], u_ca_out_311[23:21]};
assign col_out_315 = {u_ca_out_315[2:0],u_ca_out_314[11:3], u_ca_out_313[20:12], u_ca_out_312[23:21]};
assign col_out_316 = {u_ca_out_316[2:0],u_ca_out_315[11:3], u_ca_out_314[20:12], u_ca_out_313[23:21]};
assign col_out_317 = {u_ca_out_317[2:0],u_ca_out_316[11:3], u_ca_out_315[20:12], u_ca_out_314[23:21]};
assign col_out_318 = {u_ca_out_318[2:0],u_ca_out_317[11:3], u_ca_out_316[20:12], u_ca_out_315[23:21]};
assign col_out_319 = {u_ca_out_319[2:0],u_ca_out_318[11:3], u_ca_out_317[20:12], u_ca_out_316[23:21]};
assign col_out_320 = {u_ca_out_320[2:0],u_ca_out_319[11:3], u_ca_out_318[20:12], u_ca_out_317[23:21]};
assign col_out_321 = {u_ca_out_321[2:0],u_ca_out_320[11:3], u_ca_out_319[20:12], u_ca_out_318[23:21]};
assign col_out_322 = {u_ca_out_322[2:0],u_ca_out_321[11:3], u_ca_out_320[20:12], u_ca_out_319[23:21]};
assign col_out_323 = {u_ca_out_323[2:0],u_ca_out_322[11:3], u_ca_out_321[20:12], u_ca_out_320[23:21]};
assign col_out_324 = {u_ca_out_324[2:0],u_ca_out_323[11:3], u_ca_out_322[20:12], u_ca_out_321[23:21]};
assign col_out_325 = {u_ca_out_325[2:0],u_ca_out_324[11:3], u_ca_out_323[20:12], u_ca_out_322[23:21]};
assign col_out_326 = {u_ca_out_326[2:0],u_ca_out_325[11:3], u_ca_out_324[20:12], u_ca_out_323[23:21]};
assign col_out_327 = {u_ca_out_327[2:0],u_ca_out_326[11:3], u_ca_out_325[20:12], u_ca_out_324[23:21]};
assign col_out_328 = {u_ca_out_328[2:0],u_ca_out_327[11:3], u_ca_out_326[20:12], u_ca_out_325[23:21]};
assign col_out_329 = {u_ca_out_329[2:0],u_ca_out_328[11:3], u_ca_out_327[20:12], u_ca_out_326[23:21]};
assign col_out_330 = {u_ca_out_330[2:0],u_ca_out_329[11:3], u_ca_out_328[20:12], u_ca_out_327[23:21]};
assign col_out_331 = {u_ca_out_331[2:0],u_ca_out_330[11:3], u_ca_out_329[20:12], u_ca_out_328[23:21]};
assign col_out_332 = {u_ca_out_332[2:0],u_ca_out_331[11:3], u_ca_out_330[20:12], u_ca_out_329[23:21]};
assign col_out_333 = {u_ca_out_333[2:0],u_ca_out_332[11:3], u_ca_out_331[20:12], u_ca_out_330[23:21]};
assign col_out_334 = {u_ca_out_334[2:0],u_ca_out_333[11:3], u_ca_out_332[20:12], u_ca_out_331[23:21]};
assign col_out_335 = {u_ca_out_335[2:0],u_ca_out_334[11:3], u_ca_out_333[20:12], u_ca_out_332[23:21]};
assign col_out_336 = {u_ca_out_336[2:0],u_ca_out_335[11:3], u_ca_out_334[20:12], u_ca_out_333[23:21]};
assign col_out_337 = {u_ca_out_337[2:0],u_ca_out_336[11:3], u_ca_out_335[20:12], u_ca_out_334[23:21]};
assign col_out_338 = {u_ca_out_338[2:0],u_ca_out_337[11:3], u_ca_out_336[20:12], u_ca_out_335[23:21]};
assign col_out_339 = {u_ca_out_339[2:0],u_ca_out_338[11:3], u_ca_out_337[20:12], u_ca_out_336[23:21]};
assign col_out_340 = {u_ca_out_340[2:0],u_ca_out_339[11:3], u_ca_out_338[20:12], u_ca_out_337[23:21]};
assign col_out_341 = {u_ca_out_341[2:0],u_ca_out_340[11:3], u_ca_out_339[20:12], u_ca_out_338[23:21]};
assign col_out_342 = {u_ca_out_342[2:0],u_ca_out_341[11:3], u_ca_out_340[20:12], u_ca_out_339[23:21]};
assign col_out_343 = {u_ca_out_343[2:0],u_ca_out_342[11:3], u_ca_out_341[20:12], u_ca_out_340[23:21]};
assign col_out_344 = {u_ca_out_344[2:0],u_ca_out_343[11:3], u_ca_out_342[20:12], u_ca_out_341[23:21]};
assign col_out_345 = {u_ca_out_345[2:0],u_ca_out_344[11:3], u_ca_out_343[20:12], u_ca_out_342[23:21]};
assign col_out_346 = {u_ca_out_346[2:0],u_ca_out_345[11:3], u_ca_out_344[20:12], u_ca_out_343[23:21]};
assign col_out_347 = {u_ca_out_347[2:0],u_ca_out_346[11:3], u_ca_out_345[20:12], u_ca_out_344[23:21]};
assign col_out_348 = {u_ca_out_348[2:0],u_ca_out_347[11:3], u_ca_out_346[20:12], u_ca_out_345[23:21]};
assign col_out_349 = {u_ca_out_349[2:0],u_ca_out_348[11:3], u_ca_out_347[20:12], u_ca_out_346[23:21]};
assign col_out_350 = {u_ca_out_350[2:0],u_ca_out_349[11:3], u_ca_out_348[20:12], u_ca_out_347[23:21]};
assign col_out_351 = {u_ca_out_351[2:0],u_ca_out_350[11:3], u_ca_out_349[20:12], u_ca_out_348[23:21]};
assign col_out_352 = {u_ca_out_352[2:0],u_ca_out_351[11:3], u_ca_out_350[20:12], u_ca_out_349[23:21]};
assign col_out_353 = {u_ca_out_353[2:0],u_ca_out_352[11:3], u_ca_out_351[20:12], u_ca_out_350[23:21]};
assign col_out_354 = {u_ca_out_354[2:0],u_ca_out_353[11:3], u_ca_out_352[20:12], u_ca_out_351[23:21]};
assign col_out_355 = {u_ca_out_355[2:0],u_ca_out_354[11:3], u_ca_out_353[20:12], u_ca_out_352[23:21]};
assign col_out_356 = {u_ca_out_356[2:0],u_ca_out_355[11:3], u_ca_out_354[20:12], u_ca_out_353[23:21]};
assign col_out_357 = {u_ca_out_357[2:0],u_ca_out_356[11:3], u_ca_out_355[20:12], u_ca_out_354[23:21]};
assign col_out_358 = {u_ca_out_358[2:0],u_ca_out_357[11:3], u_ca_out_356[20:12], u_ca_out_355[23:21]};
assign col_out_359 = {u_ca_out_359[2:0],u_ca_out_358[11:3], u_ca_out_357[20:12], u_ca_out_356[23:21]};
assign col_out_360 = {u_ca_out_360[2:0],u_ca_out_359[11:3], u_ca_out_358[20:12], u_ca_out_357[23:21]};
assign col_out_361 = {u_ca_out_361[2:0],u_ca_out_360[11:3], u_ca_out_359[20:12], u_ca_out_358[23:21]};
assign col_out_362 = {u_ca_out_362[2:0],u_ca_out_361[11:3], u_ca_out_360[20:12], u_ca_out_359[23:21]};
assign col_out_363 = {u_ca_out_363[2:0],u_ca_out_362[11:3], u_ca_out_361[20:12], u_ca_out_360[23:21]};
assign col_out_364 = {u_ca_out_364[2:0],u_ca_out_363[11:3], u_ca_out_362[20:12], u_ca_out_361[23:21]};
assign col_out_365 = {u_ca_out_365[2:0],u_ca_out_364[11:3], u_ca_out_363[20:12], u_ca_out_362[23:21]};
assign col_out_366 = {u_ca_out_366[2:0],u_ca_out_365[11:3], u_ca_out_364[20:12], u_ca_out_363[23:21]};
assign col_out_367 = {u_ca_out_367[2:0],u_ca_out_366[11:3], u_ca_out_365[20:12], u_ca_out_364[23:21]};
assign col_out_368 = {u_ca_out_368[2:0],u_ca_out_367[11:3], u_ca_out_366[20:12], u_ca_out_365[23:21]};
assign col_out_369 = {u_ca_out_369[2:0],u_ca_out_368[11:3], u_ca_out_367[20:12], u_ca_out_366[23:21]};
assign col_out_370 = {u_ca_out_370[2:0],u_ca_out_369[11:3], u_ca_out_368[20:12], u_ca_out_367[23:21]};
assign col_out_371 = {u_ca_out_371[2:0],u_ca_out_370[11:3], u_ca_out_369[20:12], u_ca_out_368[23:21]};
assign col_out_372 = {u_ca_out_372[2:0],u_ca_out_371[11:3], u_ca_out_370[20:12], u_ca_out_369[23:21]};
assign col_out_373 = {u_ca_out_373[2:0],u_ca_out_372[11:3], u_ca_out_371[20:12], u_ca_out_370[23:21]};
assign col_out_374 = {u_ca_out_374[2:0],u_ca_out_373[11:3], u_ca_out_372[20:12], u_ca_out_371[23:21]};
assign col_out_375 = {u_ca_out_375[2:0],u_ca_out_374[11:3], u_ca_out_373[20:12], u_ca_out_372[23:21]};
assign col_out_376 = {u_ca_out_376[2:0],u_ca_out_375[11:3], u_ca_out_374[20:12], u_ca_out_373[23:21]};
assign col_out_377 = {u_ca_out_377[2:0],u_ca_out_376[11:3], u_ca_out_375[20:12], u_ca_out_374[23:21]};
assign col_out_378 = {u_ca_out_378[2:0],u_ca_out_377[11:3], u_ca_out_376[20:12], u_ca_out_375[23:21]};
assign col_out_379 = {u_ca_out_379[2:0],u_ca_out_378[11:3], u_ca_out_377[20:12], u_ca_out_376[23:21]};
assign col_out_380 = {u_ca_out_380[2:0],u_ca_out_379[11:3], u_ca_out_378[20:12], u_ca_out_377[23:21]};
assign col_out_381 = {u_ca_out_381[2:0],u_ca_out_380[11:3], u_ca_out_379[20:12], u_ca_out_378[23:21]};
assign col_out_382 = {u_ca_out_382[2:0],u_ca_out_381[11:3], u_ca_out_380[20:12], u_ca_out_379[23:21]};
assign col_out_383 = {u_ca_out_383[2:0],u_ca_out_382[11:3], u_ca_out_381[20:12], u_ca_out_380[23:21]};
assign col_out_384 = {u_ca_out_384[2:0],u_ca_out_383[11:3], u_ca_out_382[20:12], u_ca_out_381[23:21]};
assign col_out_385 = {u_ca_out_385[2:0],u_ca_out_384[11:3], u_ca_out_383[20:12], u_ca_out_382[23:21]};
assign col_out_386 = {u_ca_out_386[2:0],u_ca_out_385[11:3], u_ca_out_384[20:12], u_ca_out_383[23:21]};
assign col_out_387 = {u_ca_out_387[2:0],u_ca_out_386[11:3], u_ca_out_385[20:12], u_ca_out_384[23:21]};
assign col_out_388 = {u_ca_out_388[2:0],u_ca_out_387[11:3], u_ca_out_386[20:12], u_ca_out_385[23:21]};
assign col_out_389 = {u_ca_out_389[2:0],u_ca_out_388[11:3], u_ca_out_387[20:12], u_ca_out_386[23:21]};
assign col_out_390 = {u_ca_out_390[2:0],u_ca_out_389[11:3], u_ca_out_388[20:12], u_ca_out_387[23:21]};
assign col_out_391 = {u_ca_out_391[2:0],u_ca_out_390[11:3], u_ca_out_389[20:12], u_ca_out_388[23:21]};
assign col_out_392 = {u_ca_out_392[2:0],u_ca_out_391[11:3], u_ca_out_390[20:12], u_ca_out_389[23:21]};
assign col_out_393 = {u_ca_out_393[2:0],u_ca_out_392[11:3], u_ca_out_391[20:12], u_ca_out_390[23:21]};
assign col_out_394 = {u_ca_out_394[2:0],u_ca_out_393[11:3], u_ca_out_392[20:12], u_ca_out_391[23:21]};
assign col_out_395 = {u_ca_out_395[2:0],u_ca_out_394[11:3], u_ca_out_393[20:12], u_ca_out_392[23:21]};
assign col_out_396 = {u_ca_out_396[2:0],u_ca_out_395[11:3], u_ca_out_394[20:12], u_ca_out_393[23:21]};
assign col_out_397 = {u_ca_out_397[2:0],u_ca_out_396[11:3], u_ca_out_395[20:12], u_ca_out_394[23:21]};
assign col_out_398 = {u_ca_out_398[2:0],u_ca_out_397[11:3], u_ca_out_396[20:12], u_ca_out_395[23:21]};
assign col_out_399 = {u_ca_out_399[2:0],u_ca_out_398[11:3], u_ca_out_397[20:12], u_ca_out_396[23:21]};
assign col_out_400 = {u_ca_out_400[2:0],u_ca_out_399[11:3], u_ca_out_398[20:12], u_ca_out_397[23:21]};
assign col_out_401 = {u_ca_out_401[2:0],u_ca_out_400[11:3], u_ca_out_399[20:12], u_ca_out_398[23:21]};
assign col_out_402 = {u_ca_out_402[2:0],u_ca_out_401[11:3], u_ca_out_400[20:12], u_ca_out_399[23:21]};
assign col_out_403 = {u_ca_out_403[2:0],u_ca_out_402[11:3], u_ca_out_401[20:12], u_ca_out_400[23:21]};
assign col_out_404 = {u_ca_out_404[2:0],u_ca_out_403[11:3], u_ca_out_402[20:12], u_ca_out_401[23:21]};
assign col_out_405 = {u_ca_out_405[2:0],u_ca_out_404[11:3], u_ca_out_403[20:12], u_ca_out_402[23:21]};
assign col_out_406 = {u_ca_out_406[2:0],u_ca_out_405[11:3], u_ca_out_404[20:12], u_ca_out_403[23:21]};
assign col_out_407 = {u_ca_out_407[2:0],u_ca_out_406[11:3], u_ca_out_405[20:12], u_ca_out_404[23:21]};
assign col_out_408 = {u_ca_out_408[2:0],u_ca_out_407[11:3], u_ca_out_406[20:12], u_ca_out_405[23:21]};
assign col_out_409 = {u_ca_out_409[2:0],u_ca_out_408[11:3], u_ca_out_407[20:12], u_ca_out_406[23:21]};
assign col_out_410 = {u_ca_out_410[2:0],u_ca_out_409[11:3], u_ca_out_408[20:12], u_ca_out_407[23:21]};
assign col_out_411 = {u_ca_out_411[2:0],u_ca_out_410[11:3], u_ca_out_409[20:12], u_ca_out_408[23:21]};
assign col_out_412 = {u_ca_out_412[2:0],u_ca_out_411[11:3], u_ca_out_410[20:12], u_ca_out_409[23:21]};
assign col_out_413 = {u_ca_out_413[2:0],u_ca_out_412[11:3], u_ca_out_411[20:12], u_ca_out_410[23:21]};
assign col_out_414 = {u_ca_out_414[2:0],u_ca_out_413[11:3], u_ca_out_412[20:12], u_ca_out_411[23:21]};
assign col_out_415 = {u_ca_out_415[2:0],u_ca_out_414[11:3], u_ca_out_413[20:12], u_ca_out_412[23:21]};
assign col_out_416 = {u_ca_out_416[2:0],u_ca_out_415[11:3], u_ca_out_414[20:12], u_ca_out_413[23:21]};
assign col_out_417 = {u_ca_out_417[2:0],u_ca_out_416[11:3], u_ca_out_415[20:12], u_ca_out_414[23:21]};
assign col_out_418 = {u_ca_out_418[2:0],u_ca_out_417[11:3], u_ca_out_416[20:12], u_ca_out_415[23:21]};
assign col_out_419 = {u_ca_out_419[2:0],u_ca_out_418[11:3], u_ca_out_417[20:12], u_ca_out_416[23:21]};
assign col_out_420 = {u_ca_out_420[2:0],u_ca_out_419[11:3], u_ca_out_418[20:12], u_ca_out_417[23:21]};
assign col_out_421 = {u_ca_out_421[2:0],u_ca_out_420[11:3], u_ca_out_419[20:12], u_ca_out_418[23:21]};
assign col_out_422 = {u_ca_out_422[2:0],u_ca_out_421[11:3], u_ca_out_420[20:12], u_ca_out_419[23:21]};
assign col_out_423 = {u_ca_out_423[2:0],u_ca_out_422[11:3], u_ca_out_421[20:12], u_ca_out_420[23:21]};
assign col_out_424 = {u_ca_out_424[2:0],u_ca_out_423[11:3], u_ca_out_422[20:12], u_ca_out_421[23:21]};
assign col_out_425 = {u_ca_out_425[2:0],u_ca_out_424[11:3], u_ca_out_423[20:12], u_ca_out_422[23:21]};
assign col_out_426 = {u_ca_out_426[2:0],u_ca_out_425[11:3], u_ca_out_424[20:12], u_ca_out_423[23:21]};
assign col_out_427 = {u_ca_out_427[2:0],u_ca_out_426[11:3], u_ca_out_425[20:12], u_ca_out_424[23:21]};
assign col_out_428 = {u_ca_out_428[2:0],u_ca_out_427[11:3], u_ca_out_426[20:12], u_ca_out_425[23:21]};
assign col_out_429 = {u_ca_out_429[2:0],u_ca_out_428[11:3], u_ca_out_427[20:12], u_ca_out_426[23:21]};
assign col_out_430 = {u_ca_out_430[2:0],u_ca_out_429[11:3], u_ca_out_428[20:12], u_ca_out_427[23:21]};
assign col_out_431 = {u_ca_out_431[2:0],u_ca_out_430[11:3], u_ca_out_429[20:12], u_ca_out_428[23:21]};
assign col_out_432 = {u_ca_out_432[2:0],u_ca_out_431[11:3], u_ca_out_430[20:12], u_ca_out_429[23:21]};
assign col_out_433 = {u_ca_out_433[2:0],u_ca_out_432[11:3], u_ca_out_431[20:12], u_ca_out_430[23:21]};
assign col_out_434 = {u_ca_out_434[2:0],u_ca_out_433[11:3], u_ca_out_432[20:12], u_ca_out_431[23:21]};
assign col_out_435 = {u_ca_out_435[2:0],u_ca_out_434[11:3], u_ca_out_433[20:12], u_ca_out_432[23:21]};
assign col_out_436 = {u_ca_out_436[2:0],u_ca_out_435[11:3], u_ca_out_434[20:12], u_ca_out_433[23:21]};
assign col_out_437 = {u_ca_out_437[2:0],u_ca_out_436[11:3], u_ca_out_435[20:12], u_ca_out_434[23:21]};
assign col_out_438 = {u_ca_out_438[2:0],u_ca_out_437[11:3], u_ca_out_436[20:12], u_ca_out_435[23:21]};
assign col_out_439 = {u_ca_out_439[2:0],u_ca_out_438[11:3], u_ca_out_437[20:12], u_ca_out_436[23:21]};
assign col_out_440 = {u_ca_out_440[2:0],u_ca_out_439[11:3], u_ca_out_438[20:12], u_ca_out_437[23:21]};
assign col_out_441 = {u_ca_out_441[2:0],u_ca_out_440[11:3], u_ca_out_439[20:12], u_ca_out_438[23:21]};
assign col_out_442 = {u_ca_out_442[2:0],u_ca_out_441[11:3], u_ca_out_440[20:12], u_ca_out_439[23:21]};
assign col_out_443 = {u_ca_out_443[2:0],u_ca_out_442[11:3], u_ca_out_441[20:12], u_ca_out_440[23:21]};
assign col_out_444 = {u_ca_out_444[2:0],u_ca_out_443[11:3], u_ca_out_442[20:12], u_ca_out_441[23:21]};
assign col_out_445 = {u_ca_out_445[2:0],u_ca_out_444[11:3], u_ca_out_443[20:12], u_ca_out_442[23:21]};
assign col_out_446 = {u_ca_out_446[2:0],u_ca_out_445[11:3], u_ca_out_444[20:12], u_ca_out_443[23:21]};
assign col_out_447 = {u_ca_out_447[2:0],u_ca_out_446[11:3], u_ca_out_445[20:12], u_ca_out_444[23:21]};
assign col_out_448 = {u_ca_out_448[2:0],u_ca_out_447[11:3], u_ca_out_446[20:12], u_ca_out_445[23:21]};
assign col_out_449 = {u_ca_out_449[2:0],u_ca_out_448[11:3], u_ca_out_447[20:12], u_ca_out_446[23:21]};
assign col_out_450 = {u_ca_out_450[2:0],u_ca_out_449[11:3], u_ca_out_448[20:12], u_ca_out_447[23:21]};
assign col_out_451 = {u_ca_out_451[2:0],u_ca_out_450[11:3], u_ca_out_449[20:12], u_ca_out_448[23:21]};
assign col_out_452 = {u_ca_out_452[2:0],u_ca_out_451[11:3], u_ca_out_450[20:12], u_ca_out_449[23:21]};
assign col_out_453 = {u_ca_out_453[2:0],u_ca_out_452[11:3], u_ca_out_451[20:12], u_ca_out_450[23:21]};
assign col_out_454 = {u_ca_out_454[2:0],u_ca_out_453[11:3], u_ca_out_452[20:12], u_ca_out_451[23:21]};
assign col_out_455 = {u_ca_out_455[2:0],u_ca_out_454[11:3], u_ca_out_453[20:12], u_ca_out_452[23:21]};
assign col_out_456 = {u_ca_out_456[2:0],u_ca_out_455[11:3], u_ca_out_454[20:12], u_ca_out_453[23:21]};
assign col_out_457 = {u_ca_out_457[2:0],u_ca_out_456[11:3], u_ca_out_455[20:12], u_ca_out_454[23:21]};
assign col_out_458 = {u_ca_out_458[2:0],u_ca_out_457[11:3], u_ca_out_456[20:12], u_ca_out_455[23:21]};
assign col_out_459 = {u_ca_out_459[2:0],u_ca_out_458[11:3], u_ca_out_457[20:12], u_ca_out_456[23:21]};
assign col_out_460 = {u_ca_out_460[2:0],u_ca_out_459[11:3], u_ca_out_458[20:12], u_ca_out_457[23:21]};
assign col_out_461 = {u_ca_out_461[2:0],u_ca_out_460[11:3], u_ca_out_459[20:12], u_ca_out_458[23:21]};
assign col_out_462 = {u_ca_out_462[2:0],u_ca_out_461[11:3], u_ca_out_460[20:12], u_ca_out_459[23:21]};
assign col_out_463 = {u_ca_out_463[2:0],u_ca_out_462[11:3], u_ca_out_461[20:12], u_ca_out_460[23:21]};
assign col_out_464 = {u_ca_out_464[2:0],u_ca_out_463[11:3], u_ca_out_462[20:12], u_ca_out_461[23:21]};
assign col_out_465 = {u_ca_out_465[2:0],u_ca_out_464[11:3], u_ca_out_463[20:12], u_ca_out_462[23:21]};
assign col_out_466 = {u_ca_out_466[2:0],u_ca_out_465[11:3], u_ca_out_464[20:12], u_ca_out_463[23:21]};
assign col_out_467 = {u_ca_out_467[2:0],u_ca_out_466[11:3], u_ca_out_465[20:12], u_ca_out_464[23:21]};
assign col_out_468 = {u_ca_out_468[2:0],u_ca_out_467[11:3], u_ca_out_466[20:12], u_ca_out_465[23:21]};
assign col_out_469 = {u_ca_out_469[2:0],u_ca_out_468[11:3], u_ca_out_467[20:12], u_ca_out_466[23:21]};
assign col_out_470 = {u_ca_out_470[2:0],u_ca_out_469[11:3], u_ca_out_468[20:12], u_ca_out_467[23:21]};
assign col_out_471 = {u_ca_out_471[2:0],u_ca_out_470[11:3], u_ca_out_469[20:12], u_ca_out_468[23:21]};
assign col_out_472 = {u_ca_out_472[2:0],u_ca_out_471[11:3], u_ca_out_470[20:12], u_ca_out_469[23:21]};
assign col_out_473 = {u_ca_out_473[2:0],u_ca_out_472[11:3], u_ca_out_471[20:12], u_ca_out_470[23:21]};
assign col_out_474 = {u_ca_out_474[2:0],u_ca_out_473[11:3], u_ca_out_472[20:12], u_ca_out_471[23:21]};
assign col_out_475 = {u_ca_out_475[2:0],u_ca_out_474[11:3], u_ca_out_473[20:12], u_ca_out_472[23:21]};
assign col_out_476 = {u_ca_out_476[2:0],u_ca_out_475[11:3], u_ca_out_474[20:12], u_ca_out_473[23:21]};
assign col_out_477 = {u_ca_out_477[2:0],u_ca_out_476[11:3], u_ca_out_475[20:12], u_ca_out_474[23:21]};
assign col_out_478 = {u_ca_out_478[2:0],u_ca_out_477[11:3], u_ca_out_476[20:12], u_ca_out_475[23:21]};
assign col_out_479 = {u_ca_out_479[2:0],u_ca_out_478[11:3], u_ca_out_477[20:12], u_ca_out_476[23:21]};
assign col_out_480 = {u_ca_out_480[2:0],u_ca_out_479[11:3], u_ca_out_478[20:12], u_ca_out_477[23:21]};
assign col_out_481 = {u_ca_out_481[2:0],u_ca_out_480[11:3], u_ca_out_479[20:12], u_ca_out_478[23:21]};
assign col_out_482 = {u_ca_out_482[2:0],u_ca_out_481[11:3], u_ca_out_480[20:12], u_ca_out_479[23:21]};
assign col_out_483 = {u_ca_out_483[2:0],u_ca_out_482[11:3], u_ca_out_481[20:12], u_ca_out_480[23:21]};
assign col_out_484 = {u_ca_out_484[2:0],u_ca_out_483[11:3], u_ca_out_482[20:12], u_ca_out_481[23:21]};
assign col_out_485 = {u_ca_out_485[2:0],u_ca_out_484[11:3], u_ca_out_483[20:12], u_ca_out_482[23:21]};
assign col_out_486 = {u_ca_out_486[2:0],u_ca_out_485[11:3], u_ca_out_484[20:12], u_ca_out_483[23:21]};
assign col_out_487 = {u_ca_out_487[2:0],u_ca_out_486[11:3], u_ca_out_485[20:12], u_ca_out_484[23:21]};
assign col_out_488 = {u_ca_out_488[2:0],u_ca_out_487[11:3], u_ca_out_486[20:12], u_ca_out_485[23:21]};
assign col_out_489 = {u_ca_out_489[2:0],u_ca_out_488[11:3], u_ca_out_487[20:12], u_ca_out_486[23:21]};
assign col_out_490 = {u_ca_out_490[2:0],u_ca_out_489[11:3], u_ca_out_488[20:12], u_ca_out_487[23:21]};
assign col_out_491 = {u_ca_out_491[2:0],u_ca_out_490[11:3], u_ca_out_489[20:12], u_ca_out_488[23:21]};
assign col_out_492 = {u_ca_out_492[2:0],u_ca_out_491[11:3], u_ca_out_490[20:12], u_ca_out_489[23:21]};
assign col_out_493 = {u_ca_out_493[2:0],u_ca_out_492[11:3], u_ca_out_491[20:12], u_ca_out_490[23:21]};
assign col_out_494 = {u_ca_out_494[2:0],u_ca_out_493[11:3], u_ca_out_492[20:12], u_ca_out_491[23:21]};
assign col_out_495 = {u_ca_out_495[2:0],u_ca_out_494[11:3], u_ca_out_493[20:12], u_ca_out_492[23:21]};
assign col_out_496 = {u_ca_out_496[2:0],u_ca_out_495[11:3], u_ca_out_494[20:12], u_ca_out_493[23:21]};
assign col_out_497 = {u_ca_out_497[2:0],u_ca_out_496[11:3], u_ca_out_495[20:12], u_ca_out_494[23:21]};
assign col_out_498 = {u_ca_out_498[2:0],u_ca_out_497[11:3], u_ca_out_496[20:12], u_ca_out_495[23:21]};
assign col_out_499 = {u_ca_out_499[2:0],u_ca_out_498[11:3], u_ca_out_497[20:12], u_ca_out_496[23:21]};
assign col_out_500 = {u_ca_out_500[2:0],u_ca_out_499[11:3], u_ca_out_498[20:12], u_ca_out_497[23:21]};
assign col_out_501 = {u_ca_out_501[2:0],u_ca_out_500[11:3], u_ca_out_499[20:12], u_ca_out_498[23:21]};
assign col_out_502 = {u_ca_out_502[2:0],u_ca_out_501[11:3], u_ca_out_500[20:12], u_ca_out_499[23:21]};
assign col_out_503 = {u_ca_out_503[2:0],u_ca_out_502[11:3], u_ca_out_501[20:12], u_ca_out_500[23:21]};
assign col_out_504 = {u_ca_out_504[2:0],u_ca_out_503[11:3], u_ca_out_502[20:12], u_ca_out_501[23:21]};
assign col_out_505 = {u_ca_out_505[2:0],u_ca_out_504[11:3], u_ca_out_503[20:12], u_ca_out_502[23:21]};
assign col_out_506 = {u_ca_out_506[2:0],u_ca_out_505[11:3], u_ca_out_504[20:12], u_ca_out_503[23:21]};
assign col_out_507 = {u_ca_out_507[2:0],u_ca_out_506[11:3], u_ca_out_505[20:12], u_ca_out_504[23:21]};
assign col_out_508 = {u_ca_out_508[2:0],u_ca_out_507[11:3], u_ca_out_506[20:12], u_ca_out_505[23:21]};
assign col_out_509 = {u_ca_out_509[2:0],u_ca_out_508[11:3], u_ca_out_507[20:12], u_ca_out_506[23:21]};
assign col_out_510 = {u_ca_out_510[2:0],u_ca_out_509[11:3], u_ca_out_508[20:12], u_ca_out_507[23:21]};
assign col_out_511 = {u_ca_out_511[2:0],u_ca_out_510[11:3], u_ca_out_509[20:12], u_ca_out_508[23:21]};
assign col_out_512 = {u_ca_out_512[2:0],u_ca_out_511[11:3], u_ca_out_510[20:12], u_ca_out_509[23:21]};
assign col_out_513 = {u_ca_out_513[2:0],u_ca_out_512[11:3], u_ca_out_511[20:12], u_ca_out_510[23:21]};
assign col_out_514 = {u_ca_out_514[2:0],u_ca_out_513[11:3], u_ca_out_512[20:12], u_ca_out_511[23:21]};
assign col_out_515 = {u_ca_out_515[2:0],u_ca_out_514[11:3], u_ca_out_513[20:12], u_ca_out_512[23:21]};
assign col_out_516 = {u_ca_out_516[2:0],u_ca_out_515[11:3], u_ca_out_514[20:12], u_ca_out_513[23:21]};
assign col_out_517 = {u_ca_out_517[2:0],u_ca_out_516[11:3], u_ca_out_515[20:12], u_ca_out_514[23:21]};
assign col_out_518 = {u_ca_out_518[2:0],u_ca_out_517[11:3], u_ca_out_516[20:12], u_ca_out_515[23:21]};
assign col_out_519 = {u_ca_out_519[2:0],u_ca_out_518[11:3], u_ca_out_517[20:12], u_ca_out_516[23:21]};
assign col_out_520 = {u_ca_out_520[2:0],u_ca_out_519[11:3], u_ca_out_518[20:12], u_ca_out_517[23:21]};
assign col_out_521 = {u_ca_out_521[2:0],u_ca_out_520[11:3], u_ca_out_519[20:12], u_ca_out_518[23:21]};
assign col_out_522 = {u_ca_out_522[2:0],u_ca_out_521[11:3], u_ca_out_520[20:12], u_ca_out_519[23:21]};
assign col_out_523 = {u_ca_out_523[2:0],u_ca_out_522[11:3], u_ca_out_521[20:12], u_ca_out_520[23:21]};
assign col_out_524 = {u_ca_out_524[2:0],u_ca_out_523[11:3], u_ca_out_522[20:12], u_ca_out_521[23:21]};
assign col_out_525 = {u_ca_out_525[2:0],u_ca_out_524[11:3], u_ca_out_523[20:12], u_ca_out_522[23:21]};
assign col_out_526 = {u_ca_out_526[2:0],u_ca_out_525[11:3], u_ca_out_524[20:12], u_ca_out_523[23:21]};
assign col_out_527 = {u_ca_out_527[2:0],u_ca_out_526[11:3], u_ca_out_525[20:12], u_ca_out_524[23:21]};
assign col_out_528 = {u_ca_out_528[2:0],u_ca_out_527[11:3], u_ca_out_526[20:12], u_ca_out_525[23:21]};
assign col_out_529 = {u_ca_out_529[2:0],u_ca_out_528[11:3], u_ca_out_527[20:12], u_ca_out_526[23:21]};
assign col_out_530 = {u_ca_out_530[2:0],u_ca_out_529[11:3], u_ca_out_528[20:12], u_ca_out_527[23:21]};
assign col_out_531 = {u_ca_out_531[2:0],u_ca_out_530[11:3], u_ca_out_529[20:12], u_ca_out_528[23:21]};
assign col_out_532 = {u_ca_out_532[2:0],u_ca_out_531[11:3], u_ca_out_530[20:12], u_ca_out_529[23:21]};
assign col_out_533 = {u_ca_out_533[2:0],u_ca_out_532[11:3], u_ca_out_531[20:12], u_ca_out_530[23:21]};
assign col_out_534 = {u_ca_out_534[2:0],u_ca_out_533[11:3], u_ca_out_532[20:12], u_ca_out_531[23:21]};
assign col_out_535 = {u_ca_out_535[2:0],u_ca_out_534[11:3], u_ca_out_533[20:12], u_ca_out_532[23:21]};
assign col_out_536 = {u_ca_out_536[2:0],u_ca_out_535[11:3], u_ca_out_534[20:12], u_ca_out_533[23:21]};
assign col_out_537 = {u_ca_out_537[2:0],u_ca_out_536[11:3], u_ca_out_535[20:12], u_ca_out_534[23:21]};
assign col_out_538 = {u_ca_out_538[2:0],u_ca_out_537[11:3], u_ca_out_536[20:12], u_ca_out_535[23:21]};
assign col_out_539 = {u_ca_out_539[2:0],u_ca_out_538[11:3], u_ca_out_537[20:12], u_ca_out_536[23:21]};
assign col_out_540 = {u_ca_out_540[2:0],u_ca_out_539[11:3], u_ca_out_538[20:12], u_ca_out_537[23:21]};
assign col_out_541 = {u_ca_out_541[2:0],u_ca_out_540[11:3], u_ca_out_539[20:12], u_ca_out_538[23:21]};
assign col_out_542 = {u_ca_out_542[2:0],u_ca_out_541[11:3], u_ca_out_540[20:12], u_ca_out_539[23:21]};
assign col_out_543 = {u_ca_out_543[2:0],u_ca_out_542[11:3], u_ca_out_541[20:12], u_ca_out_540[23:21]};
assign col_out_544 = {u_ca_out_544[2:0],u_ca_out_543[11:3], u_ca_out_542[20:12], u_ca_out_541[23:21]};
assign col_out_545 = {u_ca_out_545[2:0],u_ca_out_544[11:3], u_ca_out_543[20:12], u_ca_out_542[23:21]};
assign col_out_546 = {u_ca_out_546[2:0],u_ca_out_545[11:3], u_ca_out_544[20:12], u_ca_out_543[23:21]};
assign col_out_547 = {u_ca_out_547[2:0],u_ca_out_546[11:3], u_ca_out_545[20:12], u_ca_out_544[23:21]};
assign col_out_548 = {u_ca_out_548[2:0],u_ca_out_547[11:3], u_ca_out_546[20:12], u_ca_out_545[23:21]};
assign col_out_549 = {u_ca_out_549[2:0],u_ca_out_548[11:3], u_ca_out_547[20:12], u_ca_out_546[23:21]};
assign col_out_550 = {u_ca_out_550[2:0],u_ca_out_549[11:3], u_ca_out_548[20:12], u_ca_out_547[23:21]};
assign col_out_551 = {u_ca_out_551[2:0],u_ca_out_550[11:3], u_ca_out_549[20:12], u_ca_out_548[23:21]};
assign col_out_552 = {u_ca_out_552[2:0],u_ca_out_551[11:3], u_ca_out_550[20:12], u_ca_out_549[23:21]};
assign col_out_553 = {u_ca_out_553[2:0],u_ca_out_552[11:3], u_ca_out_551[20:12], u_ca_out_550[23:21]};
assign col_out_554 = {u_ca_out_554[2:0],u_ca_out_553[11:3], u_ca_out_552[20:12], u_ca_out_551[23:21]};
assign col_out_555 = {u_ca_out_555[2:0],u_ca_out_554[11:3], u_ca_out_553[20:12], u_ca_out_552[23:21]};
assign col_out_556 = {u_ca_out_556[2:0],u_ca_out_555[11:3], u_ca_out_554[20:12], u_ca_out_553[23:21]};
assign col_out_557 = {u_ca_out_557[2:0],u_ca_out_556[11:3], u_ca_out_555[20:12], u_ca_out_554[23:21]};
assign col_out_558 = {u_ca_out_558[2:0],u_ca_out_557[11:3], u_ca_out_556[20:12], u_ca_out_555[23:21]};
assign col_out_559 = {u_ca_out_559[2:0],u_ca_out_558[11:3], u_ca_out_557[20:12], u_ca_out_556[23:21]};
assign col_out_560 = {u_ca_out_560[2:0],u_ca_out_559[11:3], u_ca_out_558[20:12], u_ca_out_557[23:21]};
assign col_out_561 = {u_ca_out_561[2:0],u_ca_out_560[11:3], u_ca_out_559[20:12], u_ca_out_558[23:21]};
assign col_out_562 = {u_ca_out_562[2:0],u_ca_out_561[11:3], u_ca_out_560[20:12], u_ca_out_559[23:21]};
assign col_out_563 = {u_ca_out_563[2:0],u_ca_out_562[11:3], u_ca_out_561[20:12], u_ca_out_560[23:21]};
assign col_out_564 = {u_ca_out_564[2:0],u_ca_out_563[11:3], u_ca_out_562[20:12], u_ca_out_561[23:21]};
assign col_out_565 = {u_ca_out_565[2:0],u_ca_out_564[11:3], u_ca_out_563[20:12], u_ca_out_562[23:21]};
assign col_out_566 = {u_ca_out_566[2:0],u_ca_out_565[11:3], u_ca_out_564[20:12], u_ca_out_563[23:21]};
assign col_out_567 = {u_ca_out_567[2:0],u_ca_out_566[11:3], u_ca_out_565[20:12], u_ca_out_564[23:21]};
assign col_out_568 = {u_ca_out_568[2:0],u_ca_out_567[11:3], u_ca_out_566[20:12], u_ca_out_565[23:21]};
assign col_out_569 = {u_ca_out_569[2:0],u_ca_out_568[11:3], u_ca_out_567[20:12], u_ca_out_566[23:21]};
assign col_out_570 = {u_ca_out_570[2:0],u_ca_out_569[11:3], u_ca_out_568[20:12], u_ca_out_567[23:21]};
assign col_out_571 = {u_ca_out_571[2:0],u_ca_out_570[11:3], u_ca_out_569[20:12], u_ca_out_568[23:21]};
assign col_out_572 = {u_ca_out_572[2:0],u_ca_out_571[11:3], u_ca_out_570[20:12], u_ca_out_569[23:21]};
assign col_out_573 = {u_ca_out_573[2:0],u_ca_out_572[11:3], u_ca_out_571[20:12], u_ca_out_570[23:21]};
assign col_out_574 = {u_ca_out_574[2:0],u_ca_out_573[11:3], u_ca_out_572[20:12], u_ca_out_571[23:21]};
assign col_out_575 = {u_ca_out_575[2:0],u_ca_out_574[11:3], u_ca_out_573[20:12], u_ca_out_572[23:21]};
assign col_out_576 = {u_ca_out_576[2:0],u_ca_out_575[11:3], u_ca_out_574[20:12], u_ca_out_573[23:21]};
assign col_out_577 = {u_ca_out_577[2:0],u_ca_out_576[11:3], u_ca_out_575[20:12], u_ca_out_574[23:21]};
assign col_out_578 = {u_ca_out_578[2:0],u_ca_out_577[11:3], u_ca_out_576[20:12], u_ca_out_575[23:21]};
assign col_out_579 = {u_ca_out_579[2:0],u_ca_out_578[11:3], u_ca_out_577[20:12], u_ca_out_576[23:21]};
assign col_out_580 = {u_ca_out_580[2:0],u_ca_out_579[11:3], u_ca_out_578[20:12], u_ca_out_577[23:21]};
assign col_out_581 = {u_ca_out_581[2:0],u_ca_out_580[11:3], u_ca_out_579[20:12], u_ca_out_578[23:21]};
assign col_out_582 = {u_ca_out_582[2:0],u_ca_out_581[11:3], u_ca_out_580[20:12], u_ca_out_579[23:21]};
assign col_out_583 = {u_ca_out_583[2:0],u_ca_out_582[11:3], u_ca_out_581[20:12], u_ca_out_580[23:21]};
assign col_out_584 = {u_ca_out_584[2:0],u_ca_out_583[11:3], u_ca_out_582[20:12], u_ca_out_581[23:21]};
assign col_out_585 = {u_ca_out_585[2:0],u_ca_out_584[11:3], u_ca_out_583[20:12], u_ca_out_582[23:21]};
assign col_out_586 = {u_ca_out_586[2:0],u_ca_out_585[11:3], u_ca_out_584[20:12], u_ca_out_583[23:21]};
assign col_out_587 = {u_ca_out_587[2:0],u_ca_out_586[11:3], u_ca_out_585[20:12], u_ca_out_584[23:21]};
assign col_out_588 = {u_ca_out_588[2:0],u_ca_out_587[11:3], u_ca_out_586[20:12], u_ca_out_585[23:21]};
assign col_out_589 = {u_ca_out_589[2:0],u_ca_out_588[11:3], u_ca_out_587[20:12], u_ca_out_586[23:21]};
assign col_out_590 = {u_ca_out_590[2:0],u_ca_out_589[11:3], u_ca_out_588[20:12], u_ca_out_587[23:21]};
assign col_out_591 = {u_ca_out_591[2:0],u_ca_out_590[11:3], u_ca_out_589[20:12], u_ca_out_588[23:21]};
assign col_out_592 = {u_ca_out_592[2:0],u_ca_out_591[11:3], u_ca_out_590[20:12], u_ca_out_589[23:21]};
assign col_out_593 = {u_ca_out_593[2:0],u_ca_out_592[11:3], u_ca_out_591[20:12], u_ca_out_590[23:21]};
assign col_out_594 = {u_ca_out_594[2:0],u_ca_out_593[11:3], u_ca_out_592[20:12], u_ca_out_591[23:21]};
assign col_out_595 = {u_ca_out_595[2:0],u_ca_out_594[11:3], u_ca_out_593[20:12], u_ca_out_592[23:21]};
assign col_out_596 = {u_ca_out_596[2:0],u_ca_out_595[11:3], u_ca_out_594[20:12], u_ca_out_593[23:21]};
assign col_out_597 = {u_ca_out_597[2:0],u_ca_out_596[11:3], u_ca_out_595[20:12], u_ca_out_594[23:21]};
assign col_out_598 = {u_ca_out_598[2:0],u_ca_out_597[11:3], u_ca_out_596[20:12], u_ca_out_595[23:21]};
assign col_out_599 = {u_ca_out_599[2:0],u_ca_out_598[11:3], u_ca_out_597[20:12], u_ca_out_596[23:21]};
assign col_out_600 = {u_ca_out_600[2:0],u_ca_out_599[11:3], u_ca_out_598[20:12], u_ca_out_597[23:21]};
assign col_out_601 = {u_ca_out_601[2:0],u_ca_out_600[11:3], u_ca_out_599[20:12], u_ca_out_598[23:21]};
assign col_out_602 = {u_ca_out_602[2:0],u_ca_out_601[11:3], u_ca_out_600[20:12], u_ca_out_599[23:21]};
assign col_out_603 = {u_ca_out_603[2:0],u_ca_out_602[11:3], u_ca_out_601[20:12], u_ca_out_600[23:21]};
assign col_out_604 = {u_ca_out_604[2:0],u_ca_out_603[11:3], u_ca_out_602[20:12], u_ca_out_601[23:21]};
assign col_out_605 = {u_ca_out_605[2:0],u_ca_out_604[11:3], u_ca_out_603[20:12], u_ca_out_602[23:21]};
assign col_out_606 = {u_ca_out_606[2:0],u_ca_out_605[11:3], u_ca_out_604[20:12], u_ca_out_603[23:21]};
assign col_out_607 = {u_ca_out_607[2:0],u_ca_out_606[11:3], u_ca_out_605[20:12], u_ca_out_604[23:21]};
assign col_out_608 = {u_ca_out_608[2:0],u_ca_out_607[11:3], u_ca_out_606[20:12], u_ca_out_605[23:21]};
assign col_out_609 = {u_ca_out_609[2:0],u_ca_out_608[11:3], u_ca_out_607[20:12], u_ca_out_606[23:21]};
assign col_out_610 = {u_ca_out_610[2:0],u_ca_out_609[11:3], u_ca_out_608[20:12], u_ca_out_607[23:21]};
assign col_out_611 = {u_ca_out_611[2:0],u_ca_out_610[11:3], u_ca_out_609[20:12], u_ca_out_608[23:21]};
assign col_out_612 = {u_ca_out_612[2:0],u_ca_out_611[11:3], u_ca_out_610[20:12], u_ca_out_609[23:21]};
assign col_out_613 = {u_ca_out_613[2:0],u_ca_out_612[11:3], u_ca_out_611[20:12], u_ca_out_610[23:21]};
assign col_out_614 = {u_ca_out_614[2:0],u_ca_out_613[11:3], u_ca_out_612[20:12], u_ca_out_611[23:21]};
assign col_out_615 = {u_ca_out_615[2:0],u_ca_out_614[11:3], u_ca_out_613[20:12], u_ca_out_612[23:21]};
assign col_out_616 = {u_ca_out_616[2:0],u_ca_out_615[11:3], u_ca_out_614[20:12], u_ca_out_613[23:21]};
assign col_out_617 = {u_ca_out_617[2:0],u_ca_out_616[11:3], u_ca_out_615[20:12], u_ca_out_614[23:21]};
assign col_out_618 = {u_ca_out_618[2:0],u_ca_out_617[11:3], u_ca_out_616[20:12], u_ca_out_615[23:21]};
assign col_out_619 = {u_ca_out_619[2:0],u_ca_out_618[11:3], u_ca_out_617[20:12], u_ca_out_616[23:21]};
assign col_out_620 = {u_ca_out_620[2:0],u_ca_out_619[11:3], u_ca_out_618[20:12], u_ca_out_617[23:21]};
assign col_out_621 = {u_ca_out_621[2:0],u_ca_out_620[11:3], u_ca_out_619[20:12], u_ca_out_618[23:21]};
assign col_out_622 = {u_ca_out_622[2:0],u_ca_out_621[11:3], u_ca_out_620[20:12], u_ca_out_619[23:21]};
assign col_out_623 = {u_ca_out_623[2:0],u_ca_out_622[11:3], u_ca_out_621[20:12], u_ca_out_620[23:21]};
assign col_out_624 = {u_ca_out_624[2:0],u_ca_out_623[11:3], u_ca_out_622[20:12], u_ca_out_621[23:21]};
assign col_out_625 = {u_ca_out_625[2:0],u_ca_out_624[11:3], u_ca_out_623[20:12], u_ca_out_622[23:21]};
assign col_out_626 = {u_ca_out_626[2:0],u_ca_out_625[11:3], u_ca_out_624[20:12], u_ca_out_623[23:21]};
assign col_out_627 = {u_ca_out_627[2:0],u_ca_out_626[11:3], u_ca_out_625[20:12], u_ca_out_624[23:21]};
assign col_out_628 = {u_ca_out_628[2:0],u_ca_out_627[11:3], u_ca_out_626[20:12], u_ca_out_625[23:21]};
assign col_out_629 = {u_ca_out_629[2:0],u_ca_out_628[11:3], u_ca_out_627[20:12], u_ca_out_626[23:21]};
assign col_out_630 = {u_ca_out_630[2:0],u_ca_out_629[11:3], u_ca_out_628[20:12], u_ca_out_627[23:21]};
assign col_out_631 = {u_ca_out_631[2:0],u_ca_out_630[11:3], u_ca_out_629[20:12], u_ca_out_628[23:21]};
assign col_out_632 = {u_ca_out_632[2:0],u_ca_out_631[11:3], u_ca_out_630[20:12], u_ca_out_629[23:21]};
assign col_out_633 = {u_ca_out_633[2:0],u_ca_out_632[11:3], u_ca_out_631[20:12], u_ca_out_630[23:21]};
assign col_out_634 = {u_ca_out_634[2:0],u_ca_out_633[11:3], u_ca_out_632[20:12], u_ca_out_631[23:21]};
assign col_out_635 = {u_ca_out_635[2:0],u_ca_out_634[11:3], u_ca_out_633[20:12], u_ca_out_632[23:21]};
assign col_out_636 = {u_ca_out_636[2:0],u_ca_out_635[11:3], u_ca_out_634[20:12], u_ca_out_633[23:21]};
assign col_out_637 = {u_ca_out_637[2:0],u_ca_out_636[11:3], u_ca_out_635[20:12], u_ca_out_634[23:21]};
assign col_out_638 = {u_ca_out_638[2:0],u_ca_out_637[11:3], u_ca_out_636[20:12], u_ca_out_635[23:21]};
assign col_out_639 = {u_ca_out_639[2:0],u_ca_out_638[11:3], u_ca_out_637[20:12], u_ca_out_636[23:21]};
assign col_out_640 = {u_ca_out_640[2:0],u_ca_out_639[11:3], u_ca_out_638[20:12], u_ca_out_637[23:21]};
assign col_out_641 = {u_ca_out_641[2:0],u_ca_out_640[11:3], u_ca_out_639[20:12], u_ca_out_638[23:21]};
assign col_out_642 = {u_ca_out_642[2:0],u_ca_out_641[11:3], u_ca_out_640[20:12], u_ca_out_639[23:21]};
assign col_out_643 = {u_ca_out_643[2:0],u_ca_out_642[11:3], u_ca_out_641[20:12], u_ca_out_640[23:21]};
assign col_out_644 = {u_ca_out_644[2:0],u_ca_out_643[11:3], u_ca_out_642[20:12], u_ca_out_641[23:21]};
assign col_out_645 = {u_ca_out_645[2:0],u_ca_out_644[11:3], u_ca_out_643[20:12], u_ca_out_642[23:21]};
assign col_out_646 = {u_ca_out_646[2:0],u_ca_out_645[11:3], u_ca_out_644[20:12], u_ca_out_643[23:21]};
assign col_out_647 = {u_ca_out_647[2:0],u_ca_out_646[11:3], u_ca_out_645[20:12], u_ca_out_644[23:21]};
assign col_out_648 = {u_ca_out_648[2:0],u_ca_out_647[11:3], u_ca_out_646[20:12], u_ca_out_645[23:21]};
assign col_out_649 = {u_ca_out_649[2:0],u_ca_out_648[11:3], u_ca_out_647[20:12], u_ca_out_646[23:21]};
assign col_out_650 = {u_ca_out_650[2:0],u_ca_out_649[11:3], u_ca_out_648[20:12], u_ca_out_647[23:21]};
assign col_out_651 = {u_ca_out_651[2:0],u_ca_out_650[11:3], u_ca_out_649[20:12], u_ca_out_648[23:21]};
assign col_out_652 = {u_ca_out_652[2:0],u_ca_out_651[11:3], u_ca_out_650[20:12], u_ca_out_649[23:21]};
assign col_out_653 = {u_ca_out_653[2:0],u_ca_out_652[11:3], u_ca_out_651[20:12], u_ca_out_650[23:21]};
assign col_out_654 = {u_ca_out_654[2:0],u_ca_out_653[11:3], u_ca_out_652[20:12], u_ca_out_651[23:21]};
assign col_out_655 = {u_ca_out_655[2:0],u_ca_out_654[11:3], u_ca_out_653[20:12], u_ca_out_652[23:21]};
assign col_out_656 = {u_ca_out_656[2:0],u_ca_out_655[11:3], u_ca_out_654[20:12], u_ca_out_653[23:21]};
assign col_out_657 = {u_ca_out_657[2:0],u_ca_out_656[11:3], u_ca_out_655[20:12], u_ca_out_654[23:21]};
assign col_out_658 = {u_ca_out_658[2:0],u_ca_out_657[11:3], u_ca_out_656[20:12], u_ca_out_655[23:21]};
assign col_out_659 = {u_ca_out_659[2:0],u_ca_out_658[11:3], u_ca_out_657[20:12], u_ca_out_656[23:21]};
assign col_out_660 = {u_ca_out_660[2:0],u_ca_out_659[11:3], u_ca_out_658[20:12], u_ca_out_657[23:21]};
assign col_out_661 = {u_ca_out_661[2:0],u_ca_out_660[11:3], u_ca_out_659[20:12], u_ca_out_658[23:21]};
assign col_out_662 = {u_ca_out_662[2:0],u_ca_out_661[11:3], u_ca_out_660[20:12], u_ca_out_659[23:21]};
assign col_out_663 = {u_ca_out_663[2:0],u_ca_out_662[11:3], u_ca_out_661[20:12], u_ca_out_660[23:21]};
assign col_out_664 = {u_ca_out_664[2:0],u_ca_out_663[11:3], u_ca_out_662[20:12], u_ca_out_661[23:21]};
assign col_out_665 = {u_ca_out_665[2:0],u_ca_out_664[11:3], u_ca_out_663[20:12], u_ca_out_662[23:21]};
assign col_out_666 = {u_ca_out_666[2:0],u_ca_out_665[11:3], u_ca_out_664[20:12], u_ca_out_663[23:21]};
assign col_out_667 = {u_ca_out_667[2:0],u_ca_out_666[11:3], u_ca_out_665[20:12], u_ca_out_664[23:21]};
assign col_out_668 = {u_ca_out_668[2:0],u_ca_out_667[11:3], u_ca_out_666[20:12], u_ca_out_665[23:21]};
assign col_out_669 = {u_ca_out_669[2:0],u_ca_out_668[11:3], u_ca_out_667[20:12], u_ca_out_666[23:21]};
assign col_out_670 = {u_ca_out_670[2:0],u_ca_out_669[11:3], u_ca_out_668[20:12], u_ca_out_667[23:21]};
assign col_out_671 = {u_ca_out_671[2:0],u_ca_out_670[11:3], u_ca_out_669[20:12], u_ca_out_668[23:21]};
assign col_out_672 = {u_ca_out_672[2:0],u_ca_out_671[11:3], u_ca_out_670[20:12], u_ca_out_669[23:21]};
assign col_out_673 = {u_ca_out_673[2:0],u_ca_out_672[11:3], u_ca_out_671[20:12], u_ca_out_670[23:21]};
assign col_out_674 = {u_ca_out_674[2:0],u_ca_out_673[11:3], u_ca_out_672[20:12], u_ca_out_671[23:21]};
assign col_out_675 = {u_ca_out_675[2:0],u_ca_out_674[11:3], u_ca_out_673[20:12], u_ca_out_672[23:21]};
assign col_out_676 = {u_ca_out_676[2:0],u_ca_out_675[11:3], u_ca_out_674[20:12], u_ca_out_673[23:21]};
assign col_out_677 = {u_ca_out_677[2:0],u_ca_out_676[11:3], u_ca_out_675[20:12], u_ca_out_674[23:21]};
assign col_out_678 = {u_ca_out_678[2:0],u_ca_out_677[11:3], u_ca_out_676[20:12], u_ca_out_675[23:21]};
assign col_out_679 = {u_ca_out_679[2:0],u_ca_out_678[11:3], u_ca_out_677[20:12], u_ca_out_676[23:21]};
assign col_out_680 = {u_ca_out_680[2:0],u_ca_out_679[11:3], u_ca_out_678[20:12], u_ca_out_677[23:21]};
assign col_out_681 = {u_ca_out_681[2:0],u_ca_out_680[11:3], u_ca_out_679[20:12], u_ca_out_678[23:21]};
assign col_out_682 = {u_ca_out_682[2:0],u_ca_out_681[11:3], u_ca_out_680[20:12], u_ca_out_679[23:21]};
assign col_out_683 = {u_ca_out_683[2:0],u_ca_out_682[11:3], u_ca_out_681[20:12], u_ca_out_680[23:21]};
assign col_out_684 = {u_ca_out_684[2:0],u_ca_out_683[11:3], u_ca_out_682[20:12], u_ca_out_681[23:21]};
assign col_out_685 = {u_ca_out_685[2:0],u_ca_out_684[11:3], u_ca_out_683[20:12], u_ca_out_682[23:21]};
assign col_out_686 = {u_ca_out_686[2:0],u_ca_out_685[11:3], u_ca_out_684[20:12], u_ca_out_683[23:21]};
assign col_out_687 = {u_ca_out_687[2:0],u_ca_out_686[11:3], u_ca_out_685[20:12], u_ca_out_684[23:21]};
assign col_out_688 = {u_ca_out_688[2:0],u_ca_out_687[11:3], u_ca_out_686[20:12], u_ca_out_685[23:21]};
assign col_out_689 = {u_ca_out_689[2:0],u_ca_out_688[11:3], u_ca_out_687[20:12], u_ca_out_686[23:21]};
assign col_out_690 = {u_ca_out_690[2:0],u_ca_out_689[11:3], u_ca_out_688[20:12], u_ca_out_687[23:21]};
assign col_out_691 = {u_ca_out_691[2:0],u_ca_out_690[11:3], u_ca_out_689[20:12], u_ca_out_688[23:21]};
assign col_out_692 = {u_ca_out_692[2:0],u_ca_out_691[11:3], u_ca_out_690[20:12], u_ca_out_689[23:21]};
assign col_out_693 = {u_ca_out_693[2:0],u_ca_out_692[11:3], u_ca_out_691[20:12], u_ca_out_690[23:21]};
assign col_out_694 = {u_ca_out_694[2:0],u_ca_out_693[11:3], u_ca_out_692[20:12], u_ca_out_691[23:21]};
assign col_out_695 = {u_ca_out_695[2:0],u_ca_out_694[11:3], u_ca_out_693[20:12], u_ca_out_692[23:21]};
assign col_out_696 = {u_ca_out_696[2:0],u_ca_out_695[11:3], u_ca_out_694[20:12], u_ca_out_693[23:21]};
assign col_out_697 = {u_ca_out_697[2:0],u_ca_out_696[11:3], u_ca_out_695[20:12], u_ca_out_694[23:21]};
assign col_out_698 = {u_ca_out_698[2:0],u_ca_out_697[11:3], u_ca_out_696[20:12], u_ca_out_695[23:21]};
assign col_out_699 = {u_ca_out_699[2:0],u_ca_out_698[11:3], u_ca_out_697[20:12], u_ca_out_696[23:21]};
assign col_out_700 = {u_ca_out_700[2:0],u_ca_out_699[11:3], u_ca_out_698[20:12], u_ca_out_697[23:21]};
assign col_out_701 = {u_ca_out_701[2:0],u_ca_out_700[11:3], u_ca_out_699[20:12], u_ca_out_698[23:21]};
assign col_out_702 = {u_ca_out_702[2:0],u_ca_out_701[11:3], u_ca_out_700[20:12], u_ca_out_699[23:21]};
assign col_out_703 = {u_ca_out_703[2:0],u_ca_out_702[11:3], u_ca_out_701[20:12], u_ca_out_700[23:21]};
assign col_out_704 = {u_ca_out_704[2:0],u_ca_out_703[11:3], u_ca_out_702[20:12], u_ca_out_701[23:21]};
assign col_out_705 = {u_ca_out_705[2:0],u_ca_out_704[11:3], u_ca_out_703[20:12], u_ca_out_702[23:21]};
assign col_out_706 = {u_ca_out_706[2:0],u_ca_out_705[11:3], u_ca_out_704[20:12], u_ca_out_703[23:21]};
assign col_out_707 = {u_ca_out_707[2:0],u_ca_out_706[11:3], u_ca_out_705[20:12], u_ca_out_704[23:21]};
assign col_out_708 = {u_ca_out_708[2:0],u_ca_out_707[11:3], u_ca_out_706[20:12], u_ca_out_705[23:21]};
assign col_out_709 = {u_ca_out_709[2:0],u_ca_out_708[11:3], u_ca_out_707[20:12], u_ca_out_706[23:21]};
assign col_out_710 = {u_ca_out_710[2:0],u_ca_out_709[11:3], u_ca_out_708[20:12], u_ca_out_707[23:21]};
assign col_out_711 = {u_ca_out_711[2:0],u_ca_out_710[11:3], u_ca_out_709[20:12], u_ca_out_708[23:21]};
assign col_out_712 = {u_ca_out_712[2:0],u_ca_out_711[11:3], u_ca_out_710[20:12], u_ca_out_709[23:21]};
assign col_out_713 = {u_ca_out_713[2:0],u_ca_out_712[11:3], u_ca_out_711[20:12], u_ca_out_710[23:21]};
assign col_out_714 = {u_ca_out_714[2:0],u_ca_out_713[11:3], u_ca_out_712[20:12], u_ca_out_711[23:21]};
assign col_out_715 = {u_ca_out_715[2:0],u_ca_out_714[11:3], u_ca_out_713[20:12], u_ca_out_712[23:21]};
assign col_out_716 = {u_ca_out_716[2:0],u_ca_out_715[11:3], u_ca_out_714[20:12], u_ca_out_713[23:21]};
assign col_out_717 = {u_ca_out_717[2:0],u_ca_out_716[11:3], u_ca_out_715[20:12], u_ca_out_714[23:21]};
assign col_out_718 = {u_ca_out_718[2:0],u_ca_out_717[11:3], u_ca_out_716[20:12], u_ca_out_715[23:21]};
assign col_out_719 = {u_ca_out_719[2:0],u_ca_out_718[11:3], u_ca_out_717[20:12], u_ca_out_716[23:21]};
assign col_out_720 = {u_ca_out_720[2:0],u_ca_out_719[11:3], u_ca_out_718[20:12], u_ca_out_717[23:21]};
assign col_out_721 = {u_ca_out_721[2:0],u_ca_out_720[11:3], u_ca_out_719[20:12], u_ca_out_718[23:21]};
assign col_out_722 = {u_ca_out_722[2:0],u_ca_out_721[11:3], u_ca_out_720[20:12], u_ca_out_719[23:21]};
assign col_out_723 = {u_ca_out_723[2:0],u_ca_out_722[11:3], u_ca_out_721[20:12], u_ca_out_720[23:21]};
assign col_out_724 = {u_ca_out_724[2:0],u_ca_out_723[11:3], u_ca_out_722[20:12], u_ca_out_721[23:21]};
assign col_out_725 = {u_ca_out_725[2:0],u_ca_out_724[11:3], u_ca_out_723[20:12], u_ca_out_722[23:21]};
assign col_out_726 = {u_ca_out_726[2:0],u_ca_out_725[11:3], u_ca_out_724[20:12], u_ca_out_723[23:21]};
assign col_out_727 = {u_ca_out_727[2:0],u_ca_out_726[11:3], u_ca_out_725[20:12], u_ca_out_724[23:21]};
assign col_out_728 = {u_ca_out_728[2:0],u_ca_out_727[11:3], u_ca_out_726[20:12], u_ca_out_725[23:21]};
assign col_out_729 = {u_ca_out_729[2:0],u_ca_out_728[11:3], u_ca_out_727[20:12], u_ca_out_726[23:21]};
assign col_out_730 = {u_ca_out_730[2:0],u_ca_out_729[11:3], u_ca_out_728[20:12], u_ca_out_727[23:21]};
assign col_out_731 = {u_ca_out_731[2:0],u_ca_out_730[11:3], u_ca_out_729[20:12], u_ca_out_728[23:21]};
assign col_out_732 = {u_ca_out_732[2:0],u_ca_out_731[11:3], u_ca_out_730[20:12], u_ca_out_729[23:21]};
assign col_out_733 = {u_ca_out_733[2:0],u_ca_out_732[11:3], u_ca_out_731[20:12], u_ca_out_730[23:21]};
assign col_out_734 = {u_ca_out_734[2:0],u_ca_out_733[11:3], u_ca_out_732[20:12], u_ca_out_731[23:21]};
assign col_out_735 = {u_ca_out_735[2:0],u_ca_out_734[11:3], u_ca_out_733[20:12], u_ca_out_732[23:21]};
assign col_out_736 = {u_ca_out_736[2:0],u_ca_out_735[11:3], u_ca_out_734[20:12], u_ca_out_733[23:21]};
assign col_out_737 = {u_ca_out_737[2:0],u_ca_out_736[11:3], u_ca_out_735[20:12], u_ca_out_734[23:21]};
assign col_out_738 = {u_ca_out_738[2:0],u_ca_out_737[11:3], u_ca_out_736[20:12], u_ca_out_735[23:21]};
assign col_out_739 = {u_ca_out_739[2:0],u_ca_out_738[11:3], u_ca_out_737[20:12], u_ca_out_736[23:21]};
assign col_out_740 = {u_ca_out_740[2:0],u_ca_out_739[11:3], u_ca_out_738[20:12], u_ca_out_737[23:21]};
assign col_out_741 = {u_ca_out_741[2:0],u_ca_out_740[11:3], u_ca_out_739[20:12], u_ca_out_738[23:21]};
assign col_out_742 = {u_ca_out_742[2:0],u_ca_out_741[11:3], u_ca_out_740[20:12], u_ca_out_739[23:21]};
assign col_out_743 = {u_ca_out_743[2:0],u_ca_out_742[11:3], u_ca_out_741[20:12], u_ca_out_740[23:21]};
assign col_out_744 = {u_ca_out_744[2:0],u_ca_out_743[11:3], u_ca_out_742[20:12], u_ca_out_741[23:21]};
assign col_out_745 = {u_ca_out_745[2:0],u_ca_out_744[11:3], u_ca_out_743[20:12], u_ca_out_742[23:21]};
assign col_out_746 = {u_ca_out_746[2:0],u_ca_out_745[11:3], u_ca_out_744[20:12], u_ca_out_743[23:21]};
assign col_out_747 = {u_ca_out_747[2:0],u_ca_out_746[11:3], u_ca_out_745[20:12], u_ca_out_744[23:21]};
assign col_out_748 = {u_ca_out_748[2:0],u_ca_out_747[11:3], u_ca_out_746[20:12], u_ca_out_745[23:21]};
assign col_out_749 = {u_ca_out_749[2:0],u_ca_out_748[11:3], u_ca_out_747[20:12], u_ca_out_746[23:21]};
assign col_out_750 = {u_ca_out_750[2:0],u_ca_out_749[11:3], u_ca_out_748[20:12], u_ca_out_747[23:21]};
assign col_out_751 = {u_ca_out_751[2:0],u_ca_out_750[11:3], u_ca_out_749[20:12], u_ca_out_748[23:21]};
assign col_out_752 = {u_ca_out_752[2:0],u_ca_out_751[11:3], u_ca_out_750[20:12], u_ca_out_749[23:21]};
assign col_out_753 = {u_ca_out_753[2:0],u_ca_out_752[11:3], u_ca_out_751[20:12], u_ca_out_750[23:21]};
assign col_out_754 = {u_ca_out_754[2:0],u_ca_out_753[11:3], u_ca_out_752[20:12], u_ca_out_751[23:21]};
assign col_out_755 = {u_ca_out_755[2:0],u_ca_out_754[11:3], u_ca_out_753[20:12], u_ca_out_752[23:21]};
assign col_out_756 = {u_ca_out_756[2:0],u_ca_out_755[11:3], u_ca_out_754[20:12], u_ca_out_753[23:21]};
assign col_out_757 = {u_ca_out_757[2:0],u_ca_out_756[11:3], u_ca_out_755[20:12], u_ca_out_754[23:21]};
assign col_out_758 = {u_ca_out_758[2:0],u_ca_out_757[11:3], u_ca_out_756[20:12], u_ca_out_755[23:21]};
assign col_out_759 = {u_ca_out_759[2:0],u_ca_out_758[11:3], u_ca_out_757[20:12], u_ca_out_756[23:21]};
assign col_out_760 = {u_ca_out_760[2:0],u_ca_out_759[11:3], u_ca_out_758[20:12], u_ca_out_757[23:21]};
assign col_out_761 = {u_ca_out_761[2:0],u_ca_out_760[11:3], u_ca_out_759[20:12], u_ca_out_758[23:21]};
assign col_out_762 = {u_ca_out_762[2:0],u_ca_out_761[11:3], u_ca_out_760[20:12], u_ca_out_759[23:21]};
assign col_out_763 = {u_ca_out_763[2:0],u_ca_out_762[11:3], u_ca_out_761[20:12], u_ca_out_760[23:21]};
assign col_out_764 = {u_ca_out_764[2:0],u_ca_out_763[11:3], u_ca_out_762[20:12], u_ca_out_761[23:21]};
assign col_out_765 = {u_ca_out_765[2:0],u_ca_out_764[11:3], u_ca_out_763[20:12], u_ca_out_762[23:21]};
assign col_out_766 = {u_ca_out_766[2:0],u_ca_out_765[11:3], u_ca_out_764[20:12], u_ca_out_763[23:21]};
assign col_out_767 = {u_ca_out_767[2:0],u_ca_out_766[11:3], u_ca_out_765[20:12], u_ca_out_764[23:21]};
assign col_out_768 = {u_ca_out_768[2:0],u_ca_out_767[11:3], u_ca_out_766[20:12], u_ca_out_765[23:21]};
assign col_out_769 = {u_ca_out_769[2:0],u_ca_out_768[11:3], u_ca_out_767[20:12], u_ca_out_766[23:21]};
assign col_out_770 = {u_ca_out_770[2:0],u_ca_out_769[11:3], u_ca_out_768[20:12], u_ca_out_767[23:21]};
assign col_out_771 = {u_ca_out_771[2:0],u_ca_out_770[11:3], u_ca_out_769[20:12], u_ca_out_768[23:21]};
assign col_out_772 = {u_ca_out_772[2:0],u_ca_out_771[11:3], u_ca_out_770[20:12], u_ca_out_769[23:21]};
assign col_out_773 = {u_ca_out_773[2:0],u_ca_out_772[11:3], u_ca_out_771[20:12], u_ca_out_770[23:21]};
assign col_out_774 = {u_ca_out_774[2:0],u_ca_out_773[11:3], u_ca_out_772[20:12], u_ca_out_771[23:21]};
assign col_out_775 = {u_ca_out_775[2:0],u_ca_out_774[11:3], u_ca_out_773[20:12], u_ca_out_772[23:21]};
assign col_out_776 = {u_ca_out_776[2:0],u_ca_out_775[11:3], u_ca_out_774[20:12], u_ca_out_773[23:21]};
assign col_out_777 = {u_ca_out_777[2:0],u_ca_out_776[11:3], u_ca_out_775[20:12], u_ca_out_774[23:21]};
assign col_out_778 = {u_ca_out_778[2:0],u_ca_out_777[11:3], u_ca_out_776[20:12], u_ca_out_775[23:21]};
assign col_out_779 = {u_ca_out_779[2:0],u_ca_out_778[11:3], u_ca_out_777[20:12], u_ca_out_776[23:21]};
assign col_out_780 = {u_ca_out_780[2:0],u_ca_out_779[11:3], u_ca_out_778[20:12], u_ca_out_777[23:21]};
assign col_out_781 = {u_ca_out_781[2:0],u_ca_out_780[11:3], u_ca_out_779[20:12], u_ca_out_778[23:21]};
assign col_out_782 = {u_ca_out_782[2:0],u_ca_out_781[11:3], u_ca_out_780[20:12], u_ca_out_779[23:21]};
assign col_out_783 = {u_ca_out_783[2:0],u_ca_out_782[11:3], u_ca_out_781[20:12], u_ca_out_780[23:21]};
assign col_out_784 = {u_ca_out_784[2:0],u_ca_out_783[11:3], u_ca_out_782[20:12], u_ca_out_781[23:21]};
assign col_out_785 = {u_ca_out_785[2:0],u_ca_out_784[11:3], u_ca_out_783[20:12], u_ca_out_782[23:21]};
assign col_out_786 = {u_ca_out_786[2:0],u_ca_out_785[11:3], u_ca_out_784[20:12], u_ca_out_783[23:21]};
assign col_out_787 = {u_ca_out_787[2:0],u_ca_out_786[11:3], u_ca_out_785[20:12], u_ca_out_784[23:21]};
assign col_out_788 = {u_ca_out_788[2:0],u_ca_out_787[11:3], u_ca_out_786[20:12], u_ca_out_785[23:21]};
assign col_out_789 = {u_ca_out_789[2:0],u_ca_out_788[11:3], u_ca_out_787[20:12], u_ca_out_786[23:21]};
assign col_out_790 = {u_ca_out_790[2:0],u_ca_out_789[11:3], u_ca_out_788[20:12], u_ca_out_787[23:21]};
assign col_out_791 = {u_ca_out_791[2:0],u_ca_out_790[11:3], u_ca_out_789[20:12], u_ca_out_788[23:21]};
assign col_out_792 = {u_ca_out_792[2:0],u_ca_out_791[11:3], u_ca_out_790[20:12], u_ca_out_789[23:21]};
assign col_out_793 = {u_ca_out_793[2:0],u_ca_out_792[11:3], u_ca_out_791[20:12], u_ca_out_790[23:21]};
assign col_out_794 = {u_ca_out_794[2:0],u_ca_out_793[11:3], u_ca_out_792[20:12], u_ca_out_791[23:21]};
assign col_out_795 = {u_ca_out_795[2:0],u_ca_out_794[11:3], u_ca_out_793[20:12], u_ca_out_792[23:21]};
assign col_out_796 = {u_ca_out_796[2:0],u_ca_out_795[11:3], u_ca_out_794[20:12], u_ca_out_793[23:21]};
assign col_out_797 = {u_ca_out_797[2:0],u_ca_out_796[11:3], u_ca_out_795[20:12], u_ca_out_794[23:21]};
assign col_out_798 = {u_ca_out_798[2:0],u_ca_out_797[11:3], u_ca_out_796[20:12], u_ca_out_795[23:21]};
assign col_out_799 = {u_ca_out_799[2:0],u_ca_out_798[11:3], u_ca_out_797[20:12], u_ca_out_796[23:21]};
assign col_out_800 = {u_ca_out_800[2:0],u_ca_out_799[11:3], u_ca_out_798[20:12], u_ca_out_797[23:21]};
assign col_out_801 = {u_ca_out_801[2:0],u_ca_out_800[11:3], u_ca_out_799[20:12], u_ca_out_798[23:21]};
assign col_out_802 = {u_ca_out_802[2:0],u_ca_out_801[11:3], u_ca_out_800[20:12], u_ca_out_799[23:21]};
assign col_out_803 = {u_ca_out_803[2:0],u_ca_out_802[11:3], u_ca_out_801[20:12], u_ca_out_800[23:21]};
assign col_out_804 = {u_ca_out_804[2:0],u_ca_out_803[11:3], u_ca_out_802[20:12], u_ca_out_801[23:21]};
assign col_out_805 = {u_ca_out_805[2:0],u_ca_out_804[11:3], u_ca_out_803[20:12], u_ca_out_802[23:21]};
assign col_out_806 = {u_ca_out_806[2:0],u_ca_out_805[11:3], u_ca_out_804[20:12], u_ca_out_803[23:21]};
assign col_out_807 = {u_ca_out_807[2:0],u_ca_out_806[11:3], u_ca_out_805[20:12], u_ca_out_804[23:21]};
assign col_out_808 = {u_ca_out_808[2:0],u_ca_out_807[11:3], u_ca_out_806[20:12], u_ca_out_805[23:21]};
assign col_out_809 = {u_ca_out_809[2:0],u_ca_out_808[11:3], u_ca_out_807[20:12], u_ca_out_806[23:21]};
assign col_out_810 = {u_ca_out_810[2:0],u_ca_out_809[11:3], u_ca_out_808[20:12], u_ca_out_807[23:21]};
assign col_out_811 = {u_ca_out_811[2:0],u_ca_out_810[11:3], u_ca_out_809[20:12], u_ca_out_808[23:21]};
assign col_out_812 = {u_ca_out_812[2:0],u_ca_out_811[11:3], u_ca_out_810[20:12], u_ca_out_809[23:21]};
assign col_out_813 = {u_ca_out_813[2:0],u_ca_out_812[11:3], u_ca_out_811[20:12], u_ca_out_810[23:21]};
assign col_out_814 = {u_ca_out_814[2:0],u_ca_out_813[11:3], u_ca_out_812[20:12], u_ca_out_811[23:21]};
assign col_out_815 = {u_ca_out_815[2:0],u_ca_out_814[11:3], u_ca_out_813[20:12], u_ca_out_812[23:21]};
assign col_out_816 = {u_ca_out_816[2:0],u_ca_out_815[11:3], u_ca_out_814[20:12], u_ca_out_813[23:21]};
assign col_out_817 = {u_ca_out_817[2:0],u_ca_out_816[11:3], u_ca_out_815[20:12], u_ca_out_814[23:21]};
assign col_out_818 = {u_ca_out_818[2:0],u_ca_out_817[11:3], u_ca_out_816[20:12], u_ca_out_815[23:21]};
assign col_out_819 = {u_ca_out_819[2:0],u_ca_out_818[11:3], u_ca_out_817[20:12], u_ca_out_816[23:21]};
assign col_out_820 = {u_ca_out_820[2:0],u_ca_out_819[11:3], u_ca_out_818[20:12], u_ca_out_817[23:21]};
assign col_out_821 = {u_ca_out_821[2:0],u_ca_out_820[11:3], u_ca_out_819[20:12], u_ca_out_818[23:21]};
assign col_out_822 = {u_ca_out_822[2:0],u_ca_out_821[11:3], u_ca_out_820[20:12], u_ca_out_819[23:21]};
assign col_out_823 = {u_ca_out_823[2:0],u_ca_out_822[11:3], u_ca_out_821[20:12], u_ca_out_820[23:21]};
assign col_out_824 = {u_ca_out_824[2:0],u_ca_out_823[11:3], u_ca_out_822[20:12], u_ca_out_821[23:21]};
assign col_out_825 = {u_ca_out_825[2:0],u_ca_out_824[11:3], u_ca_out_823[20:12], u_ca_out_822[23:21]};
assign col_out_826 = {u_ca_out_826[2:0],u_ca_out_825[11:3], u_ca_out_824[20:12], u_ca_out_823[23:21]};
assign col_out_827 = {u_ca_out_827[2:0],u_ca_out_826[11:3], u_ca_out_825[20:12], u_ca_out_824[23:21]};
assign col_out_828 = {u_ca_out_828[2:0],u_ca_out_827[11:3], u_ca_out_826[20:12], u_ca_out_825[23:21]};
assign col_out_829 = {u_ca_out_829[2:0],u_ca_out_828[11:3], u_ca_out_827[20:12], u_ca_out_826[23:21]};
assign col_out_830 = {u_ca_out_830[2:0],u_ca_out_829[11:3], u_ca_out_828[20:12], u_ca_out_827[23:21]};
assign col_out_831 = {u_ca_out_831[2:0],u_ca_out_830[11:3], u_ca_out_829[20:12], u_ca_out_828[23:21]};
assign col_out_832 = {u_ca_out_832[2:0],u_ca_out_831[11:3], u_ca_out_830[20:12], u_ca_out_829[23:21]};
assign col_out_833 = {u_ca_out_833[2:0],u_ca_out_832[11:3], u_ca_out_831[20:12], u_ca_out_830[23:21]};
assign col_out_834 = {u_ca_out_834[2:0],u_ca_out_833[11:3], u_ca_out_832[20:12], u_ca_out_831[23:21]};
assign col_out_835 = {u_ca_out_835[2:0],u_ca_out_834[11:3], u_ca_out_833[20:12], u_ca_out_832[23:21]};
assign col_out_836 = {u_ca_out_836[2:0],u_ca_out_835[11:3], u_ca_out_834[20:12], u_ca_out_833[23:21]};
assign col_out_837 = {u_ca_out_837[2:0],u_ca_out_836[11:3], u_ca_out_835[20:12], u_ca_out_834[23:21]};
assign col_out_838 = {u_ca_out_838[2:0],u_ca_out_837[11:3], u_ca_out_836[20:12], u_ca_out_835[23:21]};
assign col_out_839 = {u_ca_out_839[2:0],u_ca_out_838[11:3], u_ca_out_837[20:12], u_ca_out_836[23:21]};
assign col_out_840 = {u_ca_out_840[2:0],u_ca_out_839[11:3], u_ca_out_838[20:12], u_ca_out_837[23:21]};
assign col_out_841 = {u_ca_out_841[2:0],u_ca_out_840[11:3], u_ca_out_839[20:12], u_ca_out_838[23:21]};
assign col_out_842 = {u_ca_out_842[2:0],u_ca_out_841[11:3], u_ca_out_840[20:12], u_ca_out_839[23:21]};
assign col_out_843 = {u_ca_out_843[2:0],u_ca_out_842[11:3], u_ca_out_841[20:12], u_ca_out_840[23:21]};
assign col_out_844 = {u_ca_out_844[2:0],u_ca_out_843[11:3], u_ca_out_842[20:12], u_ca_out_841[23:21]};
assign col_out_845 = {u_ca_out_845[2:0],u_ca_out_844[11:3], u_ca_out_843[20:12], u_ca_out_842[23:21]};
assign col_out_846 = {u_ca_out_846[2:0],u_ca_out_845[11:3], u_ca_out_844[20:12], u_ca_out_843[23:21]};
assign col_out_847 = {u_ca_out_847[2:0],u_ca_out_846[11:3], u_ca_out_845[20:12], u_ca_out_844[23:21]};
assign col_out_848 = {u_ca_out_848[2:0],u_ca_out_847[11:3], u_ca_out_846[20:12], u_ca_out_845[23:21]};
assign col_out_849 = {u_ca_out_849[2:0],u_ca_out_848[11:3], u_ca_out_847[20:12], u_ca_out_846[23:21]};
assign col_out_850 = {u_ca_out_850[2:0],u_ca_out_849[11:3], u_ca_out_848[20:12], u_ca_out_847[23:21]};
assign col_out_851 = {u_ca_out_851[2:0],u_ca_out_850[11:3], u_ca_out_849[20:12], u_ca_out_848[23:21]};
assign col_out_852 = {u_ca_out_852[2:0],u_ca_out_851[11:3], u_ca_out_850[20:12], u_ca_out_849[23:21]};
assign col_out_853 = {u_ca_out_853[2:0],u_ca_out_852[11:3], u_ca_out_851[20:12], u_ca_out_850[23:21]};
assign col_out_854 = {u_ca_out_854[2:0],u_ca_out_853[11:3], u_ca_out_852[20:12], u_ca_out_851[23:21]};
assign col_out_855 = {u_ca_out_855[2:0],u_ca_out_854[11:3], u_ca_out_853[20:12], u_ca_out_852[23:21]};
assign col_out_856 = {u_ca_out_856[2:0],u_ca_out_855[11:3], u_ca_out_854[20:12], u_ca_out_853[23:21]};
assign col_out_857 = {u_ca_out_857[2:0],u_ca_out_856[11:3], u_ca_out_855[20:12], u_ca_out_854[23:21]};
assign col_out_858 = {u_ca_out_858[2:0],u_ca_out_857[11:3], u_ca_out_856[20:12], u_ca_out_855[23:21]};
assign col_out_859 = {u_ca_out_859[2:0],u_ca_out_858[11:3], u_ca_out_857[20:12], u_ca_out_856[23:21]};
assign col_out_860 = {u_ca_out_860[2:0],u_ca_out_859[11:3], u_ca_out_858[20:12], u_ca_out_857[23:21]};
assign col_out_861 = {u_ca_out_861[2:0],u_ca_out_860[11:3], u_ca_out_859[20:12], u_ca_out_858[23:21]};
assign col_out_862 = {u_ca_out_862[2:0],u_ca_out_861[11:3], u_ca_out_860[20:12], u_ca_out_859[23:21]};
assign col_out_863 = {u_ca_out_863[2:0],u_ca_out_862[11:3], u_ca_out_861[20:12], u_ca_out_860[23:21]};
assign col_out_864 = {u_ca_out_864[2:0],u_ca_out_863[11:3], u_ca_out_862[20:12], u_ca_out_861[23:21]};
assign col_out_865 = {u_ca_out_865[2:0],u_ca_out_864[11:3], u_ca_out_863[20:12], u_ca_out_862[23:21]};
assign col_out_866 = {u_ca_out_866[2:0],u_ca_out_865[11:3], u_ca_out_864[20:12], u_ca_out_863[23:21]};
assign col_out_867 = {u_ca_out_867[2:0],u_ca_out_866[11:3], u_ca_out_865[20:12], u_ca_out_864[23:21]};
assign col_out_868 = {u_ca_out_868[2:0],u_ca_out_867[11:3], u_ca_out_866[20:12], u_ca_out_865[23:21]};
assign col_out_869 = {u_ca_out_869[2:0],u_ca_out_868[11:3], u_ca_out_867[20:12], u_ca_out_866[23:21]};
assign col_out_870 = {u_ca_out_870[2:0],u_ca_out_869[11:3], u_ca_out_868[20:12], u_ca_out_867[23:21]};
assign col_out_871 = {u_ca_out_871[2:0],u_ca_out_870[11:3], u_ca_out_869[20:12], u_ca_out_868[23:21]};
assign col_out_872 = {u_ca_out_872[2:0],u_ca_out_871[11:3], u_ca_out_870[20:12], u_ca_out_869[23:21]};
assign col_out_873 = {u_ca_out_873[2:0],u_ca_out_872[11:3], u_ca_out_871[20:12], u_ca_out_870[23:21]};
assign col_out_874 = {u_ca_out_874[2:0],u_ca_out_873[11:3], u_ca_out_872[20:12], u_ca_out_871[23:21]};
assign col_out_875 = {u_ca_out_875[2:0],u_ca_out_874[11:3], u_ca_out_873[20:12], u_ca_out_872[23:21]};
assign col_out_876 = {u_ca_out_876[2:0],u_ca_out_875[11:3], u_ca_out_874[20:12], u_ca_out_873[23:21]};
assign col_out_877 = {u_ca_out_877[2:0],u_ca_out_876[11:3], u_ca_out_875[20:12], u_ca_out_874[23:21]};
assign col_out_878 = {u_ca_out_878[2:0],u_ca_out_877[11:3], u_ca_out_876[20:12], u_ca_out_875[23:21]};
assign col_out_879 = {u_ca_out_879[2:0],u_ca_out_878[11:3], u_ca_out_877[20:12], u_ca_out_876[23:21]};
assign col_out_880 = {u_ca_out_880[2:0],u_ca_out_879[11:3], u_ca_out_878[20:12], u_ca_out_877[23:21]};
assign col_out_881 = {u_ca_out_881[2:0],u_ca_out_880[11:3], u_ca_out_879[20:12], u_ca_out_878[23:21]};
assign col_out_882 = {u_ca_out_882[2:0],u_ca_out_881[11:3], u_ca_out_880[20:12], u_ca_out_879[23:21]};
assign col_out_883 = {u_ca_out_883[2:0],u_ca_out_882[11:3], u_ca_out_881[20:12], u_ca_out_880[23:21]};
assign col_out_884 = {u_ca_out_884[2:0],u_ca_out_883[11:3], u_ca_out_882[20:12], u_ca_out_881[23:21]};
assign col_out_885 = {u_ca_out_885[2:0],u_ca_out_884[11:3], u_ca_out_883[20:12], u_ca_out_882[23:21]};
assign col_out_886 = {u_ca_out_886[2:0],u_ca_out_885[11:3], u_ca_out_884[20:12], u_ca_out_883[23:21]};
assign col_out_887 = {u_ca_out_887[2:0],u_ca_out_886[11:3], u_ca_out_885[20:12], u_ca_out_884[23:21]};
assign col_out_888 = {u_ca_out_888[2:0],u_ca_out_887[11:3], u_ca_out_886[20:12], u_ca_out_885[23:21]};
assign col_out_889 = {u_ca_out_889[2:0],u_ca_out_888[11:3], u_ca_out_887[20:12], u_ca_out_886[23:21]};
assign col_out_890 = {u_ca_out_890[2:0],u_ca_out_889[11:3], u_ca_out_888[20:12], u_ca_out_887[23:21]};
assign col_out_891 = {u_ca_out_891[2:0],u_ca_out_890[11:3], u_ca_out_889[20:12], u_ca_out_888[23:21]};
assign col_out_892 = {u_ca_out_892[2:0],u_ca_out_891[11:3], u_ca_out_890[20:12], u_ca_out_889[23:21]};
assign col_out_893 = {u_ca_out_893[2:0],u_ca_out_892[11:3], u_ca_out_891[20:12], u_ca_out_890[23:21]};
assign col_out_894 = {u_ca_out_894[2:0],u_ca_out_893[11:3], u_ca_out_892[20:12], u_ca_out_891[23:21]};
assign col_out_895 = {u_ca_out_895[2:0],u_ca_out_894[11:3], u_ca_out_893[20:12], u_ca_out_892[23:21]};
assign col_out_896 = {u_ca_out_896[2:0],u_ca_out_895[11:3], u_ca_out_894[20:12], u_ca_out_893[23:21]};
assign col_out_897 = {u_ca_out_897[2:0],u_ca_out_896[11:3], u_ca_out_895[20:12], u_ca_out_894[23:21]};
assign col_out_898 = {u_ca_out_898[2:0],u_ca_out_897[11:3], u_ca_out_896[20:12], u_ca_out_895[23:21]};
assign col_out_899 = {u_ca_out_899[2:0],u_ca_out_898[11:3], u_ca_out_897[20:12], u_ca_out_896[23:21]};
assign col_out_900 = {u_ca_out_900[2:0],u_ca_out_899[11:3], u_ca_out_898[20:12], u_ca_out_897[23:21]};
assign col_out_901 = {u_ca_out_901[2:0],u_ca_out_900[11:3], u_ca_out_899[20:12], u_ca_out_898[23:21]};
assign col_out_902 = {u_ca_out_902[2:0],u_ca_out_901[11:3], u_ca_out_900[20:12], u_ca_out_899[23:21]};
assign col_out_903 = {u_ca_out_903[2:0],u_ca_out_902[11:3], u_ca_out_901[20:12], u_ca_out_900[23:21]};
assign col_out_904 = {u_ca_out_904[2:0],u_ca_out_903[11:3], u_ca_out_902[20:12], u_ca_out_901[23:21]};
assign col_out_905 = {u_ca_out_905[2:0],u_ca_out_904[11:3], u_ca_out_903[20:12], u_ca_out_902[23:21]};
assign col_out_906 = {u_ca_out_906[2:0],u_ca_out_905[11:3], u_ca_out_904[20:12], u_ca_out_903[23:21]};
assign col_out_907 = {u_ca_out_907[2:0],u_ca_out_906[11:3], u_ca_out_905[20:12], u_ca_out_904[23:21]};
assign col_out_908 = {u_ca_out_908[2:0],u_ca_out_907[11:3], u_ca_out_906[20:12], u_ca_out_905[23:21]};
assign col_out_909 = {u_ca_out_909[2:0],u_ca_out_908[11:3], u_ca_out_907[20:12], u_ca_out_906[23:21]};
assign col_out_910 = {u_ca_out_910[2:0],u_ca_out_909[11:3], u_ca_out_908[20:12], u_ca_out_907[23:21]};
assign col_out_911 = {u_ca_out_911[2:0],u_ca_out_910[11:3], u_ca_out_909[20:12], u_ca_out_908[23:21]};
assign col_out_912 = {u_ca_out_912[2:0],u_ca_out_911[11:3], u_ca_out_910[20:12], u_ca_out_909[23:21]};
assign col_out_913 = {u_ca_out_913[2:0],u_ca_out_912[11:3], u_ca_out_911[20:12], u_ca_out_910[23:21]};
assign col_out_914 = {u_ca_out_914[2:0],u_ca_out_913[11:3], u_ca_out_912[20:12], u_ca_out_911[23:21]};
assign col_out_915 = {u_ca_out_915[2:0],u_ca_out_914[11:3], u_ca_out_913[20:12], u_ca_out_912[23:21]};
assign col_out_916 = {u_ca_out_916[2:0],u_ca_out_915[11:3], u_ca_out_914[20:12], u_ca_out_913[23:21]};
assign col_out_917 = {u_ca_out_917[2:0],u_ca_out_916[11:3], u_ca_out_915[20:12], u_ca_out_914[23:21]};
assign col_out_918 = {u_ca_out_918[2:0],u_ca_out_917[11:3], u_ca_out_916[20:12], u_ca_out_915[23:21]};
assign col_out_919 = {u_ca_out_919[2:0],u_ca_out_918[11:3], u_ca_out_917[20:12], u_ca_out_916[23:21]};
assign col_out_920 = {u_ca_out_920[2:0],u_ca_out_919[11:3], u_ca_out_918[20:12], u_ca_out_917[23:21]};
assign col_out_921 = {u_ca_out_921[2:0],u_ca_out_920[11:3], u_ca_out_919[20:12], u_ca_out_918[23:21]};
assign col_out_922 = {u_ca_out_922[2:0],u_ca_out_921[11:3], u_ca_out_920[20:12], u_ca_out_919[23:21]};
assign col_out_923 = {u_ca_out_923[2:0],u_ca_out_922[11:3], u_ca_out_921[20:12], u_ca_out_920[23:21]};
assign col_out_924 = {u_ca_out_924[2:0],u_ca_out_923[11:3], u_ca_out_922[20:12], u_ca_out_921[23:21]};
assign col_out_925 = {u_ca_out_925[2:0],u_ca_out_924[11:3], u_ca_out_923[20:12], u_ca_out_922[23:21]};
assign col_out_926 = {u_ca_out_926[2:0],u_ca_out_925[11:3], u_ca_out_924[20:12], u_ca_out_923[23:21]};
assign col_out_927 = {u_ca_out_927[2:0],u_ca_out_926[11:3], u_ca_out_925[20:12], u_ca_out_924[23:21]};
assign col_out_928 = {u_ca_out_928[2:0],u_ca_out_927[11:3], u_ca_out_926[20:12], u_ca_out_925[23:21]};
assign col_out_929 = {u_ca_out_929[2:0],u_ca_out_928[11:3], u_ca_out_927[20:12], u_ca_out_926[23:21]};
assign col_out_930 = {u_ca_out_930[2:0],u_ca_out_929[11:3], u_ca_out_928[20:12], u_ca_out_927[23:21]};
assign col_out_931 = {u_ca_out_931[2:0],u_ca_out_930[11:3], u_ca_out_929[20:12], u_ca_out_928[23:21]};
assign col_out_932 = {u_ca_out_932[2:0],u_ca_out_931[11:3], u_ca_out_930[20:12], u_ca_out_929[23:21]};
assign col_out_933 = {u_ca_out_933[2:0],u_ca_out_932[11:3], u_ca_out_931[20:12], u_ca_out_930[23:21]};
assign col_out_934 = {u_ca_out_934[2:0],u_ca_out_933[11:3], u_ca_out_932[20:12], u_ca_out_931[23:21]};
assign col_out_935 = {u_ca_out_935[2:0],u_ca_out_934[11:3], u_ca_out_933[20:12], u_ca_out_932[23:21]};
assign col_out_936 = {u_ca_out_936[2:0],u_ca_out_935[11:3], u_ca_out_934[20:12], u_ca_out_933[23:21]};
assign col_out_937 = {u_ca_out_937[2:0],u_ca_out_936[11:3], u_ca_out_935[20:12], u_ca_out_934[23:21]};
assign col_out_938 = {u_ca_out_938[2:0],u_ca_out_937[11:3], u_ca_out_936[20:12], u_ca_out_935[23:21]};
assign col_out_939 = {u_ca_out_939[2:0],u_ca_out_938[11:3], u_ca_out_937[20:12], u_ca_out_936[23:21]};
assign col_out_940 = {u_ca_out_940[2:0],u_ca_out_939[11:3], u_ca_out_938[20:12], u_ca_out_937[23:21]};
assign col_out_941 = {u_ca_out_941[2:0],u_ca_out_940[11:3], u_ca_out_939[20:12], u_ca_out_938[23:21]};
assign col_out_942 = {u_ca_out_942[2:0],u_ca_out_941[11:3], u_ca_out_940[20:12], u_ca_out_939[23:21]};
assign col_out_943 = {u_ca_out_943[2:0],u_ca_out_942[11:3], u_ca_out_941[20:12], u_ca_out_940[23:21]};
assign col_out_944 = {u_ca_out_944[2:0],u_ca_out_943[11:3], u_ca_out_942[20:12], u_ca_out_941[23:21]};
assign col_out_945 = {u_ca_out_945[2:0],u_ca_out_944[11:3], u_ca_out_943[20:12], u_ca_out_942[23:21]};
assign col_out_946 = {u_ca_out_946[2:0],u_ca_out_945[11:3], u_ca_out_944[20:12], u_ca_out_943[23:21]};
assign col_out_947 = {u_ca_out_947[2:0],u_ca_out_946[11:3], u_ca_out_945[20:12], u_ca_out_944[23:21]};
assign col_out_948 = {u_ca_out_948[2:0],u_ca_out_947[11:3], u_ca_out_946[20:12], u_ca_out_945[23:21]};
assign col_out_949 = {u_ca_out_949[2:0],u_ca_out_948[11:3], u_ca_out_947[20:12], u_ca_out_946[23:21]};
assign col_out_950 = {u_ca_out_950[2:0],u_ca_out_949[11:3], u_ca_out_948[20:12], u_ca_out_947[23:21]};
assign col_out_951 = {u_ca_out_951[2:0],u_ca_out_950[11:3], u_ca_out_949[20:12], u_ca_out_948[23:21]};
assign col_out_952 = {u_ca_out_952[2:0],u_ca_out_951[11:3], u_ca_out_950[20:12], u_ca_out_949[23:21]};
assign col_out_953 = {u_ca_out_953[2:0],u_ca_out_952[11:3], u_ca_out_951[20:12], u_ca_out_950[23:21]};
assign col_out_954 = {u_ca_out_954[2:0],u_ca_out_953[11:3], u_ca_out_952[20:12], u_ca_out_951[23:21]};
assign col_out_955 = {u_ca_out_955[2:0],u_ca_out_954[11:3], u_ca_out_953[20:12], u_ca_out_952[23:21]};
assign col_out_956 = {u_ca_out_956[2:0],u_ca_out_955[11:3], u_ca_out_954[20:12], u_ca_out_953[23:21]};
assign col_out_957 = {u_ca_out_957[2:0],u_ca_out_956[11:3], u_ca_out_955[20:12], u_ca_out_954[23:21]};
assign col_out_958 = {u_ca_out_958[2:0],u_ca_out_957[11:3], u_ca_out_956[20:12], u_ca_out_955[23:21]};
assign col_out_959 = {u_ca_out_959[2:0],u_ca_out_958[11:3], u_ca_out_957[20:12], u_ca_out_956[23:21]};
assign col_out_960 = {u_ca_out_960[2:0],u_ca_out_959[11:3], u_ca_out_958[20:12], u_ca_out_957[23:21]};
assign col_out_961 = {u_ca_out_961[2:0],u_ca_out_960[11:3], u_ca_out_959[20:12], u_ca_out_958[23:21]};
assign col_out_962 = {u_ca_out_962[2:0],u_ca_out_961[11:3], u_ca_out_960[20:12], u_ca_out_959[23:21]};
assign col_out_963 = {u_ca_out_963[2:0],u_ca_out_962[11:3], u_ca_out_961[20:12], u_ca_out_960[23:21]};
assign col_out_964 = {u_ca_out_964[2:0],u_ca_out_963[11:3], u_ca_out_962[20:12], u_ca_out_961[23:21]};
assign col_out_965 = {u_ca_out_965[2:0],u_ca_out_964[11:3], u_ca_out_963[20:12], u_ca_out_962[23:21]};
assign col_out_966 = {u_ca_out_966[2:0],u_ca_out_965[11:3], u_ca_out_964[20:12], u_ca_out_963[23:21]};
assign col_out_967 = {u_ca_out_967[2:0],u_ca_out_966[11:3], u_ca_out_965[20:12], u_ca_out_964[23:21]};
assign col_out_968 = {u_ca_out_968[2:0],u_ca_out_967[11:3], u_ca_out_966[20:12], u_ca_out_965[23:21]};
assign col_out_969 = {u_ca_out_969[2:0],u_ca_out_968[11:3], u_ca_out_967[20:12], u_ca_out_966[23:21]};
assign col_out_970 = {u_ca_out_970[2:0],u_ca_out_969[11:3], u_ca_out_968[20:12], u_ca_out_967[23:21]};
assign col_out_971 = {u_ca_out_971[2:0],u_ca_out_970[11:3], u_ca_out_969[20:12], u_ca_out_968[23:21]};
assign col_out_972 = {u_ca_out_972[2:0],u_ca_out_971[11:3], u_ca_out_970[20:12], u_ca_out_969[23:21]};
assign col_out_973 = {u_ca_out_973[2:0],u_ca_out_972[11:3], u_ca_out_971[20:12], u_ca_out_970[23:21]};
assign col_out_974 = {u_ca_out_974[2:0],u_ca_out_973[11:3], u_ca_out_972[20:12], u_ca_out_971[23:21]};
assign col_out_975 = {u_ca_out_975[2:0],u_ca_out_974[11:3], u_ca_out_973[20:12], u_ca_out_972[23:21]};
assign col_out_976 = {u_ca_out_976[2:0],u_ca_out_975[11:3], u_ca_out_974[20:12], u_ca_out_973[23:21]};
assign col_out_977 = {u_ca_out_977[2:0],u_ca_out_976[11:3], u_ca_out_975[20:12], u_ca_out_974[23:21]};
assign col_out_978 = {u_ca_out_978[2:0],u_ca_out_977[11:3], u_ca_out_976[20:12], u_ca_out_975[23:21]};
assign col_out_979 = {u_ca_out_979[2:0],u_ca_out_978[11:3], u_ca_out_977[20:12], u_ca_out_976[23:21]};
assign col_out_980 = {u_ca_out_980[2:0],u_ca_out_979[11:3], u_ca_out_978[20:12], u_ca_out_977[23:21]};
assign col_out_981 = {u_ca_out_981[2:0],u_ca_out_980[11:3], u_ca_out_979[20:12], u_ca_out_978[23:21]};
assign col_out_982 = {u_ca_out_982[2:0],u_ca_out_981[11:3], u_ca_out_980[20:12], u_ca_out_979[23:21]};
assign col_out_983 = {u_ca_out_983[2:0],u_ca_out_982[11:3], u_ca_out_981[20:12], u_ca_out_980[23:21]};
assign col_out_984 = {u_ca_out_984[2:0],u_ca_out_983[11:3], u_ca_out_982[20:12], u_ca_out_981[23:21]};
assign col_out_985 = {u_ca_out_985[2:0],u_ca_out_984[11:3], u_ca_out_983[20:12], u_ca_out_982[23:21]};
assign col_out_986 = {u_ca_out_986[2:0],u_ca_out_985[11:3], u_ca_out_984[20:12], u_ca_out_983[23:21]};
assign col_out_987 = {u_ca_out_987[2:0],u_ca_out_986[11:3], u_ca_out_985[20:12], u_ca_out_984[23:21]};
assign col_out_988 = {u_ca_out_988[2:0],u_ca_out_987[11:3], u_ca_out_986[20:12], u_ca_out_985[23:21]};
assign col_out_989 = {u_ca_out_989[2:0],u_ca_out_988[11:3], u_ca_out_987[20:12], u_ca_out_986[23:21]};
assign col_out_990 = {u_ca_out_990[2:0],u_ca_out_989[11:3], u_ca_out_988[20:12], u_ca_out_987[23:21]};
assign col_out_991 = {u_ca_out_991[2:0],u_ca_out_990[11:3], u_ca_out_989[20:12], u_ca_out_988[23:21]};
assign col_out_992 = {u_ca_out_992[2:0],u_ca_out_991[11:3], u_ca_out_990[20:12], u_ca_out_989[23:21]};
assign col_out_993 = {u_ca_out_993[2:0],u_ca_out_992[11:3], u_ca_out_991[20:12], u_ca_out_990[23:21]};
assign col_out_994 = {u_ca_out_994[2:0],u_ca_out_993[11:3], u_ca_out_992[20:12], u_ca_out_991[23:21]};
assign col_out_995 = {u_ca_out_995[2:0],u_ca_out_994[11:3], u_ca_out_993[20:12], u_ca_out_992[23:21]};
assign col_out_996 = {u_ca_out_996[2:0],u_ca_out_995[11:3], u_ca_out_994[20:12], u_ca_out_993[23:21]};
assign col_out_997 = {u_ca_out_997[2:0],u_ca_out_996[11:3], u_ca_out_995[20:12], u_ca_out_994[23:21]};
assign col_out_998 = {u_ca_out_998[2:0],u_ca_out_997[11:3], u_ca_out_996[20:12], u_ca_out_995[23:21]};
assign col_out_999 = {u_ca_out_999[2:0],u_ca_out_998[11:3], u_ca_out_997[20:12], u_ca_out_996[23:21]};
assign col_out_1000 = {u_ca_out_1000[2:0],u_ca_out_999[11:3], u_ca_out_998[20:12], u_ca_out_997[23:21]};
assign col_out_1001 = {u_ca_out_1001[2:0],u_ca_out_1000[11:3], u_ca_out_999[20:12], u_ca_out_998[23:21]};
assign col_out_1002 = {u_ca_out_1002[2:0],u_ca_out_1001[11:3], u_ca_out_1000[20:12], u_ca_out_999[23:21]};
assign col_out_1003 = {u_ca_out_1003[2:0],u_ca_out_1002[11:3], u_ca_out_1001[20:12], u_ca_out_1000[23:21]};
assign col_out_1004 = {u_ca_out_1004[2:0],u_ca_out_1003[11:3], u_ca_out_1002[20:12], u_ca_out_1001[23:21]};
assign col_out_1005 = {u_ca_out_1005[2:0],u_ca_out_1004[11:3], u_ca_out_1003[20:12], u_ca_out_1002[23:21]};
assign col_out_1006 = {u_ca_out_1006[2:0],u_ca_out_1005[11:3], u_ca_out_1004[20:12], u_ca_out_1003[23:21]};
assign col_out_1007 = {u_ca_out_1007[2:0],u_ca_out_1006[11:3], u_ca_out_1005[20:12], u_ca_out_1004[23:21]};
assign col_out_1008 = {u_ca_out_1008[2:0],u_ca_out_1007[11:3], u_ca_out_1006[20:12], u_ca_out_1005[23:21]};
assign col_out_1009 = {u_ca_out_1009[2:0],u_ca_out_1008[11:3], u_ca_out_1007[20:12], u_ca_out_1006[23:21]};
assign col_out_1010 = {u_ca_out_1010[2:0],u_ca_out_1009[11:3], u_ca_out_1008[20:12], u_ca_out_1007[23:21]};
assign col_out_1011 = {u_ca_out_1011[2:0],u_ca_out_1010[11:3], u_ca_out_1009[20:12], u_ca_out_1008[23:21]};
assign col_out_1012 = {u_ca_out_1012[2:0],u_ca_out_1011[11:3], u_ca_out_1010[20:12], u_ca_out_1009[23:21]};
assign col_out_1013 = {u_ca_out_1013[2:0],u_ca_out_1012[11:3], u_ca_out_1011[20:12], u_ca_out_1010[23:21]};
assign col_out_1014 = {u_ca_out_1014[2:0],u_ca_out_1013[11:3], u_ca_out_1012[20:12], u_ca_out_1011[23:21]};
assign col_out_1015 = {u_ca_out_1015[2:0],u_ca_out_1014[11:3], u_ca_out_1013[20:12], u_ca_out_1012[23:21]};
assign col_out_1016 = {u_ca_out_1016[2:0],u_ca_out_1015[11:3], u_ca_out_1014[20:12], u_ca_out_1013[23:21]};
assign col_out_1017 = {u_ca_out_1017[2:0],u_ca_out_1016[11:3], u_ca_out_1015[20:12], u_ca_out_1014[23:21]};
assign col_out_1018 = {u_ca_out_1018[2:0],u_ca_out_1017[11:3], u_ca_out_1016[20:12], u_ca_out_1015[23:21]};
assign col_out_1019 = {u_ca_out_1019[2:0],u_ca_out_1018[11:3], u_ca_out_1017[20:12], u_ca_out_1016[23:21]};
assign col_out_1020 = {u_ca_out_1020[2:0],u_ca_out_1019[11:3], u_ca_out_1018[20:12], u_ca_out_1017[23:21]};
assign col_out_1021 = {u_ca_out_1021[2:0],u_ca_out_1020[11:3], u_ca_out_1019[20:12], u_ca_out_1018[23:21]};
assign col_out_1022 = {u_ca_out_1022[2:0],u_ca_out_1021[11:3], u_ca_out_1020[20:12], u_ca_out_1019[23:21]};
assign col_out_1023 = {u_ca_out_1023[2:0],u_ca_out_1022[11:3], u_ca_out_1021[20:12], u_ca_out_1020[23:21]};
assign col_out_1024 = {u_ca_out_1024[2:0],u_ca_out_1023[11:3], u_ca_out_1022[20:12], u_ca_out_1021[23:21]};
assign col_out_1025 = {u_ca_out_1025[2:0],u_ca_out_1024[11:3], u_ca_out_1023[20:12], u_ca_out_1022[23:21]};
assign col_out_1026 = {u_ca_out_1026[2:0],u_ca_out_1025[11:3], u_ca_out_1024[20:12], u_ca_out_1023[23:21]};
assign col_out_1027 = {u_ca_out_1027[2:0],u_ca_out_1026[11:3], u_ca_out_1025[20:12], u_ca_out_1024[23:21]};
assign col_out_1028 = {u_ca_out_1028[2:0],u_ca_out_1027[11:3], u_ca_out_1026[20:12], u_ca_out_1025[23:21]};
assign col_out_1029 = {u_ca_out_1029[2:0],u_ca_out_1028[11:3], u_ca_out_1027[20:12], u_ca_out_1026[23:21]};
assign col_out_1030 = {u_ca_out_1030[2:0],u_ca_out_1029[11:3], u_ca_out_1028[20:12], u_ca_out_1027[23:21]};
assign col_out_1031 = {u_ca_out_1031[2:0],u_ca_out_1030[11:3], u_ca_out_1029[20:12], u_ca_out_1028[23:21]};
assign col_out_1032 = {u_ca_out_1032[2:0],u_ca_out_1031[11:3], u_ca_out_1030[20:12], u_ca_out_1029[23:21]};
assign col_out_1033 = {u_ca_out_1033[2:0],u_ca_out_1032[11:3], u_ca_out_1031[20:12], u_ca_out_1030[23:21]};
assign col_out_1034 = {u_ca_out_1034[2:0],u_ca_out_1033[11:3], u_ca_out_1032[20:12], u_ca_out_1031[23:21]};
assign col_out_1035 = {u_ca_out_1035[2:0],u_ca_out_1034[11:3], u_ca_out_1033[20:12], u_ca_out_1032[23:21]};
assign col_out_1036 = {u_ca_out_1036[2:0],u_ca_out_1035[11:3], u_ca_out_1034[20:12], u_ca_out_1033[23:21]};
assign col_out_1037 = {u_ca_out_1037[2:0],u_ca_out_1036[11:3], u_ca_out_1035[20:12], u_ca_out_1034[23:21]};
assign col_out_1038 = {u_ca_out_1038[2:0],u_ca_out_1037[11:3], u_ca_out_1036[20:12], u_ca_out_1035[23:21]};
assign col_out_1039 = {u_ca_out_1039[2:0],u_ca_out_1038[11:3], u_ca_out_1037[20:12], u_ca_out_1036[23:21]};
assign col_out_1040 = {u_ca_out_1040[2:0],u_ca_out_1039[11:3], u_ca_out_1038[20:12], u_ca_out_1037[23:21]};
assign col_out_1041 = {u_ca_out_1041[2:0],u_ca_out_1040[11:3], u_ca_out_1039[20:12], u_ca_out_1038[23:21]};
assign col_out_1042 = {u_ca_out_1042[2:0],u_ca_out_1041[11:3], u_ca_out_1040[20:12], u_ca_out_1039[23:21]};
assign col_out_1043 = {u_ca_out_1043[2:0],u_ca_out_1042[11:3], u_ca_out_1041[20:12], u_ca_out_1040[23:21]};
assign col_out_1044 = {u_ca_out_1044[2:0],u_ca_out_1043[11:3], u_ca_out_1042[20:12], u_ca_out_1041[23:21]};
assign col_out_1045 = {u_ca_out_1045[2:0],u_ca_out_1044[11:3], u_ca_out_1043[20:12], u_ca_out_1042[23:21]};
assign col_out_1046 = {u_ca_out_1046[2:0],u_ca_out_1045[11:3], u_ca_out_1044[20:12], u_ca_out_1043[23:21]};
assign col_out_1047 = {u_ca_out_1047[2:0],u_ca_out_1046[11:3], u_ca_out_1045[20:12], u_ca_out_1044[23:21]};
assign col_out_1048 = {u_ca_out_1048[2:0],u_ca_out_1047[11:3], u_ca_out_1046[20:12], u_ca_out_1045[23:21]};
assign col_out_1049 = {u_ca_out_1049[2:0],u_ca_out_1048[11:3], u_ca_out_1047[20:12], u_ca_out_1046[23:21]};
assign col_out_1050 = {u_ca_out_1050[2:0],u_ca_out_1049[11:3], u_ca_out_1048[20:12], u_ca_out_1047[23:21]};
assign col_out_1051 = {u_ca_out_1051[2:0],u_ca_out_1050[11:3], u_ca_out_1049[20:12], u_ca_out_1048[23:21]};
assign col_out_1052 = {u_ca_out_1052[2:0],u_ca_out_1051[11:3], u_ca_out_1050[20:12], u_ca_out_1049[23:21]};
assign col_out_1053 = {u_ca_out_1053[2:0],u_ca_out_1052[11:3], u_ca_out_1051[20:12], u_ca_out_1050[23:21]};
assign col_out_1054 = {u_ca_out_1054[2:0],u_ca_out_1053[11:3], u_ca_out_1052[20:12], u_ca_out_1051[23:21]};
assign col_out_1055 = {u_ca_out_1055[2:0],u_ca_out_1054[11:3], u_ca_out_1053[20:12], u_ca_out_1052[23:21]};
assign col_out_1056 = {u_ca_out_1056[2:0],u_ca_out_1055[11:3], u_ca_out_1054[20:12], u_ca_out_1053[23:21]};
assign col_out_1057 = {u_ca_out_1057[2:0],u_ca_out_1056[11:3], u_ca_out_1055[20:12], u_ca_out_1054[23:21]};
assign col_out_1058 = {u_ca_out_1058[2:0],u_ca_out_1057[11:3], u_ca_out_1056[20:12], u_ca_out_1055[23:21]};
assign col_out_1059 = {u_ca_out_1059[2:0],u_ca_out_1058[11:3], u_ca_out_1057[20:12], u_ca_out_1056[23:21]};
assign col_out_1060 = {u_ca_out_1060[2:0],u_ca_out_1059[11:3], u_ca_out_1058[20:12], u_ca_out_1057[23:21]};
assign col_out_1061 = {u_ca_out_1061[2:0],u_ca_out_1060[11:3], u_ca_out_1059[20:12], u_ca_out_1058[23:21]};
assign col_out_1062 = {u_ca_out_1062[2:0],u_ca_out_1061[11:3], u_ca_out_1060[20:12], u_ca_out_1059[23:21]};
assign col_out_1063 = {u_ca_out_1063[2:0],u_ca_out_1062[11:3], u_ca_out_1061[20:12], u_ca_out_1060[23:21]};
assign col_out_1064 = {u_ca_out_1064[2:0],u_ca_out_1063[11:3], u_ca_out_1062[20:12], u_ca_out_1061[23:21]};
assign col_out_1065 = {u_ca_out_1065[2:0],u_ca_out_1064[11:3], u_ca_out_1063[20:12], u_ca_out_1062[23:21]};
assign col_out_1066 = {u_ca_out_1066[2:0],u_ca_out_1065[11:3], u_ca_out_1064[20:12], u_ca_out_1063[23:21]};
assign col_out_1067 = {u_ca_out_1067[2:0],u_ca_out_1066[11:3], u_ca_out_1065[20:12], u_ca_out_1064[23:21]};
assign col_out_1068 = {u_ca_out_1068[2:0],u_ca_out_1067[11:3], u_ca_out_1066[20:12], u_ca_out_1065[23:21]};
assign col_out_1069 = {u_ca_out_1069[2:0],u_ca_out_1068[11:3], u_ca_out_1067[20:12], u_ca_out_1066[23:21]};
assign col_out_1070 = {u_ca_out_1070[2:0],u_ca_out_1069[11:3], u_ca_out_1068[20:12], u_ca_out_1067[23:21]};
assign col_out_1071 = {u_ca_out_1071[2:0],u_ca_out_1070[11:3], u_ca_out_1069[20:12], u_ca_out_1068[23:21]};
assign col_out_1072 = {u_ca_out_1072[2:0],u_ca_out_1071[11:3], u_ca_out_1070[20:12], u_ca_out_1069[23:21]};
assign col_out_1073 = {u_ca_out_1073[2:0],u_ca_out_1072[11:3], u_ca_out_1071[20:12], u_ca_out_1070[23:21]};
assign col_out_1074 = {u_ca_out_1074[2:0],u_ca_out_1073[11:3], u_ca_out_1072[20:12], u_ca_out_1071[23:21]};
assign col_out_1075 = {u_ca_out_1075[2:0],u_ca_out_1074[11:3], u_ca_out_1073[20:12], u_ca_out_1072[23:21]};
assign col_out_1076 = {u_ca_out_1076[2:0],u_ca_out_1075[11:3], u_ca_out_1074[20:12], u_ca_out_1073[23:21]};
assign col_out_1077 = {u_ca_out_1077[2:0],u_ca_out_1076[11:3], u_ca_out_1075[20:12], u_ca_out_1074[23:21]};
assign col_out_1078 = {u_ca_out_1078[2:0],u_ca_out_1077[11:3], u_ca_out_1076[20:12], u_ca_out_1075[23:21]};
assign col_out_1079 = {u_ca_out_1079[2:0],u_ca_out_1078[11:3], u_ca_out_1077[20:12], u_ca_out_1076[23:21]};
assign col_out_1080 = {u_ca_out_1080[2:0],u_ca_out_1079[11:3], u_ca_out_1078[20:12], u_ca_out_1077[23:21]};
assign col_out_1081 = {u_ca_out_1081[2:0],u_ca_out_1080[11:3], u_ca_out_1079[20:12], u_ca_out_1078[23:21]};
assign col_out_1082 = {u_ca_out_1082[2:0],u_ca_out_1081[11:3], u_ca_out_1080[20:12], u_ca_out_1079[23:21]};
assign col_out_1083 = {u_ca_out_1083[2:0],u_ca_out_1082[11:3], u_ca_out_1081[20:12], u_ca_out_1080[23:21]};
assign col_out_1084 = {u_ca_out_1084[2:0],u_ca_out_1083[11:3], u_ca_out_1082[20:12], u_ca_out_1081[23:21]};
assign col_out_1085 = {u_ca_out_1085[2:0],u_ca_out_1084[11:3], u_ca_out_1083[20:12], u_ca_out_1082[23:21]};
assign col_out_1086 = {u_ca_out_1086[2:0],u_ca_out_1085[11:3], u_ca_out_1084[20:12], u_ca_out_1083[23:21]};
assign col_out_1087 = {u_ca_out_1087[2:0],u_ca_out_1086[11:3], u_ca_out_1085[20:12], u_ca_out_1084[23:21]};
assign col_out_1088 = {u_ca_out_1088[2:0],u_ca_out_1087[11:3], u_ca_out_1086[20:12], u_ca_out_1085[23:21]};
assign col_out_1089 = {u_ca_out_1089[2:0],u_ca_out_1088[11:3], u_ca_out_1087[20:12], u_ca_out_1086[23:21]};
assign col_out_1090 = {u_ca_out_1090[2:0],u_ca_out_1089[11:3], u_ca_out_1088[20:12], u_ca_out_1087[23:21]};
assign col_out_1091 = {u_ca_out_1091[2:0],u_ca_out_1090[11:3], u_ca_out_1089[20:12], u_ca_out_1088[23:21]};
assign col_out_1092 = {u_ca_out_1092[2:0],u_ca_out_1091[11:3], u_ca_out_1090[20:12], u_ca_out_1089[23:21]};
assign col_out_1093 = {u_ca_out_1093[2:0],u_ca_out_1092[11:3], u_ca_out_1091[20:12], u_ca_out_1090[23:21]};
assign col_out_1094 = {u_ca_out_1094[2:0],u_ca_out_1093[11:3], u_ca_out_1092[20:12], u_ca_out_1091[23:21]};
assign col_out_1095 = {u_ca_out_1095[2:0],u_ca_out_1094[11:3], u_ca_out_1093[20:12], u_ca_out_1092[23:21]};
assign col_out_1096 = {u_ca_out_1096[2:0],u_ca_out_1095[11:3], u_ca_out_1094[20:12], u_ca_out_1093[23:21]};
assign col_out_1097 = {u_ca_out_1097[2:0],u_ca_out_1096[11:3], u_ca_out_1095[20:12], u_ca_out_1094[23:21]};
assign col_out_1098 = {u_ca_out_1098[2:0],u_ca_out_1097[11:3], u_ca_out_1096[20:12], u_ca_out_1095[23:21]};
assign col_out_1099 = {u_ca_out_1099[2:0],u_ca_out_1098[11:3], u_ca_out_1097[20:12], u_ca_out_1096[23:21]};
assign col_out_1100 = {u_ca_out_1100[2:0],u_ca_out_1099[11:3], u_ca_out_1098[20:12], u_ca_out_1097[23:21]};
assign col_out_1101 = {u_ca_out_1101[2:0],u_ca_out_1100[11:3], u_ca_out_1099[20:12], u_ca_out_1098[23:21]};
assign col_out_1102 = {u_ca_out_1102[2:0],u_ca_out_1101[11:3], u_ca_out_1100[20:12], u_ca_out_1099[23:21]};
assign col_out_1103 = {u_ca_out_1103[2:0],u_ca_out_1102[11:3], u_ca_out_1101[20:12], u_ca_out_1100[23:21]};
assign col_out_1104 = {u_ca_out_1104[2:0],u_ca_out_1103[11:3], u_ca_out_1102[20:12], u_ca_out_1101[23:21]};
assign col_out_1105 = {u_ca_out_1105[2:0],u_ca_out_1104[11:3], u_ca_out_1103[20:12], u_ca_out_1102[23:21]};
assign col_out_1106 = {u_ca_out_1106[2:0],u_ca_out_1105[11:3], u_ca_out_1104[20:12], u_ca_out_1103[23:21]};
assign col_out_1107 = {u_ca_out_1107[2:0],u_ca_out_1106[11:3], u_ca_out_1105[20:12], u_ca_out_1104[23:21]};
assign col_out_1108 = {u_ca_out_1108[2:0],u_ca_out_1107[11:3], u_ca_out_1106[20:12], u_ca_out_1105[23:21]};
assign col_out_1109 = {u_ca_out_1109[2:0],u_ca_out_1108[11:3], u_ca_out_1107[20:12], u_ca_out_1106[23:21]};
assign col_out_1110 = {u_ca_out_1110[2:0],u_ca_out_1109[11:3], u_ca_out_1108[20:12], u_ca_out_1107[23:21]};
assign col_out_1111 = {u_ca_out_1111[2:0],u_ca_out_1110[11:3], u_ca_out_1109[20:12], u_ca_out_1108[23:21]};
assign col_out_1112 = {u_ca_out_1112[2:0],u_ca_out_1111[11:3], u_ca_out_1110[20:12], u_ca_out_1109[23:21]};
assign col_out_1113 = {u_ca_out_1113[2:0],u_ca_out_1112[11:3], u_ca_out_1111[20:12], u_ca_out_1110[23:21]};
assign col_out_1114 = {u_ca_out_1114[2:0],u_ca_out_1113[11:3], u_ca_out_1112[20:12], u_ca_out_1111[23:21]};
assign col_out_1115 = {u_ca_out_1115[2:0],u_ca_out_1114[11:3], u_ca_out_1113[20:12], u_ca_out_1112[23:21]};
assign col_out_1116 = {u_ca_out_1116[2:0],u_ca_out_1115[11:3], u_ca_out_1114[20:12], u_ca_out_1113[23:21]};
assign col_out_1117 = {u_ca_out_1117[2:0],u_ca_out_1116[11:3], u_ca_out_1115[20:12], u_ca_out_1114[23:21]};
assign col_out_1118 = {u_ca_out_1118[2:0],u_ca_out_1117[11:3], u_ca_out_1116[20:12], u_ca_out_1115[23:21]};
assign col_out_1119 = {u_ca_out_1119[2:0],u_ca_out_1118[11:3], u_ca_out_1117[20:12], u_ca_out_1116[23:21]};
assign col_out_1120 = {u_ca_out_1120[2:0],u_ca_out_1119[11:3], u_ca_out_1118[20:12], u_ca_out_1117[23:21]};
assign col_out_1121 = {u_ca_out_1121[2:0],u_ca_out_1120[11:3], u_ca_out_1119[20:12], u_ca_out_1118[23:21]};
assign col_out_1122 = {u_ca_out_1122[2:0],u_ca_out_1121[11:3], u_ca_out_1120[20:12], u_ca_out_1119[23:21]};
assign col_out_1123 = {u_ca_out_1123[2:0],u_ca_out_1122[11:3], u_ca_out_1121[20:12], u_ca_out_1120[23:21]};
assign col_out_1124 = {u_ca_out_1124[2:0],u_ca_out_1123[11:3], u_ca_out_1122[20:12], u_ca_out_1121[23:21]};
assign col_out_1125 = {u_ca_out_1125[2:0],u_ca_out_1124[11:3], u_ca_out_1123[20:12], u_ca_out_1122[23:21]};
assign col_out_1126 = {u_ca_out_1126[2:0],u_ca_out_1125[11:3], u_ca_out_1124[20:12], u_ca_out_1123[23:21]};
assign col_out_1127 = {u_ca_out_1127[2:0],u_ca_out_1126[11:3], u_ca_out_1125[20:12], u_ca_out_1124[23:21]};
assign col_out_1128 = {u_ca_out_1128[2:0],u_ca_out_1127[11:3], u_ca_out_1126[20:12], u_ca_out_1125[23:21]};
assign col_out_1129 = {u_ca_out_1129[2:0],u_ca_out_1128[11:3], u_ca_out_1127[20:12], u_ca_out_1126[23:21]};
assign col_out_1130 = {u_ca_out_1130[2:0],u_ca_out_1129[11:3], u_ca_out_1128[20:12], u_ca_out_1127[23:21]};
assign col_out_1131 = {u_ca_out_1131[2:0],u_ca_out_1130[11:3], u_ca_out_1129[20:12], u_ca_out_1128[23:21]};
assign col_out_1132 = {u_ca_out_1132[2:0],u_ca_out_1131[11:3], u_ca_out_1130[20:12], u_ca_out_1129[23:21]};
assign col_out_1133 = {u_ca_out_1133[2:0],u_ca_out_1132[11:3], u_ca_out_1131[20:12], u_ca_out_1130[23:21]};
assign col_out_1134 = {u_ca_out_1134[2:0],u_ca_out_1133[11:3], u_ca_out_1132[20:12], u_ca_out_1131[23:21]};
assign col_out_1135 = {u_ca_out_1135[2:0],u_ca_out_1134[11:3], u_ca_out_1133[20:12], u_ca_out_1132[23:21]};
assign col_out_1136 = {u_ca_out_1136[2:0],u_ca_out_1135[11:3], u_ca_out_1134[20:12], u_ca_out_1133[23:21]};
assign col_out_1137 = {u_ca_out_1137[2:0],u_ca_out_1136[11:3], u_ca_out_1135[20:12], u_ca_out_1134[23:21]};
assign col_out_1138 = {u_ca_out_1138[2:0],u_ca_out_1137[11:3], u_ca_out_1136[20:12], u_ca_out_1135[23:21]};
assign col_out_1139 = {u_ca_out_1139[2:0],u_ca_out_1138[11:3], u_ca_out_1137[20:12], u_ca_out_1136[23:21]};
assign col_out_1140 = {u_ca_out_1140[2:0],u_ca_out_1139[11:3], u_ca_out_1138[20:12], u_ca_out_1137[23:21]};
assign col_out_1141 = {u_ca_out_1141[2:0],u_ca_out_1140[11:3], u_ca_out_1139[20:12], u_ca_out_1138[23:21]};
assign col_out_1142 = {u_ca_out_1142[2:0],u_ca_out_1141[11:3], u_ca_out_1140[20:12], u_ca_out_1139[23:21]};
assign col_out_1143 = {u_ca_out_1143[2:0],u_ca_out_1142[11:3], u_ca_out_1141[20:12], u_ca_out_1140[23:21]};
assign col_out_1144 = {u_ca_out_1144[2:0],u_ca_out_1143[11:3], u_ca_out_1142[20:12], u_ca_out_1141[23:21]};
assign col_out_1145 = {u_ca_out_1145[2:0],u_ca_out_1144[11:3], u_ca_out_1143[20:12], u_ca_out_1142[23:21]};
assign col_out_1146 = {u_ca_out_1146[2:0],u_ca_out_1145[11:3], u_ca_out_1144[20:12], u_ca_out_1143[23:21]};
assign col_out_1147 = {u_ca_out_1147[2:0],u_ca_out_1146[11:3], u_ca_out_1145[20:12], u_ca_out_1144[23:21]};
assign col_out_1148 = {u_ca_out_1148[2:0],u_ca_out_1147[11:3], u_ca_out_1146[20:12], u_ca_out_1145[23:21]};
assign col_out_1149 = {u_ca_out_1149[2:0],u_ca_out_1148[11:3], u_ca_out_1147[20:12], u_ca_out_1146[23:21]};
assign col_out_1150 = {u_ca_out_1150[2:0],u_ca_out_1149[11:3], u_ca_out_1148[20:12], u_ca_out_1147[23:21]};
assign col_out_1151 = {u_ca_out_1151[2:0],u_ca_out_1150[11:3], u_ca_out_1149[20:12], u_ca_out_1148[23:21]};
assign col_out_1152 = {u_ca_out_1152[2:0],u_ca_out_1151[11:3], u_ca_out_1150[20:12], u_ca_out_1149[23:21]};
assign col_out_1153 = {u_ca_out_1153[2:0],u_ca_out_1152[11:3], u_ca_out_1151[20:12], u_ca_out_1150[23:21]};
assign col_out_1154 = {u_ca_out_1154[2:0],u_ca_out_1153[11:3], u_ca_out_1152[20:12], u_ca_out_1151[23:21]};
assign col_out_1155 = {u_ca_out_1155[2:0],u_ca_out_1154[11:3], u_ca_out_1153[20:12], u_ca_out_1152[23:21]};
assign col_out_1156 = {u_ca_out_1156[2:0],u_ca_out_1155[11:3], u_ca_out_1154[20:12], u_ca_out_1153[23:21]};
assign col_out_1157 = {u_ca_out_1157[2:0],u_ca_out_1156[11:3], u_ca_out_1155[20:12], u_ca_out_1154[23:21]};
assign col_out_1158 = {u_ca_out_1158[2:0],u_ca_out_1157[11:3], u_ca_out_1156[20:12], u_ca_out_1155[23:21]};
assign col_out_1159 = {u_ca_out_1159[2:0],u_ca_out_1158[11:3], u_ca_out_1157[20:12], u_ca_out_1156[23:21]};
assign col_out_1160 = {u_ca_out_1160[2:0],u_ca_out_1159[11:3], u_ca_out_1158[20:12], u_ca_out_1157[23:21]};
assign col_out_1161 = {u_ca_out_1161[2:0],u_ca_out_1160[11:3], u_ca_out_1159[20:12], u_ca_out_1158[23:21]};
assign col_out_1162 = {u_ca_out_1162[2:0],u_ca_out_1161[11:3], u_ca_out_1160[20:12], u_ca_out_1159[23:21]};
assign col_out_1163 = {u_ca_out_1163[2:0],u_ca_out_1162[11:3], u_ca_out_1161[20:12], u_ca_out_1160[23:21]};
assign col_out_1164 = {u_ca_out_1164[2:0],u_ca_out_1163[11:3], u_ca_out_1162[20:12], u_ca_out_1161[23:21]};
assign col_out_1165 = {u_ca_out_1165[2:0],u_ca_out_1164[11:3], u_ca_out_1163[20:12], u_ca_out_1162[23:21]};
assign col_out_1166 = {u_ca_out_1166[2:0],u_ca_out_1165[11:3], u_ca_out_1164[20:12], u_ca_out_1163[23:21]};
assign col_out_1167 = {u_ca_out_1167[2:0],u_ca_out_1166[11:3], u_ca_out_1165[20:12], u_ca_out_1164[23:21]};
assign col_out_1168 = {u_ca_out_1168[2:0],u_ca_out_1167[11:3], u_ca_out_1166[20:12], u_ca_out_1165[23:21]};
assign col_out_1169 = {u_ca_out_1169[2:0],u_ca_out_1168[11:3], u_ca_out_1167[20:12], u_ca_out_1166[23:21]};
assign col_out_1170 = {u_ca_out_1170[2:0],u_ca_out_1169[11:3], u_ca_out_1168[20:12], u_ca_out_1167[23:21]};
assign col_out_1171 = {u_ca_out_1171[2:0],u_ca_out_1170[11:3], u_ca_out_1169[20:12], u_ca_out_1168[23:21]};
assign col_out_1172 = {u_ca_out_1172[2:0],u_ca_out_1171[11:3], u_ca_out_1170[20:12], u_ca_out_1169[23:21]};
assign col_out_1173 = {u_ca_out_1173[2:0],u_ca_out_1172[11:3], u_ca_out_1171[20:12], u_ca_out_1170[23:21]};
assign col_out_1174 = {u_ca_out_1174[2:0],u_ca_out_1173[11:3], u_ca_out_1172[20:12], u_ca_out_1171[23:21]};
assign col_out_1175 = {u_ca_out_1175[2:0],u_ca_out_1174[11:3], u_ca_out_1173[20:12], u_ca_out_1172[23:21]};
assign col_out_1176 = {u_ca_out_1176[2:0],u_ca_out_1175[11:3], u_ca_out_1174[20:12], u_ca_out_1173[23:21]};
assign col_out_1177 = {u_ca_out_1177[2:0],u_ca_out_1176[11:3], u_ca_out_1175[20:12], u_ca_out_1174[23:21]};
assign col_out_1178 = {u_ca_out_1178[2:0],u_ca_out_1177[11:3], u_ca_out_1176[20:12], u_ca_out_1175[23:21]};
assign col_out_1179 = {u_ca_out_1179[2:0],u_ca_out_1178[11:3], u_ca_out_1177[20:12], u_ca_out_1176[23:21]};
assign col_out_1180 = {u_ca_out_1180[2:0],u_ca_out_1179[11:3], u_ca_out_1178[20:12], u_ca_out_1177[23:21]};
assign col_out_1181 = {u_ca_out_1181[2:0],u_ca_out_1180[11:3], u_ca_out_1179[20:12], u_ca_out_1178[23:21]};
assign col_out_1182 = {u_ca_out_1182[2:0],u_ca_out_1181[11:3], u_ca_out_1180[20:12], u_ca_out_1179[23:21]};
assign col_out_1183 = {u_ca_out_1183[2:0],u_ca_out_1182[11:3], u_ca_out_1181[20:12], u_ca_out_1180[23:21]};
assign col_out_1184 = {u_ca_out_1184[2:0],u_ca_out_1183[11:3], u_ca_out_1182[20:12], u_ca_out_1181[23:21]};
assign col_out_1185 = {u_ca_out_1185[2:0],u_ca_out_1184[11:3], u_ca_out_1183[20:12], u_ca_out_1182[23:21]};
assign col_out_1186 = {u_ca_out_1186[2:0],u_ca_out_1185[11:3], u_ca_out_1184[20:12], u_ca_out_1183[23:21]};
assign col_out_1187 = {u_ca_out_1187[2:0],u_ca_out_1186[11:3], u_ca_out_1185[20:12], u_ca_out_1184[23:21]};
assign col_out_1188 = {u_ca_out_1188[2:0],u_ca_out_1187[11:3], u_ca_out_1186[20:12], u_ca_out_1185[23:21]};
assign col_out_1189 = {u_ca_out_1189[2:0],u_ca_out_1188[11:3], u_ca_out_1187[20:12], u_ca_out_1186[23:21]};
assign col_out_1190 = {u_ca_out_1190[2:0],u_ca_out_1189[11:3], u_ca_out_1188[20:12], u_ca_out_1187[23:21]};
assign col_out_1191 = {u_ca_out_1191[2:0],u_ca_out_1190[11:3], u_ca_out_1189[20:12], u_ca_out_1188[23:21]};
assign col_out_1192 = {u_ca_out_1192[2:0],u_ca_out_1191[11:3], u_ca_out_1190[20:12], u_ca_out_1189[23:21]};
assign col_out_1193 = {u_ca_out_1193[2:0],u_ca_out_1192[11:3], u_ca_out_1191[20:12], u_ca_out_1190[23:21]};
assign col_out_1194 = {u_ca_out_1194[2:0],u_ca_out_1193[11:3], u_ca_out_1192[20:12], u_ca_out_1191[23:21]};
assign col_out_1195 = {u_ca_out_1195[2:0],u_ca_out_1194[11:3], u_ca_out_1193[20:12], u_ca_out_1192[23:21]};
assign col_out_1196 = {u_ca_out_1196[2:0],u_ca_out_1195[11:3], u_ca_out_1194[20:12], u_ca_out_1193[23:21]};
assign col_out_1197 = {u_ca_out_1197[2:0],u_ca_out_1196[11:3], u_ca_out_1195[20:12], u_ca_out_1194[23:21]};
assign col_out_1198 = {u_ca_out_1198[2:0],u_ca_out_1197[11:3], u_ca_out_1196[20:12], u_ca_out_1195[23:21]};
assign col_out_1199 = {u_ca_out_1199[2:0],u_ca_out_1198[11:3], u_ca_out_1197[20:12], u_ca_out_1196[23:21]};
assign col_out_1200 = {u_ca_out_1200[2:0],u_ca_out_1199[11:3], u_ca_out_1198[20:12], u_ca_out_1197[23:21]};
assign col_out_1201 = {u_ca_out_1201[2:0],u_ca_out_1200[11:3], u_ca_out_1199[20:12], u_ca_out_1198[23:21]};
assign col_out_1202 = {u_ca_out_1202[2:0],u_ca_out_1201[11:3], u_ca_out_1200[20:12], u_ca_out_1199[23:21]};
assign col_out_1203 = {u_ca_out_1203[2:0],u_ca_out_1202[11:3], u_ca_out_1201[20:12], u_ca_out_1200[23:21]};
assign col_out_1204 = {u_ca_out_1204[2:0],u_ca_out_1203[11:3], u_ca_out_1202[20:12], u_ca_out_1201[23:21]};
assign col_out_1205 = {u_ca_out_1205[2:0],u_ca_out_1204[11:3], u_ca_out_1203[20:12], u_ca_out_1202[23:21]};
assign col_out_1206 = {u_ca_out_1206[2:0],u_ca_out_1205[11:3], u_ca_out_1204[20:12], u_ca_out_1203[23:21]};
assign col_out_1207 = {u_ca_out_1207[2:0],u_ca_out_1206[11:3], u_ca_out_1205[20:12], u_ca_out_1204[23:21]};
assign col_out_1208 = {u_ca_out_1208[2:0],u_ca_out_1207[11:3], u_ca_out_1206[20:12], u_ca_out_1205[23:21]};
assign col_out_1209 = {u_ca_out_1209[2:0],u_ca_out_1208[11:3], u_ca_out_1207[20:12], u_ca_out_1206[23:21]};
assign col_out_1210 = {u_ca_out_1210[2:0],u_ca_out_1209[11:3], u_ca_out_1208[20:12], u_ca_out_1207[23:21]};
assign col_out_1211 = {u_ca_out_1211[2:0],u_ca_out_1210[11:3], u_ca_out_1209[20:12], u_ca_out_1208[23:21]};
assign col_out_1212 = {u_ca_out_1212[2:0],u_ca_out_1211[11:3], u_ca_out_1210[20:12], u_ca_out_1209[23:21]};
assign col_out_1213 = {u_ca_out_1213[2:0],u_ca_out_1212[11:3], u_ca_out_1211[20:12], u_ca_out_1210[23:21]};
assign col_out_1214 = {u_ca_out_1214[2:0],u_ca_out_1213[11:3], u_ca_out_1212[20:12], u_ca_out_1211[23:21]};
assign col_out_1215 = {u_ca_out_1215[2:0],u_ca_out_1214[11:3], u_ca_out_1213[20:12], u_ca_out_1212[23:21]};
assign col_out_1216 = {u_ca_out_1216[2:0],u_ca_out_1215[11:3], u_ca_out_1214[20:12], u_ca_out_1213[23:21]};
assign col_out_1217 = {u_ca_out_1217[2:0],u_ca_out_1216[11:3], u_ca_out_1215[20:12], u_ca_out_1214[23:21]};
assign col_out_1218 = {u_ca_out_1218[2:0],u_ca_out_1217[11:3], u_ca_out_1216[20:12], u_ca_out_1215[23:21]};
assign col_out_1219 = {u_ca_out_1219[2:0],u_ca_out_1218[11:3], u_ca_out_1217[20:12], u_ca_out_1216[23:21]};
assign col_out_1220 = {u_ca_out_1220[2:0],u_ca_out_1219[11:3], u_ca_out_1218[20:12], u_ca_out_1217[23:21]};
assign col_out_1221 = {u_ca_out_1221[2:0],u_ca_out_1220[11:3], u_ca_out_1219[20:12], u_ca_out_1218[23:21]};
assign col_out_1222 = {u_ca_out_1222[2:0],u_ca_out_1221[11:3], u_ca_out_1220[20:12], u_ca_out_1219[23:21]};
assign col_out_1223 = {u_ca_out_1223[2:0],u_ca_out_1222[11:3], u_ca_out_1221[20:12], u_ca_out_1220[23:21]};
assign col_out_1224 = {u_ca_out_1224[2:0],u_ca_out_1223[11:3], u_ca_out_1222[20:12], u_ca_out_1221[23:21]};
assign col_out_1225 = {u_ca_out_1225[2:0],u_ca_out_1224[11:3], u_ca_out_1223[20:12], u_ca_out_1222[23:21]};
assign col_out_1226 = {u_ca_out_1226[2:0],u_ca_out_1225[11:3], u_ca_out_1224[20:12], u_ca_out_1223[23:21]};
assign col_out_1227 = {u_ca_out_1227[2:0],u_ca_out_1226[11:3], u_ca_out_1225[20:12], u_ca_out_1224[23:21]};
assign col_out_1228 = {u_ca_out_1228[2:0],u_ca_out_1227[11:3], u_ca_out_1226[20:12], u_ca_out_1225[23:21]};
assign col_out_1229 = {u_ca_out_1229[2:0],u_ca_out_1228[11:3], u_ca_out_1227[20:12], u_ca_out_1226[23:21]};
assign col_out_1230 = {u_ca_out_1230[2:0],u_ca_out_1229[11:3], u_ca_out_1228[20:12], u_ca_out_1227[23:21]};
assign col_out_1231 = {u_ca_out_1231[2:0],u_ca_out_1230[11:3], u_ca_out_1229[20:12], u_ca_out_1228[23:21]};
assign col_out_1232 = {u_ca_out_1232[2:0],u_ca_out_1231[11:3], u_ca_out_1230[20:12], u_ca_out_1229[23:21]};
assign col_out_1233 = {u_ca_out_1233[2:0],u_ca_out_1232[11:3], u_ca_out_1231[20:12], u_ca_out_1230[23:21]};
assign col_out_1234 = {u_ca_out_1234[2:0],u_ca_out_1233[11:3], u_ca_out_1232[20:12], u_ca_out_1231[23:21]};
assign col_out_1235 = {u_ca_out_1235[2:0],u_ca_out_1234[11:3], u_ca_out_1233[20:12], u_ca_out_1232[23:21]};
assign col_out_1236 = {u_ca_out_1236[2:0],u_ca_out_1235[11:3], u_ca_out_1234[20:12], u_ca_out_1233[23:21]};
assign col_out_1237 = {u_ca_out_1237[2:0],u_ca_out_1236[11:3], u_ca_out_1235[20:12], u_ca_out_1234[23:21]};
assign col_out_1238 = {u_ca_out_1238[2:0],u_ca_out_1237[11:3], u_ca_out_1236[20:12], u_ca_out_1235[23:21]};
assign col_out_1239 = {u_ca_out_1239[2:0],u_ca_out_1238[11:3], u_ca_out_1237[20:12], u_ca_out_1236[23:21]};
assign col_out_1240 = {u_ca_out_1240[2:0],u_ca_out_1239[11:3], u_ca_out_1238[20:12], u_ca_out_1237[23:21]};
assign col_out_1241 = {u_ca_out_1241[2:0],u_ca_out_1240[11:3], u_ca_out_1239[20:12], u_ca_out_1238[23:21]};
assign col_out_1242 = {u_ca_out_1242[2:0],u_ca_out_1241[11:3], u_ca_out_1240[20:12], u_ca_out_1239[23:21]};
assign col_out_1243 = {u_ca_out_1243[2:0],u_ca_out_1242[11:3], u_ca_out_1241[20:12], u_ca_out_1240[23:21]};
assign col_out_1244 = {u_ca_out_1244[2:0],u_ca_out_1243[11:3], u_ca_out_1242[20:12], u_ca_out_1241[23:21]};
assign col_out_1245 = {u_ca_out_1245[2:0],u_ca_out_1244[11:3], u_ca_out_1243[20:12], u_ca_out_1242[23:21]};
assign col_out_1246 = {u_ca_out_1246[2:0],u_ca_out_1245[11:3], u_ca_out_1244[20:12], u_ca_out_1243[23:21]};
assign col_out_1247 = {u_ca_out_1247[2:0],u_ca_out_1246[11:3], u_ca_out_1245[20:12], u_ca_out_1244[23:21]};
assign col_out_1248 = {u_ca_out_1248[2:0],u_ca_out_1247[11:3], u_ca_out_1246[20:12], u_ca_out_1245[23:21]};
assign col_out_1249 = {u_ca_out_1249[2:0],u_ca_out_1248[11:3], u_ca_out_1247[20:12], u_ca_out_1246[23:21]};
assign col_out_1250 = {u_ca_out_1250[2:0],u_ca_out_1249[11:3], u_ca_out_1248[20:12], u_ca_out_1247[23:21]};
assign col_out_1251 = {u_ca_out_1251[2:0],u_ca_out_1250[11:3], u_ca_out_1249[20:12], u_ca_out_1248[23:21]};
assign col_out_1252 = {u_ca_out_1252[2:0],u_ca_out_1251[11:3], u_ca_out_1250[20:12], u_ca_out_1249[23:21]};
assign col_out_1253 = {u_ca_out_1253[2:0],u_ca_out_1252[11:3], u_ca_out_1251[20:12], u_ca_out_1250[23:21]};
assign col_out_1254 = {u_ca_out_1254[2:0],u_ca_out_1253[11:3], u_ca_out_1252[20:12], u_ca_out_1251[23:21]};
assign col_out_1255 = {u_ca_out_1255[2:0],u_ca_out_1254[11:3], u_ca_out_1253[20:12], u_ca_out_1252[23:21]};
assign col_out_1256 = {u_ca_out_1256[2:0],u_ca_out_1255[11:3], u_ca_out_1254[20:12], u_ca_out_1253[23:21]};
assign col_out_1257 = {u_ca_out_1257[2:0],u_ca_out_1256[11:3], u_ca_out_1255[20:12], u_ca_out_1254[23:21]};
assign col_out_1258 = {u_ca_out_1258[2:0],u_ca_out_1257[11:3], u_ca_out_1256[20:12], u_ca_out_1255[23:21]};
assign col_out_1259 = {u_ca_out_1259[2:0],u_ca_out_1258[11:3], u_ca_out_1257[20:12], u_ca_out_1256[23:21]};
assign col_out_1260 = {u_ca_out_1260[2:0],u_ca_out_1259[11:3], u_ca_out_1258[20:12], u_ca_out_1257[23:21]};
assign col_out_1261 = {u_ca_out_1261[2:0],u_ca_out_1260[11:3], u_ca_out_1259[20:12], u_ca_out_1258[23:21]};
assign col_out_1262 = {u_ca_out_1262[2:0],u_ca_out_1261[11:3], u_ca_out_1260[20:12], u_ca_out_1259[23:21]};
assign col_out_1263 = {u_ca_out_1263[2:0],u_ca_out_1262[11:3], u_ca_out_1261[20:12], u_ca_out_1260[23:21]};
assign col_out_1264 = {u_ca_out_1264[2:0],u_ca_out_1263[11:3], u_ca_out_1262[20:12], u_ca_out_1261[23:21]};
assign col_out_1265 = {u_ca_out_1265[2:0],u_ca_out_1264[11:3], u_ca_out_1263[20:12], u_ca_out_1262[23:21]};
assign col_out_1266 = {u_ca_out_1266[2:0],u_ca_out_1265[11:3], u_ca_out_1264[20:12], u_ca_out_1263[23:21]};
assign col_out_1267 = {u_ca_out_1267[2:0],u_ca_out_1266[11:3], u_ca_out_1265[20:12], u_ca_out_1264[23:21]};
assign col_out_1268 = {u_ca_out_1268[2:0],u_ca_out_1267[11:3], u_ca_out_1266[20:12], u_ca_out_1265[23:21]};
assign col_out_1269 = {u_ca_out_1269[2:0],u_ca_out_1268[11:3], u_ca_out_1267[20:12], u_ca_out_1266[23:21]};
assign col_out_1270 = {u_ca_out_1270[2:0],u_ca_out_1269[11:3], u_ca_out_1268[20:12], u_ca_out_1267[23:21]};
assign col_out_1271 = {u_ca_out_1271[2:0],u_ca_out_1270[11:3], u_ca_out_1269[20:12], u_ca_out_1268[23:21]};
assign col_out_1272 = {u_ca_out_1272[2:0],u_ca_out_1271[11:3], u_ca_out_1270[20:12], u_ca_out_1269[23:21]};
assign col_out_1273 = {u_ca_out_1273[2:0],u_ca_out_1272[11:3], u_ca_out_1271[20:12], u_ca_out_1270[23:21]};
assign col_out_1274 = {u_ca_out_1274[2:0],u_ca_out_1273[11:3], u_ca_out_1272[20:12], u_ca_out_1271[23:21]};
assign col_out_1275 = {u_ca_out_1275[2:0],u_ca_out_1274[11:3], u_ca_out_1273[20:12], u_ca_out_1272[23:21]};
assign col_out_1276 = {u_ca_out_1276[2:0],u_ca_out_1275[11:3], u_ca_out_1274[20:12], u_ca_out_1273[23:21]};
assign col_out_1277 = {u_ca_out_1277[2:0],u_ca_out_1276[11:3], u_ca_out_1275[20:12], u_ca_out_1274[23:21]};
assign col_out_1278 = {u_ca_out_1278[2:0],u_ca_out_1277[11:3], u_ca_out_1276[20:12], u_ca_out_1275[23:21]};
assign col_out_1279 = {u_ca_out_1279[2:0],u_ca_out_1278[11:3], u_ca_out_1277[20:12], u_ca_out_1276[23:21]};
assign col_out_1280 = {u_ca_out_1280[2:0],u_ca_out_1279[11:3], u_ca_out_1278[20:12], u_ca_out_1277[23:21]};
assign col_out_1281 = {u_ca_out_1281[2:0],u_ca_out_1280[11:3], u_ca_out_1279[20:12], u_ca_out_1278[23:21]};
assign col_out_1282 = {u_ca_out_1282[2:0],u_ca_out_1281[11:3], u_ca_out_1280[20:12], u_ca_out_1279[23:21]};
assign col_out_1283 = {{3{1'b0}}, u_ca_out_1282[11:3], u_ca_out_1281[20:12], u_ca_out_1280[23:21]};
assign col_out_1284 = {{12{1'b0}}, u_ca_out_1282[20:12], u_ca_out_1281[23:21]};
assign col_out_1285 = {{21{1'b0}}, u_ca_out_1282[23:21]};

//---------------------------------------------------------


endmodule
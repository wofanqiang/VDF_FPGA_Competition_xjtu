module xpb_5_35
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h912f150517db24abfd766457ffdf2718f19fb9dcbc3f03426e11e1e43a79a8481592c42716407c1cd00d87fef23bea4aa9adf9d482c19b78c8e5759b7cd14b0c6d1027f79e58bba2e5e52d9d01275e3b8f6677525bb00b3ac5715eb26dbd073be8ac62687e2cfa4d4973fd6fd5bfd29c5615fae23b230c1d2e7de121a3c9de58;
    5'b00010 : xpb = 1024'h71b0e4b46dc8148f2fe750d8ef6406e071c97088a306660d5e470a72c1f0a38827dd0ad5625a79ab00bcd0b70119c3caef41cbc2e2d066a5e12babd8bed0216765d11b408d207a00b93058976972f8462ac7f50c2ad9e964d5562b6a214f6be5a25132a74b90fc0d0c281400b3af7f0f5d5216e225fabb0a168c473ebeb15645;
    5'b00011 : xpb = 1024'h5232b463c3b5047262583d59dee8e6a7f1f3273489cdc8d84e7c330149679ec83a275183ae747739316c196f0ff79d4b34d59db142df31d2f971e21600cef7c25e920e897be8385e8c7b8391d1be9250c62972c5fa03c78ee53af821d4e1d08f5bf602e618f4fdcccedc2a91919f2b82648e32e210d269f6fe9aad5bd998ce32;
    5'b00100 : xpb = 1024'h32b4841319a1f45594c929dace6dc66f721cdde070952ba33eb15b8fd0de9a084c719831fa8e74c7621b62271ed576cb7a696f9fa2edfd0011b8185342cdce1d575301d26aaff6bc5fc6ae8c3a0a2c5b618af07fc92da5b8f51fc4d988743539159ad324e658ff8c919041226f8ed7f56bca4ee1fbaa18e3e6a91378f480461f;
    5'b00101 : xpb = 1024'h133653c26f8ee438c73a165bbdf2a636f246948c575c8e6e2ee6841e585595485ebbdee046a8725592caaadf2db3504bbffd418e02fcc82d29fe4e9084cca4785013f51b5977b51a3311d986a255c665fcec6e39985783e3050491913c0699e2cf3fa363b3bd014c544457b34d7e846873066ae1e681c7d0ceb779960f67be0c;
    5'b00110 : xpb = 1024'ha46568c7876a08e4c4b07ab3bdd1cd4fe3e64e69139b91b09cf8660292cf3d90744ea3075ce8ee7262d832de1fef3a9669ab3b6285be63a5f2e3c42c019def84bd241d12f7d070bd18f70723a37d24a18c52e58bf4078f1dca75f043a9c3a11eb7ec05cc31e9fb999db85523233e5704c91c65c421a4d3edfd355ab7b3319c64;
    5'b00111 : xpb = 1024'h84e73876dd56f8c7f7216734ad56ad1764100514fa62f47b8d2d8e911a4638d08698e9b5a902ec0093877b962ecd1416af3f0d50e5cd2ed30b29fa69439cc5dfb5e5105be6982f1aec42321e0bc8beac27b46345c3316d47da5abcfb5d5605c87190d60aff4dfd59606c6bb4012e0377d05881c40c7c82dae543c0d4ce191451;
    5'b01000 : xpb = 1024'h656908263343e8ab299253b59cdb8cdee439bbc0e12a57467d62b71fa1bd341098e33063f51ce98ec436c44e3daaed96f4d2df3f45dbfa00237030a6859b9c3aaea603a4d55fed78bf8d5d18741458b6c315e0ff925b4b71ea3f89b310e86a722b35a649ccb1ff1923208244df1dafead7949dc3f75431c7cd5226f1e9008c3e;
    5'b01001 : xpb = 1024'h45ead7d58930d88e5c0340368c606ca66463726cc7f1ba116d97dfae29342f50ab2d77124136e71cf4e60d064c88c7173a66b12da5eac52d3bb666e3c79a7295a766f6edc427abd692d88812dc5ff2c15e775eb96185299bfa24566ac47acf1be4da76889a1600d8e5d498d5bd0d5c5dded0b9c3e22be0b4b5608d0f03e8042b;
    5'b01010 : xpb = 1024'h266ca784df1dc8718e742cb77be54c6de48d2918aeb91cdc5dcd083cb0ab2a90bd77bdc08d50e4ab259555be5b66a0977ffa831c05f9905a53fc9d21099948f0a027ea36b2ef6a346623b30d44ab8ccbf9d8dc7330af07c60a092322780d33c59e7f46c7677a0298a888af669afd08d0e60cd5c3cd038fa19d6ef32c1ecf7c18;
    5'b01011 : xpb = 1024'h6ee7734350ab854c0e519386b6a2c3564b6dfc495807fa74e0230cb382225d0cfc2046ed96ae23956449e766a447a17c58e550a66085b876c42d35e4b981f4b98e8dd7fa1b72892396ede07acf726d6953a5a2cffd8e5f019edefda2b9f986f5824170634de04586b3cc5f778ecb543ed48f1c3b7db3e8e857d594939b6f405;
    5'b01100 : xpb = 1024'h981d8c394ce5dd00be5b7d906b49534e565699a151bf82e9bc1412af729bce18e554c895efab5e56265226755c8064626f3c4edee8c9f700352848f9c8696a5805f90577400fe4351f540ba4ae1e851224a0d17f5b88f12adf5f4e8c995c9fab40d0796eb30afea5b4b0c3674eac87e0435eeca5f2fe4aabb3fb3a6add80d25d;
    5'b01101 : xpb = 1024'h789f5be8a2d2cce3f0cc6a115ace3315d680504d3886e5b4ac493b3dfa12c958f79f0f443bc55be457016f2d6b5e3de2b4d020cd48d8c22d4d6e7f370a6840b2feb9f8c02ed7a292f29f369f166a1f1cc0024f392ab2cf54ef441b444cef0454fa7549ad806f00657764d9f82c9c34534a9b08a5ddd5f9989c09a087f8684a4a;
    5'b01110 : xpb = 1024'h59212b97f8bfbcc7233d56924a5312dd56aa06f91f4e487f9c7e63cc8189c49909e955f287df597287b0b7e57a3c1762fa63f2bba8e78d5a65b4b5744c67170df77aec091d9f60f0c5ea61997eb5b9275b63ccf2f9dcad7eff28e7fc008168feb41a19ec4dd302253a18f0890a8be0c651d724a5c8ada885841806a5134fc237;
    5'b01111 : xpb = 1024'h39a2fb474eacacaa55ae431339d7f2a4d6d3bda50615ab4a8cb38c5b0900bfd91c339ca0d3f95700b860009d8919f0e33ff7c4aa08f658877dfaebb18e65ed68f03bdf520c671f4e99358c93e7015331f6c54aacc9068ba90f0db4b3b413cda86dbeea2b1b3703e4fccd0719e87b8d39591340a5b38557726c266cc22e373a24;
    5'b10000 : xpb = 1024'h1a24caf6a4999c8d881f2f94295cd26c56fd7450ecdd0e157ce8b4e99077bb192e7de34f2013548ee90f495597f7ca63858b9698690523b4964121eed064c3c3e8fcd29afb2eddac6c80b78e4f4ced3c9226c866983069d31ef2816b67a632522763ba69e89b05a4bf811daac66b39ac604f5ca59e5d065f5434d2df491eb211;
    5'b10001 : xpb = 1024'hab53dffbbc74c139859593ec293bf985489d2e2da91c1157eafa96cdcaf163614410a7763653d0abb91cd1548a33b4ae2f39906cebc6bf2d5f26978a4d360ed0560cfa929987994f5265e52b50744b78218d3fb8f3e0750de463e01dd563398e10101cd266c7fff208f51b1a9c2b0c48b6655787d980127c82b2b400ece89069;
    5'b10010 : xpb = 1024'h8bd5afab1261b11cb806806d18c0d94cc8c6e4d98fe37422db2fbf5c52685ea1565aee24826dce39e9cc1a0c99118e2e74cd625b4bd58a5a776ccdc78f34e52b4ecdeddb884f57ad25b11025b8bfe582bceebd72c30a5337f448acd588f59e37c9b4ed11342c01b1cba931ab7a1ab8bbbda17387c457c1696ac11a1e07d00856;
    5'b10011 : xpb = 1024'h6c577f5a684ea0ffea776cee0845b91448f09b8576aad6edcb64e7ead9df59e168a534d2ce87cbc81a7b62c4a7ef67aeba613449abe455878fb30404d133bb86478ee1247717160af8fc3b20210b7f8d58503b2c92343162042d798d3c8802e18359bd50019003718e5d483c580a652ec4dd8f87af2f705652cf803b22b78043;
    5'b10100 : xpb = 1024'h4cd94f09be3b90e31ce8596ef7ca98dbc91a52315d7239b8bb9a1079615655217aef7b811aa1c9564b2aab7cb6cd412efff506380bf320b4a7f93a42133291e1404fd46d65ded468cc47661a89571997f3b1b8e6615e0f8c14124644f01a678b3cfe8d8ecef4053151115ecd35fa11a1cc19ab879a071f433adde6583d9ef830;
    5'b10101 : xpb = 1024'h2d5b1eb9142880c64f5945efe74f78a3494408dd44399c83abcf3907e8cd50618d39c22f66bbc6e47bd9f434c5ab1aaf4588d8266c01ebe1c03f707f5531683c3910c7b654a692c69f929114f1a2b3a28f1336a03087edb623f712fca3accc34f6a35dcd9c5806f113c5755e13e9be14d355c78784dece3022ec4c755886701d;
    5'b10110 : xpb = 1024'hddcee686a1570a981ca3270d6d4586ac96dbf892b00ff4e9c04619670444ba19f8408ddb2d5c472ac893cecd488f42f8b1caa14cc10b70ed885a6bc97303e9731d1baff436e512472ddbc0f59ee4dad2a74b459ffb1cbe033dbdfb4573f30deb0482e0c69bc08b0d6798beef1d96a87da91e3876fb67d1d0afab292736de80a;
    5'b10111 : xpb = 1024'h9f0c036d81f095557f4096c8d6b37f83bb0d7965e74002910a16437aaabdf3e9b516cd04c916408f7c96c4ebc6c4de7a34caa3e94ed25287a16b1c58140189a39ee1e2f6e1c70cc758c2e9ac5b15abe8b9db2bac5b61d71af94d3e66c4fc381a98f49074e7e902fe1fed895ec7993d2430a7de69aad9893a397893b41737c662;
    5'b11000 : xpb = 1024'h7f8dd31cd7dd8538b1b18349c6385f4b3b373011ce07655bfa4b6c093234ef29c76113b315303e1dad460da3d5a2b7fa7a5e75d7aee11db4b9b1529556005ffe97a2d63fd08ecb252c0e14a6c36145f3553ca9662a8bb54509320b1e788e9cc4529960b3b54d04bde2a19fefa588e99737e3fa6995b138272186f9d1321f3e4f;
    5'b11001 : xpb = 1024'h600fa2cc2dca751be4226fcab5bd3f12bb60e6bdb4cec826ea809497b9abea69d9ab5a61614a3babddf5565be480917abff247c60eefe8e1d1f788d297ff36599063c988bf568982ff593fa12bacdffdf09e271ff9b5936f1916d7d62c21016e0c3e30f282b1067da555b6808378960a3f2016698088e71409955fee4d06b63c;
    5'b11010 : xpb = 1024'h4091727b83b764ff16935c4ba5421eda3b8a9d699b962af1dab5bd264122e5a9ebf5a10fad64393a0ea49f13f35e6afb058619b46efeb40eea3dbf0fd9fe0cb48924bcd1ae1e47e0d2a46a9b93f87a088bffa4d9c8df719928fba48ddfb36617c5e301315015083d6809cd116168427d465c32696b609600f1a3c60b67ee2e29;
    5'b11011 : xpb = 1024'h2113422ad9a454e2490448cc94c6fea1bbb45415825d8dbccaeae5b4c899e0e9fe3fe7bdf97e36c83f53e7cc023c447b4b19eba2cf0d7f3c0283f54d1bfce30f81e5b01a9ce6063ea5ef9595fc4414132761229398094fc338e071459345cac17f87d1701d7909fd2abde3a23f57eef04d984e69563844edd9b22c2882d5a616;
    5'b11100 : xpb = 1024'h19511da2f9144c57b75354d844bde693bde0ac16924f087bb200e435010dc2a108a2e6c4598345670033084111a1dfb90adbd912f1c4a691aca2b8a5dfbb96a7aa6a3638badc49c793ac090648fae1dc2c2a04d67332ded48c53dfd46d82f6b392ca1aeeadd0bbced71fa331d479b6354d46a69410ff3dac1c092459dbd1e03;
    5'b11101 : xpb = 1024'h92c426df476c697178eb99a5842b05822d7dc49e2563f3ca2931f0278a8a8472261cf2935bd8b0734010b883035608463a5bb765b1dde5e1e3afa125dacd0476e7b6cb5b2a06803f5f1fee2d65b70c595229179fc2e339280e369cafb49536a721d90417690a060a36e5f7a2f3076dffaaea654b7c32fff7f03e73674186fc5b;
    5'b11110 : xpb = 1024'h7345f68e9d595954ab5c862673afe549ada77b4a0c2b5695196718b612017fb238673941a7f2ae0170c0013b1233e1c67fef895411ecb10efbf5d7631ccbdad1e077bea418ce3e9d326b1927ce02a663ed8a9559920d17521e1b696768279b50db7dd456366e07c9f99a0e33d0f71a72b226814b670aaee4d84cd9845c6e7448;
    5'b11111 : xpb = 1024'h53c7c63df3464937ddcd72a76334c5112dd131f5f2f2b960099c414499787af24ab17feff40cab8fa16f49f32111bb46c5835b4271fb7c3c143c0da05ecab12cd938b1ed0795fcfb05b64422364e406e88ec13136136f57c2e00361f1bb9fffa9522a49503d20989bc4e24c4aee6c6e5b9629d4b51e25dd1c05b3fa17755ec35;
    endcase
end

endmodule

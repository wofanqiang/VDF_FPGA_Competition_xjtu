module xpb_5_150
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h21d8277d18b2cdc784427c177399eb068d4b035c9b7e8752b214905604ee03e4683d0e9cd594d71e97cdb5239a6a3141beac1de41b657ec2e05851d2e9d65ac70e8d845d73e732bf797e445d25530fda83cbd910a4957d0f479b9f3e8d741cc1387fb935527329022ff7aae3f795e09bb2174f9884a1efeb9a81775d10b9fee0;
    5'b00010 : xpb = 1024'h43b04efa31659b8f0884f82ee733d60d1a9606b936fd0ea5642920ac09dc07c8d07a1d39ab29ae3d2f9b6a4734d462837d583bc836cafd85c0b0a3a5d3acb58e1d1b08bae7ce657ef2fc88ba4aa61fb50797b221492afa1e8f373e7d1ae8398270ff726aa4e652045fef55c7ef2bc137642e9f310943dfd73502eeba2173fdc0;
    5'b00011 : xpb = 1024'h658876774a1869568cc774465acdc113a7e10a15d27b95f8163db1020eca0bad38b72bd680be855bc7691f6acf3e93c53c0459ac52307c48a108f578bd8310552ba88d185bb5983e6c7acd176ff92f8f8b638b31edc0772dd6d2ddbba85c5643a97f2b9ff7597b068fe700abe6c1a1d31645eec98de5cfc2cf846617322dfca0;
    5'b00100 : xpb = 1024'h87609df462cb371e1109f05dce67ac1a352c0d726dfa1d4ac852415813b80f91a0f43a7356535c7a5f36d48e69a8c506fab077906d95fb0b8161474ba7596b1c3a361175cf9ccafde5f91174954c3f6a0f2f64429255f43d1e6e7cfa35d07304e1fee4d549cca408bfdeab8fde57826ec85d3e621287bfae6a05dd7442e7fb80;
    5'b00101 : xpb = 1024'ha938c5717b7e04e5954c6c7542019720c27710cf0978a49d7a66d1ae18a61376093149102be83398f70489b20412f648b95c957488fb79ce61b9991e912fc5e348c395d34383fdbd5f7755d1ba9f4f4492fb3d5336eb714c660a1c38c3448fc61a7e9e0a9c3fcd0aefd65673d5ed630a7a748dfa9729af9a048754d153a1fa60;
    5'b00110 : xpb = 1024'h1a63a798d2429de44e8970b5a5413ad5de4c10facf7f8b78ae9ea8ae6a916a526e25da3437568c28ef73ff8ebb1f16c013ee8b7281ae28459172ab934033abf8e301e58207da3337c65b978c47169aee22c21ccb4efac14af819297c968e09f523f6c5163de9fd7f990e1a78d5b31d7cddb1feb0cb80425558995129db7992d5;
    5'b00111 : xpb = 1024'h3c3bcf15eaf56babd2cbeccd18db25dc6b9714576afe12cb60b339046f7f6e36d662e8d10ceb63478741b4b255894801d29aa9569d13a70871cafd662a0a06bff18f69df7bc165f73fd9dbe96c69aac8a68df5dbf3903e5a3fb4c8bb240226b65c767e4b905d2681c905c55ccd48fe188fc94e4950223240f31ac886ec3391b5;
    5'b01000 : xpb = 1024'h5e13f69303a83973570e68e48c7510e2f8e217b4067c9a1e12c7c95a746d721b3e9ff76de2803a661f0f69d5eff379439146c73ab87925cb52234f3913e06187001cee3cefa898b6b958204691bcbaa32a59ceec9825bb69875067f9b176437794f63780e2d04f83f8fd7040c4dedeb441e09de1d4c4222c8d9c3fe3fced9095;
    5'b01001 : xpb = 1024'h7fec1e101c5b073adb50e4fc000efbe9862d1b10a1fb2170c4dc59b0795b75ffa6dd060ab8151184b6dd1ef98a5daa854ff2e51ed3dea48e327ba10bfdb6bc4e0eaa729a638fcb7632d664a3b70fca7dae25a7fd3cbb3878ceec07383eea6038cd75f0b63543788628f51b24bc74bf4ff3f7ed7a59661218281db7410da78f75;
    5'b01010 : xpb = 1024'ha1c4458d350dd5025f93611373a8e6f013781e6d3d79a8c376f0ea067e4979e40f1a14a78da9e8a34eaad41d24c7dbc70e9f0302ef44235112d3f2dee78d17151d37f6f7d776fe35ac54a900dc62da5831f1810de150b5881687a676cc5e7cfa05f5a9eb87b6a18858ecc608b40a9feba60f3d12de080203c29f2e9e1e618e55;
    5'b01011 : xpb = 1024'h12ef27b48bd26e0118d06553d6e88aa52f4d1e9903808f9eab28c106d034d0c0740ea5cb99184133471a49f9dbd3fc3e6930f900e7f6d1c8428d05539690fd2ab77646a69bcd33b01338eabb68da2601c1b86085f9600586a896b3ba9fa7f7290f6dd0f72960d1fd02248a0db3d05a5e094cadc9125e94bf16b12af6a63926ca;
    5'b01100 : xpb = 1024'h34c74f31a4853bc89d12e16b4a8275abbc9821f59eff16f15d3d515cd522d4a4dc4bb4686ead1851dee7ff1d763e2d8027dd16e5035c508b22e55726806757f1c603cb040fb4666f8cb72f188e2d35dc458439969df58295f03252f92d1c13ea47ed8a2c7bd3faff321c34f1ab663af9bb63fd61970084aab132a253b6f325aa;
    5'b01101 : xpb = 1024'h569f76aebd38099021555d82be1c60b249e325523a7d9e440f51e1b2da10d8894488c3054441ef7076b5b44110a85ec1e68934c91ec1cf4e033da8f96a3db2b8d4914f61839b992f06357375b38045b6c95012a7428affa537cdf237ba9030ab806d4361ce4724016213dfd5a2fc1b956d7b4cfa1ba274964bb419b0c7ad248a;
    5'b01110 : xpb = 1024'h78779e2bd5ead757a597d99a31b64bb8d72e28aed5fc2596c1667208defedc6dacc5d1a219d6c68f0e836964ab129003a53552ad3a274e10e395facc54140d7fe31ed3bef782cbee7fb3b7d2d8d355914d1bebb7e7207cb47f69917648044d6cb8ecfc9720ba4d03920b8ab99a91fc311f929c92a0446481e635910dd867236a;
    5'b01111 : xpb = 1024'h9a4fc5a8ee9da51f29da55b1a55036bf64792c0b717aace9737b025ee3ece0521502e03eef6b9dada6511e88457cc14563e17091558cccd3c3ee4c9f3dea6846f1ac581c6b69feadf931fc2ffe26656bd0e7c4c88bb5f9c3c70530b4d5786a2df16cb5cc732d7605c203359d9227dcccd1a9ec2b24e6546d80b7086ae921224a;
    5'b10000 : xpb = 1024'hb7aa7d045623e1de31759f2088fda74804e2c37378193c4a7b2d95f35d8372e79f77162fad9f63d9ec09464fc88e1bcbe73668f4e3f7b4af3a75f13ecee4e5c8beaa7cb2fc0342860163dea8a9db11560aea440a3c549c259143df8a8c1e45cfae4dcd814d7a67a6b3af9a291ed973f34e75ce1593ce728d4c904c370f8babf;
    5'b10001 : xpb = 1024'h2d52cf4d5e150be56759d6097c29c57b0d992f93d3001b1759c769b53ac63b12e2347fffd06ecd5c368e498896f312fe7d1f847369a4fa0dd3ffb0e6d6c4a9239a782c28a3a766e7d9948247aff0c0efe47a7d51485ac6d1a0afdd373636011e3364960d674acf7c9b32a486898377dae6feac79ddded7146f4a7c2081b2b99f;
    5'b10010 : xpb = 1024'h4f2af6ca76c7d9aceb9c5220efc3b0819ae432f06e7ea26a0bdbfa0b3fb43ef74a718e9ca603a47ace5bfeac315d44403bcba257850a78d0b45802b9c09b03eaa905b086178e99a75312c6a4d543d0ca68465661ecf043e0e84b7c75c3aa1ddf6be44f42b9bdf87ecb2a4f6a811958769915fc126280c70009cbf37d926cb87f;
    5'b10011 : xpb = 1024'h71031e478f7aa7746fdece38635d9b88282f364d09fd29bcbdf08a6144a242dbb2ae9d397b987b996629b3cfcbc77581fa77c03ba06ff79394b0548caa715eb1b79334e38b75cc66cc910b01fa96e0a4ec122f729185c0f02fe71bb4511e3aa0a46408780c312180fb21fa4e78af39124b2d4baae722b6eba44d6adaa326b75f;
    5'b10100 : xpb = 1024'h92db45c4a82d753bf4214a4fd6f7868eb57a39a9a57bb10f70051ab7499046c01aebabd6512d52b7fdf768f36631a6c3b923de1fbbd576567508a65f9447b978c620b940ff5cff26460f4f5f1fe9f07f6fde0883361b3dff7782baf2de925761dce3c1ad5ea44a832b19a532704519adfd449b436bc4a6d73ecee237b3e0b63f;
    5'b10101 : xpb = 1024'h40627ebfef20e3aad5e4e903a372a43d14f39d56b8297eaa43cf1b79b7b9d9c7fe03cfa5c9bab47f666ded01d3dc73b13b5d41db48824cda4c1b8d4434b9f8e605f08efc3b334a0acf39119ac613c28ffa4e7fb4e2a8dfe0991c836b1dbd190e65be8b9004e7af7d4516937700ad42060820bf9a01b399292e0de903bb84eb4;
    5'b10110 : xpb = 1024'h25de4f6917a4dc0231a0caa7add1154a5e9a3d3207011f3d5651820da069a180e81d4b97323082668e3493f3b7a7f87cd261f201cfeda390851a0aa72d21fa556eec8d4d379a67602671d576d1b44c038370c10bf2c00b0d512d67753f4fee521edba1ee52c1a3fa0449141b67a0b4bc12995b9224bd297e2d6255ed4c724d94;
    5'b10111 : xpb = 1024'h47b676e63057a9c9b5e346bf216b0050ebe5408ea27fa69008661263a557a565505a5a3407c5598526024917521229be910e0fe5eb53225365725c7a16f8551c7d7a11aaab819a1f9ff019d3f7075bde073c9a1c9755881c98c906b3ccc40b13575b5b23a534ccfc3440beff5f369557c4b0ab2aa95f1969c7e3cd4a5d2c4c74;
    5'b11000 : xpb = 1024'h698e9e63490a77913a25c2d69504eb57793043eb3dfe2de2ba7aa2b9aa45a949b89768d0dd5a30a3bdcffe3aec7c5b004fba2dca06b8a11645caae4d00ceafe38c0796081f68ccdf196e5e311c5a6bb88b08732d3beb052be064a5f25a3827d48fdb1458f7a7f5fe643869e356cc75f376c7fac32e010955626544a76de64b54;
    5'b11001 : xpb = 1024'h8b66c5e061bd4558be683eee089ed65e067b4747d97cb5356c8f330faf33ad2e20d4776db2ef07c2559db35e86e68c420e664bae221e1fd92623001feaa50aaa9a951a65934fff9e92eca28e41ad7b930ed44c3de080823b28004530e7ac4495c85acd8e4a1b1f00943014c74e62568f28df4a5bb2a2f940fce6bc047ea04a34;
    5'b11010 : xpb = 1024'had3eed5d7a70132042aabb057c38c16493c64aa474fb3c881ea3c365b421b1128911860a8883dee0ed6b68822150bd83cd1269923d839e9c067b51f2d47b6571a9229ec30737325e0c6ae6eb67008b6d92a0254e8515ff4a6f9be46f7520615700da86c39c8e4802c427bfab45f8372adaf699f43744e92c976833618f5a4914;
    5'b11011 : xpb = 1024'h1e69cf84d134ac1efbe7bf45df786519af9b4ad03b02236352db9a66060d07eeee06172e93f23770e5dade5ed85cddfb27a45f9036364d1336346467837f4b874360ee71cb8d67d8734f28a5f377d717226704c69d254f4901aaf1b34869db860a52adcf3e3878776d5f83b045bdf19d3e340aaa6b9b7be7eb7a2fba1731e189;
    5'b11100 : xpb = 1024'h4041f701e9e779e6802a3b5d531250203ce64e2cd680aab604f02abc0afb0bd3564325cb69870e8f7da8938272c70f3ce6507d74519bcbd6168cb63a6d55a64e51ee72cf3f749a97eccd6d0318cae6f1a632ddd741bacc58494690f1d5ddf84742d2670490aba1799d572e943d53d238f04b5a42f03d6bd385fba71727ebe069;
    5'b11101 : xpb = 1024'h621a1e7f029a47ae046cb774c6ac3b26ca31518971ff3208b704bb120fe90fb7be8034683f1be5ae157648a60d31407ea4fc9b586d014a98f6e5080d572c0115607bf72cb35bcd57664bb1603e1df6cc29feb6e7e650496790e23030635215087b522039e31eca7bcd4ed97834e9b2d4a262a9db74df5bbf207d1e7438a5df49;
    5'b11110 : xpb = 1024'h83f245fc1b4d157588af338c3a46262d577c54e60d7db95b69194b6814d7139c26bd430514b0bcccad43fdc9a79b71c063a8b93c8866c95bd73d59e041025bdc6f097b8a27430016dfc9f5bd637106a6adca8ff88ae5c676d87dcf6ef0c631c9b3d1d96f3591f37dfd46845c2c7f93705479f973f9814baabafe95d1495fde29;
    5'b11111 : xpb = 1024'ha5ca6d7933ffe33d0cf1afa3ade01133e4c75842a8fc40ae1b2ddbbe19c517808efa51a1ea4593eb4511b2ed4205a3022254d720a3cc481eb795abb32ad8b6a37d96ffe79b2a32d659483a1a88c41681319669092f7b438620196ead7e3a4e8aec5192a488051c802d3e2f402415740c0691490c7e233b9655800d2e5a19dd09;
    endcase
end

endmodule

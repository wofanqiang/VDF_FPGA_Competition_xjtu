module xpb_5_365
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h88368672c0766d92396d9172dd51a23f9711ea5a42a982d30b9652e8bec0c3b4a47f986cc1414fa6bb8f8f4ea93604e4eabc979ead6f09a7eef40820a305201e4a18b197fae8c5222d752199ce226b112169ea191e39ac6438bca5b3c1846b0e1c903cede3c00e685457ca0af1d40e591b1340fc3bbdc8205195f8fc0df99e7e;
    5'b00010 : xpb = 1024'h5fbfc78fbefea65ba7d5ab0eaa48fd2dbcadd183afdb652e994fec7bca7eda6145b6b360b85c20bed7c0df566f0df8ff715f0757382b43042d48d0e30b37cb8b1fe22e8146408cff48504091036911f14eceda99afed2bb7bbecb96cc8de338a0a18e7b216b7244321efad36ebd7f688e74ca316273033105cbc76f39310d691;
    5'b00011 : xpb = 1024'h374908acbd86df25163dc4aa7740581be249b8ad1d0d478a2709860ed63cf10de6edce54af76f1d6f3f22f5e34e5ed19f801770fc2e77c606b9d99a5736a76f7f5abab6a919854dc632b5f8838afb8d17c33cb1a41a0ab0b3f1ccd25d037fc05f7a1927649ae3a1def879062e5dbdeb8b386053012a29e0067e2f4eb18280ea4;
    5'b00100 : xpb = 1024'hed249c9bc0f17ee84a5de464437b30a07e59fd68a3f29e5b4c31fa1e1fb07ba8824e948a691c2ef10237f65fabde1347ea3e6c84da3b5bca9f26267db9d2264cb752853dcf01cb97e067e7f6df65fb1a998bb9ad3542a5ec24ce0ded791c481e52a3d3a7ca54ff8bd1f738edfdfc6e87fbf6749fe1508f0730972e29d3f46b7;
    5'b00101 : xpb = 1024'h9708d03c7c858580be136fb9218955499ef78a30cce8acb8c059728aa0bbcb6f2ca481b567d31295cbb30eb4a3f3e61969607e66fb12bf6498e66a887ea24283158dd9ebd7d8e1dbab7ba0193c18cac2cb02a5b3f18dd6c2fb09869299162f9001ba7a2860655e6111773d99d1b3d5419ad2a84639d2d110c49f6bdeab38e535;
    5'b00110 : xpb = 1024'h6e9211597b0dbe4a2c7b8954ee80b037c493715a3a1a8f144e130c1dac79e21bcddb9ca95eede3ade7e45ebc69cbda33f002ee1f85cef8c0d73b334ae6d4edefeb5756d52330a9b8c656bf10715f71a2f8679634834156167e399a4ba06ff80bef4324ec935c743bdf0f20c5cbb7bd71670c0a6025453c00cfc5e9d630501d48;
    5'b00111 : xpb = 1024'h461b52767995f7139ae3a2f0bb780b25ea2f5883a74c716fdbcca5b0b837f8c86f12b79d5608b4c60415aec42fa3ce4e76a55dd8108b321d158ffc0d4f07995cc120d3be6e887195e131de07a6a6188325cc86b514f4d56a0169ae04a7c9c087dccbcfb0c6538a16aca703f1c5bba5a133456c7a10b7a6f0daec67cdb567555b;
    5'b01000 : xpb = 1024'h1da49393781e2fdd094bbc8c886f66140fcb3fad147e53cb69863f43c3f60f751049d2914d2385de2046fecbf57bc268fd47cd909b476b7953e4c4cfb73a44c996ea50a7b9e03972fc0cfcfedbecbf6353317735a6a854bd8499c1bdaf238903ca547a74f94a9ff17a3ee71dbfbf8dd0ff7ece93fc2a11e0e612e5c53a7e8d6e;
    5'b01001 : xpb = 1024'ha5db1a0638949d6f42b94dff65c10853a6dd2a075727d69e751c922c82b6d329b4c96afe0e64d584dbd68e1a9eb1c74de804652f48b6752142d8ccf05a3f64e7e103023fb4c8fe9529821e98aa0f2a74749b614ec4e20121bd56677170a7f411e6e4b762dd0aae59ce96b128b1939c2a1a920f9037e7da0137a8dec148782bec;
    5'b01010 : xpb = 1024'h7d645b23371cd638b121679b32b86341cc791130c459b8fa02d62bbf8e74e9d6560085f2057fa69cf807de226489bb686ea6d4e7d372ae7d812d95b2c2721054b6cc7f290020c672445d3d8fdf55d154a20051cf5695807540867b2a7801bc8dd46d62271001c4349c2e9454ab978459e6cb71aa235a44f142cf5cb8cd8f63ff;
    5'b01011 : xpb = 1024'h54ed9c4035a50f021f898136ffafbe2ff214f85a318b9b55908fc5529a330082f737a0e5fc9a77b514392e2a2a61af82f54944a05e2ee7d9bf825e752aa4bbc18c95fc124b788e4f5f385c87149c7834cf65424fe848ffc8c3b68ee37f5b8509c1f60ceb42f8da0f69c67780a59b6c89b304d3c40eccafe14df5dab052a69c12;
    5'b01100 : xpb = 1024'h2c76dd5d342d47cb8df19ad2cca7191e17b0df839ebd7db11e495ee5a5f1172f986ebbd9f3b548cd306a7e31f039a39d7bebb458e8eb2135fdd7273792d7672e625f78fb96d0562c7a137b7e49e31f14fcca32d079fc7f1c46e6a29c86b54d85af7eb7af75efefea375e5aac9f9f54b97f3e35ddfa3f1ad1591c58a7d7bdd425;
    5'b01101 : xpb = 1024'h4001e7a32b58094fc59b46e999e740c3d4cc6ad0bef600cac02f878b1af2ddc39a5d6cdead019e54c9bce39b61197b8028e241173a75a923c2beff9fb0a129b3828f5e4e2281e0994ee9a757f29c5f52a2f23510baffe6fca16b6558e0f16019d076273a8e705c504f63dd899a33ce94b7797f7e5b185c16442d69f5cd50c38;
    5'b01110 : xpb = 1024'h8c36a4ecf32bee2735c745e176f0164bd45eb1074e98e2dfb7994b61706ff190de256f3aac11698c082b5d885f479c9ced4abbb02116643a2b1ff81a9e0f32b98241a77cdd10e32bc263bc0f4d4c31064b990d6a29e9aad402d35c094f93810fb9979f618ca7142d594e07e38b774b42668ad8f4216f4de1b5d8cf9b6aceaab6;
    5'b01111 : xpb = 1024'h63bfe609f1b426f0a42f5f7d43e77139f9fa9830bbcac53b4552e4f47c2e083d7f5c8a2ea32c3aa4245cad90251f90b773ed2b68abd29d966974c0dd0641de26580b24662868ab08dd3edb068292d7e678fdfdeabb9d2a2786036fc256ed498ba7204a25bf9e2a0826e5eb0f857b337232c43b0e0ce1b8d1c0ff4d92efe5e2c9;
    5'b10000 : xpb = 1024'h3b492726f03c5fba1297791910decc281f967f5a28fca796d30c7e8787ec1eea2093a5229a470bbc408dfd97eaf784d1fa8f9b21368ed6f2a7c9899f6e7489932dd4a14f73c072e5f819f9fdb7d97ec6a662ee6b4d50a97b0933837b5e47120794a8f4e9f2953fe2f47dce3b7f7f1ba1fefd9d27f85423c1cc25cb8a74fd1adc;
    5'b10001 : xpb = 1024'h12d26843eec4988380ff92b4ddd6271645326683962e89f260c6181a93aa3596c1cac0169161dcd45cbf4d9fb0cf78ec81320ad9c14b104ee61e5261d6a73500039e1e38bf183ac312f518f4ed2025a6d3c7deebdf0428ce8c63973465a0da8382319fae258c55bdc215b167798303d1cb36ff41e3c68eb1d74c4981fa1452ef;
    5'b10010 : xpb = 1024'h9b08eeb6af3b0615ba6d2427bb27c955dc4450ddd8d80cc56c5c6b03526af94b664a588352a32c7b184edcee5a057dd16beea2786eba19f6d5125a8279ac551e4db6cfd0ba00ffe5406a3a8ebb4290b7f531c904fd3dd532c5203ce8272545919ec1dc9c094c6426166d7b726b57122ae64a403e1f8456d228e2427e080df16d;
    5'b10011 : xpb = 1024'h72922fd3adc33edf28d53dc3881f244401e038074609ef20fa1604965e290ff80781737749bdfd9334802cf61fdd71ebf2911230f976535313672344e1df008b23804cba0558c7c25b455985f08937982296b9858ef15486485050a12e7f0e0d8c4a87603c437a00e4055e9e655afa5ab283a2580af6c1c23408c0758d252980;
    5'b10100 : xpb = 1024'h4a1b70f0ac4b77a8973d575f55167f32277c1f30b33bd17c87cf9e2969e726a4a8b88e6b40d8ceab50b17cfde5b56606793381e984328caf51bbec074a11abf7f949c9a350b08f9f7620787d25cfde784ffbaa0620a4d3d9cb80645a35d8d68979d332246f3a8fdbb19d41ca5f5ee28a7ebd0471f6692cb23f2f3e6d123c6193;
    5'b10101 : xpb = 1024'h21a4b20daad3b07205a570fb220dda204d18065a206db3d8158937bc75a53d5149efa95f37f39fc36ce2cd05ab8d5a20ffd5f1a20eeec60b9010b4c9b2445764cf13468c9c08577c90fb97745b1685587d609a86b258532d4eb078133d329f05675bdce8a231a5b67f3524f65962caba4af6668be1db97a24a55bc64975399a6;
    5'b10110 : xpb = 1024'ha9db38806b4a1e043f13026dff5f7c5fe429f0b4631736ab211f8aa534660105ee6f41cbf934ef6a28725c5454c35f05ea928940bc5dcfb37f04bcea55497783192bf82496f11c9ebe70b90e2938f0699eca849fd091ff91876d1dc6feb70a1383ec19d685f1b41ed38cef014b36d9136609a7881d995fc29bebb560a54d3824;
    5'b10111 : xpb = 1024'h8164799d69d256cdad7b1c09cc56d74e09c5d7ddd0491906aed92438402417b28fa65cbff04fc08244a3ac5c1a9b53207134f8f9471a090fbd5985acbd7c22efeef5750de248e47bd94bd8055e7f9749cc2f752062457ee50a9d31800610d28f7174c49ab8e8c9f9a124d22d453ac143324309a2090bcab2a71233582a647037;
    5'b11000 : xpb = 1024'h58edbaba685a8f971be335a5994e323c2f61bf073d7afb623c92bdcb4be22e5f30dd77b3e76a919a60d4fc63e073473af7d768b1d1d6426bfbae4e6f25aece5cc4bef1f72da0ac58f426f6fc93c63e29f99465a0f3f8fe388dcd45390d6a9b0b5efd6f5eebdfdfd46ebcb5593f3ea972fe7c6bbbf47e35a2b238b14faf7ba84a;
    5'b11001 : xpb = 1024'h3076fbd766e2c8608a4b4f4166458d2a54fda630aaacddbdca4c575e57a0450bd21492a7de8562b27d064c6ba64b3b557e79d86a5c927bc83a0317318de179c99a886ee078f874360f0215f3c90ce50a26f9562185ac7d8c10fd58f214c463874c861a231ed6f5af3c549885394291a2cab5cdd5dff0a092bd5f2f473492e05d;
    5'b11010 : xpb = 1024'h8003cf4656b0129f8b368dd333ce8187a998d5a17dec0195805f0f1635e5bb8734bad9bd5a033ca99379c736c232f70051c4822e74eb5247857dff3f61425367051ebc9c4503c1329dd34eafe538bea545e46a2175ffcdf942d6cab1c1e2c033a0ec4e751ce0b8a09ec7bb1334679d296ef2fefcb630b82c885ad3eb9aa1870;
    5'b11011 : xpb = 1024'h9036c36725e16ebc3220fa50108e8a5811ab77b45a8842ec639c43da221f1f6d17cb460896e1837154c72bc215593454efd8dfc194bdbecc674be81499194554ba6a9d61bf39013557525684cc75f6fb75c830bb3599a943ccea125edda29711569f01d5358e19f25e4445bc251a882bb20270ec0720d3a31a1ba63ac7a3b6ee;
    5'b11100 : xpb = 1024'h67c004842469a785a08913ebdd85e54637475eddc7ba2547f155dd6d2ddd3619b90260fc8dfc548970f87bc9db31286f767b4f7a1f79f828a5a0b0d7014bf0c190341a4b0a90c912722d757c01bc9ddba32d213bc74d2897501a2617e4fc5f8d4427ac9968852fcd2bdc28e81f1e705b7e3bd305f2933e93254224324cbaef01;
    5'b11101 : xpb = 1024'h3f4945a122f1e04f0ef12d87aa7d40345ce3460734ec07a37f0f7700399b4cc65a397bf0851725a18d29cbd1a1091c89fd1dbf32aa363184e3f57999697e9c2e65fd973455e890ef8d089473370344bbd09211bc5900a7ead34a39d0ec56280931b0575d9b7c45a7f9740c141922588b4a75351fde05a9833068a229d1d22714;
    5'b11110 : xpb = 1024'h16d286be217a19187d59472377749b22827f2d30a21de9ff0cc9109345596372fb7096e47c31f6b9a95b1bd966e110a483c02eeb34f26ae1224a425bd1b1479b3bc7141da14058cca7e3b36a6c49eb9bfdf7023ceab4273e567a4d89f3aff0851f390221ce735b82c70bef40132640bb16ae9739c97814733b8f202156e95f27;
    5'b11111 : xpb = 1024'h9f090d30e1f086aab6c6d89654c63d621991178ae4c76cd2185f637c041a27279ff02f513d73466064eaab28101715896e7cc689e2617489113e4a7c74b667b985dfc5b59c291deed558d5043a6c56ad1f60ec5608edd3a28f36f33db5345b933bc93f0fb23369eb1b63b94b04fa4f1431c1d8360535dc938d25191d64e2fda5;
    endcase
end

endmodule

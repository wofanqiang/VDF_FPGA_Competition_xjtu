module xpb_5_985
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h62dd739c4df85c98ec59bd932d9b182b0929e2a3e72eb3c9f5c7d8b3f8faa8f9c3c37ff092a4cdbe6d41e77cc4830f0bf80f904bbdf3c7fc44e09e403343bd21d5924142571fdec4219e0c72a86b5e7342870ff7a200cd2f45291c31700b9a007267d7a312cd2a8539b177156a901a2225138eb4e48bef6159968c1bab0511c7;
    5'b00010 : xpb = 1024'h150da1e2da0284690dae034f4adbe904a0ddc216f8e5c71c6db2f8123ef2a4eb843e82685b231cee3b258fb2a5a80d4d8c04f8b15934bfacd921fd222bb5059236d54dd5feaec04330a21642b7faf8b591092656b77b6d4dd4c5a66825ec916eb5c81d1c74d15c7ceca3074bdd500e1afb4d3e8778cc81926cbd9d32cd27bd23;
    5'b00011 : xpb = 1024'h77eb157f27fae101fa07c0e27877012faa07a4bae0147ae6637ad0c637ed4de548020258edc7eaaca867772f6a2b1c59841488fd172887a91e029b625ef8c2b40c678f1855ce9f07524022b560665728d390364e597c3a7d19eec29995f82b6f282ff4bf879e870226547e6147e0283d2060cd3c5d5870f3c654294e782cceea;
    5'b00100 : xpb = 1024'h2a1b43c5b40508d21b5c069e95b7d20941bb842df1cb8e38db65f0247de549d7087d04d0b64639dc764b1f654b501a9b1809f162b2697f59b243fa44576a0b246daa9babfd5d808661442c856ff5f16b22124cad6ef6da9ba98b4cd04bd922dd6b903a38e9a2b8f9d9460e97baa01c35f69a7d0ef1990324d97b3a659a4f7a46;
    5'b00101 : xpb = 1024'h8cf8b76201fd656b07b5c431c352ea344ae566d1d8fa4202d12dc8d876dff2d0cc4084c148eb079ae38d06e20fd329a7101981ae705d4755f72498848aadc846433cdcee547d5f4a82e238f818614fde64995ca510f7a7caeeb46901bbe4bcddddf811dbfc6fe37f12f785ad253036581bae0bc3d624f2863311c68145548c0d;
    5'b00110 : xpb = 1024'h3f28e5a88e078d3b290a09ede093bb0de2994644eab155554918e836bcd7eec28cbb8739116956cab170af17f0f827e8a40eea140b9e3f068b65f766831f10b6a47fe981fc0c40c991e642c827f0ea20b31b7304267247e97e50f33871c5b44c215857555e741576c5e915e397f02a50f1e7bb966a6584b74638d79867773769;
    5'b00111 : xpb = 1024'ha2065944dbffe9d41563c7810e2ed338ebc328e8d1e0091f3ee0c0eab5d297bc507f0729a40e24891eb29694b57b36f49c1e7a5fc9920702d04695a6b662cdd87a122ac4532c1f8db3844f3ad05c4893f5a282fbc8731518c37a0f69e1d14e4c93c02ef871413ffbff9a8cf90280447316fb4a4b4ef174189fcf63b4127c4930;
    5'b01000 : xpb = 1024'h5436878b680a11a436b80d3d2b6fa4128377085be3971c71b6cbe048fbca93ae10fa09a16c8c73b8ec963eca96a035363013e2c564d2feb36487f488aed41648db553757fabb010cc288590adfebe2d64424995addedb537531699a097b245bad7207471d34571f3b28c1d2f7540386bed34fa1de3320649b2f674cb349ef48c;
    5'b01001 : xpb = 1024'h666b5d1f4143974580c52f948b074ec1b2ae7cef54e2fc42eb6ffa741c28f9fd1750c19350ac2e8ba79e70077c53377c4094b2b0013f663f8c9536aa7455eb93c9843eba249e28bd18c62daef7b7d1892a6afb9f3685555e2b323d74d933d291a80b9eb3549a3eb657dad65e8002c64c36ea9f07772987ac61d85e256c19fe8;
    5'b01010 : xpb = 1024'h6944296e420c960d4466108c764b8d172454ca72dc7ce38e247ed85b3abd389995388c09c7af90a727bbce7d3c484283bc18db76be07be603da9f1aada891bdb122a852df969c14ff32a6f4d97e6db8bd52dbfb19569228527dc4008bd9ed7298ce8918e4816ce709f2f247b52904686e88238a55bfe87dc1fb411fe01c6b1af;
    5'b01011 : xpb = 1024'h1b7457b4ce16bddd65ba5648938c5df0bc08a9e5ee33f6e09c69f7b980b5348b55b38e81902ddfd6f59f76b31d6d40c5500e43dc5948b610d1eb508cd2fa644b736d91c1a0f8a2cf022e791da77675ce23afd610aae3c2a3b778ca3f737fce97d048d707aa1b00685220b4b1c5503a7fbebbe877f03f1a0d32db231523e95d0b;
    5'b01100 : xpb = 1024'h7e51cb511c0f1a76521413dbc127761bc5328c89d562aaaa9231d06d79afdd8519770e7222d2ad9562e15e2fe1f04fd1481dd428173c7e0d16cbeecd063e216d48ffd303f818819323cc85904fe1d4416636e6084ce48fd2fca1e670e38b689842b0aeaabce82aed8bd22bc72fe054a1e3cf772cd4cb096e8c71af30ceee6ed2;
    5'b01101 : xpb = 1024'h3081f997a819424673685997de6846f55ce66bfce719bdfd0a1cefcbbfa7d976d9f210e9eb50fcc530c50665c3154e12dc133c8db27d75bdab0d4daefeaf69ddaa42df979fa7631232d08f605f716e83b4b8fc67625f2ff18c3e70a7996c60068610f4241eec5ce53ec3bbfda2a0489aba0926ff690b9b9f9f98c047f1111a2e;
    5'b01110 : xpb = 1024'h935f6d33f6119edf5fc2172b0c035f2066104ea0ce4871c6ffe4c87fb8a282709db590da7df5ca839e06ede287985d1ed422ccd970713db9efedebef31f326ff7fd520d9f6c741d6546e9bd307dcccf6f7400c5f045ffd20d1678cd90977fa06f878cbc731b9876a787533130d3062bcdf1cb5b44d978b00f92f4c639c162bf5;
    5'b01111 : xpb = 1024'h458f9b7a821bc6af81165ce729442ff9fdc42e13dfff851977cfe7ddfe9a7e625e309352467419b36bea961868bd5b606818353f0bb2356a842f4ad12a646f6fe1182d6d9e5623556372a5a3176c673945c222be19da9d3f6104170fbf58f1753bd9114093bdb9622b66c3497ff056b5b5566586e1d81d320c565d7abe38d751;
    5'b10000 : xpb = 1024'ha86d0f16d01423486d701a7a56df482506ee10b7c72e38e36d97c091f795275c21f41342d918e771d92c7d952d406a6c6027c58ac9a5fd66c90fe9115da82c91b6aa6eaff57602198510b215bfd7c5ac884932b5bbdb6a6ea62d33412f648b75ae40e8e3a68ae3e765183a5eea8070d7da69f43bc6640c9365ece996693de918;
    5'b10001 : xpb = 1024'h5a9d3d5d5c1e4b188ec46036742018fe9ea1f02ad8e54c35e582dff03d8d234de26f15baa19736a1a71025cb0e6568adf41d2df064e6f5175d5147f35619750217ed7b439d04e3989414bbe5cf675feed6cb4914d1560a8d35c9bd77e54582e3f1a12e5d088f15df1809ca955d4064d0b0a3a40e5aa49ec47913faad8b609474;
    5'b10010 : xpb = 1024'hccd6ba3e82872e8b018a5f29160e9d83655cf9dea9c5f885d6dff4e83851f3fa2ea18326a1585d174f3ce00ef8a66ef881296560027ecc7f192a6d54e8abd72793087d74493c517a318c5b5def6fa31254d5f73e6d0aaabc56647ae9b267a52350173d66a9347d6cafb5acbd00058c986dd53e0eee530f58c3b0bc4ad833fd0;
    5'b10011 : xpb = 1024'h6faadf403620cf819c726385befc02033f7fb241d1cb13525335d8027c7fc83966ad9822fcba538fe235b57db40d75fb802226a1be1bb4c43673451581ce7a944ec2c9199bb3a3dbc4b6d228876258a467d46f6b88d177db0a8f63e00b321452a7694b797d60725c04acd1e13a9072ebabf0e295d3712056e5d197e058885197;
    5'b10100 : xpb = 1024'h21db0d86c22af751bdc6a941dc3cd2dcd73391b4e38226a4cb20f760c277c42b27289a9ac538a2bfb0195db39532743d14178f07595cac74cab4a3f77a3fc304b005d5ad4342855ad3badbf896f1f2e6b65685ca9e4c17f99a2bee16c1130bc0eac990f2df64a453b79e6217ad5066e4822a926867b1b287f8f8a8f77aaafcf3;
    5'b10101 : xpb = 1024'h84b88123102353eaaa2066d509d7eb07e05d7458cab0da6ec0e8d014bb726d24eaec1a8b57dd707e1d5b453059b583490c271f53175074710f954237ad838026859816ef9a62641ef558e86b3f5d5159f8dd95c2404ce528df550a48311ea5c15d316895f231ced8f14fd92d17e08106a73e211d4c3da1e9528f351325b00eba;
    5'b10110 : xpb = 1024'h36e8af699c2d7bbacb74ac912718bbe1781153cbdc67edc138d3ef73016a6916ab671d03205bbfadeb3eed663ada818aa01c87b8b2916c21a3d6a119a5f4c896e6db238341f1459e045cf23b4eeceb9c475fac2155c785476ef1947ee6ff9d2fa091ae0f543600d0a44169638aa074ff7d77d0efe07e341a65b6462a47d2ba16;
    5'b10111 : xpb = 1024'h99c62305ea25d853b7ce6a2454b3d40c813b366fc396a18b2e9bc826fa6512106f2a9cf3b3008d6c5880d4e2ff5d9096982c18047085341de8b73f59d93885b8bc6d64c59911246225fafeadf7584a0f89e6bc18f7c85276b41ab0b0570b373012f985b267032b55ddf2e078f5308f21a28b5fa4c50a237bbf4cd245f2d7cbdd;
    5'b11000 : xpb = 1024'h4bf6514c76300023d922afe071f4a4e618ef15e2d54db4dda686e785405d0e022fa59f6b7b7edc9c26647d18e0828ed82c21806a0bc62bce7cf89e3bd1a9ce291db0715940a005e134ff087e06e7e451d868d2780d42f29543b73ae70cec2e9e5659cb2bc9075d4d90e470af67f0831a78c50f77594ab5acd273e35d14fa7739;
    5'b11001 : xpb = 1024'haed3c4e8c4285cbcc57c6d739f8fbd112218f886bc7c68a79c4ec0393957b6fbf3691f5c0e23aa5a93a66495a5059de4243110b5c9b9f3cac1d93c7c04ed8b4af342b29b97bfe4a5569d14f0af5342c51aefe26faf43bfc488e057187cf7c89ec8c1a2cedbd487d2ca95e7c4d2809d3c9dd89e2c3dd6a50e2c0a6f78bfff8900;
    5'b11010 : xpb = 1024'h6103f32f5032848ce6d0b32fbcd08deab9ccd7f9ce337bfa1439df977f4fb2edb3e421d3d6a1f98a618a0ccb862a9c25b826791b64faeb7b561a9b5dfd5ed3bb5485bf2f3f4ec62465a11ec0bee2dd076971f8cec4be5fe3187ce14f32d8c00d0c21e8483dd8b9ca7d8777fb4540913574124dfed217373f3f31808fe222345c;
    5'b11011 : xpb = 1024'h13342175dc3cac5d0824f8ebda115ec45180b76cdfea8f4c8c24fef5c547aedf745f244b9f2048ba2f6db501674f9a674c1be181003be32bea5bfa3ff5d01c2bb5c8cbc2e6dda7a374a52890ce727749b7f40f2dda390001a8196b85e8b9b77b4f822dc19fdcebc230790831b800852e4a4bfdd16657c970525891a70444dfb8;
    5'b11100 : xpb = 1024'h761195122a3508f5f47eb67f07ac76ef5aaa9a10c719431681ecd7a9be4257d93822a43c31c516789caf9c7e2bd2a973442b71ccbe2fab282f3c98802913d94d8b5b0d053dfd86679643350376ddd5bcfa7b1f257c39cd30ed4287b758c5517bc1ea0564b2aa16476a2a7f4722909f506f5f8c864ae3b8d1abef1dc2af49f17f;
    5'b11101 : xpb = 1024'h2841c358b63f30c615d2fc3b24ed47c8f25e7983d8d05668f9d7f708043a53caf89da6b3fa4365a86a9344b40cf7a7b4d820da325970a2d8c37df762218521bdec9e1998e58c67e6a5473ed3866d6fff48fd358491b46d4f7cdf11ee0ea648ea054a4ade14ae483f1d1c0f7d9550934945993c58df244b02bf162ed9d16c9cdb;
    5'b11110 : xpb = 1024'h8b1f36f504378d5f022cb9ce52885ff3fb885c27bfff0a32ef9fcfbbfd34fcc4bc6126a48ce83366d7d52c30d17ab6c0d0306a7e17646ad5085e95a254c8dedfc2305adb3cac46aac6e54b462ed8ce728b84457c33b53a7ec2082e1f7eb1e2ea77b22281277b72c456cd8692ffe0ad6b6aaccb0dc3b03a6418acbaf57c71aea2;
    5'b11111 : xpb = 1024'h3d4f653b9041b52f2380ff8a6fc930cd933c3b9ad1b61d85678aef1a432cf8b67cdc291c55668296a5b8d466b29fb5026425d2e3b2a562859c9ff4844d3a27502373676ee43b2829d5e955163e6868b4da065bdb492fda9d51a4b8563492da58bb1267fa897fa4bc09bf16c972a0a16440e67ae057f0cc952bd3cc0c9e9459fe;
    endcase
end

endmodule

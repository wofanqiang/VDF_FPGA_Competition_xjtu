module xpb_5_795
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h7bbba979ed2fb95be110728eed4bb9d2247987a44fae54ded81a3042dab66981286e8ea5f50a1ae96a530dad66e38c10ff0734467bd46d36a49408afdbe6aa84d78877a38be17a7346f21ffcfc1a4ec749b09728b083d24a97280b5b4ca19529713c3846105f09a7f7ff724cec959666cfb5193ebea6bda365433dc8705bea1f;
    5'b00010 : xpb = 1024'h46ca0d9e18713deef71b6d46ca3d2c52d77d0c17c9e509463257a730026a25fa4d949fd31fedb7443547dc13ea69075799f440a6d4f60a219888d2017cfae0583ac1ba986831f7a17b4a3d575f58d95d9f5c34b8d481778478c384bbdf1887c0b370de626ff51ac2693efdbae15b06a45090539b2d021e168417008c57d56dd3;
    5'b00011 : xpb = 1024'h11d871c243b2c2820d2667fea72e9ed38a80908b441bbdad8c951e1d2a1de27372bab1004ad1539f003caa7a6dee829e34e14d072e17a70c8c7d9b531e0f162b9dfafd8d448274cfafa25ab1c29763f3f507d248f87f1cbe5a5efe1c718f7a57f5a5847ecf8b2bdcda7e8928d62076e1d16b8df79b5d7e89a2eac3503f4ef187;
    5'b00100 : xpb = 1024'h8d941b3c30e27bddee36da8d947a58a5aefa182f93ca128c64af4e6004d44bf49b293fa63fdb6e886a8fb827d4d20eaf33e8814da9ec14433111a402f9f5c0b075837530d063ef42f6947aaebeb1b2bb3eb86971a902ef08f1870977be310f8166e1bcc4dfea3584d27dfb75c2b60d48a120a7365a043c2d082e0118afaadba6;
    5'b00101 : xpb = 1024'h58a27f605c2400710441d545716bcb2661fd9ca30e00c6f3beecc54d2c88086dc04f50d36abf0ae33584868e585789f5ced58dae030db12e25066d549b09f683d8bcb825acb46c712aec980921f03d5194640701cd009442d32282d850a80218a91662e13f80469f43bd86e3b77b7d8621fbe192c85f9ca02701c3dc97245f5a;
    5'b00110 : xpb = 1024'h23b0e384876585041a4ccffd4e5d3da71501211688377b5b192a3c3a543bc4e6e575620095a2a73e007954f4dbdd053c69c29a0e5c2f4e1918fb36a63c1e2c573bf5fb1a8904e99f5f44b563852ec7e7ea0fa491f0fe397cb4bdfc38e31ef4afeb4b08fd9f1657b9b4fd1251ac40edc3a2d71bef36bafd1345d586a07e9de30e;
    5'b00111 : xpb = 1024'h9f6c8cfe74953e5ffb5d428c3ba8f779397aa8bad7e5d039f1446c7d2ef22e680de3f0a68aacc2276acc62a242c0914d68c9ce54d803bb4fbd8f3f561804d6dc137e72be14e66412a636d560814916af33c03bbaa1820bc74be607942fc089d95c874143af756161acfc849e98d6842a728c352df561bab6ab18c468eef9cd2d;
    5'b01000 : xpb = 1024'h6a7af1229fd6c2f311683d44189a69f9ec7e2d2e521c84a14b81e36a56a5eae1330a01d3b5905e8235c13108c6460c9403b6dab53125583ab18408a7b9190caf76b7b5b2f136e140da8ef2bae487a145896bd94ac57fb1012d8180f4c2377c709ebbe7600f0b727c1e3c100c8d9bf467f3676f8a63bd1b29c9ec872cd67350e1;
    5'b01001 : xpb = 1024'h35895546cb184786277337fbf58bdc7a9f81b1a1cc533908a5bf5a577e59a75a58301300e073fadd00b5ff6f49cb87da9ea3e7158a46f525a578d1f95a2d4282d9f0f8a7cd875e6f0ee7101547c62bdbdf1776dae97d563b0f1cfa5554ae6f07e0f08d7c6ea183968f7b9b7a826164a57442a9e6d2187b9ce8c049f0bdecd495;
    5'b01010 : xpb = 1024'h97b96af659cc193d7e32b3d27d4efb528536154689ed6ffffcd144a60d63d37d56242e0b579737cbaacdd5cd5103213990f375e3689210996d9b4afb4178563d2a3b9ca9d7db9d433f2d6fab04b67234c3146b0d7afb74f0b873b5e725619f23253398ce3794b100bb26e87726d4e2f51de4434073dc1007940cb4a5665849;
    5'b01011 : xpb = 1024'h7c5362e4e38985751e8ea542bfc908cd76febdb99638424ed817018780c3cd54a5c4b2d40061b22135fddb8334348f32389827bc5f3cff473e01a3fad72822db14b2b34035b956108a314d6ca71f05397e73ab93bdfecdbf87e07f1133c6f6c894616bdede969e58f8ba993563bc6b49c4d2fd81ff1a99b36cd74a7d15c24268;
    5'b01100 : xpb = 1024'h4761c7090ecb0a0834999ffa9cba7b4e2a02422d106ef6b632547874a87789cdcaeac4012b454e7c00f2a9e9b7ba0a78d385341cb85e9c3231f66d4c783c58ae77ebf6351209d33ebe896ac70a5d8fcfd41f4923e1fc72f9697bf871c63de95fd69611fb3e2caf7369fa24a35881db8745ae37de6d75fa268bab0d40fd3bc61c;
    5'b01101 : xpb = 1024'h12702b2d3a0c8e9b4aa49ab279abedcedd05c6a08aa5ab1d8c91ef61d02b4646f010d52e5628ead6cbe778503b3f85bf6e72407d1180391d25eb369e19508e81db253929ee5a506cf2e188216d9c1a6629cae6b405fa18334b1771d258b4dbf718cab8179dc2c08ddb39b0114d474bc4c689723adbd15a99aa7ed004e4b549d0;
    5'b01110 : xpb = 1024'h8e2bd4a7273c47f72bb50d4166f7a7a1017f4e44da53fffc64ac1fa4aae1afc8187f63d44b3305c0363a85fda22311d06d7974c38d54a653ca7f3f4df5373906b2adb0cd7a3bcae039d3a81e69b6692d737b7ddcb67dea7de23f7d2da55671208a06f05dae21ca35d339225e39dce22b963e8b799a78183d0fc20dcd551133ef;
    5'b01111 : xpb = 1024'h593a38cb527dcc8a41c007f943e91a21b482d2b8548ab463bee99691d2956c413da575017616a21b012f546425a88d1708668123e676433ebe74089f964b6eda15e6f3c2568c480e6e2bc578ccf4f3c3c9271b6cda7b8fb7c3daf68e37cd63b7cc3b967a0db7db504478adcc2ea252691719c5d608d378b02e95d0913c8ab7a3;
    5'b10000 : xpb = 1024'h24489cef7dbf511d57cb02b120da8ca26786572bcec168cb19270d7efa4928ba62cb862ea0fa3e75cc2422caa92e085da3538d843f97e029b268d1f1375fa4ad792036b732dcc53ca283e2d330337e5a1ed2b8fcfe7934f1a5766feeca44564f0e703c966d4dec6ab5b8393a2367c2a697f50032772ed9234d69935524043b57;
    5'b10001 : xpb = 1024'ha00446696aef0a7938db75400e2646748bffded01e6fbda9f1413dc1d4ff923b8b3a14d49604595f367730781011946ea25ac1cabb6c4d6056fcdaa113464f3250a8ae5abebe3fafe97602d02c4dcd2168835025aefd073c3c9e7b4a16e5eb787fac74dc7dacf612adb7ab870ffd590d67aa197135d596c6b2acd11d94602576;
    5'b10010 : xpb = 1024'h6b12aa8d96308f0c4ee66ff7eb17b8f53f03634398a672114b7eb4aefcb34eb4b0602601c0e7f5ba016bfede93970fb53d47ce2b148dea4b4af1a3f2b45a8505b3e1f14f9b0ebcde1dce202a8f8c57b7be2eedb5d2faac761e39f4aaa95cde0fc1e11af8dd43072d1ef736f504c2c94ae88553cda430f739d18093e17bd9a92a;
    5'b10011 : xpb = 1024'h36210eb1c172139f64f16aafc8092b75f206e7b712dd2678a5bc2b9c24670b2dd586372eebcb9214cc60cd45171c8afbd834da8b6daf87363ee66d44556ebad9171b3444775f3a0c52263d84f2cae24e13da8b45f6f851afffd56e0b3bd3d0a70415c1153cd918479036c262f988398869608e2a128c57acf05456a563532cde;
    5'b10100 : xpb = 1024'h12f72d5ecb398327afc6567a4fa9df6a50a6c2a8d13dadffff9a2894c1ac7a6faac485c16af2e6f97559bab9aa206427321e6ebc6d1242132db3695f682f0ac7a54773953afb73a867e5adf56096ce4698628d61af5f6e9e170e76bce4ac33e464a67319c6f296201764dd0ee4da9c5ea3bc88680e7b8200f2819694accb092;
    5'b10101 : xpb = 1024'h7ceb1c4fd9e3518e5c0cd7f6924657c8c983f3cedcc22fbed813d2cc26d13128231ad7020bb9495901a8a9590185925372291b3242a59157d76f3f45d2699b3151dceedcdf9131adcd707adc5223bbabb336bffecb79c9347898f2c71aec5867b7869f77acce3309f975c01ddae3402cb9f0e1c53f8e75c3746b5731bb289ab1;
    5'b10110 : xpb = 1024'h47f980740524d6217217d2ae6f37ca497c87784256f8e426325149b94e84eda14840e82f369ce5b3cc9d77bf850b0d9a0d1627929bc72e42cb640897737dd104b51631d1bbe1aedc01c89836b562464208e25d8eef776e6e5a346c27ad634afef9bb45940c6444246ab54b8bcfa8b06a3acc1c21ade9d636933f19f5a2a21e65;
    5'b10111 : xpb = 1024'h1307e49830665ab48822cd664c293cca2f8afcb5d12f988d8c8ec0a67638aa1a6d66f95c6180820e97924626089088e0a80333f2f4e8cb2dbf58d1e9149206d8184f74c698322c0a3620b59118a0d0d85e8dfb1f137513a83bcfe5883fda3d963befebb06bfa553edbf4d6f9c46e20a7bba7567e1c4536a9b212dcb98a1ba219;
    5'b11000 : xpb = 1024'h8ec38e121d96141069333ff53974f69c5404845a20dded6c64a8f0e950ef139b95d58802568a9cf801e553d36f7414f1a70a683970bd386463ecda98f078b15cefd7ec6a2413a67d7d12d58e14bb1f9fa83e9247c3f8e5f2d2f7f0e38c7bd2bfad2c23f67c595ee6d3f44946b103b70e8b5c6fbcdaebf44d17561a81fa778c38;
    5'b11001 : xpb = 1024'h59d1f23648d798a37f3e3aad1666691d070808cd9b14a1d3bee667d678a2d014bafb992f816e3952ccda2239f2f9903841f77499c9ded54f57e1a3ea918ce73053112f5f006423abb16af2e877f9aa35fdea2fd7e7f68b2cb4936a441ef2c556ef60ca12dbef70014533d4b4a5c9274c0c37aa19494754c03629dd45e1f10fec;
    5'b11010 : xpb = 1024'h24e0565a74191d3695493564f357db9dba0b8d41154b563b1923dec3a0568c8de021aa5cac51d5ad97cef0a0767f0b7edce480fa2300723a4bd66d3c32a11d03b64a7253dcb4a0d9e5c31042db3834cc5395cd680bf43066962ee3a4b169b7ee3195702f3b85811bb67360229a8e97898d12e475b7a2b53354fda009c96a93a0;
    5'b11011 : xpb = 1024'ha09bffd46148d6927659a7f3e0a3956fde8514e564f9ab19f13e0f067b0cf60f08903902a15bf0970221fe4ddd62978fdbebb5409ed4df70f06a75ec0e87c7888dd2e9f768961b4d2cb5303fd75283939d466490bc7802b12d56eefffe0b4d17a2d1a8754be48ac3ae72d26f87242df05cc7fdb4764972d6ba40ddd239c67dbf;
    5'b11100 : xpb = 1024'h6baa63f88c8a5b258c64a2abbd9507f091889958df305f814b7b85f3a2c0b2882db64a2fcc3f8cf1cd16ccb460e812d676d8c1a0f7f67c5be45f3f3daf9bfd5bf10c2cec44e6987b610d4d9a3a910e29f2f20220e075a7eb0ef2686090823faee5064e91ab7a9bde1fb25ddd7be99e2ddda33810e4a4d349d914a09621400173;
    5'b11101 : xpb = 1024'h36b8c81cb7cbdfb8a26f9d639a867a71448c1dcc596713e8a5b8fce0ca746f0152dc5b5cf723294c980b9b1ae46d8e1d11c5ce0151181946d854088f50b0332f54456fe1213715a995656af49dcf98c0489d9fb104734d24f08de1c122f93246273af4ae0b10acf890f1e94b70af0e6b5e7e726d530033bcf7e8635a08b98527;
    5'b11110 : xpb = 1024'h1c72c40e30d644bb87a981b7777ecf1f78fa23fd39dc84ffff673cdf2282b7a78026c8a2206c5a76300698167f30963acb2da61aa39b631cc48d1e0f1c46902b77eb2d5fd8792d7c9bd884f010e23569e493d412870f25ed2295b21b57024dd696f9aca6aa6be13023174b965747ea8df59acc9c15b943016bc261df03308db;
    5'b11111 : xpb = 1024'h7d82d5bad03d1da7998b0aaa64c3a6c41c0929e4234c1d2ed810a410ccde94fba070fb301710e090cd53772eced69574abba0ea8260e236870dcda90cdab13878f072a7989690d4b10afa84bfd28721de7f9d469d8f4c4a96951667d0211ba06daabd3107b05c7bafa30e706520a150faf0ec608800251d37bff63e6608ef2fa;
    endcase
end

endmodule

module xpb_5_425
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'hb30558d6a92c5fee948c87234f11b233b890193a4d0305aa0971f6fc14e07f38957403275c0ed134179e24c75539d230985a33f148665984df9db4469ac82fe3b5ba75db9ee729a6cd135ac1703b460f8359ba1ac63e12e037b6c387bf3f4c3db15a896dc2aec1b7035d736ff76156ef809ae55041cac71b89df2f9ba19bbea;
    5'b00010 : xpb = 1024'h1660ab1ad5258bfdd29190e469e236467712032749a060b5412e3edf829c0fe712ae8064eb81da2682f3c498eaa73a46130b467e290ccb309bf3b688d35905fc76b74ebb73dce534d9a26b582e0768c1f06b374358c7c25c06f6d870f7e7e987b62b512db855d836e06bae6dfeec2addf0135caa083958e3713be5f3743377d4;
    5'b00011 : xpb = 1024'h219100a83fb851fcbbda59569ed35169b29b04baee70910fe1c55e4f43ea17da9c05c0976142c739c46da6e55ffad7691c90e9bd3d9330c8e9ed91cd3d0588fab212f6192dcb57cf4673a104450b1d22e8a0d2e5052ba38a0a7244a973dbde4b9140f9c49480c45250a185a4fe62404ce81d0aff0c56055529d9d8ed2e4d33be;
    5'b00100 : xpb = 1024'h2cc15635aa4b17fba52321c8d3c46c8cee24064e9340c16a825c7dbf05381fce255d00c9d703b44d05e78931d54e748c26168cfc5219966137e76d11a6b20bf8ed6e9d76e7b9ca69b344d6b05c0ed183e0d66e86b18f84b80dedb0e1efcfd30f6c56a25b70abb06dc0d75cdbfdd855bbe026b9541072b1c6e277cbe6e866efa8;
    5'b00101 : xpb = 1024'h37f1abc314ddddfa8e6bea3b08b587b029ad07e23810f1c522f39d2ec68627c1aeb440fc4cc4a16047616b7e4aa211af2f9c303b669ffbf985e14856105e8ef728ca44d4a1a83d0420160c5c731285e4d90c0a285df365e611691d1a6bc3c7d3476c4af24cd69c89310d3412fd4e6b2ad83067a9148f5e389b15bee0a280ab92;
    5'b00110 : xpb = 1024'h432201507f70a3f977b4b2ad3da6a2d365360975dce1221fc38abc9e87d42fb5380b812ec2858e7388db4dcabff5aed23921d37a7b266191d3db239a7a0b11f56425ec325b96af9e8ce742088a163a45d141a5ca0a57471414e48952e7b7bc972281f389290188a4a1430b49fcc48099d03a15fe18ac0aaa53b3b1da5c9a677c;
    5'b00111 : xpb = 1024'h4e5256ddea0369f860fd7b1f7297bdf6a0bf0b0981b1527a6421dc0e492237a8c162c16138467b86ca55301735494bf542a776b98facc72a21d4fedee3b794f39f81939015852238f9b877b4a119eea6c977416bb6bb2842185ff58b63abb15afd979c20052c74c01178e280fc3a9608c843c4531cc8b71c0c51a4d416b42366;
    5'b01000 : xpb = 1024'h5982ac6b54962ff74a464391a788d919dc480c9d268182d504b8fb7e0a703f9c4aba0193ae07689a0bcf1263aa9ce9184c2d19f8a4332cc26fceda234d6417f1dadd3aedcf7394d36689ad60b81da307c1acdd0d631f09701bdb61c3df9fa61ed8ad44b6e15760db81aeb9b7fbb0ab77c04d72a820e5638dc4ef97cdd0cddf50;
    5'b01001 : xpb = 1024'h64b301f8bf28f5f6338f0c03dc79f43d17d10e30cb51b32fa5501aedcbbe478fd41141c623c855ad4d48f4b01ff0863b55b2bd37b8b9925abdc8b567b7109af01638e24b8962076dd35ae30ccf215768b9e278af0f82ea9e1f56cdfc5b939ae2b3c2ed4dbd824cf6f1e490eefb26c0e6b85720fd25020fff7d8d8ac78ae79b3a;
    5'b01010 : xpb = 1024'h6fe3578629bbbbf51cd7d476116b0f60535a0fc47021e38a45e73a5d8d0c4f835d6881f8998942c08ec2d6fc9544235e5f386076cd3ff7f30bc290ac20bd1dee519489a943507a08402c18b8e6250bc9b2181450bbe6cbcc22d23a34d7878fa68ed895e499ad3912621a6825fa9cd655b060cf52291ebc71362b7dc145015724;
    5'b01011 : xpb = 1024'h7b13ad13944e81f406209ce8465c2a838ee3115814f213e4e67e59cd4e5a5776e6bfc22b0f4a2fd3d03cb9490a97c08168be03b5e1c65d8b59bc6bf08a69a0ec8cf03106fd3eeca2acfd4e64fd28c02aaa4daff2684aacfa264da66d537b846a69ee3e7b75d8252dd2503f5cfa12ebc4a86a7da72d3b68e2eec970baff1b130e;
    5'b01100 : xpb = 1024'h864402a0fee147f2ef69655a7b4d45a6ca6c12ebb9c2443f8715793d0fa85f6a7017025d850b1ce711b69b957feb5da47243a6f4f64cc323a7b64734f41623eac84bd864b72d5f3d19ce8411142c748ba2834b9414ae8e2829c912a5cf6f792e4503e7125203114942861693f9890133a0742bfc31581554a76763b4b934cef8;
    5'b01101 : xpb = 1024'h9174582e69740df1d8b22dccb03e60ca05f5147f5e92749a27ac98acd0f6675df96e428ffacc09fa53307de1f53efac77bc94a340ad328bbf5b022795dc2a6e903a77fc2711bd1d7869fb9bd2b3028ec9ab8e735c1126f562d447ede4b636df220198fa92e2dfd64b2bbedcaf8ff16a2987dda513574c1c6600556ae734e8ae2;
    5'b01110 : xpb = 1024'h9ca4adbbd406d3f0c1faf63ee52f7bed417e16130362a4f4c843b81c92446f5182c582c2708cf70d94aa602e6a9297ea854eed731f598e5443a9fdbdc76f29e73f0327202b0a4471f370ef694233dd4d92ee82d76d76508430bfeb16c75762b5fb2f38400a58e98022f1c501f8752c11908788a639916e3818a349a82d6846cc;
    5'b01111 : xpb = 1024'ha7d503493e9999efab43beb11a2097107d0717a6a832d54f68dad78c539277450c1cc2f4e64de420d624427adfe6350d8ed490b233dff3ec91a3d902311bace57a5ece7de4f8b70c60422515593791ae8b241e7919da31b2343b574f434b5779d644e0d6e683d59b93279c38f7eb4180889136fb3dae1aa9d1413ca1e78202b6;
    5'b10000 : xpb = 1024'h2581380e73e2b25c9870f4c3eb76ae2471a1609778b65328b953da661ddd230922b85ae91e852a5783fe58071dbc16634400c0b25b389392efe74e85ff5bb32416b412cef562c61ba79581ed75f81de8f54c08239b7e5cf822a318d0514a9ab8252f74411e5c9297c9d8c90ff9130c631c1066df17f69eb436fb49718b95835;
    5'b10001 : xpb = 1024'hd88690e51d0f124b2cfd7be73a8860582a3179d1c5b958d2c2c5d16232bda241b82c5e107a93fb8b9b9c7cce72f5e893dc5af4a3a39eed17cf8502cc9a23e307cc6e88aa9449efc274a8dcaee63363f878a5c23e61bc6fd85a59dc581089e6f5d689fdaee10b544ecd363c7ff07463529cab4c2f59c165cfc0da790d2d3141f;
    5'b10010 : xpb = 1024'h18b8be9bbc63b7239c18a030a899a128be2c1930c12bc5e7ccc37c85e479e217a4da06137d6a2ccbfb33aa195c82fbac474b52894ec05469caf22b71334ec12eb8228fe863331196941bc3770566eaa07fbff7c5927fa82b892109fdfcfc9333387e4871ca3ba1605d093afefe7d5ba421d46317f9b8c2ceb4ab9a8a8cecd009;
    5'b10011 : xpb = 1024'h23e9142926f67d22856168a2dd8abc4bf9b51ac465fbf6426d5a9bf5a5c7ea0b2e314645f32b19df3cad8c65d1d698cf50d0f5c86346ba0218ec06b59cfb442cf37e37461d21843100ecf9231c6a9f0177f593673ee389598c9c763678f087f71393f108a6668d7bcd3f1235fdf3711319de116cfdd56f406d498d8447068bf3;
    5'b10100 : xpb = 1024'h2f1969b6918943216eaa3115127bd76f353e1c580acc269d0df1bb656715f1feb788867868ec06f27e276eb2472a35f25a56990777cd1f9a66e5e1fa06a7c72b2ed9dea3d70ff6cb6dbe2ecf336e5362702b2f08eb476a879017e26ef4e47cbaeea9999f829179973d74e96cfd69868211e7bfc201f21bb225e7807e012047dd;
    5'b10101 : xpb = 1024'h3a49bf43fc1c092057f2f987476cf29270c71debaf9c56f7ae88dad52863f9f240dfc6aadeacf405bfa150febc7dd31563dc3c468c538532b4dfbd3e70544a296a35860190fe6965da8f647b4a7207c36860caaa97ab4bb593934ea770d8717ec9bf42365ebc65b2adaac0a3fcdf9bf109f16e17060ec823de857377bb3a03c7;
    5'b10110 : xpb = 1024'h457a14d166aecf1f413bc1f97c5e0db5ac501f7f546c87524f1ffa44e9b201e5ca3706dd546de119011b334b31d170386d61df85a0d9eacb02d99882da00cd27a5912d5f4aecdc0047609a276175bc246096664c440f2ce3970ebadfeccc6642a4d4eacd3ae751ce1de097dafc55b16001fb1c6c0a2b7495972366717553bfb1;
    5'b10111 : xpb = 1024'h50aa6a5ed141951e2a848a6bb14f28d8e7d92112f93cb7acefb719b4ab0009d9538e470fca2ece2c42951597a7250d5b76e782c4b560506350d373c743ad5025e0ecd4bd04db4e9ab431cfd37879708558cc01edf0730e119a8a271868c05b067fea936417123de98e166f11fbcbc6cefa04cac10e4821074fc1596b2f6d7b9b;
    5'b11000 : xpb = 1024'h5bdabfec3bd45b1d13cd52dde64043fc236222a69e0ce807904e39246c4e11ccdce587423fefbb3f840ef7e41c78aa7e806d2603c9e6b5fb9ecd4f0bad59d3241c487c1abec9c1352103057f8f7d24e651019d8f9cd6ef3f9e059350e4b44fca5b003bfaf33d2a04fe4c4648fb41dc3df20e79161264cd79085f4c64e9873785;
    5'b11001 : xpb = 1024'h670b1579a667211bfd161b501b315f1f5eeb243a42dd186230e558942d9c19c0663cc774b5b0a852c588da3091cc47a189f2c942de6d1b93ecc72a501706562257a4237878b833cf8dd43b2ba680d94749373931493ad06da180ff8960a8448e3615e491cf6816206e821d7ffab7f1acea18276b168179eac0fd3f5ea3a0f36f;
    5'b11010 : xpb = 1024'h723b6b0710f9e71ae65ee3c250227a429a7425cde7ad48bcd17c7803eeea21b3ef9407a72b7195660702bc7d071fe4c493786c81f2f3812c3ac1059480b2d92092ffcad632a6a669faa570d7bd848da8416cd4d2f59eb19ba4fc6bc1dc9c3952112b8d28ab93023bdeb7f4b6fa2e071be221d5c01a9e265c799b32585dbaaf59;
    5'b11011 : xpb = 1024'h7d6bc0947b8cad19cfa7ac3485139565d5fd27618c7d791772139773b03829a778eb47d9a1328279487c9ec97c7381e79cfe0fc10779e6c488bae0d8ea5f5c1ece5b7233ec9519046776a683d488420939a27074a20292c9a877d7fa58902e15ec4135bf87bdee574eedcbedf9a41c8ada2b84151ebad2ce3239255217d46b43;
    5'b11100 : xpb = 1024'h889c1621e61f7318b8f074a6ba04b089118628f5314da97212aab6e37186319b0242880c16f36f8c89f68115f1c71f0aa683b3001c004c5cd6b4bc1d540bdf1d09b71991a6838b9ed447dc2feb8bf66a31d80c164e6673f7abf34432d48422d9c756de5663e8da72bf23a324f91a31f9d235326a22d77f3fead7184bd1ee272d;
    5'b11101 : xpb = 1024'h93cc6baf50b23917a2393d18eef5cbac4d0f2a88d61dd9ccb341d65332d4398e8b99c83e8cb45c9fcb706362671abc2db009563f3086b1f524ae9761bdb8621b4512c0ef6071fe39411911dc028faacb2a0da7b7faca5525af6eb06b5078179da26c86ed4013c68e2f597a5bf8904768ca3ee0bf26f42bb1a3750b458c07e317;
    5'b11110 : xpb = 1024'h9efcc13cbb44ff168b82058b23e6e6cf88982c1c7aee0a2753d8f5c2f422418214f10871027549b30cea45aedc6e5950b98ef97e450d178d72a872a62764e519806e684d1a6070d3adea478819935f2c22434359a72e3653b2ea1ca3cc6c0c617d822f841c3eb2a99f8f5192f8065cd7c2488f142b10d8235c12fe3f46219f01;
    5'b11111 : xpb = 1024'haa2d16ca25d7c51574cacdfd58d801f2c4212db01fbe3a81f4701532b57049759e4848a3783636c64e6427fb51c1f673c3149cbd59937d25c0a24dea91116817bbca0faad44ee36e1abb7d343097138d1a78defb53921781b66588dc486001255897d81af8699ec50fc528c9f77c7246ba523d692f2d849514b0f139003b5aeb;
    endcase
end

endmodule

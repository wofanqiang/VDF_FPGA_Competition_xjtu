module xpb_5_20
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h56eb5faa0a214ecdd0b7fb91254b6933eef2e17149bd01feceffa1905c8895f271ada45f24407c6341c00d5bff77fada6533f15cba5adcdb7324e9075646e1eaa240911aff6da049a21c6f76384c9f22918251566a45f92b7ec561f3055a34d3d87a9ad02738da2014149a8b4ae8a1459772fa416b24896e07e0d4904d5a27d6;
    5'b00010 : xpb = 1024'hadd6bf5414429d9ba16ff7224a96d267dde5c2e2937a03fd9dff4320b9112be4e35b48be4880f8c683801ab7feeff5b4ca67e2b974b5b9b6e649d20eac8dc3d544812235fedb40934438deec70993e452304a2acd48bf256fd8ac3e60ab469a7b0f535a04e71b4402829351695d1428b2ee5f482d64912dc0fc1a9209ab44fac;
    5'b00011 : xpb = 1024'h5414d9a85c75b7a0a7227adc5f87f44a5b62a12307bf6584ef222b5b629714cf51c06fa4a29af69b25e1e8cd1b09dfc4cb81ac300c5dc646a8cf7bb7c802310e72727ea24eb7e397d3bb4bc0100a1936c081fa6ab24bbe71c6c393de55e3fbe95a683e46c4e195d2b57de8c2e8e9bda7777f0fe1f1223f19d13302ac5f2c1117;
    5'b00100 : xpb = 1024'hab0039526697066e77da766d84d35d7e4a558294517c6783be21ccebbf1faac1c36e1403c6db72fe67a1f6291a81da9f30b59d8cc6b8a3221bf464bf1e4912f914b30fbd4e2583e175d7bb364856b85952044bc11c91b79d4588f5d15b3e30bd32e2d916ec1a6ff2c992834e33d25eed0ef20a235c46c887d913d73cac8638ed;
    5'b00101 : xpb = 1024'h513e53a6aeca20737d8cfa2799c47f60c7d260d4c5c1c90b0f44b52668a593ac31d33aea20f570d30a03c43e369bc4af31cf67035e60afb1de7a0e6839bd803242a46c299e0226e6055a2809e7c7934aef81a37efa5183b80ec1c5c9a66dc2fedc55e1bd628a518556e736fa86eada09578b2582771ff4c59a8530c870fdfa58;
    5'b00110 : xpb = 1024'ha829b350b8eb6f414e44f5b8bf0fe894b6c542460f7ecb09de4456b6c52e299ea380df494535ed364bc3d19a3613bf899703586018bb8c8d519ef76f9004621ce4e4fd449d6fc72fa77697802014326d8103f4d564977ce38d8727bcabc7f7d2b4d07c8d89c32ba56afbd185d1d37b4eeefe1fc3e2447e33a2660558be58222e;
    5'b00111 : xpb = 1024'h4e67cda5011e894653f77972d4010a773442208683c42c912f673ef16eb4128911e6062f9f4feb0aee259faf522da999981d21d6b063991d1424a118ab78cf5612d659b0ed4c6a3436f90453bf850d5f1e814c93425748fe56bff7b4f6f78a145e43853400330d37f850853224ebf66b37973b22fd1daa7163d75ee482cfe399;
    5'b01000 : xpb = 1024'ha5532d4f0b3fd81424af7503f94c73ab233501f7cd812e8ffe66e081cb3ca87b8393aa8ec390676e2fe5ad0b51a5a473fd5113336abe75f887498a2001bfb140b516eacbecba0a7dd91573c9f7d1ac81b0039de9ac9d4229d58559a7fc51bee836be2004276be7580c651fbd6fd497b0cf0a3564684233df6bb83374d02a0b6f;
    5'b01001 : xpb = 1024'h4b9147a35372f2192a61f8be0e3d958da0b1e03841c690174f89c8bc74c29165f1f8d1751daa6542d2477b206dbf8e83fe6adcaa0266828849cf33c91d341e79e30847383c96ad826897e09d974287734d80f5a78a5d0e449ebe29a047815129e03128aa9ddbc8ea99b9d369c2ed12cd17a350c3831b601d2d298d0094a1ccda;
    5'b01010 : xpb = 1024'ha27ca74d5d9440e6fb19f44f3388fec18fa4c1a98b8392161e896a4cd14b275863a675d441eae1a61407887c6d37895e639ece06bcc15f63bcf41cd0737b00648548d8533c044dcc0ab45013cf8f2695df0346fdf4a307701d838b934cdb85fdb8abc37ac514a30aadce6df50dd5b412af164b04ee3fe98b350a6190e1fbf4b0;
    5'b01011 : xpb = 1024'h48bac1a1a5c75aec00cc7809487a20a40d219fe9ffc8f39d6fac52877ad11042d20b9cba9c04df7ab66956918951736e64b8977d54696bf37f79c6798eef6d9db33a34bf8be0f0d09a36bce76f0001877c809ebbd262d38ae6bc5b8b980b183f621ecc213b84849d3b2321a160ee2f2ef7af6664091915c8f67bbb1ca673b61b;
    5'b01100 : xpb = 1024'h9fa6214bafe8a9b9d184739a6dc589d7fc14815b4985f59c3eabf417d759a63543b94119c0455bddf82963ed88c96e48c9ec88da0ec448cef29eaf80e5364f88557ac5da8b4e911a3c532c5da74ca0aa0e02f0123ca8ccb66581bd7e9d654d133a9966f162bd5ebd4f37bc2cabd6d0748f2260a5743d9f36fe5c8facf3cdddf1;
    5'b01101 : xpb = 1024'h45e43b9ff81bc3bed736f75482b6abba79915f9bbdcb57238fcedc5280df8f1fb21e68001a5f59b29a8b3202a4e35858cb065250a66c555eb524592a00aabcc1836c2246db2b341ecbd5993146bd7b9bab8047d01a6898d12eba8d76e894df54e40c6f97d92d404fdc8c6fd8feef4b90d7bb7c048f16cb74bfcde938b8459f5c;
    5'b01110 : xpb = 1024'h9ccf9b4a023d128ca7eef2e5a80214ee6884410d078859225ece7de2dd68251223cc0c5f3e9fd615dc4b3f5ea45b5333303a43ad60c7323a2849423156f19eac25acb361da98d4686df208a77f0a1abe3d02992684ae91fcad7fef69edef1428bc870a6800661a6ff0a10a6449d7ecd66f2e7645fa3b54e2c7aebdc9059fc732;
    5'b01111 : xpb = 1024'h430db59e4a702c91ada1769fbcf336d0e6011f4d7bcdbaa9aff1661d86ee0dfc9231334598b9d3ea7ead0d73c0753d4331540d23f86f3ec9eaceebda72660be5539e0fce2a75776cfd74757b1e7af5afda7ff0e4626e5e1776b8bf62391ea66a65fa130e76d5fc027df5be109cf067f2b7c791a51514812089201754ca17889d;
    5'b10000 : xpb = 1024'h99f9154854917b5f7e597230e23ea004d4f400bec58abca87ef107ade376a3ef03ded7a4bcfa504dc06d1acfbfed381d9687fe80b2ca1ba55df3d4e1c8acedcff5dea0e929e317b69f90e4f156c794d26c02423accb45742f57e21553e78db3e3e74adde9e0ed622920a589be7d909384f3a8be680390a8e9100ebe51771b073;
    5'b10001 : xpb = 1024'h40372f9c9cc49564840bf5eaf72fc1e75270deff39d01e2fd013efe88cfc8cd97243fe8b17144e2262cee8e4dc07222d97a1c7f74a72283520797e8ae4215b0923cffd5579bfbabb2f1351c4f6386fc4097f99f8aa74235dbeb6f14d89a86d7fe7e7b685147eb7b51f5f0c483af1845497d3a7459b1236cc52724570dbe971de;
    5'b10010 : xpb = 1024'h97228f46a6e5e43254c3f17c1c7b2b1b4163c070838d202e9f139178e98522cbe3f1a2ea3b54ca85a48ef640db7f1d07fcd5b95404cd0510939e67923a683cf3c6108e70792d5b04d12fc13b2e850ee69b01eb4f14ba1c893d7c53408f02a253c06251553bb791d53373a6d385da259a2f46a1870636c03a5a531a01294399b4;
    5'b10011 : xpb = 1024'h3d60a99aef18fe375a767536316c4cfdbee09eb0f7d281b5f03679b3930b0bb65256c9d0956ec85a46f0c455f7990717fdef82ca9c7511a05624113b55dcaa2cf401eadcc909fe0960b22e0ecdf5e9d8387f430cf279e8a406b52338da32349569d559fbb2277367c0c85a7fd8f2a0b677dfbce6210fec781bc4738cedbb5b1f;
    5'b10100 : xpb = 1024'h944c0944f93a4d052b2e70c756b7b631add38022418f83b4bf361b43ef93a1a8c4046e2fb9af44bd88b0d1b1f71101f26323742756cfee7bc948fa42ac238c1796427bf7c8779e5302ce9d85064288faca0194635cbfe1cf857a852bdf8c6969424ff4cbd9604d87d4dcf50b23db41fc0f52b7278c3475e623a5481d3b1582f5;
    5'b10101 : xpb = 1024'h3a8a2399416d670a30e0f4816ba8d8142b505e62b5d4e53c1059037e99198a933269951613c942922b129fc7132aec02643d3d9dee77fb0b8bcea3ebc797f950c433d8641854415792510a58a5b363ec677eec213a7fadea4eb355242abbfbaaebc2fd724fd02f1a6231a8b776f3bd1857ebd286a70da223e516a1a8ff8d4460;
    5'b10110 : xpb = 1024'h917583434b8eb5d80198f01290f441481a433fd3ff91e73adf58a50ef5a22085a41739753809bef56cd2ad2312a2e6dcc9712efaa8d2d7e6fef38cf31ddedb3b6674697f17c1e1a1346d79cede00030ef9013d77a4c5a715cd78b7173016307ec43d98427709093a76464342c1dc5e5def5eccc812322b91ecf776394ce76c36;
    5'b10111 : xpb = 1024'h37b39d9793c1cfdd074b73cca5e5632a97c01e1473d748c2307b8d499f280970127c605b9223bcca0f347b382ebcd0ecca8af871407ae476c179369c395348749465c5eb679e84a5c3efe6a27d70de00967e95358285733096b1870f7b45c2c06db0a0e8ed78eacd039af6ef14f4d97a37f7e8272d0b57cfae68cfc5115f2da1;
    5'b11000 : xpb = 1024'h8e9efd419de31eaad8036f5dcb30cc5e86b2ff85bd944ac0ff7b2ed9fbb09f62842a04bab664392d50f488942e34cbc72fbee9cdfad5c152349e1fa38f9a2a5f36a65706670c24ef660c5618b5bd7d232800e68beccb6c5c1576e902809ff794462b3bb914b1c4ed17af917a5fdd7abfcf6ae268982fe13db649a4555eb95577;
    5'b11001 : xpb = 1024'h34dd1795e61638afddb5f317e021ee41042fddc631d9ac48509e1714a536884cf28f2ba1107e3701f35656a94a4eb5d730d8b344927dcde1f723c94cab0e97986497b372b6e8c7f3f58ec2ec552e5814c57e3e49ca8b3876deafb8facbcf89d5ef9e445f8b21a67fa5044526b2f5f5dc1803fdc7b3090d7b77bafde1233116e2;
    5'b11010 : xpb = 1024'h8bc8773ff037877dae6deea9056d5774f322bf377b96ae471f9db8a501bf1e3f643cd00034beb3653516640549c6b0b1960ca4a14cd8aabd6a48b2540155798306d8448db656683d97ab32628d7af73757008fa034d131a25d751aedd129bea9c818df2fb25a809fb918dfb1fdde9721af76f8091e2d96e97f9bd271708b3eb8;
    5'b11011 : xpb = 1024'h32069194386aa182b42072631a5e7957709f9d77efdc0fce70c0a0dfab450729d2a1f6e68ed8b139d778321a65e09ac197266e17e480b74d2cce5bfd1cc9e6bc34c9a0fa06330b42272d9f362cebd228f47de75e1290fdbd26adeae61c5950eb718be7d628ca6232466d935e50f7123df81013683906c327410d2bfd35030023;
    5'b11100 : xpb = 1024'h88f1f13e428bf05084d86df43fa9e28b5f927ee9399911cd3fc0427007cd9d1c444f9b45b3192d9d19383f766558959bfc5a5f749edb94289ff345047310c8a6d70a321505a0ab8bc94a0eac6538714b860038b47cd6f6e8a5734cd921b385bf4a0682a650033c525a822de99bdfb3838f830da9a42b4c9548ee008d825d27f9;
    5'b11101 : xpb = 1024'h2f300b928abf0a558a8af1ae549b046ddd0f5d29adde735490e32aaab1538606b2b4c22c0d332b71bb9a0d8b81727fabfd7428eb3683a0b86278eead8e8535e004fb8e81557d4e9058cc7b8004a94c3d237d90725a96c3036eac1cd16ce31800f3798b4cc6731de4e7d6e195eef82e9fd81c2908bf0478d30a5f5a1946d4e964;
    5'b11110 : xpb = 1024'h861b6b3c94e059235b42ed3f79e66da1cc023e9af79b75535fe2cc3b0ddc1bf92462668b3173a7d4fd5a1ae780ea7a8662a81a47f0de7d93d59dd7b4e4cc17caa73c1f9c54eaeed9fae8eaf63cf5eb5fb4ffe1c8c4dcbc2eed717ec4723d4cd4cbf4261cedabf804fbeb7c2139e0cfe56f8f234a2a29024112402ea9942f113a;
    5'b11111 : xpb = 1024'h2c598590dd13732860f570f98ed78f84497f1cdb6be0d6dab105b475b76204e392c78d718b8da5a99fbbe8fc9d04649663c1e3be88868a239823815e00408503d52d7c08a4c791de8a6b57c9dc66c651527d3986a29c8849b6aa4ebcbd6cdf1675672ec3641bd99789402fcd8cf94b01b8283ea945022e7ed3b1883558a6d2a5;
    endcase
end

endmodule

module xpb_5_610
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h3bc1f09483730de77bb05e25814924201e068ad97b0c7b35be10b5fe965a60546433bcfa9ca60f1507119e5baa31cf0d1b241fe685449cda822d9f620043bd1fba3c2dc1dc2f8bcc71fb652022578eb69a96cd9fe6858de4c956c84c2e3df2792b641d667b4f35fa9c444db01897e0f207f52c4cb50ced67ea0b660f1123212a;
    5'b00010 : xpb = 1024'h7783e12906e61bcef760bc4b029248403c0d15b2f618f66b7c216bfd2cb4c0a8c86779f5394c1e2a0e233cb754639e1a36483fcd0a8939b5045b3ec400877a3f74785b83b85f1798e3f6ca4044af1d6d352d9b3fcd0b1bc992ad90985c7be4f256c83accf69e6bf538889b60312fc1e40fea58996a19dacfd416cc1e22464254;
    5'b00011 : xpb = 1024'h2988c67c86af4eda80ba2997381250ee89d9d5b9badd129bc5568a6100c73f52952b9770bcbaeb075d69bcc1b375c5ced5237cd6d1b0643d5e99ec7c5f8c2adba655496e4fda62043582cbdce2ae7f2dbbf6f47270a7c9da677c6e9d08f34d95324c609c124a9624e0d023151f77cacc905a603cedb6b0777b2b728aa86fd13;
    5'b00100 : xpb = 1024'h3e5a7cfc4bde02d523bc00bef4ca492f06a4283516ba4c5f7a661ea4a666d4498d867671a871bdc57ce83a27c5692b6a087657b3f25fa31e58173e29c63c7fcd74a18258c12d31ecb55391ddf08276a976563ce70d900a826fce8f35fecd27527e88e3703c73df5cea514fe16a8f5d9ed0fad25083e8586f61be1d37bbaa1e3d;
    5'b00101 : xpb = 1024'h7a1c6d90cf5110bc9f6c5ee476136d4f24aab30e91c6c7953876d4a33cc1349df1ba336c4517ccda83f9d8836f9afa77239a779a77a43ff8da44dd8bc6803ced2eddb01a9d5cbdb9274ef6fe12da056010ed0a86f4159867392557822d0b19cba9ed00d6b7c3155786959d9183273e90d8effe9d38f545d74bc98346cccd3f67;
    5'b00110 : xpb = 1024'h53118cf90d5e9db50174532e7024a1dd13b3ab7375ba25378aad14c2018e7ea52a572ee17975d60ebad3798366eb8b9daa46f9ada360c87abd33d8f8bf1855b74caa92dc9fb4c4086b0597b9c55cfe5b77ede8e4e14f93b4cef8dd3a11e69b2a6498c13824952c49c1a0462a3eef959920b4c079db6d60eef656e51550dfa26;
    5'b00111 : xpb = 1024'h40f309641448f7c2cbc7a358684b6e3def41c590b2681d8936bb874ab673483eb6d92fe8b43d6c75f2bed5f3e0a087c6f5c88f815f7aa9622e00dcf18c35427b2f06d6efa62ad80cf8abbe9bbead5e9c5215ac2e349a87201646561fcf5c5c2bd1ada979fd9888bf385e5212bc86da4b9a00785452c3c376d970d46066311b50;
    5'b01000 : xpb = 1024'h7cb4f9f897bc05aa4778017de994925e0d48506a2d7498bef4cc3d494ccda8931b0cece350e37b8af9d0744f8ad256d410ecaf67e4bf463cb02e7c538c78ff9ae94304b1825a63d96aa723bbe104ed52ecac79ce1b201504df9d1e6bfd9a4ea4fd11c6e078e7beb9d4a29fc2d51ebb3da1f5a4a107d0b0dec37c3a6f77543c7a;
    5'b01001 : xpb = 1024'h7c9a5375940dec8f822e7cc5a836f2cb9d8d812d309737d350039f230255bdf7bf82c6523630c116183d36451a61516c7f6a768475112cb81bcdc5751ea48092f2ffdc4aef8f260ca0886396a80b7d8933e4dd5751f75d8f36754bd71ad9e8bf96e521d436dfc26ea270693f5e676065b10f20b6c92411667182579ff94f739;
    5'b01010 : xpb = 1024'h438b95cbdcb3ecb073d345f1dbcc934cd7df62ec4e15eeb2f310eff0c67fbc33e02be95fc0091b26689571bffbd7e423e31ac74ecc95afa603ea7bb9522e0528e96c2b868b287e2d3c03eb598cd8468f2dd51b755ba503bdbcbe1d099feb910524d26f83bebd3221866b54440e7e56f863061e58219f2e7e51238b8910b81863;
    5'b01011 : xpb = 1024'h7f4d86606026fa97ef83a4175d15b76cf5e5edc5c92269e8b121a5ef5cda1c88445fa65a5caf2a3b6fa7101ba609b330fe3ee73551da4c8086181b1b5271c248a3a85948675809f9adff5079af2fd545c86be915422a91a28614e555ce29837e50368cea3a0c681c22afa1f4271637ea6afb4aa4d6ac1be63b2ef19821db398d;
    5'b01100 : xpb = 1024'ha62319f21abd3b6a02e8a65ce04943ba276756e6eb744a6f155a2984031cfd4a54ae5dc2f2ebac1d75a6f306cdd7173b548df35b46c190f57a67b1f17e30ab6e995525b93f698810d60b2f738ab9fcb6efdbd1c9c29f27699df1ba7423cd3654c9318270492a589383408c547ddf2b32416980f3b6dac1ddecadca2aa1bf44c;
    5'b01101 : xpb = 1024'h46242233a51ee19e1bdee88b4f4db85bc07d0047e9c3bfdcaf665896d68c3029097ea2d6cbd4c9d6de6c0d8c170f4080d06cff1c39b0b5e9d9d41a811826c7d6a3d1801d7026244d7f5c18175b032e8209948abc82af805b6335e3f3707ac5de77f7358d7fe1db83d47856756075d3a52c0bc45bf07a9985c8d642b1bb3f1576;
    5'b01110 : xpb = 1024'h81e612c82891ef85978f46b0d096dc7bde838b2164d03b126d770e956ce6907d6db25fd1687ad8ebe57dabe7c1410f8deb911f02bef552c45c01b9e3186a84f65e0daddf4c55b019f1577d377d5abd38a42b585c69350e402c8cac3f9eb8b857a35b52f3fb31117e70bca425790db4973400f0a8a58786edb2e1a8c0cc6236a0;
    5'b01111 : xpb = 1024'hcfabe06ea16c8a4483a2cff4185b94a8b1412ca0a6515d0adab0b3e503e43c9ce9d9f533afa69724d310afc8814cdd0a29b170321871f532d9019e6dddbcd64a3faa6f278f43ea150b8dfb506d687be4abd2c63c3346f144056e29112cc083e9fb7de30c5b74eeb86410af699d56f5fed1c3e130a491725567d93cb54a2f15f;
    5'b10000 : xpb = 1024'h48bcae9b6d89d68bc3ea8b24c2cedd6aa91a9da3857191066bbbc13ce698a41e32d15c4dd7a078875442a95832469cddbdbf36e9a6cbbc2dafbdb948de1f8a845e36d4b45523ca6dc2b444d5292e1674e553fa03a9b9fcf909adaadd4109fab7cb1bfb97410684e6228558a6b26d5051f5116a5fbf56048d4088f9da65c61289;
    5'b10001 : xpb = 1024'h847e9f2ff0fce4733f9ae94a4418018ac721287d007e0c3c29cc773b7cf30472970519487446879c5b5447b3dc786bead8e356d02c10590831eb58aade6347a4187302763153563a34afa9f54b85a52b7feac7a3903f8addd30473296f47ed30f68018fdbc55bae0bec9a656cb053143fd0696ac7462f1f52a945fe976e933b3;
    5'b10010 : xpb = 1024'hf934a6eb281bd91f045cf98b506de5973b1b025a612e6fa6a0073e4604ab7bef7f058ca46c61822c307a6c8a34c2a2d8fed4ed08ea225970379b8aea3d490125e5ffb895df1e4c194110c72d5016fb1267c9baaea3eebb1e6cea97ae35b3d17f2dca43a86dbf84dd44e0d27ebccec0cb621e416d924822cce304af3ff29ee72;
    5'b10011 : xpb = 1024'h4b553b0335f4cb796bf62dbe3650027991b83aff211f6230281129e2f6a518135c2415c4e36c2737ca1945244d7df93aab116eb713e6c27185a75810a4184d32189c294b3a21708e060c7192f758fe67c113694ad0c47996b02571c711992f911e40c1a1022b2e4870925ad80464ccfebe1710638e316f94b83bb103104d0f9c;
    5'b10100 : xpb = 1024'h87172b97b967d960e7a68be3b7992699afbec5d89c2bdd65e621dfe18cff7867c057d2bf8012364cd12ae37ff7afc847c6358e9d992b5f4c07d4f772a45c0a51d2d8570d1650fc5a7807d6b319b08d1e5baa36eab74a077b797c3a133fd7220a49a4df077d7a64430cd6a8881cfcadf0c60c3cb0433e5cfca2471712217030c6;
    5'b10101 : xpb = 1024'h122bd6d67aecb27f98517232288803685c4f4d8141c0b8242655dc8a70572bb4214312415291c6d338de4294be83868a7d3f869dfbbd2bdad963577669cd52c018c5502042ef8ae1d7693930a32c57a4023c0af21149684f8d467064b3ea71f146016a444800a1b0225b0f593dc468b97f278a1aa7ffed3445e3021ca9b0eb85;
    5'b10110 : xpb = 1024'h4dedc76afe5fc0671401d057a9d127887a55d85abccd3359e466928906b18c088576cf3bef37d5e83fefe0f068b555979863a6848101c8b55b90f6d86a110fdfd3017de21f1f16ae49649e50c583e65a9cd2d891f7cef634569d38b0e228646a716587aac34fd7aabe9f5d09565c49ab871cb6675d0cda9c2fee682bbad40caf;
    5'b10111 : xpb = 1024'h89afb7ff81d2ce4e8fb22e7d2b1a4ba8985c633437d9ae8fa27748879d0bec5ce9aa8c368bdde4fd47017f4c12e724a4b387c66b0646658fddbe963a6a54ccff8d3daba3fb4ea27abb600370e7db75113769a631de5484191ff400fd106656e39cc9a5113e9f0da55ae3aab96ef42a9d8f11e2b41219c80419f9ce3acbf72dd9;
    5'b11000 : xpb = 1024'h14c4633e4357a76d405d14cb9c09287744eceadcdd6e894de2ab453080639fa94a95cbb85e5d7583aeb4de60d9bae2e76a91be6b68d8321eaf4cf63e2fc6156dd32aa4b727ed31021ac165ee71573f96ddfb7a393853e4ed33be374e8479a6ca9926304e09254b127068118a8fbbe566482d301e76db583bbd95b9455437e898;
    5'b11001 : xpb = 1024'h508653d2c6cab554bc0d72f11d524c9762f375b6587b0483a0bbfb2f16bdfffdaec988b2fb038498b5c67cbc83ecb1f485b5de51ee1ccef9317a95a03009d28d8d66d279041cbcce8cbccb0e93aece4d789247d91ed972d1fd14ff9ab2b79943c48a4db48474810d0cac5f3aa853c65850225c6b2be845a3a7a11f54655b09c2;
    5'b11010 : xpb = 1024'h8c4844674a3dc33c37bdd1169e9b70b780fa008fd3877fb95eccb12dad18605212fd45ad97a993adbcd81b182e1e8101a0d9fe3873616bd3b3a83502304d8fad47a3003ae04c489afeb8302eb6065d0413291579055f00b6c66bc7e6e0f58bbcefee6b1affc3b707a8f0aceac0eba74a581788b7e0f5330b91ac8563767e2aec;
    5'b11011 : xpb = 1024'h175cefa60bc29c5ae868b7650f8a4d862d8a8838791c5a779f00add69070139e73e8852f6a292434248b7a2cf4f23f4457e3f638d5f3386285369505f5bed81b8d8ff94e0cead7225e1992ac3f822789b9bae9805f5e618ada35fe385508dba3ec4af657ca49f474be7513bbe1b362131132d62245b6c3433548706dfebee5ab;
    5'b11100 : xpb = 1024'h531ee03a8f35aa426419158a90d371a64b911311f428d5ad5d1163d526ca73f2d81c422a06cf33492b9d18889f240e517308161f5b37d53d07643467f602953b47cc270fe91a62eed014f7cc61d9b6405451b72045e3ef6fa38cc6848346ce1d17af13be45992a6f5ab9616bfa4b43051928026efac3b0ab1f53d67d0fe206d5;
    5'b11101 : xpb = 1024'h8ee0d0cf12a8b829dfc973b0121c95c669979deb6f3550e31b2219d3bd24d4473c4fff24a375425e32aeb6e44955dd5e8e2c3605e07c72178991d3c9f646525b020854d1c549eebb42105cec843144f6eee884c02c697d546ce38ed0b184c09643133124c0e86069f6fdaf1c12e323f7211d2ebbafd09e13095f3c8c210527ff;
    5'b11110 : xpb = 1024'h19f57c0dd42d9148907459fe830b72951628259414ca2ba15b56167ca07c87939d3b3ea675f4d2e49a6215f910299ba145362e06430e3ea65b2033cdbbb79ac947f54de4f1e87d42a171bf6a0dad0f7c957a58c78668de2880adc5222598107d3f6fbc618b6e9dd70c8215ed33aadebfda387c2614922e4aacfb2796a945e2be;
    5'b11111 : xpb = 1024'h55b76ca257a09f300c24b824045496b5342eb06d8fd6a6d71966cc7b36d6e7e8016efba1129ae1f9a173b454ba5b6aae605a4decc852db80dd4dd32fbbfb57e902317ba6ce18090f136d248a30049e33301126676cee6c0d4a048d6e53d602f66ad3d9c806bdd3d1a8c6639d4c42bfb1e22da872c99f1bb297068da5ba6903e8;
    endcase
end

endmodule

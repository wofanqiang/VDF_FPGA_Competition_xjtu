module xpb_5_765
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'ha401c40e013a6eff16974ca7c3a74ebaf451e34cea2161ffd8b475c8985a5ade3d1175ce78c6b638f74313d22c51013c39758546c7ca0ae26d5ed2652ed17f9c6fc5fd41efdb5ea6139cea41665555e89f258031f2b9a451f74e7c2de065722cfb095954956c6140a4f8e3db1d035ecc220599844925300ed3e322978aeba527;
    5'b00010 : xpb = 1024'h975642c64086a9356229217876f45624772dc368fecb2388338c323b7db208b476da6e242766ede34f27e85d7543f1ae0ed0e2a76ce145792a1e656c22d08a876b3cc5d53025c007149fd1e033cee7a04a4606cb58ed1b933910666106a041c7c70b207f7a0fc9f3c331e0d74236976ef531542641ff02ed6156ca2a8cf4e3e3;
    5'b00011 : xpb = 1024'h8aaac17e7fd2e36badbaf6492a415d8dfa09a3851374e5108e63eeae6309b68ab0a36679d607258da70cbce8be36e21fe42c400811f8800fe6ddf87316cf957266b38e687070216815a2b97f01487957f5668d64bf2092d47ad250942cdb1162930ce7aa5eb332a6e16addd36769d011c85d0ec83ad8d5cbeeca71bd8efe229f;
    5'b00100 : xpb = 1024'h7dff4036bf1f1da1f94ccb19dd8e64f77ce583a1281ea698e93bab2148616460ea6c5ecf84a75d37fef191740729d291b9879d68b70fbaa6a39d8b7a0acea05d622a56fbb0ba82c916a5a11dcec20b0fa08713fe25540a15bc943ac75315e0fd5f0eaed543569b59ffa3dacf8c9d08b49b88c96a33b2a8aa7c3e19509107615b;
    5'b00101 : xpb = 1024'h7153beeefe6b57d844de9fea90db6c60ffc163bd3cc86821441367942db9123724355725334794e256d665ff501cc3038ee2fac95c26f53d605d1e80fecdab485da11f8ef104e42a17a888bc9c3b9cc74ba79a978b878156fe5624fa7950b0982b10760027fa040d1ddcd7cbb1d041576eb4840c2c8c7b8909b1c0e39310a017;
    5'b00110 : xpb = 1024'h64a83da73db7920e907074bb442873ca829d43d9517229a99eeb24071310c00d5dfe4f7ae1e7cc8caebb3a8a990fb375643e582a013e2fd41d1cb187f2ccb6335917e822314f458b18ab705b69b52e7ef6c82130f1baf89840180f2d9f8b8032f7123d2b0c9d6cc03c15d4c7d70379fa41e03eae25664e67972568769519ded3;
    5'b00111 : xpb = 1024'h57fcbc5f7d03cc44dc02498bf7757b34057923f5661beb31f9c2e079f8686de397c747d09088043706a00f15e202a3e73999b58aa6556a6ad9dc448ee6cbc11e548eb0b57199a6ec19ae57fa372ec036a1e8a7ca57ee6fd981d9f960c5c64fcdc3140455f140d5735a4ed1c3fc36b29d150bf9501e4021462499100997231d8f;
    5'b01000 : xpb = 1024'h4b513b17bc50067b27941e5caac2829d885504117ac5acba549a9cecddc01bb9d19040263f283be15e84e3a12af594590ef512eb4b6ca501969bd795dacacc0950057948b1e4084d1ab13f9904a851ee4d092e63be21e71ac39be393ec011f688f15cb80d5e43e267887cec02169eb3fe837b3f21719f424b20cb79c992c5c4b;
    5'b01001 : xpb = 1024'h3ea5b9cffb9c40b17325f32d5e0f8a070b30e42d8f6f6e42af72595fc317c9900b59387bedc8738bb669b82c73e884cae450704bf083df98535b6a9ccec9d6f44b7c41dbf22e69ae1bb42737d221e3a5f829b4fd24555e5c055dcdc7123bef035b1792abba87a6d996c0cbbc469d23e2bb636e940ff3c7033f805f2f9b359b07;
    5'b01010 : xpb = 1024'h31fa38883ae87ae7beb7c7fe115c91708e0cc449a4192fcb0a4a15d2a86f7766452230d19c68ab360e4e8cb7bcdb753cb9abcdac959b1a2f101afda3c2c8e1df46f30a6f3278cb0f1cb70ed69f9b755da34a3b968a88d59d471fb7fa3876be9e271959d69f2b0f8cb4f9c8b86bd05c858e8f293608cd99e1ccf406c29d3ed9c3;
    5'b01011 : xpb = 1024'h254eb7407a34b51e0a499ccec4a998da10e8a465b8c2f1536521d2458dc7253c7eeb29274b08e2e06633614305ce65ae8f072b0d3ab254c5ccda90aab6c7ecca4269d30272c32c701db9f6756d1507154e6ac22ff0bc4cde88e1a22d5eb18e38f31b210183ce783fd332c5b49103952861bae3d801a76cc05a67ae559f48187f;
    5'b01100 : xpb = 1024'h18a335f8b980ef5455db719f77f6a04393c48481cd6cb2dbbff98eb8731ed312b8b4217cf9a91a8abe1835ce4ec156206462886ddfc98f5c899a23b1aac6f7b53de09b95b30d8dd11ebcde143a8e98ccf98b48c956efc41fcaa38c6084ec5dd3bf1ce82c6871e0f2f16bc2b0b636cdcb34e69e79fa813f9ee7db55e8a151573b;
    5'b01101 : xpb = 1024'hbf7b4b0f8cd298aa16d46702b43a7ad16a0649de21674641ad14b2b587680e8f27d19d2a849523515fd0a5997b4469239bde5ce84e0c9f34659b6b89ec602a039576428f357ef321fbfc5b308082a84a4abcf62bd233b610c657693ab272d6e8b1eaf574d1549a60fa4bfacdb6a066e0812591bf35b127d754efd7ba35a95f7;
    5'b01110 : xpb = 1024'haff978befa079889b8049317eeeaf6680af247eacc37d663f385c0f3f0d0dbc72f8e8fa12110086e0d401e2bc40547ce73336b154caad4d5b3b8891dcd97823ca91d616ae3334dd8335caff46e5d806d43d14f94afdcdfb303b3f2c18b8c9f9b862808abe281aae6b49da387f86d653a2a17f2a03c80428c493220132e463b1e;
    5'b01111 : xpb = 1024'ha34df7773953d2c0039667e8a237fdd18dce2806e0e197ec4e5d7d66d628899d695787f6cfb040186524f2b70cf83840488ec875f1c20f6c70781c24c1968d27a49429fe237daf39345f97933bd71224eef1d62e161056f44575dcf4b1c76f365229cfd6c7251399d2d6a0841da09ddcfd43ad42355a156ad6a5c7a6304f79da;
    5'b10000 : xpb = 1024'h96a2762f78a00cf64f283cb95585053b10aa0822f58b5974a93539d9bb803773a320804c7e5077c2bd09c74255eb28b21dea25d696d94a032d37af2bb5959812a00af29163c8109a35627f320950a3dc9a125cc77c43ce358737c727d8023ed11e2b9701abc87c4cf10f9d8042d3d67fd06f67e42e33e84964196f393258b896;
    5'b10001 : xpb = 1024'h89f6f4e7b7ec472c9aba118a08d20ca49385e83f0a351afd040cf64ca0d7e549dce978a22cf0af6d14ee9bcd9ede1923f34583373bf08499e9f74232a994a2fd9b81bb24a41271fb366566d0d6ca35944532e360e2774576c8f9b15afe3d0e6bea2d5e2c906be5000f489a7c68070f22a39b2286270dbb27f18d16cc3461f752;
    5'b10010 : xpb = 1024'h7d4b739ff7388162e64be65abc1f140e1661c85b1ededc855ee4b2bf862f932016b270f7db90e7176cd37058e7d10995c8a0e097e107bf30a6b6d5399d93ade896f883b7e45cd35c37684e6fa443c74bf05369fa48aabcb80abb9b8e2477de06b62f2557750f4db32d8197788d3a47c576c6dd281fe78e067f00be5f366b360e;
    5'b10011 : xpb = 1024'h709ff2583684bb9931ddbb2b6f6c1b77993da87733889e0db9bc6f326b8740f6507b694d8a311ec1c4b844e430c3fa079dfc3df8861ef9c7637668409192b8d3926f4c4b24a734bd386b360e71bd59039b73f093aede33f94c7d85c14ab2ada18230ec8259b2b6664bba9474b26d806849f297ca18c160e50c7465f2387474ca;
    5'b10100 : xpb = 1024'h63f4711075d0f5cf7d6f8ffc22b922e11c19889348325f9614942ba550deeecc8a4461a338d1566c1c9d196f79b6ea7973579b592b36345e2035fb478591c3be8de614de64f1961e396e1dad3f36eabb4694772d1511ab3a8e3f6ff470ed7d3c4e32b3ad3e561f1969f39170d7a0b90b1d1e526c119b33c399e80d853a7db386;
    5'b10101 : xpb = 1024'h5748efc8b51d3005c90164ccd6062a4a9ef568af5cdc211e6f6be81836369ca2c40d59f8e7718e167481edfac2a9daeb48b2f8b9d04d6ef4dcf58e4e7990cea9895cdd71a53bf77f3a71054c0cb07c72f1b4fdc67b45227bd0015a2797284cd71a347ad822f987cc882c8e6cfcd3f1adf04a0d0e0a7506a2275bb5183c86f242;
    5'b10110 : xpb = 1024'h4a9d6e80f4696a3c1493399d895331b421d148cb7185e2a6ca43a48b1b8e4a78fdd6524e9611c5c0cc66c2860b9ccb5d1e0e561a7564a98b99b521556d8fd99484d3a604e58658e03b73eceada2a0e2a9cd5845fe17899bd11c3445abd631c71e6364203079cf07fa6658b6922072a50c375c7b0034ed980b4cf5cab3e9030fe;
    5'b10111 : xpb = 1024'h3df1ed3933b5a47260250e6e3ca0391da4ad28e7862fa42f251b60fe00e5f84f379f4aa444b1fd6b244b9711548fbbcef369b37b1a7be4225674b45c618ee47f804a6e9825d0ba413c76d489a7a39fe247f60af947ac10fe53852e8de39dec0cb238092dec405932c49e8865473a62f396a18251fc28ac5f4243043e40996fba;
    5'b11000 : xpb = 1024'h31466bf17301dea8abb6e33eefed4087278909039ad965b77ff31d70e63da625716842f9f35235157c306b9c9d82ac40c8c510dbbf931eb913344763558def6a7bc1372b661b1ba23d79bc28751d3199f3169192addf883f954718c109d8bba77e39d058d0e3c1e5e2d785616c6d9b9669cd3cf3f5027f3dcfb6abd142a2ae76;
    5'b11001 : xpb = 1024'h249aeaa9b24e18def748b80fa33a47f0aa64e91faf83273fdacad9e3cb9553fbab313b4fa1f26cbfd4154027e6759cb29e206e3c64aa594fcff3da6a498cfa557737ffbea6657d033e7ca3c74296c3519e37182c1412ff80d70902f430138b424a3b9783b5872a990110825d91a0d4393cf8f795eddc521c5d2a536444abed32;
    5'b11010 : xpb = 1024'h17ef6961f19a531542da8ce056874f5a2d40c93bc42ce8c835a29656b0ed01d1e4fa33a55092a46a2bfa14b32f688d24737bcb9d09c193e68cb36d713d8c054072aec851e6afde643f7f8b661010550949579ec57a4676c218caed27564e5add163d5eae9a2a934c1f497f59b6d40cdc1024b237e6b624faea9dfaf746b52bee;
    5'b11011 : xpb = 1024'hb43e81a30e68d4b8e6c61b109d456c3b01ca957d8d6aa50907a52c99644afa81ec32bfaff32dc1483dee93e785b7d9648d728fdaed8ce7d49730078318b102b6e2590e526fa3fc540827304dd89e6c0f478255ee079ee035a8cd75a7c892a77e23f25d97ecdfbff3d827c55dc07457ee3506cd9df8ff7d97811a28a48be6aaa;
    5'b11100 : xpb = 1024'haf45ac283220fc4aa503ae58cd7ba57ea46e8ca4c2f80c50692ec8922e9f0a865bd4a1c977f9924d7b21fd10a4ac7ed2824cae4476a2d95fb6d1d2dd605c8fc7ddeb8e2716d59e6b541f5d4643df3ca9939da590d333925551db53885cee9ca4dd487f2e143a5d3fe27b6030f90aa44b0556065e28b527e84bf4c521d3aa0fd1;
    5'b11101 : xpb = 1024'ha29a2ae0716d3680f095832980c8ace8274a6cc0d7a1cdd8c406850513f6b85c959d9a1f2699c9f7d306d19bed9f6f4457a80ba51bba13f6739165e4545b9ab2d96256ba571fffcc552244e51158ce613ebe2c2a39670996939d3dbb83296c3fa94a4658f8ddc5f300b45d2d1e3ddcedd881c100218efac6d9686cb4d5b34e8d;
    5'b11110 : xpb = 1024'h95eea998b0b970b73c2757fa3415b451aa264cdcec4b8f611ede4177f94e6632cf669274d53a01a22aeba62736925fb62d036905c0d14e8d3050f8eb485aa59dd4d91f4d976a612d56252c83ded26018e9deb2c39f9a80d7d55f27eea9643bda754c0d83dd812ea61eed5a2943711590abad7ba21a68cda566dc1447d7bc8d49;
    5'b11111 : xpb = 1024'h89432850f005aaed87b92ccae762bbbb2d022cf900f550e979b5fdeadea61409092f8aca83da394c82d07ab27f855028025ec66665e88923ed108bf23c59b088d04fe7e0d7b4c28e57281422ac4bf1d094ff395d05cdf81917211221cf9f0b75414dd4aec22497593d26572568a44e337ed936441342a083f44fbbdad9c5cc05;
    endcase
end

endmodule

module xpb_5_540
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'ha7b334298820e6a3487245609c72617693f62fc29bd2cf4b558b8484bf2ed0172de1a80a5e310580a1cf109a54c0888a64b5c6951baef87df745a080233c7dc3bf7924afede7608fd858aa3d2acaeba77cc9556985fd50963b8ca4e6e78ac7cb77e2c3ddcd45a73252a32d3df65dee44e986641b6b5d210fc628eb819a47fa52;
    5'b00010 : xpb = 1024'h9eb922fd4e53987dc5df12ea288a7b9bb6765c54622dfe1f2d3a4fb3cb5af326587ad29bf23b8c72a43fe1edc623004a6551654414ab20b03dec01a20ba686d60aa314b12c3dc3da9e1751d7bcba131e058db13a7f74741bc18cb7d314eaed04c0bdf591e9c255d71e86739cf4ebb6608432e954866ee4ef45e25bfeabad8e39;
    5'b00011 : xpb = 1024'h95bf11d114864a58434be073b4a295c0d8f688e628892cf304e91ae2d78716358313fd2d86461364a6b0b3413785780a65ed03f30da748e2849262c3f4108fe855cd04b26a94272563d5f9724ea93a948e520d0b78eb97a1478ccabf424b123e09992746063f047bea69b9fbf3797e7c1edf6e8da180a8cec59bcc7bbd132220;
    5'b00100 : xpb = 1024'h8cc500a4dab8fc32c0b8adfd40baafe5fb76b577eee45bc6dc97e611e3b33944adad27bf1a509a56a9218494a8e7efca6688a2a206a37114cb38c3e5dc7a98faa0f6f4b3a8ea8a702994a10ce098620b171668dc7262bb26cd8cddab6fab3777527458fa22bbb320b64d005af2074697b98bf3c6bc926cae45553cf8ce78b607;
    5'b00101 : xpb = 1024'h83caef78a0ebae0d3e257b86ccd2ca0b1df6e209b53f8a9ab446b140efdf5c53d8465250ae5b2148ab9255e81a4a678a67244150ff9f994711df2507c4e4a20cec20e4b4e740edbaef5348a7728789819fdac4ad6bd9deac538cf0979d0b5cb09b4f8aae3f3861c5823046b9f0950eb3543878ffd7a4308dc50ead75dfde49ee;
    5'b00110 : xpb = 1024'h7ad0de4c671e5fe7bb92491058eae43040770e9b7b9ab96e8bf57c6ffc0b7f6302df7ce24265a83aae03273b8bacdf4a67bfdffff89bc17958858629ad4eab1f374ad4b625975105b511f0420476b0f8289f207e65510231d98d0383ca6b81e9e42abc625bb5106a4e138d18ef22d6ceeee4fe38f2b5f46d44c81df2f143ddd5;
    5'b00111 : xpb = 1024'h71d6cd202d5111c238ff1699e502fe5562f73b2d41f5e84263a4479f0837a2722d78a773d6702f2cb073f88efd0f570a685b7eaef197e9ab9f2be74b95b8b4318274c4b763edb4507ad097dc9665d86eb1637c4f5ec825b75f8d166ff7cba7232d05ee167831bf0f19f6d377edb09eea899183720dc7b84cc4818e7002a971bc;
    5'b01000 : xpb = 1024'h68dcbbf3f383c39cb66be423711b187a857767bf085117163b5312ce1463c5815811d2056a7ab61eb2e4c9e26e71ceca68f71d5dea9411dde5d2486d7e22bd43cd9eb4b8a244179b408f3f772854ffe53a27d820583f493ce58d295c252bcc5c75e11fca94ae6db3e5da19d6ec3e6706243e08ab28d97c2c443afeed140f05a3;
    5'b01001 : xpb = 1024'h5fe2aac7b9b6757733d8b1acfd33329fa7f79450ceac45ea1301ddfd208fe89082aafc96fe853d10b5559b35dfd4468a6992bc0ce3903a102c78a98f668cc65618c8a4b9e09a7ae6064de711ba44275bc2ec33f151b66cc26b8d3c48528bf195bebc517eb12b1c58b1bd6035eacc2f21beea8de443eb400bc3f46f6a2574998a;
    5'b01010 : xpb = 1024'h56e8999b7fe92751b1457f36894b4cc4ca77c0e2950774bdeab0a92c2cbc0b9fad442728928fc402b7c66c895136be4a6a2e5abbdc8c6242731f0ab14ef6cf6863f294bb1ef0de30cc0c8eac4c334ed24bb08fc24b2d9047f18d4f347fec16cf07978332cda7cafd7da0a694e959f73d5997131d5efd03eb43addfe736da2d71;
    5'b01011 : xpb = 1024'h4dee886f461bd92c2eb24cc0156366e9ecf7ed745b62a391c25f745b38e82eaed7dd51ba269a4af4ba373ddcc299360a6ac9f96ad5888a74b9c56bd33760d87aaf1c84bc5d47417b91cb3646de227648d474eb9344a4b3cd778d6220ad4c3c085072b4e6ea2479a24983ecf3e7e7bf58f44398567a0ec7cac3675064483fc158;
    5'b01100 : xpb = 1024'h44f477430c4e8b06ac1f1a49a17b810f0f781a0621bdd2659a0e3f8a451451be02767c4bbaa4d1e6bca80f3033fbadca6b659819ce84b2a7006bccf51fcae18cfa4674bd9b9da4c65789dde170119dbf5d3947643e1bd752fd8d750cdaac6141994de69b06a1284715673352e67587748ef01d8f95208baa4320c0e159a5553f;
    5'b01101 : xpb = 1024'h3bfa6616d2813ce1298be7d32d939b3431f84697e819013971bd0ab9514074cd2d0fa6dd4eaf58d8bf18e083a55e258a6c0136c8c780dad947122e170834ea9f457064bed9f408111d48857c0200c535e5fda3353792fad8838d87f9080c867ae229184f231dd6ebe14a79b1e5034f90299ca2c8b0324f89c2da315e6b0ae926;
    5'b01110 : xpb = 1024'h330054ea98b3eebba6f8b55cb9abb55954787329ae74300d496bd5e85d6c97dc57a8d16ee2b9dfcac189b1d716c09d4a6c9cd577c07d030b8db88f38f09ef3b1909a54c0184a6b5be3072d1693efecac6ec1ff06310a1e5e098d9ae5356cabb42b044a033f9a8590ad2dc010e39117abc4492801cb4413694293a1db7c707d0d;
    5'b01111 : xpb = 1024'h2a0643be5ee6a096246582e645c3cf7e76f89fbb74cf5ee1211aa1176998baeb8241fc0076c466bcc3fa832a8823150a6d387426b9792b3dd45ef05ad908fcc3dbc444c156a0cea6a8c5d4b125df1422f7865ad72a8141e38f8dadd162ccd0ed73df7bb75c1734357911066fe21edfc75ef5ad3ae655d748c24d12588dd610f4;
    5'b10000 : xpb = 1024'h210c329225195270a1d2506fd1dbe9a39978cc4d3b2a8db4f8c96c4675c4ddfaacdb26920aceedaec66b547df9858cca6dd412d5b27553701b05517cc17305d626ee34c294f731f16e847c4bb7ce3b99804ab6a823f86569158dc0bd902cf626bcbaad6b7893e2da44f44ccee0aca7e2f9a2327401679b28420682d59f3ba4db;
    5'b10001 : xpb = 1024'h18122165eb4c044b1f3f1df95df403c8bbf8f8df0185bc88d078377581f10109d77451239ed974a0c8dc25d16ae8048a6e6fb184ab717ba261abb29ea9dd0ee8721824c3d34d953c344323e649bd6310090f12791d6f88ee9b8dd3a9bd8d1b600595df1f9510917f10d7932ddf3a6ffe944eb7ad1c795f07c1bff352b0a138c2;
    5'b10010 : xpb = 1024'hf181039b17eb6259cabeb82ea0c1dedde792570c7e0eb5ca82702a48e1d2419020d7bb532e3fb92cb4cf724dc4a7c4a6f0b5033a46da3d4a85213c0924717fabd4214c511a3f886fa01cb80dbac8a8691d36e4a16e6ac74218de695eaed40994e7110d3b18d4023dcbad98cddc8381a2efb3ce6378b22e7417963cfc206cca9;
    5'b10011 : xpb = 1024'h61dff0d77b168001a18b90c7624381300f952028e3c1a307fd5cdd39a4947282ca6a646c6ee8284cdbdc8784dacf40a6fa6eee29d69cc06eef874e27ab1210d086c04c64ffa5bd1bfc0731b6d9bb1fd1a97ca1b105dcff9a78df982184d65d2974c4287ce09eec8a89e1febdc560035c9a7c21f529ce6c6c132d44cd36c6090;
    5'b10100 : xpb = 1024'hadd13336ffd24ea3628afe6d1296998994ef81c52a0ee97bd56152585978173f5a884e51251f88056f8cd912a26d7c94d45cb577b918c484e63e15629ded9ed0c7e529763de1bc6198191d5898669da497611f84965b208fe31a9e68ffd82d9e0f2f06659b4f95fafb414d29d2b3ee7ab32e263abdfa07d6875bbfce6db45ae2;
    5'b10101 : xpb = 1024'ha4d7220ac605007ddff7cbf69eaeb3aeb76fae56f06a184fad101d8765a43a4e852178e2b92a0ef771fdaa6613cff454d4f85426b214ecb72ce476848657a7e3130f19777c381fac5dd7c4f32a55c51b20257b558fd24415691ab1552d3852d7580a3819b7cc449fc7249388d141b6964ddaab73d90bcbb60715304b7f19eec9;
    5'b10110 : xpb = 1024'h9bdd10de8c37b2585d6499802ac6cdd3d9efdae8b6c5472384bee8b671d05d5dafbaa3744d3495e9746e7bb985326c14d593f2d5ab1114e9738ad7a66ec1b0f55e390978ba8e82f723966c8dbc44ec91a8e9d7268949679aef1ac4415a987810a0e569cdd448f3449307d9e7cfcf7eb1e88730acf41d8f9586cea0c8907f82b0;
    5'b10111 : xpb = 1024'h92e2ffb2526a6432dad16709b6dee7f8fc70077a7d2075f75c6db3e57dfc806cda53ce05e13f1cdb76df4d0cf694e3d4d62f9184a40d3d1bba3138c8572bba07a962f979f8e4e641e95514284e34140831ae32f782c08b20751ad72d87f89d49e9c09b81f0c5a1e95eeb2046ce5d46cd8333b5e60f2f537506881145a1e51697;
    5'b11000 : xpb = 1024'h89e8ee86189d160d583e349342f7021e1ef0340c437ba4cb341c7f148a28a37c04ecf8977549a3cd79501e6067f75b94d6cb30339d09654e00d799ea3f95c319f48ce97b373b498caf13bbc2e0233b7eba728ec87c37aea5fb1aea19b558c283329bcd360d42508e2ace66a5cceb0ee91de03b1f2a411754864181c2b34aaa7e;
    5'b11001 : xpb = 1024'h80eedd59decfc7e7d5ab021ccf0f1c434170609e09d6d39f0bcb4a439654c68b2f86232909542abf7bc0efb3d959d354d766cee296058d80477dfb0c27ffcc2c3fb6d97c7591acd774d2635d721262f54336ea9975aed22b811afd05e2b8e7bc7b76feea29beff32f6b1ad04cb78d704b88cc0584552db3405faf23fc4b03e65;
    5'b11010 : xpb = 1024'h77f4cc2da50279c25317cfa65b27366863f08d2fd0320272e37a1572a280e99a5a1f4dba9d5eb1b17e31c1074abc4b14d8026d918f01b5b28e245c2e1069d53e8ae0c97db3e810223a910af804018a6bcbfb466a6f25f5b1071b0ff210190cf5c452309e463badd7c294f363ca069f205339459160649f1385b462bcd615d24c;
    5'b11011 : xpb = 1024'h6efabb016b352b9cd0849d2fe73f508d8670b9c1968d3146bb28e0a1aead0ca984b8784c316938a380a2925abc1ec2d4d89e0c4087fddde4d4cabd4ff8d3de50d60ab97ef23e736d004fb29295f0b1e254bfa23b689d19368d1b22de3d79322f0d2d625262b85c7c8e7839c2c894673bede5caca7b7662f3056dd339e77b6633;
    5'b11100 : xpb = 1024'h6600a9d53167dd774df16ab973576ab2a8f0e6535ce8601a92d7abd0bad92fb8af51a2ddc573bf95831363ae2d813a94d939aaef80fa06171b711e71e13de7632134a9803094d6b7c60e5a2d27dfd958dd83fe0c62143cbc131b35ca6ad95768560894067f350b215a5b8021c7222f5788925003968826d2852743b6f8e0fa1a;
    5'b11101 : xpb = 1024'h5d0698a8f79a8f51cb5e3842ff6f84d7cb7112e523438eee6a8676ffc70552c7d9eacd6f597e4687858435019ee3b254d9d5499e79f62e4962177f93c9a7f0756c5e99816eeb3a028bcd01c7b9cf00cf664859dd5b8b6041991b48b698397ca19ee3c5ba9bb1b9c6263ec680c5aff773233ed53cb199eab204e0b4340a468e01;
    5'b11110 : xpb = 1024'h540c877cbdcd412c48cb05cc8b879efcedf13f76e99ebdc24235422ed33175d70483f800ed88cd7987f5065510462a14da70e84d72f2567ba8bde0b5b211f987b7888982ad419d4d518ba9624bbe2845ef0cb5ae550283c71f1b5ba2c599a1dae7bef76eb82e686af2220cdfc43dbf8ebdeb5a75ccabae91849a24b11bac21e8;
    5'b11111 : xpb = 1024'h4b12765083fff306c637d356179fb92210716c08aff9ec9619e40d5ddf5d98e62f1d22928193546b8a65d7a881a8a1d4db0c86fc6bee7eadef6441d79a7c029a02b27983eb980098174a50fcddad4fbc77d1117f4e79a74ca51b6e8ef2f9c714309a2922d4ab170fbe05533ec2cb87aa5897dfaee7bd72710453952e2d11b5cf;
    endcase
end

endmodule

module compressor_array_3_2_1024
(
    input  [2:0] col_in_0,
    input  [2:0] col_in_1,
    input  [2:0] col_in_2,
    input  [2:0] col_in_3,
    input  [2:0] col_in_4,
    input  [2:0] col_in_5,
    input  [2:0] col_in_6,
    input  [2:0] col_in_7,
    input  [2:0] col_in_8,
    input  [2:0] col_in_9,
    input  [2:0] col_in_10,
    input  [2:0] col_in_11,
    input  [2:0] col_in_12,
    input  [2:0] col_in_13,
    input  [2:0] col_in_14,
    input  [2:0] col_in_15,
    input  [2:0] col_in_16,
    input  [2:0] col_in_17,
    input  [2:0] col_in_18,
    input  [2:0] col_in_19,
    input  [2:0] col_in_20,
    input  [2:0] col_in_21,
    input  [2:0] col_in_22,
    input  [2:0] col_in_23,
    input  [2:0] col_in_24,
    input  [2:0] col_in_25,
    input  [2:0] col_in_26,
    input  [2:0] col_in_27,
    input  [2:0] col_in_28,
    input  [2:0] col_in_29,
    input  [2:0] col_in_30,
    input  [2:0] col_in_31,
    input  [2:0] col_in_32,
    input  [2:0] col_in_33,
    input  [2:0] col_in_34,
    input  [2:0] col_in_35,
    input  [2:0] col_in_36,
    input  [2:0] col_in_37,
    input  [2:0] col_in_38,
    input  [2:0] col_in_39,
    input  [2:0] col_in_40,
    input  [2:0] col_in_41,
    input  [2:0] col_in_42,
    input  [2:0] col_in_43,
    input  [2:0] col_in_44,
    input  [2:0] col_in_45,
    input  [2:0] col_in_46,
    input  [2:0] col_in_47,
    input  [2:0] col_in_48,
    input  [2:0] col_in_49,
    input  [2:0] col_in_50,
    input  [2:0] col_in_51,
    input  [2:0] col_in_52,
    input  [2:0] col_in_53,
    input  [2:0] col_in_54,
    input  [2:0] col_in_55,
    input  [2:0] col_in_56,
    input  [2:0] col_in_57,
    input  [2:0] col_in_58,
    input  [2:0] col_in_59,
    input  [2:0] col_in_60,
    input  [2:0] col_in_61,
    input  [2:0] col_in_62,
    input  [2:0] col_in_63,
    input  [2:0] col_in_64,
    input  [2:0] col_in_65,
    input  [2:0] col_in_66,
    input  [2:0] col_in_67,
    input  [2:0] col_in_68,
    input  [2:0] col_in_69,
    input  [2:0] col_in_70,
    input  [2:0] col_in_71,
    input  [2:0] col_in_72,
    input  [2:0] col_in_73,
    input  [2:0] col_in_74,
    input  [2:0] col_in_75,
    input  [2:0] col_in_76,
    input  [2:0] col_in_77,
    input  [2:0] col_in_78,
    input  [2:0] col_in_79,
    input  [2:0] col_in_80,
    input  [2:0] col_in_81,
    input  [2:0] col_in_82,
    input  [2:0] col_in_83,
    input  [2:0] col_in_84,
    input  [2:0] col_in_85,
    input  [2:0] col_in_86,
    input  [2:0] col_in_87,
    input  [2:0] col_in_88,
    input  [2:0] col_in_89,
    input  [2:0] col_in_90,
    input  [2:0] col_in_91,
    input  [2:0] col_in_92,
    input  [2:0] col_in_93,
    input  [2:0] col_in_94,
    input  [2:0] col_in_95,
    input  [2:0] col_in_96,
    input  [2:0] col_in_97,
    input  [2:0] col_in_98,
    input  [2:0] col_in_99,
    input  [2:0] col_in_100,
    input  [2:0] col_in_101,
    input  [2:0] col_in_102,
    input  [2:0] col_in_103,
    input  [2:0] col_in_104,
    input  [2:0] col_in_105,
    input  [2:0] col_in_106,
    input  [2:0] col_in_107,
    input  [2:0] col_in_108,
    input  [2:0] col_in_109,
    input  [2:0] col_in_110,
    input  [2:0] col_in_111,
    input  [2:0] col_in_112,
    input  [2:0] col_in_113,
    input  [2:0] col_in_114,
    input  [2:0] col_in_115,
    input  [2:0] col_in_116,
    input  [2:0] col_in_117,
    input  [2:0] col_in_118,
    input  [2:0] col_in_119,
    input  [2:0] col_in_120,
    input  [2:0] col_in_121,
    input  [2:0] col_in_122,
    input  [2:0] col_in_123,
    input  [2:0] col_in_124,
    input  [2:0] col_in_125,
    input  [2:0] col_in_126,
    input  [2:0] col_in_127,
    input  [2:0] col_in_128,
    input  [2:0] col_in_129,
    input  [2:0] col_in_130,
    input  [2:0] col_in_131,
    input  [2:0] col_in_132,
    input  [2:0] col_in_133,
    input  [2:0] col_in_134,
    input  [2:0] col_in_135,
    input  [2:0] col_in_136,
    input  [2:0] col_in_137,
    input  [2:0] col_in_138,
    input  [2:0] col_in_139,
    input  [2:0] col_in_140,
    input  [2:0] col_in_141,
    input  [2:0] col_in_142,
    input  [2:0] col_in_143,
    input  [2:0] col_in_144,
    input  [2:0] col_in_145,
    input  [2:0] col_in_146,
    input  [2:0] col_in_147,
    input  [2:0] col_in_148,
    input  [2:0] col_in_149,
    input  [2:0] col_in_150,
    input  [2:0] col_in_151,
    input  [2:0] col_in_152,
    input  [2:0] col_in_153,
    input  [2:0] col_in_154,
    input  [2:0] col_in_155,
    input  [2:0] col_in_156,
    input  [2:0] col_in_157,
    input  [2:0] col_in_158,
    input  [2:0] col_in_159,
    input  [2:0] col_in_160,
    input  [2:0] col_in_161,
    input  [2:0] col_in_162,
    input  [2:0] col_in_163,
    input  [2:0] col_in_164,
    input  [2:0] col_in_165,
    input  [2:0] col_in_166,
    input  [2:0] col_in_167,
    input  [2:0] col_in_168,
    input  [2:0] col_in_169,
    input  [2:0] col_in_170,
    input  [2:0] col_in_171,
    input  [2:0] col_in_172,
    input  [2:0] col_in_173,
    input  [2:0] col_in_174,
    input  [2:0] col_in_175,
    input  [2:0] col_in_176,
    input  [2:0] col_in_177,
    input  [2:0] col_in_178,
    input  [2:0] col_in_179,
    input  [2:0] col_in_180,
    input  [2:0] col_in_181,
    input  [2:0] col_in_182,
    input  [2:0] col_in_183,
    input  [2:0] col_in_184,
    input  [2:0] col_in_185,
    input  [2:0] col_in_186,
    input  [2:0] col_in_187,
    input  [2:0] col_in_188,
    input  [2:0] col_in_189,
    input  [2:0] col_in_190,
    input  [2:0] col_in_191,
    input  [2:0] col_in_192,
    input  [2:0] col_in_193,
    input  [2:0] col_in_194,
    input  [2:0] col_in_195,
    input  [2:0] col_in_196,
    input  [2:0] col_in_197,
    input  [2:0] col_in_198,
    input  [2:0] col_in_199,
    input  [2:0] col_in_200,
    input  [2:0] col_in_201,
    input  [2:0] col_in_202,
    input  [2:0] col_in_203,
    input  [2:0] col_in_204,
    input  [2:0] col_in_205,
    input  [2:0] col_in_206,
    input  [2:0] col_in_207,
    input  [2:0] col_in_208,
    input  [2:0] col_in_209,
    input  [2:0] col_in_210,
    input  [2:0] col_in_211,
    input  [2:0] col_in_212,
    input  [2:0] col_in_213,
    input  [2:0] col_in_214,
    input  [2:0] col_in_215,
    input  [2:0] col_in_216,
    input  [2:0] col_in_217,
    input  [2:0] col_in_218,
    input  [2:0] col_in_219,
    input  [2:0] col_in_220,
    input  [2:0] col_in_221,
    input  [2:0] col_in_222,
    input  [2:0] col_in_223,
    input  [2:0] col_in_224,
    input  [2:0] col_in_225,
    input  [2:0] col_in_226,
    input  [2:0] col_in_227,
    input  [2:0] col_in_228,
    input  [2:0] col_in_229,
    input  [2:0] col_in_230,
    input  [2:0] col_in_231,
    input  [2:0] col_in_232,
    input  [2:0] col_in_233,
    input  [2:0] col_in_234,
    input  [2:0] col_in_235,
    input  [2:0] col_in_236,
    input  [2:0] col_in_237,
    input  [2:0] col_in_238,
    input  [2:0] col_in_239,
    input  [2:0] col_in_240,
    input  [2:0] col_in_241,
    input  [2:0] col_in_242,
    input  [2:0] col_in_243,
    input  [2:0] col_in_244,
    input  [2:0] col_in_245,
    input  [2:0] col_in_246,
    input  [2:0] col_in_247,
    input  [2:0] col_in_248,
    input  [2:0] col_in_249,
    input  [2:0] col_in_250,
    input  [2:0] col_in_251,
    input  [2:0] col_in_252,
    input  [2:0] col_in_253,
    input  [2:0] col_in_254,
    input  [2:0] col_in_255,
    input  [2:0] col_in_256,
    input  [2:0] col_in_257,
    input  [2:0] col_in_258,
    input  [2:0] col_in_259,
    input  [2:0] col_in_260,
    input  [2:0] col_in_261,
    input  [2:0] col_in_262,
    input  [2:0] col_in_263,
    input  [2:0] col_in_264,
    input  [2:0] col_in_265,
    input  [2:0] col_in_266,
    input  [2:0] col_in_267,
    input  [2:0] col_in_268,
    input  [2:0] col_in_269,
    input  [2:0] col_in_270,
    input  [2:0] col_in_271,
    input  [2:0] col_in_272,
    input  [2:0] col_in_273,
    input  [2:0] col_in_274,
    input  [2:0] col_in_275,
    input  [2:0] col_in_276,
    input  [2:0] col_in_277,
    input  [2:0] col_in_278,
    input  [2:0] col_in_279,
    input  [2:0] col_in_280,
    input  [2:0] col_in_281,
    input  [2:0] col_in_282,
    input  [2:0] col_in_283,
    input  [2:0] col_in_284,
    input  [2:0] col_in_285,
    input  [2:0] col_in_286,
    input  [2:0] col_in_287,
    input  [2:0] col_in_288,
    input  [2:0] col_in_289,
    input  [2:0] col_in_290,
    input  [2:0] col_in_291,
    input  [2:0] col_in_292,
    input  [2:0] col_in_293,
    input  [2:0] col_in_294,
    input  [2:0] col_in_295,
    input  [2:0] col_in_296,
    input  [2:0] col_in_297,
    input  [2:0] col_in_298,
    input  [2:0] col_in_299,
    input  [2:0] col_in_300,
    input  [2:0] col_in_301,
    input  [2:0] col_in_302,
    input  [2:0] col_in_303,
    input  [2:0] col_in_304,
    input  [2:0] col_in_305,
    input  [2:0] col_in_306,
    input  [2:0] col_in_307,
    input  [2:0] col_in_308,
    input  [2:0] col_in_309,
    input  [2:0] col_in_310,
    input  [2:0] col_in_311,
    input  [2:0] col_in_312,
    input  [2:0] col_in_313,
    input  [2:0] col_in_314,
    input  [2:0] col_in_315,
    input  [2:0] col_in_316,
    input  [2:0] col_in_317,
    input  [2:0] col_in_318,
    input  [2:0] col_in_319,
    input  [2:0] col_in_320,
    input  [2:0] col_in_321,
    input  [2:0] col_in_322,
    input  [2:0] col_in_323,
    input  [2:0] col_in_324,
    input  [2:0] col_in_325,
    input  [2:0] col_in_326,
    input  [2:0] col_in_327,
    input  [2:0] col_in_328,
    input  [2:0] col_in_329,
    input  [2:0] col_in_330,
    input  [2:0] col_in_331,
    input  [2:0] col_in_332,
    input  [2:0] col_in_333,
    input  [2:0] col_in_334,
    input  [2:0] col_in_335,
    input  [2:0] col_in_336,
    input  [2:0] col_in_337,
    input  [2:0] col_in_338,
    input  [2:0] col_in_339,
    input  [2:0] col_in_340,
    input  [2:0] col_in_341,
    input  [2:0] col_in_342,
    input  [2:0] col_in_343,
    input  [2:0] col_in_344,
    input  [2:0] col_in_345,
    input  [2:0] col_in_346,
    input  [2:0] col_in_347,
    input  [2:0] col_in_348,
    input  [2:0] col_in_349,
    input  [2:0] col_in_350,
    input  [2:0] col_in_351,
    input  [2:0] col_in_352,
    input  [2:0] col_in_353,
    input  [2:0] col_in_354,
    input  [2:0] col_in_355,
    input  [2:0] col_in_356,
    input  [2:0] col_in_357,
    input  [2:0] col_in_358,
    input  [2:0] col_in_359,
    input  [2:0] col_in_360,
    input  [2:0] col_in_361,
    input  [2:0] col_in_362,
    input  [2:0] col_in_363,
    input  [2:0] col_in_364,
    input  [2:0] col_in_365,
    input  [2:0] col_in_366,
    input  [2:0] col_in_367,
    input  [2:0] col_in_368,
    input  [2:0] col_in_369,
    input  [2:0] col_in_370,
    input  [2:0] col_in_371,
    input  [2:0] col_in_372,
    input  [2:0] col_in_373,
    input  [2:0] col_in_374,
    input  [2:0] col_in_375,
    input  [2:0] col_in_376,
    input  [2:0] col_in_377,
    input  [2:0] col_in_378,
    input  [2:0] col_in_379,
    input  [2:0] col_in_380,
    input  [2:0] col_in_381,
    input  [2:0] col_in_382,
    input  [2:0] col_in_383,
    input  [2:0] col_in_384,
    input  [2:0] col_in_385,
    input  [2:0] col_in_386,
    input  [2:0] col_in_387,
    input  [2:0] col_in_388,
    input  [2:0] col_in_389,
    input  [2:0] col_in_390,
    input  [2:0] col_in_391,
    input  [2:0] col_in_392,
    input  [2:0] col_in_393,
    input  [2:0] col_in_394,
    input  [2:0] col_in_395,
    input  [2:0] col_in_396,
    input  [2:0] col_in_397,
    input  [2:0] col_in_398,
    input  [2:0] col_in_399,
    input  [2:0] col_in_400,
    input  [2:0] col_in_401,
    input  [2:0] col_in_402,
    input  [2:0] col_in_403,
    input  [2:0] col_in_404,
    input  [2:0] col_in_405,
    input  [2:0] col_in_406,
    input  [2:0] col_in_407,
    input  [2:0] col_in_408,
    input  [2:0] col_in_409,
    input  [2:0] col_in_410,
    input  [2:0] col_in_411,
    input  [2:0] col_in_412,
    input  [2:0] col_in_413,
    input  [2:0] col_in_414,
    input  [2:0] col_in_415,
    input  [2:0] col_in_416,
    input  [2:0] col_in_417,
    input  [2:0] col_in_418,
    input  [2:0] col_in_419,
    input  [2:0] col_in_420,
    input  [2:0] col_in_421,
    input  [2:0] col_in_422,
    input  [2:0] col_in_423,
    input  [2:0] col_in_424,
    input  [2:0] col_in_425,
    input  [2:0] col_in_426,
    input  [2:0] col_in_427,
    input  [2:0] col_in_428,
    input  [2:0] col_in_429,
    input  [2:0] col_in_430,
    input  [2:0] col_in_431,
    input  [2:0] col_in_432,
    input  [2:0] col_in_433,
    input  [2:0] col_in_434,
    input  [2:0] col_in_435,
    input  [2:0] col_in_436,
    input  [2:0] col_in_437,
    input  [2:0] col_in_438,
    input  [2:0] col_in_439,
    input  [2:0] col_in_440,
    input  [2:0] col_in_441,
    input  [2:0] col_in_442,
    input  [2:0] col_in_443,
    input  [2:0] col_in_444,
    input  [2:0] col_in_445,
    input  [2:0] col_in_446,
    input  [2:0] col_in_447,
    input  [2:0] col_in_448,
    input  [2:0] col_in_449,
    input  [2:0] col_in_450,
    input  [2:0] col_in_451,
    input  [2:0] col_in_452,
    input  [2:0] col_in_453,
    input  [2:0] col_in_454,
    input  [2:0] col_in_455,
    input  [2:0] col_in_456,
    input  [2:0] col_in_457,
    input  [2:0] col_in_458,
    input  [2:0] col_in_459,
    input  [2:0] col_in_460,
    input  [2:0] col_in_461,
    input  [2:0] col_in_462,
    input  [2:0] col_in_463,
    input  [2:0] col_in_464,
    input  [2:0] col_in_465,
    input  [2:0] col_in_466,
    input  [2:0] col_in_467,
    input  [2:0] col_in_468,
    input  [2:0] col_in_469,
    input  [2:0] col_in_470,
    input  [2:0] col_in_471,
    input  [2:0] col_in_472,
    input  [2:0] col_in_473,
    input  [2:0] col_in_474,
    input  [2:0] col_in_475,
    input  [2:0] col_in_476,
    input  [2:0] col_in_477,
    input  [2:0] col_in_478,
    input  [2:0] col_in_479,
    input  [2:0] col_in_480,
    input  [2:0] col_in_481,
    input  [2:0] col_in_482,
    input  [2:0] col_in_483,
    input  [2:0] col_in_484,
    input  [2:0] col_in_485,
    input  [2:0] col_in_486,
    input  [2:0] col_in_487,
    input  [2:0] col_in_488,
    input  [2:0] col_in_489,
    input  [2:0] col_in_490,
    input  [2:0] col_in_491,
    input  [2:0] col_in_492,
    input  [2:0] col_in_493,
    input  [2:0] col_in_494,
    input  [2:0] col_in_495,
    input  [2:0] col_in_496,
    input  [2:0] col_in_497,
    input  [2:0] col_in_498,
    input  [2:0] col_in_499,
    input  [2:0] col_in_500,
    input  [2:0] col_in_501,
    input  [2:0] col_in_502,
    input  [2:0] col_in_503,
    input  [2:0] col_in_504,
    input  [2:0] col_in_505,
    input  [2:0] col_in_506,
    input  [2:0] col_in_507,
    input  [2:0] col_in_508,
    input  [2:0] col_in_509,
    input  [2:0] col_in_510,
    input  [2:0] col_in_511,
    input  [2:0] col_in_512,
    input  [2:0] col_in_513,
    input  [2:0] col_in_514,
    input  [2:0] col_in_515,
    input  [2:0] col_in_516,
    input  [2:0] col_in_517,
    input  [2:0] col_in_518,
    input  [2:0] col_in_519,
    input  [2:0] col_in_520,
    input  [2:0] col_in_521,
    input  [2:0] col_in_522,
    input  [2:0] col_in_523,
    input  [2:0] col_in_524,
    input  [2:0] col_in_525,
    input  [2:0] col_in_526,
    input  [2:0] col_in_527,
    input  [2:0] col_in_528,
    input  [2:0] col_in_529,
    input  [2:0] col_in_530,
    input  [2:0] col_in_531,
    input  [2:0] col_in_532,
    input  [2:0] col_in_533,
    input  [2:0] col_in_534,
    input  [2:0] col_in_535,
    input  [2:0] col_in_536,
    input  [2:0] col_in_537,
    input  [2:0] col_in_538,
    input  [2:0] col_in_539,
    input  [2:0] col_in_540,
    input  [2:0] col_in_541,
    input  [2:0] col_in_542,
    input  [2:0] col_in_543,
    input  [2:0] col_in_544,
    input  [2:0] col_in_545,
    input  [2:0] col_in_546,
    input  [2:0] col_in_547,
    input  [2:0] col_in_548,
    input  [2:0] col_in_549,
    input  [2:0] col_in_550,
    input  [2:0] col_in_551,
    input  [2:0] col_in_552,
    input  [2:0] col_in_553,
    input  [2:0] col_in_554,
    input  [2:0] col_in_555,
    input  [2:0] col_in_556,
    input  [2:0] col_in_557,
    input  [2:0] col_in_558,
    input  [2:0] col_in_559,
    input  [2:0] col_in_560,
    input  [2:0] col_in_561,
    input  [2:0] col_in_562,
    input  [2:0] col_in_563,
    input  [2:0] col_in_564,
    input  [2:0] col_in_565,
    input  [2:0] col_in_566,
    input  [2:0] col_in_567,
    input  [2:0] col_in_568,
    input  [2:0] col_in_569,
    input  [2:0] col_in_570,
    input  [2:0] col_in_571,
    input  [2:0] col_in_572,
    input  [2:0] col_in_573,
    input  [2:0] col_in_574,
    input  [2:0] col_in_575,
    input  [2:0] col_in_576,
    input  [2:0] col_in_577,
    input  [2:0] col_in_578,
    input  [2:0] col_in_579,
    input  [2:0] col_in_580,
    input  [2:0] col_in_581,
    input  [2:0] col_in_582,
    input  [2:0] col_in_583,
    input  [2:0] col_in_584,
    input  [2:0] col_in_585,
    input  [2:0] col_in_586,
    input  [2:0] col_in_587,
    input  [2:0] col_in_588,
    input  [2:0] col_in_589,
    input  [2:0] col_in_590,
    input  [2:0] col_in_591,
    input  [2:0] col_in_592,
    input  [2:0] col_in_593,
    input  [2:0] col_in_594,
    input  [2:0] col_in_595,
    input  [2:0] col_in_596,
    input  [2:0] col_in_597,
    input  [2:0] col_in_598,
    input  [2:0] col_in_599,
    input  [2:0] col_in_600,
    input  [2:0] col_in_601,
    input  [2:0] col_in_602,
    input  [2:0] col_in_603,
    input  [2:0] col_in_604,
    input  [2:0] col_in_605,
    input  [2:0] col_in_606,
    input  [2:0] col_in_607,
    input  [2:0] col_in_608,
    input  [2:0] col_in_609,
    input  [2:0] col_in_610,
    input  [2:0] col_in_611,
    input  [2:0] col_in_612,
    input  [2:0] col_in_613,
    input  [2:0] col_in_614,
    input  [2:0] col_in_615,
    input  [2:0] col_in_616,
    input  [2:0] col_in_617,
    input  [2:0] col_in_618,
    input  [2:0] col_in_619,
    input  [2:0] col_in_620,
    input  [2:0] col_in_621,
    input  [2:0] col_in_622,
    input  [2:0] col_in_623,
    input  [2:0] col_in_624,
    input  [2:0] col_in_625,
    input  [2:0] col_in_626,
    input  [2:0] col_in_627,
    input  [2:0] col_in_628,
    input  [2:0] col_in_629,
    input  [2:0] col_in_630,
    input  [2:0] col_in_631,
    input  [2:0] col_in_632,
    input  [2:0] col_in_633,
    input  [2:0] col_in_634,
    input  [2:0] col_in_635,
    input  [2:0] col_in_636,
    input  [2:0] col_in_637,
    input  [2:0] col_in_638,
    input  [2:0] col_in_639,
    input  [2:0] col_in_640,
    input  [2:0] col_in_641,
    input  [2:0] col_in_642,
    input  [2:0] col_in_643,
    input  [2:0] col_in_644,
    input  [2:0] col_in_645,
    input  [2:0] col_in_646,
    input  [2:0] col_in_647,
    input  [2:0] col_in_648,
    input  [2:0] col_in_649,
    input  [2:0] col_in_650,
    input  [2:0] col_in_651,
    input  [2:0] col_in_652,
    input  [2:0] col_in_653,
    input  [2:0] col_in_654,
    input  [2:0] col_in_655,
    input  [2:0] col_in_656,
    input  [2:0] col_in_657,
    input  [2:0] col_in_658,
    input  [2:0] col_in_659,
    input  [2:0] col_in_660,
    input  [2:0] col_in_661,
    input  [2:0] col_in_662,
    input  [2:0] col_in_663,
    input  [2:0] col_in_664,
    input  [2:0] col_in_665,
    input  [2:0] col_in_666,
    input  [2:0] col_in_667,
    input  [2:0] col_in_668,
    input  [2:0] col_in_669,
    input  [2:0] col_in_670,
    input  [2:0] col_in_671,
    input  [2:0] col_in_672,
    input  [2:0] col_in_673,
    input  [2:0] col_in_674,
    input  [2:0] col_in_675,
    input  [2:0] col_in_676,
    input  [2:0] col_in_677,
    input  [2:0] col_in_678,
    input  [2:0] col_in_679,
    input  [2:0] col_in_680,
    input  [2:0] col_in_681,
    input  [2:0] col_in_682,
    input  [2:0] col_in_683,
    input  [2:0] col_in_684,
    input  [2:0] col_in_685,
    input  [2:0] col_in_686,
    input  [2:0] col_in_687,
    input  [2:0] col_in_688,
    input  [2:0] col_in_689,
    input  [2:0] col_in_690,
    input  [2:0] col_in_691,
    input  [2:0] col_in_692,
    input  [2:0] col_in_693,
    input  [2:0] col_in_694,
    input  [2:0] col_in_695,
    input  [2:0] col_in_696,
    input  [2:0] col_in_697,
    input  [2:0] col_in_698,
    input  [2:0] col_in_699,
    input  [2:0] col_in_700,
    input  [2:0] col_in_701,
    input  [2:0] col_in_702,
    input  [2:0] col_in_703,
    input  [2:0] col_in_704,
    input  [2:0] col_in_705,
    input  [2:0] col_in_706,
    input  [2:0] col_in_707,
    input  [2:0] col_in_708,
    input  [2:0] col_in_709,
    input  [2:0] col_in_710,
    input  [2:0] col_in_711,
    input  [2:0] col_in_712,
    input  [2:0] col_in_713,
    input  [2:0] col_in_714,
    input  [2:0] col_in_715,
    input  [2:0] col_in_716,
    input  [2:0] col_in_717,
    input  [2:0] col_in_718,
    input  [2:0] col_in_719,
    input  [2:0] col_in_720,
    input  [2:0] col_in_721,
    input  [2:0] col_in_722,
    input  [2:0] col_in_723,
    input  [2:0] col_in_724,
    input  [2:0] col_in_725,
    input  [2:0] col_in_726,
    input  [2:0] col_in_727,
    input  [2:0] col_in_728,
    input  [2:0] col_in_729,
    input  [2:0] col_in_730,
    input  [2:0] col_in_731,
    input  [2:0] col_in_732,
    input  [2:0] col_in_733,
    input  [2:0] col_in_734,
    input  [2:0] col_in_735,
    input  [2:0] col_in_736,
    input  [2:0] col_in_737,
    input  [2:0] col_in_738,
    input  [2:0] col_in_739,
    input  [2:0] col_in_740,
    input  [2:0] col_in_741,
    input  [2:0] col_in_742,
    input  [2:0] col_in_743,
    input  [2:0] col_in_744,
    input  [2:0] col_in_745,
    input  [2:0] col_in_746,
    input  [2:0] col_in_747,
    input  [2:0] col_in_748,
    input  [2:0] col_in_749,
    input  [2:0] col_in_750,
    input  [2:0] col_in_751,
    input  [2:0] col_in_752,
    input  [2:0] col_in_753,
    input  [2:0] col_in_754,
    input  [2:0] col_in_755,
    input  [2:0] col_in_756,
    input  [2:0] col_in_757,
    input  [2:0] col_in_758,
    input  [2:0] col_in_759,
    input  [2:0] col_in_760,
    input  [2:0] col_in_761,
    input  [2:0] col_in_762,
    input  [2:0] col_in_763,
    input  [2:0] col_in_764,
    input  [2:0] col_in_765,
    input  [2:0] col_in_766,
    input  [2:0] col_in_767,
    input  [2:0] col_in_768,
    input  [2:0] col_in_769,
    input  [2:0] col_in_770,
    input  [2:0] col_in_771,
    input  [2:0] col_in_772,
    input  [2:0] col_in_773,
    input  [2:0] col_in_774,
    input  [2:0] col_in_775,
    input  [2:0] col_in_776,
    input  [2:0] col_in_777,
    input  [2:0] col_in_778,
    input  [2:0] col_in_779,
    input  [2:0] col_in_780,
    input  [2:0] col_in_781,
    input  [2:0] col_in_782,
    input  [2:0] col_in_783,
    input  [2:0] col_in_784,
    input  [2:0] col_in_785,
    input  [2:0] col_in_786,
    input  [2:0] col_in_787,
    input  [2:0] col_in_788,
    input  [2:0] col_in_789,
    input  [2:0] col_in_790,
    input  [2:0] col_in_791,
    input  [2:0] col_in_792,
    input  [2:0] col_in_793,
    input  [2:0] col_in_794,
    input  [2:0] col_in_795,
    input  [2:0] col_in_796,
    input  [2:0] col_in_797,
    input  [2:0] col_in_798,
    input  [2:0] col_in_799,
    input  [2:0] col_in_800,
    input  [2:0] col_in_801,
    input  [2:0] col_in_802,
    input  [2:0] col_in_803,
    input  [2:0] col_in_804,
    input  [2:0] col_in_805,
    input  [2:0] col_in_806,
    input  [2:0] col_in_807,
    input  [2:0] col_in_808,
    input  [2:0] col_in_809,
    input  [2:0] col_in_810,
    input  [2:0] col_in_811,
    input  [2:0] col_in_812,
    input  [2:0] col_in_813,
    input  [2:0] col_in_814,
    input  [2:0] col_in_815,
    input  [2:0] col_in_816,
    input  [2:0] col_in_817,
    input  [2:0] col_in_818,
    input  [2:0] col_in_819,
    input  [2:0] col_in_820,
    input  [2:0] col_in_821,
    input  [2:0] col_in_822,
    input  [2:0] col_in_823,
    input  [2:0] col_in_824,
    input  [2:0] col_in_825,
    input  [2:0] col_in_826,
    input  [2:0] col_in_827,
    input  [2:0] col_in_828,
    input  [2:0] col_in_829,
    input  [2:0] col_in_830,
    input  [2:0] col_in_831,
    input  [2:0] col_in_832,
    input  [2:0] col_in_833,
    input  [2:0] col_in_834,
    input  [2:0] col_in_835,
    input  [2:0] col_in_836,
    input  [2:0] col_in_837,
    input  [2:0] col_in_838,
    input  [2:0] col_in_839,
    input  [2:0] col_in_840,
    input  [2:0] col_in_841,
    input  [2:0] col_in_842,
    input  [2:0] col_in_843,
    input  [2:0] col_in_844,
    input  [2:0] col_in_845,
    input  [2:0] col_in_846,
    input  [2:0] col_in_847,
    input  [2:0] col_in_848,
    input  [2:0] col_in_849,
    input  [2:0] col_in_850,
    input  [2:0] col_in_851,
    input  [2:0] col_in_852,
    input  [2:0] col_in_853,
    input  [2:0] col_in_854,
    input  [2:0] col_in_855,
    input  [2:0] col_in_856,
    input  [2:0] col_in_857,
    input  [2:0] col_in_858,
    input  [2:0] col_in_859,
    input  [2:0] col_in_860,
    input  [2:0] col_in_861,
    input  [2:0] col_in_862,
    input  [2:0] col_in_863,
    input  [2:0] col_in_864,
    input  [2:0] col_in_865,
    input  [2:0] col_in_866,
    input  [2:0] col_in_867,
    input  [2:0] col_in_868,
    input  [2:0] col_in_869,
    input  [2:0] col_in_870,
    input  [2:0] col_in_871,
    input  [2:0] col_in_872,
    input  [2:0] col_in_873,
    input  [2:0] col_in_874,
    input  [2:0] col_in_875,
    input  [2:0] col_in_876,
    input  [2:0] col_in_877,
    input  [2:0] col_in_878,
    input  [2:0] col_in_879,
    input  [2:0] col_in_880,
    input  [2:0] col_in_881,
    input  [2:0] col_in_882,
    input  [2:0] col_in_883,
    input  [2:0] col_in_884,
    input  [2:0] col_in_885,
    input  [2:0] col_in_886,
    input  [2:0] col_in_887,
    input  [2:0] col_in_888,
    input  [2:0] col_in_889,
    input  [2:0] col_in_890,
    input  [2:0] col_in_891,
    input  [2:0] col_in_892,
    input  [2:0] col_in_893,
    input  [2:0] col_in_894,
    input  [2:0] col_in_895,
    input  [2:0] col_in_896,
    input  [2:0] col_in_897,
    input  [2:0] col_in_898,
    input  [2:0] col_in_899,
    input  [2:0] col_in_900,
    input  [2:0] col_in_901,
    input  [2:0] col_in_902,
    input  [2:0] col_in_903,
    input  [2:0] col_in_904,
    input  [2:0] col_in_905,
    input  [2:0] col_in_906,
    input  [2:0] col_in_907,
    input  [2:0] col_in_908,
    input  [2:0] col_in_909,
    input  [2:0] col_in_910,
    input  [2:0] col_in_911,
    input  [2:0] col_in_912,
    input  [2:0] col_in_913,
    input  [2:0] col_in_914,
    input  [2:0] col_in_915,
    input  [2:0] col_in_916,
    input  [2:0] col_in_917,
    input  [2:0] col_in_918,
    input  [2:0] col_in_919,
    input  [2:0] col_in_920,
    input  [2:0] col_in_921,
    input  [2:0] col_in_922,
    input  [2:0] col_in_923,
    input  [2:0] col_in_924,
    input  [2:0] col_in_925,
    input  [2:0] col_in_926,
    input  [2:0] col_in_927,
    input  [2:0] col_in_928,
    input  [2:0] col_in_929,
    input  [2:0] col_in_930,
    input  [2:0] col_in_931,
    input  [2:0] col_in_932,
    input  [2:0] col_in_933,
    input  [2:0] col_in_934,
    input  [2:0] col_in_935,
    input  [2:0] col_in_936,
    input  [2:0] col_in_937,
    input  [2:0] col_in_938,
    input  [2:0] col_in_939,
    input  [2:0] col_in_940,
    input  [2:0] col_in_941,
    input  [2:0] col_in_942,
    input  [2:0] col_in_943,
    input  [2:0] col_in_944,
    input  [2:0] col_in_945,
    input  [2:0] col_in_946,
    input  [2:0] col_in_947,
    input  [2:0] col_in_948,
    input  [2:0] col_in_949,
    input  [2:0] col_in_950,
    input  [2:0] col_in_951,
    input  [2:0] col_in_952,
    input  [2:0] col_in_953,
    input  [2:0] col_in_954,
    input  [2:0] col_in_955,
    input  [2:0] col_in_956,
    input  [2:0] col_in_957,
    input  [2:0] col_in_958,
    input  [2:0] col_in_959,
    input  [2:0] col_in_960,
    input  [2:0] col_in_961,
    input  [2:0] col_in_962,
    input  [2:0] col_in_963,
    input  [2:0] col_in_964,
    input  [2:0] col_in_965,
    input  [2:0] col_in_966,
    input  [2:0] col_in_967,
    input  [2:0] col_in_968,
    input  [2:0] col_in_969,
    input  [2:0] col_in_970,
    input  [2:0] col_in_971,
    input  [2:0] col_in_972,
    input  [2:0] col_in_973,
    input  [2:0] col_in_974,
    input  [2:0] col_in_975,
    input  [2:0] col_in_976,
    input  [2:0] col_in_977,
    input  [2:0] col_in_978,
    input  [2:0] col_in_979,
    input  [2:0] col_in_980,
    input  [2:0] col_in_981,
    input  [2:0] col_in_982,
    input  [2:0] col_in_983,
    input  [2:0] col_in_984,
    input  [2:0] col_in_985,
    input  [2:0] col_in_986,
    input  [2:0] col_in_987,
    input  [2:0] col_in_988,
    input  [2:0] col_in_989,
    input  [2:0] col_in_990,
    input  [2:0] col_in_991,
    input  [2:0] col_in_992,
    input  [2:0] col_in_993,
    input  [2:0] col_in_994,
    input  [2:0] col_in_995,
    input  [2:0] col_in_996,
    input  [2:0] col_in_997,
    input  [2:0] col_in_998,
    input  [2:0] col_in_999,
    input  [2:0] col_in_1000,
    input  [2:0] col_in_1001,
    input  [2:0] col_in_1002,
    input  [2:0] col_in_1003,
    input  [2:0] col_in_1004,
    input  [2:0] col_in_1005,
    input  [2:0] col_in_1006,
    input  [2:0] col_in_1007,
    input  [2:0] col_in_1008,
    input  [2:0] col_in_1009,
    input  [2:0] col_in_1010,
    input  [2:0] col_in_1011,
    input  [2:0] col_in_1012,
    input  [2:0] col_in_1013,
    input  [2:0] col_in_1014,
    input  [2:0] col_in_1015,
    input  [2:0] col_in_1016,
    input  [2:0] col_in_1017,
    input  [2:0] col_in_1018,
    input  [2:0] col_in_1019,
    input  [2:0] col_in_1020,
    input  [2:0] col_in_1021,
    input  [2:0] col_in_1022,
    input  [2:0] col_in_1023,

    output [1:0] col_out_0,
    output [1:0] col_out_1,
    output [1:0] col_out_2,
    output [1:0] col_out_3,
    output [1:0] col_out_4,
    output [1:0] col_out_5,
    output [1:0] col_out_6,
    output [1:0] col_out_7,
    output [1:0] col_out_8,
    output [1:0] col_out_9,
    output [1:0] col_out_10,
    output [1:0] col_out_11,
    output [1:0] col_out_12,
    output [1:0] col_out_13,
    output [1:0] col_out_14,
    output [1:0] col_out_15,
    output [1:0] col_out_16,
    output [1:0] col_out_17,
    output [1:0] col_out_18,
    output [1:0] col_out_19,
    output [1:0] col_out_20,
    output [1:0] col_out_21,
    output [1:0] col_out_22,
    output [1:0] col_out_23,
    output [1:0] col_out_24,
    output [1:0] col_out_25,
    output [1:0] col_out_26,
    output [1:0] col_out_27,
    output [1:0] col_out_28,
    output [1:0] col_out_29,
    output [1:0] col_out_30,
    output [1:0] col_out_31,
    output [1:0] col_out_32,
    output [1:0] col_out_33,
    output [1:0] col_out_34,
    output [1:0] col_out_35,
    output [1:0] col_out_36,
    output [1:0] col_out_37,
    output [1:0] col_out_38,
    output [1:0] col_out_39,
    output [1:0] col_out_40,
    output [1:0] col_out_41,
    output [1:0] col_out_42,
    output [1:0] col_out_43,
    output [1:0] col_out_44,
    output [1:0] col_out_45,
    output [1:0] col_out_46,
    output [1:0] col_out_47,
    output [1:0] col_out_48,
    output [1:0] col_out_49,
    output [1:0] col_out_50,
    output [1:0] col_out_51,
    output [1:0] col_out_52,
    output [1:0] col_out_53,
    output [1:0] col_out_54,
    output [1:0] col_out_55,
    output [1:0] col_out_56,
    output [1:0] col_out_57,
    output [1:0] col_out_58,
    output [1:0] col_out_59,
    output [1:0] col_out_60,
    output [1:0] col_out_61,
    output [1:0] col_out_62,
    output [1:0] col_out_63,
    output [1:0] col_out_64,
    output [1:0] col_out_65,
    output [1:0] col_out_66,
    output [1:0] col_out_67,
    output [1:0] col_out_68,
    output [1:0] col_out_69,
    output [1:0] col_out_70,
    output [1:0] col_out_71,
    output [1:0] col_out_72,
    output [1:0] col_out_73,
    output [1:0] col_out_74,
    output [1:0] col_out_75,
    output [1:0] col_out_76,
    output [1:0] col_out_77,
    output [1:0] col_out_78,
    output [1:0] col_out_79,
    output [1:0] col_out_80,
    output [1:0] col_out_81,
    output [1:0] col_out_82,
    output [1:0] col_out_83,
    output [1:0] col_out_84,
    output [1:0] col_out_85,
    output [1:0] col_out_86,
    output [1:0] col_out_87,
    output [1:0] col_out_88,
    output [1:0] col_out_89,
    output [1:0] col_out_90,
    output [1:0] col_out_91,
    output [1:0] col_out_92,
    output [1:0] col_out_93,
    output [1:0] col_out_94,
    output [1:0] col_out_95,
    output [1:0] col_out_96,
    output [1:0] col_out_97,
    output [1:0] col_out_98,
    output [1:0] col_out_99,
    output [1:0] col_out_100,
    output [1:0] col_out_101,
    output [1:0] col_out_102,
    output [1:0] col_out_103,
    output [1:0] col_out_104,
    output [1:0] col_out_105,
    output [1:0] col_out_106,
    output [1:0] col_out_107,
    output [1:0] col_out_108,
    output [1:0] col_out_109,
    output [1:0] col_out_110,
    output [1:0] col_out_111,
    output [1:0] col_out_112,
    output [1:0] col_out_113,
    output [1:0] col_out_114,
    output [1:0] col_out_115,
    output [1:0] col_out_116,
    output [1:0] col_out_117,
    output [1:0] col_out_118,
    output [1:0] col_out_119,
    output [1:0] col_out_120,
    output [1:0] col_out_121,
    output [1:0] col_out_122,
    output [1:0] col_out_123,
    output [1:0] col_out_124,
    output [1:0] col_out_125,
    output [1:0] col_out_126,
    output [1:0] col_out_127,
    output [1:0] col_out_128,
    output [1:0] col_out_129,
    output [1:0] col_out_130,
    output [1:0] col_out_131,
    output [1:0] col_out_132,
    output [1:0] col_out_133,
    output [1:0] col_out_134,
    output [1:0] col_out_135,
    output [1:0] col_out_136,
    output [1:0] col_out_137,
    output [1:0] col_out_138,
    output [1:0] col_out_139,
    output [1:0] col_out_140,
    output [1:0] col_out_141,
    output [1:0] col_out_142,
    output [1:0] col_out_143,
    output [1:0] col_out_144,
    output [1:0] col_out_145,
    output [1:0] col_out_146,
    output [1:0] col_out_147,
    output [1:0] col_out_148,
    output [1:0] col_out_149,
    output [1:0] col_out_150,
    output [1:0] col_out_151,
    output [1:0] col_out_152,
    output [1:0] col_out_153,
    output [1:0] col_out_154,
    output [1:0] col_out_155,
    output [1:0] col_out_156,
    output [1:0] col_out_157,
    output [1:0] col_out_158,
    output [1:0] col_out_159,
    output [1:0] col_out_160,
    output [1:0] col_out_161,
    output [1:0] col_out_162,
    output [1:0] col_out_163,
    output [1:0] col_out_164,
    output [1:0] col_out_165,
    output [1:0] col_out_166,
    output [1:0] col_out_167,
    output [1:0] col_out_168,
    output [1:0] col_out_169,
    output [1:0] col_out_170,
    output [1:0] col_out_171,
    output [1:0] col_out_172,
    output [1:0] col_out_173,
    output [1:0] col_out_174,
    output [1:0] col_out_175,
    output [1:0] col_out_176,
    output [1:0] col_out_177,
    output [1:0] col_out_178,
    output [1:0] col_out_179,
    output [1:0] col_out_180,
    output [1:0] col_out_181,
    output [1:0] col_out_182,
    output [1:0] col_out_183,
    output [1:0] col_out_184,
    output [1:0] col_out_185,
    output [1:0] col_out_186,
    output [1:0] col_out_187,
    output [1:0] col_out_188,
    output [1:0] col_out_189,
    output [1:0] col_out_190,
    output [1:0] col_out_191,
    output [1:0] col_out_192,
    output [1:0] col_out_193,
    output [1:0] col_out_194,
    output [1:0] col_out_195,
    output [1:0] col_out_196,
    output [1:0] col_out_197,
    output [1:0] col_out_198,
    output [1:0] col_out_199,
    output [1:0] col_out_200,
    output [1:0] col_out_201,
    output [1:0] col_out_202,
    output [1:0] col_out_203,
    output [1:0] col_out_204,
    output [1:0] col_out_205,
    output [1:0] col_out_206,
    output [1:0] col_out_207,
    output [1:0] col_out_208,
    output [1:0] col_out_209,
    output [1:0] col_out_210,
    output [1:0] col_out_211,
    output [1:0] col_out_212,
    output [1:0] col_out_213,
    output [1:0] col_out_214,
    output [1:0] col_out_215,
    output [1:0] col_out_216,
    output [1:0] col_out_217,
    output [1:0] col_out_218,
    output [1:0] col_out_219,
    output [1:0] col_out_220,
    output [1:0] col_out_221,
    output [1:0] col_out_222,
    output [1:0] col_out_223,
    output [1:0] col_out_224,
    output [1:0] col_out_225,
    output [1:0] col_out_226,
    output [1:0] col_out_227,
    output [1:0] col_out_228,
    output [1:0] col_out_229,
    output [1:0] col_out_230,
    output [1:0] col_out_231,
    output [1:0] col_out_232,
    output [1:0] col_out_233,
    output [1:0] col_out_234,
    output [1:0] col_out_235,
    output [1:0] col_out_236,
    output [1:0] col_out_237,
    output [1:0] col_out_238,
    output [1:0] col_out_239,
    output [1:0] col_out_240,
    output [1:0] col_out_241,
    output [1:0] col_out_242,
    output [1:0] col_out_243,
    output [1:0] col_out_244,
    output [1:0] col_out_245,
    output [1:0] col_out_246,
    output [1:0] col_out_247,
    output [1:0] col_out_248,
    output [1:0] col_out_249,
    output [1:0] col_out_250,
    output [1:0] col_out_251,
    output [1:0] col_out_252,
    output [1:0] col_out_253,
    output [1:0] col_out_254,
    output [1:0] col_out_255,
    output [1:0] col_out_256,
    output [1:0] col_out_257,
    output [1:0] col_out_258,
    output [1:0] col_out_259,
    output [1:0] col_out_260,
    output [1:0] col_out_261,
    output [1:0] col_out_262,
    output [1:0] col_out_263,
    output [1:0] col_out_264,
    output [1:0] col_out_265,
    output [1:0] col_out_266,
    output [1:0] col_out_267,
    output [1:0] col_out_268,
    output [1:0] col_out_269,
    output [1:0] col_out_270,
    output [1:0] col_out_271,
    output [1:0] col_out_272,
    output [1:0] col_out_273,
    output [1:0] col_out_274,
    output [1:0] col_out_275,
    output [1:0] col_out_276,
    output [1:0] col_out_277,
    output [1:0] col_out_278,
    output [1:0] col_out_279,
    output [1:0] col_out_280,
    output [1:0] col_out_281,
    output [1:0] col_out_282,
    output [1:0] col_out_283,
    output [1:0] col_out_284,
    output [1:0] col_out_285,
    output [1:0] col_out_286,
    output [1:0] col_out_287,
    output [1:0] col_out_288,
    output [1:0] col_out_289,
    output [1:0] col_out_290,
    output [1:0] col_out_291,
    output [1:0] col_out_292,
    output [1:0] col_out_293,
    output [1:0] col_out_294,
    output [1:0] col_out_295,
    output [1:0] col_out_296,
    output [1:0] col_out_297,
    output [1:0] col_out_298,
    output [1:0] col_out_299,
    output [1:0] col_out_300,
    output [1:0] col_out_301,
    output [1:0] col_out_302,
    output [1:0] col_out_303,
    output [1:0] col_out_304,
    output [1:0] col_out_305,
    output [1:0] col_out_306,
    output [1:0] col_out_307,
    output [1:0] col_out_308,
    output [1:0] col_out_309,
    output [1:0] col_out_310,
    output [1:0] col_out_311,
    output [1:0] col_out_312,
    output [1:0] col_out_313,
    output [1:0] col_out_314,
    output [1:0] col_out_315,
    output [1:0] col_out_316,
    output [1:0] col_out_317,
    output [1:0] col_out_318,
    output [1:0] col_out_319,
    output [1:0] col_out_320,
    output [1:0] col_out_321,
    output [1:0] col_out_322,
    output [1:0] col_out_323,
    output [1:0] col_out_324,
    output [1:0] col_out_325,
    output [1:0] col_out_326,
    output [1:0] col_out_327,
    output [1:0] col_out_328,
    output [1:0] col_out_329,
    output [1:0] col_out_330,
    output [1:0] col_out_331,
    output [1:0] col_out_332,
    output [1:0] col_out_333,
    output [1:0] col_out_334,
    output [1:0] col_out_335,
    output [1:0] col_out_336,
    output [1:0] col_out_337,
    output [1:0] col_out_338,
    output [1:0] col_out_339,
    output [1:0] col_out_340,
    output [1:0] col_out_341,
    output [1:0] col_out_342,
    output [1:0] col_out_343,
    output [1:0] col_out_344,
    output [1:0] col_out_345,
    output [1:0] col_out_346,
    output [1:0] col_out_347,
    output [1:0] col_out_348,
    output [1:0] col_out_349,
    output [1:0] col_out_350,
    output [1:0] col_out_351,
    output [1:0] col_out_352,
    output [1:0] col_out_353,
    output [1:0] col_out_354,
    output [1:0] col_out_355,
    output [1:0] col_out_356,
    output [1:0] col_out_357,
    output [1:0] col_out_358,
    output [1:0] col_out_359,
    output [1:0] col_out_360,
    output [1:0] col_out_361,
    output [1:0] col_out_362,
    output [1:0] col_out_363,
    output [1:0] col_out_364,
    output [1:0] col_out_365,
    output [1:0] col_out_366,
    output [1:0] col_out_367,
    output [1:0] col_out_368,
    output [1:0] col_out_369,
    output [1:0] col_out_370,
    output [1:0] col_out_371,
    output [1:0] col_out_372,
    output [1:0] col_out_373,
    output [1:0] col_out_374,
    output [1:0] col_out_375,
    output [1:0] col_out_376,
    output [1:0] col_out_377,
    output [1:0] col_out_378,
    output [1:0] col_out_379,
    output [1:0] col_out_380,
    output [1:0] col_out_381,
    output [1:0] col_out_382,
    output [1:0] col_out_383,
    output [1:0] col_out_384,
    output [1:0] col_out_385,
    output [1:0] col_out_386,
    output [1:0] col_out_387,
    output [1:0] col_out_388,
    output [1:0] col_out_389,
    output [1:0] col_out_390,
    output [1:0] col_out_391,
    output [1:0] col_out_392,
    output [1:0] col_out_393,
    output [1:0] col_out_394,
    output [1:0] col_out_395,
    output [1:0] col_out_396,
    output [1:0] col_out_397,
    output [1:0] col_out_398,
    output [1:0] col_out_399,
    output [1:0] col_out_400,
    output [1:0] col_out_401,
    output [1:0] col_out_402,
    output [1:0] col_out_403,
    output [1:0] col_out_404,
    output [1:0] col_out_405,
    output [1:0] col_out_406,
    output [1:0] col_out_407,
    output [1:0] col_out_408,
    output [1:0] col_out_409,
    output [1:0] col_out_410,
    output [1:0] col_out_411,
    output [1:0] col_out_412,
    output [1:0] col_out_413,
    output [1:0] col_out_414,
    output [1:0] col_out_415,
    output [1:0] col_out_416,
    output [1:0] col_out_417,
    output [1:0] col_out_418,
    output [1:0] col_out_419,
    output [1:0] col_out_420,
    output [1:0] col_out_421,
    output [1:0] col_out_422,
    output [1:0] col_out_423,
    output [1:0] col_out_424,
    output [1:0] col_out_425,
    output [1:0] col_out_426,
    output [1:0] col_out_427,
    output [1:0] col_out_428,
    output [1:0] col_out_429,
    output [1:0] col_out_430,
    output [1:0] col_out_431,
    output [1:0] col_out_432,
    output [1:0] col_out_433,
    output [1:0] col_out_434,
    output [1:0] col_out_435,
    output [1:0] col_out_436,
    output [1:0] col_out_437,
    output [1:0] col_out_438,
    output [1:0] col_out_439,
    output [1:0] col_out_440,
    output [1:0] col_out_441,
    output [1:0] col_out_442,
    output [1:0] col_out_443,
    output [1:0] col_out_444,
    output [1:0] col_out_445,
    output [1:0] col_out_446,
    output [1:0] col_out_447,
    output [1:0] col_out_448,
    output [1:0] col_out_449,
    output [1:0] col_out_450,
    output [1:0] col_out_451,
    output [1:0] col_out_452,
    output [1:0] col_out_453,
    output [1:0] col_out_454,
    output [1:0] col_out_455,
    output [1:0] col_out_456,
    output [1:0] col_out_457,
    output [1:0] col_out_458,
    output [1:0] col_out_459,
    output [1:0] col_out_460,
    output [1:0] col_out_461,
    output [1:0] col_out_462,
    output [1:0] col_out_463,
    output [1:0] col_out_464,
    output [1:0] col_out_465,
    output [1:0] col_out_466,
    output [1:0] col_out_467,
    output [1:0] col_out_468,
    output [1:0] col_out_469,
    output [1:0] col_out_470,
    output [1:0] col_out_471,
    output [1:0] col_out_472,
    output [1:0] col_out_473,
    output [1:0] col_out_474,
    output [1:0] col_out_475,
    output [1:0] col_out_476,
    output [1:0] col_out_477,
    output [1:0] col_out_478,
    output [1:0] col_out_479,
    output [1:0] col_out_480,
    output [1:0] col_out_481,
    output [1:0] col_out_482,
    output [1:0] col_out_483,
    output [1:0] col_out_484,
    output [1:0] col_out_485,
    output [1:0] col_out_486,
    output [1:0] col_out_487,
    output [1:0] col_out_488,
    output [1:0] col_out_489,
    output [1:0] col_out_490,
    output [1:0] col_out_491,
    output [1:0] col_out_492,
    output [1:0] col_out_493,
    output [1:0] col_out_494,
    output [1:0] col_out_495,
    output [1:0] col_out_496,
    output [1:0] col_out_497,
    output [1:0] col_out_498,
    output [1:0] col_out_499,
    output [1:0] col_out_500,
    output [1:0] col_out_501,
    output [1:0] col_out_502,
    output [1:0] col_out_503,
    output [1:0] col_out_504,
    output [1:0] col_out_505,
    output [1:0] col_out_506,
    output [1:0] col_out_507,
    output [1:0] col_out_508,
    output [1:0] col_out_509,
    output [1:0] col_out_510,
    output [1:0] col_out_511,
    output [1:0] col_out_512,
    output [1:0] col_out_513,
    output [1:0] col_out_514,
    output [1:0] col_out_515,
    output [1:0] col_out_516,
    output [1:0] col_out_517,
    output [1:0] col_out_518,
    output [1:0] col_out_519,
    output [1:0] col_out_520,
    output [1:0] col_out_521,
    output [1:0] col_out_522,
    output [1:0] col_out_523,
    output [1:0] col_out_524,
    output [1:0] col_out_525,
    output [1:0] col_out_526,
    output [1:0] col_out_527,
    output [1:0] col_out_528,
    output [1:0] col_out_529,
    output [1:0] col_out_530,
    output [1:0] col_out_531,
    output [1:0] col_out_532,
    output [1:0] col_out_533,
    output [1:0] col_out_534,
    output [1:0] col_out_535,
    output [1:0] col_out_536,
    output [1:0] col_out_537,
    output [1:0] col_out_538,
    output [1:0] col_out_539,
    output [1:0] col_out_540,
    output [1:0] col_out_541,
    output [1:0] col_out_542,
    output [1:0] col_out_543,
    output [1:0] col_out_544,
    output [1:0] col_out_545,
    output [1:0] col_out_546,
    output [1:0] col_out_547,
    output [1:0] col_out_548,
    output [1:0] col_out_549,
    output [1:0] col_out_550,
    output [1:0] col_out_551,
    output [1:0] col_out_552,
    output [1:0] col_out_553,
    output [1:0] col_out_554,
    output [1:0] col_out_555,
    output [1:0] col_out_556,
    output [1:0] col_out_557,
    output [1:0] col_out_558,
    output [1:0] col_out_559,
    output [1:0] col_out_560,
    output [1:0] col_out_561,
    output [1:0] col_out_562,
    output [1:0] col_out_563,
    output [1:0] col_out_564,
    output [1:0] col_out_565,
    output [1:0] col_out_566,
    output [1:0] col_out_567,
    output [1:0] col_out_568,
    output [1:0] col_out_569,
    output [1:0] col_out_570,
    output [1:0] col_out_571,
    output [1:0] col_out_572,
    output [1:0] col_out_573,
    output [1:0] col_out_574,
    output [1:0] col_out_575,
    output [1:0] col_out_576,
    output [1:0] col_out_577,
    output [1:0] col_out_578,
    output [1:0] col_out_579,
    output [1:0] col_out_580,
    output [1:0] col_out_581,
    output [1:0] col_out_582,
    output [1:0] col_out_583,
    output [1:0] col_out_584,
    output [1:0] col_out_585,
    output [1:0] col_out_586,
    output [1:0] col_out_587,
    output [1:0] col_out_588,
    output [1:0] col_out_589,
    output [1:0] col_out_590,
    output [1:0] col_out_591,
    output [1:0] col_out_592,
    output [1:0] col_out_593,
    output [1:0] col_out_594,
    output [1:0] col_out_595,
    output [1:0] col_out_596,
    output [1:0] col_out_597,
    output [1:0] col_out_598,
    output [1:0] col_out_599,
    output [1:0] col_out_600,
    output [1:0] col_out_601,
    output [1:0] col_out_602,
    output [1:0] col_out_603,
    output [1:0] col_out_604,
    output [1:0] col_out_605,
    output [1:0] col_out_606,
    output [1:0] col_out_607,
    output [1:0] col_out_608,
    output [1:0] col_out_609,
    output [1:0] col_out_610,
    output [1:0] col_out_611,
    output [1:0] col_out_612,
    output [1:0] col_out_613,
    output [1:0] col_out_614,
    output [1:0] col_out_615,
    output [1:0] col_out_616,
    output [1:0] col_out_617,
    output [1:0] col_out_618,
    output [1:0] col_out_619,
    output [1:0] col_out_620,
    output [1:0] col_out_621,
    output [1:0] col_out_622,
    output [1:0] col_out_623,
    output [1:0] col_out_624,
    output [1:0] col_out_625,
    output [1:0] col_out_626,
    output [1:0] col_out_627,
    output [1:0] col_out_628,
    output [1:0] col_out_629,
    output [1:0] col_out_630,
    output [1:0] col_out_631,
    output [1:0] col_out_632,
    output [1:0] col_out_633,
    output [1:0] col_out_634,
    output [1:0] col_out_635,
    output [1:0] col_out_636,
    output [1:0] col_out_637,
    output [1:0] col_out_638,
    output [1:0] col_out_639,
    output [1:0] col_out_640,
    output [1:0] col_out_641,
    output [1:0] col_out_642,
    output [1:0] col_out_643,
    output [1:0] col_out_644,
    output [1:0] col_out_645,
    output [1:0] col_out_646,
    output [1:0] col_out_647,
    output [1:0] col_out_648,
    output [1:0] col_out_649,
    output [1:0] col_out_650,
    output [1:0] col_out_651,
    output [1:0] col_out_652,
    output [1:0] col_out_653,
    output [1:0] col_out_654,
    output [1:0] col_out_655,
    output [1:0] col_out_656,
    output [1:0] col_out_657,
    output [1:0] col_out_658,
    output [1:0] col_out_659,
    output [1:0] col_out_660,
    output [1:0] col_out_661,
    output [1:0] col_out_662,
    output [1:0] col_out_663,
    output [1:0] col_out_664,
    output [1:0] col_out_665,
    output [1:0] col_out_666,
    output [1:0] col_out_667,
    output [1:0] col_out_668,
    output [1:0] col_out_669,
    output [1:0] col_out_670,
    output [1:0] col_out_671,
    output [1:0] col_out_672,
    output [1:0] col_out_673,
    output [1:0] col_out_674,
    output [1:0] col_out_675,
    output [1:0] col_out_676,
    output [1:0] col_out_677,
    output [1:0] col_out_678,
    output [1:0] col_out_679,
    output [1:0] col_out_680,
    output [1:0] col_out_681,
    output [1:0] col_out_682,
    output [1:0] col_out_683,
    output [1:0] col_out_684,
    output [1:0] col_out_685,
    output [1:0] col_out_686,
    output [1:0] col_out_687,
    output [1:0] col_out_688,
    output [1:0] col_out_689,
    output [1:0] col_out_690,
    output [1:0] col_out_691,
    output [1:0] col_out_692,
    output [1:0] col_out_693,
    output [1:0] col_out_694,
    output [1:0] col_out_695,
    output [1:0] col_out_696,
    output [1:0] col_out_697,
    output [1:0] col_out_698,
    output [1:0] col_out_699,
    output [1:0] col_out_700,
    output [1:0] col_out_701,
    output [1:0] col_out_702,
    output [1:0] col_out_703,
    output [1:0] col_out_704,
    output [1:0] col_out_705,
    output [1:0] col_out_706,
    output [1:0] col_out_707,
    output [1:0] col_out_708,
    output [1:0] col_out_709,
    output [1:0] col_out_710,
    output [1:0] col_out_711,
    output [1:0] col_out_712,
    output [1:0] col_out_713,
    output [1:0] col_out_714,
    output [1:0] col_out_715,
    output [1:0] col_out_716,
    output [1:0] col_out_717,
    output [1:0] col_out_718,
    output [1:0] col_out_719,
    output [1:0] col_out_720,
    output [1:0] col_out_721,
    output [1:0] col_out_722,
    output [1:0] col_out_723,
    output [1:0] col_out_724,
    output [1:0] col_out_725,
    output [1:0] col_out_726,
    output [1:0] col_out_727,
    output [1:0] col_out_728,
    output [1:0] col_out_729,
    output [1:0] col_out_730,
    output [1:0] col_out_731,
    output [1:0] col_out_732,
    output [1:0] col_out_733,
    output [1:0] col_out_734,
    output [1:0] col_out_735,
    output [1:0] col_out_736,
    output [1:0] col_out_737,
    output [1:0] col_out_738,
    output [1:0] col_out_739,
    output [1:0] col_out_740,
    output [1:0] col_out_741,
    output [1:0] col_out_742,
    output [1:0] col_out_743,
    output [1:0] col_out_744,
    output [1:0] col_out_745,
    output [1:0] col_out_746,
    output [1:0] col_out_747,
    output [1:0] col_out_748,
    output [1:0] col_out_749,
    output [1:0] col_out_750,
    output [1:0] col_out_751,
    output [1:0] col_out_752,
    output [1:0] col_out_753,
    output [1:0] col_out_754,
    output [1:0] col_out_755,
    output [1:0] col_out_756,
    output [1:0] col_out_757,
    output [1:0] col_out_758,
    output [1:0] col_out_759,
    output [1:0] col_out_760,
    output [1:0] col_out_761,
    output [1:0] col_out_762,
    output [1:0] col_out_763,
    output [1:0] col_out_764,
    output [1:0] col_out_765,
    output [1:0] col_out_766,
    output [1:0] col_out_767,
    output [1:0] col_out_768,
    output [1:0] col_out_769,
    output [1:0] col_out_770,
    output [1:0] col_out_771,
    output [1:0] col_out_772,
    output [1:0] col_out_773,
    output [1:0] col_out_774,
    output [1:0] col_out_775,
    output [1:0] col_out_776,
    output [1:0] col_out_777,
    output [1:0] col_out_778,
    output [1:0] col_out_779,
    output [1:0] col_out_780,
    output [1:0] col_out_781,
    output [1:0] col_out_782,
    output [1:0] col_out_783,
    output [1:0] col_out_784,
    output [1:0] col_out_785,
    output [1:0] col_out_786,
    output [1:0] col_out_787,
    output [1:0] col_out_788,
    output [1:0] col_out_789,
    output [1:0] col_out_790,
    output [1:0] col_out_791,
    output [1:0] col_out_792,
    output [1:0] col_out_793,
    output [1:0] col_out_794,
    output [1:0] col_out_795,
    output [1:0] col_out_796,
    output [1:0] col_out_797,
    output [1:0] col_out_798,
    output [1:0] col_out_799,
    output [1:0] col_out_800,
    output [1:0] col_out_801,
    output [1:0] col_out_802,
    output [1:0] col_out_803,
    output [1:0] col_out_804,
    output [1:0] col_out_805,
    output [1:0] col_out_806,
    output [1:0] col_out_807,
    output [1:0] col_out_808,
    output [1:0] col_out_809,
    output [1:0] col_out_810,
    output [1:0] col_out_811,
    output [1:0] col_out_812,
    output [1:0] col_out_813,
    output [1:0] col_out_814,
    output [1:0] col_out_815,
    output [1:0] col_out_816,
    output [1:0] col_out_817,
    output [1:0] col_out_818,
    output [1:0] col_out_819,
    output [1:0] col_out_820,
    output [1:0] col_out_821,
    output [1:0] col_out_822,
    output [1:0] col_out_823,
    output [1:0] col_out_824,
    output [1:0] col_out_825,
    output [1:0] col_out_826,
    output [1:0] col_out_827,
    output [1:0] col_out_828,
    output [1:0] col_out_829,
    output [1:0] col_out_830,
    output [1:0] col_out_831,
    output [1:0] col_out_832,
    output [1:0] col_out_833,
    output [1:0] col_out_834,
    output [1:0] col_out_835,
    output [1:0] col_out_836,
    output [1:0] col_out_837,
    output [1:0] col_out_838,
    output [1:0] col_out_839,
    output [1:0] col_out_840,
    output [1:0] col_out_841,
    output [1:0] col_out_842,
    output [1:0] col_out_843,
    output [1:0] col_out_844,
    output [1:0] col_out_845,
    output [1:0] col_out_846,
    output [1:0] col_out_847,
    output [1:0] col_out_848,
    output [1:0] col_out_849,
    output [1:0] col_out_850,
    output [1:0] col_out_851,
    output [1:0] col_out_852,
    output [1:0] col_out_853,
    output [1:0] col_out_854,
    output [1:0] col_out_855,
    output [1:0] col_out_856,
    output [1:0] col_out_857,
    output [1:0] col_out_858,
    output [1:0] col_out_859,
    output [1:0] col_out_860,
    output [1:0] col_out_861,
    output [1:0] col_out_862,
    output [1:0] col_out_863,
    output [1:0] col_out_864,
    output [1:0] col_out_865,
    output [1:0] col_out_866,
    output [1:0] col_out_867,
    output [1:0] col_out_868,
    output [1:0] col_out_869,
    output [1:0] col_out_870,
    output [1:0] col_out_871,
    output [1:0] col_out_872,
    output [1:0] col_out_873,
    output [1:0] col_out_874,
    output [1:0] col_out_875,
    output [1:0] col_out_876,
    output [1:0] col_out_877,
    output [1:0] col_out_878,
    output [1:0] col_out_879,
    output [1:0] col_out_880,
    output [1:0] col_out_881,
    output [1:0] col_out_882,
    output [1:0] col_out_883,
    output [1:0] col_out_884,
    output [1:0] col_out_885,
    output [1:0] col_out_886,
    output [1:0] col_out_887,
    output [1:0] col_out_888,
    output [1:0] col_out_889,
    output [1:0] col_out_890,
    output [1:0] col_out_891,
    output [1:0] col_out_892,
    output [1:0] col_out_893,
    output [1:0] col_out_894,
    output [1:0] col_out_895,
    output [1:0] col_out_896,
    output [1:0] col_out_897,
    output [1:0] col_out_898,
    output [1:0] col_out_899,
    output [1:0] col_out_900,
    output [1:0] col_out_901,
    output [1:0] col_out_902,
    output [1:0] col_out_903,
    output [1:0] col_out_904,
    output [1:0] col_out_905,
    output [1:0] col_out_906,
    output [1:0] col_out_907,
    output [1:0] col_out_908,
    output [1:0] col_out_909,
    output [1:0] col_out_910,
    output [1:0] col_out_911,
    output [1:0] col_out_912,
    output [1:0] col_out_913,
    output [1:0] col_out_914,
    output [1:0] col_out_915,
    output [1:0] col_out_916,
    output [1:0] col_out_917,
    output [1:0] col_out_918,
    output [1:0] col_out_919,
    output [1:0] col_out_920,
    output [1:0] col_out_921,
    output [1:0] col_out_922,
    output [1:0] col_out_923,
    output [1:0] col_out_924,
    output [1:0] col_out_925,
    output [1:0] col_out_926,
    output [1:0] col_out_927,
    output [1:0] col_out_928,
    output [1:0] col_out_929,
    output [1:0] col_out_930,
    output [1:0] col_out_931,
    output [1:0] col_out_932,
    output [1:0] col_out_933,
    output [1:0] col_out_934,
    output [1:0] col_out_935,
    output [1:0] col_out_936,
    output [1:0] col_out_937,
    output [1:0] col_out_938,
    output [1:0] col_out_939,
    output [1:0] col_out_940,
    output [1:0] col_out_941,
    output [1:0] col_out_942,
    output [1:0] col_out_943,
    output [1:0] col_out_944,
    output [1:0] col_out_945,
    output [1:0] col_out_946,
    output [1:0] col_out_947,
    output [1:0] col_out_948,
    output [1:0] col_out_949,
    output [1:0] col_out_950,
    output [1:0] col_out_951,
    output [1:0] col_out_952,
    output [1:0] col_out_953,
    output [1:0] col_out_954,
    output [1:0] col_out_955,
    output [1:0] col_out_956,
    output [1:0] col_out_957,
    output [1:0] col_out_958,
    output [1:0] col_out_959,
    output [1:0] col_out_960,
    output [1:0] col_out_961,
    output [1:0] col_out_962,
    output [1:0] col_out_963,
    output [1:0] col_out_964,
    output [1:0] col_out_965,
    output [1:0] col_out_966,
    output [1:0] col_out_967,
    output [1:0] col_out_968,
    output [1:0] col_out_969,
    output [1:0] col_out_970,
    output [1:0] col_out_971,
    output [1:0] col_out_972,
    output [1:0] col_out_973,
    output [1:0] col_out_974,
    output [1:0] col_out_975,
    output [1:0] col_out_976,
    output [1:0] col_out_977,
    output [1:0] col_out_978,
    output [1:0] col_out_979,
    output [1:0] col_out_980,
    output [1:0] col_out_981,
    output [1:0] col_out_982,
    output [1:0] col_out_983,
    output [1:0] col_out_984,
    output [1:0] col_out_985,
    output [1:0] col_out_986,
    output [1:0] col_out_987,
    output [1:0] col_out_988,
    output [1:0] col_out_989,
    output [1:0] col_out_990,
    output [1:0] col_out_991,
    output [1:0] col_out_992,
    output [1:0] col_out_993,
    output [1:0] col_out_994,
    output [1:0] col_out_995,
    output [1:0] col_out_996,
    output [1:0] col_out_997,
    output [1:0] col_out_998,
    output [1:0] col_out_999,
    output [1:0] col_out_1000,
    output [1:0] col_out_1001,
    output [1:0] col_out_1002,
    output [1:0] col_out_1003,
    output [1:0] col_out_1004,
    output [1:0] col_out_1005,
    output [1:0] col_out_1006,
    output [1:0] col_out_1007,
    output [1:0] col_out_1008,
    output [1:0] col_out_1009,
    output [1:0] col_out_1010,
    output [1:0] col_out_1011,
    output [1:0] col_out_1012,
    output [1:0] col_out_1013,
    output [1:0] col_out_1014,
    output [1:0] col_out_1015,
    output [1:0] col_out_1016,
    output [1:0] col_out_1017,
    output [1:0] col_out_1018,
    output [1:0] col_out_1019,
    output [1:0] col_out_1020,
    output [1:0] col_out_1021,
    output [1:0] col_out_1022,
    output [1:0] col_out_1023,
    output [1:0] col_out_1024
);



//--compressor_array input and output----------------------

wire [2:0] u_ca_in_0;
wire [2:0] u_ca_in_1;
wire [2:0] u_ca_in_2;
wire [2:0] u_ca_in_3;
wire [2:0] u_ca_in_4;
wire [2:0] u_ca_in_5;
wire [2:0] u_ca_in_6;
wire [2:0] u_ca_in_7;
wire [2:0] u_ca_in_8;
wire [2:0] u_ca_in_9;
wire [2:0] u_ca_in_10;
wire [2:0] u_ca_in_11;
wire [2:0] u_ca_in_12;
wire [2:0] u_ca_in_13;
wire [2:0] u_ca_in_14;
wire [2:0] u_ca_in_15;
wire [2:0] u_ca_in_16;
wire [2:0] u_ca_in_17;
wire [2:0] u_ca_in_18;
wire [2:0] u_ca_in_19;
wire [2:0] u_ca_in_20;
wire [2:0] u_ca_in_21;
wire [2:0] u_ca_in_22;
wire [2:0] u_ca_in_23;
wire [2:0] u_ca_in_24;
wire [2:0] u_ca_in_25;
wire [2:0] u_ca_in_26;
wire [2:0] u_ca_in_27;
wire [2:0] u_ca_in_28;
wire [2:0] u_ca_in_29;
wire [2:0] u_ca_in_30;
wire [2:0] u_ca_in_31;
wire [2:0] u_ca_in_32;
wire [2:0] u_ca_in_33;
wire [2:0] u_ca_in_34;
wire [2:0] u_ca_in_35;
wire [2:0] u_ca_in_36;
wire [2:0] u_ca_in_37;
wire [2:0] u_ca_in_38;
wire [2:0] u_ca_in_39;
wire [2:0] u_ca_in_40;
wire [2:0] u_ca_in_41;
wire [2:0] u_ca_in_42;
wire [2:0] u_ca_in_43;
wire [2:0] u_ca_in_44;
wire [2:0] u_ca_in_45;
wire [2:0] u_ca_in_46;
wire [2:0] u_ca_in_47;
wire [2:0] u_ca_in_48;
wire [2:0] u_ca_in_49;
wire [2:0] u_ca_in_50;
wire [2:0] u_ca_in_51;
wire [2:0] u_ca_in_52;
wire [2:0] u_ca_in_53;
wire [2:0] u_ca_in_54;
wire [2:0] u_ca_in_55;
wire [2:0] u_ca_in_56;
wire [2:0] u_ca_in_57;
wire [2:0] u_ca_in_58;
wire [2:0] u_ca_in_59;
wire [2:0] u_ca_in_60;
wire [2:0] u_ca_in_61;
wire [2:0] u_ca_in_62;
wire [2:0] u_ca_in_63;
wire [2:0] u_ca_in_64;
wire [2:0] u_ca_in_65;
wire [2:0] u_ca_in_66;
wire [2:0] u_ca_in_67;
wire [2:0] u_ca_in_68;
wire [2:0] u_ca_in_69;
wire [2:0] u_ca_in_70;
wire [2:0] u_ca_in_71;
wire [2:0] u_ca_in_72;
wire [2:0] u_ca_in_73;
wire [2:0] u_ca_in_74;
wire [2:0] u_ca_in_75;
wire [2:0] u_ca_in_76;
wire [2:0] u_ca_in_77;
wire [2:0] u_ca_in_78;
wire [2:0] u_ca_in_79;
wire [2:0] u_ca_in_80;
wire [2:0] u_ca_in_81;
wire [2:0] u_ca_in_82;
wire [2:0] u_ca_in_83;
wire [2:0] u_ca_in_84;
wire [2:0] u_ca_in_85;
wire [2:0] u_ca_in_86;
wire [2:0] u_ca_in_87;
wire [2:0] u_ca_in_88;
wire [2:0] u_ca_in_89;
wire [2:0] u_ca_in_90;
wire [2:0] u_ca_in_91;
wire [2:0] u_ca_in_92;
wire [2:0] u_ca_in_93;
wire [2:0] u_ca_in_94;
wire [2:0] u_ca_in_95;
wire [2:0] u_ca_in_96;
wire [2:0] u_ca_in_97;
wire [2:0] u_ca_in_98;
wire [2:0] u_ca_in_99;
wire [2:0] u_ca_in_100;
wire [2:0] u_ca_in_101;
wire [2:0] u_ca_in_102;
wire [2:0] u_ca_in_103;
wire [2:0] u_ca_in_104;
wire [2:0] u_ca_in_105;
wire [2:0] u_ca_in_106;
wire [2:0] u_ca_in_107;
wire [2:0] u_ca_in_108;
wire [2:0] u_ca_in_109;
wire [2:0] u_ca_in_110;
wire [2:0] u_ca_in_111;
wire [2:0] u_ca_in_112;
wire [2:0] u_ca_in_113;
wire [2:0] u_ca_in_114;
wire [2:0] u_ca_in_115;
wire [2:0] u_ca_in_116;
wire [2:0] u_ca_in_117;
wire [2:0] u_ca_in_118;
wire [2:0] u_ca_in_119;
wire [2:0] u_ca_in_120;
wire [2:0] u_ca_in_121;
wire [2:0] u_ca_in_122;
wire [2:0] u_ca_in_123;
wire [2:0] u_ca_in_124;
wire [2:0] u_ca_in_125;
wire [2:0] u_ca_in_126;
wire [2:0] u_ca_in_127;
wire [2:0] u_ca_in_128;
wire [2:0] u_ca_in_129;
wire [2:0] u_ca_in_130;
wire [2:0] u_ca_in_131;
wire [2:0] u_ca_in_132;
wire [2:0] u_ca_in_133;
wire [2:0] u_ca_in_134;
wire [2:0] u_ca_in_135;
wire [2:0] u_ca_in_136;
wire [2:0] u_ca_in_137;
wire [2:0] u_ca_in_138;
wire [2:0] u_ca_in_139;
wire [2:0] u_ca_in_140;
wire [2:0] u_ca_in_141;
wire [2:0] u_ca_in_142;
wire [2:0] u_ca_in_143;
wire [2:0] u_ca_in_144;
wire [2:0] u_ca_in_145;
wire [2:0] u_ca_in_146;
wire [2:0] u_ca_in_147;
wire [2:0] u_ca_in_148;
wire [2:0] u_ca_in_149;
wire [2:0] u_ca_in_150;
wire [2:0] u_ca_in_151;
wire [2:0] u_ca_in_152;
wire [2:0] u_ca_in_153;
wire [2:0] u_ca_in_154;
wire [2:0] u_ca_in_155;
wire [2:0] u_ca_in_156;
wire [2:0] u_ca_in_157;
wire [2:0] u_ca_in_158;
wire [2:0] u_ca_in_159;
wire [2:0] u_ca_in_160;
wire [2:0] u_ca_in_161;
wire [2:0] u_ca_in_162;
wire [2:0] u_ca_in_163;
wire [2:0] u_ca_in_164;
wire [2:0] u_ca_in_165;
wire [2:0] u_ca_in_166;
wire [2:0] u_ca_in_167;
wire [2:0] u_ca_in_168;
wire [2:0] u_ca_in_169;
wire [2:0] u_ca_in_170;
wire [2:0] u_ca_in_171;
wire [2:0] u_ca_in_172;
wire [2:0] u_ca_in_173;
wire [2:0] u_ca_in_174;
wire [2:0] u_ca_in_175;
wire [2:0] u_ca_in_176;
wire [2:0] u_ca_in_177;
wire [2:0] u_ca_in_178;
wire [2:0] u_ca_in_179;
wire [2:0] u_ca_in_180;
wire [2:0] u_ca_in_181;
wire [2:0] u_ca_in_182;
wire [2:0] u_ca_in_183;
wire [2:0] u_ca_in_184;
wire [2:0] u_ca_in_185;
wire [2:0] u_ca_in_186;
wire [2:0] u_ca_in_187;
wire [2:0] u_ca_in_188;
wire [2:0] u_ca_in_189;
wire [2:0] u_ca_in_190;
wire [2:0] u_ca_in_191;
wire [2:0] u_ca_in_192;
wire [2:0] u_ca_in_193;
wire [2:0] u_ca_in_194;
wire [2:0] u_ca_in_195;
wire [2:0] u_ca_in_196;
wire [2:0] u_ca_in_197;
wire [2:0] u_ca_in_198;
wire [2:0] u_ca_in_199;
wire [2:0] u_ca_in_200;
wire [2:0] u_ca_in_201;
wire [2:0] u_ca_in_202;
wire [2:0] u_ca_in_203;
wire [2:0] u_ca_in_204;
wire [2:0] u_ca_in_205;
wire [2:0] u_ca_in_206;
wire [2:0] u_ca_in_207;
wire [2:0] u_ca_in_208;
wire [2:0] u_ca_in_209;
wire [2:0] u_ca_in_210;
wire [2:0] u_ca_in_211;
wire [2:0] u_ca_in_212;
wire [2:0] u_ca_in_213;
wire [2:0] u_ca_in_214;
wire [2:0] u_ca_in_215;
wire [2:0] u_ca_in_216;
wire [2:0] u_ca_in_217;
wire [2:0] u_ca_in_218;
wire [2:0] u_ca_in_219;
wire [2:0] u_ca_in_220;
wire [2:0] u_ca_in_221;
wire [2:0] u_ca_in_222;
wire [2:0] u_ca_in_223;
wire [2:0] u_ca_in_224;
wire [2:0] u_ca_in_225;
wire [2:0] u_ca_in_226;
wire [2:0] u_ca_in_227;
wire [2:0] u_ca_in_228;
wire [2:0] u_ca_in_229;
wire [2:0] u_ca_in_230;
wire [2:0] u_ca_in_231;
wire [2:0] u_ca_in_232;
wire [2:0] u_ca_in_233;
wire [2:0] u_ca_in_234;
wire [2:0] u_ca_in_235;
wire [2:0] u_ca_in_236;
wire [2:0] u_ca_in_237;
wire [2:0] u_ca_in_238;
wire [2:0] u_ca_in_239;
wire [2:0] u_ca_in_240;
wire [2:0] u_ca_in_241;
wire [2:0] u_ca_in_242;
wire [2:0] u_ca_in_243;
wire [2:0] u_ca_in_244;
wire [2:0] u_ca_in_245;
wire [2:0] u_ca_in_246;
wire [2:0] u_ca_in_247;
wire [2:0] u_ca_in_248;
wire [2:0] u_ca_in_249;
wire [2:0] u_ca_in_250;
wire [2:0] u_ca_in_251;
wire [2:0] u_ca_in_252;
wire [2:0] u_ca_in_253;
wire [2:0] u_ca_in_254;
wire [2:0] u_ca_in_255;
wire [2:0] u_ca_in_256;
wire [2:0] u_ca_in_257;
wire [2:0] u_ca_in_258;
wire [2:0] u_ca_in_259;
wire [2:0] u_ca_in_260;
wire [2:0] u_ca_in_261;
wire [2:0] u_ca_in_262;
wire [2:0] u_ca_in_263;
wire [2:0] u_ca_in_264;
wire [2:0] u_ca_in_265;
wire [2:0] u_ca_in_266;
wire [2:0] u_ca_in_267;
wire [2:0] u_ca_in_268;
wire [2:0] u_ca_in_269;
wire [2:0] u_ca_in_270;
wire [2:0] u_ca_in_271;
wire [2:0] u_ca_in_272;
wire [2:0] u_ca_in_273;
wire [2:0] u_ca_in_274;
wire [2:0] u_ca_in_275;
wire [2:0] u_ca_in_276;
wire [2:0] u_ca_in_277;
wire [2:0] u_ca_in_278;
wire [2:0] u_ca_in_279;
wire [2:0] u_ca_in_280;
wire [2:0] u_ca_in_281;
wire [2:0] u_ca_in_282;
wire [2:0] u_ca_in_283;
wire [2:0] u_ca_in_284;
wire [2:0] u_ca_in_285;
wire [2:0] u_ca_in_286;
wire [2:0] u_ca_in_287;
wire [2:0] u_ca_in_288;
wire [2:0] u_ca_in_289;
wire [2:0] u_ca_in_290;
wire [2:0] u_ca_in_291;
wire [2:0] u_ca_in_292;
wire [2:0] u_ca_in_293;
wire [2:0] u_ca_in_294;
wire [2:0] u_ca_in_295;
wire [2:0] u_ca_in_296;
wire [2:0] u_ca_in_297;
wire [2:0] u_ca_in_298;
wire [2:0] u_ca_in_299;
wire [2:0] u_ca_in_300;
wire [2:0] u_ca_in_301;
wire [2:0] u_ca_in_302;
wire [2:0] u_ca_in_303;
wire [2:0] u_ca_in_304;
wire [2:0] u_ca_in_305;
wire [2:0] u_ca_in_306;
wire [2:0] u_ca_in_307;
wire [2:0] u_ca_in_308;
wire [2:0] u_ca_in_309;
wire [2:0] u_ca_in_310;
wire [2:0] u_ca_in_311;
wire [2:0] u_ca_in_312;
wire [2:0] u_ca_in_313;
wire [2:0] u_ca_in_314;
wire [2:0] u_ca_in_315;
wire [2:0] u_ca_in_316;
wire [2:0] u_ca_in_317;
wire [2:0] u_ca_in_318;
wire [2:0] u_ca_in_319;
wire [2:0] u_ca_in_320;
wire [2:0] u_ca_in_321;
wire [2:0] u_ca_in_322;
wire [2:0] u_ca_in_323;
wire [2:0] u_ca_in_324;
wire [2:0] u_ca_in_325;
wire [2:0] u_ca_in_326;
wire [2:0] u_ca_in_327;
wire [2:0] u_ca_in_328;
wire [2:0] u_ca_in_329;
wire [2:0] u_ca_in_330;
wire [2:0] u_ca_in_331;
wire [2:0] u_ca_in_332;
wire [2:0] u_ca_in_333;
wire [2:0] u_ca_in_334;
wire [2:0] u_ca_in_335;
wire [2:0] u_ca_in_336;
wire [2:0] u_ca_in_337;
wire [2:0] u_ca_in_338;
wire [2:0] u_ca_in_339;
wire [2:0] u_ca_in_340;
wire [2:0] u_ca_in_341;
wire [2:0] u_ca_in_342;
wire [2:0] u_ca_in_343;
wire [2:0] u_ca_in_344;
wire [2:0] u_ca_in_345;
wire [2:0] u_ca_in_346;
wire [2:0] u_ca_in_347;
wire [2:0] u_ca_in_348;
wire [2:0] u_ca_in_349;
wire [2:0] u_ca_in_350;
wire [2:0] u_ca_in_351;
wire [2:0] u_ca_in_352;
wire [2:0] u_ca_in_353;
wire [2:0] u_ca_in_354;
wire [2:0] u_ca_in_355;
wire [2:0] u_ca_in_356;
wire [2:0] u_ca_in_357;
wire [2:0] u_ca_in_358;
wire [2:0] u_ca_in_359;
wire [2:0] u_ca_in_360;
wire [2:0] u_ca_in_361;
wire [2:0] u_ca_in_362;
wire [2:0] u_ca_in_363;
wire [2:0] u_ca_in_364;
wire [2:0] u_ca_in_365;
wire [2:0] u_ca_in_366;
wire [2:0] u_ca_in_367;
wire [2:0] u_ca_in_368;
wire [2:0] u_ca_in_369;
wire [2:0] u_ca_in_370;
wire [2:0] u_ca_in_371;
wire [2:0] u_ca_in_372;
wire [2:0] u_ca_in_373;
wire [2:0] u_ca_in_374;
wire [2:0] u_ca_in_375;
wire [2:0] u_ca_in_376;
wire [2:0] u_ca_in_377;
wire [2:0] u_ca_in_378;
wire [2:0] u_ca_in_379;
wire [2:0] u_ca_in_380;
wire [2:0] u_ca_in_381;
wire [2:0] u_ca_in_382;
wire [2:0] u_ca_in_383;
wire [2:0] u_ca_in_384;
wire [2:0] u_ca_in_385;
wire [2:0] u_ca_in_386;
wire [2:0] u_ca_in_387;
wire [2:0] u_ca_in_388;
wire [2:0] u_ca_in_389;
wire [2:0] u_ca_in_390;
wire [2:0] u_ca_in_391;
wire [2:0] u_ca_in_392;
wire [2:0] u_ca_in_393;
wire [2:0] u_ca_in_394;
wire [2:0] u_ca_in_395;
wire [2:0] u_ca_in_396;
wire [2:0] u_ca_in_397;
wire [2:0] u_ca_in_398;
wire [2:0] u_ca_in_399;
wire [2:0] u_ca_in_400;
wire [2:0] u_ca_in_401;
wire [2:0] u_ca_in_402;
wire [2:0] u_ca_in_403;
wire [2:0] u_ca_in_404;
wire [2:0] u_ca_in_405;
wire [2:0] u_ca_in_406;
wire [2:0] u_ca_in_407;
wire [2:0] u_ca_in_408;
wire [2:0] u_ca_in_409;
wire [2:0] u_ca_in_410;
wire [2:0] u_ca_in_411;
wire [2:0] u_ca_in_412;
wire [2:0] u_ca_in_413;
wire [2:0] u_ca_in_414;
wire [2:0] u_ca_in_415;
wire [2:0] u_ca_in_416;
wire [2:0] u_ca_in_417;
wire [2:0] u_ca_in_418;
wire [2:0] u_ca_in_419;
wire [2:0] u_ca_in_420;
wire [2:0] u_ca_in_421;
wire [2:0] u_ca_in_422;
wire [2:0] u_ca_in_423;
wire [2:0] u_ca_in_424;
wire [2:0] u_ca_in_425;
wire [2:0] u_ca_in_426;
wire [2:0] u_ca_in_427;
wire [2:0] u_ca_in_428;
wire [2:0] u_ca_in_429;
wire [2:0] u_ca_in_430;
wire [2:0] u_ca_in_431;
wire [2:0] u_ca_in_432;
wire [2:0] u_ca_in_433;
wire [2:0] u_ca_in_434;
wire [2:0] u_ca_in_435;
wire [2:0] u_ca_in_436;
wire [2:0] u_ca_in_437;
wire [2:0] u_ca_in_438;
wire [2:0] u_ca_in_439;
wire [2:0] u_ca_in_440;
wire [2:0] u_ca_in_441;
wire [2:0] u_ca_in_442;
wire [2:0] u_ca_in_443;
wire [2:0] u_ca_in_444;
wire [2:0] u_ca_in_445;
wire [2:0] u_ca_in_446;
wire [2:0] u_ca_in_447;
wire [2:0] u_ca_in_448;
wire [2:0] u_ca_in_449;
wire [2:0] u_ca_in_450;
wire [2:0] u_ca_in_451;
wire [2:0] u_ca_in_452;
wire [2:0] u_ca_in_453;
wire [2:0] u_ca_in_454;
wire [2:0] u_ca_in_455;
wire [2:0] u_ca_in_456;
wire [2:0] u_ca_in_457;
wire [2:0] u_ca_in_458;
wire [2:0] u_ca_in_459;
wire [2:0] u_ca_in_460;
wire [2:0] u_ca_in_461;
wire [2:0] u_ca_in_462;
wire [2:0] u_ca_in_463;
wire [2:0] u_ca_in_464;
wire [2:0] u_ca_in_465;
wire [2:0] u_ca_in_466;
wire [2:0] u_ca_in_467;
wire [2:0] u_ca_in_468;
wire [2:0] u_ca_in_469;
wire [2:0] u_ca_in_470;
wire [2:0] u_ca_in_471;
wire [2:0] u_ca_in_472;
wire [2:0] u_ca_in_473;
wire [2:0] u_ca_in_474;
wire [2:0] u_ca_in_475;
wire [2:0] u_ca_in_476;
wire [2:0] u_ca_in_477;
wire [2:0] u_ca_in_478;
wire [2:0] u_ca_in_479;
wire [2:0] u_ca_in_480;
wire [2:0] u_ca_in_481;
wire [2:0] u_ca_in_482;
wire [2:0] u_ca_in_483;
wire [2:0] u_ca_in_484;
wire [2:0] u_ca_in_485;
wire [2:0] u_ca_in_486;
wire [2:0] u_ca_in_487;
wire [2:0] u_ca_in_488;
wire [2:0] u_ca_in_489;
wire [2:0] u_ca_in_490;
wire [2:0] u_ca_in_491;
wire [2:0] u_ca_in_492;
wire [2:0] u_ca_in_493;
wire [2:0] u_ca_in_494;
wire [2:0] u_ca_in_495;
wire [2:0] u_ca_in_496;
wire [2:0] u_ca_in_497;
wire [2:0] u_ca_in_498;
wire [2:0] u_ca_in_499;
wire [2:0] u_ca_in_500;
wire [2:0] u_ca_in_501;
wire [2:0] u_ca_in_502;
wire [2:0] u_ca_in_503;
wire [2:0] u_ca_in_504;
wire [2:0] u_ca_in_505;
wire [2:0] u_ca_in_506;
wire [2:0] u_ca_in_507;
wire [2:0] u_ca_in_508;
wire [2:0] u_ca_in_509;
wire [2:0] u_ca_in_510;
wire [2:0] u_ca_in_511;
wire [2:0] u_ca_in_512;
wire [2:0] u_ca_in_513;
wire [2:0] u_ca_in_514;
wire [2:0] u_ca_in_515;
wire [2:0] u_ca_in_516;
wire [2:0] u_ca_in_517;
wire [2:0] u_ca_in_518;
wire [2:0] u_ca_in_519;
wire [2:0] u_ca_in_520;
wire [2:0] u_ca_in_521;
wire [2:0] u_ca_in_522;
wire [2:0] u_ca_in_523;
wire [2:0] u_ca_in_524;
wire [2:0] u_ca_in_525;
wire [2:0] u_ca_in_526;
wire [2:0] u_ca_in_527;
wire [2:0] u_ca_in_528;
wire [2:0] u_ca_in_529;
wire [2:0] u_ca_in_530;
wire [2:0] u_ca_in_531;
wire [2:0] u_ca_in_532;
wire [2:0] u_ca_in_533;
wire [2:0] u_ca_in_534;
wire [2:0] u_ca_in_535;
wire [2:0] u_ca_in_536;
wire [2:0] u_ca_in_537;
wire [2:0] u_ca_in_538;
wire [2:0] u_ca_in_539;
wire [2:0] u_ca_in_540;
wire [2:0] u_ca_in_541;
wire [2:0] u_ca_in_542;
wire [2:0] u_ca_in_543;
wire [2:0] u_ca_in_544;
wire [2:0] u_ca_in_545;
wire [2:0] u_ca_in_546;
wire [2:0] u_ca_in_547;
wire [2:0] u_ca_in_548;
wire [2:0] u_ca_in_549;
wire [2:0] u_ca_in_550;
wire [2:0] u_ca_in_551;
wire [2:0] u_ca_in_552;
wire [2:0] u_ca_in_553;
wire [2:0] u_ca_in_554;
wire [2:0] u_ca_in_555;
wire [2:0] u_ca_in_556;
wire [2:0] u_ca_in_557;
wire [2:0] u_ca_in_558;
wire [2:0] u_ca_in_559;
wire [2:0] u_ca_in_560;
wire [2:0] u_ca_in_561;
wire [2:0] u_ca_in_562;
wire [2:0] u_ca_in_563;
wire [2:0] u_ca_in_564;
wire [2:0] u_ca_in_565;
wire [2:0] u_ca_in_566;
wire [2:0] u_ca_in_567;
wire [2:0] u_ca_in_568;
wire [2:0] u_ca_in_569;
wire [2:0] u_ca_in_570;
wire [2:0] u_ca_in_571;
wire [2:0] u_ca_in_572;
wire [2:0] u_ca_in_573;
wire [2:0] u_ca_in_574;
wire [2:0] u_ca_in_575;
wire [2:0] u_ca_in_576;
wire [2:0] u_ca_in_577;
wire [2:0] u_ca_in_578;
wire [2:0] u_ca_in_579;
wire [2:0] u_ca_in_580;
wire [2:0] u_ca_in_581;
wire [2:0] u_ca_in_582;
wire [2:0] u_ca_in_583;
wire [2:0] u_ca_in_584;
wire [2:0] u_ca_in_585;
wire [2:0] u_ca_in_586;
wire [2:0] u_ca_in_587;
wire [2:0] u_ca_in_588;
wire [2:0] u_ca_in_589;
wire [2:0] u_ca_in_590;
wire [2:0] u_ca_in_591;
wire [2:0] u_ca_in_592;
wire [2:0] u_ca_in_593;
wire [2:0] u_ca_in_594;
wire [2:0] u_ca_in_595;
wire [2:0] u_ca_in_596;
wire [2:0] u_ca_in_597;
wire [2:0] u_ca_in_598;
wire [2:0] u_ca_in_599;
wire [2:0] u_ca_in_600;
wire [2:0] u_ca_in_601;
wire [2:0] u_ca_in_602;
wire [2:0] u_ca_in_603;
wire [2:0] u_ca_in_604;
wire [2:0] u_ca_in_605;
wire [2:0] u_ca_in_606;
wire [2:0] u_ca_in_607;
wire [2:0] u_ca_in_608;
wire [2:0] u_ca_in_609;
wire [2:0] u_ca_in_610;
wire [2:0] u_ca_in_611;
wire [2:0] u_ca_in_612;
wire [2:0] u_ca_in_613;
wire [2:0] u_ca_in_614;
wire [2:0] u_ca_in_615;
wire [2:0] u_ca_in_616;
wire [2:0] u_ca_in_617;
wire [2:0] u_ca_in_618;
wire [2:0] u_ca_in_619;
wire [2:0] u_ca_in_620;
wire [2:0] u_ca_in_621;
wire [2:0] u_ca_in_622;
wire [2:0] u_ca_in_623;
wire [2:0] u_ca_in_624;
wire [2:0] u_ca_in_625;
wire [2:0] u_ca_in_626;
wire [2:0] u_ca_in_627;
wire [2:0] u_ca_in_628;
wire [2:0] u_ca_in_629;
wire [2:0] u_ca_in_630;
wire [2:0] u_ca_in_631;
wire [2:0] u_ca_in_632;
wire [2:0] u_ca_in_633;
wire [2:0] u_ca_in_634;
wire [2:0] u_ca_in_635;
wire [2:0] u_ca_in_636;
wire [2:0] u_ca_in_637;
wire [2:0] u_ca_in_638;
wire [2:0] u_ca_in_639;
wire [2:0] u_ca_in_640;
wire [2:0] u_ca_in_641;
wire [2:0] u_ca_in_642;
wire [2:0] u_ca_in_643;
wire [2:0] u_ca_in_644;
wire [2:0] u_ca_in_645;
wire [2:0] u_ca_in_646;
wire [2:0] u_ca_in_647;
wire [2:0] u_ca_in_648;
wire [2:0] u_ca_in_649;
wire [2:0] u_ca_in_650;
wire [2:0] u_ca_in_651;
wire [2:0] u_ca_in_652;
wire [2:0] u_ca_in_653;
wire [2:0] u_ca_in_654;
wire [2:0] u_ca_in_655;
wire [2:0] u_ca_in_656;
wire [2:0] u_ca_in_657;
wire [2:0] u_ca_in_658;
wire [2:0] u_ca_in_659;
wire [2:0] u_ca_in_660;
wire [2:0] u_ca_in_661;
wire [2:0] u_ca_in_662;
wire [2:0] u_ca_in_663;
wire [2:0] u_ca_in_664;
wire [2:0] u_ca_in_665;
wire [2:0] u_ca_in_666;
wire [2:0] u_ca_in_667;
wire [2:0] u_ca_in_668;
wire [2:0] u_ca_in_669;
wire [2:0] u_ca_in_670;
wire [2:0] u_ca_in_671;
wire [2:0] u_ca_in_672;
wire [2:0] u_ca_in_673;
wire [2:0] u_ca_in_674;
wire [2:0] u_ca_in_675;
wire [2:0] u_ca_in_676;
wire [2:0] u_ca_in_677;
wire [2:0] u_ca_in_678;
wire [2:0] u_ca_in_679;
wire [2:0] u_ca_in_680;
wire [2:0] u_ca_in_681;
wire [2:0] u_ca_in_682;
wire [2:0] u_ca_in_683;
wire [2:0] u_ca_in_684;
wire [2:0] u_ca_in_685;
wire [2:0] u_ca_in_686;
wire [2:0] u_ca_in_687;
wire [2:0] u_ca_in_688;
wire [2:0] u_ca_in_689;
wire [2:0] u_ca_in_690;
wire [2:0] u_ca_in_691;
wire [2:0] u_ca_in_692;
wire [2:0] u_ca_in_693;
wire [2:0] u_ca_in_694;
wire [2:0] u_ca_in_695;
wire [2:0] u_ca_in_696;
wire [2:0] u_ca_in_697;
wire [2:0] u_ca_in_698;
wire [2:0] u_ca_in_699;
wire [2:0] u_ca_in_700;
wire [2:0] u_ca_in_701;
wire [2:0] u_ca_in_702;
wire [2:0] u_ca_in_703;
wire [2:0] u_ca_in_704;
wire [2:0] u_ca_in_705;
wire [2:0] u_ca_in_706;
wire [2:0] u_ca_in_707;
wire [2:0] u_ca_in_708;
wire [2:0] u_ca_in_709;
wire [2:0] u_ca_in_710;
wire [2:0] u_ca_in_711;
wire [2:0] u_ca_in_712;
wire [2:0] u_ca_in_713;
wire [2:0] u_ca_in_714;
wire [2:0] u_ca_in_715;
wire [2:0] u_ca_in_716;
wire [2:0] u_ca_in_717;
wire [2:0] u_ca_in_718;
wire [2:0] u_ca_in_719;
wire [2:0] u_ca_in_720;
wire [2:0] u_ca_in_721;
wire [2:0] u_ca_in_722;
wire [2:0] u_ca_in_723;
wire [2:0] u_ca_in_724;
wire [2:0] u_ca_in_725;
wire [2:0] u_ca_in_726;
wire [2:0] u_ca_in_727;
wire [2:0] u_ca_in_728;
wire [2:0] u_ca_in_729;
wire [2:0] u_ca_in_730;
wire [2:0] u_ca_in_731;
wire [2:0] u_ca_in_732;
wire [2:0] u_ca_in_733;
wire [2:0] u_ca_in_734;
wire [2:0] u_ca_in_735;
wire [2:0] u_ca_in_736;
wire [2:0] u_ca_in_737;
wire [2:0] u_ca_in_738;
wire [2:0] u_ca_in_739;
wire [2:0] u_ca_in_740;
wire [2:0] u_ca_in_741;
wire [2:0] u_ca_in_742;
wire [2:0] u_ca_in_743;
wire [2:0] u_ca_in_744;
wire [2:0] u_ca_in_745;
wire [2:0] u_ca_in_746;
wire [2:0] u_ca_in_747;
wire [2:0] u_ca_in_748;
wire [2:0] u_ca_in_749;
wire [2:0] u_ca_in_750;
wire [2:0] u_ca_in_751;
wire [2:0] u_ca_in_752;
wire [2:0] u_ca_in_753;
wire [2:0] u_ca_in_754;
wire [2:0] u_ca_in_755;
wire [2:0] u_ca_in_756;
wire [2:0] u_ca_in_757;
wire [2:0] u_ca_in_758;
wire [2:0] u_ca_in_759;
wire [2:0] u_ca_in_760;
wire [2:0] u_ca_in_761;
wire [2:0] u_ca_in_762;
wire [2:0] u_ca_in_763;
wire [2:0] u_ca_in_764;
wire [2:0] u_ca_in_765;
wire [2:0] u_ca_in_766;
wire [2:0] u_ca_in_767;
wire [2:0] u_ca_in_768;
wire [2:0] u_ca_in_769;
wire [2:0] u_ca_in_770;
wire [2:0] u_ca_in_771;
wire [2:0] u_ca_in_772;
wire [2:0] u_ca_in_773;
wire [2:0] u_ca_in_774;
wire [2:0] u_ca_in_775;
wire [2:0] u_ca_in_776;
wire [2:0] u_ca_in_777;
wire [2:0] u_ca_in_778;
wire [2:0] u_ca_in_779;
wire [2:0] u_ca_in_780;
wire [2:0] u_ca_in_781;
wire [2:0] u_ca_in_782;
wire [2:0] u_ca_in_783;
wire [2:0] u_ca_in_784;
wire [2:0] u_ca_in_785;
wire [2:0] u_ca_in_786;
wire [2:0] u_ca_in_787;
wire [2:0] u_ca_in_788;
wire [2:0] u_ca_in_789;
wire [2:0] u_ca_in_790;
wire [2:0] u_ca_in_791;
wire [2:0] u_ca_in_792;
wire [2:0] u_ca_in_793;
wire [2:0] u_ca_in_794;
wire [2:0] u_ca_in_795;
wire [2:0] u_ca_in_796;
wire [2:0] u_ca_in_797;
wire [2:0] u_ca_in_798;
wire [2:0] u_ca_in_799;
wire [2:0] u_ca_in_800;
wire [2:0] u_ca_in_801;
wire [2:0] u_ca_in_802;
wire [2:0] u_ca_in_803;
wire [2:0] u_ca_in_804;
wire [2:0] u_ca_in_805;
wire [2:0] u_ca_in_806;
wire [2:0] u_ca_in_807;
wire [2:0] u_ca_in_808;
wire [2:0] u_ca_in_809;
wire [2:0] u_ca_in_810;
wire [2:0] u_ca_in_811;
wire [2:0] u_ca_in_812;
wire [2:0] u_ca_in_813;
wire [2:0] u_ca_in_814;
wire [2:0] u_ca_in_815;
wire [2:0] u_ca_in_816;
wire [2:0] u_ca_in_817;
wire [2:0] u_ca_in_818;
wire [2:0] u_ca_in_819;
wire [2:0] u_ca_in_820;
wire [2:0] u_ca_in_821;
wire [2:0] u_ca_in_822;
wire [2:0] u_ca_in_823;
wire [2:0] u_ca_in_824;
wire [2:0] u_ca_in_825;
wire [2:0] u_ca_in_826;
wire [2:0] u_ca_in_827;
wire [2:0] u_ca_in_828;
wire [2:0] u_ca_in_829;
wire [2:0] u_ca_in_830;
wire [2:0] u_ca_in_831;
wire [2:0] u_ca_in_832;
wire [2:0] u_ca_in_833;
wire [2:0] u_ca_in_834;
wire [2:0] u_ca_in_835;
wire [2:0] u_ca_in_836;
wire [2:0] u_ca_in_837;
wire [2:0] u_ca_in_838;
wire [2:0] u_ca_in_839;
wire [2:0] u_ca_in_840;
wire [2:0] u_ca_in_841;
wire [2:0] u_ca_in_842;
wire [2:0] u_ca_in_843;
wire [2:0] u_ca_in_844;
wire [2:0] u_ca_in_845;
wire [2:0] u_ca_in_846;
wire [2:0] u_ca_in_847;
wire [2:0] u_ca_in_848;
wire [2:0] u_ca_in_849;
wire [2:0] u_ca_in_850;
wire [2:0] u_ca_in_851;
wire [2:0] u_ca_in_852;
wire [2:0] u_ca_in_853;
wire [2:0] u_ca_in_854;
wire [2:0] u_ca_in_855;
wire [2:0] u_ca_in_856;
wire [2:0] u_ca_in_857;
wire [2:0] u_ca_in_858;
wire [2:0] u_ca_in_859;
wire [2:0] u_ca_in_860;
wire [2:0] u_ca_in_861;
wire [2:0] u_ca_in_862;
wire [2:0] u_ca_in_863;
wire [2:0] u_ca_in_864;
wire [2:0] u_ca_in_865;
wire [2:0] u_ca_in_866;
wire [2:0] u_ca_in_867;
wire [2:0] u_ca_in_868;
wire [2:0] u_ca_in_869;
wire [2:0] u_ca_in_870;
wire [2:0] u_ca_in_871;
wire [2:0] u_ca_in_872;
wire [2:0] u_ca_in_873;
wire [2:0] u_ca_in_874;
wire [2:0] u_ca_in_875;
wire [2:0] u_ca_in_876;
wire [2:0] u_ca_in_877;
wire [2:0] u_ca_in_878;
wire [2:0] u_ca_in_879;
wire [2:0] u_ca_in_880;
wire [2:0] u_ca_in_881;
wire [2:0] u_ca_in_882;
wire [2:0] u_ca_in_883;
wire [2:0] u_ca_in_884;
wire [2:0] u_ca_in_885;
wire [2:0] u_ca_in_886;
wire [2:0] u_ca_in_887;
wire [2:0] u_ca_in_888;
wire [2:0] u_ca_in_889;
wire [2:0] u_ca_in_890;
wire [2:0] u_ca_in_891;
wire [2:0] u_ca_in_892;
wire [2:0] u_ca_in_893;
wire [2:0] u_ca_in_894;
wire [2:0] u_ca_in_895;
wire [2:0] u_ca_in_896;
wire [2:0] u_ca_in_897;
wire [2:0] u_ca_in_898;
wire [2:0] u_ca_in_899;
wire [2:0] u_ca_in_900;
wire [2:0] u_ca_in_901;
wire [2:0] u_ca_in_902;
wire [2:0] u_ca_in_903;
wire [2:0] u_ca_in_904;
wire [2:0] u_ca_in_905;
wire [2:0] u_ca_in_906;
wire [2:0] u_ca_in_907;
wire [2:0] u_ca_in_908;
wire [2:0] u_ca_in_909;
wire [2:0] u_ca_in_910;
wire [2:0] u_ca_in_911;
wire [2:0] u_ca_in_912;
wire [2:0] u_ca_in_913;
wire [2:0] u_ca_in_914;
wire [2:0] u_ca_in_915;
wire [2:0] u_ca_in_916;
wire [2:0] u_ca_in_917;
wire [2:0] u_ca_in_918;
wire [2:0] u_ca_in_919;
wire [2:0] u_ca_in_920;
wire [2:0] u_ca_in_921;
wire [2:0] u_ca_in_922;
wire [2:0] u_ca_in_923;
wire [2:0] u_ca_in_924;
wire [2:0] u_ca_in_925;
wire [2:0] u_ca_in_926;
wire [2:0] u_ca_in_927;
wire [2:0] u_ca_in_928;
wire [2:0] u_ca_in_929;
wire [2:0] u_ca_in_930;
wire [2:0] u_ca_in_931;
wire [2:0] u_ca_in_932;
wire [2:0] u_ca_in_933;
wire [2:0] u_ca_in_934;
wire [2:0] u_ca_in_935;
wire [2:0] u_ca_in_936;
wire [2:0] u_ca_in_937;
wire [2:0] u_ca_in_938;
wire [2:0] u_ca_in_939;
wire [2:0] u_ca_in_940;
wire [2:0] u_ca_in_941;
wire [2:0] u_ca_in_942;
wire [2:0] u_ca_in_943;
wire [2:0] u_ca_in_944;
wire [2:0] u_ca_in_945;
wire [2:0] u_ca_in_946;
wire [2:0] u_ca_in_947;
wire [2:0] u_ca_in_948;
wire [2:0] u_ca_in_949;
wire [2:0] u_ca_in_950;
wire [2:0] u_ca_in_951;
wire [2:0] u_ca_in_952;
wire [2:0] u_ca_in_953;
wire [2:0] u_ca_in_954;
wire [2:0] u_ca_in_955;
wire [2:0] u_ca_in_956;
wire [2:0] u_ca_in_957;
wire [2:0] u_ca_in_958;
wire [2:0] u_ca_in_959;
wire [2:0] u_ca_in_960;
wire [2:0] u_ca_in_961;
wire [2:0] u_ca_in_962;
wire [2:0] u_ca_in_963;
wire [2:0] u_ca_in_964;
wire [2:0] u_ca_in_965;
wire [2:0] u_ca_in_966;
wire [2:0] u_ca_in_967;
wire [2:0] u_ca_in_968;
wire [2:0] u_ca_in_969;
wire [2:0] u_ca_in_970;
wire [2:0] u_ca_in_971;
wire [2:0] u_ca_in_972;
wire [2:0] u_ca_in_973;
wire [2:0] u_ca_in_974;
wire [2:0] u_ca_in_975;
wire [2:0] u_ca_in_976;
wire [2:0] u_ca_in_977;
wire [2:0] u_ca_in_978;
wire [2:0] u_ca_in_979;
wire [2:0] u_ca_in_980;
wire [2:0] u_ca_in_981;
wire [2:0] u_ca_in_982;
wire [2:0] u_ca_in_983;
wire [2:0] u_ca_in_984;
wire [2:0] u_ca_in_985;
wire [2:0] u_ca_in_986;
wire [2:0] u_ca_in_987;
wire [2:0] u_ca_in_988;
wire [2:0] u_ca_in_989;
wire [2:0] u_ca_in_990;
wire [2:0] u_ca_in_991;
wire [2:0] u_ca_in_992;
wire [2:0] u_ca_in_993;
wire [2:0] u_ca_in_994;
wire [2:0] u_ca_in_995;
wire [2:0] u_ca_in_996;
wire [2:0] u_ca_in_997;
wire [2:0] u_ca_in_998;
wire [2:0] u_ca_in_999;
wire [2:0] u_ca_in_1000;
wire [2:0] u_ca_in_1001;
wire [2:0] u_ca_in_1002;
wire [2:0] u_ca_in_1003;
wire [2:0] u_ca_in_1004;
wire [2:0] u_ca_in_1005;
wire [2:0] u_ca_in_1006;
wire [2:0] u_ca_in_1007;
wire [2:0] u_ca_in_1008;
wire [2:0] u_ca_in_1009;
wire [2:0] u_ca_in_1010;
wire [2:0] u_ca_in_1011;
wire [2:0] u_ca_in_1012;
wire [2:0] u_ca_in_1013;
wire [2:0] u_ca_in_1014;
wire [2:0] u_ca_in_1015;
wire [2:0] u_ca_in_1016;
wire [2:0] u_ca_in_1017;
wire [2:0] u_ca_in_1018;
wire [2:0] u_ca_in_1019;
wire [2:0] u_ca_in_1020;
wire [2:0] u_ca_in_1021;
wire [2:0] u_ca_in_1022;
wire [2:0] u_ca_in_1023;


wire [1:0] u_ca_out_0;
wire [1:0] u_ca_out_1;
wire [1:0] u_ca_out_2;
wire [1:0] u_ca_out_3;
wire [1:0] u_ca_out_4;
wire [1:0] u_ca_out_5;
wire [1:0] u_ca_out_6;
wire [1:0] u_ca_out_7;
wire [1:0] u_ca_out_8;
wire [1:0] u_ca_out_9;
wire [1:0] u_ca_out_10;
wire [1:0] u_ca_out_11;
wire [1:0] u_ca_out_12;
wire [1:0] u_ca_out_13;
wire [1:0] u_ca_out_14;
wire [1:0] u_ca_out_15;
wire [1:0] u_ca_out_16;
wire [1:0] u_ca_out_17;
wire [1:0] u_ca_out_18;
wire [1:0] u_ca_out_19;
wire [1:0] u_ca_out_20;
wire [1:0] u_ca_out_21;
wire [1:0] u_ca_out_22;
wire [1:0] u_ca_out_23;
wire [1:0] u_ca_out_24;
wire [1:0] u_ca_out_25;
wire [1:0] u_ca_out_26;
wire [1:0] u_ca_out_27;
wire [1:0] u_ca_out_28;
wire [1:0] u_ca_out_29;
wire [1:0] u_ca_out_30;
wire [1:0] u_ca_out_31;
wire [1:0] u_ca_out_32;
wire [1:0] u_ca_out_33;
wire [1:0] u_ca_out_34;
wire [1:0] u_ca_out_35;
wire [1:0] u_ca_out_36;
wire [1:0] u_ca_out_37;
wire [1:0] u_ca_out_38;
wire [1:0] u_ca_out_39;
wire [1:0] u_ca_out_40;
wire [1:0] u_ca_out_41;
wire [1:0] u_ca_out_42;
wire [1:0] u_ca_out_43;
wire [1:0] u_ca_out_44;
wire [1:0] u_ca_out_45;
wire [1:0] u_ca_out_46;
wire [1:0] u_ca_out_47;
wire [1:0] u_ca_out_48;
wire [1:0] u_ca_out_49;
wire [1:0] u_ca_out_50;
wire [1:0] u_ca_out_51;
wire [1:0] u_ca_out_52;
wire [1:0] u_ca_out_53;
wire [1:0] u_ca_out_54;
wire [1:0] u_ca_out_55;
wire [1:0] u_ca_out_56;
wire [1:0] u_ca_out_57;
wire [1:0] u_ca_out_58;
wire [1:0] u_ca_out_59;
wire [1:0] u_ca_out_60;
wire [1:0] u_ca_out_61;
wire [1:0] u_ca_out_62;
wire [1:0] u_ca_out_63;
wire [1:0] u_ca_out_64;
wire [1:0] u_ca_out_65;
wire [1:0] u_ca_out_66;
wire [1:0] u_ca_out_67;
wire [1:0] u_ca_out_68;
wire [1:0] u_ca_out_69;
wire [1:0] u_ca_out_70;
wire [1:0] u_ca_out_71;
wire [1:0] u_ca_out_72;
wire [1:0] u_ca_out_73;
wire [1:0] u_ca_out_74;
wire [1:0] u_ca_out_75;
wire [1:0] u_ca_out_76;
wire [1:0] u_ca_out_77;
wire [1:0] u_ca_out_78;
wire [1:0] u_ca_out_79;
wire [1:0] u_ca_out_80;
wire [1:0] u_ca_out_81;
wire [1:0] u_ca_out_82;
wire [1:0] u_ca_out_83;
wire [1:0] u_ca_out_84;
wire [1:0] u_ca_out_85;
wire [1:0] u_ca_out_86;
wire [1:0] u_ca_out_87;
wire [1:0] u_ca_out_88;
wire [1:0] u_ca_out_89;
wire [1:0] u_ca_out_90;
wire [1:0] u_ca_out_91;
wire [1:0] u_ca_out_92;
wire [1:0] u_ca_out_93;
wire [1:0] u_ca_out_94;
wire [1:0] u_ca_out_95;
wire [1:0] u_ca_out_96;
wire [1:0] u_ca_out_97;
wire [1:0] u_ca_out_98;
wire [1:0] u_ca_out_99;
wire [1:0] u_ca_out_100;
wire [1:0] u_ca_out_101;
wire [1:0] u_ca_out_102;
wire [1:0] u_ca_out_103;
wire [1:0] u_ca_out_104;
wire [1:0] u_ca_out_105;
wire [1:0] u_ca_out_106;
wire [1:0] u_ca_out_107;
wire [1:0] u_ca_out_108;
wire [1:0] u_ca_out_109;
wire [1:0] u_ca_out_110;
wire [1:0] u_ca_out_111;
wire [1:0] u_ca_out_112;
wire [1:0] u_ca_out_113;
wire [1:0] u_ca_out_114;
wire [1:0] u_ca_out_115;
wire [1:0] u_ca_out_116;
wire [1:0] u_ca_out_117;
wire [1:0] u_ca_out_118;
wire [1:0] u_ca_out_119;
wire [1:0] u_ca_out_120;
wire [1:0] u_ca_out_121;
wire [1:0] u_ca_out_122;
wire [1:0] u_ca_out_123;
wire [1:0] u_ca_out_124;
wire [1:0] u_ca_out_125;
wire [1:0] u_ca_out_126;
wire [1:0] u_ca_out_127;
wire [1:0] u_ca_out_128;
wire [1:0] u_ca_out_129;
wire [1:0] u_ca_out_130;
wire [1:0] u_ca_out_131;
wire [1:0] u_ca_out_132;
wire [1:0] u_ca_out_133;
wire [1:0] u_ca_out_134;
wire [1:0] u_ca_out_135;
wire [1:0] u_ca_out_136;
wire [1:0] u_ca_out_137;
wire [1:0] u_ca_out_138;
wire [1:0] u_ca_out_139;
wire [1:0] u_ca_out_140;
wire [1:0] u_ca_out_141;
wire [1:0] u_ca_out_142;
wire [1:0] u_ca_out_143;
wire [1:0] u_ca_out_144;
wire [1:0] u_ca_out_145;
wire [1:0] u_ca_out_146;
wire [1:0] u_ca_out_147;
wire [1:0] u_ca_out_148;
wire [1:0] u_ca_out_149;
wire [1:0] u_ca_out_150;
wire [1:0] u_ca_out_151;
wire [1:0] u_ca_out_152;
wire [1:0] u_ca_out_153;
wire [1:0] u_ca_out_154;
wire [1:0] u_ca_out_155;
wire [1:0] u_ca_out_156;
wire [1:0] u_ca_out_157;
wire [1:0] u_ca_out_158;
wire [1:0] u_ca_out_159;
wire [1:0] u_ca_out_160;
wire [1:0] u_ca_out_161;
wire [1:0] u_ca_out_162;
wire [1:0] u_ca_out_163;
wire [1:0] u_ca_out_164;
wire [1:0] u_ca_out_165;
wire [1:0] u_ca_out_166;
wire [1:0] u_ca_out_167;
wire [1:0] u_ca_out_168;
wire [1:0] u_ca_out_169;
wire [1:0] u_ca_out_170;
wire [1:0] u_ca_out_171;
wire [1:0] u_ca_out_172;
wire [1:0] u_ca_out_173;
wire [1:0] u_ca_out_174;
wire [1:0] u_ca_out_175;
wire [1:0] u_ca_out_176;
wire [1:0] u_ca_out_177;
wire [1:0] u_ca_out_178;
wire [1:0] u_ca_out_179;
wire [1:0] u_ca_out_180;
wire [1:0] u_ca_out_181;
wire [1:0] u_ca_out_182;
wire [1:0] u_ca_out_183;
wire [1:0] u_ca_out_184;
wire [1:0] u_ca_out_185;
wire [1:0] u_ca_out_186;
wire [1:0] u_ca_out_187;
wire [1:0] u_ca_out_188;
wire [1:0] u_ca_out_189;
wire [1:0] u_ca_out_190;
wire [1:0] u_ca_out_191;
wire [1:0] u_ca_out_192;
wire [1:0] u_ca_out_193;
wire [1:0] u_ca_out_194;
wire [1:0] u_ca_out_195;
wire [1:0] u_ca_out_196;
wire [1:0] u_ca_out_197;
wire [1:0] u_ca_out_198;
wire [1:0] u_ca_out_199;
wire [1:0] u_ca_out_200;
wire [1:0] u_ca_out_201;
wire [1:0] u_ca_out_202;
wire [1:0] u_ca_out_203;
wire [1:0] u_ca_out_204;
wire [1:0] u_ca_out_205;
wire [1:0] u_ca_out_206;
wire [1:0] u_ca_out_207;
wire [1:0] u_ca_out_208;
wire [1:0] u_ca_out_209;
wire [1:0] u_ca_out_210;
wire [1:0] u_ca_out_211;
wire [1:0] u_ca_out_212;
wire [1:0] u_ca_out_213;
wire [1:0] u_ca_out_214;
wire [1:0] u_ca_out_215;
wire [1:0] u_ca_out_216;
wire [1:0] u_ca_out_217;
wire [1:0] u_ca_out_218;
wire [1:0] u_ca_out_219;
wire [1:0] u_ca_out_220;
wire [1:0] u_ca_out_221;
wire [1:0] u_ca_out_222;
wire [1:0] u_ca_out_223;
wire [1:0] u_ca_out_224;
wire [1:0] u_ca_out_225;
wire [1:0] u_ca_out_226;
wire [1:0] u_ca_out_227;
wire [1:0] u_ca_out_228;
wire [1:0] u_ca_out_229;
wire [1:0] u_ca_out_230;
wire [1:0] u_ca_out_231;
wire [1:0] u_ca_out_232;
wire [1:0] u_ca_out_233;
wire [1:0] u_ca_out_234;
wire [1:0] u_ca_out_235;
wire [1:0] u_ca_out_236;
wire [1:0] u_ca_out_237;
wire [1:0] u_ca_out_238;
wire [1:0] u_ca_out_239;
wire [1:0] u_ca_out_240;
wire [1:0] u_ca_out_241;
wire [1:0] u_ca_out_242;
wire [1:0] u_ca_out_243;
wire [1:0] u_ca_out_244;
wire [1:0] u_ca_out_245;
wire [1:0] u_ca_out_246;
wire [1:0] u_ca_out_247;
wire [1:0] u_ca_out_248;
wire [1:0] u_ca_out_249;
wire [1:0] u_ca_out_250;
wire [1:0] u_ca_out_251;
wire [1:0] u_ca_out_252;
wire [1:0] u_ca_out_253;
wire [1:0] u_ca_out_254;
wire [1:0] u_ca_out_255;
wire [1:0] u_ca_out_256;
wire [1:0] u_ca_out_257;
wire [1:0] u_ca_out_258;
wire [1:0] u_ca_out_259;
wire [1:0] u_ca_out_260;
wire [1:0] u_ca_out_261;
wire [1:0] u_ca_out_262;
wire [1:0] u_ca_out_263;
wire [1:0] u_ca_out_264;
wire [1:0] u_ca_out_265;
wire [1:0] u_ca_out_266;
wire [1:0] u_ca_out_267;
wire [1:0] u_ca_out_268;
wire [1:0] u_ca_out_269;
wire [1:0] u_ca_out_270;
wire [1:0] u_ca_out_271;
wire [1:0] u_ca_out_272;
wire [1:0] u_ca_out_273;
wire [1:0] u_ca_out_274;
wire [1:0] u_ca_out_275;
wire [1:0] u_ca_out_276;
wire [1:0] u_ca_out_277;
wire [1:0] u_ca_out_278;
wire [1:0] u_ca_out_279;
wire [1:0] u_ca_out_280;
wire [1:0] u_ca_out_281;
wire [1:0] u_ca_out_282;
wire [1:0] u_ca_out_283;
wire [1:0] u_ca_out_284;
wire [1:0] u_ca_out_285;
wire [1:0] u_ca_out_286;
wire [1:0] u_ca_out_287;
wire [1:0] u_ca_out_288;
wire [1:0] u_ca_out_289;
wire [1:0] u_ca_out_290;
wire [1:0] u_ca_out_291;
wire [1:0] u_ca_out_292;
wire [1:0] u_ca_out_293;
wire [1:0] u_ca_out_294;
wire [1:0] u_ca_out_295;
wire [1:0] u_ca_out_296;
wire [1:0] u_ca_out_297;
wire [1:0] u_ca_out_298;
wire [1:0] u_ca_out_299;
wire [1:0] u_ca_out_300;
wire [1:0] u_ca_out_301;
wire [1:0] u_ca_out_302;
wire [1:0] u_ca_out_303;
wire [1:0] u_ca_out_304;
wire [1:0] u_ca_out_305;
wire [1:0] u_ca_out_306;
wire [1:0] u_ca_out_307;
wire [1:0] u_ca_out_308;
wire [1:0] u_ca_out_309;
wire [1:0] u_ca_out_310;
wire [1:0] u_ca_out_311;
wire [1:0] u_ca_out_312;
wire [1:0] u_ca_out_313;
wire [1:0] u_ca_out_314;
wire [1:0] u_ca_out_315;
wire [1:0] u_ca_out_316;
wire [1:0] u_ca_out_317;
wire [1:0] u_ca_out_318;
wire [1:0] u_ca_out_319;
wire [1:0] u_ca_out_320;
wire [1:0] u_ca_out_321;
wire [1:0] u_ca_out_322;
wire [1:0] u_ca_out_323;
wire [1:0] u_ca_out_324;
wire [1:0] u_ca_out_325;
wire [1:0] u_ca_out_326;
wire [1:0] u_ca_out_327;
wire [1:0] u_ca_out_328;
wire [1:0] u_ca_out_329;
wire [1:0] u_ca_out_330;
wire [1:0] u_ca_out_331;
wire [1:0] u_ca_out_332;
wire [1:0] u_ca_out_333;
wire [1:0] u_ca_out_334;
wire [1:0] u_ca_out_335;
wire [1:0] u_ca_out_336;
wire [1:0] u_ca_out_337;
wire [1:0] u_ca_out_338;
wire [1:0] u_ca_out_339;
wire [1:0] u_ca_out_340;
wire [1:0] u_ca_out_341;
wire [1:0] u_ca_out_342;
wire [1:0] u_ca_out_343;
wire [1:0] u_ca_out_344;
wire [1:0] u_ca_out_345;
wire [1:0] u_ca_out_346;
wire [1:0] u_ca_out_347;
wire [1:0] u_ca_out_348;
wire [1:0] u_ca_out_349;
wire [1:0] u_ca_out_350;
wire [1:0] u_ca_out_351;
wire [1:0] u_ca_out_352;
wire [1:0] u_ca_out_353;
wire [1:0] u_ca_out_354;
wire [1:0] u_ca_out_355;
wire [1:0] u_ca_out_356;
wire [1:0] u_ca_out_357;
wire [1:0] u_ca_out_358;
wire [1:0] u_ca_out_359;
wire [1:0] u_ca_out_360;
wire [1:0] u_ca_out_361;
wire [1:0] u_ca_out_362;
wire [1:0] u_ca_out_363;
wire [1:0] u_ca_out_364;
wire [1:0] u_ca_out_365;
wire [1:0] u_ca_out_366;
wire [1:0] u_ca_out_367;
wire [1:0] u_ca_out_368;
wire [1:0] u_ca_out_369;
wire [1:0] u_ca_out_370;
wire [1:0] u_ca_out_371;
wire [1:0] u_ca_out_372;
wire [1:0] u_ca_out_373;
wire [1:0] u_ca_out_374;
wire [1:0] u_ca_out_375;
wire [1:0] u_ca_out_376;
wire [1:0] u_ca_out_377;
wire [1:0] u_ca_out_378;
wire [1:0] u_ca_out_379;
wire [1:0] u_ca_out_380;
wire [1:0] u_ca_out_381;
wire [1:0] u_ca_out_382;
wire [1:0] u_ca_out_383;
wire [1:0] u_ca_out_384;
wire [1:0] u_ca_out_385;
wire [1:0] u_ca_out_386;
wire [1:0] u_ca_out_387;
wire [1:0] u_ca_out_388;
wire [1:0] u_ca_out_389;
wire [1:0] u_ca_out_390;
wire [1:0] u_ca_out_391;
wire [1:0] u_ca_out_392;
wire [1:0] u_ca_out_393;
wire [1:0] u_ca_out_394;
wire [1:0] u_ca_out_395;
wire [1:0] u_ca_out_396;
wire [1:0] u_ca_out_397;
wire [1:0] u_ca_out_398;
wire [1:0] u_ca_out_399;
wire [1:0] u_ca_out_400;
wire [1:0] u_ca_out_401;
wire [1:0] u_ca_out_402;
wire [1:0] u_ca_out_403;
wire [1:0] u_ca_out_404;
wire [1:0] u_ca_out_405;
wire [1:0] u_ca_out_406;
wire [1:0] u_ca_out_407;
wire [1:0] u_ca_out_408;
wire [1:0] u_ca_out_409;
wire [1:0] u_ca_out_410;
wire [1:0] u_ca_out_411;
wire [1:0] u_ca_out_412;
wire [1:0] u_ca_out_413;
wire [1:0] u_ca_out_414;
wire [1:0] u_ca_out_415;
wire [1:0] u_ca_out_416;
wire [1:0] u_ca_out_417;
wire [1:0] u_ca_out_418;
wire [1:0] u_ca_out_419;
wire [1:0] u_ca_out_420;
wire [1:0] u_ca_out_421;
wire [1:0] u_ca_out_422;
wire [1:0] u_ca_out_423;
wire [1:0] u_ca_out_424;
wire [1:0] u_ca_out_425;
wire [1:0] u_ca_out_426;
wire [1:0] u_ca_out_427;
wire [1:0] u_ca_out_428;
wire [1:0] u_ca_out_429;
wire [1:0] u_ca_out_430;
wire [1:0] u_ca_out_431;
wire [1:0] u_ca_out_432;
wire [1:0] u_ca_out_433;
wire [1:0] u_ca_out_434;
wire [1:0] u_ca_out_435;
wire [1:0] u_ca_out_436;
wire [1:0] u_ca_out_437;
wire [1:0] u_ca_out_438;
wire [1:0] u_ca_out_439;
wire [1:0] u_ca_out_440;
wire [1:0] u_ca_out_441;
wire [1:0] u_ca_out_442;
wire [1:0] u_ca_out_443;
wire [1:0] u_ca_out_444;
wire [1:0] u_ca_out_445;
wire [1:0] u_ca_out_446;
wire [1:0] u_ca_out_447;
wire [1:0] u_ca_out_448;
wire [1:0] u_ca_out_449;
wire [1:0] u_ca_out_450;
wire [1:0] u_ca_out_451;
wire [1:0] u_ca_out_452;
wire [1:0] u_ca_out_453;
wire [1:0] u_ca_out_454;
wire [1:0] u_ca_out_455;
wire [1:0] u_ca_out_456;
wire [1:0] u_ca_out_457;
wire [1:0] u_ca_out_458;
wire [1:0] u_ca_out_459;
wire [1:0] u_ca_out_460;
wire [1:0] u_ca_out_461;
wire [1:0] u_ca_out_462;
wire [1:0] u_ca_out_463;
wire [1:0] u_ca_out_464;
wire [1:0] u_ca_out_465;
wire [1:0] u_ca_out_466;
wire [1:0] u_ca_out_467;
wire [1:0] u_ca_out_468;
wire [1:0] u_ca_out_469;
wire [1:0] u_ca_out_470;
wire [1:0] u_ca_out_471;
wire [1:0] u_ca_out_472;
wire [1:0] u_ca_out_473;
wire [1:0] u_ca_out_474;
wire [1:0] u_ca_out_475;
wire [1:0] u_ca_out_476;
wire [1:0] u_ca_out_477;
wire [1:0] u_ca_out_478;
wire [1:0] u_ca_out_479;
wire [1:0] u_ca_out_480;
wire [1:0] u_ca_out_481;
wire [1:0] u_ca_out_482;
wire [1:0] u_ca_out_483;
wire [1:0] u_ca_out_484;
wire [1:0] u_ca_out_485;
wire [1:0] u_ca_out_486;
wire [1:0] u_ca_out_487;
wire [1:0] u_ca_out_488;
wire [1:0] u_ca_out_489;
wire [1:0] u_ca_out_490;
wire [1:0] u_ca_out_491;
wire [1:0] u_ca_out_492;
wire [1:0] u_ca_out_493;
wire [1:0] u_ca_out_494;
wire [1:0] u_ca_out_495;
wire [1:0] u_ca_out_496;
wire [1:0] u_ca_out_497;
wire [1:0] u_ca_out_498;
wire [1:0] u_ca_out_499;
wire [1:0] u_ca_out_500;
wire [1:0] u_ca_out_501;
wire [1:0] u_ca_out_502;
wire [1:0] u_ca_out_503;
wire [1:0] u_ca_out_504;
wire [1:0] u_ca_out_505;
wire [1:0] u_ca_out_506;
wire [1:0] u_ca_out_507;
wire [1:0] u_ca_out_508;
wire [1:0] u_ca_out_509;
wire [1:0] u_ca_out_510;
wire [1:0] u_ca_out_511;
wire [1:0] u_ca_out_512;
wire [1:0] u_ca_out_513;
wire [1:0] u_ca_out_514;
wire [1:0] u_ca_out_515;
wire [1:0] u_ca_out_516;
wire [1:0] u_ca_out_517;
wire [1:0] u_ca_out_518;
wire [1:0] u_ca_out_519;
wire [1:0] u_ca_out_520;
wire [1:0] u_ca_out_521;
wire [1:0] u_ca_out_522;
wire [1:0] u_ca_out_523;
wire [1:0] u_ca_out_524;
wire [1:0] u_ca_out_525;
wire [1:0] u_ca_out_526;
wire [1:0] u_ca_out_527;
wire [1:0] u_ca_out_528;
wire [1:0] u_ca_out_529;
wire [1:0] u_ca_out_530;
wire [1:0] u_ca_out_531;
wire [1:0] u_ca_out_532;
wire [1:0] u_ca_out_533;
wire [1:0] u_ca_out_534;
wire [1:0] u_ca_out_535;
wire [1:0] u_ca_out_536;
wire [1:0] u_ca_out_537;
wire [1:0] u_ca_out_538;
wire [1:0] u_ca_out_539;
wire [1:0] u_ca_out_540;
wire [1:0] u_ca_out_541;
wire [1:0] u_ca_out_542;
wire [1:0] u_ca_out_543;
wire [1:0] u_ca_out_544;
wire [1:0] u_ca_out_545;
wire [1:0] u_ca_out_546;
wire [1:0] u_ca_out_547;
wire [1:0] u_ca_out_548;
wire [1:0] u_ca_out_549;
wire [1:0] u_ca_out_550;
wire [1:0] u_ca_out_551;
wire [1:0] u_ca_out_552;
wire [1:0] u_ca_out_553;
wire [1:0] u_ca_out_554;
wire [1:0] u_ca_out_555;
wire [1:0] u_ca_out_556;
wire [1:0] u_ca_out_557;
wire [1:0] u_ca_out_558;
wire [1:0] u_ca_out_559;
wire [1:0] u_ca_out_560;
wire [1:0] u_ca_out_561;
wire [1:0] u_ca_out_562;
wire [1:0] u_ca_out_563;
wire [1:0] u_ca_out_564;
wire [1:0] u_ca_out_565;
wire [1:0] u_ca_out_566;
wire [1:0] u_ca_out_567;
wire [1:0] u_ca_out_568;
wire [1:0] u_ca_out_569;
wire [1:0] u_ca_out_570;
wire [1:0] u_ca_out_571;
wire [1:0] u_ca_out_572;
wire [1:0] u_ca_out_573;
wire [1:0] u_ca_out_574;
wire [1:0] u_ca_out_575;
wire [1:0] u_ca_out_576;
wire [1:0] u_ca_out_577;
wire [1:0] u_ca_out_578;
wire [1:0] u_ca_out_579;
wire [1:0] u_ca_out_580;
wire [1:0] u_ca_out_581;
wire [1:0] u_ca_out_582;
wire [1:0] u_ca_out_583;
wire [1:0] u_ca_out_584;
wire [1:0] u_ca_out_585;
wire [1:0] u_ca_out_586;
wire [1:0] u_ca_out_587;
wire [1:0] u_ca_out_588;
wire [1:0] u_ca_out_589;
wire [1:0] u_ca_out_590;
wire [1:0] u_ca_out_591;
wire [1:0] u_ca_out_592;
wire [1:0] u_ca_out_593;
wire [1:0] u_ca_out_594;
wire [1:0] u_ca_out_595;
wire [1:0] u_ca_out_596;
wire [1:0] u_ca_out_597;
wire [1:0] u_ca_out_598;
wire [1:0] u_ca_out_599;
wire [1:0] u_ca_out_600;
wire [1:0] u_ca_out_601;
wire [1:0] u_ca_out_602;
wire [1:0] u_ca_out_603;
wire [1:0] u_ca_out_604;
wire [1:0] u_ca_out_605;
wire [1:0] u_ca_out_606;
wire [1:0] u_ca_out_607;
wire [1:0] u_ca_out_608;
wire [1:0] u_ca_out_609;
wire [1:0] u_ca_out_610;
wire [1:0] u_ca_out_611;
wire [1:0] u_ca_out_612;
wire [1:0] u_ca_out_613;
wire [1:0] u_ca_out_614;
wire [1:0] u_ca_out_615;
wire [1:0] u_ca_out_616;
wire [1:0] u_ca_out_617;
wire [1:0] u_ca_out_618;
wire [1:0] u_ca_out_619;
wire [1:0] u_ca_out_620;
wire [1:0] u_ca_out_621;
wire [1:0] u_ca_out_622;
wire [1:0] u_ca_out_623;
wire [1:0] u_ca_out_624;
wire [1:0] u_ca_out_625;
wire [1:0] u_ca_out_626;
wire [1:0] u_ca_out_627;
wire [1:0] u_ca_out_628;
wire [1:0] u_ca_out_629;
wire [1:0] u_ca_out_630;
wire [1:0] u_ca_out_631;
wire [1:0] u_ca_out_632;
wire [1:0] u_ca_out_633;
wire [1:0] u_ca_out_634;
wire [1:0] u_ca_out_635;
wire [1:0] u_ca_out_636;
wire [1:0] u_ca_out_637;
wire [1:0] u_ca_out_638;
wire [1:0] u_ca_out_639;
wire [1:0] u_ca_out_640;
wire [1:0] u_ca_out_641;
wire [1:0] u_ca_out_642;
wire [1:0] u_ca_out_643;
wire [1:0] u_ca_out_644;
wire [1:0] u_ca_out_645;
wire [1:0] u_ca_out_646;
wire [1:0] u_ca_out_647;
wire [1:0] u_ca_out_648;
wire [1:0] u_ca_out_649;
wire [1:0] u_ca_out_650;
wire [1:0] u_ca_out_651;
wire [1:0] u_ca_out_652;
wire [1:0] u_ca_out_653;
wire [1:0] u_ca_out_654;
wire [1:0] u_ca_out_655;
wire [1:0] u_ca_out_656;
wire [1:0] u_ca_out_657;
wire [1:0] u_ca_out_658;
wire [1:0] u_ca_out_659;
wire [1:0] u_ca_out_660;
wire [1:0] u_ca_out_661;
wire [1:0] u_ca_out_662;
wire [1:0] u_ca_out_663;
wire [1:0] u_ca_out_664;
wire [1:0] u_ca_out_665;
wire [1:0] u_ca_out_666;
wire [1:0] u_ca_out_667;
wire [1:0] u_ca_out_668;
wire [1:0] u_ca_out_669;
wire [1:0] u_ca_out_670;
wire [1:0] u_ca_out_671;
wire [1:0] u_ca_out_672;
wire [1:0] u_ca_out_673;
wire [1:0] u_ca_out_674;
wire [1:0] u_ca_out_675;
wire [1:0] u_ca_out_676;
wire [1:0] u_ca_out_677;
wire [1:0] u_ca_out_678;
wire [1:0] u_ca_out_679;
wire [1:0] u_ca_out_680;
wire [1:0] u_ca_out_681;
wire [1:0] u_ca_out_682;
wire [1:0] u_ca_out_683;
wire [1:0] u_ca_out_684;
wire [1:0] u_ca_out_685;
wire [1:0] u_ca_out_686;
wire [1:0] u_ca_out_687;
wire [1:0] u_ca_out_688;
wire [1:0] u_ca_out_689;
wire [1:0] u_ca_out_690;
wire [1:0] u_ca_out_691;
wire [1:0] u_ca_out_692;
wire [1:0] u_ca_out_693;
wire [1:0] u_ca_out_694;
wire [1:0] u_ca_out_695;
wire [1:0] u_ca_out_696;
wire [1:0] u_ca_out_697;
wire [1:0] u_ca_out_698;
wire [1:0] u_ca_out_699;
wire [1:0] u_ca_out_700;
wire [1:0] u_ca_out_701;
wire [1:0] u_ca_out_702;
wire [1:0] u_ca_out_703;
wire [1:0] u_ca_out_704;
wire [1:0] u_ca_out_705;
wire [1:0] u_ca_out_706;
wire [1:0] u_ca_out_707;
wire [1:0] u_ca_out_708;
wire [1:0] u_ca_out_709;
wire [1:0] u_ca_out_710;
wire [1:0] u_ca_out_711;
wire [1:0] u_ca_out_712;
wire [1:0] u_ca_out_713;
wire [1:0] u_ca_out_714;
wire [1:0] u_ca_out_715;
wire [1:0] u_ca_out_716;
wire [1:0] u_ca_out_717;
wire [1:0] u_ca_out_718;
wire [1:0] u_ca_out_719;
wire [1:0] u_ca_out_720;
wire [1:0] u_ca_out_721;
wire [1:0] u_ca_out_722;
wire [1:0] u_ca_out_723;
wire [1:0] u_ca_out_724;
wire [1:0] u_ca_out_725;
wire [1:0] u_ca_out_726;
wire [1:0] u_ca_out_727;
wire [1:0] u_ca_out_728;
wire [1:0] u_ca_out_729;
wire [1:0] u_ca_out_730;
wire [1:0] u_ca_out_731;
wire [1:0] u_ca_out_732;
wire [1:0] u_ca_out_733;
wire [1:0] u_ca_out_734;
wire [1:0] u_ca_out_735;
wire [1:0] u_ca_out_736;
wire [1:0] u_ca_out_737;
wire [1:0] u_ca_out_738;
wire [1:0] u_ca_out_739;
wire [1:0] u_ca_out_740;
wire [1:0] u_ca_out_741;
wire [1:0] u_ca_out_742;
wire [1:0] u_ca_out_743;
wire [1:0] u_ca_out_744;
wire [1:0] u_ca_out_745;
wire [1:0] u_ca_out_746;
wire [1:0] u_ca_out_747;
wire [1:0] u_ca_out_748;
wire [1:0] u_ca_out_749;
wire [1:0] u_ca_out_750;
wire [1:0] u_ca_out_751;
wire [1:0] u_ca_out_752;
wire [1:0] u_ca_out_753;
wire [1:0] u_ca_out_754;
wire [1:0] u_ca_out_755;
wire [1:0] u_ca_out_756;
wire [1:0] u_ca_out_757;
wire [1:0] u_ca_out_758;
wire [1:0] u_ca_out_759;
wire [1:0] u_ca_out_760;
wire [1:0] u_ca_out_761;
wire [1:0] u_ca_out_762;
wire [1:0] u_ca_out_763;
wire [1:0] u_ca_out_764;
wire [1:0] u_ca_out_765;
wire [1:0] u_ca_out_766;
wire [1:0] u_ca_out_767;
wire [1:0] u_ca_out_768;
wire [1:0] u_ca_out_769;
wire [1:0] u_ca_out_770;
wire [1:0] u_ca_out_771;
wire [1:0] u_ca_out_772;
wire [1:0] u_ca_out_773;
wire [1:0] u_ca_out_774;
wire [1:0] u_ca_out_775;
wire [1:0] u_ca_out_776;
wire [1:0] u_ca_out_777;
wire [1:0] u_ca_out_778;
wire [1:0] u_ca_out_779;
wire [1:0] u_ca_out_780;
wire [1:0] u_ca_out_781;
wire [1:0] u_ca_out_782;
wire [1:0] u_ca_out_783;
wire [1:0] u_ca_out_784;
wire [1:0] u_ca_out_785;
wire [1:0] u_ca_out_786;
wire [1:0] u_ca_out_787;
wire [1:0] u_ca_out_788;
wire [1:0] u_ca_out_789;
wire [1:0] u_ca_out_790;
wire [1:0] u_ca_out_791;
wire [1:0] u_ca_out_792;
wire [1:0] u_ca_out_793;
wire [1:0] u_ca_out_794;
wire [1:0] u_ca_out_795;
wire [1:0] u_ca_out_796;
wire [1:0] u_ca_out_797;
wire [1:0] u_ca_out_798;
wire [1:0] u_ca_out_799;
wire [1:0] u_ca_out_800;
wire [1:0] u_ca_out_801;
wire [1:0] u_ca_out_802;
wire [1:0] u_ca_out_803;
wire [1:0] u_ca_out_804;
wire [1:0] u_ca_out_805;
wire [1:0] u_ca_out_806;
wire [1:0] u_ca_out_807;
wire [1:0] u_ca_out_808;
wire [1:0] u_ca_out_809;
wire [1:0] u_ca_out_810;
wire [1:0] u_ca_out_811;
wire [1:0] u_ca_out_812;
wire [1:0] u_ca_out_813;
wire [1:0] u_ca_out_814;
wire [1:0] u_ca_out_815;
wire [1:0] u_ca_out_816;
wire [1:0] u_ca_out_817;
wire [1:0] u_ca_out_818;
wire [1:0] u_ca_out_819;
wire [1:0] u_ca_out_820;
wire [1:0] u_ca_out_821;
wire [1:0] u_ca_out_822;
wire [1:0] u_ca_out_823;
wire [1:0] u_ca_out_824;
wire [1:0] u_ca_out_825;
wire [1:0] u_ca_out_826;
wire [1:0] u_ca_out_827;
wire [1:0] u_ca_out_828;
wire [1:0] u_ca_out_829;
wire [1:0] u_ca_out_830;
wire [1:0] u_ca_out_831;
wire [1:0] u_ca_out_832;
wire [1:0] u_ca_out_833;
wire [1:0] u_ca_out_834;
wire [1:0] u_ca_out_835;
wire [1:0] u_ca_out_836;
wire [1:0] u_ca_out_837;
wire [1:0] u_ca_out_838;
wire [1:0] u_ca_out_839;
wire [1:0] u_ca_out_840;
wire [1:0] u_ca_out_841;
wire [1:0] u_ca_out_842;
wire [1:0] u_ca_out_843;
wire [1:0] u_ca_out_844;
wire [1:0] u_ca_out_845;
wire [1:0] u_ca_out_846;
wire [1:0] u_ca_out_847;
wire [1:0] u_ca_out_848;
wire [1:0] u_ca_out_849;
wire [1:0] u_ca_out_850;
wire [1:0] u_ca_out_851;
wire [1:0] u_ca_out_852;
wire [1:0] u_ca_out_853;
wire [1:0] u_ca_out_854;
wire [1:0] u_ca_out_855;
wire [1:0] u_ca_out_856;
wire [1:0] u_ca_out_857;
wire [1:0] u_ca_out_858;
wire [1:0] u_ca_out_859;
wire [1:0] u_ca_out_860;
wire [1:0] u_ca_out_861;
wire [1:0] u_ca_out_862;
wire [1:0] u_ca_out_863;
wire [1:0] u_ca_out_864;
wire [1:0] u_ca_out_865;
wire [1:0] u_ca_out_866;
wire [1:0] u_ca_out_867;
wire [1:0] u_ca_out_868;
wire [1:0] u_ca_out_869;
wire [1:0] u_ca_out_870;
wire [1:0] u_ca_out_871;
wire [1:0] u_ca_out_872;
wire [1:0] u_ca_out_873;
wire [1:0] u_ca_out_874;
wire [1:0] u_ca_out_875;
wire [1:0] u_ca_out_876;
wire [1:0] u_ca_out_877;
wire [1:0] u_ca_out_878;
wire [1:0] u_ca_out_879;
wire [1:0] u_ca_out_880;
wire [1:0] u_ca_out_881;
wire [1:0] u_ca_out_882;
wire [1:0] u_ca_out_883;
wire [1:0] u_ca_out_884;
wire [1:0] u_ca_out_885;
wire [1:0] u_ca_out_886;
wire [1:0] u_ca_out_887;
wire [1:0] u_ca_out_888;
wire [1:0] u_ca_out_889;
wire [1:0] u_ca_out_890;
wire [1:0] u_ca_out_891;
wire [1:0] u_ca_out_892;
wire [1:0] u_ca_out_893;
wire [1:0] u_ca_out_894;
wire [1:0] u_ca_out_895;
wire [1:0] u_ca_out_896;
wire [1:0] u_ca_out_897;
wire [1:0] u_ca_out_898;
wire [1:0] u_ca_out_899;
wire [1:0] u_ca_out_900;
wire [1:0] u_ca_out_901;
wire [1:0] u_ca_out_902;
wire [1:0] u_ca_out_903;
wire [1:0] u_ca_out_904;
wire [1:0] u_ca_out_905;
wire [1:0] u_ca_out_906;
wire [1:0] u_ca_out_907;
wire [1:0] u_ca_out_908;
wire [1:0] u_ca_out_909;
wire [1:0] u_ca_out_910;
wire [1:0] u_ca_out_911;
wire [1:0] u_ca_out_912;
wire [1:0] u_ca_out_913;
wire [1:0] u_ca_out_914;
wire [1:0] u_ca_out_915;
wire [1:0] u_ca_out_916;
wire [1:0] u_ca_out_917;
wire [1:0] u_ca_out_918;
wire [1:0] u_ca_out_919;
wire [1:0] u_ca_out_920;
wire [1:0] u_ca_out_921;
wire [1:0] u_ca_out_922;
wire [1:0] u_ca_out_923;
wire [1:0] u_ca_out_924;
wire [1:0] u_ca_out_925;
wire [1:0] u_ca_out_926;
wire [1:0] u_ca_out_927;
wire [1:0] u_ca_out_928;
wire [1:0] u_ca_out_929;
wire [1:0] u_ca_out_930;
wire [1:0] u_ca_out_931;
wire [1:0] u_ca_out_932;
wire [1:0] u_ca_out_933;
wire [1:0] u_ca_out_934;
wire [1:0] u_ca_out_935;
wire [1:0] u_ca_out_936;
wire [1:0] u_ca_out_937;
wire [1:0] u_ca_out_938;
wire [1:0] u_ca_out_939;
wire [1:0] u_ca_out_940;
wire [1:0] u_ca_out_941;
wire [1:0] u_ca_out_942;
wire [1:0] u_ca_out_943;
wire [1:0] u_ca_out_944;
wire [1:0] u_ca_out_945;
wire [1:0] u_ca_out_946;
wire [1:0] u_ca_out_947;
wire [1:0] u_ca_out_948;
wire [1:0] u_ca_out_949;
wire [1:0] u_ca_out_950;
wire [1:0] u_ca_out_951;
wire [1:0] u_ca_out_952;
wire [1:0] u_ca_out_953;
wire [1:0] u_ca_out_954;
wire [1:0] u_ca_out_955;
wire [1:0] u_ca_out_956;
wire [1:0] u_ca_out_957;
wire [1:0] u_ca_out_958;
wire [1:0] u_ca_out_959;
wire [1:0] u_ca_out_960;
wire [1:0] u_ca_out_961;
wire [1:0] u_ca_out_962;
wire [1:0] u_ca_out_963;
wire [1:0] u_ca_out_964;
wire [1:0] u_ca_out_965;
wire [1:0] u_ca_out_966;
wire [1:0] u_ca_out_967;
wire [1:0] u_ca_out_968;
wire [1:0] u_ca_out_969;
wire [1:0] u_ca_out_970;
wire [1:0] u_ca_out_971;
wire [1:0] u_ca_out_972;
wire [1:0] u_ca_out_973;
wire [1:0] u_ca_out_974;
wire [1:0] u_ca_out_975;
wire [1:0] u_ca_out_976;
wire [1:0] u_ca_out_977;
wire [1:0] u_ca_out_978;
wire [1:0] u_ca_out_979;
wire [1:0] u_ca_out_980;
wire [1:0] u_ca_out_981;
wire [1:0] u_ca_out_982;
wire [1:0] u_ca_out_983;
wire [1:0] u_ca_out_984;
wire [1:0] u_ca_out_985;
wire [1:0] u_ca_out_986;
wire [1:0] u_ca_out_987;
wire [1:0] u_ca_out_988;
wire [1:0] u_ca_out_989;
wire [1:0] u_ca_out_990;
wire [1:0] u_ca_out_991;
wire [1:0] u_ca_out_992;
wire [1:0] u_ca_out_993;
wire [1:0] u_ca_out_994;
wire [1:0] u_ca_out_995;
wire [1:0] u_ca_out_996;
wire [1:0] u_ca_out_997;
wire [1:0] u_ca_out_998;
wire [1:0] u_ca_out_999;
wire [1:0] u_ca_out_1000;
wire [1:0] u_ca_out_1001;
wire [1:0] u_ca_out_1002;
wire [1:0] u_ca_out_1003;
wire [1:0] u_ca_out_1004;
wire [1:0] u_ca_out_1005;
wire [1:0] u_ca_out_1006;
wire [1:0] u_ca_out_1007;
wire [1:0] u_ca_out_1008;
wire [1:0] u_ca_out_1009;
wire [1:0] u_ca_out_1010;
wire [1:0] u_ca_out_1011;
wire [1:0] u_ca_out_1012;
wire [1:0] u_ca_out_1013;
wire [1:0] u_ca_out_1014;
wire [1:0] u_ca_out_1015;
wire [1:0] u_ca_out_1016;
wire [1:0] u_ca_out_1017;
wire [1:0] u_ca_out_1018;
wire [1:0] u_ca_out_1019;
wire [1:0] u_ca_out_1020;
wire [1:0] u_ca_out_1021;
wire [1:0] u_ca_out_1022;
wire [1:0] u_ca_out_1023;

assign u_ca_in_0 = col_in_0;
assign u_ca_in_1 = col_in_1;
assign u_ca_in_2 = col_in_2;
assign u_ca_in_3 = col_in_3;
assign u_ca_in_4 = col_in_4;
assign u_ca_in_5 = col_in_5;
assign u_ca_in_6 = col_in_6;
assign u_ca_in_7 = col_in_7;
assign u_ca_in_8 = col_in_8;
assign u_ca_in_9 = col_in_9;
assign u_ca_in_10 = col_in_10;
assign u_ca_in_11 = col_in_11;
assign u_ca_in_12 = col_in_12;
assign u_ca_in_13 = col_in_13;
assign u_ca_in_14 = col_in_14;
assign u_ca_in_15 = col_in_15;
assign u_ca_in_16 = col_in_16;
assign u_ca_in_17 = col_in_17;
assign u_ca_in_18 = col_in_18;
assign u_ca_in_19 = col_in_19;
assign u_ca_in_20 = col_in_20;
assign u_ca_in_21 = col_in_21;
assign u_ca_in_22 = col_in_22;
assign u_ca_in_23 = col_in_23;
assign u_ca_in_24 = col_in_24;
assign u_ca_in_25 = col_in_25;
assign u_ca_in_26 = col_in_26;
assign u_ca_in_27 = col_in_27;
assign u_ca_in_28 = col_in_28;
assign u_ca_in_29 = col_in_29;
assign u_ca_in_30 = col_in_30;
assign u_ca_in_31 = col_in_31;
assign u_ca_in_32 = col_in_32;
assign u_ca_in_33 = col_in_33;
assign u_ca_in_34 = col_in_34;
assign u_ca_in_35 = col_in_35;
assign u_ca_in_36 = col_in_36;
assign u_ca_in_37 = col_in_37;
assign u_ca_in_38 = col_in_38;
assign u_ca_in_39 = col_in_39;
assign u_ca_in_40 = col_in_40;
assign u_ca_in_41 = col_in_41;
assign u_ca_in_42 = col_in_42;
assign u_ca_in_43 = col_in_43;
assign u_ca_in_44 = col_in_44;
assign u_ca_in_45 = col_in_45;
assign u_ca_in_46 = col_in_46;
assign u_ca_in_47 = col_in_47;
assign u_ca_in_48 = col_in_48;
assign u_ca_in_49 = col_in_49;
assign u_ca_in_50 = col_in_50;
assign u_ca_in_51 = col_in_51;
assign u_ca_in_52 = col_in_52;
assign u_ca_in_53 = col_in_53;
assign u_ca_in_54 = col_in_54;
assign u_ca_in_55 = col_in_55;
assign u_ca_in_56 = col_in_56;
assign u_ca_in_57 = col_in_57;
assign u_ca_in_58 = col_in_58;
assign u_ca_in_59 = col_in_59;
assign u_ca_in_60 = col_in_60;
assign u_ca_in_61 = col_in_61;
assign u_ca_in_62 = col_in_62;
assign u_ca_in_63 = col_in_63;
assign u_ca_in_64 = col_in_64;
assign u_ca_in_65 = col_in_65;
assign u_ca_in_66 = col_in_66;
assign u_ca_in_67 = col_in_67;
assign u_ca_in_68 = col_in_68;
assign u_ca_in_69 = col_in_69;
assign u_ca_in_70 = col_in_70;
assign u_ca_in_71 = col_in_71;
assign u_ca_in_72 = col_in_72;
assign u_ca_in_73 = col_in_73;
assign u_ca_in_74 = col_in_74;
assign u_ca_in_75 = col_in_75;
assign u_ca_in_76 = col_in_76;
assign u_ca_in_77 = col_in_77;
assign u_ca_in_78 = col_in_78;
assign u_ca_in_79 = col_in_79;
assign u_ca_in_80 = col_in_80;
assign u_ca_in_81 = col_in_81;
assign u_ca_in_82 = col_in_82;
assign u_ca_in_83 = col_in_83;
assign u_ca_in_84 = col_in_84;
assign u_ca_in_85 = col_in_85;
assign u_ca_in_86 = col_in_86;
assign u_ca_in_87 = col_in_87;
assign u_ca_in_88 = col_in_88;
assign u_ca_in_89 = col_in_89;
assign u_ca_in_90 = col_in_90;
assign u_ca_in_91 = col_in_91;
assign u_ca_in_92 = col_in_92;
assign u_ca_in_93 = col_in_93;
assign u_ca_in_94 = col_in_94;
assign u_ca_in_95 = col_in_95;
assign u_ca_in_96 = col_in_96;
assign u_ca_in_97 = col_in_97;
assign u_ca_in_98 = col_in_98;
assign u_ca_in_99 = col_in_99;
assign u_ca_in_100 = col_in_100;
assign u_ca_in_101 = col_in_101;
assign u_ca_in_102 = col_in_102;
assign u_ca_in_103 = col_in_103;
assign u_ca_in_104 = col_in_104;
assign u_ca_in_105 = col_in_105;
assign u_ca_in_106 = col_in_106;
assign u_ca_in_107 = col_in_107;
assign u_ca_in_108 = col_in_108;
assign u_ca_in_109 = col_in_109;
assign u_ca_in_110 = col_in_110;
assign u_ca_in_111 = col_in_111;
assign u_ca_in_112 = col_in_112;
assign u_ca_in_113 = col_in_113;
assign u_ca_in_114 = col_in_114;
assign u_ca_in_115 = col_in_115;
assign u_ca_in_116 = col_in_116;
assign u_ca_in_117 = col_in_117;
assign u_ca_in_118 = col_in_118;
assign u_ca_in_119 = col_in_119;
assign u_ca_in_120 = col_in_120;
assign u_ca_in_121 = col_in_121;
assign u_ca_in_122 = col_in_122;
assign u_ca_in_123 = col_in_123;
assign u_ca_in_124 = col_in_124;
assign u_ca_in_125 = col_in_125;
assign u_ca_in_126 = col_in_126;
assign u_ca_in_127 = col_in_127;
assign u_ca_in_128 = col_in_128;
assign u_ca_in_129 = col_in_129;
assign u_ca_in_130 = col_in_130;
assign u_ca_in_131 = col_in_131;
assign u_ca_in_132 = col_in_132;
assign u_ca_in_133 = col_in_133;
assign u_ca_in_134 = col_in_134;
assign u_ca_in_135 = col_in_135;
assign u_ca_in_136 = col_in_136;
assign u_ca_in_137 = col_in_137;
assign u_ca_in_138 = col_in_138;
assign u_ca_in_139 = col_in_139;
assign u_ca_in_140 = col_in_140;
assign u_ca_in_141 = col_in_141;
assign u_ca_in_142 = col_in_142;
assign u_ca_in_143 = col_in_143;
assign u_ca_in_144 = col_in_144;
assign u_ca_in_145 = col_in_145;
assign u_ca_in_146 = col_in_146;
assign u_ca_in_147 = col_in_147;
assign u_ca_in_148 = col_in_148;
assign u_ca_in_149 = col_in_149;
assign u_ca_in_150 = col_in_150;
assign u_ca_in_151 = col_in_151;
assign u_ca_in_152 = col_in_152;
assign u_ca_in_153 = col_in_153;
assign u_ca_in_154 = col_in_154;
assign u_ca_in_155 = col_in_155;
assign u_ca_in_156 = col_in_156;
assign u_ca_in_157 = col_in_157;
assign u_ca_in_158 = col_in_158;
assign u_ca_in_159 = col_in_159;
assign u_ca_in_160 = col_in_160;
assign u_ca_in_161 = col_in_161;
assign u_ca_in_162 = col_in_162;
assign u_ca_in_163 = col_in_163;
assign u_ca_in_164 = col_in_164;
assign u_ca_in_165 = col_in_165;
assign u_ca_in_166 = col_in_166;
assign u_ca_in_167 = col_in_167;
assign u_ca_in_168 = col_in_168;
assign u_ca_in_169 = col_in_169;
assign u_ca_in_170 = col_in_170;
assign u_ca_in_171 = col_in_171;
assign u_ca_in_172 = col_in_172;
assign u_ca_in_173 = col_in_173;
assign u_ca_in_174 = col_in_174;
assign u_ca_in_175 = col_in_175;
assign u_ca_in_176 = col_in_176;
assign u_ca_in_177 = col_in_177;
assign u_ca_in_178 = col_in_178;
assign u_ca_in_179 = col_in_179;
assign u_ca_in_180 = col_in_180;
assign u_ca_in_181 = col_in_181;
assign u_ca_in_182 = col_in_182;
assign u_ca_in_183 = col_in_183;
assign u_ca_in_184 = col_in_184;
assign u_ca_in_185 = col_in_185;
assign u_ca_in_186 = col_in_186;
assign u_ca_in_187 = col_in_187;
assign u_ca_in_188 = col_in_188;
assign u_ca_in_189 = col_in_189;
assign u_ca_in_190 = col_in_190;
assign u_ca_in_191 = col_in_191;
assign u_ca_in_192 = col_in_192;
assign u_ca_in_193 = col_in_193;
assign u_ca_in_194 = col_in_194;
assign u_ca_in_195 = col_in_195;
assign u_ca_in_196 = col_in_196;
assign u_ca_in_197 = col_in_197;
assign u_ca_in_198 = col_in_198;
assign u_ca_in_199 = col_in_199;
assign u_ca_in_200 = col_in_200;
assign u_ca_in_201 = col_in_201;
assign u_ca_in_202 = col_in_202;
assign u_ca_in_203 = col_in_203;
assign u_ca_in_204 = col_in_204;
assign u_ca_in_205 = col_in_205;
assign u_ca_in_206 = col_in_206;
assign u_ca_in_207 = col_in_207;
assign u_ca_in_208 = col_in_208;
assign u_ca_in_209 = col_in_209;
assign u_ca_in_210 = col_in_210;
assign u_ca_in_211 = col_in_211;
assign u_ca_in_212 = col_in_212;
assign u_ca_in_213 = col_in_213;
assign u_ca_in_214 = col_in_214;
assign u_ca_in_215 = col_in_215;
assign u_ca_in_216 = col_in_216;
assign u_ca_in_217 = col_in_217;
assign u_ca_in_218 = col_in_218;
assign u_ca_in_219 = col_in_219;
assign u_ca_in_220 = col_in_220;
assign u_ca_in_221 = col_in_221;
assign u_ca_in_222 = col_in_222;
assign u_ca_in_223 = col_in_223;
assign u_ca_in_224 = col_in_224;
assign u_ca_in_225 = col_in_225;
assign u_ca_in_226 = col_in_226;
assign u_ca_in_227 = col_in_227;
assign u_ca_in_228 = col_in_228;
assign u_ca_in_229 = col_in_229;
assign u_ca_in_230 = col_in_230;
assign u_ca_in_231 = col_in_231;
assign u_ca_in_232 = col_in_232;
assign u_ca_in_233 = col_in_233;
assign u_ca_in_234 = col_in_234;
assign u_ca_in_235 = col_in_235;
assign u_ca_in_236 = col_in_236;
assign u_ca_in_237 = col_in_237;
assign u_ca_in_238 = col_in_238;
assign u_ca_in_239 = col_in_239;
assign u_ca_in_240 = col_in_240;
assign u_ca_in_241 = col_in_241;
assign u_ca_in_242 = col_in_242;
assign u_ca_in_243 = col_in_243;
assign u_ca_in_244 = col_in_244;
assign u_ca_in_245 = col_in_245;
assign u_ca_in_246 = col_in_246;
assign u_ca_in_247 = col_in_247;
assign u_ca_in_248 = col_in_248;
assign u_ca_in_249 = col_in_249;
assign u_ca_in_250 = col_in_250;
assign u_ca_in_251 = col_in_251;
assign u_ca_in_252 = col_in_252;
assign u_ca_in_253 = col_in_253;
assign u_ca_in_254 = col_in_254;
assign u_ca_in_255 = col_in_255;
assign u_ca_in_256 = col_in_256;
assign u_ca_in_257 = col_in_257;
assign u_ca_in_258 = col_in_258;
assign u_ca_in_259 = col_in_259;
assign u_ca_in_260 = col_in_260;
assign u_ca_in_261 = col_in_261;
assign u_ca_in_262 = col_in_262;
assign u_ca_in_263 = col_in_263;
assign u_ca_in_264 = col_in_264;
assign u_ca_in_265 = col_in_265;
assign u_ca_in_266 = col_in_266;
assign u_ca_in_267 = col_in_267;
assign u_ca_in_268 = col_in_268;
assign u_ca_in_269 = col_in_269;
assign u_ca_in_270 = col_in_270;
assign u_ca_in_271 = col_in_271;
assign u_ca_in_272 = col_in_272;
assign u_ca_in_273 = col_in_273;
assign u_ca_in_274 = col_in_274;
assign u_ca_in_275 = col_in_275;
assign u_ca_in_276 = col_in_276;
assign u_ca_in_277 = col_in_277;
assign u_ca_in_278 = col_in_278;
assign u_ca_in_279 = col_in_279;
assign u_ca_in_280 = col_in_280;
assign u_ca_in_281 = col_in_281;
assign u_ca_in_282 = col_in_282;
assign u_ca_in_283 = col_in_283;
assign u_ca_in_284 = col_in_284;
assign u_ca_in_285 = col_in_285;
assign u_ca_in_286 = col_in_286;
assign u_ca_in_287 = col_in_287;
assign u_ca_in_288 = col_in_288;
assign u_ca_in_289 = col_in_289;
assign u_ca_in_290 = col_in_290;
assign u_ca_in_291 = col_in_291;
assign u_ca_in_292 = col_in_292;
assign u_ca_in_293 = col_in_293;
assign u_ca_in_294 = col_in_294;
assign u_ca_in_295 = col_in_295;
assign u_ca_in_296 = col_in_296;
assign u_ca_in_297 = col_in_297;
assign u_ca_in_298 = col_in_298;
assign u_ca_in_299 = col_in_299;
assign u_ca_in_300 = col_in_300;
assign u_ca_in_301 = col_in_301;
assign u_ca_in_302 = col_in_302;
assign u_ca_in_303 = col_in_303;
assign u_ca_in_304 = col_in_304;
assign u_ca_in_305 = col_in_305;
assign u_ca_in_306 = col_in_306;
assign u_ca_in_307 = col_in_307;
assign u_ca_in_308 = col_in_308;
assign u_ca_in_309 = col_in_309;
assign u_ca_in_310 = col_in_310;
assign u_ca_in_311 = col_in_311;
assign u_ca_in_312 = col_in_312;
assign u_ca_in_313 = col_in_313;
assign u_ca_in_314 = col_in_314;
assign u_ca_in_315 = col_in_315;
assign u_ca_in_316 = col_in_316;
assign u_ca_in_317 = col_in_317;
assign u_ca_in_318 = col_in_318;
assign u_ca_in_319 = col_in_319;
assign u_ca_in_320 = col_in_320;
assign u_ca_in_321 = col_in_321;
assign u_ca_in_322 = col_in_322;
assign u_ca_in_323 = col_in_323;
assign u_ca_in_324 = col_in_324;
assign u_ca_in_325 = col_in_325;
assign u_ca_in_326 = col_in_326;
assign u_ca_in_327 = col_in_327;
assign u_ca_in_328 = col_in_328;
assign u_ca_in_329 = col_in_329;
assign u_ca_in_330 = col_in_330;
assign u_ca_in_331 = col_in_331;
assign u_ca_in_332 = col_in_332;
assign u_ca_in_333 = col_in_333;
assign u_ca_in_334 = col_in_334;
assign u_ca_in_335 = col_in_335;
assign u_ca_in_336 = col_in_336;
assign u_ca_in_337 = col_in_337;
assign u_ca_in_338 = col_in_338;
assign u_ca_in_339 = col_in_339;
assign u_ca_in_340 = col_in_340;
assign u_ca_in_341 = col_in_341;
assign u_ca_in_342 = col_in_342;
assign u_ca_in_343 = col_in_343;
assign u_ca_in_344 = col_in_344;
assign u_ca_in_345 = col_in_345;
assign u_ca_in_346 = col_in_346;
assign u_ca_in_347 = col_in_347;
assign u_ca_in_348 = col_in_348;
assign u_ca_in_349 = col_in_349;
assign u_ca_in_350 = col_in_350;
assign u_ca_in_351 = col_in_351;
assign u_ca_in_352 = col_in_352;
assign u_ca_in_353 = col_in_353;
assign u_ca_in_354 = col_in_354;
assign u_ca_in_355 = col_in_355;
assign u_ca_in_356 = col_in_356;
assign u_ca_in_357 = col_in_357;
assign u_ca_in_358 = col_in_358;
assign u_ca_in_359 = col_in_359;
assign u_ca_in_360 = col_in_360;
assign u_ca_in_361 = col_in_361;
assign u_ca_in_362 = col_in_362;
assign u_ca_in_363 = col_in_363;
assign u_ca_in_364 = col_in_364;
assign u_ca_in_365 = col_in_365;
assign u_ca_in_366 = col_in_366;
assign u_ca_in_367 = col_in_367;
assign u_ca_in_368 = col_in_368;
assign u_ca_in_369 = col_in_369;
assign u_ca_in_370 = col_in_370;
assign u_ca_in_371 = col_in_371;
assign u_ca_in_372 = col_in_372;
assign u_ca_in_373 = col_in_373;
assign u_ca_in_374 = col_in_374;
assign u_ca_in_375 = col_in_375;
assign u_ca_in_376 = col_in_376;
assign u_ca_in_377 = col_in_377;
assign u_ca_in_378 = col_in_378;
assign u_ca_in_379 = col_in_379;
assign u_ca_in_380 = col_in_380;
assign u_ca_in_381 = col_in_381;
assign u_ca_in_382 = col_in_382;
assign u_ca_in_383 = col_in_383;
assign u_ca_in_384 = col_in_384;
assign u_ca_in_385 = col_in_385;
assign u_ca_in_386 = col_in_386;
assign u_ca_in_387 = col_in_387;
assign u_ca_in_388 = col_in_388;
assign u_ca_in_389 = col_in_389;
assign u_ca_in_390 = col_in_390;
assign u_ca_in_391 = col_in_391;
assign u_ca_in_392 = col_in_392;
assign u_ca_in_393 = col_in_393;
assign u_ca_in_394 = col_in_394;
assign u_ca_in_395 = col_in_395;
assign u_ca_in_396 = col_in_396;
assign u_ca_in_397 = col_in_397;
assign u_ca_in_398 = col_in_398;
assign u_ca_in_399 = col_in_399;
assign u_ca_in_400 = col_in_400;
assign u_ca_in_401 = col_in_401;
assign u_ca_in_402 = col_in_402;
assign u_ca_in_403 = col_in_403;
assign u_ca_in_404 = col_in_404;
assign u_ca_in_405 = col_in_405;
assign u_ca_in_406 = col_in_406;
assign u_ca_in_407 = col_in_407;
assign u_ca_in_408 = col_in_408;
assign u_ca_in_409 = col_in_409;
assign u_ca_in_410 = col_in_410;
assign u_ca_in_411 = col_in_411;
assign u_ca_in_412 = col_in_412;
assign u_ca_in_413 = col_in_413;
assign u_ca_in_414 = col_in_414;
assign u_ca_in_415 = col_in_415;
assign u_ca_in_416 = col_in_416;
assign u_ca_in_417 = col_in_417;
assign u_ca_in_418 = col_in_418;
assign u_ca_in_419 = col_in_419;
assign u_ca_in_420 = col_in_420;
assign u_ca_in_421 = col_in_421;
assign u_ca_in_422 = col_in_422;
assign u_ca_in_423 = col_in_423;
assign u_ca_in_424 = col_in_424;
assign u_ca_in_425 = col_in_425;
assign u_ca_in_426 = col_in_426;
assign u_ca_in_427 = col_in_427;
assign u_ca_in_428 = col_in_428;
assign u_ca_in_429 = col_in_429;
assign u_ca_in_430 = col_in_430;
assign u_ca_in_431 = col_in_431;
assign u_ca_in_432 = col_in_432;
assign u_ca_in_433 = col_in_433;
assign u_ca_in_434 = col_in_434;
assign u_ca_in_435 = col_in_435;
assign u_ca_in_436 = col_in_436;
assign u_ca_in_437 = col_in_437;
assign u_ca_in_438 = col_in_438;
assign u_ca_in_439 = col_in_439;
assign u_ca_in_440 = col_in_440;
assign u_ca_in_441 = col_in_441;
assign u_ca_in_442 = col_in_442;
assign u_ca_in_443 = col_in_443;
assign u_ca_in_444 = col_in_444;
assign u_ca_in_445 = col_in_445;
assign u_ca_in_446 = col_in_446;
assign u_ca_in_447 = col_in_447;
assign u_ca_in_448 = col_in_448;
assign u_ca_in_449 = col_in_449;
assign u_ca_in_450 = col_in_450;
assign u_ca_in_451 = col_in_451;
assign u_ca_in_452 = col_in_452;
assign u_ca_in_453 = col_in_453;
assign u_ca_in_454 = col_in_454;
assign u_ca_in_455 = col_in_455;
assign u_ca_in_456 = col_in_456;
assign u_ca_in_457 = col_in_457;
assign u_ca_in_458 = col_in_458;
assign u_ca_in_459 = col_in_459;
assign u_ca_in_460 = col_in_460;
assign u_ca_in_461 = col_in_461;
assign u_ca_in_462 = col_in_462;
assign u_ca_in_463 = col_in_463;
assign u_ca_in_464 = col_in_464;
assign u_ca_in_465 = col_in_465;
assign u_ca_in_466 = col_in_466;
assign u_ca_in_467 = col_in_467;
assign u_ca_in_468 = col_in_468;
assign u_ca_in_469 = col_in_469;
assign u_ca_in_470 = col_in_470;
assign u_ca_in_471 = col_in_471;
assign u_ca_in_472 = col_in_472;
assign u_ca_in_473 = col_in_473;
assign u_ca_in_474 = col_in_474;
assign u_ca_in_475 = col_in_475;
assign u_ca_in_476 = col_in_476;
assign u_ca_in_477 = col_in_477;
assign u_ca_in_478 = col_in_478;
assign u_ca_in_479 = col_in_479;
assign u_ca_in_480 = col_in_480;
assign u_ca_in_481 = col_in_481;
assign u_ca_in_482 = col_in_482;
assign u_ca_in_483 = col_in_483;
assign u_ca_in_484 = col_in_484;
assign u_ca_in_485 = col_in_485;
assign u_ca_in_486 = col_in_486;
assign u_ca_in_487 = col_in_487;
assign u_ca_in_488 = col_in_488;
assign u_ca_in_489 = col_in_489;
assign u_ca_in_490 = col_in_490;
assign u_ca_in_491 = col_in_491;
assign u_ca_in_492 = col_in_492;
assign u_ca_in_493 = col_in_493;
assign u_ca_in_494 = col_in_494;
assign u_ca_in_495 = col_in_495;
assign u_ca_in_496 = col_in_496;
assign u_ca_in_497 = col_in_497;
assign u_ca_in_498 = col_in_498;
assign u_ca_in_499 = col_in_499;
assign u_ca_in_500 = col_in_500;
assign u_ca_in_501 = col_in_501;
assign u_ca_in_502 = col_in_502;
assign u_ca_in_503 = col_in_503;
assign u_ca_in_504 = col_in_504;
assign u_ca_in_505 = col_in_505;
assign u_ca_in_506 = col_in_506;
assign u_ca_in_507 = col_in_507;
assign u_ca_in_508 = col_in_508;
assign u_ca_in_509 = col_in_509;
assign u_ca_in_510 = col_in_510;
assign u_ca_in_511 = col_in_511;
assign u_ca_in_512 = col_in_512;
assign u_ca_in_513 = col_in_513;
assign u_ca_in_514 = col_in_514;
assign u_ca_in_515 = col_in_515;
assign u_ca_in_516 = col_in_516;
assign u_ca_in_517 = col_in_517;
assign u_ca_in_518 = col_in_518;
assign u_ca_in_519 = col_in_519;
assign u_ca_in_520 = col_in_520;
assign u_ca_in_521 = col_in_521;
assign u_ca_in_522 = col_in_522;
assign u_ca_in_523 = col_in_523;
assign u_ca_in_524 = col_in_524;
assign u_ca_in_525 = col_in_525;
assign u_ca_in_526 = col_in_526;
assign u_ca_in_527 = col_in_527;
assign u_ca_in_528 = col_in_528;
assign u_ca_in_529 = col_in_529;
assign u_ca_in_530 = col_in_530;
assign u_ca_in_531 = col_in_531;
assign u_ca_in_532 = col_in_532;
assign u_ca_in_533 = col_in_533;
assign u_ca_in_534 = col_in_534;
assign u_ca_in_535 = col_in_535;
assign u_ca_in_536 = col_in_536;
assign u_ca_in_537 = col_in_537;
assign u_ca_in_538 = col_in_538;
assign u_ca_in_539 = col_in_539;
assign u_ca_in_540 = col_in_540;
assign u_ca_in_541 = col_in_541;
assign u_ca_in_542 = col_in_542;
assign u_ca_in_543 = col_in_543;
assign u_ca_in_544 = col_in_544;
assign u_ca_in_545 = col_in_545;
assign u_ca_in_546 = col_in_546;
assign u_ca_in_547 = col_in_547;
assign u_ca_in_548 = col_in_548;
assign u_ca_in_549 = col_in_549;
assign u_ca_in_550 = col_in_550;
assign u_ca_in_551 = col_in_551;
assign u_ca_in_552 = col_in_552;
assign u_ca_in_553 = col_in_553;
assign u_ca_in_554 = col_in_554;
assign u_ca_in_555 = col_in_555;
assign u_ca_in_556 = col_in_556;
assign u_ca_in_557 = col_in_557;
assign u_ca_in_558 = col_in_558;
assign u_ca_in_559 = col_in_559;
assign u_ca_in_560 = col_in_560;
assign u_ca_in_561 = col_in_561;
assign u_ca_in_562 = col_in_562;
assign u_ca_in_563 = col_in_563;
assign u_ca_in_564 = col_in_564;
assign u_ca_in_565 = col_in_565;
assign u_ca_in_566 = col_in_566;
assign u_ca_in_567 = col_in_567;
assign u_ca_in_568 = col_in_568;
assign u_ca_in_569 = col_in_569;
assign u_ca_in_570 = col_in_570;
assign u_ca_in_571 = col_in_571;
assign u_ca_in_572 = col_in_572;
assign u_ca_in_573 = col_in_573;
assign u_ca_in_574 = col_in_574;
assign u_ca_in_575 = col_in_575;
assign u_ca_in_576 = col_in_576;
assign u_ca_in_577 = col_in_577;
assign u_ca_in_578 = col_in_578;
assign u_ca_in_579 = col_in_579;
assign u_ca_in_580 = col_in_580;
assign u_ca_in_581 = col_in_581;
assign u_ca_in_582 = col_in_582;
assign u_ca_in_583 = col_in_583;
assign u_ca_in_584 = col_in_584;
assign u_ca_in_585 = col_in_585;
assign u_ca_in_586 = col_in_586;
assign u_ca_in_587 = col_in_587;
assign u_ca_in_588 = col_in_588;
assign u_ca_in_589 = col_in_589;
assign u_ca_in_590 = col_in_590;
assign u_ca_in_591 = col_in_591;
assign u_ca_in_592 = col_in_592;
assign u_ca_in_593 = col_in_593;
assign u_ca_in_594 = col_in_594;
assign u_ca_in_595 = col_in_595;
assign u_ca_in_596 = col_in_596;
assign u_ca_in_597 = col_in_597;
assign u_ca_in_598 = col_in_598;
assign u_ca_in_599 = col_in_599;
assign u_ca_in_600 = col_in_600;
assign u_ca_in_601 = col_in_601;
assign u_ca_in_602 = col_in_602;
assign u_ca_in_603 = col_in_603;
assign u_ca_in_604 = col_in_604;
assign u_ca_in_605 = col_in_605;
assign u_ca_in_606 = col_in_606;
assign u_ca_in_607 = col_in_607;
assign u_ca_in_608 = col_in_608;
assign u_ca_in_609 = col_in_609;
assign u_ca_in_610 = col_in_610;
assign u_ca_in_611 = col_in_611;
assign u_ca_in_612 = col_in_612;
assign u_ca_in_613 = col_in_613;
assign u_ca_in_614 = col_in_614;
assign u_ca_in_615 = col_in_615;
assign u_ca_in_616 = col_in_616;
assign u_ca_in_617 = col_in_617;
assign u_ca_in_618 = col_in_618;
assign u_ca_in_619 = col_in_619;
assign u_ca_in_620 = col_in_620;
assign u_ca_in_621 = col_in_621;
assign u_ca_in_622 = col_in_622;
assign u_ca_in_623 = col_in_623;
assign u_ca_in_624 = col_in_624;
assign u_ca_in_625 = col_in_625;
assign u_ca_in_626 = col_in_626;
assign u_ca_in_627 = col_in_627;
assign u_ca_in_628 = col_in_628;
assign u_ca_in_629 = col_in_629;
assign u_ca_in_630 = col_in_630;
assign u_ca_in_631 = col_in_631;
assign u_ca_in_632 = col_in_632;
assign u_ca_in_633 = col_in_633;
assign u_ca_in_634 = col_in_634;
assign u_ca_in_635 = col_in_635;
assign u_ca_in_636 = col_in_636;
assign u_ca_in_637 = col_in_637;
assign u_ca_in_638 = col_in_638;
assign u_ca_in_639 = col_in_639;
assign u_ca_in_640 = col_in_640;
assign u_ca_in_641 = col_in_641;
assign u_ca_in_642 = col_in_642;
assign u_ca_in_643 = col_in_643;
assign u_ca_in_644 = col_in_644;
assign u_ca_in_645 = col_in_645;
assign u_ca_in_646 = col_in_646;
assign u_ca_in_647 = col_in_647;
assign u_ca_in_648 = col_in_648;
assign u_ca_in_649 = col_in_649;
assign u_ca_in_650 = col_in_650;
assign u_ca_in_651 = col_in_651;
assign u_ca_in_652 = col_in_652;
assign u_ca_in_653 = col_in_653;
assign u_ca_in_654 = col_in_654;
assign u_ca_in_655 = col_in_655;
assign u_ca_in_656 = col_in_656;
assign u_ca_in_657 = col_in_657;
assign u_ca_in_658 = col_in_658;
assign u_ca_in_659 = col_in_659;
assign u_ca_in_660 = col_in_660;
assign u_ca_in_661 = col_in_661;
assign u_ca_in_662 = col_in_662;
assign u_ca_in_663 = col_in_663;
assign u_ca_in_664 = col_in_664;
assign u_ca_in_665 = col_in_665;
assign u_ca_in_666 = col_in_666;
assign u_ca_in_667 = col_in_667;
assign u_ca_in_668 = col_in_668;
assign u_ca_in_669 = col_in_669;
assign u_ca_in_670 = col_in_670;
assign u_ca_in_671 = col_in_671;
assign u_ca_in_672 = col_in_672;
assign u_ca_in_673 = col_in_673;
assign u_ca_in_674 = col_in_674;
assign u_ca_in_675 = col_in_675;
assign u_ca_in_676 = col_in_676;
assign u_ca_in_677 = col_in_677;
assign u_ca_in_678 = col_in_678;
assign u_ca_in_679 = col_in_679;
assign u_ca_in_680 = col_in_680;
assign u_ca_in_681 = col_in_681;
assign u_ca_in_682 = col_in_682;
assign u_ca_in_683 = col_in_683;
assign u_ca_in_684 = col_in_684;
assign u_ca_in_685 = col_in_685;
assign u_ca_in_686 = col_in_686;
assign u_ca_in_687 = col_in_687;
assign u_ca_in_688 = col_in_688;
assign u_ca_in_689 = col_in_689;
assign u_ca_in_690 = col_in_690;
assign u_ca_in_691 = col_in_691;
assign u_ca_in_692 = col_in_692;
assign u_ca_in_693 = col_in_693;
assign u_ca_in_694 = col_in_694;
assign u_ca_in_695 = col_in_695;
assign u_ca_in_696 = col_in_696;
assign u_ca_in_697 = col_in_697;
assign u_ca_in_698 = col_in_698;
assign u_ca_in_699 = col_in_699;
assign u_ca_in_700 = col_in_700;
assign u_ca_in_701 = col_in_701;
assign u_ca_in_702 = col_in_702;
assign u_ca_in_703 = col_in_703;
assign u_ca_in_704 = col_in_704;
assign u_ca_in_705 = col_in_705;
assign u_ca_in_706 = col_in_706;
assign u_ca_in_707 = col_in_707;
assign u_ca_in_708 = col_in_708;
assign u_ca_in_709 = col_in_709;
assign u_ca_in_710 = col_in_710;
assign u_ca_in_711 = col_in_711;
assign u_ca_in_712 = col_in_712;
assign u_ca_in_713 = col_in_713;
assign u_ca_in_714 = col_in_714;
assign u_ca_in_715 = col_in_715;
assign u_ca_in_716 = col_in_716;
assign u_ca_in_717 = col_in_717;
assign u_ca_in_718 = col_in_718;
assign u_ca_in_719 = col_in_719;
assign u_ca_in_720 = col_in_720;
assign u_ca_in_721 = col_in_721;
assign u_ca_in_722 = col_in_722;
assign u_ca_in_723 = col_in_723;
assign u_ca_in_724 = col_in_724;
assign u_ca_in_725 = col_in_725;
assign u_ca_in_726 = col_in_726;
assign u_ca_in_727 = col_in_727;
assign u_ca_in_728 = col_in_728;
assign u_ca_in_729 = col_in_729;
assign u_ca_in_730 = col_in_730;
assign u_ca_in_731 = col_in_731;
assign u_ca_in_732 = col_in_732;
assign u_ca_in_733 = col_in_733;
assign u_ca_in_734 = col_in_734;
assign u_ca_in_735 = col_in_735;
assign u_ca_in_736 = col_in_736;
assign u_ca_in_737 = col_in_737;
assign u_ca_in_738 = col_in_738;
assign u_ca_in_739 = col_in_739;
assign u_ca_in_740 = col_in_740;
assign u_ca_in_741 = col_in_741;
assign u_ca_in_742 = col_in_742;
assign u_ca_in_743 = col_in_743;
assign u_ca_in_744 = col_in_744;
assign u_ca_in_745 = col_in_745;
assign u_ca_in_746 = col_in_746;
assign u_ca_in_747 = col_in_747;
assign u_ca_in_748 = col_in_748;
assign u_ca_in_749 = col_in_749;
assign u_ca_in_750 = col_in_750;
assign u_ca_in_751 = col_in_751;
assign u_ca_in_752 = col_in_752;
assign u_ca_in_753 = col_in_753;
assign u_ca_in_754 = col_in_754;
assign u_ca_in_755 = col_in_755;
assign u_ca_in_756 = col_in_756;
assign u_ca_in_757 = col_in_757;
assign u_ca_in_758 = col_in_758;
assign u_ca_in_759 = col_in_759;
assign u_ca_in_760 = col_in_760;
assign u_ca_in_761 = col_in_761;
assign u_ca_in_762 = col_in_762;
assign u_ca_in_763 = col_in_763;
assign u_ca_in_764 = col_in_764;
assign u_ca_in_765 = col_in_765;
assign u_ca_in_766 = col_in_766;
assign u_ca_in_767 = col_in_767;
assign u_ca_in_768 = col_in_768;
assign u_ca_in_769 = col_in_769;
assign u_ca_in_770 = col_in_770;
assign u_ca_in_771 = col_in_771;
assign u_ca_in_772 = col_in_772;
assign u_ca_in_773 = col_in_773;
assign u_ca_in_774 = col_in_774;
assign u_ca_in_775 = col_in_775;
assign u_ca_in_776 = col_in_776;
assign u_ca_in_777 = col_in_777;
assign u_ca_in_778 = col_in_778;
assign u_ca_in_779 = col_in_779;
assign u_ca_in_780 = col_in_780;
assign u_ca_in_781 = col_in_781;
assign u_ca_in_782 = col_in_782;
assign u_ca_in_783 = col_in_783;
assign u_ca_in_784 = col_in_784;
assign u_ca_in_785 = col_in_785;
assign u_ca_in_786 = col_in_786;
assign u_ca_in_787 = col_in_787;
assign u_ca_in_788 = col_in_788;
assign u_ca_in_789 = col_in_789;
assign u_ca_in_790 = col_in_790;
assign u_ca_in_791 = col_in_791;
assign u_ca_in_792 = col_in_792;
assign u_ca_in_793 = col_in_793;
assign u_ca_in_794 = col_in_794;
assign u_ca_in_795 = col_in_795;
assign u_ca_in_796 = col_in_796;
assign u_ca_in_797 = col_in_797;
assign u_ca_in_798 = col_in_798;
assign u_ca_in_799 = col_in_799;
assign u_ca_in_800 = col_in_800;
assign u_ca_in_801 = col_in_801;
assign u_ca_in_802 = col_in_802;
assign u_ca_in_803 = col_in_803;
assign u_ca_in_804 = col_in_804;
assign u_ca_in_805 = col_in_805;
assign u_ca_in_806 = col_in_806;
assign u_ca_in_807 = col_in_807;
assign u_ca_in_808 = col_in_808;
assign u_ca_in_809 = col_in_809;
assign u_ca_in_810 = col_in_810;
assign u_ca_in_811 = col_in_811;
assign u_ca_in_812 = col_in_812;
assign u_ca_in_813 = col_in_813;
assign u_ca_in_814 = col_in_814;
assign u_ca_in_815 = col_in_815;
assign u_ca_in_816 = col_in_816;
assign u_ca_in_817 = col_in_817;
assign u_ca_in_818 = col_in_818;
assign u_ca_in_819 = col_in_819;
assign u_ca_in_820 = col_in_820;
assign u_ca_in_821 = col_in_821;
assign u_ca_in_822 = col_in_822;
assign u_ca_in_823 = col_in_823;
assign u_ca_in_824 = col_in_824;
assign u_ca_in_825 = col_in_825;
assign u_ca_in_826 = col_in_826;
assign u_ca_in_827 = col_in_827;
assign u_ca_in_828 = col_in_828;
assign u_ca_in_829 = col_in_829;
assign u_ca_in_830 = col_in_830;
assign u_ca_in_831 = col_in_831;
assign u_ca_in_832 = col_in_832;
assign u_ca_in_833 = col_in_833;
assign u_ca_in_834 = col_in_834;
assign u_ca_in_835 = col_in_835;
assign u_ca_in_836 = col_in_836;
assign u_ca_in_837 = col_in_837;
assign u_ca_in_838 = col_in_838;
assign u_ca_in_839 = col_in_839;
assign u_ca_in_840 = col_in_840;
assign u_ca_in_841 = col_in_841;
assign u_ca_in_842 = col_in_842;
assign u_ca_in_843 = col_in_843;
assign u_ca_in_844 = col_in_844;
assign u_ca_in_845 = col_in_845;
assign u_ca_in_846 = col_in_846;
assign u_ca_in_847 = col_in_847;
assign u_ca_in_848 = col_in_848;
assign u_ca_in_849 = col_in_849;
assign u_ca_in_850 = col_in_850;
assign u_ca_in_851 = col_in_851;
assign u_ca_in_852 = col_in_852;
assign u_ca_in_853 = col_in_853;
assign u_ca_in_854 = col_in_854;
assign u_ca_in_855 = col_in_855;
assign u_ca_in_856 = col_in_856;
assign u_ca_in_857 = col_in_857;
assign u_ca_in_858 = col_in_858;
assign u_ca_in_859 = col_in_859;
assign u_ca_in_860 = col_in_860;
assign u_ca_in_861 = col_in_861;
assign u_ca_in_862 = col_in_862;
assign u_ca_in_863 = col_in_863;
assign u_ca_in_864 = col_in_864;
assign u_ca_in_865 = col_in_865;
assign u_ca_in_866 = col_in_866;
assign u_ca_in_867 = col_in_867;
assign u_ca_in_868 = col_in_868;
assign u_ca_in_869 = col_in_869;
assign u_ca_in_870 = col_in_870;
assign u_ca_in_871 = col_in_871;
assign u_ca_in_872 = col_in_872;
assign u_ca_in_873 = col_in_873;
assign u_ca_in_874 = col_in_874;
assign u_ca_in_875 = col_in_875;
assign u_ca_in_876 = col_in_876;
assign u_ca_in_877 = col_in_877;
assign u_ca_in_878 = col_in_878;
assign u_ca_in_879 = col_in_879;
assign u_ca_in_880 = col_in_880;
assign u_ca_in_881 = col_in_881;
assign u_ca_in_882 = col_in_882;
assign u_ca_in_883 = col_in_883;
assign u_ca_in_884 = col_in_884;
assign u_ca_in_885 = col_in_885;
assign u_ca_in_886 = col_in_886;
assign u_ca_in_887 = col_in_887;
assign u_ca_in_888 = col_in_888;
assign u_ca_in_889 = col_in_889;
assign u_ca_in_890 = col_in_890;
assign u_ca_in_891 = col_in_891;
assign u_ca_in_892 = col_in_892;
assign u_ca_in_893 = col_in_893;
assign u_ca_in_894 = col_in_894;
assign u_ca_in_895 = col_in_895;
assign u_ca_in_896 = col_in_896;
assign u_ca_in_897 = col_in_897;
assign u_ca_in_898 = col_in_898;
assign u_ca_in_899 = col_in_899;
assign u_ca_in_900 = col_in_900;
assign u_ca_in_901 = col_in_901;
assign u_ca_in_902 = col_in_902;
assign u_ca_in_903 = col_in_903;
assign u_ca_in_904 = col_in_904;
assign u_ca_in_905 = col_in_905;
assign u_ca_in_906 = col_in_906;
assign u_ca_in_907 = col_in_907;
assign u_ca_in_908 = col_in_908;
assign u_ca_in_909 = col_in_909;
assign u_ca_in_910 = col_in_910;
assign u_ca_in_911 = col_in_911;
assign u_ca_in_912 = col_in_912;
assign u_ca_in_913 = col_in_913;
assign u_ca_in_914 = col_in_914;
assign u_ca_in_915 = col_in_915;
assign u_ca_in_916 = col_in_916;
assign u_ca_in_917 = col_in_917;
assign u_ca_in_918 = col_in_918;
assign u_ca_in_919 = col_in_919;
assign u_ca_in_920 = col_in_920;
assign u_ca_in_921 = col_in_921;
assign u_ca_in_922 = col_in_922;
assign u_ca_in_923 = col_in_923;
assign u_ca_in_924 = col_in_924;
assign u_ca_in_925 = col_in_925;
assign u_ca_in_926 = col_in_926;
assign u_ca_in_927 = col_in_927;
assign u_ca_in_928 = col_in_928;
assign u_ca_in_929 = col_in_929;
assign u_ca_in_930 = col_in_930;
assign u_ca_in_931 = col_in_931;
assign u_ca_in_932 = col_in_932;
assign u_ca_in_933 = col_in_933;
assign u_ca_in_934 = col_in_934;
assign u_ca_in_935 = col_in_935;
assign u_ca_in_936 = col_in_936;
assign u_ca_in_937 = col_in_937;
assign u_ca_in_938 = col_in_938;
assign u_ca_in_939 = col_in_939;
assign u_ca_in_940 = col_in_940;
assign u_ca_in_941 = col_in_941;
assign u_ca_in_942 = col_in_942;
assign u_ca_in_943 = col_in_943;
assign u_ca_in_944 = col_in_944;
assign u_ca_in_945 = col_in_945;
assign u_ca_in_946 = col_in_946;
assign u_ca_in_947 = col_in_947;
assign u_ca_in_948 = col_in_948;
assign u_ca_in_949 = col_in_949;
assign u_ca_in_950 = col_in_950;
assign u_ca_in_951 = col_in_951;
assign u_ca_in_952 = col_in_952;
assign u_ca_in_953 = col_in_953;
assign u_ca_in_954 = col_in_954;
assign u_ca_in_955 = col_in_955;
assign u_ca_in_956 = col_in_956;
assign u_ca_in_957 = col_in_957;
assign u_ca_in_958 = col_in_958;
assign u_ca_in_959 = col_in_959;
assign u_ca_in_960 = col_in_960;
assign u_ca_in_961 = col_in_961;
assign u_ca_in_962 = col_in_962;
assign u_ca_in_963 = col_in_963;
assign u_ca_in_964 = col_in_964;
assign u_ca_in_965 = col_in_965;
assign u_ca_in_966 = col_in_966;
assign u_ca_in_967 = col_in_967;
assign u_ca_in_968 = col_in_968;
assign u_ca_in_969 = col_in_969;
assign u_ca_in_970 = col_in_970;
assign u_ca_in_971 = col_in_971;
assign u_ca_in_972 = col_in_972;
assign u_ca_in_973 = col_in_973;
assign u_ca_in_974 = col_in_974;
assign u_ca_in_975 = col_in_975;
assign u_ca_in_976 = col_in_976;
assign u_ca_in_977 = col_in_977;
assign u_ca_in_978 = col_in_978;
assign u_ca_in_979 = col_in_979;
assign u_ca_in_980 = col_in_980;
assign u_ca_in_981 = col_in_981;
assign u_ca_in_982 = col_in_982;
assign u_ca_in_983 = col_in_983;
assign u_ca_in_984 = col_in_984;
assign u_ca_in_985 = col_in_985;
assign u_ca_in_986 = col_in_986;
assign u_ca_in_987 = col_in_987;
assign u_ca_in_988 = col_in_988;
assign u_ca_in_989 = col_in_989;
assign u_ca_in_990 = col_in_990;
assign u_ca_in_991 = col_in_991;
assign u_ca_in_992 = col_in_992;
assign u_ca_in_993 = col_in_993;
assign u_ca_in_994 = col_in_994;
assign u_ca_in_995 = col_in_995;
assign u_ca_in_996 = col_in_996;
assign u_ca_in_997 = col_in_997;
assign u_ca_in_998 = col_in_998;
assign u_ca_in_999 = col_in_999;
assign u_ca_in_1000 = col_in_1000;
assign u_ca_in_1001 = col_in_1001;
assign u_ca_in_1002 = col_in_1002;
assign u_ca_in_1003 = col_in_1003;
assign u_ca_in_1004 = col_in_1004;
assign u_ca_in_1005 = col_in_1005;
assign u_ca_in_1006 = col_in_1006;
assign u_ca_in_1007 = col_in_1007;
assign u_ca_in_1008 = col_in_1008;
assign u_ca_in_1009 = col_in_1009;
assign u_ca_in_1010 = col_in_1010;
assign u_ca_in_1011 = col_in_1011;
assign u_ca_in_1012 = col_in_1012;
assign u_ca_in_1013 = col_in_1013;
assign u_ca_in_1014 = col_in_1014;
assign u_ca_in_1015 = col_in_1015;
assign u_ca_in_1016 = col_in_1016;
assign u_ca_in_1017 = col_in_1017;
assign u_ca_in_1018 = col_in_1018;
assign u_ca_in_1019 = col_in_1019;
assign u_ca_in_1020 = col_in_1020;
assign u_ca_in_1021 = col_in_1021;
assign u_ca_in_1022 = col_in_1022;
assign u_ca_in_1023 = col_in_1023;

//---------------------------------------------------------



//--compressor_array---------------------------------------
compressor_3_2 u_ca_3_2_0(.d_in(u_ca_in_0), .d_out(u_ca_out_0));
compressor_3_2 u_ca_3_2_1(.d_in(u_ca_in_1), .d_out(u_ca_out_1));
compressor_3_2 u_ca_3_2_2(.d_in(u_ca_in_2), .d_out(u_ca_out_2));
compressor_3_2 u_ca_3_2_3(.d_in(u_ca_in_3), .d_out(u_ca_out_3));
compressor_3_2 u_ca_3_2_4(.d_in(u_ca_in_4), .d_out(u_ca_out_4));
compressor_3_2 u_ca_3_2_5(.d_in(u_ca_in_5), .d_out(u_ca_out_5));
compressor_3_2 u_ca_3_2_6(.d_in(u_ca_in_6), .d_out(u_ca_out_6));
compressor_3_2 u_ca_3_2_7(.d_in(u_ca_in_7), .d_out(u_ca_out_7));
compressor_3_2 u_ca_3_2_8(.d_in(u_ca_in_8), .d_out(u_ca_out_8));
compressor_3_2 u_ca_3_2_9(.d_in(u_ca_in_9), .d_out(u_ca_out_9));
compressor_3_2 u_ca_3_2_10(.d_in(u_ca_in_10), .d_out(u_ca_out_10));
compressor_3_2 u_ca_3_2_11(.d_in(u_ca_in_11), .d_out(u_ca_out_11));
compressor_3_2 u_ca_3_2_12(.d_in(u_ca_in_12), .d_out(u_ca_out_12));
compressor_3_2 u_ca_3_2_13(.d_in(u_ca_in_13), .d_out(u_ca_out_13));
compressor_3_2 u_ca_3_2_14(.d_in(u_ca_in_14), .d_out(u_ca_out_14));
compressor_3_2 u_ca_3_2_15(.d_in(u_ca_in_15), .d_out(u_ca_out_15));
compressor_3_2 u_ca_3_2_16(.d_in(u_ca_in_16), .d_out(u_ca_out_16));
compressor_3_2 u_ca_3_2_17(.d_in(u_ca_in_17), .d_out(u_ca_out_17));
compressor_3_2 u_ca_3_2_18(.d_in(u_ca_in_18), .d_out(u_ca_out_18));
compressor_3_2 u_ca_3_2_19(.d_in(u_ca_in_19), .d_out(u_ca_out_19));
compressor_3_2 u_ca_3_2_20(.d_in(u_ca_in_20), .d_out(u_ca_out_20));
compressor_3_2 u_ca_3_2_21(.d_in(u_ca_in_21), .d_out(u_ca_out_21));
compressor_3_2 u_ca_3_2_22(.d_in(u_ca_in_22), .d_out(u_ca_out_22));
compressor_3_2 u_ca_3_2_23(.d_in(u_ca_in_23), .d_out(u_ca_out_23));
compressor_3_2 u_ca_3_2_24(.d_in(u_ca_in_24), .d_out(u_ca_out_24));
compressor_3_2 u_ca_3_2_25(.d_in(u_ca_in_25), .d_out(u_ca_out_25));
compressor_3_2 u_ca_3_2_26(.d_in(u_ca_in_26), .d_out(u_ca_out_26));
compressor_3_2 u_ca_3_2_27(.d_in(u_ca_in_27), .d_out(u_ca_out_27));
compressor_3_2 u_ca_3_2_28(.d_in(u_ca_in_28), .d_out(u_ca_out_28));
compressor_3_2 u_ca_3_2_29(.d_in(u_ca_in_29), .d_out(u_ca_out_29));
compressor_3_2 u_ca_3_2_30(.d_in(u_ca_in_30), .d_out(u_ca_out_30));
compressor_3_2 u_ca_3_2_31(.d_in(u_ca_in_31), .d_out(u_ca_out_31));
compressor_3_2 u_ca_3_2_32(.d_in(u_ca_in_32), .d_out(u_ca_out_32));
compressor_3_2 u_ca_3_2_33(.d_in(u_ca_in_33), .d_out(u_ca_out_33));
compressor_3_2 u_ca_3_2_34(.d_in(u_ca_in_34), .d_out(u_ca_out_34));
compressor_3_2 u_ca_3_2_35(.d_in(u_ca_in_35), .d_out(u_ca_out_35));
compressor_3_2 u_ca_3_2_36(.d_in(u_ca_in_36), .d_out(u_ca_out_36));
compressor_3_2 u_ca_3_2_37(.d_in(u_ca_in_37), .d_out(u_ca_out_37));
compressor_3_2 u_ca_3_2_38(.d_in(u_ca_in_38), .d_out(u_ca_out_38));
compressor_3_2 u_ca_3_2_39(.d_in(u_ca_in_39), .d_out(u_ca_out_39));
compressor_3_2 u_ca_3_2_40(.d_in(u_ca_in_40), .d_out(u_ca_out_40));
compressor_3_2 u_ca_3_2_41(.d_in(u_ca_in_41), .d_out(u_ca_out_41));
compressor_3_2 u_ca_3_2_42(.d_in(u_ca_in_42), .d_out(u_ca_out_42));
compressor_3_2 u_ca_3_2_43(.d_in(u_ca_in_43), .d_out(u_ca_out_43));
compressor_3_2 u_ca_3_2_44(.d_in(u_ca_in_44), .d_out(u_ca_out_44));
compressor_3_2 u_ca_3_2_45(.d_in(u_ca_in_45), .d_out(u_ca_out_45));
compressor_3_2 u_ca_3_2_46(.d_in(u_ca_in_46), .d_out(u_ca_out_46));
compressor_3_2 u_ca_3_2_47(.d_in(u_ca_in_47), .d_out(u_ca_out_47));
compressor_3_2 u_ca_3_2_48(.d_in(u_ca_in_48), .d_out(u_ca_out_48));
compressor_3_2 u_ca_3_2_49(.d_in(u_ca_in_49), .d_out(u_ca_out_49));
compressor_3_2 u_ca_3_2_50(.d_in(u_ca_in_50), .d_out(u_ca_out_50));
compressor_3_2 u_ca_3_2_51(.d_in(u_ca_in_51), .d_out(u_ca_out_51));
compressor_3_2 u_ca_3_2_52(.d_in(u_ca_in_52), .d_out(u_ca_out_52));
compressor_3_2 u_ca_3_2_53(.d_in(u_ca_in_53), .d_out(u_ca_out_53));
compressor_3_2 u_ca_3_2_54(.d_in(u_ca_in_54), .d_out(u_ca_out_54));
compressor_3_2 u_ca_3_2_55(.d_in(u_ca_in_55), .d_out(u_ca_out_55));
compressor_3_2 u_ca_3_2_56(.d_in(u_ca_in_56), .d_out(u_ca_out_56));
compressor_3_2 u_ca_3_2_57(.d_in(u_ca_in_57), .d_out(u_ca_out_57));
compressor_3_2 u_ca_3_2_58(.d_in(u_ca_in_58), .d_out(u_ca_out_58));
compressor_3_2 u_ca_3_2_59(.d_in(u_ca_in_59), .d_out(u_ca_out_59));
compressor_3_2 u_ca_3_2_60(.d_in(u_ca_in_60), .d_out(u_ca_out_60));
compressor_3_2 u_ca_3_2_61(.d_in(u_ca_in_61), .d_out(u_ca_out_61));
compressor_3_2 u_ca_3_2_62(.d_in(u_ca_in_62), .d_out(u_ca_out_62));
compressor_3_2 u_ca_3_2_63(.d_in(u_ca_in_63), .d_out(u_ca_out_63));
compressor_3_2 u_ca_3_2_64(.d_in(u_ca_in_64), .d_out(u_ca_out_64));
compressor_3_2 u_ca_3_2_65(.d_in(u_ca_in_65), .d_out(u_ca_out_65));
compressor_3_2 u_ca_3_2_66(.d_in(u_ca_in_66), .d_out(u_ca_out_66));
compressor_3_2 u_ca_3_2_67(.d_in(u_ca_in_67), .d_out(u_ca_out_67));
compressor_3_2 u_ca_3_2_68(.d_in(u_ca_in_68), .d_out(u_ca_out_68));
compressor_3_2 u_ca_3_2_69(.d_in(u_ca_in_69), .d_out(u_ca_out_69));
compressor_3_2 u_ca_3_2_70(.d_in(u_ca_in_70), .d_out(u_ca_out_70));
compressor_3_2 u_ca_3_2_71(.d_in(u_ca_in_71), .d_out(u_ca_out_71));
compressor_3_2 u_ca_3_2_72(.d_in(u_ca_in_72), .d_out(u_ca_out_72));
compressor_3_2 u_ca_3_2_73(.d_in(u_ca_in_73), .d_out(u_ca_out_73));
compressor_3_2 u_ca_3_2_74(.d_in(u_ca_in_74), .d_out(u_ca_out_74));
compressor_3_2 u_ca_3_2_75(.d_in(u_ca_in_75), .d_out(u_ca_out_75));
compressor_3_2 u_ca_3_2_76(.d_in(u_ca_in_76), .d_out(u_ca_out_76));
compressor_3_2 u_ca_3_2_77(.d_in(u_ca_in_77), .d_out(u_ca_out_77));
compressor_3_2 u_ca_3_2_78(.d_in(u_ca_in_78), .d_out(u_ca_out_78));
compressor_3_2 u_ca_3_2_79(.d_in(u_ca_in_79), .d_out(u_ca_out_79));
compressor_3_2 u_ca_3_2_80(.d_in(u_ca_in_80), .d_out(u_ca_out_80));
compressor_3_2 u_ca_3_2_81(.d_in(u_ca_in_81), .d_out(u_ca_out_81));
compressor_3_2 u_ca_3_2_82(.d_in(u_ca_in_82), .d_out(u_ca_out_82));
compressor_3_2 u_ca_3_2_83(.d_in(u_ca_in_83), .d_out(u_ca_out_83));
compressor_3_2 u_ca_3_2_84(.d_in(u_ca_in_84), .d_out(u_ca_out_84));
compressor_3_2 u_ca_3_2_85(.d_in(u_ca_in_85), .d_out(u_ca_out_85));
compressor_3_2 u_ca_3_2_86(.d_in(u_ca_in_86), .d_out(u_ca_out_86));
compressor_3_2 u_ca_3_2_87(.d_in(u_ca_in_87), .d_out(u_ca_out_87));
compressor_3_2 u_ca_3_2_88(.d_in(u_ca_in_88), .d_out(u_ca_out_88));
compressor_3_2 u_ca_3_2_89(.d_in(u_ca_in_89), .d_out(u_ca_out_89));
compressor_3_2 u_ca_3_2_90(.d_in(u_ca_in_90), .d_out(u_ca_out_90));
compressor_3_2 u_ca_3_2_91(.d_in(u_ca_in_91), .d_out(u_ca_out_91));
compressor_3_2 u_ca_3_2_92(.d_in(u_ca_in_92), .d_out(u_ca_out_92));
compressor_3_2 u_ca_3_2_93(.d_in(u_ca_in_93), .d_out(u_ca_out_93));
compressor_3_2 u_ca_3_2_94(.d_in(u_ca_in_94), .d_out(u_ca_out_94));
compressor_3_2 u_ca_3_2_95(.d_in(u_ca_in_95), .d_out(u_ca_out_95));
compressor_3_2 u_ca_3_2_96(.d_in(u_ca_in_96), .d_out(u_ca_out_96));
compressor_3_2 u_ca_3_2_97(.d_in(u_ca_in_97), .d_out(u_ca_out_97));
compressor_3_2 u_ca_3_2_98(.d_in(u_ca_in_98), .d_out(u_ca_out_98));
compressor_3_2 u_ca_3_2_99(.d_in(u_ca_in_99), .d_out(u_ca_out_99));
compressor_3_2 u_ca_3_2_100(.d_in(u_ca_in_100), .d_out(u_ca_out_100));
compressor_3_2 u_ca_3_2_101(.d_in(u_ca_in_101), .d_out(u_ca_out_101));
compressor_3_2 u_ca_3_2_102(.d_in(u_ca_in_102), .d_out(u_ca_out_102));
compressor_3_2 u_ca_3_2_103(.d_in(u_ca_in_103), .d_out(u_ca_out_103));
compressor_3_2 u_ca_3_2_104(.d_in(u_ca_in_104), .d_out(u_ca_out_104));
compressor_3_2 u_ca_3_2_105(.d_in(u_ca_in_105), .d_out(u_ca_out_105));
compressor_3_2 u_ca_3_2_106(.d_in(u_ca_in_106), .d_out(u_ca_out_106));
compressor_3_2 u_ca_3_2_107(.d_in(u_ca_in_107), .d_out(u_ca_out_107));
compressor_3_2 u_ca_3_2_108(.d_in(u_ca_in_108), .d_out(u_ca_out_108));
compressor_3_2 u_ca_3_2_109(.d_in(u_ca_in_109), .d_out(u_ca_out_109));
compressor_3_2 u_ca_3_2_110(.d_in(u_ca_in_110), .d_out(u_ca_out_110));
compressor_3_2 u_ca_3_2_111(.d_in(u_ca_in_111), .d_out(u_ca_out_111));
compressor_3_2 u_ca_3_2_112(.d_in(u_ca_in_112), .d_out(u_ca_out_112));
compressor_3_2 u_ca_3_2_113(.d_in(u_ca_in_113), .d_out(u_ca_out_113));
compressor_3_2 u_ca_3_2_114(.d_in(u_ca_in_114), .d_out(u_ca_out_114));
compressor_3_2 u_ca_3_2_115(.d_in(u_ca_in_115), .d_out(u_ca_out_115));
compressor_3_2 u_ca_3_2_116(.d_in(u_ca_in_116), .d_out(u_ca_out_116));
compressor_3_2 u_ca_3_2_117(.d_in(u_ca_in_117), .d_out(u_ca_out_117));
compressor_3_2 u_ca_3_2_118(.d_in(u_ca_in_118), .d_out(u_ca_out_118));
compressor_3_2 u_ca_3_2_119(.d_in(u_ca_in_119), .d_out(u_ca_out_119));
compressor_3_2 u_ca_3_2_120(.d_in(u_ca_in_120), .d_out(u_ca_out_120));
compressor_3_2 u_ca_3_2_121(.d_in(u_ca_in_121), .d_out(u_ca_out_121));
compressor_3_2 u_ca_3_2_122(.d_in(u_ca_in_122), .d_out(u_ca_out_122));
compressor_3_2 u_ca_3_2_123(.d_in(u_ca_in_123), .d_out(u_ca_out_123));
compressor_3_2 u_ca_3_2_124(.d_in(u_ca_in_124), .d_out(u_ca_out_124));
compressor_3_2 u_ca_3_2_125(.d_in(u_ca_in_125), .d_out(u_ca_out_125));
compressor_3_2 u_ca_3_2_126(.d_in(u_ca_in_126), .d_out(u_ca_out_126));
compressor_3_2 u_ca_3_2_127(.d_in(u_ca_in_127), .d_out(u_ca_out_127));
compressor_3_2 u_ca_3_2_128(.d_in(u_ca_in_128), .d_out(u_ca_out_128));
compressor_3_2 u_ca_3_2_129(.d_in(u_ca_in_129), .d_out(u_ca_out_129));
compressor_3_2 u_ca_3_2_130(.d_in(u_ca_in_130), .d_out(u_ca_out_130));
compressor_3_2 u_ca_3_2_131(.d_in(u_ca_in_131), .d_out(u_ca_out_131));
compressor_3_2 u_ca_3_2_132(.d_in(u_ca_in_132), .d_out(u_ca_out_132));
compressor_3_2 u_ca_3_2_133(.d_in(u_ca_in_133), .d_out(u_ca_out_133));
compressor_3_2 u_ca_3_2_134(.d_in(u_ca_in_134), .d_out(u_ca_out_134));
compressor_3_2 u_ca_3_2_135(.d_in(u_ca_in_135), .d_out(u_ca_out_135));
compressor_3_2 u_ca_3_2_136(.d_in(u_ca_in_136), .d_out(u_ca_out_136));
compressor_3_2 u_ca_3_2_137(.d_in(u_ca_in_137), .d_out(u_ca_out_137));
compressor_3_2 u_ca_3_2_138(.d_in(u_ca_in_138), .d_out(u_ca_out_138));
compressor_3_2 u_ca_3_2_139(.d_in(u_ca_in_139), .d_out(u_ca_out_139));
compressor_3_2 u_ca_3_2_140(.d_in(u_ca_in_140), .d_out(u_ca_out_140));
compressor_3_2 u_ca_3_2_141(.d_in(u_ca_in_141), .d_out(u_ca_out_141));
compressor_3_2 u_ca_3_2_142(.d_in(u_ca_in_142), .d_out(u_ca_out_142));
compressor_3_2 u_ca_3_2_143(.d_in(u_ca_in_143), .d_out(u_ca_out_143));
compressor_3_2 u_ca_3_2_144(.d_in(u_ca_in_144), .d_out(u_ca_out_144));
compressor_3_2 u_ca_3_2_145(.d_in(u_ca_in_145), .d_out(u_ca_out_145));
compressor_3_2 u_ca_3_2_146(.d_in(u_ca_in_146), .d_out(u_ca_out_146));
compressor_3_2 u_ca_3_2_147(.d_in(u_ca_in_147), .d_out(u_ca_out_147));
compressor_3_2 u_ca_3_2_148(.d_in(u_ca_in_148), .d_out(u_ca_out_148));
compressor_3_2 u_ca_3_2_149(.d_in(u_ca_in_149), .d_out(u_ca_out_149));
compressor_3_2 u_ca_3_2_150(.d_in(u_ca_in_150), .d_out(u_ca_out_150));
compressor_3_2 u_ca_3_2_151(.d_in(u_ca_in_151), .d_out(u_ca_out_151));
compressor_3_2 u_ca_3_2_152(.d_in(u_ca_in_152), .d_out(u_ca_out_152));
compressor_3_2 u_ca_3_2_153(.d_in(u_ca_in_153), .d_out(u_ca_out_153));
compressor_3_2 u_ca_3_2_154(.d_in(u_ca_in_154), .d_out(u_ca_out_154));
compressor_3_2 u_ca_3_2_155(.d_in(u_ca_in_155), .d_out(u_ca_out_155));
compressor_3_2 u_ca_3_2_156(.d_in(u_ca_in_156), .d_out(u_ca_out_156));
compressor_3_2 u_ca_3_2_157(.d_in(u_ca_in_157), .d_out(u_ca_out_157));
compressor_3_2 u_ca_3_2_158(.d_in(u_ca_in_158), .d_out(u_ca_out_158));
compressor_3_2 u_ca_3_2_159(.d_in(u_ca_in_159), .d_out(u_ca_out_159));
compressor_3_2 u_ca_3_2_160(.d_in(u_ca_in_160), .d_out(u_ca_out_160));
compressor_3_2 u_ca_3_2_161(.d_in(u_ca_in_161), .d_out(u_ca_out_161));
compressor_3_2 u_ca_3_2_162(.d_in(u_ca_in_162), .d_out(u_ca_out_162));
compressor_3_2 u_ca_3_2_163(.d_in(u_ca_in_163), .d_out(u_ca_out_163));
compressor_3_2 u_ca_3_2_164(.d_in(u_ca_in_164), .d_out(u_ca_out_164));
compressor_3_2 u_ca_3_2_165(.d_in(u_ca_in_165), .d_out(u_ca_out_165));
compressor_3_2 u_ca_3_2_166(.d_in(u_ca_in_166), .d_out(u_ca_out_166));
compressor_3_2 u_ca_3_2_167(.d_in(u_ca_in_167), .d_out(u_ca_out_167));
compressor_3_2 u_ca_3_2_168(.d_in(u_ca_in_168), .d_out(u_ca_out_168));
compressor_3_2 u_ca_3_2_169(.d_in(u_ca_in_169), .d_out(u_ca_out_169));
compressor_3_2 u_ca_3_2_170(.d_in(u_ca_in_170), .d_out(u_ca_out_170));
compressor_3_2 u_ca_3_2_171(.d_in(u_ca_in_171), .d_out(u_ca_out_171));
compressor_3_2 u_ca_3_2_172(.d_in(u_ca_in_172), .d_out(u_ca_out_172));
compressor_3_2 u_ca_3_2_173(.d_in(u_ca_in_173), .d_out(u_ca_out_173));
compressor_3_2 u_ca_3_2_174(.d_in(u_ca_in_174), .d_out(u_ca_out_174));
compressor_3_2 u_ca_3_2_175(.d_in(u_ca_in_175), .d_out(u_ca_out_175));
compressor_3_2 u_ca_3_2_176(.d_in(u_ca_in_176), .d_out(u_ca_out_176));
compressor_3_2 u_ca_3_2_177(.d_in(u_ca_in_177), .d_out(u_ca_out_177));
compressor_3_2 u_ca_3_2_178(.d_in(u_ca_in_178), .d_out(u_ca_out_178));
compressor_3_2 u_ca_3_2_179(.d_in(u_ca_in_179), .d_out(u_ca_out_179));
compressor_3_2 u_ca_3_2_180(.d_in(u_ca_in_180), .d_out(u_ca_out_180));
compressor_3_2 u_ca_3_2_181(.d_in(u_ca_in_181), .d_out(u_ca_out_181));
compressor_3_2 u_ca_3_2_182(.d_in(u_ca_in_182), .d_out(u_ca_out_182));
compressor_3_2 u_ca_3_2_183(.d_in(u_ca_in_183), .d_out(u_ca_out_183));
compressor_3_2 u_ca_3_2_184(.d_in(u_ca_in_184), .d_out(u_ca_out_184));
compressor_3_2 u_ca_3_2_185(.d_in(u_ca_in_185), .d_out(u_ca_out_185));
compressor_3_2 u_ca_3_2_186(.d_in(u_ca_in_186), .d_out(u_ca_out_186));
compressor_3_2 u_ca_3_2_187(.d_in(u_ca_in_187), .d_out(u_ca_out_187));
compressor_3_2 u_ca_3_2_188(.d_in(u_ca_in_188), .d_out(u_ca_out_188));
compressor_3_2 u_ca_3_2_189(.d_in(u_ca_in_189), .d_out(u_ca_out_189));
compressor_3_2 u_ca_3_2_190(.d_in(u_ca_in_190), .d_out(u_ca_out_190));
compressor_3_2 u_ca_3_2_191(.d_in(u_ca_in_191), .d_out(u_ca_out_191));
compressor_3_2 u_ca_3_2_192(.d_in(u_ca_in_192), .d_out(u_ca_out_192));
compressor_3_2 u_ca_3_2_193(.d_in(u_ca_in_193), .d_out(u_ca_out_193));
compressor_3_2 u_ca_3_2_194(.d_in(u_ca_in_194), .d_out(u_ca_out_194));
compressor_3_2 u_ca_3_2_195(.d_in(u_ca_in_195), .d_out(u_ca_out_195));
compressor_3_2 u_ca_3_2_196(.d_in(u_ca_in_196), .d_out(u_ca_out_196));
compressor_3_2 u_ca_3_2_197(.d_in(u_ca_in_197), .d_out(u_ca_out_197));
compressor_3_2 u_ca_3_2_198(.d_in(u_ca_in_198), .d_out(u_ca_out_198));
compressor_3_2 u_ca_3_2_199(.d_in(u_ca_in_199), .d_out(u_ca_out_199));
compressor_3_2 u_ca_3_2_200(.d_in(u_ca_in_200), .d_out(u_ca_out_200));
compressor_3_2 u_ca_3_2_201(.d_in(u_ca_in_201), .d_out(u_ca_out_201));
compressor_3_2 u_ca_3_2_202(.d_in(u_ca_in_202), .d_out(u_ca_out_202));
compressor_3_2 u_ca_3_2_203(.d_in(u_ca_in_203), .d_out(u_ca_out_203));
compressor_3_2 u_ca_3_2_204(.d_in(u_ca_in_204), .d_out(u_ca_out_204));
compressor_3_2 u_ca_3_2_205(.d_in(u_ca_in_205), .d_out(u_ca_out_205));
compressor_3_2 u_ca_3_2_206(.d_in(u_ca_in_206), .d_out(u_ca_out_206));
compressor_3_2 u_ca_3_2_207(.d_in(u_ca_in_207), .d_out(u_ca_out_207));
compressor_3_2 u_ca_3_2_208(.d_in(u_ca_in_208), .d_out(u_ca_out_208));
compressor_3_2 u_ca_3_2_209(.d_in(u_ca_in_209), .d_out(u_ca_out_209));
compressor_3_2 u_ca_3_2_210(.d_in(u_ca_in_210), .d_out(u_ca_out_210));
compressor_3_2 u_ca_3_2_211(.d_in(u_ca_in_211), .d_out(u_ca_out_211));
compressor_3_2 u_ca_3_2_212(.d_in(u_ca_in_212), .d_out(u_ca_out_212));
compressor_3_2 u_ca_3_2_213(.d_in(u_ca_in_213), .d_out(u_ca_out_213));
compressor_3_2 u_ca_3_2_214(.d_in(u_ca_in_214), .d_out(u_ca_out_214));
compressor_3_2 u_ca_3_2_215(.d_in(u_ca_in_215), .d_out(u_ca_out_215));
compressor_3_2 u_ca_3_2_216(.d_in(u_ca_in_216), .d_out(u_ca_out_216));
compressor_3_2 u_ca_3_2_217(.d_in(u_ca_in_217), .d_out(u_ca_out_217));
compressor_3_2 u_ca_3_2_218(.d_in(u_ca_in_218), .d_out(u_ca_out_218));
compressor_3_2 u_ca_3_2_219(.d_in(u_ca_in_219), .d_out(u_ca_out_219));
compressor_3_2 u_ca_3_2_220(.d_in(u_ca_in_220), .d_out(u_ca_out_220));
compressor_3_2 u_ca_3_2_221(.d_in(u_ca_in_221), .d_out(u_ca_out_221));
compressor_3_2 u_ca_3_2_222(.d_in(u_ca_in_222), .d_out(u_ca_out_222));
compressor_3_2 u_ca_3_2_223(.d_in(u_ca_in_223), .d_out(u_ca_out_223));
compressor_3_2 u_ca_3_2_224(.d_in(u_ca_in_224), .d_out(u_ca_out_224));
compressor_3_2 u_ca_3_2_225(.d_in(u_ca_in_225), .d_out(u_ca_out_225));
compressor_3_2 u_ca_3_2_226(.d_in(u_ca_in_226), .d_out(u_ca_out_226));
compressor_3_2 u_ca_3_2_227(.d_in(u_ca_in_227), .d_out(u_ca_out_227));
compressor_3_2 u_ca_3_2_228(.d_in(u_ca_in_228), .d_out(u_ca_out_228));
compressor_3_2 u_ca_3_2_229(.d_in(u_ca_in_229), .d_out(u_ca_out_229));
compressor_3_2 u_ca_3_2_230(.d_in(u_ca_in_230), .d_out(u_ca_out_230));
compressor_3_2 u_ca_3_2_231(.d_in(u_ca_in_231), .d_out(u_ca_out_231));
compressor_3_2 u_ca_3_2_232(.d_in(u_ca_in_232), .d_out(u_ca_out_232));
compressor_3_2 u_ca_3_2_233(.d_in(u_ca_in_233), .d_out(u_ca_out_233));
compressor_3_2 u_ca_3_2_234(.d_in(u_ca_in_234), .d_out(u_ca_out_234));
compressor_3_2 u_ca_3_2_235(.d_in(u_ca_in_235), .d_out(u_ca_out_235));
compressor_3_2 u_ca_3_2_236(.d_in(u_ca_in_236), .d_out(u_ca_out_236));
compressor_3_2 u_ca_3_2_237(.d_in(u_ca_in_237), .d_out(u_ca_out_237));
compressor_3_2 u_ca_3_2_238(.d_in(u_ca_in_238), .d_out(u_ca_out_238));
compressor_3_2 u_ca_3_2_239(.d_in(u_ca_in_239), .d_out(u_ca_out_239));
compressor_3_2 u_ca_3_2_240(.d_in(u_ca_in_240), .d_out(u_ca_out_240));
compressor_3_2 u_ca_3_2_241(.d_in(u_ca_in_241), .d_out(u_ca_out_241));
compressor_3_2 u_ca_3_2_242(.d_in(u_ca_in_242), .d_out(u_ca_out_242));
compressor_3_2 u_ca_3_2_243(.d_in(u_ca_in_243), .d_out(u_ca_out_243));
compressor_3_2 u_ca_3_2_244(.d_in(u_ca_in_244), .d_out(u_ca_out_244));
compressor_3_2 u_ca_3_2_245(.d_in(u_ca_in_245), .d_out(u_ca_out_245));
compressor_3_2 u_ca_3_2_246(.d_in(u_ca_in_246), .d_out(u_ca_out_246));
compressor_3_2 u_ca_3_2_247(.d_in(u_ca_in_247), .d_out(u_ca_out_247));
compressor_3_2 u_ca_3_2_248(.d_in(u_ca_in_248), .d_out(u_ca_out_248));
compressor_3_2 u_ca_3_2_249(.d_in(u_ca_in_249), .d_out(u_ca_out_249));
compressor_3_2 u_ca_3_2_250(.d_in(u_ca_in_250), .d_out(u_ca_out_250));
compressor_3_2 u_ca_3_2_251(.d_in(u_ca_in_251), .d_out(u_ca_out_251));
compressor_3_2 u_ca_3_2_252(.d_in(u_ca_in_252), .d_out(u_ca_out_252));
compressor_3_2 u_ca_3_2_253(.d_in(u_ca_in_253), .d_out(u_ca_out_253));
compressor_3_2 u_ca_3_2_254(.d_in(u_ca_in_254), .d_out(u_ca_out_254));
compressor_3_2 u_ca_3_2_255(.d_in(u_ca_in_255), .d_out(u_ca_out_255));
compressor_3_2 u_ca_3_2_256(.d_in(u_ca_in_256), .d_out(u_ca_out_256));
compressor_3_2 u_ca_3_2_257(.d_in(u_ca_in_257), .d_out(u_ca_out_257));
compressor_3_2 u_ca_3_2_258(.d_in(u_ca_in_258), .d_out(u_ca_out_258));
compressor_3_2 u_ca_3_2_259(.d_in(u_ca_in_259), .d_out(u_ca_out_259));
compressor_3_2 u_ca_3_2_260(.d_in(u_ca_in_260), .d_out(u_ca_out_260));
compressor_3_2 u_ca_3_2_261(.d_in(u_ca_in_261), .d_out(u_ca_out_261));
compressor_3_2 u_ca_3_2_262(.d_in(u_ca_in_262), .d_out(u_ca_out_262));
compressor_3_2 u_ca_3_2_263(.d_in(u_ca_in_263), .d_out(u_ca_out_263));
compressor_3_2 u_ca_3_2_264(.d_in(u_ca_in_264), .d_out(u_ca_out_264));
compressor_3_2 u_ca_3_2_265(.d_in(u_ca_in_265), .d_out(u_ca_out_265));
compressor_3_2 u_ca_3_2_266(.d_in(u_ca_in_266), .d_out(u_ca_out_266));
compressor_3_2 u_ca_3_2_267(.d_in(u_ca_in_267), .d_out(u_ca_out_267));
compressor_3_2 u_ca_3_2_268(.d_in(u_ca_in_268), .d_out(u_ca_out_268));
compressor_3_2 u_ca_3_2_269(.d_in(u_ca_in_269), .d_out(u_ca_out_269));
compressor_3_2 u_ca_3_2_270(.d_in(u_ca_in_270), .d_out(u_ca_out_270));
compressor_3_2 u_ca_3_2_271(.d_in(u_ca_in_271), .d_out(u_ca_out_271));
compressor_3_2 u_ca_3_2_272(.d_in(u_ca_in_272), .d_out(u_ca_out_272));
compressor_3_2 u_ca_3_2_273(.d_in(u_ca_in_273), .d_out(u_ca_out_273));
compressor_3_2 u_ca_3_2_274(.d_in(u_ca_in_274), .d_out(u_ca_out_274));
compressor_3_2 u_ca_3_2_275(.d_in(u_ca_in_275), .d_out(u_ca_out_275));
compressor_3_2 u_ca_3_2_276(.d_in(u_ca_in_276), .d_out(u_ca_out_276));
compressor_3_2 u_ca_3_2_277(.d_in(u_ca_in_277), .d_out(u_ca_out_277));
compressor_3_2 u_ca_3_2_278(.d_in(u_ca_in_278), .d_out(u_ca_out_278));
compressor_3_2 u_ca_3_2_279(.d_in(u_ca_in_279), .d_out(u_ca_out_279));
compressor_3_2 u_ca_3_2_280(.d_in(u_ca_in_280), .d_out(u_ca_out_280));
compressor_3_2 u_ca_3_2_281(.d_in(u_ca_in_281), .d_out(u_ca_out_281));
compressor_3_2 u_ca_3_2_282(.d_in(u_ca_in_282), .d_out(u_ca_out_282));
compressor_3_2 u_ca_3_2_283(.d_in(u_ca_in_283), .d_out(u_ca_out_283));
compressor_3_2 u_ca_3_2_284(.d_in(u_ca_in_284), .d_out(u_ca_out_284));
compressor_3_2 u_ca_3_2_285(.d_in(u_ca_in_285), .d_out(u_ca_out_285));
compressor_3_2 u_ca_3_2_286(.d_in(u_ca_in_286), .d_out(u_ca_out_286));
compressor_3_2 u_ca_3_2_287(.d_in(u_ca_in_287), .d_out(u_ca_out_287));
compressor_3_2 u_ca_3_2_288(.d_in(u_ca_in_288), .d_out(u_ca_out_288));
compressor_3_2 u_ca_3_2_289(.d_in(u_ca_in_289), .d_out(u_ca_out_289));
compressor_3_2 u_ca_3_2_290(.d_in(u_ca_in_290), .d_out(u_ca_out_290));
compressor_3_2 u_ca_3_2_291(.d_in(u_ca_in_291), .d_out(u_ca_out_291));
compressor_3_2 u_ca_3_2_292(.d_in(u_ca_in_292), .d_out(u_ca_out_292));
compressor_3_2 u_ca_3_2_293(.d_in(u_ca_in_293), .d_out(u_ca_out_293));
compressor_3_2 u_ca_3_2_294(.d_in(u_ca_in_294), .d_out(u_ca_out_294));
compressor_3_2 u_ca_3_2_295(.d_in(u_ca_in_295), .d_out(u_ca_out_295));
compressor_3_2 u_ca_3_2_296(.d_in(u_ca_in_296), .d_out(u_ca_out_296));
compressor_3_2 u_ca_3_2_297(.d_in(u_ca_in_297), .d_out(u_ca_out_297));
compressor_3_2 u_ca_3_2_298(.d_in(u_ca_in_298), .d_out(u_ca_out_298));
compressor_3_2 u_ca_3_2_299(.d_in(u_ca_in_299), .d_out(u_ca_out_299));
compressor_3_2 u_ca_3_2_300(.d_in(u_ca_in_300), .d_out(u_ca_out_300));
compressor_3_2 u_ca_3_2_301(.d_in(u_ca_in_301), .d_out(u_ca_out_301));
compressor_3_2 u_ca_3_2_302(.d_in(u_ca_in_302), .d_out(u_ca_out_302));
compressor_3_2 u_ca_3_2_303(.d_in(u_ca_in_303), .d_out(u_ca_out_303));
compressor_3_2 u_ca_3_2_304(.d_in(u_ca_in_304), .d_out(u_ca_out_304));
compressor_3_2 u_ca_3_2_305(.d_in(u_ca_in_305), .d_out(u_ca_out_305));
compressor_3_2 u_ca_3_2_306(.d_in(u_ca_in_306), .d_out(u_ca_out_306));
compressor_3_2 u_ca_3_2_307(.d_in(u_ca_in_307), .d_out(u_ca_out_307));
compressor_3_2 u_ca_3_2_308(.d_in(u_ca_in_308), .d_out(u_ca_out_308));
compressor_3_2 u_ca_3_2_309(.d_in(u_ca_in_309), .d_out(u_ca_out_309));
compressor_3_2 u_ca_3_2_310(.d_in(u_ca_in_310), .d_out(u_ca_out_310));
compressor_3_2 u_ca_3_2_311(.d_in(u_ca_in_311), .d_out(u_ca_out_311));
compressor_3_2 u_ca_3_2_312(.d_in(u_ca_in_312), .d_out(u_ca_out_312));
compressor_3_2 u_ca_3_2_313(.d_in(u_ca_in_313), .d_out(u_ca_out_313));
compressor_3_2 u_ca_3_2_314(.d_in(u_ca_in_314), .d_out(u_ca_out_314));
compressor_3_2 u_ca_3_2_315(.d_in(u_ca_in_315), .d_out(u_ca_out_315));
compressor_3_2 u_ca_3_2_316(.d_in(u_ca_in_316), .d_out(u_ca_out_316));
compressor_3_2 u_ca_3_2_317(.d_in(u_ca_in_317), .d_out(u_ca_out_317));
compressor_3_2 u_ca_3_2_318(.d_in(u_ca_in_318), .d_out(u_ca_out_318));
compressor_3_2 u_ca_3_2_319(.d_in(u_ca_in_319), .d_out(u_ca_out_319));
compressor_3_2 u_ca_3_2_320(.d_in(u_ca_in_320), .d_out(u_ca_out_320));
compressor_3_2 u_ca_3_2_321(.d_in(u_ca_in_321), .d_out(u_ca_out_321));
compressor_3_2 u_ca_3_2_322(.d_in(u_ca_in_322), .d_out(u_ca_out_322));
compressor_3_2 u_ca_3_2_323(.d_in(u_ca_in_323), .d_out(u_ca_out_323));
compressor_3_2 u_ca_3_2_324(.d_in(u_ca_in_324), .d_out(u_ca_out_324));
compressor_3_2 u_ca_3_2_325(.d_in(u_ca_in_325), .d_out(u_ca_out_325));
compressor_3_2 u_ca_3_2_326(.d_in(u_ca_in_326), .d_out(u_ca_out_326));
compressor_3_2 u_ca_3_2_327(.d_in(u_ca_in_327), .d_out(u_ca_out_327));
compressor_3_2 u_ca_3_2_328(.d_in(u_ca_in_328), .d_out(u_ca_out_328));
compressor_3_2 u_ca_3_2_329(.d_in(u_ca_in_329), .d_out(u_ca_out_329));
compressor_3_2 u_ca_3_2_330(.d_in(u_ca_in_330), .d_out(u_ca_out_330));
compressor_3_2 u_ca_3_2_331(.d_in(u_ca_in_331), .d_out(u_ca_out_331));
compressor_3_2 u_ca_3_2_332(.d_in(u_ca_in_332), .d_out(u_ca_out_332));
compressor_3_2 u_ca_3_2_333(.d_in(u_ca_in_333), .d_out(u_ca_out_333));
compressor_3_2 u_ca_3_2_334(.d_in(u_ca_in_334), .d_out(u_ca_out_334));
compressor_3_2 u_ca_3_2_335(.d_in(u_ca_in_335), .d_out(u_ca_out_335));
compressor_3_2 u_ca_3_2_336(.d_in(u_ca_in_336), .d_out(u_ca_out_336));
compressor_3_2 u_ca_3_2_337(.d_in(u_ca_in_337), .d_out(u_ca_out_337));
compressor_3_2 u_ca_3_2_338(.d_in(u_ca_in_338), .d_out(u_ca_out_338));
compressor_3_2 u_ca_3_2_339(.d_in(u_ca_in_339), .d_out(u_ca_out_339));
compressor_3_2 u_ca_3_2_340(.d_in(u_ca_in_340), .d_out(u_ca_out_340));
compressor_3_2 u_ca_3_2_341(.d_in(u_ca_in_341), .d_out(u_ca_out_341));
compressor_3_2 u_ca_3_2_342(.d_in(u_ca_in_342), .d_out(u_ca_out_342));
compressor_3_2 u_ca_3_2_343(.d_in(u_ca_in_343), .d_out(u_ca_out_343));
compressor_3_2 u_ca_3_2_344(.d_in(u_ca_in_344), .d_out(u_ca_out_344));
compressor_3_2 u_ca_3_2_345(.d_in(u_ca_in_345), .d_out(u_ca_out_345));
compressor_3_2 u_ca_3_2_346(.d_in(u_ca_in_346), .d_out(u_ca_out_346));
compressor_3_2 u_ca_3_2_347(.d_in(u_ca_in_347), .d_out(u_ca_out_347));
compressor_3_2 u_ca_3_2_348(.d_in(u_ca_in_348), .d_out(u_ca_out_348));
compressor_3_2 u_ca_3_2_349(.d_in(u_ca_in_349), .d_out(u_ca_out_349));
compressor_3_2 u_ca_3_2_350(.d_in(u_ca_in_350), .d_out(u_ca_out_350));
compressor_3_2 u_ca_3_2_351(.d_in(u_ca_in_351), .d_out(u_ca_out_351));
compressor_3_2 u_ca_3_2_352(.d_in(u_ca_in_352), .d_out(u_ca_out_352));
compressor_3_2 u_ca_3_2_353(.d_in(u_ca_in_353), .d_out(u_ca_out_353));
compressor_3_2 u_ca_3_2_354(.d_in(u_ca_in_354), .d_out(u_ca_out_354));
compressor_3_2 u_ca_3_2_355(.d_in(u_ca_in_355), .d_out(u_ca_out_355));
compressor_3_2 u_ca_3_2_356(.d_in(u_ca_in_356), .d_out(u_ca_out_356));
compressor_3_2 u_ca_3_2_357(.d_in(u_ca_in_357), .d_out(u_ca_out_357));
compressor_3_2 u_ca_3_2_358(.d_in(u_ca_in_358), .d_out(u_ca_out_358));
compressor_3_2 u_ca_3_2_359(.d_in(u_ca_in_359), .d_out(u_ca_out_359));
compressor_3_2 u_ca_3_2_360(.d_in(u_ca_in_360), .d_out(u_ca_out_360));
compressor_3_2 u_ca_3_2_361(.d_in(u_ca_in_361), .d_out(u_ca_out_361));
compressor_3_2 u_ca_3_2_362(.d_in(u_ca_in_362), .d_out(u_ca_out_362));
compressor_3_2 u_ca_3_2_363(.d_in(u_ca_in_363), .d_out(u_ca_out_363));
compressor_3_2 u_ca_3_2_364(.d_in(u_ca_in_364), .d_out(u_ca_out_364));
compressor_3_2 u_ca_3_2_365(.d_in(u_ca_in_365), .d_out(u_ca_out_365));
compressor_3_2 u_ca_3_2_366(.d_in(u_ca_in_366), .d_out(u_ca_out_366));
compressor_3_2 u_ca_3_2_367(.d_in(u_ca_in_367), .d_out(u_ca_out_367));
compressor_3_2 u_ca_3_2_368(.d_in(u_ca_in_368), .d_out(u_ca_out_368));
compressor_3_2 u_ca_3_2_369(.d_in(u_ca_in_369), .d_out(u_ca_out_369));
compressor_3_2 u_ca_3_2_370(.d_in(u_ca_in_370), .d_out(u_ca_out_370));
compressor_3_2 u_ca_3_2_371(.d_in(u_ca_in_371), .d_out(u_ca_out_371));
compressor_3_2 u_ca_3_2_372(.d_in(u_ca_in_372), .d_out(u_ca_out_372));
compressor_3_2 u_ca_3_2_373(.d_in(u_ca_in_373), .d_out(u_ca_out_373));
compressor_3_2 u_ca_3_2_374(.d_in(u_ca_in_374), .d_out(u_ca_out_374));
compressor_3_2 u_ca_3_2_375(.d_in(u_ca_in_375), .d_out(u_ca_out_375));
compressor_3_2 u_ca_3_2_376(.d_in(u_ca_in_376), .d_out(u_ca_out_376));
compressor_3_2 u_ca_3_2_377(.d_in(u_ca_in_377), .d_out(u_ca_out_377));
compressor_3_2 u_ca_3_2_378(.d_in(u_ca_in_378), .d_out(u_ca_out_378));
compressor_3_2 u_ca_3_2_379(.d_in(u_ca_in_379), .d_out(u_ca_out_379));
compressor_3_2 u_ca_3_2_380(.d_in(u_ca_in_380), .d_out(u_ca_out_380));
compressor_3_2 u_ca_3_2_381(.d_in(u_ca_in_381), .d_out(u_ca_out_381));
compressor_3_2 u_ca_3_2_382(.d_in(u_ca_in_382), .d_out(u_ca_out_382));
compressor_3_2 u_ca_3_2_383(.d_in(u_ca_in_383), .d_out(u_ca_out_383));
compressor_3_2 u_ca_3_2_384(.d_in(u_ca_in_384), .d_out(u_ca_out_384));
compressor_3_2 u_ca_3_2_385(.d_in(u_ca_in_385), .d_out(u_ca_out_385));
compressor_3_2 u_ca_3_2_386(.d_in(u_ca_in_386), .d_out(u_ca_out_386));
compressor_3_2 u_ca_3_2_387(.d_in(u_ca_in_387), .d_out(u_ca_out_387));
compressor_3_2 u_ca_3_2_388(.d_in(u_ca_in_388), .d_out(u_ca_out_388));
compressor_3_2 u_ca_3_2_389(.d_in(u_ca_in_389), .d_out(u_ca_out_389));
compressor_3_2 u_ca_3_2_390(.d_in(u_ca_in_390), .d_out(u_ca_out_390));
compressor_3_2 u_ca_3_2_391(.d_in(u_ca_in_391), .d_out(u_ca_out_391));
compressor_3_2 u_ca_3_2_392(.d_in(u_ca_in_392), .d_out(u_ca_out_392));
compressor_3_2 u_ca_3_2_393(.d_in(u_ca_in_393), .d_out(u_ca_out_393));
compressor_3_2 u_ca_3_2_394(.d_in(u_ca_in_394), .d_out(u_ca_out_394));
compressor_3_2 u_ca_3_2_395(.d_in(u_ca_in_395), .d_out(u_ca_out_395));
compressor_3_2 u_ca_3_2_396(.d_in(u_ca_in_396), .d_out(u_ca_out_396));
compressor_3_2 u_ca_3_2_397(.d_in(u_ca_in_397), .d_out(u_ca_out_397));
compressor_3_2 u_ca_3_2_398(.d_in(u_ca_in_398), .d_out(u_ca_out_398));
compressor_3_2 u_ca_3_2_399(.d_in(u_ca_in_399), .d_out(u_ca_out_399));
compressor_3_2 u_ca_3_2_400(.d_in(u_ca_in_400), .d_out(u_ca_out_400));
compressor_3_2 u_ca_3_2_401(.d_in(u_ca_in_401), .d_out(u_ca_out_401));
compressor_3_2 u_ca_3_2_402(.d_in(u_ca_in_402), .d_out(u_ca_out_402));
compressor_3_2 u_ca_3_2_403(.d_in(u_ca_in_403), .d_out(u_ca_out_403));
compressor_3_2 u_ca_3_2_404(.d_in(u_ca_in_404), .d_out(u_ca_out_404));
compressor_3_2 u_ca_3_2_405(.d_in(u_ca_in_405), .d_out(u_ca_out_405));
compressor_3_2 u_ca_3_2_406(.d_in(u_ca_in_406), .d_out(u_ca_out_406));
compressor_3_2 u_ca_3_2_407(.d_in(u_ca_in_407), .d_out(u_ca_out_407));
compressor_3_2 u_ca_3_2_408(.d_in(u_ca_in_408), .d_out(u_ca_out_408));
compressor_3_2 u_ca_3_2_409(.d_in(u_ca_in_409), .d_out(u_ca_out_409));
compressor_3_2 u_ca_3_2_410(.d_in(u_ca_in_410), .d_out(u_ca_out_410));
compressor_3_2 u_ca_3_2_411(.d_in(u_ca_in_411), .d_out(u_ca_out_411));
compressor_3_2 u_ca_3_2_412(.d_in(u_ca_in_412), .d_out(u_ca_out_412));
compressor_3_2 u_ca_3_2_413(.d_in(u_ca_in_413), .d_out(u_ca_out_413));
compressor_3_2 u_ca_3_2_414(.d_in(u_ca_in_414), .d_out(u_ca_out_414));
compressor_3_2 u_ca_3_2_415(.d_in(u_ca_in_415), .d_out(u_ca_out_415));
compressor_3_2 u_ca_3_2_416(.d_in(u_ca_in_416), .d_out(u_ca_out_416));
compressor_3_2 u_ca_3_2_417(.d_in(u_ca_in_417), .d_out(u_ca_out_417));
compressor_3_2 u_ca_3_2_418(.d_in(u_ca_in_418), .d_out(u_ca_out_418));
compressor_3_2 u_ca_3_2_419(.d_in(u_ca_in_419), .d_out(u_ca_out_419));
compressor_3_2 u_ca_3_2_420(.d_in(u_ca_in_420), .d_out(u_ca_out_420));
compressor_3_2 u_ca_3_2_421(.d_in(u_ca_in_421), .d_out(u_ca_out_421));
compressor_3_2 u_ca_3_2_422(.d_in(u_ca_in_422), .d_out(u_ca_out_422));
compressor_3_2 u_ca_3_2_423(.d_in(u_ca_in_423), .d_out(u_ca_out_423));
compressor_3_2 u_ca_3_2_424(.d_in(u_ca_in_424), .d_out(u_ca_out_424));
compressor_3_2 u_ca_3_2_425(.d_in(u_ca_in_425), .d_out(u_ca_out_425));
compressor_3_2 u_ca_3_2_426(.d_in(u_ca_in_426), .d_out(u_ca_out_426));
compressor_3_2 u_ca_3_2_427(.d_in(u_ca_in_427), .d_out(u_ca_out_427));
compressor_3_2 u_ca_3_2_428(.d_in(u_ca_in_428), .d_out(u_ca_out_428));
compressor_3_2 u_ca_3_2_429(.d_in(u_ca_in_429), .d_out(u_ca_out_429));
compressor_3_2 u_ca_3_2_430(.d_in(u_ca_in_430), .d_out(u_ca_out_430));
compressor_3_2 u_ca_3_2_431(.d_in(u_ca_in_431), .d_out(u_ca_out_431));
compressor_3_2 u_ca_3_2_432(.d_in(u_ca_in_432), .d_out(u_ca_out_432));
compressor_3_2 u_ca_3_2_433(.d_in(u_ca_in_433), .d_out(u_ca_out_433));
compressor_3_2 u_ca_3_2_434(.d_in(u_ca_in_434), .d_out(u_ca_out_434));
compressor_3_2 u_ca_3_2_435(.d_in(u_ca_in_435), .d_out(u_ca_out_435));
compressor_3_2 u_ca_3_2_436(.d_in(u_ca_in_436), .d_out(u_ca_out_436));
compressor_3_2 u_ca_3_2_437(.d_in(u_ca_in_437), .d_out(u_ca_out_437));
compressor_3_2 u_ca_3_2_438(.d_in(u_ca_in_438), .d_out(u_ca_out_438));
compressor_3_2 u_ca_3_2_439(.d_in(u_ca_in_439), .d_out(u_ca_out_439));
compressor_3_2 u_ca_3_2_440(.d_in(u_ca_in_440), .d_out(u_ca_out_440));
compressor_3_2 u_ca_3_2_441(.d_in(u_ca_in_441), .d_out(u_ca_out_441));
compressor_3_2 u_ca_3_2_442(.d_in(u_ca_in_442), .d_out(u_ca_out_442));
compressor_3_2 u_ca_3_2_443(.d_in(u_ca_in_443), .d_out(u_ca_out_443));
compressor_3_2 u_ca_3_2_444(.d_in(u_ca_in_444), .d_out(u_ca_out_444));
compressor_3_2 u_ca_3_2_445(.d_in(u_ca_in_445), .d_out(u_ca_out_445));
compressor_3_2 u_ca_3_2_446(.d_in(u_ca_in_446), .d_out(u_ca_out_446));
compressor_3_2 u_ca_3_2_447(.d_in(u_ca_in_447), .d_out(u_ca_out_447));
compressor_3_2 u_ca_3_2_448(.d_in(u_ca_in_448), .d_out(u_ca_out_448));
compressor_3_2 u_ca_3_2_449(.d_in(u_ca_in_449), .d_out(u_ca_out_449));
compressor_3_2 u_ca_3_2_450(.d_in(u_ca_in_450), .d_out(u_ca_out_450));
compressor_3_2 u_ca_3_2_451(.d_in(u_ca_in_451), .d_out(u_ca_out_451));
compressor_3_2 u_ca_3_2_452(.d_in(u_ca_in_452), .d_out(u_ca_out_452));
compressor_3_2 u_ca_3_2_453(.d_in(u_ca_in_453), .d_out(u_ca_out_453));
compressor_3_2 u_ca_3_2_454(.d_in(u_ca_in_454), .d_out(u_ca_out_454));
compressor_3_2 u_ca_3_2_455(.d_in(u_ca_in_455), .d_out(u_ca_out_455));
compressor_3_2 u_ca_3_2_456(.d_in(u_ca_in_456), .d_out(u_ca_out_456));
compressor_3_2 u_ca_3_2_457(.d_in(u_ca_in_457), .d_out(u_ca_out_457));
compressor_3_2 u_ca_3_2_458(.d_in(u_ca_in_458), .d_out(u_ca_out_458));
compressor_3_2 u_ca_3_2_459(.d_in(u_ca_in_459), .d_out(u_ca_out_459));
compressor_3_2 u_ca_3_2_460(.d_in(u_ca_in_460), .d_out(u_ca_out_460));
compressor_3_2 u_ca_3_2_461(.d_in(u_ca_in_461), .d_out(u_ca_out_461));
compressor_3_2 u_ca_3_2_462(.d_in(u_ca_in_462), .d_out(u_ca_out_462));
compressor_3_2 u_ca_3_2_463(.d_in(u_ca_in_463), .d_out(u_ca_out_463));
compressor_3_2 u_ca_3_2_464(.d_in(u_ca_in_464), .d_out(u_ca_out_464));
compressor_3_2 u_ca_3_2_465(.d_in(u_ca_in_465), .d_out(u_ca_out_465));
compressor_3_2 u_ca_3_2_466(.d_in(u_ca_in_466), .d_out(u_ca_out_466));
compressor_3_2 u_ca_3_2_467(.d_in(u_ca_in_467), .d_out(u_ca_out_467));
compressor_3_2 u_ca_3_2_468(.d_in(u_ca_in_468), .d_out(u_ca_out_468));
compressor_3_2 u_ca_3_2_469(.d_in(u_ca_in_469), .d_out(u_ca_out_469));
compressor_3_2 u_ca_3_2_470(.d_in(u_ca_in_470), .d_out(u_ca_out_470));
compressor_3_2 u_ca_3_2_471(.d_in(u_ca_in_471), .d_out(u_ca_out_471));
compressor_3_2 u_ca_3_2_472(.d_in(u_ca_in_472), .d_out(u_ca_out_472));
compressor_3_2 u_ca_3_2_473(.d_in(u_ca_in_473), .d_out(u_ca_out_473));
compressor_3_2 u_ca_3_2_474(.d_in(u_ca_in_474), .d_out(u_ca_out_474));
compressor_3_2 u_ca_3_2_475(.d_in(u_ca_in_475), .d_out(u_ca_out_475));
compressor_3_2 u_ca_3_2_476(.d_in(u_ca_in_476), .d_out(u_ca_out_476));
compressor_3_2 u_ca_3_2_477(.d_in(u_ca_in_477), .d_out(u_ca_out_477));
compressor_3_2 u_ca_3_2_478(.d_in(u_ca_in_478), .d_out(u_ca_out_478));
compressor_3_2 u_ca_3_2_479(.d_in(u_ca_in_479), .d_out(u_ca_out_479));
compressor_3_2 u_ca_3_2_480(.d_in(u_ca_in_480), .d_out(u_ca_out_480));
compressor_3_2 u_ca_3_2_481(.d_in(u_ca_in_481), .d_out(u_ca_out_481));
compressor_3_2 u_ca_3_2_482(.d_in(u_ca_in_482), .d_out(u_ca_out_482));
compressor_3_2 u_ca_3_2_483(.d_in(u_ca_in_483), .d_out(u_ca_out_483));
compressor_3_2 u_ca_3_2_484(.d_in(u_ca_in_484), .d_out(u_ca_out_484));
compressor_3_2 u_ca_3_2_485(.d_in(u_ca_in_485), .d_out(u_ca_out_485));
compressor_3_2 u_ca_3_2_486(.d_in(u_ca_in_486), .d_out(u_ca_out_486));
compressor_3_2 u_ca_3_2_487(.d_in(u_ca_in_487), .d_out(u_ca_out_487));
compressor_3_2 u_ca_3_2_488(.d_in(u_ca_in_488), .d_out(u_ca_out_488));
compressor_3_2 u_ca_3_2_489(.d_in(u_ca_in_489), .d_out(u_ca_out_489));
compressor_3_2 u_ca_3_2_490(.d_in(u_ca_in_490), .d_out(u_ca_out_490));
compressor_3_2 u_ca_3_2_491(.d_in(u_ca_in_491), .d_out(u_ca_out_491));
compressor_3_2 u_ca_3_2_492(.d_in(u_ca_in_492), .d_out(u_ca_out_492));
compressor_3_2 u_ca_3_2_493(.d_in(u_ca_in_493), .d_out(u_ca_out_493));
compressor_3_2 u_ca_3_2_494(.d_in(u_ca_in_494), .d_out(u_ca_out_494));
compressor_3_2 u_ca_3_2_495(.d_in(u_ca_in_495), .d_out(u_ca_out_495));
compressor_3_2 u_ca_3_2_496(.d_in(u_ca_in_496), .d_out(u_ca_out_496));
compressor_3_2 u_ca_3_2_497(.d_in(u_ca_in_497), .d_out(u_ca_out_497));
compressor_3_2 u_ca_3_2_498(.d_in(u_ca_in_498), .d_out(u_ca_out_498));
compressor_3_2 u_ca_3_2_499(.d_in(u_ca_in_499), .d_out(u_ca_out_499));
compressor_3_2 u_ca_3_2_500(.d_in(u_ca_in_500), .d_out(u_ca_out_500));
compressor_3_2 u_ca_3_2_501(.d_in(u_ca_in_501), .d_out(u_ca_out_501));
compressor_3_2 u_ca_3_2_502(.d_in(u_ca_in_502), .d_out(u_ca_out_502));
compressor_3_2 u_ca_3_2_503(.d_in(u_ca_in_503), .d_out(u_ca_out_503));
compressor_3_2 u_ca_3_2_504(.d_in(u_ca_in_504), .d_out(u_ca_out_504));
compressor_3_2 u_ca_3_2_505(.d_in(u_ca_in_505), .d_out(u_ca_out_505));
compressor_3_2 u_ca_3_2_506(.d_in(u_ca_in_506), .d_out(u_ca_out_506));
compressor_3_2 u_ca_3_2_507(.d_in(u_ca_in_507), .d_out(u_ca_out_507));
compressor_3_2 u_ca_3_2_508(.d_in(u_ca_in_508), .d_out(u_ca_out_508));
compressor_3_2 u_ca_3_2_509(.d_in(u_ca_in_509), .d_out(u_ca_out_509));
compressor_3_2 u_ca_3_2_510(.d_in(u_ca_in_510), .d_out(u_ca_out_510));
compressor_3_2 u_ca_3_2_511(.d_in(u_ca_in_511), .d_out(u_ca_out_511));
compressor_3_2 u_ca_3_2_512(.d_in(u_ca_in_512), .d_out(u_ca_out_512));
compressor_3_2 u_ca_3_2_513(.d_in(u_ca_in_513), .d_out(u_ca_out_513));
compressor_3_2 u_ca_3_2_514(.d_in(u_ca_in_514), .d_out(u_ca_out_514));
compressor_3_2 u_ca_3_2_515(.d_in(u_ca_in_515), .d_out(u_ca_out_515));
compressor_3_2 u_ca_3_2_516(.d_in(u_ca_in_516), .d_out(u_ca_out_516));
compressor_3_2 u_ca_3_2_517(.d_in(u_ca_in_517), .d_out(u_ca_out_517));
compressor_3_2 u_ca_3_2_518(.d_in(u_ca_in_518), .d_out(u_ca_out_518));
compressor_3_2 u_ca_3_2_519(.d_in(u_ca_in_519), .d_out(u_ca_out_519));
compressor_3_2 u_ca_3_2_520(.d_in(u_ca_in_520), .d_out(u_ca_out_520));
compressor_3_2 u_ca_3_2_521(.d_in(u_ca_in_521), .d_out(u_ca_out_521));
compressor_3_2 u_ca_3_2_522(.d_in(u_ca_in_522), .d_out(u_ca_out_522));
compressor_3_2 u_ca_3_2_523(.d_in(u_ca_in_523), .d_out(u_ca_out_523));
compressor_3_2 u_ca_3_2_524(.d_in(u_ca_in_524), .d_out(u_ca_out_524));
compressor_3_2 u_ca_3_2_525(.d_in(u_ca_in_525), .d_out(u_ca_out_525));
compressor_3_2 u_ca_3_2_526(.d_in(u_ca_in_526), .d_out(u_ca_out_526));
compressor_3_2 u_ca_3_2_527(.d_in(u_ca_in_527), .d_out(u_ca_out_527));
compressor_3_2 u_ca_3_2_528(.d_in(u_ca_in_528), .d_out(u_ca_out_528));
compressor_3_2 u_ca_3_2_529(.d_in(u_ca_in_529), .d_out(u_ca_out_529));
compressor_3_2 u_ca_3_2_530(.d_in(u_ca_in_530), .d_out(u_ca_out_530));
compressor_3_2 u_ca_3_2_531(.d_in(u_ca_in_531), .d_out(u_ca_out_531));
compressor_3_2 u_ca_3_2_532(.d_in(u_ca_in_532), .d_out(u_ca_out_532));
compressor_3_2 u_ca_3_2_533(.d_in(u_ca_in_533), .d_out(u_ca_out_533));
compressor_3_2 u_ca_3_2_534(.d_in(u_ca_in_534), .d_out(u_ca_out_534));
compressor_3_2 u_ca_3_2_535(.d_in(u_ca_in_535), .d_out(u_ca_out_535));
compressor_3_2 u_ca_3_2_536(.d_in(u_ca_in_536), .d_out(u_ca_out_536));
compressor_3_2 u_ca_3_2_537(.d_in(u_ca_in_537), .d_out(u_ca_out_537));
compressor_3_2 u_ca_3_2_538(.d_in(u_ca_in_538), .d_out(u_ca_out_538));
compressor_3_2 u_ca_3_2_539(.d_in(u_ca_in_539), .d_out(u_ca_out_539));
compressor_3_2 u_ca_3_2_540(.d_in(u_ca_in_540), .d_out(u_ca_out_540));
compressor_3_2 u_ca_3_2_541(.d_in(u_ca_in_541), .d_out(u_ca_out_541));
compressor_3_2 u_ca_3_2_542(.d_in(u_ca_in_542), .d_out(u_ca_out_542));
compressor_3_2 u_ca_3_2_543(.d_in(u_ca_in_543), .d_out(u_ca_out_543));
compressor_3_2 u_ca_3_2_544(.d_in(u_ca_in_544), .d_out(u_ca_out_544));
compressor_3_2 u_ca_3_2_545(.d_in(u_ca_in_545), .d_out(u_ca_out_545));
compressor_3_2 u_ca_3_2_546(.d_in(u_ca_in_546), .d_out(u_ca_out_546));
compressor_3_2 u_ca_3_2_547(.d_in(u_ca_in_547), .d_out(u_ca_out_547));
compressor_3_2 u_ca_3_2_548(.d_in(u_ca_in_548), .d_out(u_ca_out_548));
compressor_3_2 u_ca_3_2_549(.d_in(u_ca_in_549), .d_out(u_ca_out_549));
compressor_3_2 u_ca_3_2_550(.d_in(u_ca_in_550), .d_out(u_ca_out_550));
compressor_3_2 u_ca_3_2_551(.d_in(u_ca_in_551), .d_out(u_ca_out_551));
compressor_3_2 u_ca_3_2_552(.d_in(u_ca_in_552), .d_out(u_ca_out_552));
compressor_3_2 u_ca_3_2_553(.d_in(u_ca_in_553), .d_out(u_ca_out_553));
compressor_3_2 u_ca_3_2_554(.d_in(u_ca_in_554), .d_out(u_ca_out_554));
compressor_3_2 u_ca_3_2_555(.d_in(u_ca_in_555), .d_out(u_ca_out_555));
compressor_3_2 u_ca_3_2_556(.d_in(u_ca_in_556), .d_out(u_ca_out_556));
compressor_3_2 u_ca_3_2_557(.d_in(u_ca_in_557), .d_out(u_ca_out_557));
compressor_3_2 u_ca_3_2_558(.d_in(u_ca_in_558), .d_out(u_ca_out_558));
compressor_3_2 u_ca_3_2_559(.d_in(u_ca_in_559), .d_out(u_ca_out_559));
compressor_3_2 u_ca_3_2_560(.d_in(u_ca_in_560), .d_out(u_ca_out_560));
compressor_3_2 u_ca_3_2_561(.d_in(u_ca_in_561), .d_out(u_ca_out_561));
compressor_3_2 u_ca_3_2_562(.d_in(u_ca_in_562), .d_out(u_ca_out_562));
compressor_3_2 u_ca_3_2_563(.d_in(u_ca_in_563), .d_out(u_ca_out_563));
compressor_3_2 u_ca_3_2_564(.d_in(u_ca_in_564), .d_out(u_ca_out_564));
compressor_3_2 u_ca_3_2_565(.d_in(u_ca_in_565), .d_out(u_ca_out_565));
compressor_3_2 u_ca_3_2_566(.d_in(u_ca_in_566), .d_out(u_ca_out_566));
compressor_3_2 u_ca_3_2_567(.d_in(u_ca_in_567), .d_out(u_ca_out_567));
compressor_3_2 u_ca_3_2_568(.d_in(u_ca_in_568), .d_out(u_ca_out_568));
compressor_3_2 u_ca_3_2_569(.d_in(u_ca_in_569), .d_out(u_ca_out_569));
compressor_3_2 u_ca_3_2_570(.d_in(u_ca_in_570), .d_out(u_ca_out_570));
compressor_3_2 u_ca_3_2_571(.d_in(u_ca_in_571), .d_out(u_ca_out_571));
compressor_3_2 u_ca_3_2_572(.d_in(u_ca_in_572), .d_out(u_ca_out_572));
compressor_3_2 u_ca_3_2_573(.d_in(u_ca_in_573), .d_out(u_ca_out_573));
compressor_3_2 u_ca_3_2_574(.d_in(u_ca_in_574), .d_out(u_ca_out_574));
compressor_3_2 u_ca_3_2_575(.d_in(u_ca_in_575), .d_out(u_ca_out_575));
compressor_3_2 u_ca_3_2_576(.d_in(u_ca_in_576), .d_out(u_ca_out_576));
compressor_3_2 u_ca_3_2_577(.d_in(u_ca_in_577), .d_out(u_ca_out_577));
compressor_3_2 u_ca_3_2_578(.d_in(u_ca_in_578), .d_out(u_ca_out_578));
compressor_3_2 u_ca_3_2_579(.d_in(u_ca_in_579), .d_out(u_ca_out_579));
compressor_3_2 u_ca_3_2_580(.d_in(u_ca_in_580), .d_out(u_ca_out_580));
compressor_3_2 u_ca_3_2_581(.d_in(u_ca_in_581), .d_out(u_ca_out_581));
compressor_3_2 u_ca_3_2_582(.d_in(u_ca_in_582), .d_out(u_ca_out_582));
compressor_3_2 u_ca_3_2_583(.d_in(u_ca_in_583), .d_out(u_ca_out_583));
compressor_3_2 u_ca_3_2_584(.d_in(u_ca_in_584), .d_out(u_ca_out_584));
compressor_3_2 u_ca_3_2_585(.d_in(u_ca_in_585), .d_out(u_ca_out_585));
compressor_3_2 u_ca_3_2_586(.d_in(u_ca_in_586), .d_out(u_ca_out_586));
compressor_3_2 u_ca_3_2_587(.d_in(u_ca_in_587), .d_out(u_ca_out_587));
compressor_3_2 u_ca_3_2_588(.d_in(u_ca_in_588), .d_out(u_ca_out_588));
compressor_3_2 u_ca_3_2_589(.d_in(u_ca_in_589), .d_out(u_ca_out_589));
compressor_3_2 u_ca_3_2_590(.d_in(u_ca_in_590), .d_out(u_ca_out_590));
compressor_3_2 u_ca_3_2_591(.d_in(u_ca_in_591), .d_out(u_ca_out_591));
compressor_3_2 u_ca_3_2_592(.d_in(u_ca_in_592), .d_out(u_ca_out_592));
compressor_3_2 u_ca_3_2_593(.d_in(u_ca_in_593), .d_out(u_ca_out_593));
compressor_3_2 u_ca_3_2_594(.d_in(u_ca_in_594), .d_out(u_ca_out_594));
compressor_3_2 u_ca_3_2_595(.d_in(u_ca_in_595), .d_out(u_ca_out_595));
compressor_3_2 u_ca_3_2_596(.d_in(u_ca_in_596), .d_out(u_ca_out_596));
compressor_3_2 u_ca_3_2_597(.d_in(u_ca_in_597), .d_out(u_ca_out_597));
compressor_3_2 u_ca_3_2_598(.d_in(u_ca_in_598), .d_out(u_ca_out_598));
compressor_3_2 u_ca_3_2_599(.d_in(u_ca_in_599), .d_out(u_ca_out_599));
compressor_3_2 u_ca_3_2_600(.d_in(u_ca_in_600), .d_out(u_ca_out_600));
compressor_3_2 u_ca_3_2_601(.d_in(u_ca_in_601), .d_out(u_ca_out_601));
compressor_3_2 u_ca_3_2_602(.d_in(u_ca_in_602), .d_out(u_ca_out_602));
compressor_3_2 u_ca_3_2_603(.d_in(u_ca_in_603), .d_out(u_ca_out_603));
compressor_3_2 u_ca_3_2_604(.d_in(u_ca_in_604), .d_out(u_ca_out_604));
compressor_3_2 u_ca_3_2_605(.d_in(u_ca_in_605), .d_out(u_ca_out_605));
compressor_3_2 u_ca_3_2_606(.d_in(u_ca_in_606), .d_out(u_ca_out_606));
compressor_3_2 u_ca_3_2_607(.d_in(u_ca_in_607), .d_out(u_ca_out_607));
compressor_3_2 u_ca_3_2_608(.d_in(u_ca_in_608), .d_out(u_ca_out_608));
compressor_3_2 u_ca_3_2_609(.d_in(u_ca_in_609), .d_out(u_ca_out_609));
compressor_3_2 u_ca_3_2_610(.d_in(u_ca_in_610), .d_out(u_ca_out_610));
compressor_3_2 u_ca_3_2_611(.d_in(u_ca_in_611), .d_out(u_ca_out_611));
compressor_3_2 u_ca_3_2_612(.d_in(u_ca_in_612), .d_out(u_ca_out_612));
compressor_3_2 u_ca_3_2_613(.d_in(u_ca_in_613), .d_out(u_ca_out_613));
compressor_3_2 u_ca_3_2_614(.d_in(u_ca_in_614), .d_out(u_ca_out_614));
compressor_3_2 u_ca_3_2_615(.d_in(u_ca_in_615), .d_out(u_ca_out_615));
compressor_3_2 u_ca_3_2_616(.d_in(u_ca_in_616), .d_out(u_ca_out_616));
compressor_3_2 u_ca_3_2_617(.d_in(u_ca_in_617), .d_out(u_ca_out_617));
compressor_3_2 u_ca_3_2_618(.d_in(u_ca_in_618), .d_out(u_ca_out_618));
compressor_3_2 u_ca_3_2_619(.d_in(u_ca_in_619), .d_out(u_ca_out_619));
compressor_3_2 u_ca_3_2_620(.d_in(u_ca_in_620), .d_out(u_ca_out_620));
compressor_3_2 u_ca_3_2_621(.d_in(u_ca_in_621), .d_out(u_ca_out_621));
compressor_3_2 u_ca_3_2_622(.d_in(u_ca_in_622), .d_out(u_ca_out_622));
compressor_3_2 u_ca_3_2_623(.d_in(u_ca_in_623), .d_out(u_ca_out_623));
compressor_3_2 u_ca_3_2_624(.d_in(u_ca_in_624), .d_out(u_ca_out_624));
compressor_3_2 u_ca_3_2_625(.d_in(u_ca_in_625), .d_out(u_ca_out_625));
compressor_3_2 u_ca_3_2_626(.d_in(u_ca_in_626), .d_out(u_ca_out_626));
compressor_3_2 u_ca_3_2_627(.d_in(u_ca_in_627), .d_out(u_ca_out_627));
compressor_3_2 u_ca_3_2_628(.d_in(u_ca_in_628), .d_out(u_ca_out_628));
compressor_3_2 u_ca_3_2_629(.d_in(u_ca_in_629), .d_out(u_ca_out_629));
compressor_3_2 u_ca_3_2_630(.d_in(u_ca_in_630), .d_out(u_ca_out_630));
compressor_3_2 u_ca_3_2_631(.d_in(u_ca_in_631), .d_out(u_ca_out_631));
compressor_3_2 u_ca_3_2_632(.d_in(u_ca_in_632), .d_out(u_ca_out_632));
compressor_3_2 u_ca_3_2_633(.d_in(u_ca_in_633), .d_out(u_ca_out_633));
compressor_3_2 u_ca_3_2_634(.d_in(u_ca_in_634), .d_out(u_ca_out_634));
compressor_3_2 u_ca_3_2_635(.d_in(u_ca_in_635), .d_out(u_ca_out_635));
compressor_3_2 u_ca_3_2_636(.d_in(u_ca_in_636), .d_out(u_ca_out_636));
compressor_3_2 u_ca_3_2_637(.d_in(u_ca_in_637), .d_out(u_ca_out_637));
compressor_3_2 u_ca_3_2_638(.d_in(u_ca_in_638), .d_out(u_ca_out_638));
compressor_3_2 u_ca_3_2_639(.d_in(u_ca_in_639), .d_out(u_ca_out_639));
compressor_3_2 u_ca_3_2_640(.d_in(u_ca_in_640), .d_out(u_ca_out_640));
compressor_3_2 u_ca_3_2_641(.d_in(u_ca_in_641), .d_out(u_ca_out_641));
compressor_3_2 u_ca_3_2_642(.d_in(u_ca_in_642), .d_out(u_ca_out_642));
compressor_3_2 u_ca_3_2_643(.d_in(u_ca_in_643), .d_out(u_ca_out_643));
compressor_3_2 u_ca_3_2_644(.d_in(u_ca_in_644), .d_out(u_ca_out_644));
compressor_3_2 u_ca_3_2_645(.d_in(u_ca_in_645), .d_out(u_ca_out_645));
compressor_3_2 u_ca_3_2_646(.d_in(u_ca_in_646), .d_out(u_ca_out_646));
compressor_3_2 u_ca_3_2_647(.d_in(u_ca_in_647), .d_out(u_ca_out_647));
compressor_3_2 u_ca_3_2_648(.d_in(u_ca_in_648), .d_out(u_ca_out_648));
compressor_3_2 u_ca_3_2_649(.d_in(u_ca_in_649), .d_out(u_ca_out_649));
compressor_3_2 u_ca_3_2_650(.d_in(u_ca_in_650), .d_out(u_ca_out_650));
compressor_3_2 u_ca_3_2_651(.d_in(u_ca_in_651), .d_out(u_ca_out_651));
compressor_3_2 u_ca_3_2_652(.d_in(u_ca_in_652), .d_out(u_ca_out_652));
compressor_3_2 u_ca_3_2_653(.d_in(u_ca_in_653), .d_out(u_ca_out_653));
compressor_3_2 u_ca_3_2_654(.d_in(u_ca_in_654), .d_out(u_ca_out_654));
compressor_3_2 u_ca_3_2_655(.d_in(u_ca_in_655), .d_out(u_ca_out_655));
compressor_3_2 u_ca_3_2_656(.d_in(u_ca_in_656), .d_out(u_ca_out_656));
compressor_3_2 u_ca_3_2_657(.d_in(u_ca_in_657), .d_out(u_ca_out_657));
compressor_3_2 u_ca_3_2_658(.d_in(u_ca_in_658), .d_out(u_ca_out_658));
compressor_3_2 u_ca_3_2_659(.d_in(u_ca_in_659), .d_out(u_ca_out_659));
compressor_3_2 u_ca_3_2_660(.d_in(u_ca_in_660), .d_out(u_ca_out_660));
compressor_3_2 u_ca_3_2_661(.d_in(u_ca_in_661), .d_out(u_ca_out_661));
compressor_3_2 u_ca_3_2_662(.d_in(u_ca_in_662), .d_out(u_ca_out_662));
compressor_3_2 u_ca_3_2_663(.d_in(u_ca_in_663), .d_out(u_ca_out_663));
compressor_3_2 u_ca_3_2_664(.d_in(u_ca_in_664), .d_out(u_ca_out_664));
compressor_3_2 u_ca_3_2_665(.d_in(u_ca_in_665), .d_out(u_ca_out_665));
compressor_3_2 u_ca_3_2_666(.d_in(u_ca_in_666), .d_out(u_ca_out_666));
compressor_3_2 u_ca_3_2_667(.d_in(u_ca_in_667), .d_out(u_ca_out_667));
compressor_3_2 u_ca_3_2_668(.d_in(u_ca_in_668), .d_out(u_ca_out_668));
compressor_3_2 u_ca_3_2_669(.d_in(u_ca_in_669), .d_out(u_ca_out_669));
compressor_3_2 u_ca_3_2_670(.d_in(u_ca_in_670), .d_out(u_ca_out_670));
compressor_3_2 u_ca_3_2_671(.d_in(u_ca_in_671), .d_out(u_ca_out_671));
compressor_3_2 u_ca_3_2_672(.d_in(u_ca_in_672), .d_out(u_ca_out_672));
compressor_3_2 u_ca_3_2_673(.d_in(u_ca_in_673), .d_out(u_ca_out_673));
compressor_3_2 u_ca_3_2_674(.d_in(u_ca_in_674), .d_out(u_ca_out_674));
compressor_3_2 u_ca_3_2_675(.d_in(u_ca_in_675), .d_out(u_ca_out_675));
compressor_3_2 u_ca_3_2_676(.d_in(u_ca_in_676), .d_out(u_ca_out_676));
compressor_3_2 u_ca_3_2_677(.d_in(u_ca_in_677), .d_out(u_ca_out_677));
compressor_3_2 u_ca_3_2_678(.d_in(u_ca_in_678), .d_out(u_ca_out_678));
compressor_3_2 u_ca_3_2_679(.d_in(u_ca_in_679), .d_out(u_ca_out_679));
compressor_3_2 u_ca_3_2_680(.d_in(u_ca_in_680), .d_out(u_ca_out_680));
compressor_3_2 u_ca_3_2_681(.d_in(u_ca_in_681), .d_out(u_ca_out_681));
compressor_3_2 u_ca_3_2_682(.d_in(u_ca_in_682), .d_out(u_ca_out_682));
compressor_3_2 u_ca_3_2_683(.d_in(u_ca_in_683), .d_out(u_ca_out_683));
compressor_3_2 u_ca_3_2_684(.d_in(u_ca_in_684), .d_out(u_ca_out_684));
compressor_3_2 u_ca_3_2_685(.d_in(u_ca_in_685), .d_out(u_ca_out_685));
compressor_3_2 u_ca_3_2_686(.d_in(u_ca_in_686), .d_out(u_ca_out_686));
compressor_3_2 u_ca_3_2_687(.d_in(u_ca_in_687), .d_out(u_ca_out_687));
compressor_3_2 u_ca_3_2_688(.d_in(u_ca_in_688), .d_out(u_ca_out_688));
compressor_3_2 u_ca_3_2_689(.d_in(u_ca_in_689), .d_out(u_ca_out_689));
compressor_3_2 u_ca_3_2_690(.d_in(u_ca_in_690), .d_out(u_ca_out_690));
compressor_3_2 u_ca_3_2_691(.d_in(u_ca_in_691), .d_out(u_ca_out_691));
compressor_3_2 u_ca_3_2_692(.d_in(u_ca_in_692), .d_out(u_ca_out_692));
compressor_3_2 u_ca_3_2_693(.d_in(u_ca_in_693), .d_out(u_ca_out_693));
compressor_3_2 u_ca_3_2_694(.d_in(u_ca_in_694), .d_out(u_ca_out_694));
compressor_3_2 u_ca_3_2_695(.d_in(u_ca_in_695), .d_out(u_ca_out_695));
compressor_3_2 u_ca_3_2_696(.d_in(u_ca_in_696), .d_out(u_ca_out_696));
compressor_3_2 u_ca_3_2_697(.d_in(u_ca_in_697), .d_out(u_ca_out_697));
compressor_3_2 u_ca_3_2_698(.d_in(u_ca_in_698), .d_out(u_ca_out_698));
compressor_3_2 u_ca_3_2_699(.d_in(u_ca_in_699), .d_out(u_ca_out_699));
compressor_3_2 u_ca_3_2_700(.d_in(u_ca_in_700), .d_out(u_ca_out_700));
compressor_3_2 u_ca_3_2_701(.d_in(u_ca_in_701), .d_out(u_ca_out_701));
compressor_3_2 u_ca_3_2_702(.d_in(u_ca_in_702), .d_out(u_ca_out_702));
compressor_3_2 u_ca_3_2_703(.d_in(u_ca_in_703), .d_out(u_ca_out_703));
compressor_3_2 u_ca_3_2_704(.d_in(u_ca_in_704), .d_out(u_ca_out_704));
compressor_3_2 u_ca_3_2_705(.d_in(u_ca_in_705), .d_out(u_ca_out_705));
compressor_3_2 u_ca_3_2_706(.d_in(u_ca_in_706), .d_out(u_ca_out_706));
compressor_3_2 u_ca_3_2_707(.d_in(u_ca_in_707), .d_out(u_ca_out_707));
compressor_3_2 u_ca_3_2_708(.d_in(u_ca_in_708), .d_out(u_ca_out_708));
compressor_3_2 u_ca_3_2_709(.d_in(u_ca_in_709), .d_out(u_ca_out_709));
compressor_3_2 u_ca_3_2_710(.d_in(u_ca_in_710), .d_out(u_ca_out_710));
compressor_3_2 u_ca_3_2_711(.d_in(u_ca_in_711), .d_out(u_ca_out_711));
compressor_3_2 u_ca_3_2_712(.d_in(u_ca_in_712), .d_out(u_ca_out_712));
compressor_3_2 u_ca_3_2_713(.d_in(u_ca_in_713), .d_out(u_ca_out_713));
compressor_3_2 u_ca_3_2_714(.d_in(u_ca_in_714), .d_out(u_ca_out_714));
compressor_3_2 u_ca_3_2_715(.d_in(u_ca_in_715), .d_out(u_ca_out_715));
compressor_3_2 u_ca_3_2_716(.d_in(u_ca_in_716), .d_out(u_ca_out_716));
compressor_3_2 u_ca_3_2_717(.d_in(u_ca_in_717), .d_out(u_ca_out_717));
compressor_3_2 u_ca_3_2_718(.d_in(u_ca_in_718), .d_out(u_ca_out_718));
compressor_3_2 u_ca_3_2_719(.d_in(u_ca_in_719), .d_out(u_ca_out_719));
compressor_3_2 u_ca_3_2_720(.d_in(u_ca_in_720), .d_out(u_ca_out_720));
compressor_3_2 u_ca_3_2_721(.d_in(u_ca_in_721), .d_out(u_ca_out_721));
compressor_3_2 u_ca_3_2_722(.d_in(u_ca_in_722), .d_out(u_ca_out_722));
compressor_3_2 u_ca_3_2_723(.d_in(u_ca_in_723), .d_out(u_ca_out_723));
compressor_3_2 u_ca_3_2_724(.d_in(u_ca_in_724), .d_out(u_ca_out_724));
compressor_3_2 u_ca_3_2_725(.d_in(u_ca_in_725), .d_out(u_ca_out_725));
compressor_3_2 u_ca_3_2_726(.d_in(u_ca_in_726), .d_out(u_ca_out_726));
compressor_3_2 u_ca_3_2_727(.d_in(u_ca_in_727), .d_out(u_ca_out_727));
compressor_3_2 u_ca_3_2_728(.d_in(u_ca_in_728), .d_out(u_ca_out_728));
compressor_3_2 u_ca_3_2_729(.d_in(u_ca_in_729), .d_out(u_ca_out_729));
compressor_3_2 u_ca_3_2_730(.d_in(u_ca_in_730), .d_out(u_ca_out_730));
compressor_3_2 u_ca_3_2_731(.d_in(u_ca_in_731), .d_out(u_ca_out_731));
compressor_3_2 u_ca_3_2_732(.d_in(u_ca_in_732), .d_out(u_ca_out_732));
compressor_3_2 u_ca_3_2_733(.d_in(u_ca_in_733), .d_out(u_ca_out_733));
compressor_3_2 u_ca_3_2_734(.d_in(u_ca_in_734), .d_out(u_ca_out_734));
compressor_3_2 u_ca_3_2_735(.d_in(u_ca_in_735), .d_out(u_ca_out_735));
compressor_3_2 u_ca_3_2_736(.d_in(u_ca_in_736), .d_out(u_ca_out_736));
compressor_3_2 u_ca_3_2_737(.d_in(u_ca_in_737), .d_out(u_ca_out_737));
compressor_3_2 u_ca_3_2_738(.d_in(u_ca_in_738), .d_out(u_ca_out_738));
compressor_3_2 u_ca_3_2_739(.d_in(u_ca_in_739), .d_out(u_ca_out_739));
compressor_3_2 u_ca_3_2_740(.d_in(u_ca_in_740), .d_out(u_ca_out_740));
compressor_3_2 u_ca_3_2_741(.d_in(u_ca_in_741), .d_out(u_ca_out_741));
compressor_3_2 u_ca_3_2_742(.d_in(u_ca_in_742), .d_out(u_ca_out_742));
compressor_3_2 u_ca_3_2_743(.d_in(u_ca_in_743), .d_out(u_ca_out_743));
compressor_3_2 u_ca_3_2_744(.d_in(u_ca_in_744), .d_out(u_ca_out_744));
compressor_3_2 u_ca_3_2_745(.d_in(u_ca_in_745), .d_out(u_ca_out_745));
compressor_3_2 u_ca_3_2_746(.d_in(u_ca_in_746), .d_out(u_ca_out_746));
compressor_3_2 u_ca_3_2_747(.d_in(u_ca_in_747), .d_out(u_ca_out_747));
compressor_3_2 u_ca_3_2_748(.d_in(u_ca_in_748), .d_out(u_ca_out_748));
compressor_3_2 u_ca_3_2_749(.d_in(u_ca_in_749), .d_out(u_ca_out_749));
compressor_3_2 u_ca_3_2_750(.d_in(u_ca_in_750), .d_out(u_ca_out_750));
compressor_3_2 u_ca_3_2_751(.d_in(u_ca_in_751), .d_out(u_ca_out_751));
compressor_3_2 u_ca_3_2_752(.d_in(u_ca_in_752), .d_out(u_ca_out_752));
compressor_3_2 u_ca_3_2_753(.d_in(u_ca_in_753), .d_out(u_ca_out_753));
compressor_3_2 u_ca_3_2_754(.d_in(u_ca_in_754), .d_out(u_ca_out_754));
compressor_3_2 u_ca_3_2_755(.d_in(u_ca_in_755), .d_out(u_ca_out_755));
compressor_3_2 u_ca_3_2_756(.d_in(u_ca_in_756), .d_out(u_ca_out_756));
compressor_3_2 u_ca_3_2_757(.d_in(u_ca_in_757), .d_out(u_ca_out_757));
compressor_3_2 u_ca_3_2_758(.d_in(u_ca_in_758), .d_out(u_ca_out_758));
compressor_3_2 u_ca_3_2_759(.d_in(u_ca_in_759), .d_out(u_ca_out_759));
compressor_3_2 u_ca_3_2_760(.d_in(u_ca_in_760), .d_out(u_ca_out_760));
compressor_3_2 u_ca_3_2_761(.d_in(u_ca_in_761), .d_out(u_ca_out_761));
compressor_3_2 u_ca_3_2_762(.d_in(u_ca_in_762), .d_out(u_ca_out_762));
compressor_3_2 u_ca_3_2_763(.d_in(u_ca_in_763), .d_out(u_ca_out_763));
compressor_3_2 u_ca_3_2_764(.d_in(u_ca_in_764), .d_out(u_ca_out_764));
compressor_3_2 u_ca_3_2_765(.d_in(u_ca_in_765), .d_out(u_ca_out_765));
compressor_3_2 u_ca_3_2_766(.d_in(u_ca_in_766), .d_out(u_ca_out_766));
compressor_3_2 u_ca_3_2_767(.d_in(u_ca_in_767), .d_out(u_ca_out_767));
compressor_3_2 u_ca_3_2_768(.d_in(u_ca_in_768), .d_out(u_ca_out_768));
compressor_3_2 u_ca_3_2_769(.d_in(u_ca_in_769), .d_out(u_ca_out_769));
compressor_3_2 u_ca_3_2_770(.d_in(u_ca_in_770), .d_out(u_ca_out_770));
compressor_3_2 u_ca_3_2_771(.d_in(u_ca_in_771), .d_out(u_ca_out_771));
compressor_3_2 u_ca_3_2_772(.d_in(u_ca_in_772), .d_out(u_ca_out_772));
compressor_3_2 u_ca_3_2_773(.d_in(u_ca_in_773), .d_out(u_ca_out_773));
compressor_3_2 u_ca_3_2_774(.d_in(u_ca_in_774), .d_out(u_ca_out_774));
compressor_3_2 u_ca_3_2_775(.d_in(u_ca_in_775), .d_out(u_ca_out_775));
compressor_3_2 u_ca_3_2_776(.d_in(u_ca_in_776), .d_out(u_ca_out_776));
compressor_3_2 u_ca_3_2_777(.d_in(u_ca_in_777), .d_out(u_ca_out_777));
compressor_3_2 u_ca_3_2_778(.d_in(u_ca_in_778), .d_out(u_ca_out_778));
compressor_3_2 u_ca_3_2_779(.d_in(u_ca_in_779), .d_out(u_ca_out_779));
compressor_3_2 u_ca_3_2_780(.d_in(u_ca_in_780), .d_out(u_ca_out_780));
compressor_3_2 u_ca_3_2_781(.d_in(u_ca_in_781), .d_out(u_ca_out_781));
compressor_3_2 u_ca_3_2_782(.d_in(u_ca_in_782), .d_out(u_ca_out_782));
compressor_3_2 u_ca_3_2_783(.d_in(u_ca_in_783), .d_out(u_ca_out_783));
compressor_3_2 u_ca_3_2_784(.d_in(u_ca_in_784), .d_out(u_ca_out_784));
compressor_3_2 u_ca_3_2_785(.d_in(u_ca_in_785), .d_out(u_ca_out_785));
compressor_3_2 u_ca_3_2_786(.d_in(u_ca_in_786), .d_out(u_ca_out_786));
compressor_3_2 u_ca_3_2_787(.d_in(u_ca_in_787), .d_out(u_ca_out_787));
compressor_3_2 u_ca_3_2_788(.d_in(u_ca_in_788), .d_out(u_ca_out_788));
compressor_3_2 u_ca_3_2_789(.d_in(u_ca_in_789), .d_out(u_ca_out_789));
compressor_3_2 u_ca_3_2_790(.d_in(u_ca_in_790), .d_out(u_ca_out_790));
compressor_3_2 u_ca_3_2_791(.d_in(u_ca_in_791), .d_out(u_ca_out_791));
compressor_3_2 u_ca_3_2_792(.d_in(u_ca_in_792), .d_out(u_ca_out_792));
compressor_3_2 u_ca_3_2_793(.d_in(u_ca_in_793), .d_out(u_ca_out_793));
compressor_3_2 u_ca_3_2_794(.d_in(u_ca_in_794), .d_out(u_ca_out_794));
compressor_3_2 u_ca_3_2_795(.d_in(u_ca_in_795), .d_out(u_ca_out_795));
compressor_3_2 u_ca_3_2_796(.d_in(u_ca_in_796), .d_out(u_ca_out_796));
compressor_3_2 u_ca_3_2_797(.d_in(u_ca_in_797), .d_out(u_ca_out_797));
compressor_3_2 u_ca_3_2_798(.d_in(u_ca_in_798), .d_out(u_ca_out_798));
compressor_3_2 u_ca_3_2_799(.d_in(u_ca_in_799), .d_out(u_ca_out_799));
compressor_3_2 u_ca_3_2_800(.d_in(u_ca_in_800), .d_out(u_ca_out_800));
compressor_3_2 u_ca_3_2_801(.d_in(u_ca_in_801), .d_out(u_ca_out_801));
compressor_3_2 u_ca_3_2_802(.d_in(u_ca_in_802), .d_out(u_ca_out_802));
compressor_3_2 u_ca_3_2_803(.d_in(u_ca_in_803), .d_out(u_ca_out_803));
compressor_3_2 u_ca_3_2_804(.d_in(u_ca_in_804), .d_out(u_ca_out_804));
compressor_3_2 u_ca_3_2_805(.d_in(u_ca_in_805), .d_out(u_ca_out_805));
compressor_3_2 u_ca_3_2_806(.d_in(u_ca_in_806), .d_out(u_ca_out_806));
compressor_3_2 u_ca_3_2_807(.d_in(u_ca_in_807), .d_out(u_ca_out_807));
compressor_3_2 u_ca_3_2_808(.d_in(u_ca_in_808), .d_out(u_ca_out_808));
compressor_3_2 u_ca_3_2_809(.d_in(u_ca_in_809), .d_out(u_ca_out_809));
compressor_3_2 u_ca_3_2_810(.d_in(u_ca_in_810), .d_out(u_ca_out_810));
compressor_3_2 u_ca_3_2_811(.d_in(u_ca_in_811), .d_out(u_ca_out_811));
compressor_3_2 u_ca_3_2_812(.d_in(u_ca_in_812), .d_out(u_ca_out_812));
compressor_3_2 u_ca_3_2_813(.d_in(u_ca_in_813), .d_out(u_ca_out_813));
compressor_3_2 u_ca_3_2_814(.d_in(u_ca_in_814), .d_out(u_ca_out_814));
compressor_3_2 u_ca_3_2_815(.d_in(u_ca_in_815), .d_out(u_ca_out_815));
compressor_3_2 u_ca_3_2_816(.d_in(u_ca_in_816), .d_out(u_ca_out_816));
compressor_3_2 u_ca_3_2_817(.d_in(u_ca_in_817), .d_out(u_ca_out_817));
compressor_3_2 u_ca_3_2_818(.d_in(u_ca_in_818), .d_out(u_ca_out_818));
compressor_3_2 u_ca_3_2_819(.d_in(u_ca_in_819), .d_out(u_ca_out_819));
compressor_3_2 u_ca_3_2_820(.d_in(u_ca_in_820), .d_out(u_ca_out_820));
compressor_3_2 u_ca_3_2_821(.d_in(u_ca_in_821), .d_out(u_ca_out_821));
compressor_3_2 u_ca_3_2_822(.d_in(u_ca_in_822), .d_out(u_ca_out_822));
compressor_3_2 u_ca_3_2_823(.d_in(u_ca_in_823), .d_out(u_ca_out_823));
compressor_3_2 u_ca_3_2_824(.d_in(u_ca_in_824), .d_out(u_ca_out_824));
compressor_3_2 u_ca_3_2_825(.d_in(u_ca_in_825), .d_out(u_ca_out_825));
compressor_3_2 u_ca_3_2_826(.d_in(u_ca_in_826), .d_out(u_ca_out_826));
compressor_3_2 u_ca_3_2_827(.d_in(u_ca_in_827), .d_out(u_ca_out_827));
compressor_3_2 u_ca_3_2_828(.d_in(u_ca_in_828), .d_out(u_ca_out_828));
compressor_3_2 u_ca_3_2_829(.d_in(u_ca_in_829), .d_out(u_ca_out_829));
compressor_3_2 u_ca_3_2_830(.d_in(u_ca_in_830), .d_out(u_ca_out_830));
compressor_3_2 u_ca_3_2_831(.d_in(u_ca_in_831), .d_out(u_ca_out_831));
compressor_3_2 u_ca_3_2_832(.d_in(u_ca_in_832), .d_out(u_ca_out_832));
compressor_3_2 u_ca_3_2_833(.d_in(u_ca_in_833), .d_out(u_ca_out_833));
compressor_3_2 u_ca_3_2_834(.d_in(u_ca_in_834), .d_out(u_ca_out_834));
compressor_3_2 u_ca_3_2_835(.d_in(u_ca_in_835), .d_out(u_ca_out_835));
compressor_3_2 u_ca_3_2_836(.d_in(u_ca_in_836), .d_out(u_ca_out_836));
compressor_3_2 u_ca_3_2_837(.d_in(u_ca_in_837), .d_out(u_ca_out_837));
compressor_3_2 u_ca_3_2_838(.d_in(u_ca_in_838), .d_out(u_ca_out_838));
compressor_3_2 u_ca_3_2_839(.d_in(u_ca_in_839), .d_out(u_ca_out_839));
compressor_3_2 u_ca_3_2_840(.d_in(u_ca_in_840), .d_out(u_ca_out_840));
compressor_3_2 u_ca_3_2_841(.d_in(u_ca_in_841), .d_out(u_ca_out_841));
compressor_3_2 u_ca_3_2_842(.d_in(u_ca_in_842), .d_out(u_ca_out_842));
compressor_3_2 u_ca_3_2_843(.d_in(u_ca_in_843), .d_out(u_ca_out_843));
compressor_3_2 u_ca_3_2_844(.d_in(u_ca_in_844), .d_out(u_ca_out_844));
compressor_3_2 u_ca_3_2_845(.d_in(u_ca_in_845), .d_out(u_ca_out_845));
compressor_3_2 u_ca_3_2_846(.d_in(u_ca_in_846), .d_out(u_ca_out_846));
compressor_3_2 u_ca_3_2_847(.d_in(u_ca_in_847), .d_out(u_ca_out_847));
compressor_3_2 u_ca_3_2_848(.d_in(u_ca_in_848), .d_out(u_ca_out_848));
compressor_3_2 u_ca_3_2_849(.d_in(u_ca_in_849), .d_out(u_ca_out_849));
compressor_3_2 u_ca_3_2_850(.d_in(u_ca_in_850), .d_out(u_ca_out_850));
compressor_3_2 u_ca_3_2_851(.d_in(u_ca_in_851), .d_out(u_ca_out_851));
compressor_3_2 u_ca_3_2_852(.d_in(u_ca_in_852), .d_out(u_ca_out_852));
compressor_3_2 u_ca_3_2_853(.d_in(u_ca_in_853), .d_out(u_ca_out_853));
compressor_3_2 u_ca_3_2_854(.d_in(u_ca_in_854), .d_out(u_ca_out_854));
compressor_3_2 u_ca_3_2_855(.d_in(u_ca_in_855), .d_out(u_ca_out_855));
compressor_3_2 u_ca_3_2_856(.d_in(u_ca_in_856), .d_out(u_ca_out_856));
compressor_3_2 u_ca_3_2_857(.d_in(u_ca_in_857), .d_out(u_ca_out_857));
compressor_3_2 u_ca_3_2_858(.d_in(u_ca_in_858), .d_out(u_ca_out_858));
compressor_3_2 u_ca_3_2_859(.d_in(u_ca_in_859), .d_out(u_ca_out_859));
compressor_3_2 u_ca_3_2_860(.d_in(u_ca_in_860), .d_out(u_ca_out_860));
compressor_3_2 u_ca_3_2_861(.d_in(u_ca_in_861), .d_out(u_ca_out_861));
compressor_3_2 u_ca_3_2_862(.d_in(u_ca_in_862), .d_out(u_ca_out_862));
compressor_3_2 u_ca_3_2_863(.d_in(u_ca_in_863), .d_out(u_ca_out_863));
compressor_3_2 u_ca_3_2_864(.d_in(u_ca_in_864), .d_out(u_ca_out_864));
compressor_3_2 u_ca_3_2_865(.d_in(u_ca_in_865), .d_out(u_ca_out_865));
compressor_3_2 u_ca_3_2_866(.d_in(u_ca_in_866), .d_out(u_ca_out_866));
compressor_3_2 u_ca_3_2_867(.d_in(u_ca_in_867), .d_out(u_ca_out_867));
compressor_3_2 u_ca_3_2_868(.d_in(u_ca_in_868), .d_out(u_ca_out_868));
compressor_3_2 u_ca_3_2_869(.d_in(u_ca_in_869), .d_out(u_ca_out_869));
compressor_3_2 u_ca_3_2_870(.d_in(u_ca_in_870), .d_out(u_ca_out_870));
compressor_3_2 u_ca_3_2_871(.d_in(u_ca_in_871), .d_out(u_ca_out_871));
compressor_3_2 u_ca_3_2_872(.d_in(u_ca_in_872), .d_out(u_ca_out_872));
compressor_3_2 u_ca_3_2_873(.d_in(u_ca_in_873), .d_out(u_ca_out_873));
compressor_3_2 u_ca_3_2_874(.d_in(u_ca_in_874), .d_out(u_ca_out_874));
compressor_3_2 u_ca_3_2_875(.d_in(u_ca_in_875), .d_out(u_ca_out_875));
compressor_3_2 u_ca_3_2_876(.d_in(u_ca_in_876), .d_out(u_ca_out_876));
compressor_3_2 u_ca_3_2_877(.d_in(u_ca_in_877), .d_out(u_ca_out_877));
compressor_3_2 u_ca_3_2_878(.d_in(u_ca_in_878), .d_out(u_ca_out_878));
compressor_3_2 u_ca_3_2_879(.d_in(u_ca_in_879), .d_out(u_ca_out_879));
compressor_3_2 u_ca_3_2_880(.d_in(u_ca_in_880), .d_out(u_ca_out_880));
compressor_3_2 u_ca_3_2_881(.d_in(u_ca_in_881), .d_out(u_ca_out_881));
compressor_3_2 u_ca_3_2_882(.d_in(u_ca_in_882), .d_out(u_ca_out_882));
compressor_3_2 u_ca_3_2_883(.d_in(u_ca_in_883), .d_out(u_ca_out_883));
compressor_3_2 u_ca_3_2_884(.d_in(u_ca_in_884), .d_out(u_ca_out_884));
compressor_3_2 u_ca_3_2_885(.d_in(u_ca_in_885), .d_out(u_ca_out_885));
compressor_3_2 u_ca_3_2_886(.d_in(u_ca_in_886), .d_out(u_ca_out_886));
compressor_3_2 u_ca_3_2_887(.d_in(u_ca_in_887), .d_out(u_ca_out_887));
compressor_3_2 u_ca_3_2_888(.d_in(u_ca_in_888), .d_out(u_ca_out_888));
compressor_3_2 u_ca_3_2_889(.d_in(u_ca_in_889), .d_out(u_ca_out_889));
compressor_3_2 u_ca_3_2_890(.d_in(u_ca_in_890), .d_out(u_ca_out_890));
compressor_3_2 u_ca_3_2_891(.d_in(u_ca_in_891), .d_out(u_ca_out_891));
compressor_3_2 u_ca_3_2_892(.d_in(u_ca_in_892), .d_out(u_ca_out_892));
compressor_3_2 u_ca_3_2_893(.d_in(u_ca_in_893), .d_out(u_ca_out_893));
compressor_3_2 u_ca_3_2_894(.d_in(u_ca_in_894), .d_out(u_ca_out_894));
compressor_3_2 u_ca_3_2_895(.d_in(u_ca_in_895), .d_out(u_ca_out_895));
compressor_3_2 u_ca_3_2_896(.d_in(u_ca_in_896), .d_out(u_ca_out_896));
compressor_3_2 u_ca_3_2_897(.d_in(u_ca_in_897), .d_out(u_ca_out_897));
compressor_3_2 u_ca_3_2_898(.d_in(u_ca_in_898), .d_out(u_ca_out_898));
compressor_3_2 u_ca_3_2_899(.d_in(u_ca_in_899), .d_out(u_ca_out_899));
compressor_3_2 u_ca_3_2_900(.d_in(u_ca_in_900), .d_out(u_ca_out_900));
compressor_3_2 u_ca_3_2_901(.d_in(u_ca_in_901), .d_out(u_ca_out_901));
compressor_3_2 u_ca_3_2_902(.d_in(u_ca_in_902), .d_out(u_ca_out_902));
compressor_3_2 u_ca_3_2_903(.d_in(u_ca_in_903), .d_out(u_ca_out_903));
compressor_3_2 u_ca_3_2_904(.d_in(u_ca_in_904), .d_out(u_ca_out_904));
compressor_3_2 u_ca_3_2_905(.d_in(u_ca_in_905), .d_out(u_ca_out_905));
compressor_3_2 u_ca_3_2_906(.d_in(u_ca_in_906), .d_out(u_ca_out_906));
compressor_3_2 u_ca_3_2_907(.d_in(u_ca_in_907), .d_out(u_ca_out_907));
compressor_3_2 u_ca_3_2_908(.d_in(u_ca_in_908), .d_out(u_ca_out_908));
compressor_3_2 u_ca_3_2_909(.d_in(u_ca_in_909), .d_out(u_ca_out_909));
compressor_3_2 u_ca_3_2_910(.d_in(u_ca_in_910), .d_out(u_ca_out_910));
compressor_3_2 u_ca_3_2_911(.d_in(u_ca_in_911), .d_out(u_ca_out_911));
compressor_3_2 u_ca_3_2_912(.d_in(u_ca_in_912), .d_out(u_ca_out_912));
compressor_3_2 u_ca_3_2_913(.d_in(u_ca_in_913), .d_out(u_ca_out_913));
compressor_3_2 u_ca_3_2_914(.d_in(u_ca_in_914), .d_out(u_ca_out_914));
compressor_3_2 u_ca_3_2_915(.d_in(u_ca_in_915), .d_out(u_ca_out_915));
compressor_3_2 u_ca_3_2_916(.d_in(u_ca_in_916), .d_out(u_ca_out_916));
compressor_3_2 u_ca_3_2_917(.d_in(u_ca_in_917), .d_out(u_ca_out_917));
compressor_3_2 u_ca_3_2_918(.d_in(u_ca_in_918), .d_out(u_ca_out_918));
compressor_3_2 u_ca_3_2_919(.d_in(u_ca_in_919), .d_out(u_ca_out_919));
compressor_3_2 u_ca_3_2_920(.d_in(u_ca_in_920), .d_out(u_ca_out_920));
compressor_3_2 u_ca_3_2_921(.d_in(u_ca_in_921), .d_out(u_ca_out_921));
compressor_3_2 u_ca_3_2_922(.d_in(u_ca_in_922), .d_out(u_ca_out_922));
compressor_3_2 u_ca_3_2_923(.d_in(u_ca_in_923), .d_out(u_ca_out_923));
compressor_3_2 u_ca_3_2_924(.d_in(u_ca_in_924), .d_out(u_ca_out_924));
compressor_3_2 u_ca_3_2_925(.d_in(u_ca_in_925), .d_out(u_ca_out_925));
compressor_3_2 u_ca_3_2_926(.d_in(u_ca_in_926), .d_out(u_ca_out_926));
compressor_3_2 u_ca_3_2_927(.d_in(u_ca_in_927), .d_out(u_ca_out_927));
compressor_3_2 u_ca_3_2_928(.d_in(u_ca_in_928), .d_out(u_ca_out_928));
compressor_3_2 u_ca_3_2_929(.d_in(u_ca_in_929), .d_out(u_ca_out_929));
compressor_3_2 u_ca_3_2_930(.d_in(u_ca_in_930), .d_out(u_ca_out_930));
compressor_3_2 u_ca_3_2_931(.d_in(u_ca_in_931), .d_out(u_ca_out_931));
compressor_3_2 u_ca_3_2_932(.d_in(u_ca_in_932), .d_out(u_ca_out_932));
compressor_3_2 u_ca_3_2_933(.d_in(u_ca_in_933), .d_out(u_ca_out_933));
compressor_3_2 u_ca_3_2_934(.d_in(u_ca_in_934), .d_out(u_ca_out_934));
compressor_3_2 u_ca_3_2_935(.d_in(u_ca_in_935), .d_out(u_ca_out_935));
compressor_3_2 u_ca_3_2_936(.d_in(u_ca_in_936), .d_out(u_ca_out_936));
compressor_3_2 u_ca_3_2_937(.d_in(u_ca_in_937), .d_out(u_ca_out_937));
compressor_3_2 u_ca_3_2_938(.d_in(u_ca_in_938), .d_out(u_ca_out_938));
compressor_3_2 u_ca_3_2_939(.d_in(u_ca_in_939), .d_out(u_ca_out_939));
compressor_3_2 u_ca_3_2_940(.d_in(u_ca_in_940), .d_out(u_ca_out_940));
compressor_3_2 u_ca_3_2_941(.d_in(u_ca_in_941), .d_out(u_ca_out_941));
compressor_3_2 u_ca_3_2_942(.d_in(u_ca_in_942), .d_out(u_ca_out_942));
compressor_3_2 u_ca_3_2_943(.d_in(u_ca_in_943), .d_out(u_ca_out_943));
compressor_3_2 u_ca_3_2_944(.d_in(u_ca_in_944), .d_out(u_ca_out_944));
compressor_3_2 u_ca_3_2_945(.d_in(u_ca_in_945), .d_out(u_ca_out_945));
compressor_3_2 u_ca_3_2_946(.d_in(u_ca_in_946), .d_out(u_ca_out_946));
compressor_3_2 u_ca_3_2_947(.d_in(u_ca_in_947), .d_out(u_ca_out_947));
compressor_3_2 u_ca_3_2_948(.d_in(u_ca_in_948), .d_out(u_ca_out_948));
compressor_3_2 u_ca_3_2_949(.d_in(u_ca_in_949), .d_out(u_ca_out_949));
compressor_3_2 u_ca_3_2_950(.d_in(u_ca_in_950), .d_out(u_ca_out_950));
compressor_3_2 u_ca_3_2_951(.d_in(u_ca_in_951), .d_out(u_ca_out_951));
compressor_3_2 u_ca_3_2_952(.d_in(u_ca_in_952), .d_out(u_ca_out_952));
compressor_3_2 u_ca_3_2_953(.d_in(u_ca_in_953), .d_out(u_ca_out_953));
compressor_3_2 u_ca_3_2_954(.d_in(u_ca_in_954), .d_out(u_ca_out_954));
compressor_3_2 u_ca_3_2_955(.d_in(u_ca_in_955), .d_out(u_ca_out_955));
compressor_3_2 u_ca_3_2_956(.d_in(u_ca_in_956), .d_out(u_ca_out_956));
compressor_3_2 u_ca_3_2_957(.d_in(u_ca_in_957), .d_out(u_ca_out_957));
compressor_3_2 u_ca_3_2_958(.d_in(u_ca_in_958), .d_out(u_ca_out_958));
compressor_3_2 u_ca_3_2_959(.d_in(u_ca_in_959), .d_out(u_ca_out_959));
compressor_3_2 u_ca_3_2_960(.d_in(u_ca_in_960), .d_out(u_ca_out_960));
compressor_3_2 u_ca_3_2_961(.d_in(u_ca_in_961), .d_out(u_ca_out_961));
compressor_3_2 u_ca_3_2_962(.d_in(u_ca_in_962), .d_out(u_ca_out_962));
compressor_3_2 u_ca_3_2_963(.d_in(u_ca_in_963), .d_out(u_ca_out_963));
compressor_3_2 u_ca_3_2_964(.d_in(u_ca_in_964), .d_out(u_ca_out_964));
compressor_3_2 u_ca_3_2_965(.d_in(u_ca_in_965), .d_out(u_ca_out_965));
compressor_3_2 u_ca_3_2_966(.d_in(u_ca_in_966), .d_out(u_ca_out_966));
compressor_3_2 u_ca_3_2_967(.d_in(u_ca_in_967), .d_out(u_ca_out_967));
compressor_3_2 u_ca_3_2_968(.d_in(u_ca_in_968), .d_out(u_ca_out_968));
compressor_3_2 u_ca_3_2_969(.d_in(u_ca_in_969), .d_out(u_ca_out_969));
compressor_3_2 u_ca_3_2_970(.d_in(u_ca_in_970), .d_out(u_ca_out_970));
compressor_3_2 u_ca_3_2_971(.d_in(u_ca_in_971), .d_out(u_ca_out_971));
compressor_3_2 u_ca_3_2_972(.d_in(u_ca_in_972), .d_out(u_ca_out_972));
compressor_3_2 u_ca_3_2_973(.d_in(u_ca_in_973), .d_out(u_ca_out_973));
compressor_3_2 u_ca_3_2_974(.d_in(u_ca_in_974), .d_out(u_ca_out_974));
compressor_3_2 u_ca_3_2_975(.d_in(u_ca_in_975), .d_out(u_ca_out_975));
compressor_3_2 u_ca_3_2_976(.d_in(u_ca_in_976), .d_out(u_ca_out_976));
compressor_3_2 u_ca_3_2_977(.d_in(u_ca_in_977), .d_out(u_ca_out_977));
compressor_3_2 u_ca_3_2_978(.d_in(u_ca_in_978), .d_out(u_ca_out_978));
compressor_3_2 u_ca_3_2_979(.d_in(u_ca_in_979), .d_out(u_ca_out_979));
compressor_3_2 u_ca_3_2_980(.d_in(u_ca_in_980), .d_out(u_ca_out_980));
compressor_3_2 u_ca_3_2_981(.d_in(u_ca_in_981), .d_out(u_ca_out_981));
compressor_3_2 u_ca_3_2_982(.d_in(u_ca_in_982), .d_out(u_ca_out_982));
compressor_3_2 u_ca_3_2_983(.d_in(u_ca_in_983), .d_out(u_ca_out_983));
compressor_3_2 u_ca_3_2_984(.d_in(u_ca_in_984), .d_out(u_ca_out_984));
compressor_3_2 u_ca_3_2_985(.d_in(u_ca_in_985), .d_out(u_ca_out_985));
compressor_3_2 u_ca_3_2_986(.d_in(u_ca_in_986), .d_out(u_ca_out_986));
compressor_3_2 u_ca_3_2_987(.d_in(u_ca_in_987), .d_out(u_ca_out_987));
compressor_3_2 u_ca_3_2_988(.d_in(u_ca_in_988), .d_out(u_ca_out_988));
compressor_3_2 u_ca_3_2_989(.d_in(u_ca_in_989), .d_out(u_ca_out_989));
compressor_3_2 u_ca_3_2_990(.d_in(u_ca_in_990), .d_out(u_ca_out_990));
compressor_3_2 u_ca_3_2_991(.d_in(u_ca_in_991), .d_out(u_ca_out_991));
compressor_3_2 u_ca_3_2_992(.d_in(u_ca_in_992), .d_out(u_ca_out_992));
compressor_3_2 u_ca_3_2_993(.d_in(u_ca_in_993), .d_out(u_ca_out_993));
compressor_3_2 u_ca_3_2_994(.d_in(u_ca_in_994), .d_out(u_ca_out_994));
compressor_3_2 u_ca_3_2_995(.d_in(u_ca_in_995), .d_out(u_ca_out_995));
compressor_3_2 u_ca_3_2_996(.d_in(u_ca_in_996), .d_out(u_ca_out_996));
compressor_3_2 u_ca_3_2_997(.d_in(u_ca_in_997), .d_out(u_ca_out_997));
compressor_3_2 u_ca_3_2_998(.d_in(u_ca_in_998), .d_out(u_ca_out_998));
compressor_3_2 u_ca_3_2_999(.d_in(u_ca_in_999), .d_out(u_ca_out_999));
compressor_3_2 u_ca_3_2_1000(.d_in(u_ca_in_1000), .d_out(u_ca_out_1000));
compressor_3_2 u_ca_3_2_1001(.d_in(u_ca_in_1001), .d_out(u_ca_out_1001));
compressor_3_2 u_ca_3_2_1002(.d_in(u_ca_in_1002), .d_out(u_ca_out_1002));
compressor_3_2 u_ca_3_2_1003(.d_in(u_ca_in_1003), .d_out(u_ca_out_1003));
compressor_3_2 u_ca_3_2_1004(.d_in(u_ca_in_1004), .d_out(u_ca_out_1004));
compressor_3_2 u_ca_3_2_1005(.d_in(u_ca_in_1005), .d_out(u_ca_out_1005));
compressor_3_2 u_ca_3_2_1006(.d_in(u_ca_in_1006), .d_out(u_ca_out_1006));
compressor_3_2 u_ca_3_2_1007(.d_in(u_ca_in_1007), .d_out(u_ca_out_1007));
compressor_3_2 u_ca_3_2_1008(.d_in(u_ca_in_1008), .d_out(u_ca_out_1008));
compressor_3_2 u_ca_3_2_1009(.d_in(u_ca_in_1009), .d_out(u_ca_out_1009));
compressor_3_2 u_ca_3_2_1010(.d_in(u_ca_in_1010), .d_out(u_ca_out_1010));
compressor_3_2 u_ca_3_2_1011(.d_in(u_ca_in_1011), .d_out(u_ca_out_1011));
compressor_3_2 u_ca_3_2_1012(.d_in(u_ca_in_1012), .d_out(u_ca_out_1012));
compressor_3_2 u_ca_3_2_1013(.d_in(u_ca_in_1013), .d_out(u_ca_out_1013));
compressor_3_2 u_ca_3_2_1014(.d_in(u_ca_in_1014), .d_out(u_ca_out_1014));
compressor_3_2 u_ca_3_2_1015(.d_in(u_ca_in_1015), .d_out(u_ca_out_1015));
compressor_3_2 u_ca_3_2_1016(.d_in(u_ca_in_1016), .d_out(u_ca_out_1016));
compressor_3_2 u_ca_3_2_1017(.d_in(u_ca_in_1017), .d_out(u_ca_out_1017));
compressor_3_2 u_ca_3_2_1018(.d_in(u_ca_in_1018), .d_out(u_ca_out_1018));
compressor_3_2 u_ca_3_2_1019(.d_in(u_ca_in_1019), .d_out(u_ca_out_1019));
compressor_3_2 u_ca_3_2_1020(.d_in(u_ca_in_1020), .d_out(u_ca_out_1020));
compressor_3_2 u_ca_3_2_1021(.d_in(u_ca_in_1021), .d_out(u_ca_out_1021));
compressor_3_2 u_ca_3_2_1022(.d_in(u_ca_in_1022), .d_out(u_ca_out_1022));
compressor_3_2 u_ca_3_2_1023(.d_in(u_ca_in_1023), .d_out(u_ca_out_1023));

//---------------------------------------------------------



//--output-------------------------------------------------

assign col_out_0 = {{1{1'b0}}, u_ca_out_0[0:0]};
assign col_out_1 = {u_ca_out_1[0:0], u_ca_out_0[1:1]};
assign col_out_2 = {u_ca_out_2[0:0], u_ca_out_1[1:1]};
assign col_out_3 = {u_ca_out_3[0:0], u_ca_out_2[1:1]};
assign col_out_4 = {u_ca_out_4[0:0], u_ca_out_3[1:1]};
assign col_out_5 = {u_ca_out_5[0:0], u_ca_out_4[1:1]};
assign col_out_6 = {u_ca_out_6[0:0], u_ca_out_5[1:1]};
assign col_out_7 = {u_ca_out_7[0:0], u_ca_out_6[1:1]};
assign col_out_8 = {u_ca_out_8[0:0], u_ca_out_7[1:1]};
assign col_out_9 = {u_ca_out_9[0:0], u_ca_out_8[1:1]};
assign col_out_10 = {u_ca_out_10[0:0], u_ca_out_9[1:1]};
assign col_out_11 = {u_ca_out_11[0:0], u_ca_out_10[1:1]};
assign col_out_12 = {u_ca_out_12[0:0], u_ca_out_11[1:1]};
assign col_out_13 = {u_ca_out_13[0:0], u_ca_out_12[1:1]};
assign col_out_14 = {u_ca_out_14[0:0], u_ca_out_13[1:1]};
assign col_out_15 = {u_ca_out_15[0:0], u_ca_out_14[1:1]};
assign col_out_16 = {u_ca_out_16[0:0], u_ca_out_15[1:1]};
assign col_out_17 = {u_ca_out_17[0:0], u_ca_out_16[1:1]};
assign col_out_18 = {u_ca_out_18[0:0], u_ca_out_17[1:1]};
assign col_out_19 = {u_ca_out_19[0:0], u_ca_out_18[1:1]};
assign col_out_20 = {u_ca_out_20[0:0], u_ca_out_19[1:1]};
assign col_out_21 = {u_ca_out_21[0:0], u_ca_out_20[1:1]};
assign col_out_22 = {u_ca_out_22[0:0], u_ca_out_21[1:1]};
assign col_out_23 = {u_ca_out_23[0:0], u_ca_out_22[1:1]};
assign col_out_24 = {u_ca_out_24[0:0], u_ca_out_23[1:1]};
assign col_out_25 = {u_ca_out_25[0:0], u_ca_out_24[1:1]};
assign col_out_26 = {u_ca_out_26[0:0], u_ca_out_25[1:1]};
assign col_out_27 = {u_ca_out_27[0:0], u_ca_out_26[1:1]};
assign col_out_28 = {u_ca_out_28[0:0], u_ca_out_27[1:1]};
assign col_out_29 = {u_ca_out_29[0:0], u_ca_out_28[1:1]};
assign col_out_30 = {u_ca_out_30[0:0], u_ca_out_29[1:1]};
assign col_out_31 = {u_ca_out_31[0:0], u_ca_out_30[1:1]};
assign col_out_32 = {u_ca_out_32[0:0], u_ca_out_31[1:1]};
assign col_out_33 = {u_ca_out_33[0:0], u_ca_out_32[1:1]};
assign col_out_34 = {u_ca_out_34[0:0], u_ca_out_33[1:1]};
assign col_out_35 = {u_ca_out_35[0:0], u_ca_out_34[1:1]};
assign col_out_36 = {u_ca_out_36[0:0], u_ca_out_35[1:1]};
assign col_out_37 = {u_ca_out_37[0:0], u_ca_out_36[1:1]};
assign col_out_38 = {u_ca_out_38[0:0], u_ca_out_37[1:1]};
assign col_out_39 = {u_ca_out_39[0:0], u_ca_out_38[1:1]};
assign col_out_40 = {u_ca_out_40[0:0], u_ca_out_39[1:1]};
assign col_out_41 = {u_ca_out_41[0:0], u_ca_out_40[1:1]};
assign col_out_42 = {u_ca_out_42[0:0], u_ca_out_41[1:1]};
assign col_out_43 = {u_ca_out_43[0:0], u_ca_out_42[1:1]};
assign col_out_44 = {u_ca_out_44[0:0], u_ca_out_43[1:1]};
assign col_out_45 = {u_ca_out_45[0:0], u_ca_out_44[1:1]};
assign col_out_46 = {u_ca_out_46[0:0], u_ca_out_45[1:1]};
assign col_out_47 = {u_ca_out_47[0:0], u_ca_out_46[1:1]};
assign col_out_48 = {u_ca_out_48[0:0], u_ca_out_47[1:1]};
assign col_out_49 = {u_ca_out_49[0:0], u_ca_out_48[1:1]};
assign col_out_50 = {u_ca_out_50[0:0], u_ca_out_49[1:1]};
assign col_out_51 = {u_ca_out_51[0:0], u_ca_out_50[1:1]};
assign col_out_52 = {u_ca_out_52[0:0], u_ca_out_51[1:1]};
assign col_out_53 = {u_ca_out_53[0:0], u_ca_out_52[1:1]};
assign col_out_54 = {u_ca_out_54[0:0], u_ca_out_53[1:1]};
assign col_out_55 = {u_ca_out_55[0:0], u_ca_out_54[1:1]};
assign col_out_56 = {u_ca_out_56[0:0], u_ca_out_55[1:1]};
assign col_out_57 = {u_ca_out_57[0:0], u_ca_out_56[1:1]};
assign col_out_58 = {u_ca_out_58[0:0], u_ca_out_57[1:1]};
assign col_out_59 = {u_ca_out_59[0:0], u_ca_out_58[1:1]};
assign col_out_60 = {u_ca_out_60[0:0], u_ca_out_59[1:1]};
assign col_out_61 = {u_ca_out_61[0:0], u_ca_out_60[1:1]};
assign col_out_62 = {u_ca_out_62[0:0], u_ca_out_61[1:1]};
assign col_out_63 = {u_ca_out_63[0:0], u_ca_out_62[1:1]};
assign col_out_64 = {u_ca_out_64[0:0], u_ca_out_63[1:1]};
assign col_out_65 = {u_ca_out_65[0:0], u_ca_out_64[1:1]};
assign col_out_66 = {u_ca_out_66[0:0], u_ca_out_65[1:1]};
assign col_out_67 = {u_ca_out_67[0:0], u_ca_out_66[1:1]};
assign col_out_68 = {u_ca_out_68[0:0], u_ca_out_67[1:1]};
assign col_out_69 = {u_ca_out_69[0:0], u_ca_out_68[1:1]};
assign col_out_70 = {u_ca_out_70[0:0], u_ca_out_69[1:1]};
assign col_out_71 = {u_ca_out_71[0:0], u_ca_out_70[1:1]};
assign col_out_72 = {u_ca_out_72[0:0], u_ca_out_71[1:1]};
assign col_out_73 = {u_ca_out_73[0:0], u_ca_out_72[1:1]};
assign col_out_74 = {u_ca_out_74[0:0], u_ca_out_73[1:1]};
assign col_out_75 = {u_ca_out_75[0:0], u_ca_out_74[1:1]};
assign col_out_76 = {u_ca_out_76[0:0], u_ca_out_75[1:1]};
assign col_out_77 = {u_ca_out_77[0:0], u_ca_out_76[1:1]};
assign col_out_78 = {u_ca_out_78[0:0], u_ca_out_77[1:1]};
assign col_out_79 = {u_ca_out_79[0:0], u_ca_out_78[1:1]};
assign col_out_80 = {u_ca_out_80[0:0], u_ca_out_79[1:1]};
assign col_out_81 = {u_ca_out_81[0:0], u_ca_out_80[1:1]};
assign col_out_82 = {u_ca_out_82[0:0], u_ca_out_81[1:1]};
assign col_out_83 = {u_ca_out_83[0:0], u_ca_out_82[1:1]};
assign col_out_84 = {u_ca_out_84[0:0], u_ca_out_83[1:1]};
assign col_out_85 = {u_ca_out_85[0:0], u_ca_out_84[1:1]};
assign col_out_86 = {u_ca_out_86[0:0], u_ca_out_85[1:1]};
assign col_out_87 = {u_ca_out_87[0:0], u_ca_out_86[1:1]};
assign col_out_88 = {u_ca_out_88[0:0], u_ca_out_87[1:1]};
assign col_out_89 = {u_ca_out_89[0:0], u_ca_out_88[1:1]};
assign col_out_90 = {u_ca_out_90[0:0], u_ca_out_89[1:1]};
assign col_out_91 = {u_ca_out_91[0:0], u_ca_out_90[1:1]};
assign col_out_92 = {u_ca_out_92[0:0], u_ca_out_91[1:1]};
assign col_out_93 = {u_ca_out_93[0:0], u_ca_out_92[1:1]};
assign col_out_94 = {u_ca_out_94[0:0], u_ca_out_93[1:1]};
assign col_out_95 = {u_ca_out_95[0:0], u_ca_out_94[1:1]};
assign col_out_96 = {u_ca_out_96[0:0], u_ca_out_95[1:1]};
assign col_out_97 = {u_ca_out_97[0:0], u_ca_out_96[1:1]};
assign col_out_98 = {u_ca_out_98[0:0], u_ca_out_97[1:1]};
assign col_out_99 = {u_ca_out_99[0:0], u_ca_out_98[1:1]};
assign col_out_100 = {u_ca_out_100[0:0], u_ca_out_99[1:1]};
assign col_out_101 = {u_ca_out_101[0:0], u_ca_out_100[1:1]};
assign col_out_102 = {u_ca_out_102[0:0], u_ca_out_101[1:1]};
assign col_out_103 = {u_ca_out_103[0:0], u_ca_out_102[1:1]};
assign col_out_104 = {u_ca_out_104[0:0], u_ca_out_103[1:1]};
assign col_out_105 = {u_ca_out_105[0:0], u_ca_out_104[1:1]};
assign col_out_106 = {u_ca_out_106[0:0], u_ca_out_105[1:1]};
assign col_out_107 = {u_ca_out_107[0:0], u_ca_out_106[1:1]};
assign col_out_108 = {u_ca_out_108[0:0], u_ca_out_107[1:1]};
assign col_out_109 = {u_ca_out_109[0:0], u_ca_out_108[1:1]};
assign col_out_110 = {u_ca_out_110[0:0], u_ca_out_109[1:1]};
assign col_out_111 = {u_ca_out_111[0:0], u_ca_out_110[1:1]};
assign col_out_112 = {u_ca_out_112[0:0], u_ca_out_111[1:1]};
assign col_out_113 = {u_ca_out_113[0:0], u_ca_out_112[1:1]};
assign col_out_114 = {u_ca_out_114[0:0], u_ca_out_113[1:1]};
assign col_out_115 = {u_ca_out_115[0:0], u_ca_out_114[1:1]};
assign col_out_116 = {u_ca_out_116[0:0], u_ca_out_115[1:1]};
assign col_out_117 = {u_ca_out_117[0:0], u_ca_out_116[1:1]};
assign col_out_118 = {u_ca_out_118[0:0], u_ca_out_117[1:1]};
assign col_out_119 = {u_ca_out_119[0:0], u_ca_out_118[1:1]};
assign col_out_120 = {u_ca_out_120[0:0], u_ca_out_119[1:1]};
assign col_out_121 = {u_ca_out_121[0:0], u_ca_out_120[1:1]};
assign col_out_122 = {u_ca_out_122[0:0], u_ca_out_121[1:1]};
assign col_out_123 = {u_ca_out_123[0:0], u_ca_out_122[1:1]};
assign col_out_124 = {u_ca_out_124[0:0], u_ca_out_123[1:1]};
assign col_out_125 = {u_ca_out_125[0:0], u_ca_out_124[1:1]};
assign col_out_126 = {u_ca_out_126[0:0], u_ca_out_125[1:1]};
assign col_out_127 = {u_ca_out_127[0:0], u_ca_out_126[1:1]};
assign col_out_128 = {u_ca_out_128[0:0], u_ca_out_127[1:1]};
assign col_out_129 = {u_ca_out_129[0:0], u_ca_out_128[1:1]};
assign col_out_130 = {u_ca_out_130[0:0], u_ca_out_129[1:1]};
assign col_out_131 = {u_ca_out_131[0:0], u_ca_out_130[1:1]};
assign col_out_132 = {u_ca_out_132[0:0], u_ca_out_131[1:1]};
assign col_out_133 = {u_ca_out_133[0:0], u_ca_out_132[1:1]};
assign col_out_134 = {u_ca_out_134[0:0], u_ca_out_133[1:1]};
assign col_out_135 = {u_ca_out_135[0:0], u_ca_out_134[1:1]};
assign col_out_136 = {u_ca_out_136[0:0], u_ca_out_135[1:1]};
assign col_out_137 = {u_ca_out_137[0:0], u_ca_out_136[1:1]};
assign col_out_138 = {u_ca_out_138[0:0], u_ca_out_137[1:1]};
assign col_out_139 = {u_ca_out_139[0:0], u_ca_out_138[1:1]};
assign col_out_140 = {u_ca_out_140[0:0], u_ca_out_139[1:1]};
assign col_out_141 = {u_ca_out_141[0:0], u_ca_out_140[1:1]};
assign col_out_142 = {u_ca_out_142[0:0], u_ca_out_141[1:1]};
assign col_out_143 = {u_ca_out_143[0:0], u_ca_out_142[1:1]};
assign col_out_144 = {u_ca_out_144[0:0], u_ca_out_143[1:1]};
assign col_out_145 = {u_ca_out_145[0:0], u_ca_out_144[1:1]};
assign col_out_146 = {u_ca_out_146[0:0], u_ca_out_145[1:1]};
assign col_out_147 = {u_ca_out_147[0:0], u_ca_out_146[1:1]};
assign col_out_148 = {u_ca_out_148[0:0], u_ca_out_147[1:1]};
assign col_out_149 = {u_ca_out_149[0:0], u_ca_out_148[1:1]};
assign col_out_150 = {u_ca_out_150[0:0], u_ca_out_149[1:1]};
assign col_out_151 = {u_ca_out_151[0:0], u_ca_out_150[1:1]};
assign col_out_152 = {u_ca_out_152[0:0], u_ca_out_151[1:1]};
assign col_out_153 = {u_ca_out_153[0:0], u_ca_out_152[1:1]};
assign col_out_154 = {u_ca_out_154[0:0], u_ca_out_153[1:1]};
assign col_out_155 = {u_ca_out_155[0:0], u_ca_out_154[1:1]};
assign col_out_156 = {u_ca_out_156[0:0], u_ca_out_155[1:1]};
assign col_out_157 = {u_ca_out_157[0:0], u_ca_out_156[1:1]};
assign col_out_158 = {u_ca_out_158[0:0], u_ca_out_157[1:1]};
assign col_out_159 = {u_ca_out_159[0:0], u_ca_out_158[1:1]};
assign col_out_160 = {u_ca_out_160[0:0], u_ca_out_159[1:1]};
assign col_out_161 = {u_ca_out_161[0:0], u_ca_out_160[1:1]};
assign col_out_162 = {u_ca_out_162[0:0], u_ca_out_161[1:1]};
assign col_out_163 = {u_ca_out_163[0:0], u_ca_out_162[1:1]};
assign col_out_164 = {u_ca_out_164[0:0], u_ca_out_163[1:1]};
assign col_out_165 = {u_ca_out_165[0:0], u_ca_out_164[1:1]};
assign col_out_166 = {u_ca_out_166[0:0], u_ca_out_165[1:1]};
assign col_out_167 = {u_ca_out_167[0:0], u_ca_out_166[1:1]};
assign col_out_168 = {u_ca_out_168[0:0], u_ca_out_167[1:1]};
assign col_out_169 = {u_ca_out_169[0:0], u_ca_out_168[1:1]};
assign col_out_170 = {u_ca_out_170[0:0], u_ca_out_169[1:1]};
assign col_out_171 = {u_ca_out_171[0:0], u_ca_out_170[1:1]};
assign col_out_172 = {u_ca_out_172[0:0], u_ca_out_171[1:1]};
assign col_out_173 = {u_ca_out_173[0:0], u_ca_out_172[1:1]};
assign col_out_174 = {u_ca_out_174[0:0], u_ca_out_173[1:1]};
assign col_out_175 = {u_ca_out_175[0:0], u_ca_out_174[1:1]};
assign col_out_176 = {u_ca_out_176[0:0], u_ca_out_175[1:1]};
assign col_out_177 = {u_ca_out_177[0:0], u_ca_out_176[1:1]};
assign col_out_178 = {u_ca_out_178[0:0], u_ca_out_177[1:1]};
assign col_out_179 = {u_ca_out_179[0:0], u_ca_out_178[1:1]};
assign col_out_180 = {u_ca_out_180[0:0], u_ca_out_179[1:1]};
assign col_out_181 = {u_ca_out_181[0:0], u_ca_out_180[1:1]};
assign col_out_182 = {u_ca_out_182[0:0], u_ca_out_181[1:1]};
assign col_out_183 = {u_ca_out_183[0:0], u_ca_out_182[1:1]};
assign col_out_184 = {u_ca_out_184[0:0], u_ca_out_183[1:1]};
assign col_out_185 = {u_ca_out_185[0:0], u_ca_out_184[1:1]};
assign col_out_186 = {u_ca_out_186[0:0], u_ca_out_185[1:1]};
assign col_out_187 = {u_ca_out_187[0:0], u_ca_out_186[1:1]};
assign col_out_188 = {u_ca_out_188[0:0], u_ca_out_187[1:1]};
assign col_out_189 = {u_ca_out_189[0:0], u_ca_out_188[1:1]};
assign col_out_190 = {u_ca_out_190[0:0], u_ca_out_189[1:1]};
assign col_out_191 = {u_ca_out_191[0:0], u_ca_out_190[1:1]};
assign col_out_192 = {u_ca_out_192[0:0], u_ca_out_191[1:1]};
assign col_out_193 = {u_ca_out_193[0:0], u_ca_out_192[1:1]};
assign col_out_194 = {u_ca_out_194[0:0], u_ca_out_193[1:1]};
assign col_out_195 = {u_ca_out_195[0:0], u_ca_out_194[1:1]};
assign col_out_196 = {u_ca_out_196[0:0], u_ca_out_195[1:1]};
assign col_out_197 = {u_ca_out_197[0:0], u_ca_out_196[1:1]};
assign col_out_198 = {u_ca_out_198[0:0], u_ca_out_197[1:1]};
assign col_out_199 = {u_ca_out_199[0:0], u_ca_out_198[1:1]};
assign col_out_200 = {u_ca_out_200[0:0], u_ca_out_199[1:1]};
assign col_out_201 = {u_ca_out_201[0:0], u_ca_out_200[1:1]};
assign col_out_202 = {u_ca_out_202[0:0], u_ca_out_201[1:1]};
assign col_out_203 = {u_ca_out_203[0:0], u_ca_out_202[1:1]};
assign col_out_204 = {u_ca_out_204[0:0], u_ca_out_203[1:1]};
assign col_out_205 = {u_ca_out_205[0:0], u_ca_out_204[1:1]};
assign col_out_206 = {u_ca_out_206[0:0], u_ca_out_205[1:1]};
assign col_out_207 = {u_ca_out_207[0:0], u_ca_out_206[1:1]};
assign col_out_208 = {u_ca_out_208[0:0], u_ca_out_207[1:1]};
assign col_out_209 = {u_ca_out_209[0:0], u_ca_out_208[1:1]};
assign col_out_210 = {u_ca_out_210[0:0], u_ca_out_209[1:1]};
assign col_out_211 = {u_ca_out_211[0:0], u_ca_out_210[1:1]};
assign col_out_212 = {u_ca_out_212[0:0], u_ca_out_211[1:1]};
assign col_out_213 = {u_ca_out_213[0:0], u_ca_out_212[1:1]};
assign col_out_214 = {u_ca_out_214[0:0], u_ca_out_213[1:1]};
assign col_out_215 = {u_ca_out_215[0:0], u_ca_out_214[1:1]};
assign col_out_216 = {u_ca_out_216[0:0], u_ca_out_215[1:1]};
assign col_out_217 = {u_ca_out_217[0:0], u_ca_out_216[1:1]};
assign col_out_218 = {u_ca_out_218[0:0], u_ca_out_217[1:1]};
assign col_out_219 = {u_ca_out_219[0:0], u_ca_out_218[1:1]};
assign col_out_220 = {u_ca_out_220[0:0], u_ca_out_219[1:1]};
assign col_out_221 = {u_ca_out_221[0:0], u_ca_out_220[1:1]};
assign col_out_222 = {u_ca_out_222[0:0], u_ca_out_221[1:1]};
assign col_out_223 = {u_ca_out_223[0:0], u_ca_out_222[1:1]};
assign col_out_224 = {u_ca_out_224[0:0], u_ca_out_223[1:1]};
assign col_out_225 = {u_ca_out_225[0:0], u_ca_out_224[1:1]};
assign col_out_226 = {u_ca_out_226[0:0], u_ca_out_225[1:1]};
assign col_out_227 = {u_ca_out_227[0:0], u_ca_out_226[1:1]};
assign col_out_228 = {u_ca_out_228[0:0], u_ca_out_227[1:1]};
assign col_out_229 = {u_ca_out_229[0:0], u_ca_out_228[1:1]};
assign col_out_230 = {u_ca_out_230[0:0], u_ca_out_229[1:1]};
assign col_out_231 = {u_ca_out_231[0:0], u_ca_out_230[1:1]};
assign col_out_232 = {u_ca_out_232[0:0], u_ca_out_231[1:1]};
assign col_out_233 = {u_ca_out_233[0:0], u_ca_out_232[1:1]};
assign col_out_234 = {u_ca_out_234[0:0], u_ca_out_233[1:1]};
assign col_out_235 = {u_ca_out_235[0:0], u_ca_out_234[1:1]};
assign col_out_236 = {u_ca_out_236[0:0], u_ca_out_235[1:1]};
assign col_out_237 = {u_ca_out_237[0:0], u_ca_out_236[1:1]};
assign col_out_238 = {u_ca_out_238[0:0], u_ca_out_237[1:1]};
assign col_out_239 = {u_ca_out_239[0:0], u_ca_out_238[1:1]};
assign col_out_240 = {u_ca_out_240[0:0], u_ca_out_239[1:1]};
assign col_out_241 = {u_ca_out_241[0:0], u_ca_out_240[1:1]};
assign col_out_242 = {u_ca_out_242[0:0], u_ca_out_241[1:1]};
assign col_out_243 = {u_ca_out_243[0:0], u_ca_out_242[1:1]};
assign col_out_244 = {u_ca_out_244[0:0], u_ca_out_243[1:1]};
assign col_out_245 = {u_ca_out_245[0:0], u_ca_out_244[1:1]};
assign col_out_246 = {u_ca_out_246[0:0], u_ca_out_245[1:1]};
assign col_out_247 = {u_ca_out_247[0:0], u_ca_out_246[1:1]};
assign col_out_248 = {u_ca_out_248[0:0], u_ca_out_247[1:1]};
assign col_out_249 = {u_ca_out_249[0:0], u_ca_out_248[1:1]};
assign col_out_250 = {u_ca_out_250[0:0], u_ca_out_249[1:1]};
assign col_out_251 = {u_ca_out_251[0:0], u_ca_out_250[1:1]};
assign col_out_252 = {u_ca_out_252[0:0], u_ca_out_251[1:1]};
assign col_out_253 = {u_ca_out_253[0:0], u_ca_out_252[1:1]};
assign col_out_254 = {u_ca_out_254[0:0], u_ca_out_253[1:1]};
assign col_out_255 = {u_ca_out_255[0:0], u_ca_out_254[1:1]};
assign col_out_256 = {u_ca_out_256[0:0], u_ca_out_255[1:1]};
assign col_out_257 = {u_ca_out_257[0:0], u_ca_out_256[1:1]};
assign col_out_258 = {u_ca_out_258[0:0], u_ca_out_257[1:1]};
assign col_out_259 = {u_ca_out_259[0:0], u_ca_out_258[1:1]};
assign col_out_260 = {u_ca_out_260[0:0], u_ca_out_259[1:1]};
assign col_out_261 = {u_ca_out_261[0:0], u_ca_out_260[1:1]};
assign col_out_262 = {u_ca_out_262[0:0], u_ca_out_261[1:1]};
assign col_out_263 = {u_ca_out_263[0:0], u_ca_out_262[1:1]};
assign col_out_264 = {u_ca_out_264[0:0], u_ca_out_263[1:1]};
assign col_out_265 = {u_ca_out_265[0:0], u_ca_out_264[1:1]};
assign col_out_266 = {u_ca_out_266[0:0], u_ca_out_265[1:1]};
assign col_out_267 = {u_ca_out_267[0:0], u_ca_out_266[1:1]};
assign col_out_268 = {u_ca_out_268[0:0], u_ca_out_267[1:1]};
assign col_out_269 = {u_ca_out_269[0:0], u_ca_out_268[1:1]};
assign col_out_270 = {u_ca_out_270[0:0], u_ca_out_269[1:1]};
assign col_out_271 = {u_ca_out_271[0:0], u_ca_out_270[1:1]};
assign col_out_272 = {u_ca_out_272[0:0], u_ca_out_271[1:1]};
assign col_out_273 = {u_ca_out_273[0:0], u_ca_out_272[1:1]};
assign col_out_274 = {u_ca_out_274[0:0], u_ca_out_273[1:1]};
assign col_out_275 = {u_ca_out_275[0:0], u_ca_out_274[1:1]};
assign col_out_276 = {u_ca_out_276[0:0], u_ca_out_275[1:1]};
assign col_out_277 = {u_ca_out_277[0:0], u_ca_out_276[1:1]};
assign col_out_278 = {u_ca_out_278[0:0], u_ca_out_277[1:1]};
assign col_out_279 = {u_ca_out_279[0:0], u_ca_out_278[1:1]};
assign col_out_280 = {u_ca_out_280[0:0], u_ca_out_279[1:1]};
assign col_out_281 = {u_ca_out_281[0:0], u_ca_out_280[1:1]};
assign col_out_282 = {u_ca_out_282[0:0], u_ca_out_281[1:1]};
assign col_out_283 = {u_ca_out_283[0:0], u_ca_out_282[1:1]};
assign col_out_284 = {u_ca_out_284[0:0], u_ca_out_283[1:1]};
assign col_out_285 = {u_ca_out_285[0:0], u_ca_out_284[1:1]};
assign col_out_286 = {u_ca_out_286[0:0], u_ca_out_285[1:1]};
assign col_out_287 = {u_ca_out_287[0:0], u_ca_out_286[1:1]};
assign col_out_288 = {u_ca_out_288[0:0], u_ca_out_287[1:1]};
assign col_out_289 = {u_ca_out_289[0:0], u_ca_out_288[1:1]};
assign col_out_290 = {u_ca_out_290[0:0], u_ca_out_289[1:1]};
assign col_out_291 = {u_ca_out_291[0:0], u_ca_out_290[1:1]};
assign col_out_292 = {u_ca_out_292[0:0], u_ca_out_291[1:1]};
assign col_out_293 = {u_ca_out_293[0:0], u_ca_out_292[1:1]};
assign col_out_294 = {u_ca_out_294[0:0], u_ca_out_293[1:1]};
assign col_out_295 = {u_ca_out_295[0:0], u_ca_out_294[1:1]};
assign col_out_296 = {u_ca_out_296[0:0], u_ca_out_295[1:1]};
assign col_out_297 = {u_ca_out_297[0:0], u_ca_out_296[1:1]};
assign col_out_298 = {u_ca_out_298[0:0], u_ca_out_297[1:1]};
assign col_out_299 = {u_ca_out_299[0:0], u_ca_out_298[1:1]};
assign col_out_300 = {u_ca_out_300[0:0], u_ca_out_299[1:1]};
assign col_out_301 = {u_ca_out_301[0:0], u_ca_out_300[1:1]};
assign col_out_302 = {u_ca_out_302[0:0], u_ca_out_301[1:1]};
assign col_out_303 = {u_ca_out_303[0:0], u_ca_out_302[1:1]};
assign col_out_304 = {u_ca_out_304[0:0], u_ca_out_303[1:1]};
assign col_out_305 = {u_ca_out_305[0:0], u_ca_out_304[1:1]};
assign col_out_306 = {u_ca_out_306[0:0], u_ca_out_305[1:1]};
assign col_out_307 = {u_ca_out_307[0:0], u_ca_out_306[1:1]};
assign col_out_308 = {u_ca_out_308[0:0], u_ca_out_307[1:1]};
assign col_out_309 = {u_ca_out_309[0:0], u_ca_out_308[1:1]};
assign col_out_310 = {u_ca_out_310[0:0], u_ca_out_309[1:1]};
assign col_out_311 = {u_ca_out_311[0:0], u_ca_out_310[1:1]};
assign col_out_312 = {u_ca_out_312[0:0], u_ca_out_311[1:1]};
assign col_out_313 = {u_ca_out_313[0:0], u_ca_out_312[1:1]};
assign col_out_314 = {u_ca_out_314[0:0], u_ca_out_313[1:1]};
assign col_out_315 = {u_ca_out_315[0:0], u_ca_out_314[1:1]};
assign col_out_316 = {u_ca_out_316[0:0], u_ca_out_315[1:1]};
assign col_out_317 = {u_ca_out_317[0:0], u_ca_out_316[1:1]};
assign col_out_318 = {u_ca_out_318[0:0], u_ca_out_317[1:1]};
assign col_out_319 = {u_ca_out_319[0:0], u_ca_out_318[1:1]};
assign col_out_320 = {u_ca_out_320[0:0], u_ca_out_319[1:1]};
assign col_out_321 = {u_ca_out_321[0:0], u_ca_out_320[1:1]};
assign col_out_322 = {u_ca_out_322[0:0], u_ca_out_321[1:1]};
assign col_out_323 = {u_ca_out_323[0:0], u_ca_out_322[1:1]};
assign col_out_324 = {u_ca_out_324[0:0], u_ca_out_323[1:1]};
assign col_out_325 = {u_ca_out_325[0:0], u_ca_out_324[1:1]};
assign col_out_326 = {u_ca_out_326[0:0], u_ca_out_325[1:1]};
assign col_out_327 = {u_ca_out_327[0:0], u_ca_out_326[1:1]};
assign col_out_328 = {u_ca_out_328[0:0], u_ca_out_327[1:1]};
assign col_out_329 = {u_ca_out_329[0:0], u_ca_out_328[1:1]};
assign col_out_330 = {u_ca_out_330[0:0], u_ca_out_329[1:1]};
assign col_out_331 = {u_ca_out_331[0:0], u_ca_out_330[1:1]};
assign col_out_332 = {u_ca_out_332[0:0], u_ca_out_331[1:1]};
assign col_out_333 = {u_ca_out_333[0:0], u_ca_out_332[1:1]};
assign col_out_334 = {u_ca_out_334[0:0], u_ca_out_333[1:1]};
assign col_out_335 = {u_ca_out_335[0:0], u_ca_out_334[1:1]};
assign col_out_336 = {u_ca_out_336[0:0], u_ca_out_335[1:1]};
assign col_out_337 = {u_ca_out_337[0:0], u_ca_out_336[1:1]};
assign col_out_338 = {u_ca_out_338[0:0], u_ca_out_337[1:1]};
assign col_out_339 = {u_ca_out_339[0:0], u_ca_out_338[1:1]};
assign col_out_340 = {u_ca_out_340[0:0], u_ca_out_339[1:1]};
assign col_out_341 = {u_ca_out_341[0:0], u_ca_out_340[1:1]};
assign col_out_342 = {u_ca_out_342[0:0], u_ca_out_341[1:1]};
assign col_out_343 = {u_ca_out_343[0:0], u_ca_out_342[1:1]};
assign col_out_344 = {u_ca_out_344[0:0], u_ca_out_343[1:1]};
assign col_out_345 = {u_ca_out_345[0:0], u_ca_out_344[1:1]};
assign col_out_346 = {u_ca_out_346[0:0], u_ca_out_345[1:1]};
assign col_out_347 = {u_ca_out_347[0:0], u_ca_out_346[1:1]};
assign col_out_348 = {u_ca_out_348[0:0], u_ca_out_347[1:1]};
assign col_out_349 = {u_ca_out_349[0:0], u_ca_out_348[1:1]};
assign col_out_350 = {u_ca_out_350[0:0], u_ca_out_349[1:1]};
assign col_out_351 = {u_ca_out_351[0:0], u_ca_out_350[1:1]};
assign col_out_352 = {u_ca_out_352[0:0], u_ca_out_351[1:1]};
assign col_out_353 = {u_ca_out_353[0:0], u_ca_out_352[1:1]};
assign col_out_354 = {u_ca_out_354[0:0], u_ca_out_353[1:1]};
assign col_out_355 = {u_ca_out_355[0:0], u_ca_out_354[1:1]};
assign col_out_356 = {u_ca_out_356[0:0], u_ca_out_355[1:1]};
assign col_out_357 = {u_ca_out_357[0:0], u_ca_out_356[1:1]};
assign col_out_358 = {u_ca_out_358[0:0], u_ca_out_357[1:1]};
assign col_out_359 = {u_ca_out_359[0:0], u_ca_out_358[1:1]};
assign col_out_360 = {u_ca_out_360[0:0], u_ca_out_359[1:1]};
assign col_out_361 = {u_ca_out_361[0:0], u_ca_out_360[1:1]};
assign col_out_362 = {u_ca_out_362[0:0], u_ca_out_361[1:1]};
assign col_out_363 = {u_ca_out_363[0:0], u_ca_out_362[1:1]};
assign col_out_364 = {u_ca_out_364[0:0], u_ca_out_363[1:1]};
assign col_out_365 = {u_ca_out_365[0:0], u_ca_out_364[1:1]};
assign col_out_366 = {u_ca_out_366[0:0], u_ca_out_365[1:1]};
assign col_out_367 = {u_ca_out_367[0:0], u_ca_out_366[1:1]};
assign col_out_368 = {u_ca_out_368[0:0], u_ca_out_367[1:1]};
assign col_out_369 = {u_ca_out_369[0:0], u_ca_out_368[1:1]};
assign col_out_370 = {u_ca_out_370[0:0], u_ca_out_369[1:1]};
assign col_out_371 = {u_ca_out_371[0:0], u_ca_out_370[1:1]};
assign col_out_372 = {u_ca_out_372[0:0], u_ca_out_371[1:1]};
assign col_out_373 = {u_ca_out_373[0:0], u_ca_out_372[1:1]};
assign col_out_374 = {u_ca_out_374[0:0], u_ca_out_373[1:1]};
assign col_out_375 = {u_ca_out_375[0:0], u_ca_out_374[1:1]};
assign col_out_376 = {u_ca_out_376[0:0], u_ca_out_375[1:1]};
assign col_out_377 = {u_ca_out_377[0:0], u_ca_out_376[1:1]};
assign col_out_378 = {u_ca_out_378[0:0], u_ca_out_377[1:1]};
assign col_out_379 = {u_ca_out_379[0:0], u_ca_out_378[1:1]};
assign col_out_380 = {u_ca_out_380[0:0], u_ca_out_379[1:1]};
assign col_out_381 = {u_ca_out_381[0:0], u_ca_out_380[1:1]};
assign col_out_382 = {u_ca_out_382[0:0], u_ca_out_381[1:1]};
assign col_out_383 = {u_ca_out_383[0:0], u_ca_out_382[1:1]};
assign col_out_384 = {u_ca_out_384[0:0], u_ca_out_383[1:1]};
assign col_out_385 = {u_ca_out_385[0:0], u_ca_out_384[1:1]};
assign col_out_386 = {u_ca_out_386[0:0], u_ca_out_385[1:1]};
assign col_out_387 = {u_ca_out_387[0:0], u_ca_out_386[1:1]};
assign col_out_388 = {u_ca_out_388[0:0], u_ca_out_387[1:1]};
assign col_out_389 = {u_ca_out_389[0:0], u_ca_out_388[1:1]};
assign col_out_390 = {u_ca_out_390[0:0], u_ca_out_389[1:1]};
assign col_out_391 = {u_ca_out_391[0:0], u_ca_out_390[1:1]};
assign col_out_392 = {u_ca_out_392[0:0], u_ca_out_391[1:1]};
assign col_out_393 = {u_ca_out_393[0:0], u_ca_out_392[1:1]};
assign col_out_394 = {u_ca_out_394[0:0], u_ca_out_393[1:1]};
assign col_out_395 = {u_ca_out_395[0:0], u_ca_out_394[1:1]};
assign col_out_396 = {u_ca_out_396[0:0], u_ca_out_395[1:1]};
assign col_out_397 = {u_ca_out_397[0:0], u_ca_out_396[1:1]};
assign col_out_398 = {u_ca_out_398[0:0], u_ca_out_397[1:1]};
assign col_out_399 = {u_ca_out_399[0:0], u_ca_out_398[1:1]};
assign col_out_400 = {u_ca_out_400[0:0], u_ca_out_399[1:1]};
assign col_out_401 = {u_ca_out_401[0:0], u_ca_out_400[1:1]};
assign col_out_402 = {u_ca_out_402[0:0], u_ca_out_401[1:1]};
assign col_out_403 = {u_ca_out_403[0:0], u_ca_out_402[1:1]};
assign col_out_404 = {u_ca_out_404[0:0], u_ca_out_403[1:1]};
assign col_out_405 = {u_ca_out_405[0:0], u_ca_out_404[1:1]};
assign col_out_406 = {u_ca_out_406[0:0], u_ca_out_405[1:1]};
assign col_out_407 = {u_ca_out_407[0:0], u_ca_out_406[1:1]};
assign col_out_408 = {u_ca_out_408[0:0], u_ca_out_407[1:1]};
assign col_out_409 = {u_ca_out_409[0:0], u_ca_out_408[1:1]};
assign col_out_410 = {u_ca_out_410[0:0], u_ca_out_409[1:1]};
assign col_out_411 = {u_ca_out_411[0:0], u_ca_out_410[1:1]};
assign col_out_412 = {u_ca_out_412[0:0], u_ca_out_411[1:1]};
assign col_out_413 = {u_ca_out_413[0:0], u_ca_out_412[1:1]};
assign col_out_414 = {u_ca_out_414[0:0], u_ca_out_413[1:1]};
assign col_out_415 = {u_ca_out_415[0:0], u_ca_out_414[1:1]};
assign col_out_416 = {u_ca_out_416[0:0], u_ca_out_415[1:1]};
assign col_out_417 = {u_ca_out_417[0:0], u_ca_out_416[1:1]};
assign col_out_418 = {u_ca_out_418[0:0], u_ca_out_417[1:1]};
assign col_out_419 = {u_ca_out_419[0:0], u_ca_out_418[1:1]};
assign col_out_420 = {u_ca_out_420[0:0], u_ca_out_419[1:1]};
assign col_out_421 = {u_ca_out_421[0:0], u_ca_out_420[1:1]};
assign col_out_422 = {u_ca_out_422[0:0], u_ca_out_421[1:1]};
assign col_out_423 = {u_ca_out_423[0:0], u_ca_out_422[1:1]};
assign col_out_424 = {u_ca_out_424[0:0], u_ca_out_423[1:1]};
assign col_out_425 = {u_ca_out_425[0:0], u_ca_out_424[1:1]};
assign col_out_426 = {u_ca_out_426[0:0], u_ca_out_425[1:1]};
assign col_out_427 = {u_ca_out_427[0:0], u_ca_out_426[1:1]};
assign col_out_428 = {u_ca_out_428[0:0], u_ca_out_427[1:1]};
assign col_out_429 = {u_ca_out_429[0:0], u_ca_out_428[1:1]};
assign col_out_430 = {u_ca_out_430[0:0], u_ca_out_429[1:1]};
assign col_out_431 = {u_ca_out_431[0:0], u_ca_out_430[1:1]};
assign col_out_432 = {u_ca_out_432[0:0], u_ca_out_431[1:1]};
assign col_out_433 = {u_ca_out_433[0:0], u_ca_out_432[1:1]};
assign col_out_434 = {u_ca_out_434[0:0], u_ca_out_433[1:1]};
assign col_out_435 = {u_ca_out_435[0:0], u_ca_out_434[1:1]};
assign col_out_436 = {u_ca_out_436[0:0], u_ca_out_435[1:1]};
assign col_out_437 = {u_ca_out_437[0:0], u_ca_out_436[1:1]};
assign col_out_438 = {u_ca_out_438[0:0], u_ca_out_437[1:1]};
assign col_out_439 = {u_ca_out_439[0:0], u_ca_out_438[1:1]};
assign col_out_440 = {u_ca_out_440[0:0], u_ca_out_439[1:1]};
assign col_out_441 = {u_ca_out_441[0:0], u_ca_out_440[1:1]};
assign col_out_442 = {u_ca_out_442[0:0], u_ca_out_441[1:1]};
assign col_out_443 = {u_ca_out_443[0:0], u_ca_out_442[1:1]};
assign col_out_444 = {u_ca_out_444[0:0], u_ca_out_443[1:1]};
assign col_out_445 = {u_ca_out_445[0:0], u_ca_out_444[1:1]};
assign col_out_446 = {u_ca_out_446[0:0], u_ca_out_445[1:1]};
assign col_out_447 = {u_ca_out_447[0:0], u_ca_out_446[1:1]};
assign col_out_448 = {u_ca_out_448[0:0], u_ca_out_447[1:1]};
assign col_out_449 = {u_ca_out_449[0:0], u_ca_out_448[1:1]};
assign col_out_450 = {u_ca_out_450[0:0], u_ca_out_449[1:1]};
assign col_out_451 = {u_ca_out_451[0:0], u_ca_out_450[1:1]};
assign col_out_452 = {u_ca_out_452[0:0], u_ca_out_451[1:1]};
assign col_out_453 = {u_ca_out_453[0:0], u_ca_out_452[1:1]};
assign col_out_454 = {u_ca_out_454[0:0], u_ca_out_453[1:1]};
assign col_out_455 = {u_ca_out_455[0:0], u_ca_out_454[1:1]};
assign col_out_456 = {u_ca_out_456[0:0], u_ca_out_455[1:1]};
assign col_out_457 = {u_ca_out_457[0:0], u_ca_out_456[1:1]};
assign col_out_458 = {u_ca_out_458[0:0], u_ca_out_457[1:1]};
assign col_out_459 = {u_ca_out_459[0:0], u_ca_out_458[1:1]};
assign col_out_460 = {u_ca_out_460[0:0], u_ca_out_459[1:1]};
assign col_out_461 = {u_ca_out_461[0:0], u_ca_out_460[1:1]};
assign col_out_462 = {u_ca_out_462[0:0], u_ca_out_461[1:1]};
assign col_out_463 = {u_ca_out_463[0:0], u_ca_out_462[1:1]};
assign col_out_464 = {u_ca_out_464[0:0], u_ca_out_463[1:1]};
assign col_out_465 = {u_ca_out_465[0:0], u_ca_out_464[1:1]};
assign col_out_466 = {u_ca_out_466[0:0], u_ca_out_465[1:1]};
assign col_out_467 = {u_ca_out_467[0:0], u_ca_out_466[1:1]};
assign col_out_468 = {u_ca_out_468[0:0], u_ca_out_467[1:1]};
assign col_out_469 = {u_ca_out_469[0:0], u_ca_out_468[1:1]};
assign col_out_470 = {u_ca_out_470[0:0], u_ca_out_469[1:1]};
assign col_out_471 = {u_ca_out_471[0:0], u_ca_out_470[1:1]};
assign col_out_472 = {u_ca_out_472[0:0], u_ca_out_471[1:1]};
assign col_out_473 = {u_ca_out_473[0:0], u_ca_out_472[1:1]};
assign col_out_474 = {u_ca_out_474[0:0], u_ca_out_473[1:1]};
assign col_out_475 = {u_ca_out_475[0:0], u_ca_out_474[1:1]};
assign col_out_476 = {u_ca_out_476[0:0], u_ca_out_475[1:1]};
assign col_out_477 = {u_ca_out_477[0:0], u_ca_out_476[1:1]};
assign col_out_478 = {u_ca_out_478[0:0], u_ca_out_477[1:1]};
assign col_out_479 = {u_ca_out_479[0:0], u_ca_out_478[1:1]};
assign col_out_480 = {u_ca_out_480[0:0], u_ca_out_479[1:1]};
assign col_out_481 = {u_ca_out_481[0:0], u_ca_out_480[1:1]};
assign col_out_482 = {u_ca_out_482[0:0], u_ca_out_481[1:1]};
assign col_out_483 = {u_ca_out_483[0:0], u_ca_out_482[1:1]};
assign col_out_484 = {u_ca_out_484[0:0], u_ca_out_483[1:1]};
assign col_out_485 = {u_ca_out_485[0:0], u_ca_out_484[1:1]};
assign col_out_486 = {u_ca_out_486[0:0], u_ca_out_485[1:1]};
assign col_out_487 = {u_ca_out_487[0:0], u_ca_out_486[1:1]};
assign col_out_488 = {u_ca_out_488[0:0], u_ca_out_487[1:1]};
assign col_out_489 = {u_ca_out_489[0:0], u_ca_out_488[1:1]};
assign col_out_490 = {u_ca_out_490[0:0], u_ca_out_489[1:1]};
assign col_out_491 = {u_ca_out_491[0:0], u_ca_out_490[1:1]};
assign col_out_492 = {u_ca_out_492[0:0], u_ca_out_491[1:1]};
assign col_out_493 = {u_ca_out_493[0:0], u_ca_out_492[1:1]};
assign col_out_494 = {u_ca_out_494[0:0], u_ca_out_493[1:1]};
assign col_out_495 = {u_ca_out_495[0:0], u_ca_out_494[1:1]};
assign col_out_496 = {u_ca_out_496[0:0], u_ca_out_495[1:1]};
assign col_out_497 = {u_ca_out_497[0:0], u_ca_out_496[1:1]};
assign col_out_498 = {u_ca_out_498[0:0], u_ca_out_497[1:1]};
assign col_out_499 = {u_ca_out_499[0:0], u_ca_out_498[1:1]};
assign col_out_500 = {u_ca_out_500[0:0], u_ca_out_499[1:1]};
assign col_out_501 = {u_ca_out_501[0:0], u_ca_out_500[1:1]};
assign col_out_502 = {u_ca_out_502[0:0], u_ca_out_501[1:1]};
assign col_out_503 = {u_ca_out_503[0:0], u_ca_out_502[1:1]};
assign col_out_504 = {u_ca_out_504[0:0], u_ca_out_503[1:1]};
assign col_out_505 = {u_ca_out_505[0:0], u_ca_out_504[1:1]};
assign col_out_506 = {u_ca_out_506[0:0], u_ca_out_505[1:1]};
assign col_out_507 = {u_ca_out_507[0:0], u_ca_out_506[1:1]};
assign col_out_508 = {u_ca_out_508[0:0], u_ca_out_507[1:1]};
assign col_out_509 = {u_ca_out_509[0:0], u_ca_out_508[1:1]};
assign col_out_510 = {u_ca_out_510[0:0], u_ca_out_509[1:1]};
assign col_out_511 = {u_ca_out_511[0:0], u_ca_out_510[1:1]};
assign col_out_512 = {u_ca_out_512[0:0], u_ca_out_511[1:1]};
assign col_out_513 = {u_ca_out_513[0:0], u_ca_out_512[1:1]};
assign col_out_514 = {u_ca_out_514[0:0], u_ca_out_513[1:1]};
assign col_out_515 = {u_ca_out_515[0:0], u_ca_out_514[1:1]};
assign col_out_516 = {u_ca_out_516[0:0], u_ca_out_515[1:1]};
assign col_out_517 = {u_ca_out_517[0:0], u_ca_out_516[1:1]};
assign col_out_518 = {u_ca_out_518[0:0], u_ca_out_517[1:1]};
assign col_out_519 = {u_ca_out_519[0:0], u_ca_out_518[1:1]};
assign col_out_520 = {u_ca_out_520[0:0], u_ca_out_519[1:1]};
assign col_out_521 = {u_ca_out_521[0:0], u_ca_out_520[1:1]};
assign col_out_522 = {u_ca_out_522[0:0], u_ca_out_521[1:1]};
assign col_out_523 = {u_ca_out_523[0:0], u_ca_out_522[1:1]};
assign col_out_524 = {u_ca_out_524[0:0], u_ca_out_523[1:1]};
assign col_out_525 = {u_ca_out_525[0:0], u_ca_out_524[1:1]};
assign col_out_526 = {u_ca_out_526[0:0], u_ca_out_525[1:1]};
assign col_out_527 = {u_ca_out_527[0:0], u_ca_out_526[1:1]};
assign col_out_528 = {u_ca_out_528[0:0], u_ca_out_527[1:1]};
assign col_out_529 = {u_ca_out_529[0:0], u_ca_out_528[1:1]};
assign col_out_530 = {u_ca_out_530[0:0], u_ca_out_529[1:1]};
assign col_out_531 = {u_ca_out_531[0:0], u_ca_out_530[1:1]};
assign col_out_532 = {u_ca_out_532[0:0], u_ca_out_531[1:1]};
assign col_out_533 = {u_ca_out_533[0:0], u_ca_out_532[1:1]};
assign col_out_534 = {u_ca_out_534[0:0], u_ca_out_533[1:1]};
assign col_out_535 = {u_ca_out_535[0:0], u_ca_out_534[1:1]};
assign col_out_536 = {u_ca_out_536[0:0], u_ca_out_535[1:1]};
assign col_out_537 = {u_ca_out_537[0:0], u_ca_out_536[1:1]};
assign col_out_538 = {u_ca_out_538[0:0], u_ca_out_537[1:1]};
assign col_out_539 = {u_ca_out_539[0:0], u_ca_out_538[1:1]};
assign col_out_540 = {u_ca_out_540[0:0], u_ca_out_539[1:1]};
assign col_out_541 = {u_ca_out_541[0:0], u_ca_out_540[1:1]};
assign col_out_542 = {u_ca_out_542[0:0], u_ca_out_541[1:1]};
assign col_out_543 = {u_ca_out_543[0:0], u_ca_out_542[1:1]};
assign col_out_544 = {u_ca_out_544[0:0], u_ca_out_543[1:1]};
assign col_out_545 = {u_ca_out_545[0:0], u_ca_out_544[1:1]};
assign col_out_546 = {u_ca_out_546[0:0], u_ca_out_545[1:1]};
assign col_out_547 = {u_ca_out_547[0:0], u_ca_out_546[1:1]};
assign col_out_548 = {u_ca_out_548[0:0], u_ca_out_547[1:1]};
assign col_out_549 = {u_ca_out_549[0:0], u_ca_out_548[1:1]};
assign col_out_550 = {u_ca_out_550[0:0], u_ca_out_549[1:1]};
assign col_out_551 = {u_ca_out_551[0:0], u_ca_out_550[1:1]};
assign col_out_552 = {u_ca_out_552[0:0], u_ca_out_551[1:1]};
assign col_out_553 = {u_ca_out_553[0:0], u_ca_out_552[1:1]};
assign col_out_554 = {u_ca_out_554[0:0], u_ca_out_553[1:1]};
assign col_out_555 = {u_ca_out_555[0:0], u_ca_out_554[1:1]};
assign col_out_556 = {u_ca_out_556[0:0], u_ca_out_555[1:1]};
assign col_out_557 = {u_ca_out_557[0:0], u_ca_out_556[1:1]};
assign col_out_558 = {u_ca_out_558[0:0], u_ca_out_557[1:1]};
assign col_out_559 = {u_ca_out_559[0:0], u_ca_out_558[1:1]};
assign col_out_560 = {u_ca_out_560[0:0], u_ca_out_559[1:1]};
assign col_out_561 = {u_ca_out_561[0:0], u_ca_out_560[1:1]};
assign col_out_562 = {u_ca_out_562[0:0], u_ca_out_561[1:1]};
assign col_out_563 = {u_ca_out_563[0:0], u_ca_out_562[1:1]};
assign col_out_564 = {u_ca_out_564[0:0], u_ca_out_563[1:1]};
assign col_out_565 = {u_ca_out_565[0:0], u_ca_out_564[1:1]};
assign col_out_566 = {u_ca_out_566[0:0], u_ca_out_565[1:1]};
assign col_out_567 = {u_ca_out_567[0:0], u_ca_out_566[1:1]};
assign col_out_568 = {u_ca_out_568[0:0], u_ca_out_567[1:1]};
assign col_out_569 = {u_ca_out_569[0:0], u_ca_out_568[1:1]};
assign col_out_570 = {u_ca_out_570[0:0], u_ca_out_569[1:1]};
assign col_out_571 = {u_ca_out_571[0:0], u_ca_out_570[1:1]};
assign col_out_572 = {u_ca_out_572[0:0], u_ca_out_571[1:1]};
assign col_out_573 = {u_ca_out_573[0:0], u_ca_out_572[1:1]};
assign col_out_574 = {u_ca_out_574[0:0], u_ca_out_573[1:1]};
assign col_out_575 = {u_ca_out_575[0:0], u_ca_out_574[1:1]};
assign col_out_576 = {u_ca_out_576[0:0], u_ca_out_575[1:1]};
assign col_out_577 = {u_ca_out_577[0:0], u_ca_out_576[1:1]};
assign col_out_578 = {u_ca_out_578[0:0], u_ca_out_577[1:1]};
assign col_out_579 = {u_ca_out_579[0:0], u_ca_out_578[1:1]};
assign col_out_580 = {u_ca_out_580[0:0], u_ca_out_579[1:1]};
assign col_out_581 = {u_ca_out_581[0:0], u_ca_out_580[1:1]};
assign col_out_582 = {u_ca_out_582[0:0], u_ca_out_581[1:1]};
assign col_out_583 = {u_ca_out_583[0:0], u_ca_out_582[1:1]};
assign col_out_584 = {u_ca_out_584[0:0], u_ca_out_583[1:1]};
assign col_out_585 = {u_ca_out_585[0:0], u_ca_out_584[1:1]};
assign col_out_586 = {u_ca_out_586[0:0], u_ca_out_585[1:1]};
assign col_out_587 = {u_ca_out_587[0:0], u_ca_out_586[1:1]};
assign col_out_588 = {u_ca_out_588[0:0], u_ca_out_587[1:1]};
assign col_out_589 = {u_ca_out_589[0:0], u_ca_out_588[1:1]};
assign col_out_590 = {u_ca_out_590[0:0], u_ca_out_589[1:1]};
assign col_out_591 = {u_ca_out_591[0:0], u_ca_out_590[1:1]};
assign col_out_592 = {u_ca_out_592[0:0], u_ca_out_591[1:1]};
assign col_out_593 = {u_ca_out_593[0:0], u_ca_out_592[1:1]};
assign col_out_594 = {u_ca_out_594[0:0], u_ca_out_593[1:1]};
assign col_out_595 = {u_ca_out_595[0:0], u_ca_out_594[1:1]};
assign col_out_596 = {u_ca_out_596[0:0], u_ca_out_595[1:1]};
assign col_out_597 = {u_ca_out_597[0:0], u_ca_out_596[1:1]};
assign col_out_598 = {u_ca_out_598[0:0], u_ca_out_597[1:1]};
assign col_out_599 = {u_ca_out_599[0:0], u_ca_out_598[1:1]};
assign col_out_600 = {u_ca_out_600[0:0], u_ca_out_599[1:1]};
assign col_out_601 = {u_ca_out_601[0:0], u_ca_out_600[1:1]};
assign col_out_602 = {u_ca_out_602[0:0], u_ca_out_601[1:1]};
assign col_out_603 = {u_ca_out_603[0:0], u_ca_out_602[1:1]};
assign col_out_604 = {u_ca_out_604[0:0], u_ca_out_603[1:1]};
assign col_out_605 = {u_ca_out_605[0:0], u_ca_out_604[1:1]};
assign col_out_606 = {u_ca_out_606[0:0], u_ca_out_605[1:1]};
assign col_out_607 = {u_ca_out_607[0:0], u_ca_out_606[1:1]};
assign col_out_608 = {u_ca_out_608[0:0], u_ca_out_607[1:1]};
assign col_out_609 = {u_ca_out_609[0:0], u_ca_out_608[1:1]};
assign col_out_610 = {u_ca_out_610[0:0], u_ca_out_609[1:1]};
assign col_out_611 = {u_ca_out_611[0:0], u_ca_out_610[1:1]};
assign col_out_612 = {u_ca_out_612[0:0], u_ca_out_611[1:1]};
assign col_out_613 = {u_ca_out_613[0:0], u_ca_out_612[1:1]};
assign col_out_614 = {u_ca_out_614[0:0], u_ca_out_613[1:1]};
assign col_out_615 = {u_ca_out_615[0:0], u_ca_out_614[1:1]};
assign col_out_616 = {u_ca_out_616[0:0], u_ca_out_615[1:1]};
assign col_out_617 = {u_ca_out_617[0:0], u_ca_out_616[1:1]};
assign col_out_618 = {u_ca_out_618[0:0], u_ca_out_617[1:1]};
assign col_out_619 = {u_ca_out_619[0:0], u_ca_out_618[1:1]};
assign col_out_620 = {u_ca_out_620[0:0], u_ca_out_619[1:1]};
assign col_out_621 = {u_ca_out_621[0:0], u_ca_out_620[1:1]};
assign col_out_622 = {u_ca_out_622[0:0], u_ca_out_621[1:1]};
assign col_out_623 = {u_ca_out_623[0:0], u_ca_out_622[1:1]};
assign col_out_624 = {u_ca_out_624[0:0], u_ca_out_623[1:1]};
assign col_out_625 = {u_ca_out_625[0:0], u_ca_out_624[1:1]};
assign col_out_626 = {u_ca_out_626[0:0], u_ca_out_625[1:1]};
assign col_out_627 = {u_ca_out_627[0:0], u_ca_out_626[1:1]};
assign col_out_628 = {u_ca_out_628[0:0], u_ca_out_627[1:1]};
assign col_out_629 = {u_ca_out_629[0:0], u_ca_out_628[1:1]};
assign col_out_630 = {u_ca_out_630[0:0], u_ca_out_629[1:1]};
assign col_out_631 = {u_ca_out_631[0:0], u_ca_out_630[1:1]};
assign col_out_632 = {u_ca_out_632[0:0], u_ca_out_631[1:1]};
assign col_out_633 = {u_ca_out_633[0:0], u_ca_out_632[1:1]};
assign col_out_634 = {u_ca_out_634[0:0], u_ca_out_633[1:1]};
assign col_out_635 = {u_ca_out_635[0:0], u_ca_out_634[1:1]};
assign col_out_636 = {u_ca_out_636[0:0], u_ca_out_635[1:1]};
assign col_out_637 = {u_ca_out_637[0:0], u_ca_out_636[1:1]};
assign col_out_638 = {u_ca_out_638[0:0], u_ca_out_637[1:1]};
assign col_out_639 = {u_ca_out_639[0:0], u_ca_out_638[1:1]};
assign col_out_640 = {u_ca_out_640[0:0], u_ca_out_639[1:1]};
assign col_out_641 = {u_ca_out_641[0:0], u_ca_out_640[1:1]};
assign col_out_642 = {u_ca_out_642[0:0], u_ca_out_641[1:1]};
assign col_out_643 = {u_ca_out_643[0:0], u_ca_out_642[1:1]};
assign col_out_644 = {u_ca_out_644[0:0], u_ca_out_643[1:1]};
assign col_out_645 = {u_ca_out_645[0:0], u_ca_out_644[1:1]};
assign col_out_646 = {u_ca_out_646[0:0], u_ca_out_645[1:1]};
assign col_out_647 = {u_ca_out_647[0:0], u_ca_out_646[1:1]};
assign col_out_648 = {u_ca_out_648[0:0], u_ca_out_647[1:1]};
assign col_out_649 = {u_ca_out_649[0:0], u_ca_out_648[1:1]};
assign col_out_650 = {u_ca_out_650[0:0], u_ca_out_649[1:1]};
assign col_out_651 = {u_ca_out_651[0:0], u_ca_out_650[1:1]};
assign col_out_652 = {u_ca_out_652[0:0], u_ca_out_651[1:1]};
assign col_out_653 = {u_ca_out_653[0:0], u_ca_out_652[1:1]};
assign col_out_654 = {u_ca_out_654[0:0], u_ca_out_653[1:1]};
assign col_out_655 = {u_ca_out_655[0:0], u_ca_out_654[1:1]};
assign col_out_656 = {u_ca_out_656[0:0], u_ca_out_655[1:1]};
assign col_out_657 = {u_ca_out_657[0:0], u_ca_out_656[1:1]};
assign col_out_658 = {u_ca_out_658[0:0], u_ca_out_657[1:1]};
assign col_out_659 = {u_ca_out_659[0:0], u_ca_out_658[1:1]};
assign col_out_660 = {u_ca_out_660[0:0], u_ca_out_659[1:1]};
assign col_out_661 = {u_ca_out_661[0:0], u_ca_out_660[1:1]};
assign col_out_662 = {u_ca_out_662[0:0], u_ca_out_661[1:1]};
assign col_out_663 = {u_ca_out_663[0:0], u_ca_out_662[1:1]};
assign col_out_664 = {u_ca_out_664[0:0], u_ca_out_663[1:1]};
assign col_out_665 = {u_ca_out_665[0:0], u_ca_out_664[1:1]};
assign col_out_666 = {u_ca_out_666[0:0], u_ca_out_665[1:1]};
assign col_out_667 = {u_ca_out_667[0:0], u_ca_out_666[1:1]};
assign col_out_668 = {u_ca_out_668[0:0], u_ca_out_667[1:1]};
assign col_out_669 = {u_ca_out_669[0:0], u_ca_out_668[1:1]};
assign col_out_670 = {u_ca_out_670[0:0], u_ca_out_669[1:1]};
assign col_out_671 = {u_ca_out_671[0:0], u_ca_out_670[1:1]};
assign col_out_672 = {u_ca_out_672[0:0], u_ca_out_671[1:1]};
assign col_out_673 = {u_ca_out_673[0:0], u_ca_out_672[1:1]};
assign col_out_674 = {u_ca_out_674[0:0], u_ca_out_673[1:1]};
assign col_out_675 = {u_ca_out_675[0:0], u_ca_out_674[1:1]};
assign col_out_676 = {u_ca_out_676[0:0], u_ca_out_675[1:1]};
assign col_out_677 = {u_ca_out_677[0:0], u_ca_out_676[1:1]};
assign col_out_678 = {u_ca_out_678[0:0], u_ca_out_677[1:1]};
assign col_out_679 = {u_ca_out_679[0:0], u_ca_out_678[1:1]};
assign col_out_680 = {u_ca_out_680[0:0], u_ca_out_679[1:1]};
assign col_out_681 = {u_ca_out_681[0:0], u_ca_out_680[1:1]};
assign col_out_682 = {u_ca_out_682[0:0], u_ca_out_681[1:1]};
assign col_out_683 = {u_ca_out_683[0:0], u_ca_out_682[1:1]};
assign col_out_684 = {u_ca_out_684[0:0], u_ca_out_683[1:1]};
assign col_out_685 = {u_ca_out_685[0:0], u_ca_out_684[1:1]};
assign col_out_686 = {u_ca_out_686[0:0], u_ca_out_685[1:1]};
assign col_out_687 = {u_ca_out_687[0:0], u_ca_out_686[1:1]};
assign col_out_688 = {u_ca_out_688[0:0], u_ca_out_687[1:1]};
assign col_out_689 = {u_ca_out_689[0:0], u_ca_out_688[1:1]};
assign col_out_690 = {u_ca_out_690[0:0], u_ca_out_689[1:1]};
assign col_out_691 = {u_ca_out_691[0:0], u_ca_out_690[1:1]};
assign col_out_692 = {u_ca_out_692[0:0], u_ca_out_691[1:1]};
assign col_out_693 = {u_ca_out_693[0:0], u_ca_out_692[1:1]};
assign col_out_694 = {u_ca_out_694[0:0], u_ca_out_693[1:1]};
assign col_out_695 = {u_ca_out_695[0:0], u_ca_out_694[1:1]};
assign col_out_696 = {u_ca_out_696[0:0], u_ca_out_695[1:1]};
assign col_out_697 = {u_ca_out_697[0:0], u_ca_out_696[1:1]};
assign col_out_698 = {u_ca_out_698[0:0], u_ca_out_697[1:1]};
assign col_out_699 = {u_ca_out_699[0:0], u_ca_out_698[1:1]};
assign col_out_700 = {u_ca_out_700[0:0], u_ca_out_699[1:1]};
assign col_out_701 = {u_ca_out_701[0:0], u_ca_out_700[1:1]};
assign col_out_702 = {u_ca_out_702[0:0], u_ca_out_701[1:1]};
assign col_out_703 = {u_ca_out_703[0:0], u_ca_out_702[1:1]};
assign col_out_704 = {u_ca_out_704[0:0], u_ca_out_703[1:1]};
assign col_out_705 = {u_ca_out_705[0:0], u_ca_out_704[1:1]};
assign col_out_706 = {u_ca_out_706[0:0], u_ca_out_705[1:1]};
assign col_out_707 = {u_ca_out_707[0:0], u_ca_out_706[1:1]};
assign col_out_708 = {u_ca_out_708[0:0], u_ca_out_707[1:1]};
assign col_out_709 = {u_ca_out_709[0:0], u_ca_out_708[1:1]};
assign col_out_710 = {u_ca_out_710[0:0], u_ca_out_709[1:1]};
assign col_out_711 = {u_ca_out_711[0:0], u_ca_out_710[1:1]};
assign col_out_712 = {u_ca_out_712[0:0], u_ca_out_711[1:1]};
assign col_out_713 = {u_ca_out_713[0:0], u_ca_out_712[1:1]};
assign col_out_714 = {u_ca_out_714[0:0], u_ca_out_713[1:1]};
assign col_out_715 = {u_ca_out_715[0:0], u_ca_out_714[1:1]};
assign col_out_716 = {u_ca_out_716[0:0], u_ca_out_715[1:1]};
assign col_out_717 = {u_ca_out_717[0:0], u_ca_out_716[1:1]};
assign col_out_718 = {u_ca_out_718[0:0], u_ca_out_717[1:1]};
assign col_out_719 = {u_ca_out_719[0:0], u_ca_out_718[1:1]};
assign col_out_720 = {u_ca_out_720[0:0], u_ca_out_719[1:1]};
assign col_out_721 = {u_ca_out_721[0:0], u_ca_out_720[1:1]};
assign col_out_722 = {u_ca_out_722[0:0], u_ca_out_721[1:1]};
assign col_out_723 = {u_ca_out_723[0:0], u_ca_out_722[1:1]};
assign col_out_724 = {u_ca_out_724[0:0], u_ca_out_723[1:1]};
assign col_out_725 = {u_ca_out_725[0:0], u_ca_out_724[1:1]};
assign col_out_726 = {u_ca_out_726[0:0], u_ca_out_725[1:1]};
assign col_out_727 = {u_ca_out_727[0:0], u_ca_out_726[1:1]};
assign col_out_728 = {u_ca_out_728[0:0], u_ca_out_727[1:1]};
assign col_out_729 = {u_ca_out_729[0:0], u_ca_out_728[1:1]};
assign col_out_730 = {u_ca_out_730[0:0], u_ca_out_729[1:1]};
assign col_out_731 = {u_ca_out_731[0:0], u_ca_out_730[1:1]};
assign col_out_732 = {u_ca_out_732[0:0], u_ca_out_731[1:1]};
assign col_out_733 = {u_ca_out_733[0:0], u_ca_out_732[1:1]};
assign col_out_734 = {u_ca_out_734[0:0], u_ca_out_733[1:1]};
assign col_out_735 = {u_ca_out_735[0:0], u_ca_out_734[1:1]};
assign col_out_736 = {u_ca_out_736[0:0], u_ca_out_735[1:1]};
assign col_out_737 = {u_ca_out_737[0:0], u_ca_out_736[1:1]};
assign col_out_738 = {u_ca_out_738[0:0], u_ca_out_737[1:1]};
assign col_out_739 = {u_ca_out_739[0:0], u_ca_out_738[1:1]};
assign col_out_740 = {u_ca_out_740[0:0], u_ca_out_739[1:1]};
assign col_out_741 = {u_ca_out_741[0:0], u_ca_out_740[1:1]};
assign col_out_742 = {u_ca_out_742[0:0], u_ca_out_741[1:1]};
assign col_out_743 = {u_ca_out_743[0:0], u_ca_out_742[1:1]};
assign col_out_744 = {u_ca_out_744[0:0], u_ca_out_743[1:1]};
assign col_out_745 = {u_ca_out_745[0:0], u_ca_out_744[1:1]};
assign col_out_746 = {u_ca_out_746[0:0], u_ca_out_745[1:1]};
assign col_out_747 = {u_ca_out_747[0:0], u_ca_out_746[1:1]};
assign col_out_748 = {u_ca_out_748[0:0], u_ca_out_747[1:1]};
assign col_out_749 = {u_ca_out_749[0:0], u_ca_out_748[1:1]};
assign col_out_750 = {u_ca_out_750[0:0], u_ca_out_749[1:1]};
assign col_out_751 = {u_ca_out_751[0:0], u_ca_out_750[1:1]};
assign col_out_752 = {u_ca_out_752[0:0], u_ca_out_751[1:1]};
assign col_out_753 = {u_ca_out_753[0:0], u_ca_out_752[1:1]};
assign col_out_754 = {u_ca_out_754[0:0], u_ca_out_753[1:1]};
assign col_out_755 = {u_ca_out_755[0:0], u_ca_out_754[1:1]};
assign col_out_756 = {u_ca_out_756[0:0], u_ca_out_755[1:1]};
assign col_out_757 = {u_ca_out_757[0:0], u_ca_out_756[1:1]};
assign col_out_758 = {u_ca_out_758[0:0], u_ca_out_757[1:1]};
assign col_out_759 = {u_ca_out_759[0:0], u_ca_out_758[1:1]};
assign col_out_760 = {u_ca_out_760[0:0], u_ca_out_759[1:1]};
assign col_out_761 = {u_ca_out_761[0:0], u_ca_out_760[1:1]};
assign col_out_762 = {u_ca_out_762[0:0], u_ca_out_761[1:1]};
assign col_out_763 = {u_ca_out_763[0:0], u_ca_out_762[1:1]};
assign col_out_764 = {u_ca_out_764[0:0], u_ca_out_763[1:1]};
assign col_out_765 = {u_ca_out_765[0:0], u_ca_out_764[1:1]};
assign col_out_766 = {u_ca_out_766[0:0], u_ca_out_765[1:1]};
assign col_out_767 = {u_ca_out_767[0:0], u_ca_out_766[1:1]};
assign col_out_768 = {u_ca_out_768[0:0], u_ca_out_767[1:1]};
assign col_out_769 = {u_ca_out_769[0:0], u_ca_out_768[1:1]};
assign col_out_770 = {u_ca_out_770[0:0], u_ca_out_769[1:1]};
assign col_out_771 = {u_ca_out_771[0:0], u_ca_out_770[1:1]};
assign col_out_772 = {u_ca_out_772[0:0], u_ca_out_771[1:1]};
assign col_out_773 = {u_ca_out_773[0:0], u_ca_out_772[1:1]};
assign col_out_774 = {u_ca_out_774[0:0], u_ca_out_773[1:1]};
assign col_out_775 = {u_ca_out_775[0:0], u_ca_out_774[1:1]};
assign col_out_776 = {u_ca_out_776[0:0], u_ca_out_775[1:1]};
assign col_out_777 = {u_ca_out_777[0:0], u_ca_out_776[1:1]};
assign col_out_778 = {u_ca_out_778[0:0], u_ca_out_777[1:1]};
assign col_out_779 = {u_ca_out_779[0:0], u_ca_out_778[1:1]};
assign col_out_780 = {u_ca_out_780[0:0], u_ca_out_779[1:1]};
assign col_out_781 = {u_ca_out_781[0:0], u_ca_out_780[1:1]};
assign col_out_782 = {u_ca_out_782[0:0], u_ca_out_781[1:1]};
assign col_out_783 = {u_ca_out_783[0:0], u_ca_out_782[1:1]};
assign col_out_784 = {u_ca_out_784[0:0], u_ca_out_783[1:1]};
assign col_out_785 = {u_ca_out_785[0:0], u_ca_out_784[1:1]};
assign col_out_786 = {u_ca_out_786[0:0], u_ca_out_785[1:1]};
assign col_out_787 = {u_ca_out_787[0:0], u_ca_out_786[1:1]};
assign col_out_788 = {u_ca_out_788[0:0], u_ca_out_787[1:1]};
assign col_out_789 = {u_ca_out_789[0:0], u_ca_out_788[1:1]};
assign col_out_790 = {u_ca_out_790[0:0], u_ca_out_789[1:1]};
assign col_out_791 = {u_ca_out_791[0:0], u_ca_out_790[1:1]};
assign col_out_792 = {u_ca_out_792[0:0], u_ca_out_791[1:1]};
assign col_out_793 = {u_ca_out_793[0:0], u_ca_out_792[1:1]};
assign col_out_794 = {u_ca_out_794[0:0], u_ca_out_793[1:1]};
assign col_out_795 = {u_ca_out_795[0:0], u_ca_out_794[1:1]};
assign col_out_796 = {u_ca_out_796[0:0], u_ca_out_795[1:1]};
assign col_out_797 = {u_ca_out_797[0:0], u_ca_out_796[1:1]};
assign col_out_798 = {u_ca_out_798[0:0], u_ca_out_797[1:1]};
assign col_out_799 = {u_ca_out_799[0:0], u_ca_out_798[1:1]};
assign col_out_800 = {u_ca_out_800[0:0], u_ca_out_799[1:1]};
assign col_out_801 = {u_ca_out_801[0:0], u_ca_out_800[1:1]};
assign col_out_802 = {u_ca_out_802[0:0], u_ca_out_801[1:1]};
assign col_out_803 = {u_ca_out_803[0:0], u_ca_out_802[1:1]};
assign col_out_804 = {u_ca_out_804[0:0], u_ca_out_803[1:1]};
assign col_out_805 = {u_ca_out_805[0:0], u_ca_out_804[1:1]};
assign col_out_806 = {u_ca_out_806[0:0], u_ca_out_805[1:1]};
assign col_out_807 = {u_ca_out_807[0:0], u_ca_out_806[1:1]};
assign col_out_808 = {u_ca_out_808[0:0], u_ca_out_807[1:1]};
assign col_out_809 = {u_ca_out_809[0:0], u_ca_out_808[1:1]};
assign col_out_810 = {u_ca_out_810[0:0], u_ca_out_809[1:1]};
assign col_out_811 = {u_ca_out_811[0:0], u_ca_out_810[1:1]};
assign col_out_812 = {u_ca_out_812[0:0], u_ca_out_811[1:1]};
assign col_out_813 = {u_ca_out_813[0:0], u_ca_out_812[1:1]};
assign col_out_814 = {u_ca_out_814[0:0], u_ca_out_813[1:1]};
assign col_out_815 = {u_ca_out_815[0:0], u_ca_out_814[1:1]};
assign col_out_816 = {u_ca_out_816[0:0], u_ca_out_815[1:1]};
assign col_out_817 = {u_ca_out_817[0:0], u_ca_out_816[1:1]};
assign col_out_818 = {u_ca_out_818[0:0], u_ca_out_817[1:1]};
assign col_out_819 = {u_ca_out_819[0:0], u_ca_out_818[1:1]};
assign col_out_820 = {u_ca_out_820[0:0], u_ca_out_819[1:1]};
assign col_out_821 = {u_ca_out_821[0:0], u_ca_out_820[1:1]};
assign col_out_822 = {u_ca_out_822[0:0], u_ca_out_821[1:1]};
assign col_out_823 = {u_ca_out_823[0:0], u_ca_out_822[1:1]};
assign col_out_824 = {u_ca_out_824[0:0], u_ca_out_823[1:1]};
assign col_out_825 = {u_ca_out_825[0:0], u_ca_out_824[1:1]};
assign col_out_826 = {u_ca_out_826[0:0], u_ca_out_825[1:1]};
assign col_out_827 = {u_ca_out_827[0:0], u_ca_out_826[1:1]};
assign col_out_828 = {u_ca_out_828[0:0], u_ca_out_827[1:1]};
assign col_out_829 = {u_ca_out_829[0:0], u_ca_out_828[1:1]};
assign col_out_830 = {u_ca_out_830[0:0], u_ca_out_829[1:1]};
assign col_out_831 = {u_ca_out_831[0:0], u_ca_out_830[1:1]};
assign col_out_832 = {u_ca_out_832[0:0], u_ca_out_831[1:1]};
assign col_out_833 = {u_ca_out_833[0:0], u_ca_out_832[1:1]};
assign col_out_834 = {u_ca_out_834[0:0], u_ca_out_833[1:1]};
assign col_out_835 = {u_ca_out_835[0:0], u_ca_out_834[1:1]};
assign col_out_836 = {u_ca_out_836[0:0], u_ca_out_835[1:1]};
assign col_out_837 = {u_ca_out_837[0:0], u_ca_out_836[1:1]};
assign col_out_838 = {u_ca_out_838[0:0], u_ca_out_837[1:1]};
assign col_out_839 = {u_ca_out_839[0:0], u_ca_out_838[1:1]};
assign col_out_840 = {u_ca_out_840[0:0], u_ca_out_839[1:1]};
assign col_out_841 = {u_ca_out_841[0:0], u_ca_out_840[1:1]};
assign col_out_842 = {u_ca_out_842[0:0], u_ca_out_841[1:1]};
assign col_out_843 = {u_ca_out_843[0:0], u_ca_out_842[1:1]};
assign col_out_844 = {u_ca_out_844[0:0], u_ca_out_843[1:1]};
assign col_out_845 = {u_ca_out_845[0:0], u_ca_out_844[1:1]};
assign col_out_846 = {u_ca_out_846[0:0], u_ca_out_845[1:1]};
assign col_out_847 = {u_ca_out_847[0:0], u_ca_out_846[1:1]};
assign col_out_848 = {u_ca_out_848[0:0], u_ca_out_847[1:1]};
assign col_out_849 = {u_ca_out_849[0:0], u_ca_out_848[1:1]};
assign col_out_850 = {u_ca_out_850[0:0], u_ca_out_849[1:1]};
assign col_out_851 = {u_ca_out_851[0:0], u_ca_out_850[1:1]};
assign col_out_852 = {u_ca_out_852[0:0], u_ca_out_851[1:1]};
assign col_out_853 = {u_ca_out_853[0:0], u_ca_out_852[1:1]};
assign col_out_854 = {u_ca_out_854[0:0], u_ca_out_853[1:1]};
assign col_out_855 = {u_ca_out_855[0:0], u_ca_out_854[1:1]};
assign col_out_856 = {u_ca_out_856[0:0], u_ca_out_855[1:1]};
assign col_out_857 = {u_ca_out_857[0:0], u_ca_out_856[1:1]};
assign col_out_858 = {u_ca_out_858[0:0], u_ca_out_857[1:1]};
assign col_out_859 = {u_ca_out_859[0:0], u_ca_out_858[1:1]};
assign col_out_860 = {u_ca_out_860[0:0], u_ca_out_859[1:1]};
assign col_out_861 = {u_ca_out_861[0:0], u_ca_out_860[1:1]};
assign col_out_862 = {u_ca_out_862[0:0], u_ca_out_861[1:1]};
assign col_out_863 = {u_ca_out_863[0:0], u_ca_out_862[1:1]};
assign col_out_864 = {u_ca_out_864[0:0], u_ca_out_863[1:1]};
assign col_out_865 = {u_ca_out_865[0:0], u_ca_out_864[1:1]};
assign col_out_866 = {u_ca_out_866[0:0], u_ca_out_865[1:1]};
assign col_out_867 = {u_ca_out_867[0:0], u_ca_out_866[1:1]};
assign col_out_868 = {u_ca_out_868[0:0], u_ca_out_867[1:1]};
assign col_out_869 = {u_ca_out_869[0:0], u_ca_out_868[1:1]};
assign col_out_870 = {u_ca_out_870[0:0], u_ca_out_869[1:1]};
assign col_out_871 = {u_ca_out_871[0:0], u_ca_out_870[1:1]};
assign col_out_872 = {u_ca_out_872[0:0], u_ca_out_871[1:1]};
assign col_out_873 = {u_ca_out_873[0:0], u_ca_out_872[1:1]};
assign col_out_874 = {u_ca_out_874[0:0], u_ca_out_873[1:1]};
assign col_out_875 = {u_ca_out_875[0:0], u_ca_out_874[1:1]};
assign col_out_876 = {u_ca_out_876[0:0], u_ca_out_875[1:1]};
assign col_out_877 = {u_ca_out_877[0:0], u_ca_out_876[1:1]};
assign col_out_878 = {u_ca_out_878[0:0], u_ca_out_877[1:1]};
assign col_out_879 = {u_ca_out_879[0:0], u_ca_out_878[1:1]};
assign col_out_880 = {u_ca_out_880[0:0], u_ca_out_879[1:1]};
assign col_out_881 = {u_ca_out_881[0:0], u_ca_out_880[1:1]};
assign col_out_882 = {u_ca_out_882[0:0], u_ca_out_881[1:1]};
assign col_out_883 = {u_ca_out_883[0:0], u_ca_out_882[1:1]};
assign col_out_884 = {u_ca_out_884[0:0], u_ca_out_883[1:1]};
assign col_out_885 = {u_ca_out_885[0:0], u_ca_out_884[1:1]};
assign col_out_886 = {u_ca_out_886[0:0], u_ca_out_885[1:1]};
assign col_out_887 = {u_ca_out_887[0:0], u_ca_out_886[1:1]};
assign col_out_888 = {u_ca_out_888[0:0], u_ca_out_887[1:1]};
assign col_out_889 = {u_ca_out_889[0:0], u_ca_out_888[1:1]};
assign col_out_890 = {u_ca_out_890[0:0], u_ca_out_889[1:1]};
assign col_out_891 = {u_ca_out_891[0:0], u_ca_out_890[1:1]};
assign col_out_892 = {u_ca_out_892[0:0], u_ca_out_891[1:1]};
assign col_out_893 = {u_ca_out_893[0:0], u_ca_out_892[1:1]};
assign col_out_894 = {u_ca_out_894[0:0], u_ca_out_893[1:1]};
assign col_out_895 = {u_ca_out_895[0:0], u_ca_out_894[1:1]};
assign col_out_896 = {u_ca_out_896[0:0], u_ca_out_895[1:1]};
assign col_out_897 = {u_ca_out_897[0:0], u_ca_out_896[1:1]};
assign col_out_898 = {u_ca_out_898[0:0], u_ca_out_897[1:1]};
assign col_out_899 = {u_ca_out_899[0:0], u_ca_out_898[1:1]};
assign col_out_900 = {u_ca_out_900[0:0], u_ca_out_899[1:1]};
assign col_out_901 = {u_ca_out_901[0:0], u_ca_out_900[1:1]};
assign col_out_902 = {u_ca_out_902[0:0], u_ca_out_901[1:1]};
assign col_out_903 = {u_ca_out_903[0:0], u_ca_out_902[1:1]};
assign col_out_904 = {u_ca_out_904[0:0], u_ca_out_903[1:1]};
assign col_out_905 = {u_ca_out_905[0:0], u_ca_out_904[1:1]};
assign col_out_906 = {u_ca_out_906[0:0], u_ca_out_905[1:1]};
assign col_out_907 = {u_ca_out_907[0:0], u_ca_out_906[1:1]};
assign col_out_908 = {u_ca_out_908[0:0], u_ca_out_907[1:1]};
assign col_out_909 = {u_ca_out_909[0:0], u_ca_out_908[1:1]};
assign col_out_910 = {u_ca_out_910[0:0], u_ca_out_909[1:1]};
assign col_out_911 = {u_ca_out_911[0:0], u_ca_out_910[1:1]};
assign col_out_912 = {u_ca_out_912[0:0], u_ca_out_911[1:1]};
assign col_out_913 = {u_ca_out_913[0:0], u_ca_out_912[1:1]};
assign col_out_914 = {u_ca_out_914[0:0], u_ca_out_913[1:1]};
assign col_out_915 = {u_ca_out_915[0:0], u_ca_out_914[1:1]};
assign col_out_916 = {u_ca_out_916[0:0], u_ca_out_915[1:1]};
assign col_out_917 = {u_ca_out_917[0:0], u_ca_out_916[1:1]};
assign col_out_918 = {u_ca_out_918[0:0], u_ca_out_917[1:1]};
assign col_out_919 = {u_ca_out_919[0:0], u_ca_out_918[1:1]};
assign col_out_920 = {u_ca_out_920[0:0], u_ca_out_919[1:1]};
assign col_out_921 = {u_ca_out_921[0:0], u_ca_out_920[1:1]};
assign col_out_922 = {u_ca_out_922[0:0], u_ca_out_921[1:1]};
assign col_out_923 = {u_ca_out_923[0:0], u_ca_out_922[1:1]};
assign col_out_924 = {u_ca_out_924[0:0], u_ca_out_923[1:1]};
assign col_out_925 = {u_ca_out_925[0:0], u_ca_out_924[1:1]};
assign col_out_926 = {u_ca_out_926[0:0], u_ca_out_925[1:1]};
assign col_out_927 = {u_ca_out_927[0:0], u_ca_out_926[1:1]};
assign col_out_928 = {u_ca_out_928[0:0], u_ca_out_927[1:1]};
assign col_out_929 = {u_ca_out_929[0:0], u_ca_out_928[1:1]};
assign col_out_930 = {u_ca_out_930[0:0], u_ca_out_929[1:1]};
assign col_out_931 = {u_ca_out_931[0:0], u_ca_out_930[1:1]};
assign col_out_932 = {u_ca_out_932[0:0], u_ca_out_931[1:1]};
assign col_out_933 = {u_ca_out_933[0:0], u_ca_out_932[1:1]};
assign col_out_934 = {u_ca_out_934[0:0], u_ca_out_933[1:1]};
assign col_out_935 = {u_ca_out_935[0:0], u_ca_out_934[1:1]};
assign col_out_936 = {u_ca_out_936[0:0], u_ca_out_935[1:1]};
assign col_out_937 = {u_ca_out_937[0:0], u_ca_out_936[1:1]};
assign col_out_938 = {u_ca_out_938[0:0], u_ca_out_937[1:1]};
assign col_out_939 = {u_ca_out_939[0:0], u_ca_out_938[1:1]};
assign col_out_940 = {u_ca_out_940[0:0], u_ca_out_939[1:1]};
assign col_out_941 = {u_ca_out_941[0:0], u_ca_out_940[1:1]};
assign col_out_942 = {u_ca_out_942[0:0], u_ca_out_941[1:1]};
assign col_out_943 = {u_ca_out_943[0:0], u_ca_out_942[1:1]};
assign col_out_944 = {u_ca_out_944[0:0], u_ca_out_943[1:1]};
assign col_out_945 = {u_ca_out_945[0:0], u_ca_out_944[1:1]};
assign col_out_946 = {u_ca_out_946[0:0], u_ca_out_945[1:1]};
assign col_out_947 = {u_ca_out_947[0:0], u_ca_out_946[1:1]};
assign col_out_948 = {u_ca_out_948[0:0], u_ca_out_947[1:1]};
assign col_out_949 = {u_ca_out_949[0:0], u_ca_out_948[1:1]};
assign col_out_950 = {u_ca_out_950[0:0], u_ca_out_949[1:1]};
assign col_out_951 = {u_ca_out_951[0:0], u_ca_out_950[1:1]};
assign col_out_952 = {u_ca_out_952[0:0], u_ca_out_951[1:1]};
assign col_out_953 = {u_ca_out_953[0:0], u_ca_out_952[1:1]};
assign col_out_954 = {u_ca_out_954[0:0], u_ca_out_953[1:1]};
assign col_out_955 = {u_ca_out_955[0:0], u_ca_out_954[1:1]};
assign col_out_956 = {u_ca_out_956[0:0], u_ca_out_955[1:1]};
assign col_out_957 = {u_ca_out_957[0:0], u_ca_out_956[1:1]};
assign col_out_958 = {u_ca_out_958[0:0], u_ca_out_957[1:1]};
assign col_out_959 = {u_ca_out_959[0:0], u_ca_out_958[1:1]};
assign col_out_960 = {u_ca_out_960[0:0], u_ca_out_959[1:1]};
assign col_out_961 = {u_ca_out_961[0:0], u_ca_out_960[1:1]};
assign col_out_962 = {u_ca_out_962[0:0], u_ca_out_961[1:1]};
assign col_out_963 = {u_ca_out_963[0:0], u_ca_out_962[1:1]};
assign col_out_964 = {u_ca_out_964[0:0], u_ca_out_963[1:1]};
assign col_out_965 = {u_ca_out_965[0:0], u_ca_out_964[1:1]};
assign col_out_966 = {u_ca_out_966[0:0], u_ca_out_965[1:1]};
assign col_out_967 = {u_ca_out_967[0:0], u_ca_out_966[1:1]};
assign col_out_968 = {u_ca_out_968[0:0], u_ca_out_967[1:1]};
assign col_out_969 = {u_ca_out_969[0:0], u_ca_out_968[1:1]};
assign col_out_970 = {u_ca_out_970[0:0], u_ca_out_969[1:1]};
assign col_out_971 = {u_ca_out_971[0:0], u_ca_out_970[1:1]};
assign col_out_972 = {u_ca_out_972[0:0], u_ca_out_971[1:1]};
assign col_out_973 = {u_ca_out_973[0:0], u_ca_out_972[1:1]};
assign col_out_974 = {u_ca_out_974[0:0], u_ca_out_973[1:1]};
assign col_out_975 = {u_ca_out_975[0:0], u_ca_out_974[1:1]};
assign col_out_976 = {u_ca_out_976[0:0], u_ca_out_975[1:1]};
assign col_out_977 = {u_ca_out_977[0:0], u_ca_out_976[1:1]};
assign col_out_978 = {u_ca_out_978[0:0], u_ca_out_977[1:1]};
assign col_out_979 = {u_ca_out_979[0:0], u_ca_out_978[1:1]};
assign col_out_980 = {u_ca_out_980[0:0], u_ca_out_979[1:1]};
assign col_out_981 = {u_ca_out_981[0:0], u_ca_out_980[1:1]};
assign col_out_982 = {u_ca_out_982[0:0], u_ca_out_981[1:1]};
assign col_out_983 = {u_ca_out_983[0:0], u_ca_out_982[1:1]};
assign col_out_984 = {u_ca_out_984[0:0], u_ca_out_983[1:1]};
assign col_out_985 = {u_ca_out_985[0:0], u_ca_out_984[1:1]};
assign col_out_986 = {u_ca_out_986[0:0], u_ca_out_985[1:1]};
assign col_out_987 = {u_ca_out_987[0:0], u_ca_out_986[1:1]};
assign col_out_988 = {u_ca_out_988[0:0], u_ca_out_987[1:1]};
assign col_out_989 = {u_ca_out_989[0:0], u_ca_out_988[1:1]};
assign col_out_990 = {u_ca_out_990[0:0], u_ca_out_989[1:1]};
assign col_out_991 = {u_ca_out_991[0:0], u_ca_out_990[1:1]};
assign col_out_992 = {u_ca_out_992[0:0], u_ca_out_991[1:1]};
assign col_out_993 = {u_ca_out_993[0:0], u_ca_out_992[1:1]};
assign col_out_994 = {u_ca_out_994[0:0], u_ca_out_993[1:1]};
assign col_out_995 = {u_ca_out_995[0:0], u_ca_out_994[1:1]};
assign col_out_996 = {u_ca_out_996[0:0], u_ca_out_995[1:1]};
assign col_out_997 = {u_ca_out_997[0:0], u_ca_out_996[1:1]};
assign col_out_998 = {u_ca_out_998[0:0], u_ca_out_997[1:1]};
assign col_out_999 = {u_ca_out_999[0:0], u_ca_out_998[1:1]};
assign col_out_1000 = {u_ca_out_1000[0:0], u_ca_out_999[1:1]};
assign col_out_1001 = {u_ca_out_1001[0:0], u_ca_out_1000[1:1]};
assign col_out_1002 = {u_ca_out_1002[0:0], u_ca_out_1001[1:1]};
assign col_out_1003 = {u_ca_out_1003[0:0], u_ca_out_1002[1:1]};
assign col_out_1004 = {u_ca_out_1004[0:0], u_ca_out_1003[1:1]};
assign col_out_1005 = {u_ca_out_1005[0:0], u_ca_out_1004[1:1]};
assign col_out_1006 = {u_ca_out_1006[0:0], u_ca_out_1005[1:1]};
assign col_out_1007 = {u_ca_out_1007[0:0], u_ca_out_1006[1:1]};
assign col_out_1008 = {u_ca_out_1008[0:0], u_ca_out_1007[1:1]};
assign col_out_1009 = {u_ca_out_1009[0:0], u_ca_out_1008[1:1]};
assign col_out_1010 = {u_ca_out_1010[0:0], u_ca_out_1009[1:1]};
assign col_out_1011 = {u_ca_out_1011[0:0], u_ca_out_1010[1:1]};
assign col_out_1012 = {u_ca_out_1012[0:0], u_ca_out_1011[1:1]};
assign col_out_1013 = {u_ca_out_1013[0:0], u_ca_out_1012[1:1]};
assign col_out_1014 = {u_ca_out_1014[0:0], u_ca_out_1013[1:1]};
assign col_out_1015 = {u_ca_out_1015[0:0], u_ca_out_1014[1:1]};
assign col_out_1016 = {u_ca_out_1016[0:0], u_ca_out_1015[1:1]};
assign col_out_1017 = {u_ca_out_1017[0:0], u_ca_out_1016[1:1]};
assign col_out_1018 = {u_ca_out_1018[0:0], u_ca_out_1017[1:1]};
assign col_out_1019 = {u_ca_out_1019[0:0], u_ca_out_1018[1:1]};
assign col_out_1020 = {u_ca_out_1020[0:0], u_ca_out_1019[1:1]};
assign col_out_1021 = {u_ca_out_1021[0:0], u_ca_out_1020[1:1]};
assign col_out_1022 = {u_ca_out_1022[0:0], u_ca_out_1021[1:1]};
assign col_out_1023 = {u_ca_out_1023[0:0], u_ca_out_1022[1:1]};
assign col_out_1024 = {{1{1'b0}}, u_ca_out_1023[1:1]};

//---------------------------------------------------------


endmodule
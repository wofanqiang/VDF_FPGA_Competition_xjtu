module xpb_5_730
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h8c3035b3abaae12befcbe1b7c9003413c0a2bbc3d959414d052b41a6119ca515fe32060a626e128d49186ee501a50b8f2c575b81368f4c25d63eb0743916b20795b8a9a8f256694175fd30f9dfc72c1cc63b3885ab24fbf64ea22c85ca5d4efa0fbc51ded585a1df55cd3099ffd160fe5abf4fad633236b7831a894d2ae71f84;
    5'b00010 : xpb = 1024'h67b3261195678d8f14924b9881a620d60fcf7456dd3ae2228c79c9f670369d23f91b8e9bfab5a68bf2d29e831fec0653f4948f1c4a6bc7fffbde218a375aef5db7221ea3351bd53dd9605f5126b2940898717772c9c3cadbe7b7c710da8ffb61f0711193fa424b3124da7a5507d29bd366a4c0787619103ebfc59795ccebd89d;
    5'b00011 : xpb = 1024'h4336166f7f2439f23958b5793a4c0d985efc2ce9e11c82f813c85246ced09531f405172d92fd3a8a9c8cce213e330118bcd1c2b75e4843da217d92a0359f2cb3d88b939d77e1413a3cc38da86d9dfbf46aa7b65fe86299c180cd619beac2a7c9d125d1491efef482f3e7c4100fd3d6a8728a314388ffe9c5fc70a5de6ef091b6;
    5'b00100 : xpb = 1024'h1eb906cd68e0e6555e1f1f59f2f1fa5aae28e57ce4fe23cd9b16da972d6a8d3feeee9fbf2b44ce894646fdbf5c79fbdd850ef6527224bfb4471d03b633e36a09f9f50897baa6ad36a026bbffb48963e03cddf54d070168a719e2fc26faf55431b1da90fe43bb9dd4c2f50dcb17d5117d7e6fa20e9be6c34d391bb42710f54acf;
    5'b00101 : xpb = 1024'haae93c81148bc7814deb0111bbf22e6e6ecba140be57651aa0421c3d3f073255ed20a5c98db2e1168f5f6ca45e1f076cb16651d3a8b40bda1d5bb42a6cfa1c118fadb240acfd16781623ecf994508ffd03192dd2b226649d688528acc552a32bc196e2dd19413fb418c23e6517a6727bd92ef1bbff18fa04bc363d743bdc6a53;
    5'b00110 : xpb = 1024'h866c2cdefe4873e472b16af274981b30bdf859d3c23905f02790a48d9da12a63e80a2e5b25fa751539199c427c66023179a3856ebc9087b442fb25406b3e5967b117273aefc2827479871b50db3bf7e8d54f6cbfd0c53383019ac337d5854f93a24ba2923dfde905e7cf88201fa7ad50e514628711ffd38bf8e14bbcdde1236c;
    5'b00111 : xpb = 1024'h61ef1d3ce80520479777d4d32d3e07f30d251266c61aa6c5aedf2cddfc3b2271e2f3b6ecbe420913e2d3cbe09aacfcf641e0b909d06d038e689a9656698296bdd2809c353287ee70dcea49a822275fd4a785abacef6402689ab05dc2e5b7fbfb8300624762ba9257b6dcd1db27a8e825f0f9d35224e6ad13358c5a057fe5dc85;
    5'b01000 : xpb = 1024'h3d720d9ad1c1ccaabc3e3eb3e5e3f4b55c51caf9c9fc479b362db52e5ad51a7fdddd3f7e56899d128c8dfb7eb8f3f7bb0a1deca4e4497f688e3a076c67c6d413f3ea112f754d5a6d404d77ff6912c7c079bbea9a0e02d14e33c5f84df5eaa86363b521fc87773ba985ea1b962faa22fafcdf441d37cd869a7237684e21ea959e;
    5'b01001 : xpb = 1024'h18f4fdf8bb7e790de104a8949e89e177ab7e838ccddde870bd7c3d7eb96f128dd8c6c80feed1311136482b1cd73af27fd25b203ff825fb42b3d97882660b116a15538629b812c669a3b0a656affe2fac4bf229872ca1a033ccdb92d9061d54cb4469e1b1ac33e4fb54f7655137ab5dd008c4b4e84ab46021aee27696c3ef4eb7;
    5'b01010 : xpb = 1024'ha52533ac67295a39d0d08a4c678a158b6c213f50a73729bdc2a77f24cb0bb7a3d6f8ce1a513f439e7f609a01d8dffe0efeb27bc12eb547688a1828f69f21c371ab0c2fd2aa692fab19add7508fc55bc9122d620cd7c69c2a1b7dbf5ed07aa3c55426339081b986daaac495eb377cbece63840495ade696d931fcffe3eed66e3b;
    5'b01011 : xpb = 1024'h80a8240a50e6069cf596f42d2030024dbb4df7e3ab18ca9349f6077529a5afb1d1e256abe986d79d291ac99ff726f8d3c6efaf5c4291c342afb79a0c9d6600c7cc75a4cced2e9ba77d1105a7d6b0c3b4e463a0f9f6656b0fb49359e9e0ad502d34daf345a676302c79d1dfa63f7df9a36f697560c0cd70606ea80e2c90db2754;
    5'b01100 : xpb = 1024'h5c2b14683aa2b3001a5d5e0dd8d5ef100a7ab076aefa6b68d1448fc5883fa7bfcccbdf3d81ce6b9bd2d4f93e156df3988f2ce2f7566e3f1cd5570b229baa3e1deddf19c72ff407a3e07433ff1d9c2ba0b699dfe7150439f54da8f474f0dffc95158fb2facb32d97e48df2961477f34787b4ee62bd3b449e7ab531c7532dfe06d;
    5'b01101 : xpb = 1024'h37ae04c6245f5f633f23c7ee917bdbd259a76909b2dc0c3e58931815e6d99fcdc7b567cf1a15ff9a7c8f28dc33b4ee5d576a16926a4abaf6faf67c3899ee7b740f488ec172b973a043d762566487938c88d01ed433a308dae6be8f000112a8fcf64472afefef82d017ec731c4f806f4d873456f6e69b236ee7fe2abdd4e49986;
    5'b01110 : xpb = 1024'h1330f5240e1c0bc663ea31cf4a21c894a8d4219cb6bdad13dfe1a066457397dbc29ef060b25d93992649587a51fbe9221fa74a2d7e2736d12095ed4e9832b8ca30b203bbb57edf9ca73a90adab72fb785b065dc15241d7c07fd4298b11455564d6f9326514ac2c21e6f9bcd75781aa229319c7c1f981fcf624a9390676e9529f;
    5'b01111 : xpb = 1024'h9f612ad7b9c6ecf253b613871321fca86976dd609016ee60e50ce20c57103cf1c0d0f66b14cba6266f61c75f53a0f4b14bfea5aeb4b682f6f6d49dc2d1496ad1c66aad64a7d548de1d37c1a78b3a279521419646fd66d3b6ce765610dba2a45ee6b58443ea31ce013cc6ed7157530b20edd9176f5cb433ada7c3c253a1d07223;
    5'b10000 : xpb = 1024'h7ae41b35a3839955787c7d67cbc7e96ab8a395f393f88f366c5b6a5cb5aa34ffbbba7efcad133a25191bf6fd71e7ef76143bd949c892fed11c740ed8cf8da827e7d4225eea9ab4da809aeffed2258f80f377d5341c05a29c678bf09bebd550c6c76a43f90eee77530bd4372c5f5445f5f9be883a6f9b0d34e46ed09c43d52b3c;
    5'b10001 : xpb = 1024'h56670b938d4045b89d42e748846dd62d07d04e8697da300bf3a9f2ad14442d0db6a4078e455ace23c2d6269b902eea3adc790ce4dc6f7aab42137feecdd1e57e093d97592d6020d6e3fe1e561910f76cc5ae14213aa4718200a18b26fc07fd2ea81f03ae33ab20a4dae180e7675580cb05a3f9058281e6bc2119dee4e5d9e455;
    5'b10010 : xpb = 1024'h31e9fbf176fcf21bc20951293d13c2ef56fd07199bbbd0e17af87afd72de251bb18d901fdda262226c905639ae75e4ffa4b6407ff04bf68567b2f104cc1622d42aa70c5370258cd347614cad5ffc5f5897e4530e5943406799b725b20c3aa99688d3c3635867c9f6a9eecaa26f56bba0118969d09568c0435dc4ed2d87de9d6e;
    5'b10011 : xpb = 1024'hd6cec4f60b99e7ee6cfbb09f5b9afb1a629bfac9f9d71b70247034dd1781d29ac7718b175e9f621164a85d7ccbcdfc46cf3741b0428725f8d52621aca5a602a4c10814db2eaf8cfaac47b04a6e7c7446a1a91fb77e20f4d32ccc03d1c6d55fe698883187d24734878fc145d7757f6751d6eda9ba84f99ca9a6ffb7629e35687;
    5'b10100 : xpb = 1024'h999d22030c647faad69b9cc1beb9e3c566cc7b7078f6b304077244f3e314c23faaa91ebbd85808ae5f62f4bcce61eb53994acf9c3ab7be856391128f03711231e1c92af6a541621120c1abfe86aef3613055ca8123070b43816eecc2e6caa4f87944d4f752aa1527cec944f777295773782e2a490b81d0821d8a84c354ca760b;
    5'b10101 : xpb = 1024'h75201260f6212c0dfb6206a2775fd087b5f934037cd853d98ec0cd4441aeba4da592a74d709f9cad091d245aeca8e618618803374e943a5f893083a501b54f8803329ff0e806ce0d8424da55cd9a5b4d028c096e41a5da291a84874df6fd516059f994ac7766be799dd68eb27f2a924884139b141e68aa095a35930bf6cf2f24;
    5'b10110 : xpb = 1024'h50a302bedfddd871202870833005bd4a0525ec9680b9f4af160f5594a048b25ba07c2fdf08e730abb2d753f90aefe0dd29c536d26270b639aecff4bafff98cde249c14eb2acc3a09e78808ad1485c338d4c2485b6044a90eb39a21d9072ffdc83aae54619c2367cb6ce3d86d872bcd1d8ff90bdf314f839096e0a15498d3e83d;
    5'b10111 : xpb = 1024'h2c25f31cc99a84d444eeda63e8abaa0c5452a529849b95849d5ddde4fee2aa699b65b870a12ec4aa5c9183972936dba1f2026a6d764d3213d46f65d0fe3dca34460589e56d91a6064aeb37045b712b24a6f887487ee377f44cafbc641762aa301b631416c0e0111d3bf122288f2d07f29bde7caa44365d17d38baf9d3ad8a156;
    5'b11000 : xpb = 1024'h7a8e37ab357313769b54444a15196cea37f5dbc887d365a24ac66355d7ca277964f4102397658a9064bb335477dd666ba3f9e088a29adedfa0ed6e6fc82078a676efedfb0571202ae4e655ba25c9310792ec6359d8246d9e5c556ef27955697fc17d3cbe59cba6f0afe6be3972e42c7a7c3ed75571d369f1036bde5dcdd5a6f;
    5'b11001 : xpb = 1024'h93d9192e5f021263598125fc6a51cae26422198061d677a729d7a7db6f19478d9481470c9be46b364f64221a4922e1f5e696f989c0b8fa13d04d875b3598b991fd27a888a2ad7b44244b96558223bf2d3f69febb48a742d034678374f1f2a5920bd425aabb225c4e60cb9c7d96ffa3c602833d22ba4f6d569351473307c479f3;
    5'b11010 : xpb = 1024'h6f5c098c48bebec67e478fdd22f7b7a4b34ed21365b8187cb126302bcdb33f9b8f6acf9e342bff34f91e51b86769dcbaaed42d24d49575edf5ecf87133dcf6e81e911d82e572e74087aec4acc90f271911a03da8674611b5cd7d1e00022551f9ec88e55fdfdf05a02fd8e6389f00de9b0e68adedcd3646ddcffc557ba9c9330c;
    5'b11011 : xpb = 1024'h4adef9ea327b6b29a30df9bddb9da467027b8aa66999b9523874b87c2c4d37a98a54582fcc739333a2d8815685b0d77f771160bfe871f1c81b8c69873221343e3ffa927d2838533ceb11f3040ffa8f04e3d67c9585e4e09b6692b88b1257fe61cd3da515049baef1fee62ff3a70219701a4e1eb8e01d20650ca763c44bcdec25;
    5'b11100 : xpb = 1024'h2661ea481c38178cc7d4639e9443912951a843396d7b5a27bfc340cc8ae72fb7853de0c164bb27324c92b0f4a3f7d2443f4e945afc4e6da2412bda9d30657194616407776afdbf394e75215b56e5f6f0b60cbb82a483af80ffa85316228aaac9adf264ca29585843cdf379aeaf03544526338f83f303f9ec4952720cedd2a53e;
    5'b11101 : xpb = 1024'h1e4daa605f4c3efec9acd7f4ce97deba0d4fbcc715cfafd4711c91ce98127c580276952fd02bb30f64ce092c23ecd09078bc7f6102ae97c66cb4bb32ea9aeea82cd7c71adc32b35b1d84fb29dd15edc8842fa6fc3227e6698bdeda132bd57318ea7247f4e1501959d00c369b7048f1a3219004f05ead37385fd80558fd75e57;
    5'b11110 : xpb = 1024'h8e151059b19fa51bdc66af3715e9b1ff6177b7904ab63c4a4c3d0ac2fb1dccdb7e596f5d5f70cdbe3f654f77c3e3d89833e3237746ba35a23d09fc2767c060f21886261aa019947727d580ac7d988af94e7e32f56e477a5ce7601a26fd1aa62b9e63765e239aa374f2cdf403b6d5f0188cd84ffc691d0a2b091809a2babe7ddb;
    5'b11111 : xpb = 1024'h699800b79b5c517f012d1917ce8f9ec1b0a470234e97dd1fd38b931359b7c4e97942f7eef7b861bce91f7f15e22ad35cfc2057125a96b17c62a96d3d66049e4839ef9b14e2df00738b38af03c483f2e520b471e28ce649428075b4b20d4d52937f18361348574cc6c1db3dbebed72aed98bdc0c77c03e3b245c317eb5cc336f4;
    endcase
end

endmodule

module xpb_5_65
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h583019cc46a450483932806bcf28fb3c63c9b96523e56544cea3630d5d897f68f6532066820e1a4c00cdea8ba869536e6184f135d43ef2a21ee9c0827b16f439a74f7d8947ded073e710111b1d5555db3f3b8c19212c1843a1ee55eb73265b793a2efb88c751b8acc50e8fc404ff207554470b9b4dc71f89c641636291349459;
    5'b00010 : xpb = 1024'hb06033988d48a090726500d79e51f678c79372ca47caca899d46c61abb12fed1eca640cd041c3498019bd51750d2a6dcc309e26ba87de5443dd38104f62de8734e9efb128fbda0e7ce2022363aaaabb67e7718324258308743dcabd6e64cb6f2745df7118ea371598a1d1f8809fe40eaa88e17369b8e3f138c82c6c5226928b2;
    5'b00011 : xpb = 1024'h57e3080f11febc0fe092096c5d20aa63b9e728fe96388f56ee0d6fd26599d132dfb0e3babc03d055630b805c15dde980c074abbb5a0a079aac1e0229367267fb819f43ed280b7416a29630aebf243d60c9adaab2d6fe1bba303e6fc79f486fd97f856070a52c3178c86bc86d172d3b36adfb43ef990a016d0c54af232abb56a0;
    5'b00100 : xpb = 1024'hb01321db58a30c5819c489d82c49a5a01db0e263ba1df49bbcb0d2dfc323509bd60404213e11eaa163d96ae7be473cef21f99cf12e48fa3ccb07c2abb1895c3528eec1766fea448a89a641c9dc79933c08e936cbf82a33fdd22cc5b3126ecb52b9b45bf96c7dea258d7a58311c2c5bac02424f8ae6d120f6d2961285bbefeaf9;
    5'b00101 : xpb = 1024'h5795f651dd5927d787f1926ceb18598b10049898088bb9690d777c976daa22fcc90ea70ef5f9865ec549162c83527f931f646640dfd51c93395243cff1cddbbd5bef0a51083817b95e1c504260f324e6541fc94c8cd01f30be8e89a3cb6a8439c4dbc5588306aa44cbc90116295b55f807af7c43e44ce3505267fae3c44218e7;
    5'b00110 : xpb = 1024'hafc6101e23fd781fc12412d8ba4154c773ce51fd2c711eaddc1adfa4cb33a265bf61c7757807a0aac61700b82bbbd30180e95776b4140f35583c04526ce4cff7033e87da5016e82d452c615d7e487ac1935b5565adfc3774607cdf8f3e90dfb2ff0ac0e14a5862f190d790da2e5a766d5bf687df321402da18a95e465576ad40;
    5'b00111 : xpb = 1024'h5748e494a8b3939f2f511b6d791008b2662208317adee37b2ce1895c75ba74c6b26c6a632fef3c682786abfcf0c715a57e5420c665a0318bc6868576ad294f7f363ed0b4e864bb5c19a26fd602c20c6bde91e7e642a222a74cdea37ff78c989a0a322a4060e12310cf2639bf3b8970b96163b4982f8fc533987b46a45dc8db2e;
    5'b01000 : xpb = 1024'haf78fe60ef57e3e768839bd9483903eec9ebc1969ec448bffb84ec69d343f42fa8bf8ac9b1fd56b42854968899306913dfd911fc39df242de57045f9284043b8dd8e4e3e30438bd000b280f1201762471dcd73ff63ce3aeaeeccf96b6ab2f413446125c92832dbbd9434c9834088912eb5aac0337d56e4bd5ebcaa06eefd6f87;
    5'b01001 : xpb = 1024'h56fbd2d7740dff66d6b0a46e0707b7d9bc3f77caed320d8d4c4b96217dcac6909bca2db769e4f27189c441cd5e3babb7dd43db4beb6b468453bac71d6884c341108e9718c8915efed5288f69a490f3f16904067ff874261ddb2ebd5c23aeacfa4f888f283ebb9bdcd28372684db78b7abb17ecec7ad2a716de8e9264f74f9d75;
    5'b01010 : xpb = 1024'haf2beca3bab24faf0fe324d9d630b31620093130111772d21aeef92edb5445f9921d4e1debf30cbd8a922c5906a4ff263ec8cc81bfaa392672a4879fe39bb77ab7de14a210702f72bc38a084c1e649cca83f929919a03e617d1d134796d5087389b78ab1060d54899792022c52b6abf00f5ef887c899c6a0a4cff5c7888431ce;
    5'b01011 : xpb = 1024'h56aec11a3f686b2e7e102d6e94ff6701125ce7645f85379f6bb5a2e685db185a8527f10ba3daa87aec01d79dcbb041ca3c3395d171365b7ce0ef08c423e03702eade5d7ca8be02a190aeaefd465fdb76f3762519ae462994697ed7384fd0c15a94def4101c9614a8d5e0ab115fe5a63c14cc2540c61588fa24a1de2590d65fbc;
    5'b01100 : xpb = 1024'haededae6860cbb76b742adda6428623d7626a0c9836a9ce43a5905f3e36497c37b7b117225e8c2c6eccfc229741995389db8870745754e1effd8c9469ef72b3c922ddb05f09cd31577bec01863b5315232b1b132cf7241d80b6d2d23c2f71cd3cf0def98e3e7cd559aef3ad564e4c6b1691330dc13dca883eae34188220af415;
    5'b01101 : xpb = 1024'h5661af5d0ac2d6f6256fb66f22f71628687a56fdd1d861b18b1fafab8deb6a246e85b45fddd05e844e3f6d6e3924d7dc9b235056f70170756e234a6adf3baac4c52e23e088eaa6444c34ce90e82ec2fc7de843b364182d0af7cef1147bf2d5bada3558f7fa708d74d93de3ba7213c0fd6e805d9511586add6ab529e62a5d2203;
    5'b01110 : xpb = 1024'hae91c9295167273e5ea236daf2201164cc441062f5bdc6f659c312b8eb74e98d64d8d4c65fde78d04f0d57f9e18e2b4afca8418ccb4063178d0d0aed5a529efe6c7da169d0c976b83344dfac058418d7bd23cfcc8544454e99bd46ffef19313414645480c1c246219e4c737e7712e172c2c769305f1f8a6730f68d48bb91b65c;
    5'b01111 : xpb = 1024'h56149d9fd61d42bdcccf3f6fb0eec54fbe97c697442b8bc3aa89bc7095fbbbee57e377b417c6148db07d033ea6996deefa130adc7ccc856dfb578c119a971e869f7dea44691749e707baee2489fdaa82085a624d19ea3081861f0af0a814ea1b1f8bbddfd84b0640dc9b1c638441dbbec83495e95c9b4cc0b0c875a6c3e3e44a;
    5'b10000 : xpb = 1024'hae44b76c1cc193060601bfdb8017c08c22617ffc6810f108792d1f7df3853b574e36981a99d42ed9b14aedca4f02c15d5b97fc12510b78101a414c9415ae12c046cd67cdb0f61a5aeecaff3fa753005d4795ee663b1648c5280d60dc1b3b459459bab9689f9cbeeda1a9ac278940fc341c7ba184aa626c4a7709d909551878a3;
    5'b10001 : xpb = 1024'h55c78be2a177ae85742ec8703ee6747714b53630b67eb5d5c9f3c9359e0c0db841413b0851bbca9712ba990f140e04015902c56202979a66888bcdb855f2924879cdb0a84943ed89c3410db82bcc920792cc80e6cfbc33f8146f24ccd436fe7b64e222c7b6257f0cdff8550c966ff68021e8ce3da7de2ea3f6dbc1675d6aa691;
    5'b10010 : xpb = 1024'hadf7a5aee81bfecdad6148dc0e0f6fb3787eef95da641b1a98972c42fb958d2137945b6ed3c9e4e31388839abc77576fba87b697d6d68d08a7758e3ad1098682211d2e319122bdfdaa511ed34921e7e2d2080cfff0e84c3bb65d7ab8475d59f49f111e507d7737b9a506e4d09b6f16f5762fd9d8f5a54e2dbd1d24c9ee9f3aea;
    5'b10011 : xpb = 1024'h557a7a256cd21a4d1b8e5170ccde239e6ad2a5ca28d1dfe7e95dd5faa61c5f822a9efe5c8bb180a074f82edf81829a13b7f27fe78862af5f15c00f5f114e060a541d770c2970912c7ec72d4bcd9b798d1d3e9f80858e376ea2bf3ea9005912dbaa3887af93fff7d8e3558db5a89e11417b9d0691f32110873cef0d27f6f168d8;
    5'b10100 : xpb = 1024'hadaa93f1b3766a9554c0d1dc9c071edace9c5f2f4cb7452cb801390803a5deeb20f21ec30dbf9aec75c6196b29ebed821977711d5ca1a20134a9cfe18c64fa43fb6cf495714f61a065d73e66eaf0cf685c7a2b99a6ba4fb244ad9494737f6e54e46783385b51b085a8641d79ad9d31b6cfe4122d40e830110330708a8825fd31;
    5'b10101 : xpb = 1024'h552d6868382c8614c2edda715ad5d2c5c0f015639b2509fa08c7e2bfae2cb14c13fcc1b0c5a736a9d735c4afeef7302616e23a6d0e2dc457a2f45105cca979cc2e6d3d70099d34cf3a4d4cdf6f6a6112a7b0be1a3b603ae5310f58852c7b273bef8eec9771da70a4e6b2c65ebacc2c02d5513ee63e63f26a830258e890782b1f;
    5'b10110 : xpb = 1024'had5d82347ed0d65cfc205add29fece0224b9cec8bf0a6f3ed76b45cd0bb630b50a4fe21747b550f5d803af3b9760839478672ba2e26cb6f9c1de118847c06e05d5bcbaf9517c0543215d5dfa8cbfb6ede6ec4a335c8c5328d2fdae709fa182b529bde820392c2951abc15622bfcb4c7829984a818c2b11f44943bc4b21acbf78;
    5'b10111 : xpb = 1024'h54e056ab0386f1dc6a4d6371e8cd81ed170d84fd0d78340c2831ef84b63d0315fd5a8504ff9cecb339735a805c6bc63875d1f4f293f8d950302892ac8804ed8e08bd03d3e9c9d871f5d36c73113948983222dcb3f1323e5bbf5f7261589d3b9c34e5517f4fb4e970ea0fff07ccfa46c42f05773a89a6d44dc915a4a929feed66;
    5'b11000 : xpb = 1024'had1070774a2b4224a37fe3ddb7f67d297ad73e62315d9950f6d5529213c6827ef3ada56b81ab06ff3a41450c04d519a6d756e6286837cbf24f12532f031be1c7b00c815d31a8a8e5dce37d8e2e8e9e73715e68cd125e569f614dc84ccbc397156f144d081706a21daf1e8ecbd1f96739834c82d5d76df3d78f57080bbb3381bf;
    5'b11001 : xpb = 1024'h549344edcee15da411acec7276c531146d2af4967fcb5e1e479bfc49be4d54dfe6b848593992a2bc9bb0f050c9e05c4ad4c1af7819c3ee48bd5cd4534360614fe30cca37c9f67c14b1598c06b308301dbc94fb4da70441d24daf8c3d84bf4ffc7a3bb6672d8f623ced6d37b0df28618588b9af8ed4e9b6310f28f069c385afad;
    5'b11010 : xpb = 1024'hacc35eba1585adec4adf6cde45ee2c50d0f4adfba3b0c363163f5f571bd6d448dd0b68bfbba0bd089c7edadc7249afb93646a0adee02e0eadc4694d5be7755898a5c47c111d54c8898699d21d05d85f8fbd08766c8305a15ef9de228f7e5ab75b46ab1eff4e11ae9b27bc774e42781fadd00bb2a22b0d5bad56a53cc54ba4406;
    5'b11011 : xpb = 1024'h544633309a3bc96bb90c757304bce03bc348642ff21e88306706090ec65da6a9d0160bad738858c5fdee86213754f25d33b169fd9f8f03414a9115f9febbd511bd5c909baa231fb76cdfab9a54d717a3470719e75cd64548dbffa619b0e1645cbf921b4f0b69db08f0ca7059f1567c46e26de7e3202c9814553c3c2a5d0c71f4;
    5'b11100 : xpb = 1024'hac764cfce0e019b3f23ef5ded3e5db7827121d951603ed7535a96c1c23e72612c6692c13f5967311febc70acdfbe45cb95365b3373cdf5e3697ad67c79d2c94b64ac0e24f201f02b53efbcb5722c6d7e8642a6007e025d8c7dedfc052407bfd5f9c116d7d2bb93b5b5d9001df6559cbc36b4f37e6df3b79e1b7d9f8cee41064d;
    5'b11101 : xpb = 1024'h53f9217365963533606bfe7392b48f631965d3c96471b242867015d3ce6df873b973cf01ad7e0ecf602c1bf1a4c9886f92a12483255a1839d7c557a0ba1748d397ac56ff8a4fc35a2865cb2df6a5ff28d179388112a848bf6a4fbff5dd0378bd04e88036e94453d4f427a903038497083c2220376b6f79f79b4f87eaf693343b;
    5'b11110 : xpb = 1024'hac293b3fac3a857b999e7edf61dd8a9f7d2f8d2e88571787551378e12bf777dcafc6ef682f8c291b60fa067d4d32dbddf42615b8f9990adbf6af1823352e3d0d3efbd488d22e93ce0f75dc4913fb550410b4c49a33d461030c3e15e15029d4363f177bbfb0960c81b93638c70883b77d90692bd2b93699816190eb4d87c7c894;
    5'b11111 : xpb = 1024'h53ac0fb630f0a0fb07cb877420ac3e8a6f834362d6c4dc54a5da2298d67e4a3da2d19255e773c4d8c269b1c2123e1e81f190df08ab252d3264f999477572bc9571fc1d636a7c66fce3ebeac19874e6ae5beb571ac87a4c35f89fd9d209258d1d4a3ee51ec71ecca0f784e1ac15b2b1c995d6588bb6b25bdae162d3ab9019f682;
    endcase
end

endmodule

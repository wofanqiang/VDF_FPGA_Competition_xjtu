module xpb_4_5
(
    input [4:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    4'b0000 : xpb = 1024'h0;
    4'b0001 : xpb = 1024'h40dd8a97273283eb8504775b0fc72f5d9ccb6d39a4812a876256b299d584e88f68f9744bad15425f5d10a1432518fba2034cd4a5c3de926643629d116e2f081d19c4889c73f27d96a85386c88882bf34271b2696bfe3e6ff60bdc4f28c56c9bb8ca3bc823be35691c98483ef78992493d4d9f3559275415357f7e52f675198c6;
    4'b0010 : xpb = 1024'h81bb152e4e6507d70a08eeb61f8e5ebb3996da734902550ec4ad6533ab09d11ed1f2e8975a2a84beba2142864a31f7440699a94b87bd24cc86c53a22dc5e103a33891138e7e4fb2d50a70d9111057e684e364d2d7fc7cdfec17b89e518ad93771947790477c6ad23930907def1324927a9b3e6ab24ea82a6afefca5ecea3318c;
    4'b0011 : xpb = 1024'h11eb5a6fb3a956f9c407ee3a1efb46c764ec447c180bdf1ea9275e77cd8c0ca637a3df6a3d19488f77d3a4828bece21ba5cc560b28e8e6e7198897d60fbaa3a5d8fe6526ac467b7ee66091b700ac796b814c7a2bb32587ed6cacbcdcead9baa076e3a35d02e10b27d5cda4ef71fb47922fb3fb1e671466c9c1783489ad1263e7;
    4'b0100 : xpb = 1024'h52c8e506dadbdae5490c65952ec2762501b7b1b5bc8d09a60b7e1111a310f535a09d53b5ea2e8aeed4e445c5b105ddbda9192ab0ecc7794d5ceb34e77de9abc2f2c2edc32038f9158eb4187f892f389fa867a0c273096eeccd6a81cf7730845c03875fdf3ec461b99f5228deea946c26048dee73f989a81d197019b91463fcad;
    4'b0101 : xpb = 1024'h93a66f9e020e5ed0ce10dcf03e89a5829e831eef610e342d6dd4c3ab7895ddc50996c8019743cd4e31f4e708d61ed95fac65ff56b0a60bb3a04dd1f8ec18b3e00c87765f942b76ac37079f4811b1f7d3cf82c75932ed55ec2e2846c203874e17902b1c617aa7b84b68d6acce632d90b9d967e1c98bfee9707167fee87bb59573;
    4'b0110 : xpb = 1024'h23d6b4df6752adf3880fdc743df68d8ec9d888f83017be3d524ebcef9b18194c6f47bed47a32911eefa7490517d9c4374b98ac1651d1cdce33112fac1f75474bb1fcca4d588cf6fdccc1236e0158f2d70298f457664b0fdad95979b9d5b37540edc746ba05c2164fab9b49dee3f68f245f67f63cce28cd9382f069135a24c7ce;
    4'b0111 : xpb = 1024'h64b43f768e8531df0d1453cf4dbdbcec66a3f631d498e8c4b4a56f89709d01dbd84133202747d37e4cb7ea483cf2bfd94ee580bc15b060347673ccbd8da44f68cbc152e9cc7f74947514aa3689dbb20b29b41aee262ef6da3a173eac620a3efc7a6b033c41a56ce1751fcdce5c8fb3b83441e992609e0ee6dae84e42c1766094;
    4'b1000 : xpb = 1024'ha591ca0db5b7b5ca9218cb2a5d84ec4a036f636b791a134c16fc22234621ea6b413aa76bd45d15dda9c88b8b620bbb7b52325561d98ef29ab9d669cefbd35785e585db864071f22b1d6830ff125e713f50cf4184e612ddd99ad5039eee6108b8070ebfbe7d88c3733ea451bdd528d84c091bdce7f313503a32e0337228c7f95a;
    4'b1001 : xpb = 1024'h35c20f4f1afc04ed4c17caae5cf1d4562ec4cd7448239d5bfb761b6768a425f2a6eb9e3eb74bd9ae677aed87a3c6a652f16502217abab4b54c99c7822f2feaf18afb2f7404d3727cb321b52502056c4283e56e83197097c846063696c08d2fe164aaea1708a321778168eece55f1d6b68f1bf15b353d345d44689d9d07372bb5;
    4'b1010 : xpb = 1024'h769f99e6422e88d8d11c42096cb903b3cb903aadeca4c7e35dccce013e290e820fe5128a64611c0dc48b8ecac8dfa1f4f4b1d6c73e99471b8ffc64939d5ef30ea4bfb81078c5f0135b753bed8a882b76ab009519d9547ec7a6c3fb894ce3f99cf14ea699448678094aed72bdce8afb4a63f5e4b0c7b275b09c6082cc6e88c47b;
    4'b1011 : xpb = 1024'h6cfdf27a772d7fb8b1b418d6c25ebbff6e5a4b6bbae51f34246c74560ab4a097596095d474fdfde823df0c70a9a8ccc93e48386dfc5093622bfc246d0bb867a4a350bfe3d277064f12ec0137a2f2679de16c2180cb238b651f52e811f1020c64eead0f1cfa0d60d8db20fce4f53f9b4e9f5f92409dc59d3ade8ecf74cf7f6d6;
    4'b1100 : xpb = 1024'h47ad69becea55be7101fb8e87bed1b1d93b111f0602f7c7aa49d79df36303298de8f7da8f465223ddf4e920a2fb3886e9731582ca3a39b9c66225f583eea8e9763f9949ab119edfb998246dc02b1e5ae0531e8aecc961fb5b2b2f373ab66ea81db8e8d740b842c9f573693bdc7ed1e48becfec799c519b2705e0d226b4498f9c;
    4'b1101 : xpb = 1024'h888af455f5d7dfd2952430438bb44a7b307c7f2a04b0a70206f42c790bb51b284788f1f4a17a649d3c5f334d54cc84109a7e2cd267822e02a984fc69ad1996b47dbe1d37250c6b9241d5cda48b34a4e22c4d0f458c7a06b51370b86637bdb43d683249f64767833120bb17ad408642dc93a9dfcf2ec6dc7a5dd8b7561b9b2862;
    4'b1110 : xpb = 1024'h18bb39975b1c2ef54f232fc78b2132875bd1e932d3ba3111eb6e25bd2e3756afad39e8c78469286dfa11954996876ee839b0d99208adf01d3c485a1ce0762a2023337124e96debe3d78f51ca7adb9fe55f633c43bfd7c0a3bea1eb5e09e9db66c5ce744ed281e135637fb4bdc14f414719a9f44270f0c09d6f612180fa0a5abd;
    4'b1111 : xpb = 1024'h5998c42e824eb2e0d427a7229ae861e4f89d566c783b5b994dc4d85703bc3f3f16335d13317e6acd5722368cbba06a8a3cfdae37cc8c82837faaf72e4ea5323d3cf7f9c15d60697a7fe2d893035e5f19867e62da7fbba7a31f5fb0509640a522527230d10e6537c72d0438ad39e865daee83e798036601f0c75906b0615bf383;
    endcase
end

endmodule

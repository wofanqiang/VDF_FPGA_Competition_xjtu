module xpb_5_640
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h66f836b8eef38ab264f733f3d01559bdea2a2be09e7d7d47edeb2fddc4fe7c8eb26a666855e73dbadf5393b15f0636b3b3de1d2d162596d000d9b2bf83298767b95da057f77cda78c4f0ba4fbd8c2c77651b3d8050604159dc6c07650b4450616af2595ae214bc870bd60442de99d79094d8ff0eba7c8a4ecccd3c390237266d;
    5'b00010 : xpb = 1024'h1d43281c1bf8e09bfee8f0108fd06c2a62de549067835a185df9a665d6fa4c15618c4f57e1a7fce71f48e81bdaae5c9d03a2127409985d5451142620cb809a1dfe6c0c013f68b7ac774771fce23c94bdd6318168143a55a3034b7ccf5c5dfe30a6dd208c1360808090ec21a6c56388f7dad81f3b24adb76d532afd6d7b8be66f;
    5'b00011 : xpb = 1024'h843b5ed50aec6b4e63e024045fe5c5e84d0880710600d7604be4d6439bf8c8a413f6b5c0378f3aa1fe9c7bcd39b49350b7802fa11fbdf42451edd8e04eaa2185b7c9ac5936e592253c382c4c9fc8c1353b4cbee8649a96fcdfb7843467a24e9211cf79e6f5753d079cc225e9a3fd60886fb11e49df2a41bc1ff839a67dc30cdc;
    5'b00100 : xpb = 1024'h3a86503837f1c137fdd1e0211fa0d854c5bca920cf06b430bbf34ccbadf4982ac3189eafc34ff9ce3e91d037b55cb93a074424e81330baa8a2284c419701343bfcd818027ed16f58ee8ee3f9c479297bac6302d02874ab460696f99eb8bbfc614dba411826c1010121d8434d8ac711efb5b03e76495b6edaa655fadaf717ccde;
    5'b00101 : xpb = 1024'ha17e86f126e54bea62c91414efb63212afe6d5016d843178a9de7ca972f314b975830518193737891de563e91462efedbb22421529565178a301ff011a2abba3b635b85a764e49d1b37f9e49820555f3117e405078d4ec9fe3030103c4004cc2b8ac9a7308d5bd882dae47906960e9804a893d8503d7f92973233713f94ef34b;
    5'b00110 : xpb = 1024'h57c9785453eaa1d3fcbad031af71447f289afdb1368a0e4919ecf33184eee44024a4ee07a4f7f6b55ddab853900b15d70ae6375c1cc917fcf33c72626281ce59fb442403be3a270565d655f6a6b5be39829484383caf00e909e2766e1519fa91f49761a43a218181b2c464f4502a9ae790885db16e092647f980f84872a3b34d;
    5'b00111 : xpb = 1024'he1469b780eff7bd96ac8c4e6f2c56eba14f2660ff8feb1989fb69b996eab3c6d3c6d6f730b8b5e19dd00cbe0bb33bc05aaa2ca3103bde814376e5c3aad8e11040528fad06260439182d0da3cb66267ff3aac8200089153230c1ebd86633a861308228d56b6d457b37da825836f44c4ed6877dddd83a53667fdeb97cebf8734f;
    5'b01000 : xpb = 1024'h750ca0706fe3826ffba3c0423f41b0a98b7952419e0d686177e699975be9305586313d5f869ff39c7d23a06f6ab972740e8849d026617551445098832e026877f9b03004fda2deb1dd1dc7f388f252f758c605a050e9568c0d2df33d7177f8c29b7482304d82020243b0869b158e23df6b607cec92b6ddb54cabf5b5ee2f99bc;
    5'b01001 : xpb = 1024'h2b5791d39ce8d85995957c5efefcc316042d7af167134531e7f5101f6de4ffdc3553264f1260b2c8bd18f4d9e661985d5e4c3f1719d43bd5948b0be476597b2e3ebe9bae458ebbe58f747fa0ada2bb3dc9dc498814c36ad5340d68a7c291a691d75f49617ecdc5fbc8c6a3fefc57d546b15f9d18fce80ad3d309b6ea678459be;
    5'b01010 : xpb = 1024'h924fc88c8bdc630bfa8cb052cf121cd3ee57a6d20590c279d5e03ffd32e37c6ae7bd8cb76847f0839c6c888b4567cf11122a5c442ff9d2a59564bea3f9830295f81c3c063d0b965e546539f06b2ee7b52ef787086523ac2f1079700ccdd5f6f34251a2bc60e28282d49ca841daf1acd746389c27b76495229fd6f32369bb802b;
    5'b01011 : xpb = 1024'h489ab9efb8e1b8f5947e6c6f8ecd2f40670bcf81ce969f4a45eeb68544df4bf196df75a6f408afafdc61dcf5c10ff4fa61ee518b236c9929e59f320541da154c3d2aa7af84f7739206bbf19d8fdf4ffba00dcaf028fdc0783758e5771eefa4c27e3c69ed922e467c59b2c5a5c1bb5e3e8c37bc542195c2412634b457e310402d;
    5'b01100 : xpb = 1024'haf92f0a8a7d543a7f975a0635ee288fe5135fb626d141c9233d9e66309ddc8804949dc0f49efed6abbb570a720162bae15cc6eb839922ff9e678e4c4c5039cb3f68848077c744e0acbacabed4d6b7c7305290870795e01d213c4ecdc2a33f523e92ec348744303036588c9e8a05535cf2110bb62dc124c8ff301f090e547669a;
    5'b01101 : xpb = 1024'h65dde20bd4da999193675c801e9d9b6ac9ea24123619f962a3e85ceb1bd99806f86bc4fed5b0ac96fbaac5119bbe5197659063ff2d04f67e36b358260d5aaf6a3b96b3b0c4602b3e7e03639a721be4b9763f4c583d38161b3aa462467b4da2f325198a79a58ec6fcea9ee74c871ee736670fdb8f464379ae795fb1c55e9c269c;
    5'b01110 : xpb = 1024'h1c28d36f01dfef7b2d59189cde58add7429e4cc1ff1fd63313f6d3732dd5678da78dadee61716bc33ba0197c17667780b55459462077bd0286edcb8755b1c22080a51f5a0c4c0872305a1b4796cc4cffe755904001122a646183d7b0cc6750c2610451aad6da8af66fb504b06de8989dad0efbbbb074a6ccffbd72f9d7f0e69e;
    5'b01111 : xpb = 1024'h83210a27f0d37a2d92504c90ae6e07952cc878a29d9d537b01e20350f2d3e41c59f81456b758a97e1af3ad2d766cae3469327673369d53d287c77e46d8db49883a02bfb203c8e2eaf54ad597545879774c70cdc051726bbe3defdf15d7aba123cbf6ab05b8ef477d7b8b08f34c82702e41e7faca6af1311bcc8aaf32da280d0b;
    5'b10000 : xpb = 1024'h396bfb8b1dd8d0172c4208ad6e291a01a57ca15266a3304b71f079d904cfb3a30919fd46431968aa5ae90197f214d41db8f66bba2a101a56d801f1a821325c3e7f112b5b4bb4c01ea7a18d447908e1bdbd8711a8154c800764cf548028c54ef307e17236ea3b0b7700a12657334c219587e71af6d5225e3a52e87067537ccd0d;
    5'b10001 : xpb = 1024'ha06432440ccc5ac991393ca13e3e73bf8fa6cd330520ad935fdba9b6c9ce3031bb8463ae9900a6653a3c9549511b0ad16cd488e74035b126d8dba467a45be3a6386ecbb343319a976c92479436950e3522a24f2865acc161413b5be534099f5472d3cb91cc4fc7fe0c772a9a11e5f9261cc01a058f9ee8891fb5aca055b3f37a;
    5'b10010 : xpb = 1024'h56af23a739d1b0b32b2af8bdfdf9862c085af5e2ce268a63cfea203edbc9ffb86aa64c9e24c165917a31e9b3ccc330babc987e2e33a877ab291617c8ecb2f65c7d7d375c8b1d77cb1ee8ff415b45767b93b893102986d5aa681ad14f85234d23aebe92c2fd9b8bf7918d47fdf8afaa8d62bf3a31f9d015a7a6136dd4cf08b37c;
    5'b10011 : xpb = 1024'hcfa150a66d7069cc51cb4dabdb49898810f1e92972c67343ff896c6edc5cf3f19c8358db08224bdba273e1e486b56a40c5c7375271b3e2f79508b2a350a0912c28ba305d30954fed13fb6ee7ff5dec204ced6f7ed60e9f38efa46b9d63cfaf2eaa959f42ee74ff116a36561df795bf4a8be5a5e640142c62c712f09485d737e;
    5'b10100 : xpb = 1024'h73f24bc355ca914f2a13e8ce8dc9f2566b394a7335a9e47c2de3c6a4b2c44bcdcc329bf606696278997ad1cfa7718d57c03a90a23d40d4ff7a2a3de9b833907a7be9435dca862f779630713e3d820b3969ea14783dc12b4d6b664e1ee1814b54559bb34f10fc0c78227969a4be1333853d97596d1e7dcd14f93e6b424a9499eb;
    5'b10101 : xpb = 1024'h2a3d3d2682cfe738c405a4eb4d8504c2e3ed7322feafc14c9df23d2cc4c01b547b5484e5922a21a4d970263a2319b3410ffe85e930b39b83ca64b14b008aa330c0f7af0712720cab488728eb6232737fdb005860019b3f969245c389329af92391867a804247d071a78f8708a4dce4ec8396799988aefa337f9c2c76c3e959ed;
    5'b10110 : xpb = 1024'h913573df71c371eb28fcd8df1d9a5e80ce179f039d2d3e948bdd6d0a89be97e32dbeeb4de8115f5fb8c3b9eb821fe9f4c3dca31646d93253cb3e640a83b42a987a554f5f09eee7240d77e33b1fbe9ff7401b95e051fb80f06eb1caee3ddf4984fc78d3db245c8cf8b3658b4b8376bc7d186f78a8432b84824c6968afc620805a;
    5'b10111 : xpb = 1024'h478065429ec8c7d4c2ee94fbdd5570ed46cbc7b366331b64fbebe3929bba6769dce0d43d73d21e8bf8b90e55fdc80fde13a0985d3a4bf8d81b78d76bcc0b3d4ebf63bb0851dac457bfce9ae8446f083db131d9c815d59539959140588ef8f75438639b0c55a850f2387ba8af6a406de45e6e98d4ad5cb1a0d2c729e43f75405c;
    5'b11000 : xpb = 1024'hae789bfb8dbc528727e5c8efad6acaab30f5f39404b098ace9d7137060b8e3f88f4b3aa5c9b95c46d80ca2075cce4691c77eb58a50718fa81c528a2b4f34c4b678c15b6049579ed084bf553801fb34b5164d17486635d69371fd47bd9a3d47b5a355f46737bd0d794451acf248da4574f34797e367d93bef9f94661d41ac66c9;
    5'b11001 : xpb = 1024'h64c38d5ebac1a870c1d7850c6d25dd17a9aa1c43cdb6757d59e589f872b4b37f3e6d2395557a1b731801f671d8766c7b1742aad143e4562c6c8cfd8c978bd76cbdcfc70991437c0437160ce526ab9cfb87635b302a0feadc98dcbd27eb56f584df40bb986908d172c967ca562fa3f6dc3946b80fd20a690e25f22751bb0126cb;
    5'b11010 : xpb = 1024'h1b0e7ec1e7c6fe5a5bc941292ce0ef84225e44f396bc524dc9f4008084b08305ed8f0c84e13ada9f57f74adc541e92646706a01837571cb0bcc770eddfe2ea2302de32b2d92f5937e96cc4924b5c0541f8799f17ede9ff25bfbc32923c70a3541b2b82c99a54956c4e7de7ba166da8437f45d83c3c3b962cac4fe8863455e6cd;
    5'b11011 : xpb = 1024'h8206b57ad6ba890cc0c0751cfcf649420c8870d43539cf95b7df305e49aeff949ff972ed3722185a374ade8db324c9181ae4bd454d7cb380bda123ad630c718abc3bd30ad0ac33b0ae5d7ee208e831b95d94dc983e4a407f9c2839f747b4f3b5861ddc247c6951f35a53ebfcf5077fd4141ed74af6b8207b791d24bf368d0d3a;
    5'b11100 : xpb = 1024'h3851a6de03bfdef65ab23139bcb15bae853c9983fe3fac6627eda6e65baacf1b4f1b5bdcc2e2d786774032f82eccef016aa8b28c40ef7a050ddb970eab638441014a3eb4189810e460b4368f2d9899ffceab2080022454c8c307af6198cea184c208a355adb515ecdf6a0960dbd1313b5a1df77760e94d99ff7ae5f3afe1cd3c;
    5'b11101 : xpb = 1024'h9f49dd96f2b369a8bfa9652d8cc6b56c6f66c5649cbd29ae15d8d6c420a94baa0185c24518ca15415693c6a98dd325b51e86cfb9571510d50eb549ce2e8d0ba8baa7df0c1014eb5d25a4f0deeb24c67733c65e00528496229f73b6c6a412f1e62cfafcb08fc9d273eb400da3ba6b08cbeef6f6861b65d7e8cc48222cb218f3a9;
    5'b11110 : xpb = 1024'h5594cefa1fb8bf92599b214a4c81c7d8e81aee1465c3067e85e74d4c32a51b30b0a7ab34a48ad46d96891b14097b4b9e6e4ac5004a87d7595eefbd2f76e41e5effb64ab55800c890d7fba88c0fd52ebda4dca1e8165eaa6bc6532c30f52c9fb568e5c3e1c115966d70562b07a134ba3334f616b28597050752a5e3612b6db3ab;
    5'b11111 : xpb = 1024'hbdfc05d4cbe157bf38cdd670c3cda4560cf16c42ec8e34ef5f5c3d444a0eab75fc99424304b9399d67e6f7e85237187be0eba473dfa9dddaf2a3090bf3b311544c4b65e9feca5c48a5260393485970415f2e5cfda38beb4ed32a19b46464d84a4d08b12f2615a66f56c486b87fe6b9a7af536deefc83225d903a495a4c273ad;
    endcase
end

endmodule

module xpb_5_955
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'he9d422a168158799cd8201fb2e18f32274f542ea2fa1164b54c84fbb38ceb8f2f034341d01fa21d4e1c3471e13a6e0c8cb54e15835655a59cacb48980a7cfbb47e9d5ba8694c23caca23365d103afc68b1fa34647ebace69e1c9a1a8a94d86c9134aaa059af51d2724f53358fb842053215f9540bb3db346343ef448ae06301;
    5'b00010 : xpb = 1024'h1d3a84542d02b0f339b0403f65c31e644e9ea85d45f422c96a9909f76719d71e5e068683a03f443a9c3868e3c274dc19196a9c2b06acab4b39596913014f9f768fd3ab750d298479594466cba2075f8d163f468c8fd759cd3c3934351529b0d922695540b35ea3a4e49ea66b1f70840a642bf2a81767b668c687de8915c0c602;
    5'b00011 : xpb = 1024'h2bd7c67e4384096cd688605f18a4ad9675edfc8be8ee342e1fe58ef31aa6c2ad8d09c9c5705ee657ea549d55a3af4a25a61fea408a0300f0d6061d9c81f76f31d7bd812f93be46b605e69a31730b0f53a15ee9d2d7c306b3da55ce4f9fbe8945b39dffe10d0df57756edf9a0af28c60f9641ebfc231b919d29cbcdcda0a12903;
    5'b00100 : xpb = 1024'h3a7508a85a0561e67360807ecb863cc89d3d50ba8be84592d53213eece33ae3cbc0d0d07407e88753870d1c784e9b83232d538560d59569672b2d226029f3eed1fa756ea1a5308f2b288cd97440ebf1a2c7e8d191faeb39a7872686a2a5361b244d2aa8166bd4749c93d4cd63ee10814c857e5502ecf6cd18d0fbd122b818c04;
    5'b00101 : xpb = 1024'h49124ad27086ba601038a09e7e67cbfac48ca4e92ee256f78a7e98ea81c099cbeb105049109e2a92868d06396624263ebf8a866b90afac3c0f5f86af83470ea867912ca4a0e7cb2f5f2b00fd15126ee0b79e305f679a6081168f0284b4e83a1ed6075521c06c991c3b8ca00bce994a19fa6ddea43a834805f053ac56b661ef05;
    5'b00110 : xpb = 1024'h57af8cfc870812d9ad10c0be31495b2cebdbf917d1dc685c3fcb1de6354d855b1a13938ae0bdccafd4a93aab475e944b4c3fd481140601e1ac0c3b3903eede63af7b025f277c8d6c0bcd3462e6161ea742bdd3a5af860d67b4ab9c9f3f7d128b673bffc21a1beaeeaddbf3415e518c1f2c83d7f84637233a53979b9b41425206;
    5'b00111 : xpb = 1024'h664ccf269d896b5349e8e0dde42aea5f132b4d4674d679c0f517a2e1e8da70ea4916d6ccb0dd6ecd22c56f1d28990257d8f52296975c578748b8efc28496ae1ef764d819ae114fa8b86f67c8b719ce6dcddd76ebf771ba4e52c836b9ca11eaf7f870aa6273cb3cc1202b4676ee09ce245e99d14c51eafe6eb6db8adfcc22b507;
    5'b01000 : xpb = 1024'h74ea1150b40ac3cce6c100fd970c79913a7aa17517d08b25aa6427dd9c675c79781a1a0e80fd10ea70e1a38f09d3706465aa70ac1ab2ad2ce565a44c053e7dda3f4eadd434a611e565119b2e881d7e3458fd1a323f5d6734f0e4d0d454a6c36489a55502cd7a8e93927a99ac7dc2102990afcaa05d9ed9a31a1f7a2457031808;
    5'b01001 : xpb = 1024'h8387537aca8c1c468399211d49ee08c361c9f5a3baca9c8a5fb0acd94ff44808a71d5d50511cb307befdd800eb0dde70f25fbec19e0902d2821258d585e64d958738838ebb3ad42211b3ce9459212dfae41cbd788749141b8f016aeedf3b9bd11ad9ffa32729e06604c9ece20d7a522ec2c5c3f46952b4d77d636968e1e37b09;
    5'b01010 : xpb = 1024'h922495a4e10d74c02071413cfccf97f5891949d25dc4adef14fd31d503813397d620a092213c55250d1a0c72cc484c7d7f150cd7215f58781ebf0d5f068e1d50cf22594941cf965ebe5601fa2a24ddc16f3c60becf34c1022d1e050969d0743dac0eaa4380d93238771940179d329433f4dbbd487506900be0a758ad6cc3de0a;
    5'b01011 : xpb = 1024'ha0c1d7cef78ecd39bd49615cafb12727b0689e0100bebf53ca49b6d0b70e1f270523e3d3f15bf7425b3640e4ad82ba8a0bca5aeca4b5ae1dbb6bc1e88735ed0c170c2f03c864589b6af8355ffb288d87fa5c040517206de8cb3a9f23f4654caa3d4354e3da88840ae968934d2cead63926f1b69c80ba6b4043eb47f1f7a4410b;
    5'b01100 : xpb = 1024'haf5f19f90e1025b35a21817c6292b659d7b7f22fa3b8d0b87f963bcc6a9b0ab634272715c17b995fa95275568ebd2896987fa902280c03c35818767207ddbcc75ef604be4ef91ad8179a68c5cc2c3d4e857ba74b5f0c1acf6957393e7efa2516ce77ff843437d5dd5bb7e682bca3183e5907aff08c6e4674a72f37368284a40c;
    5'b01101 : xpb = 1024'hd4f16cd62a349642bf429c50519fe3a8d91432d713b41a5b70607726b25493d5fe1ecdec774bcee58106a818c9985d8c11acf3188af891d4425eb9d4db317d13290a5ca25fcdfcfb1a29989045428e41c9650f91a719aa551e7415e4f645af130a517fadd1e2f22474752d9548b341a3c43ca6247d6c478c403ab768482a0a2;
    5'b01110 : xpb = 1024'h1bec58f77924a1ddc8cc49e4b7fb8d6cb4e0975c1435530a6c528c6e1eb234cc8ee5302097945f0ba62c9ef36dd3f3e54dd01d470c05dec2e0d2a026ce5ae78c7a7a7b84ac91a20c5e44cceed557d8aaa7b5f43f625d478bf003db78d9f9335dc1d9c29b36cd80f4b996a60ee443761f6e59c3b6538a9fad27479abb0f6303a3;
    5'b01111 : xpb = 1024'h2a899b218fa5fa5765a46a046add1c9edc2feb8ab72f646f219f1169d23f205bbde8736267b40128f448d3654f0e61f1da856b5c8f5c34687d7f54b04f02b747c264513f332664490ae70054a65b887132d59785aa48f4728e207593648e0bca530e6d3b907cd2c72be5f94473fbb824a06fbd0a5f3e7ae18a8b89ff9a4366a4;
    5'b10000 : xpb = 1024'h3926dd4ba62752d1027c8a241dbeabd1037f3fb95a2975d3d6eb966585cc0beaecebb6a437d3a346426507d73048cffe673ab97212b28a0e1a2c0939cfaa87030a4e26f9b9bb2685b78933ba775f3837bdf53acbf234a1592c3d0fadef22e436e44317dbea2c24999e354c7a03b3fa29d285b65e6af25615edcf79442523c9a5;
    5'b10001 : xpb = 1024'h47c41f75bca8ab4a9f54aa43d0a03b032ace93e7fd2387388c381b613958f77a1beef9e607f3456390813c4911833e0af3f007879608dfb3b6d8bdc3505256be5237fcb4404fe8c2642b67204862e7fe4914de123a204e3fca59a9c879b7bca37577c27c43db766c10849faf936c3c2f049bafb276a6314a51136888b0042ca6;
    5'b10010 : xpb = 1024'h5661619fd32a03c43c2cca638381ca35521de816a01d989d4184a05cece5e3094af23d27d812e780de9d70baf2bdac1780a5559d195f35595385724cd0fa26799a21d26ec6e4aaff10cd9a86196697c4d4348158820bfb26687643e3044c951006ac6d1c9d8ac83e82d3f2e523247e3436b1a906825a0c7eb45757cd3ae48fa7;
    5'b10011 : xpb = 1024'h64fea3c9e9ab5c3dd904ea8336635967796d3c454317aa01f6d12558a072ce9879f58069a832899e2cb9a52cd3f81a240d5aa3b29cb58afef03226d651a1f634e20ba8294d796d3bbd6fcdebea6a478b5f54249ec9f7a80d0692ddfd8ee16d7c97e117bcf73a1a10f523461ab2dcc03968c7a25a8e0de7b3179b4711c5c4f2a8;
    5'b10100 : xpb = 1024'h739be5f4002cb4b775dd0aa2e944e899a0bc9073e611bb66ac1daa5453ffba27a8f8c3ab78522bbb7ad5d99eb53288309a0ff1c8200be0a48cdedb5fd249c5f029f57de3d40e2f786a120151bb6df751ea73c7e511e354f3a4af7818197645e92915c25d50e96be3677299504295023e9add9bae99c1c2e77adf365650a555a9;
    5'b10101 : xpb = 1024'h8239281e16ae0d3112b52ac29c2677cbc80be4a2890bcccb616a2f50078ca5b6d7fc06ed4871cdd8c8f20e10966cf63d26c53fdda362364a298b8fe952f195ab71df539e5aa2f1b516b434b78c71a71875936b2b59cf01da42cc1232a40b1e55ba4a6cfdaa98bdb5d9c1ec85d24d4443ccf39502a5759e1bde23259adb85b8aa;
    5'b10110 : xpb = 1024'h90d66a482d2f65aaaf8d4ae24f0806fdef5b38d12c05de3016b6b44bbb19914606ff4a2f18916ff6170e428277a76449b37a8df326b88befc6384472d3996566b9c92958e137b3f1c356681d5d7556df00b30e71a1baaec0e0e8ac4d2e9ff6c24b7f179e04480f884c113fbb62058648ff098e56b1297950416714df66661bab;
    5'b10111 : xpb = 1024'h9f73ac7243b0be244c656b0201e9963016aa8cffceffef94cc0339476ea67cd536028d70e8b11213652a76f458e1d256402fdc08aa0ee19562e4f8fc5441352201b2ff1367cc762e6ff89b832e7906a58bd2b1b7e9a65ba77f054667b934cf2edcb3c23e5df7615abe6092f0f1bdc84e311f87aabcdd5484a4ab0423f1467eac;
    5'b11000 : xpb = 1024'hae10ee9c5a32169de93d8b21b4cb25623df9e12e71fa00f9814fbe43223368646505d0b2b8d0b430b346ab663a1c4062cce52a1e2d65373aff91ad85d4e904dd499cd4cdee61386b1c9acee8ff7cb66c16f254fe3192088e1d21e08243c9a79b6de86cdeb7a6b32d30afe62681760a53633580fec8912fb907eef3687c26e1ad;
    5'b11001 : xpb = 1024'hc00eb70aec53a4ebb10336a57526d42f3d3322c3f7c71e6b8bf89e922bda6eb90c0967bbec9d7bf6204a09137f89da4f580504d8e08bc94eb9f22b11abe5fe71d3775d9c564fd62b6a2ffac37a4a201ae0cfeabecf7886405b1e8a21433dd75d0158555608d0c721c3f527d195e262f46719b7083f9adbd24c367a87e24de43;
    5'b11010 : xpb = 1024'h1a9e2d9ac54692c857e8538a0a33fc751b22865ae276834b6e0c0ee4d64a927abfc3d9bd8ee979dcb020d50319330bb182359e63115f123a884bd73a9b662fa265214b944bf9bf9f6345331208a851c8392ca1f234e3354aa3ce82bc9ec8b5e2614a2ff5ba3c5e448e8ea5b2a9166834788794c48fad88f1880756ed09054144;
    5'b11011 : xpb = 1024'h293b6fc4dbc7eb41f4c073a9bd158ba74271da89857094b0235893e089d77e09eec71cff5f091bf9fe3d0974fa6d79be0eeaec7894b567e024f88bc41c0dff5dad0b214ed28e81dc0fe76677d9ac018ec44c45387ccee23141eb1cd7295d8e4ef27eda9613ebb01700ddf8e838ceaa39aa9d8e189b616425eb4b463193e5a445;
    5'b11100 : xpb = 1024'h37d8b1eef24943bb919893c96ff71ad969c12eb8286aa614d8a518dc3d6469991dca60412f28be174c593de6dba7e7ca9ba03a8e180bbd85c1a5404d9cb5cf18f4f4f70959234418bc8999ddaaafb1554f6be87ec4ba8f17e007b6f1b3f266bb83b385366d9b01e9732d4c1dc886ec3edcb3876ca7153f5a4e8f35761ec60746;
    5'b11101 : xpb = 1024'h4675f41908ca9c352e70b3e922d8aa0b911082e6cb64b7798df19dd7f0f155284ccda382ff4860349a757258bce255d7285588a39b62132b5e51f4d71d5d9ed43cdeccc3dfb80655692bcd437bb3611bda8b8bc50ca63bfe7e24510c3e873f2814e82fd6c74a53bbe57c9f53583f2e440ec980c0b2c91a8eb1d324baa9a66a47;
    5'b11110 : xpb = 1024'h551336431f4bf4aecb48d408d5ba393db85fd7156e5ec8de433e22d3a47e40b77bd0e6c4cf680251e891a6ca9e1cc3e3b50ad6b91eb868d0fafea9609e056e8f84c8a27e664cc89215ce00a94cb710e265ab2f0b5491e8e51c40eb26c91c1794a61cda7720f9a58e57cbf288e7f7704940df7a14be7cf5c3151713ff3486cd48;
    5'b11111 : xpb = 1024'h63b0786d35cd4d286820f428889bc86fdfaf2b441158da42f88aa7cf580b2c46aad42a069f87a46f36addb3c7f5731f041c024cea20ebe7697ab5dea1ead3e4accb27838ece18acec270340f1dbac0a8f0cad2519c7d95cbba5d854153b0f001375185177aa8f760ca1b45be77afb24e72f57368ca30d0f7785b0343bf673049;
    endcase
end

endmodule

module xpb_5_390
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h22e55ec576d8e4dfa8bf75928d4acbc0dc9c04b28a76a9c0ed9860f3367292eb847c7bfc43fbeb38f6f8d6c5ed657f35840e24edd5a8e86006c5a2628c38a88f1454607833170bb41d41345baad1c06a4da0f9ccfd82c56a437b854d270b6d3c8a62c508c9652476308562d58e29b9b02c2dd8a0674f7fb4a952fb24820c349d;
    5'b00010 : xpb = 1024'h45cabd8aedb1c9bf517eeb251a959781b938096514ed5381db30c1e66ce525d708f8f7f887f7d671edf1ad8bdacafe6b081c49dbab51d0c00d8b44c51871511e28a8c0f0662e17683a8268b755a380d49b41f399fb058ad486f70a9a4e16da7914c58a1192ca48ec610ac5ab1c537360585bb140ce9eff6952a5f6490418693a;
    5'b00011 : xpb = 1024'h68b01c50648aae9efa3e60b7a7e0634295d40e179f63fd42c8c922d9a357b8c28d7573f4cbf3c1aae4ea8451c8307da08c2a6ec980fab9201450e727a4a9f9ad3cfd21689945231c57c39d130075413ee8e2ed66f888503eca728fe7752247b59f284f1a5c2f6d6291902880aa7d2d10848989e135ee7f1dfbf8f16d86249dd7;
    5'b00100 : xpb = 1024'h8b957b15db63937ea2fdd64a352b2f03727012ca29daa703b66183ccd9ca4bae11f1eff10feface3dbe35b17b595fcd6103893b756a3a1801b16898a30e2a23c515181e0cc5c2ed07504d16eab4701a93683e733f60b15a90dee15349c2db4f2298b1423259491d8c2158b5638a6e6c0b0b762819d3dfed2a54bec920830d274;
    5'b00101 : xpb = 1024'hae7ad9db523c785e4bbd4bdcc275fac44f0c177cb45150c4a3f9e4c0103cde99966e6bed53eb981cd2dc31dda2fb7c0b9446b8a52c4c89e021dc2becbd1b4acb65a5e258ff733a84924605ca5618c2138424e100f38ddb1351699a81c339222eb3edd92beef9b64ef29aee2bc6d0a070dce53b22048d7e874e9ee7b68a3d0711;
    5'b00110 : xpb = 1024'h20b2f34b07272875297749983f667f33ba3218fe69505a0e13b58c5d93acc47d17a26a70cdc104c72a76c95cad02ea76b43ab5acdf42a1f478028ef10e817ea905ab0e2282f948f39ced3783680ebe4cddc0e135648a736cdf588dd43019ecd90f490c0b0795e2379c606a225d2a33f7ba3934e01b91a10bb18267d68366d543;
    5'b00111 : xpb = 1024'h439852107e000d54d236bf2accb14af496ce1db0f3c703cf014ded50ca1f57689c1ee66d11bcf000216fa0229a6869ac3848da9ab4eb8a547ec831539aba273819ff6e9ab61054a7ba2e6bdf12e07eb72b61db02620d38d722d4132157255a1599abd113d0fb06adcce5ccf7eb53eda7e6670d8082e120c05ad562fb057309e0;
    5'b01000 : xpb = 1024'h667db0d5f4d8f2347af634bd59fc16b5736a22637e3dad8feee64e440091ea54209b626955b8db39186876e887cde8e1bc56ff888a9472b4858dd3b626f2cfc72e53cf12e927605bd76fa03abdb23f217902d4cf5f8ffe41664f986e7e30c752240e961c9a602b23fd6b2fcd797da7581294e620ea30a07504285e1f877f3e7d;
    5'b01001 : xpb = 1024'h89630f9b6bb1d71423b5aa4fe746e2765006271608b45750dc7eaf3737047d3fa517de6599b4c6720f614dae7533681740652476603d5b148c537618b32b785642a82f8b1c3e6c0ff4b0d4966883ff8bc6a3ce9c5d12c3aba9cb1dbba53c348eae715b2563c54f9a2df092a307a761083ec2bec151802029ad7b5944098b731a;
    5'b01010 : xpb = 1024'hac486e60e28abbf3cc751fe27491ae372ca22bc8932b0111ca17102a6d77102b29945a61ddb0b1ab065a24746298e74cc473496435e643749319187b3f6420e556fc90034f5577c411f208f21355bff61444c8695a958915ed46a308cc47a1cb38d4202e2d2a74105e75f57895d11ab86af09761b8cf9fde56ce54688b97a7b7;
    5'b01011 : xpb = 1024'h1e8087d097756c0aaa2f1d9df18232a697c82d4a482a0a5b39d2b7c7f0e6f60eaac858e557861e555df4bbf36ca055b7e467466be8dc5b88e93f7b7f90ca54c2f701bbccd2db86331c993aab254bbc2f6de0c89dcb92216f7b35965b39286c75942f530d45c69ff9083b716f2c2aae3f4844911fcfd3c262b9b1d48884c175e9;
    5'b01100 : xpb = 1024'h4165e6960e4e50ea52ee93307eccfe67746431fcd2a0b41c276b18bb275988fa2f44d4e19b82098e54ed92b95a05d4ed68756b59be8543e8f0051de21d02fd520b561c4505f291e739da6f06d01d7c99bb81c26ac914e6d9beb11ba86033d9b21e9218160f2bc46f38c0d444ba5467ef747269c0372342176304cfad06cdaa86;
    5'b01101 : xpb = 1024'h644b455b852735c9fbae08c30c17ca28510036af5d175ddd150379ae5dcc1be5b3c150dddf7df4c74be6697f476b5422ec839047942e2c48f6cac044a93ba5e11faa7cbd39099d9b571ba3627aef3d040922bc37c697ac44022ca0f5873f46eea8f4dd1ed890e8e56946371a487e219fa0a042609e72c1cc0c57cad188d9df23;
    5'b01110 : xpb = 1024'h8730a420fc001aa9a46d7e55996295e92d9c3b61e78e079e029bdaa1943eaed1383dccda2379e00042df404534d0d3587091b53569d714a8fd9062a735744e7033fedd356c20a94f745cd7be25c0fd6e56c3b604c41a71ae45a82642ae4ab42b3357a227a1f60d5b99cb99efd6a7db4fccce1b0105c24180b5aac5f60ae613c0;
    5'b01111 : xpb = 1024'haa1602e672d8ff894d2cf3e826ad61aa0a3840147204b15ef0343b94cab141bcbcba48d66775cb3939d8170b2236528df49fda233f7ffd0904560509c1acf6ff48533dad9f37b503919e0c19d092bdd8a464afd1c19d37188923ab8fd5562167bdba67306b5b31d1ca50fcc564d194fff8fbf3a16d11c1355efdc11a8cf2485d;
    5'b10000 : xpb = 1024'h1c4e1c5627c3afa02ae6f1a3a39de619755e41962703baa85fefe3324e2127a03dee4759e14b37e39172ae8a2c3dc0f91493d72af276151d5a7c680e13132adce858697722bdc3729c453dd2e288ba11fe00b0063299cf7217129ee24236ec1219159a0f83f75dba741678bbfb2b2886d64fed5f8415e3b9c1e1413a861c168f;
    5'b10001 : xpb = 1024'h3f337b1b9e9c947fd3a6673630e8b1da51fa4648b17a64694d8844258493ba8bc26ac3562547231c886b855019a3402e98a1fc18c81efd7d61420a709f4bd36bfcacc9ef55d4cf26b986722e8d5a7a7c4ba1a9d3301c94dc5a8e242f6942594ea3785f184d5c8230a49bdb918954e237027dc5ffeb65636e6b343c5f08284b2c;
    5'b10010 : xpb = 1024'h6218d9e11575795f7c65dcc8be337d9b2e964afb3bf10e2a3b20a518bb064d7746e73f5269430e557f645c160708bf641cb021069dc7e5dd6807acd32b847bfb11012a6788ebdadad6c7a68a382c3ae69942a3a02d9f5a469e09a97c904dc68b2ddb242116c1a6a6d5213e67177e9be72eab9ea052b4e323148737838a347fc9;
    5'b10011 : xpb = 1024'h84fe38a68c4e5e3f2525525b4b7e495c0b324fadc667b7eb28b9060bf178e062cb63bb4ead3ef98e765d32dbf46e3e99a0be45f47370ce3d6ecd4f35b7bd248a25558adfbc02e68ef408dae5e2fdfb50e6e39d6d2b221fb0e1852ec9b75933c7b83de929e026cb1d05a6a13ca5a855975ad97740ba0462d7bdda32a80c40b466;
    5'b10100 : xpb = 1024'ha7e3976c0327431ecde4c7edd8c9151ce7ce546050de61ac165166ff27eb734e4fe0374af13ae4c76d5609a1e1d3bdcf24cc6ae24919b69d7592f19843f5cd1939a9eb57ef19f243114a0f418dcfbbbb3484973a28a4e51b2500b416de64a10442a0ae32a98bef93362c041233d20f4787074fe12153e28c672d2dcc8e4ce903;
    5'b10101 : xpb = 1024'h1a1bb0dbb811f335ab9ec5a955b9998c52f455e205dd6af5860d0e9cab5b5931d11435ce6b105171c4f0a120ebdb2c3a44c067e9fc0fceb1cbb9549c955c00f6d9af172172a000b21bf140fa9fc5b7f48e20976e99a17d74b2efa7694b456bae9dfbe111c2281b7bdff18008ca2ba2ce645b499f38580510ca10adec8776b735;
    5'b10110 : xpb = 1024'h3d010fa12eead815545e3b3be304654d2f905a94905414b673a56f8fe1cdec1d5590b1caaf0c3caabbe977e6d940ab6fc8ce8cd7d1b8b711d27ef6ff2194a985ee037799a5b70c66393275564a97785edbc1913b972442def66b2cb67250d8eb285ea61a8b8d3ff21076e2de58555c7e9089223f9fa784c57363a9110982ebd2;
    5'b10111 : xpb = 1024'h5fe66e66a5c3bcf4fd1db0ce704f310e0c2c5f471acabe77613dd08318407f08da0d2dc6f30827e3b2e24eacc6a62aa54cdcb1c5a7619f71d9449961adcd52150257d811d8ce181a5673a9b1f56938c929628b0894a7084939e6b203995c4627b2c16b2354f2646840fc45b3e67f162ebcb6fae006f7047a1cb6a4358b8f206f;
    5'b11000 : xpb = 1024'h82cbcd2c1c9ca1d4a5dd2660fd99fccee8c863f9a54168384ed631764eb311f45e89a9c33704131ca9db2572b40ba9dad0ead6b37d0a87d1e00a3bc43a05faa416ac388a0be523ce73b4de0da03af933770384d59229cdb37d623750c067b3643d24302c1e5788de7181a88974a8cfdee8e4d3806e46842ec6099f5a0d9b550c;
    5'b11001 : xpb = 1024'ha5b12bf1937586b44e9c9bf38ae4c88fc56468ac2fb811f93c6e92698525a4dfe30625bf7afffe55a0d3fc38a171291054f8fba152b37031e6cfde26c63ea3332b0099023efc2f8290f612694b0cb99dc4a47ea28fac931dc0ddbc9de77320a0c786f534e7bcad54a2070b5f02d2898f1512ac20d59603e36f5c9a7e8fa789a9;
    5'b11010 : xpb = 1024'h17e94561486036cb2c5699af07d54cff308a6a2de4b71b42ac2a3a0708958ac3643a2442f4d56afff86e93b7ab78977b74ecf8a905a988463cf6412b17a4d710cb05c4cbc2823df19b9d44225d02b5d71e407ed700a92b774eccaff05453eb4b22e228140058d93d4bcc8755992c1d15f266a5deec9a2667d2401a9e88d157db;
    5'b11011 : xpb = 1024'h3acea426bf391baad5160f41952018c00d266ee06f2dc50399c29afa3f081daee8b6a03f38d15638ef676a7d98de16b0f8fb1d96db5270a643bbe38da3dd7f9fdf5a2543f59949a5b8de787e07d476416be178a3fe2bf0e19248353d7b5f5887ad44ed1cc9bdfdb37c51ea2b2755d6c61e947e7f53e9a61c7b9315c30add8c78;
    5'b11100 : xpb = 1024'h5db402ec3612008a7dd584d4226ae480e9c27392f9a46ec4875afbed757ab09a6d331c3b7ccd4171e6604143864395e67d094284b0fb59064a8185f03016282ef3ae85bc28b05559d61facd9b2a636abb9827270fbaeb64bd5c3ba8aa26ac5c437a7b22593232229acd74d00b57f90764ac2571fbb3925d124e610e78ce9c115;
    5'b11101 : xpb = 1024'h809961b1aceae56a2694fa66afb5b041c65e7845841b188574f35ce0abed4385f1af9837c0c92caadd59180973a9151c0117677286a4416651472852bc4ed0be0802e6345bc7610df360e1355d77f71607236c3df9317bb6193f3fd7c9763300c20a772e5c88469fdd5cafd643a94a2676f02fc02288a585ce390c0c0ef5f5b2;
    5'b11110 : xpb = 1024'ha37ec07723c3ca49cf546ff93d007c02a2fa7cf80e91c246628bbdd3e25fd671762c143404c517e3d451eecf610e945185258c605c4d29c6580ccab54887794d1c5746ac8ede6cc210a215910849b78054c4660af6b441205cbac524f081a03d4c6d3c3725ed6b160de212abd1d303d6a31e086089d8253a778c073091022a4f;
    5'b11111 : xpb = 1024'h15b6d9e6d8ae7a60ad0e6db4b9f100720e207e79c390cb8fd247657165cfbc54f76012b77e9a848e2bec864e6b1602bca51989680f4341daae332db999edad2abc5c727612647b311b49474a1a3fb3b9ae60663f67b0d979eaa9b8775d626ae7a7c86f163e8996feb7a78ea2682c975d8072021ea0dc47beda6f87508a2bf881;
    endcase
end

endmodule

module xpb_5_175
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h9f3da7e808fb60854d2b6648b6eae4e794ea52fabbce67585b59442e28ca912b2387b7b74ed52ac3a322f9d01d0f3030c5b6665011a46a91a5eb49f81a11691d7ce92d2a2e82995f6bcc2c49f298a4c3c2014e6b492f8018706fcb2acf44bc1ee57dafd47c02f6931d144196cbf1491d3ab4149e44f9d7f0a7a767a198da2d5;
    5'b00010 : xpb = 1024'h13e7b4fd011f6c10a9a56cc916dd5c9cf29d4a5f5779cceb0b6b2885c51952256470f6f6e9daa55874645f3a03a1e60618b6ccca02348d5234bd693f03422d23af9d25a545d0532bed7985893e531498784029cd6925f0030e0df96559e89783dcafb5fa8f805ed263a28832d97e2923a7568293c89f3afe14f4ecf4331b45aa;
    5'b00011 : xpb = 1024'h1ddb8f7b81af2218fe78232da24c0aeb6bebef8f0336b3609120bcc8a7a5fb3816a972725ec7f804ae968ed70572d9092512332f034ed3fb4f1c1dde84e343b5876bb877e8b87cc1e436484ddd7c9ee4b4603eb41db8e8049514f61806dce345cb0790f7d7408e3b9573cc4c463d3db57b01c3ddaceed87d1f6f636e4ca8e87f;
    5'b00100 : xpb = 1024'h27cf69fa023ed821534ad9922dbab939e53a94beaef399d616d6510b8a32a44ac8e1ededd3b54ab0e8c8be740743cc0c316d999404691aa4697ad27e06845a475f3a4b4a8ba0a657daf30b127ca62930f080539ad24be0061c1bf2cab3d12f07b95f6bf51f00bda4c7451065b2fc52474ead0527913e75fc29e9d9e866368b54;
    5'b00101 : xpb = 1024'h31c3447882ce8e29a81d8ff6b92967885e8939ee5ab0804b9c8be54e6cbf4d5d7b1a696948a29d5d22faee110914bf0f3dc8fff90583614d83d9871d882570d93708de1d2e88cfedd1afcdd71bcfb37d2ca0688186ded807a322ef7d60c57ac9a7b746f266c0ed0df916547f1fbb66d922584671758e137b346450627fc42e29;
    5'b00110 : xpb = 1024'h3bb71ef7035e4431fcf0465b449815d6d7d7df1e066d66c1224179914f4bf6702d52e4e4bd8ff0095d2d1dae0ae5b2124a24665e069da7f69e383bbd09c6876b0ed770efd170f983c86c909bbaf93dc968c07d683b71d0092a29ec300db9c68b960f21efae811c772ae798988c7a7b6af60387bb59ddb0fa3edec6dc9951d0fe;
    5'b00111 : xpb = 1024'h45aaf97583edfa3a51c2fcbfd006c4255126844db22a4d36a7f70dd431d89f82df8b6060327d42b5975f4d4b0cb6a515567fccc307b7ee9fb896f05c8b679dfce6a603c274592319bf2953605a22c815a4e0924ef004c80ab130e8e2baae124d8466fcecf6414be05cb8dcb1f9398ffcc9aec9053e2d4e7949593d56b2df73d3;
    5'b01000 : xpb = 1024'h4f9ed3f4047db042a695b3245b757273ca75297d5de733ac2daca2171465489591c3dbdba76a9561d1917ce80e87981862db332808d23548d2f5a4fc0d08b48ebe74969517414cafb5e61624f94c5261e100a735a497c00c3837e59567a25e0f72bed7ea3e017b498e8a20cb65f8a48e9d5a0a4f227cebf853d3b3d0cc6d16a8;
    5'b01001 : xpb = 1024'h5992ae72850d664afb686988e6e420c243c3cead09a41a21b3623659f6f1f1a843fc57571c57e80e0bc3ac8510588b1b6f36998d09ec7bf1ed54599b8ea9cb2096432967ba297645aca2d8e99875dcae1d20bc1c592ab80dbf3ee2481496a9d16116b2e785c1aab2c05b64e4d2b7b92071054b9906cc89775e4e2a4ae5fab97d;
    5'b01010 : xpb = 1024'h638688f1059d1c53503b1fed7252cf10bd1273dcb56100973917ca9cd97e9abaf634d2d291453aba45f5dc2212297e1e7b91fff20b06c29b07b30e3b104ae1b26e11bc3a5d119fdba35f9bae379f66fa5940d1030dbdb00f4645defac18af5934f6e8de4cd81da1bf22ca8fe3f76cdb244b08ce2eb1c26f668c8a0c4ff885c52;
    5'b01011 : xpb = 1024'h6d7a636f862cd25ba50dd651fdc17d5f3661190c611de70cbecd5edfbc0b43cda86d4e4e06328d6680280bbf13fa712187ed66570c2109442211c2da91ebf84445e04f0cfff9c9719a1c5e72d6c8f1469560e5e9c250a810cd4cdbad6e7f41553dc668e21542098523fded17ac35e244185bce2ccf6bc4757343173f1915ff27;
    5'b01100 : xpb = 1024'h776e3dee06bc8863f9e08cb689302badafafbe3c0cdacd824482f3229e97ece05aa5c9c97b1fe012ba5a3b5c15cb64249448ccbc0d3b4fed3c70777a138d0ed61daee1dfa2e1f30790d9213775f27b92d180fad076e3a0125453d8601b738d172c1e43df5d0238ee55cf313118f4f6d5ec070f76b3bb61f47dbd8db932a3a1fc;
    5'b01101 : xpb = 1024'h8162186c874c3e6c4eb3431b149ed9fc28fe636bb897b3f7ca388765812495f30cde4544f00d32bef48c6af9179c5727a0a433210e55969656cf2c19952e2567f57d74b245ca1c9d8795e3fc151c05df0da10fb72b769813db5ad512c867d8d91a761edca4c2685787a0754a85b40b67bfb250c0980aff73883804334c3144d1;
    5'b01110 : xpb = 1024'h8b55f2eb07dbf474a385f97fa00d884aa24d089b64549a6d4fee1ba863b13f05bf16c0c064fa856b2ebe9a96196d4a2aacff99860f6fdd3f712de0b916cf3bf9cd4c0784e8b246337e52a6c0b445902b49c1249de00990156261d1c5755c249b08cdf9d9ec8297c0b971b963f2731ff9935d920a7c5a9cf292b27aad65bee7a6;
    5'b01111 : xpb = 1024'h9549cd69886baa7cf858afe42b7c36991b9badcb101180e2d5a3afeb463de818714f3c3bd9e7d81768f0ca331b3e3d2db95affeb108a23e88b8c95589870528ba51a9a578b9a6fc9750f6985536f1a7785e13984949c8816e968ce782250705cf725d4d73442c729eb42fd7d5f32348b6708d35460aa3a719d2cf1277f4c8a7b;
    5'b10000 : xpb = 1024'h9f3da7e808fb60854d2b6648b6eae4e794ea52fabbce67585b59442e28ca912b2387b7b74ed52ac3a322f9d01d0f3030c5b6665011a46a91a5eb49f81a11691d7ce92d2a2e82995f6bcc2c49f298a4c3c2014e6b492f8018706fcb2acf44bc1ee57dafd47c02f6931d144196cbf1491d3ab4149e44f9d7f0a7a767a198da2d50;
    5'b10001 : xpb = 1024'ha9318266898b168da1fe1cad425993360e38f82a678b4dcde10ed8710b573a3dd5c03332c3c27d6fdd55296d1ee02333d211ccb512beb13ac049fe979bb27faf54b7bffcd16ac2f56288ef0e91c22f0ffe216351fdc27819f776c7dd7c3907e0d3d58ad1c3c325fc4ee585b038b05daf0e5f55e82949756fb221de1bb267d025;
    5'b10010 : xpb = 1024'h278178f482c97cd2bcb5b3abd6dfa3316119a293dd093cbe8e7b35e3ae1364884b031356e89518d782919c33d53056c7a530b33f12627982a0973d8e281218fb8371e20c4c1ef4646abaf30980ff52b463c7ea025cf430ac8f132956f02b1109325d3a55aba5cd7f9f6e2eaad9f4c179330b84fbd4db5be762cd99143130c8f;
    5'b10011 : xpb = 1024'hc6bf20dc8bc4dd5809e119f48dca8818f603f58e98d7a416e9d47a11d6ddf5b36e8acb0e376a439b25b49603f23f86f86ae7198f2406e4144682878642238219005b0f367aa18dc3d6871f537397f77825c9386da623b0c4ff82f481bf6fcd2817daea2a27a8c412bc827041a5e60a966dbf999a19d533d80a7500b5ca0af64;
    5'b10100 : xpb = 1024'h165fcc8c494c03ddd570c803d44b56d008aee488954a60b6f452dbe3fffa886de921282c5863f6e5ec8d78fd40f4eb729309d7fdf35ab4ea5ec6dd17e5c34eb367d443c60a924272342534b9d66309c3be7ca86d8ef5330dd6ff2bfac8eb48946fd5899fea3abbaa5d996b1d871d753b3a873ae385ecf0bc8b21c685762e5239;
    5'b10101 : xpb = 1024'h2053a70ac9dbb9e62a437e685fba051e81fd89b84107472c7a087026e28731809b59a3a7cd51499226bfa89a42c5de759f653e62f474fb93792591b7676465453fa2d698ad7a6c082ae1f77e758c940ffa9cbd5443882b0f5e0628ad75df94565e2d649d31faeb138f6aaf36f3dc89cd0e327c2d6a3c8e3b959c3cff8fbbf50e;
    5'b10110 : xpb = 1024'h2a4781894a6b6fee7f1634cceb28b36cfb4c2ee7ecc42da1ffbe0469c513da934d921f23423e9c3e60f1d8374496d178abc0a4c7f58f423c93844656e9057bd71771696b5062959e219eba4314b61e5c36bcd23af81b2310e50d256022d3e0184c853f9a79bb1a7cc13bf350609b9e5ee1ddbd774e8c2bbaa016b379a94997e3;
    5'b10111 : xpb = 1024'h343b5c07cafb25f6d3e8eb31769761bb749ad41798811417857398aca7a083a5ffca9a9eb72beeea9b2407d44667c47bb81c0b2cf6a988e5ade2faf66aa69268ef3ffc3df34abf34185b7d07b3dfa8a872dce721acae1b126c142212cfc82bda3add1a97c17b49e5f30d3769cd5ab2f0b588fec132dbc939aa9129f3c2d73ab8;
    5'b11000 : xpb = 1024'h3e2f36864b8adbff28bba19602061009ede97947443dfa8d0b292cef8a2d2cb8b203161a2c194196d55637714838b77ec4777191f7c3cf8ec841af95ec47a8fac70e8f109632e8ca0f183fcc530932f4aefcfc0861411313f31b1ec57cbc779c2934f595093b794f24de7b833a19c7828934400b172b66b8b50ba06ddc64dd8d;
    5'b11001 : xpb = 1024'h48231104cc1a92077d8e57fa8d74be5867381e76effae10290dec1326cb9d5cb643b9195a10694430f88670e4a09aa81d0d2d7f6f8de1637e2a064356de8bf8c9edd21e3391b126005d50290f232bd40eb1d10ef15d40b157a221b7829b0c35e178cd09250fba8b856afbf9ca6d8dc145cdf8154fb7b0437bf8616e7f5f28062;
    5'b11010 : xpb = 1024'h5216eb834caa480fd2610e5f18e36ca6e086c3a69bb7c778169455754f467ede16740d1115f3e6ef49ba96ab4bda9d84dd2e3e5bf9f85ce0fcff18d4ef89d61e76abb4b5dc033bf5fc91c555915c478d273d25d5ca6703170129182ad6a50f2005e4ab8f98bbd821888103b61397f0a6308ac29edfcaa1b6ca008d620f802337;
    5'b11011 : xpb = 1024'h5c0ac601cd39fe182733c4c3a4521af559d568d64774aded9c49e9b831d327f0c8ac888c8ae1399b83ecc6484dab9087e989a4c0fb12a38a175dcd74712aecb04e7a47887eeb658bf34e881a3085d1d9635d3abc7ef9fb18883014dd83995ae1f43c868ce07c078aba5247cf80570538043603e8c41a3f35d47b03dc290dc60c;
    5'b11100 : xpb = 1024'h65fea0804dc9b4207c067b282fc0c943d3240e05f331946321ff7dfb145fd1037ae50407ffce8c47be1ef5e54f7c838af5e50b25fc2cea3331bc8213f2cc03422648da5b21d38f21ea0b4adecfaf5c259f7d4fa3338cf31a0f371190308da6a3e294618a283c36f3ec238be8ed1619c9d7e14532a869dcb4def57a56429b68e1;
    5'b11101 : xpb = 1024'h6ff27afece596a28d0d9318cbb2f77924c72b3359eee7ad8a7b5123df6ec7a162d1d7f8374bbdef3f8512582514d768e0240718afd4730dc4c1b36b3746d19d3fe176d2dc4bbb8b7e0c80da36ed8e671db9d6489e81feb1b963e0e42dd81f265d0ec3c876ffc665d1df4d00259d52e5bab8c867c8cb97a33e96ff0d05c290bb6;
    5'b11110 : xpb = 1024'h79e6557d4ee9203125abe7f1469e25e0c5c158654aab614e2d6aa680d9792328df55fafee9a931a03283551f531e69910e9bd7effe6177856679eb52f60e3065d5e6000067a3e24dd784d0680e0270be17bd79709cb2e31d1d450af58a763e27bf441784b7bc95c64fc6141bc69442ed7f37c7c6710917b2f3ea674a75b6ae8b;
    5'b11111 : xpb = 1024'h83da2ffbcf78d6397a7e9e55d20cd42f3f0ffd94f66847c3b3203ac3bc05cc3b918e767a5e96844c6cb584bc54ef5c941af73e54ff7bbe2e80d89ff277af46f7adb492d30a8c0be3ce41932cad2bfb0a53dd8e575145db1ea44c07a8376a89e9ad9bf281ff7cc52f819758353353577f52e309105558b531fe64ddc48f445160;
    endcase
end

endmodule

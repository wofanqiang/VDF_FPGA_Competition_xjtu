module xpb_5_215
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h5a5aa6466bf4f17107cc73e286fba0d8106104b062ce38e4da557123322025d763f04bc53163974e95bd3e39da9b3f8ff974a7e93b1bd702686c7e026605d9c624dbd75748a747c557771a00fb3268c61bd6d02969548b81d9acaf70d912528fad41bf96b03cbd3c8c457ccb5146e219a56d80e70c6c01424424ce1480c6da28;
    5'b00010 : xpb = 1024'h408073715fbae1944936fedfd9cfa5eaf4c062ff024d15236ce28f0b13d9ea6c4981a1198a0b00e8c1c3d2cd1d86e558ecf27ec5384ddb92039bca691393edad56879ffe1bd92459c54315f5d890d5b43a8a6ba4622e9f2fdcccce6f7fa028d2b7bed03afb081eb91cb12b7aabd9e09fc0122ebc88ca55441da212478ab4de5;
    5'b00011 : xpb = 1024'h5e62ad7d81f09f8a4c5fe3d084989b36bfad0ae052f30a3711239a13e35dc47e288865d6ca04475d21d97b66ac73ade58843cfd58ea0b4bb88a63aa8f73f18a0fa4451572a64da0af3cb4b6058bb76215f7f76e3af777574d7797c57d10c551cd8bdac9a5fed3f281e108f82fc048023a16ea3d2d4f8a69685feef38f972280d;
    5'b00100 : xpb = 1024'h8100e6e2bf75c328926dfdbfb39f4bd5e980c5fe049a2a46d9c51e1627b3d4d893034233141601d18387a59a3b0dcab1d9e4fd8a709bb724073794d22727db5aad0f3ffc37b248b38a862bebb121ab687514d748c45d3e5fb9999cdeff4051a56f7da075f6103d72396256f557b3c13f80245d791194aa883b44248f1569bca;
    5'b00101 : xpb = 1024'h626ab4b497ec4da390f353be823595956ef911104317db8947f1c304949b6324ed207fe862a4f76badf5b8937e4c1c3b1712f7c1e2259274a8dff74f8878577bcfaccb570c226c50901f7cbfb644837ca3281d9df59a5f67d546493ec90657aa0439999e0f9dc113afdba23aa6c21e2d9d6fc6be9d854beac7d9105d721d75f2;
    5'b00110 : xpb = 1024'hc1815a541f30a4bcdba4fc9f8d6ef1c0de4128fd06e73f6a46a7ad213b8dbf44dc84e34c9e2102ba454b78675894b00ac6d77c4fa8e992b60ad35f3b3abbc9080396dffa538b6d0d4fc941e189b2811caf9f42ed268bdd8f96666b4e7ee07a78273c70b0f1185c2b56138270038da1df40368c359a5effcc58e636d6a01e9af;
    5'b00111 : xpb = 1024'h6672bbebade7fbbcd586c3ac7fd28ff41e451740333cacdb7ebfebf545d901cbb1b899f9fb45a77a3a11f5c050248a90a5e21fae35aa702dc919b3f619b19656a5154556eddffe962c73ae1f13cd90d7e6d0c4583bbd495ad3131625c1005a372fb586a1bf4e42ff41a6b4f2517fbc379970e9aa6611f13f09b33181eac8c3d7;
    5'b01000 : xpb = 1024'h10201cdc57eeb865124dbfb7f673e97abd3018bfc0934548db38a3c2c4f67a9b126068466282c03a3070f4b34761b9563b3c9fb14e1376e480e6f29a44e4fb6b55a1e7ff86f649167150c57d7624356d0ea29ae9188ba7cbf733339bdfe80a34adefb40ebec207ae472c4adeaaf67827f0048baf2232955107688491e2ad3794;
    5'b01001 : xpb = 1024'h6a7ac322c3e3a9d61a1a339a7d6f8a52cd911d7023617e2db58e14e5f716a0727650b40b93e65788c62e32ed21fcf8e634b1479a892f4de6e953709caaead5317a7dbf56cf9d90dbc8c7df7e71569e332a796b1281e0334dd0dfe30cb8fa5cc45b3173a56efec4ead371c7a9fc3d5a4195720c962e9e96934b8d52a6637411bc;
    5'b01010 : xpb = 1024'h142824136dea667e56e12fa5f410e3d96c7c1eefb0b8169b1206ccb376341941d6f88257fb237048bc8d31e0193a27abca0bc79da198549da120af40d61e3a462b0a61ff68b3db5c0da4f6dcd3ad42c8524b41a35eae91bef5000082d7e20cc1d96ba1126e728999d8f75d9655b41631ec05ae9aeabf3aa54942a5b65b588579;
    5'b01011 : xpb = 1024'h6e82ca59d9df57ef5eada3887b0c84b17cdd23a013864f7fec5c3dd6a8543f193ae8ce1d2c870797524a7019f3d5673bc3806f86dcb42ba0098d2d433c24140c4fe63956b15b2321651c10ddcedfab8e6e2211ccc8031d40ceacaff3b0f45f5186ad60a91eaf46d6653cda61a6faf84b91732f81f72b3be78d6773cadc1f5fa1;
    5'b01100 : xpb = 1024'h18302b4a83e614979b749f93f1adde381bc8251fa0dce7ed48d4f5a42771b7e89b909c6993c4205748a96f0ceb12960158daef89f51d3256c15a6be7675779210072dbff4a716da1a9f9283c3136502395f3e85da4d17bb1f2cccd69cfdc0f4f04e78e161e230b856ac2704e0071b43be806d186b34bdff98b1cc6dad403d35e;
    5'b01101 : xpb = 1024'h728ad190efdb0608a341137678a97f102c2929d003ab20d2232a66c75991ddbfff80e82ec527b7a5de66ad46c5add591524f97733039095929c6e9e9cd5d52e7254eb3569318b5670170423d2c68b8e9b1cab8870e260733cc797cdaa8ee61deb2294dacce5fc8c1f707ed1951b896558d74526dbfb7e13bcf4194ef54caad86;
    5'b01110 : xpb = 1024'h1c38328199e1c2b0e0080f81ef4ad896cb142b4f9101b93f7fa31e94d8af568f6028b67b2c64d065d4c5ac39bceb0456e7aa177648a2100fe194288df890b7fbd5db55ff2c2effe7464d599b8ebf5d7ed99c8f17eaf465a4f0999a50c7d611dc30637b19cdd38d70fc8d8305ab2f5245e407f4727bd8854dccf6e7ff4caf2143;
    5'b01111 : xpb = 1024'h7692d8c805d6b421e7d483647646796edb752ffff3cff22459f88fb80acf7c66c41902405dc867b46a82ea73978643e6e11ebf5f83bde7124a00a6905e9691c1fab72d5674d647ac9dc4739c89f1c644f5735f415448f126ca4649c1a0e8646bdda53ab07e104aad88d2ffd0fc76345f8975755988448690111bb613cd75fb6b;
    5'b10000 : xpb = 1024'h204039b8afdd70ca249b7f6fece7d2f57a60317f81268a91b671478589ecf53624c0d08cc505807460e1e9668ec372ac76793f629c26edc901cde53489c9f6d6ab43cfff0dec922ce2a18afaec486ada1d4535d231174f97ee666737bfd014695bdf681d7d840f5c8e5895bd55ecf04fe009175e44652aa20ed10923c55a6f28;
    5'b10001 : xpb = 1024'h7a9adfff1bd2623b2c67f35273e373cd8ac1362fe3f4c37690c6b8a8bc0d1b0d88b11c51f66917c2f69f27a0695eb23c6fede74bd742c4cb6a3a6336efcfd09cd01fa7565693d9f23a18a4fbe77ad3a0391c05fb9a6bdb19c81316a898e266f9092127b42dc0cc991a9e1288a733d2698576984550d12be452f5d73846214950;
    5'b10010 : xpb = 1024'h244840efc5d91ee3692eef5dea84cd5429ac37af714b5be3ed3f70763b2a93dce958ea9e5da63082ecfe2693609be1020548674eefabcb822207a1db1b0335b180ac49feefaa24727ef5bc5a49d1783560eddc8c773a398aec33341eb7ca16f6875b55212d3491482023a87500aa8e59dc0a3a4a0cf1cff650ab2a483e05bd0d;
    5'b10011 : xpb = 1024'h7ea2e73631ce105470fb634071806e2c3a0d3c5fd41994c8c794e1996d4ab9b44d4936638f09c7d182bb64cd3b372091febd0f382ac7a2848a741fdd81090f77a588215638516c37d66cd65b4503e0fb7cc4acb5e08ec50cc5dfe38f90dc6986349d14b7dd714e84ac69254051f170738177bb31195dd13894cff85cbecc9735;
    5'b10100 : xpb = 1024'h28504826dbd4ccfcadc25f4be821c7b2d8f83ddf61702d36240d9966ec683283adf104aff646e091791a63c032744f5794178f3b4330a93b42415e81ac3c748c5614c3fed167b6b81b49edb9a75a8590a4968346bd5d237dea000105afc41983b2d74224dce51333b1eebb2cab682c63d80b5d35d57e754a92854b6cb6b10af2;
    5'b10101 : xpb = 1024'h82aaee6d47c9be6db58ed32e6f1d688ae959428fc43e661afe630a8a1e88585b11e1507527aa77e00ed7a1fa0d0f8ee78d8c37247e4c803daaaddc8412424e527af09b561a0efe7d72c107baa28cee56c06d537026b1aeffc3acb07688d66c13601901bb8d21d0703e3437f7fcaf0e7d7d78de1ce1ea768cd6aa19813777e51a;
    5'b10110 : xpb = 1024'h2c584f5df1d07b15f255cf39e5bec2118844440f5194fe885adbc2579da5d12a72891ec18ee790a00536a0ed044cbdad22e6b72796b586f4627b1b283d75b3672b7d3dfeb32548fdb79e1f1904e392ebe83f2a0103800d70e7cccdeca7be1c10de532f288c95951f43b9cde45625ca6dd40c80219e0b1a9ed45f6c912f5c58d7;
    5'b10111 : xpb = 1024'h86b2f5a45dc56c86fa22431c6cba62e998a548bfb463376d3531337acfc5f701d6796a86c04b27ee9af3df26dee7fd3d1c5b5f10d1d15df6cae7992aa37b8d2d50591555fbcc90c30f15391a0015fbb20415fa2a6cd498f2c1797d5d80d06ea08b94eebf3cd2525bcfff4aafa76cac87797a0108aa771be118843aa5b02332ff;
    5'b11000 : xpb = 1024'h3060569507cc292f36e93f27e35bbc7037904a3f41b9cfda91a9eb484ee36fd1372138d3278840ae9152de19d6252c02b1b5df13ea3a64ad82b4d7ceceaef24200e5b7fe94e2db4353f25078626ca0472be7d0bb49a2f763e5999ad39fb81e9e09cf1c2c3c46170ad584e09c00e36877d00da30d6697bff316398db5a807a6bc;
    5'b11001 : xpb = 1024'h8abafcdb73c11aa03eb5b30a6a575d4847f14eefa48808bf6bff5c6b810395a89b11849858ebd7fd27101c53b0c06b92ab2a86fd25563bafeb2155d134b4cc0825c18f55dd8a2308ab696a795d9f090d47bea0e4b2f782e5bf464a4478ca712db710dbc2ec82d44761ca5d67522a4a91757b23f47303c1355a5e5bca28ce80e4;
    5'b11010 : xpb = 1024'h34685dcc1dc7d7487b7caf15e0f8b6cee6dc506f31dea12cc878143900210e77fbb952e4c028f0bd1d6f1b46a7fd9a58408507003dbf4266a2ee94755fe8311cd64e31fe76a06d88f04681d7bff5ada26f9077758fc5e156e36667ba97b2212b354b092febf698f6674ff353aba10681cc0ec5f92f2465475813aeda20b2f4a1;
    5'b11011 : xpb = 1024'h8ec3041289bcc8b9834922f867f457a6f73d551f94acda11a2cd855c3241344f5fa99ea9f18c880bb32c59808298d9e839f9aee978db19690b5b1277c5ee0ae2fb2a0955bf47b54e47bd9bd8bb2816688b67479ef91a6cd8bd13172b70c473bae28cc8c69c335632f395701efce7e89b717c46e03b9066899c387ceea179cec9;
    5'b11100 : xpb = 1024'h3870650333c38561c0101f03de95b12d9628569f2203727eff463d29b15ead1ec0516cf658c9a0cba98b587379d608adcf542eec9144201fc328511bf1216ff7abb6abfe585dffce8c9ab3371d7ebafdb3391e2fd5e8cb49e13334a18fac23b860c6f6339ba71ae1f91b060b565ea48bc80fe8e4f7b10a9b99edcffe995e4286;
    5'b11101 : xpb = 1024'h92cb0b499fb876d2c7dc92e665915205a6895b4f84d1ab63d99bae4ce37ed2f62441b8bb8a2d381a3f4896ad5471483dc8c8d6d5cc5ff7222b94cf1e572749bdd0928355a1054793e411cd3818b123c3cf0fee593f3d56cbbadfe41268be76480e08b5ca4be3d81e856082d6a7a586a56d7d69cc041d0bddde129e131a251cae;
    5'b11110 : xpb = 1024'h3c786c3a49bf337b04a38ef1dc32ab8c45745ccf122843d13614661a629c4bc584e98707f16a50da35a795a04bae77035e2356d8e4c8fdd8e3620dc2825aaed2811f25fe3a1b921428eee4967b07c858f6e1c4ea1c0bb53cdf00018887a626458c42e3374b579ccd8ae618c3011c4295c4110bd0c03dafefdbc7f1231209906b;
    5'b11111 : xpb = 1024'h96d31280b5b424ec0c7002d4632e4c6455d5617f74f67cb61069d73d94bc719ce8d9d2cd22cde828cb64d3da2649b6935797fec21fe4d4db4bce8bc4e8608898a5fafd5582c2d9d98065fe97763a311f12b89513856040beb8acb0f960b878d53984a2cdfb945a0a172b958e526324af697e8cb7cca9b1321fecbf3792d06a93;
    endcase
end

endmodule

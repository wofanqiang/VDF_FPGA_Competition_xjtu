module xpb_5_335
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'hfcb6443ee8def236b4e17ac653e5c4e11fde1f45d3e14d29306a7a5f3fa8bf541188add86dc64a76d2118a1fba5407031cb39b614184e6141f93cfa41803a3375ceca9c3972e8eee9b75d70aaf7178d37896586a9f7709b985610c5f33c407533a1012d44dde9c196a95551da422bd79d49c320d6108b2c940c95f238bf31d6;
    5'b00010 : xpb = 1024'h1f96c887dd1bde46d69c2f58ca7cb89c23fbc3e8ba7c29a5260d4f4be7f517ea823115bb0db8c94eda423143f74a80e06396736c28309cc283f279f483007466eb9d953872e5d1ddd36ebae155ee2f1a6f12cb0d53eee13730ac218be67880ea6742025a89bbd3832d52aaa3b48457af3a938641ac21165928192be4717e63ac;
    5'b00011 : xpb = 1024'h2f622ccbcba9cd6a41ea47052fbb14ea35f9a5dd17ba3e77b913f6f1dbefa3dfc349a09894952df6476349e5f2efc1509561ad223c48eb23c5ebb6eec480ae9a616c5fd4ac58baccbd26185200e546a7a69c3093fde651d2c9023251d9b4c15f9ae30387ce99bd44c3fbfff58ec68386d7dd49628231a185bc25c1d6aa3d9582;
    5'b00100 : xpb = 1024'h3f2d910fba37bc8dad385eb194f9713847f787d174f8534a4c1a9e97cfea2fd504622b761b71929db4846287ee9501c0c72ce6d85061398507e4f3e90600e8cdd73b2a70e5cba3bba6dd75c2abdc5e34de25961aa7ddc26e61584317ccf101d4ce8404b51377a7065aa555476908af5e75270c8358422cb2503257c8e2fcc758;
    5'b00101 : xpb = 1024'h4ef8f553a8c5abb11886765dfa37cd8659f569c5d236681cdf21463dc3e4bbca457ab653a24df74521a57b29ea3a4230f8f8208e647987e649de30e3478123014d09f50d1f3e8caa9094d33356d375c215aefba151d53309f9ae53ddc02d424a022505e2585590c7f14eaa99434adb361270cfa42e52b7dee43eedbb1bbbf92e;
    5'b00110 : xpb = 1024'h5ec4599797539ad483d48e0a5f7629d46bf34bba2f747cef7227ede3b7df47bf86934131292a5bec8ec693cbe5df82a12ac35a447891d6478bd76ddd89015d34c2d8bfa958b175997a4c30a401ca8d4f4d386127fbcca3a5920464a3b36982bf35c6070f9d337a8987f7ffeb1d8d070dafba92c50463430b784b83ad547b2b04;
    5'b00111 : xpb = 1024'h6e8fbddb85e189f7ef22a5b6c4b486227df12dae8cb291c2052e9589abd9d3b4c7abcc0eb006c093fbe7ac6de184c3115c8e93fa8caa24a8cdd0aad7ca81976838a78a4592245e8864038e14acc1a4dc84c1c6aea5c414412a5a7569a6a5c3346967083ce211644b1ea1553cf7cf32e54d0455e5da73ce380c58199f8d3a5cda;
    5'b01000 : xpb = 1024'h7e5b221f746f791b5a70bd6329f2e2708fef0fa2e9f0a69498353d2f9fd45faa08c456ec36e3253b6908c50fdd2a03818e59cdb0a0c2730a0fc9e7d20c01d19bae7654e1cb9747774dbaeb8557b8bc69bc4b2c354fbb84dcc2b0862f99e203a99d08096a26ef4e0cb54aaa8ed2115ebcea4e1906b0845964a064af91c5f98eb0;
    5'b01001 : xpb = 1024'h8e26866362fd683ec5bed50f8f313ebea1ecf197472ebb672b3be4d593ceeb9f49dce1c9bdbf89e2d629ddb1d8cf43f1c0250766b4dac16b51c324cc4d820bcf24451f7e050a3066377248f602afd3f6f3d491bbf9b2f5785b0696f58d1e441ed0a90a976bcd37ce4bf3ffe0ac538a948797dc278694e49134714583feb8c086;
    5'b01010 : xpb = 1024'h9df1eaa7518b5762310cecbbf46f9b0cb3ead38ba46cd039be428c7b87c977948af56ca7449bee8a434af653d4748461f1f0411cc8f30fcc93bc61c68f0246029a13ea1a3e7d19552129a666ada6eb842b5df742a3aa6613f35ca7bb805a8494044a0bc4b0ab218fe29d55328695b66c24e19f485ca56fbdc87ddb763777f25c;
    5'b01011 : xpb = 1024'hadbd4eeb401946859c5b046859adf75ac5e8b58001aae50c514934217bc40389cc0df784cb785331b06c0ef5d019c4d223bb7ad2dd0b5e2dd5b59ec0d08280360fe2b4b677f002440ae103d7589e031162e75cc94da1d6af8bb2b8817396c50937eb0cf1f5890b517946aa8460d7e243c22b626932b5faea5c8a716870372432;
    5'b01100 : xpb = 1024'hcdb6dd96cb900e03ca3a43dae920c57667094438971596766732271bcbbe27709de04e9882e394a7e2ee850e860f477f16c8ca2ce70dc43670f9c5cd73045b811624aa401d1edede1fe5ea56ab9566da66bc8b76b131a3a6e7c374caca862ec3c847bf5899dfc85893018f74349e7f2109b46a7b87b28e6aa278c562013ef9d;
    5'b01101 : xpb = 1024'h1ca6d21d5b46f003a7f1bbea13d068a5786e7637e6af6e39f979ca17b0b66e6c4af68fc70f0a9df1eb5000f2e40634e82337c658e2892aa4a908d95718b07feb873115403b44d6dccbb5bc1615b06dfaddf52e3e150a8ad606d248129fe4a36170257d22ce7be6471fd96e491d8c13c9ade509c88e8bb4133e34224858d32173;
    5'b01110 : xpb = 1024'h2c72366149d4df27133fd396790ec4f38a6c582c43ed830c8c8071bda4b0fa618c0f1aa495e7029958711994dfab75585503000ef6a17905eb0216515a30ba1efcffdfdc74b7bfcbb56d1986c0a78588157e93c4bf01fb719f2858d89320e3d6a3c67e501359d008b682c39af7ce3fa14b2ecce9649c3f3fd240b83a91925349;
    5'b01111 : xpb = 1024'h3c3d9aa53862ce4a7e8deb42de4d21419c6a3a20a12b97df1f87196398ab8656cd27a5821cc36740c5923236db50b5c886ce39c50ab9c7672cfb534b9bb0f45272ceaa78ae2aa8ba9f2476f76b9e9d154d07f94b68f96c0d377e699e865d244bd7677f7d5837b9ca4d2c18ecd2106b78e878900a3aacca6c664d4e2cca51851f;
    5'b10000 : xpb = 1024'h4c08fee926f0bd6de9dc02ef438b7d8fae681c14fe69acb1b28dc1098ca6124c0e40305fa39fcbe832b34ad8d6f5f638b899737b1ed215c86ef49045dd312e85e89d7514e79d91a988dbd4681695b4a284915ed212f0dca8cfd47a64799964c10b0880aa9d15a38be3d56e3eac52975085c2532b10bd5598fa59e41f0310b6f5;
    5'b10001 : xpb = 1024'h5bd4632d157eac91552a1a9ba8c9d9ddc065fe095ba7c184459468af80a09e414f58bb3d2a7c308f9fd4637ad29b36a8ea64ad3132ea6429b0edcd401eb168b95e6c3fb121107a98729331d8c18ccc2fbc1ac458bce84d44682a8b2a6cd5a5363ea981d7e1f38d4d7a7ec3908694c328230c164be6cde0c58e667a113bcfe8cb;
    5'b10010 : xpb = 1024'h6b9fc771040c9bb4c07832480e08362bd263dffdb8e5d656d89b1055749b2a369071461ab15895370cf57c1cce4077191c2fe6e74702b28af2e70a3a6031a2ecd43b0a4d5a8363875c4a8f496c83e3bcf3a429df66dfbde000809bf06011e5ab724a830526d1770f112818e260d6eeffc055d96cbcde6bf222731003748f1aa1;
    5'b10011 : xpb = 1024'h7b6b2bb4f29a8ad82bc649f473469279e461c1f21623eb296ba1b7fb6895b62bd189d0f83834f9de7a1694bec9e5b7894dfb209d5b1b00ec34e04734a1b1dd204a09d4e993f64c764601ecba177afb4a2b2d8f6610d72e7b98d6acb6534e2620a5eb84326baf60d0a7d16e343b191ad75d9f9c8d92eef71eb67fa5f5ad4e4c77;
    5'b10100 : xpb = 1024'h8b368ff8e12879fb971461a0d884eec7f65fa3e67361fffbfea85fa15c90422112a25bd5bf115e85e737ad60c58af7f97fc65a536f334f4d76d9842ee3321753bfd89f85cd6935652fb94a2ac27212d762b6f4ecbace9f17312cbd7c468a6695d98c855fb08d4a923e7ac386155b46aefae95fae68ff824b4a8c3be7e60d7e4d;
    5'b10101 : xpb = 1024'h9b01f43ccfb6691f0262794d3dc34b16085d85dad0a014ce91af0747508ace1653bae6b345edc32d5458c602c1303869b1919409834b9daeb8d2c12924b2518735a76a2206dc1e541970a79b6d692a649a405a7364c60fb2c982ce4239c6a70b0d2d868cf56b3453d52418d7ef9d7286983322cf3f100d77de98d1da1eccb023;
    5'b10110 : xpb = 1024'haacd5880be4458426db090f9a301a7641a5b67cf2dde29a124b5aeed44855a0b94d37190ccca27d4c179dea4bcd578d9e35ccdbf9763ec0ffacbfe2366328bbaab7634be404f07430328050c186041f1d1c9bffa0ebd804e61d8df082d02e78040ce87ba3a491e156bcd6e29c9df9e5e357ce5f0152098a472a567cc578be1f9;
    5'b10111 : xpb = 1024'h9eb776eeae4129d0df930cef7e5bc60bae34692b5a49dfc39df9d3d857d38f8d2a37ef589800ded8f3cb7ffd51ca87fb10ddf8f88c96a258c25fbbf6ce0513cacf5caabca30f2ecda455fda2a7b954e154e2be82c2ec3d944a25dd3661485634567f6bdce5e0f497bb6dc9cac51a40c83ecca2e9ae5c6a0c04282ba0768ad64;
    5'b11000 : xpb = 1024'h19b6dbb2d97201c07947487b5d2418aecce1288712e2b2cecce644e37977c4ee13bc09d3105c7294fc5dd0a1d0c1e8efe2d919459ce1b886ce1f38b9ae608b7022c4954803a3dbdbc3fcbd4ad572acdb4cd7916ed6263474dcf86e995950c5d87908f7eb133bf90b126031ee8693cfe421368d4f70f651cd544f18ac4027df3a;
    5'b11001 : xpb = 1024'h29823ff6c7fff0e3e4956027c26274fcdedf0a7b7020c7a15fecec896d7250e354d494b09738d73c697ee943cc67296014a452fbb0fa06e8101875b3efe0c5a398935fe43d16c4caadb41abb8069c4688460f6f5801da510754e7f5f4c8d064daca9f9185819e2cca909874060d5fbbbbe8050704706dcf9e85bae9e78e71110;
    5'b11010 : xpb = 1024'h394da43ab68de0074fe377d427a0d14af0dcec6fcd5edc73f2f3942f616cdcd895ed1f8e1e153be3d6a001e5c80c69d0466f8cb1c51255495211b2ae3160ffd70e622a807689adb9976b782c2b60dbf5bbea5c7c2a1515ac0da490253fc946c2e04afa459cf7cc8e3fb2dc923b1827935bca13911d1768267c684490b1a642e6;
    5'b11011 : xpb = 1024'h4919087ea51bcf2abb318f808cdf2d9902dace642a9cf14685fa3bd5556768cdd705aa6ba4f1a08b43c11a87c3b1aa40783ac667d92aa3aa940aefa872e13a0a8430f51caffc96a88122d59cd657f382f373c202d40c8647a5faa0eb3305873813ebfb72e1d5b64fd65c31e4155a536af913d6b1f327f3531074da82ea6574bc;
    5'b11100 : xpb = 1024'h58e46cc293a9be4e267fa72cf21d89e714d8b05887db06191900e37b4961f4c3181e35492bce0532b0e23329bf56eab0aa06001ded42f20bd6042ca2b461743df9ffbfb8e96f7f976ada330d814f0b102afd27897e03f6e33e50b1b12641c7ad478cfca026b3a0116d058735ef9c7f42965d99d2c9387e7fa48170752324a692;
    5'b11101 : xpb = 1024'h68afd1068237ad7191cdbed9575be63526d6924ce5191aebac078b213d5c80b85936c026b2aa69da1e034bcbbafc2b20dbd139d4015b406d17fd699cf5e1ae716fce8a5522e268865491907e2c46229d62868d1027fb677ed6a6c277197e08227b2dfdcd6b9189d303aedc87c9deab1a33a75cf39f4909ac388e06675be3d868;
    5'b11110 : xpb = 1024'h787b354a70c59c94fd1bd685bc9a428338d4744142572fbe3f0e32c731570cad9a4f4b043986ce818b24646db6a16b910d9c738a15738ece59f6a6973761e8a4e59d54f15c5551753e48edeed73d3a2a9a0ff296d1f2d81a6efcd33d0cba4897aecefefab06f73949a5831d9a420d6f1d0f12014755994d8cc9a9c5994a30a3e;
    5'b11111 : xpb = 1024'h8846998e5f538bb86869ee3221d89ed14ad256359f954490d214da6d255198a2db67d5e1c0633328f8457d0fb246ac013f67ad40298bdd2f9befe39178e222d85b6c1f8d95c83a6428004b5f823451b7d199581d7bea48b60752e402fff6890ce2700027f54d5d563101872b7e6302c96e3ae3354b6a200560a7324bcd623c14;
    endcase
end

endmodule

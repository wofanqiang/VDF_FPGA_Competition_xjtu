module xpb_5_500
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h8161751d699a0e02d8122eec870b47098e38f9a12884613e2143e137aa812ebf4424a18f41b0ff29024d583a1f83c9a38dbf63b3e7128576e8b2023e466bb6e0baea2374a6942ac490b11a2195653812ced61588bcb60ab5150083e1dff110acd34d1276e8a7d183fc0a10d705e6f1cb0e739284f41c281ad5381cc13320140f;
    5'b00010 : xpb = 1024'h5215a4e51145e73ce51ee601fdbc46c1aafbf0117b912204c4ab0919a1ffb0768500c5a5b93b7fc3653c712d5ba9827cb7649f81ab723aa220c4c51e5204f9100185123a9d9758440ec831a091eeabf4a9a73178ece5e859747475c905b77ec7779292c42086aa7a71543acf13fdbd6cce0d462797ecf3056400be7ddd5dc1b3;
    5'b00011 : xpb = 1024'h22c9d4acb8f1c076f22b9d17746d4679c7bee681ce9de2cb681230fb997e322dc5dce9bc30c6005dc82b8a2097cf3b55e109db4f6fd1efcd58d787fe5d9e3b3f48200100949a85c38cdf491f8e781fd684784d691d15c5fdd3e867b02b7dece21bd8131158658370e69e64c72214890e8da6f9ca3bbdbdeff2c9603a879b6f57;
    5'b00100 : xpb = 1024'ha42b49ca228bce79ca3dcc03fb788d8355f7e022f72244098956123343ff60ed0a018b4b7276ff86ca78e25ab75304f96ec93f0356e4754441898a3ca409f220030a24753b2eb0881d90634123dd57e9534e62f1d9cbd0b2e8e8eb920b6efd8eef252588410d54f4e2a8759e27fb7ad99c1a8c4f2fd9e60ac8017cfbbabb8366;
    5'b00101 : xpb = 1024'h74df7991ca37a7b3d74a831972298d3b72bad6934a2f04d02cbd3a153b7de2a44addaf61ea0180212d67fb4df378bdd2986e7ad11b442a6f799c4d1cafa3344f49a5133b3231de079ba77ac02066cbcb2e1f7ee209fbae57485cdd7931356ba9936aa5d578ec2deb57f29f963612467b5bb43ff1d3aab0f556ca1eb864f9310a;
    5'b00110 : xpb = 1024'h4593a95971e380ede4573a2ee8da8cf38f7dcd039d3bc596d02461f732fc645b8bb9d378618c00bb905714412f9e76abc213b69edfa3df9ab1af0ffcbb3c767e9040020129350b8719be923f1cf03fad08f09ad23a2b8bfba7d0cf6056fbd9c437b02622b0cb06e1cd3cc98e4429121d1b4df394777b7bdfe592c0750f36deae;
    5'b00111 : xpb = 1024'h1647d921198f5a27f163f1445f8b8cabac40c373f048865d738b89d92a7ae612cc95f78ed9168155f3462d346bc42f84ebb8f26ca40394c5e9c1d2dcc6d5b8add6daf0c72038390697d5a9be1979b38ee3c1b6c26a5b69a00744c1477cc247dedbf5a66fe8a9dfd84286f386523fddbedae7a7371b4c46ca745b6231b9748c52;
    5'b01000 : xpb = 1024'h97a94e3e8329682ac9762030e696d3b53a79bd1518cce79b94cf6b10d4fc14d210ba991e1ac7807ef593856e8b47f928797856208b161a3cd273d51b0d416f8e91c5143bc6cc63cb2886c3dfaedeeba1b297cc4b271174551c4545295cb3588baf42b8e6d151b15c3e91045d5826cf89e95b39bc0f686ee549937ef2ec94a061;
    5'b01001 : xpb = 1024'h685d7e062ad54164d682d7465d47d36d573cb3856bd9a862383692f2cc7a96895196bd349252011958829e61c76db201a31d91ee4f75cf680a8697fb18dab1bdd8600301bdcf914aa69ddb5eab685f838d68e83b574151f97bb937108279c6a65388393409308a52b3db2e55663d9b2ba8f4ed5eb33939cfd85c20af96d24e05;
    5'b01010 : xpb = 1024'h3911adcdd2811a9ee38f8e5bd3f8d32573ffa9f5bee66928db9dbad4c3f918409272e14b09dc81b3bb71b75503936adaccc2cdbc13d5849342995adb2473f3ed1efaf1c7b4d2beca24b4f2dda7f1d365683a042b87712f9ddb2d28f7a84034c0f7cdb981410f63492925584d745466cd688ea101570a04ba6724c26c410ffba9;
    5'b01011 : xpb = 1024'h9c5dd957a2cf3d8f09c45714aa9d2dd90c2a06611f329ef7f04e2b6bb7799f7d34f05618167024e1e60d0483fb923b3f6680989d83539be7aac1dbb300d361c6595e08dabd5ec49a2cc0a5ca47b4747430b201bb7a10d423aa11adece06a2db9c1339ce78ee3c3f9e6f8245826b326f282854a3fadacfa4f5ed6428eb4da94d;
    5'b01100 : xpb = 1024'h8b2752b2e3c701dbc8ae745dd1b519e71efb9a073a778b2da048c3ee65f8c8b71773a6f0c318017720ae28825f3ced5784276d3dbf47bf35635e1ff97678ecfd20800402526a170e337d247e39e07f5a11e135a4745717f74fa19ec0adf7b3886f604c4561960dc39a79931c8852243a369be728eef6f7bfcb2580ea1e6dbd5c;
    5'b01101 : xpb = 1024'h5bdb827a8b72db15d5bb2b734866199f3bbe90778d844bf443afebd05d774a6e584fcb073aa28211839d41759b62a630adcca90b83a774609b70e2d982122f2c671af2c8496d448db1943bfd3669f33becb25194a486f59baf1590a7d3be21a313a5cc929974e6ba0fc3bd149668efdbf6359acb92c7c2aa59ee22a6c8ab6b00;
    5'b01110 : xpb = 1024'h2c8fb242331eb44fe2c7e288bf171957588186e7e0910cbae71713b254f5cc25992bef1db22d02abe68c5a68d7885f09d771e4d94807298bd383a5b98dab715badb5e18e4070720d2fab537c32f3671dc7836d84d4b6d3400e89828ef9848fbdb7eb4cdfd153bfb0850de70ca47fbb7db5cf4e6e36988d94e8b6c46372e918a4;
    5'b01111 : xpb = 1024'hadf1275f9cb8c252bada117546226060e6ba808909156df9085af4e9ff76fae4dd5090acf3de01d4e8d9b2a2f70c28ad6531488d2f19af02bc35a7f7d417283c68a00502e7049cd1c05c6d9dc8589f309659830d916cddf5238a0670d975a06a8b385f56b9fb91348117f7e3aa66ad48c442e0f32ab4b5afbdeee124a6092cb3;
    5'b10000 : xpb = 1024'h7ea5572744649b8cc7e6c88abcd36019037d76f95c222ebfabc21ccbf6f57c9c1e2cb4c36b68826f4bc8cb963331e1868ed6845af379642df4486ad7dfb06a6baf3af3c8de07ca513e73851cc4e21312712a9efdc19cbb9982fdf857ff3c0e852f7ddfa3f1da6a2af66221dbb87d78ea83dc9495ce85809a4cb782e15046da57;
    5'b10001 : xpb = 1024'h4f5986eeec1074c6d4f37fa033845fd120406d69af2eef864f2944adee73fe535f08d8d9e2f30309aeb7e4896f579a5fb87bc028b7d919592c5b2db7eb49ac9af5d5e28ed50af7d0bc8a9c9bc16b86f44bfbbaedf1cc993de271ea3f25027c9fd3c35ff129b943216bac4bd3c694448c4376483872564b84db80249dfa8487fb;
    5'b10010 : xpb = 1024'h200db6b693bc4e00e20036b5aa355f893d0363da023bb04cf2906c8fe5f2800a9fe4fcf05a7d83a411a6fd7cab7d5338e220fbf67c38ce84646df097f6e2eeca3c70d154cc0e25503aa1b41abdf4fad626ccd6de21fc76e241e5dc264ac8eaba7808e03e61981c17e0f675cbd4ab102e030ffbdb1627166f6a48c65aa4c2359f;
    5'b10011 : xpb = 1024'ha16f2bd3fd565c03ba1265a23140a692cb3c5d7b2ac0118b13d44dc79073aec9e4099e7f9c2e82cd13f455b6cb011cdc6fe05faa634b53fb4d1ff2d63d4ea5aaf75af4c972a25014cb52ce3c535a32e8f5a2ec66deb2819756e660082ab9fb674b55f2b54a3fed9bdd0086a2da9201f911838e600a433e8a3f80e31bd7e249ae;
    5'b10100 : xpb = 1024'h72235b9ba502353dc71f1cb7a7f1a64ae7ff53eb7dccd251b73b75a987f2308124e5c29613b9036776e36eaa0726d5b599859b7827ab09268532b5b648e7e7da3df5e38f69a57d944969e5bb4fe3a6cad07408570ee25f3bb65a51ef50806981ef9b7302821ec692524ab09ae8a8cd9ad11d4202ae140974ce4984d8821ff752;
    5'b10101 : xpb = 1024'h42d78b634cae0e77d42bd3cd1ea2a60304c24a5bd0d993185aa29d8b7f70b23865c1e6ac8b438401d9d2879d434c8e8ec32ad745ec0abe51bd45789654812a098490d25560a8ab13c780fd3a4c6d1aacab4524473f123ce015ce43d67646d79c93e0f34fb9fd9f88c794da92f6bf993c90b6f5a551e4d45f5d1226952c5da4f6;
    5'b10110 : xpb = 1024'h138bbb2af459e7b1e1388ae29553a5bb218540cc23e653defe09c56d76ef33efa69e0ac302ce049c3cc1a0907f724767ecd01313b06a737cf5583b76601a6c38cb2bc11b57abd893459814b948f68e8e861640376f421a84754235bd9c0d45b73826739cf1dc787f3cdf048b04d664de5050a947f5b59f49ebdac851d69b529a;
    5'b10111 : xpb = 1024'h94ed30485df3f5b4b94ab9cf1c5eecc4afbe3a6d4c6ab51d1f4da6a5217062aeeac2ac52447f03c53f0ef8ca9ef6110b7a8f76c7977cf8f3de0a3db4a68623198615e48ffe400357d6492edade5bc6a154ec55c02bf825398a42b99f7bfe56640b738613da844a0338e915620abd56a95ec43bcce9d1c764c112e51309bb66a9;
    5'b11000 : xpb = 1024'h65a16010059fceeec65770e4930fec7ccc8130dd9f7775e3c2b4ce8718eee4662b9ed068bc09845fa1fe11bddb1bc9e4a434b2955bdcae1f161d0094b21f6548ccb0d355f54330d754604659dae53a832fbd71b05c2802dde9b6ab86a1c4c47eafb90661126322f9ae333f5a18d4224b1e5def6f8da2924f4fdb86cfb3f9144d;
    5'b11001 : xpb = 1024'h36558fd7ad4ba828d36427fa09c0ec34e944274df28436aa661bf669106d661d6c7af47f339404fa04ed2ab1174182bdcdd9ee63203c634a4e2fc374bdb8a778134bc21bec465e56d2775dd8d76eae650a8e8da08c57e082492a9d6dc78b329953fe86ae4a41fbf0237d695226eaedecddf7a31231735d39dea4288c5e36c1f1;
    5'b11010 : xpb = 1024'h709bf9f54f78162e070df0f8071ebed06071dbe4590f77109831e4b07ebe7d4ad571895ab1e859467dc43a453673b96f77f2a30e49c187586428654c951e9a759e6b0e1e3498bd6508e7557d3f82246e55fa990bc87be26a89e8f54ed51a0b3f84406fb8220d4e698c7934a3501b98e9d9156b4d54428246d6cca4908746f95;
    5'b11011 : xpb = 1024'h886b34bcbe918f65b8830dfc077d32f69440175f6e1558af2ac6ff82b26d1693f17bba24eccf84bd6a299bde72eb053a853e8de4cbae9dec6ef488930fbda08814d0d45689ddb69ae13f8f79695d5a59b435bf19793dc8dbbd9f1336cd42b160cb9119726ac8a66a94d1a4213ae8ab59ac04e939c960503f42a4e70a3b9483a4;
    5'b11100 : xpb = 1024'h591f6484663d689fc58fc5117e2e32aeb1030dcfc1221975ce2e2764a9eb984b3257de3b645a0557cd18b4d1af10be13aee3c9b2900e5317a7074b731b56e2b75b6bc31c80e0e41a5f56a6f865e6ce3b8f06db09a96da6801d13051df3091f7b6fd699bfa2a77f610a1bce1948ff76fb6b9e9cdc6d311b29d16d88c6e5d23148;
    5'b11101 : xpb = 1024'h29d3944c0de941d9d29c7c26f4df3266cdc60440142eda3c71954f46a16a1a0273340251dbe485f23007cdc4eb3676ecd8890580546e0842df1a0e5326f024e6a206b1e277e41199dd6dbe776270421d69d7f6f9d99d84247c86f70518cf8d96141c1a0cda8658577f65f8115716429d2b38507f1101e61460362a83900fdeec;
    5'b11110 : xpb = 1024'hab35096977834fdcaaaeab137bea79705bfefde13cb33b7a92d9307e4beb48c1b758a3e11d95851b325525ff0aba4090664869343b808db9c7cc10916d5bdbc75cf0d5571e783c5e6e1ed898f7d57a3038ae0c8296538ed991877ae6f8c09e42e7692c83c32e29db7b7008e85cfd346839abe304051e0e2f356e4744c32ff2fb;
    5'b11111 : xpb = 1024'h7be939311f2f2916b7bb6228f29b792878c1f4518fbffc41364058604369ca78f834c7f7952005b595443ef246dff9698feda501ffe042e4ffded37178f51df6a38bc41d157b69ddec35f017f45eee12137f2872c6836c7df0fb6cce1e870c5d8baeacd0fb0d02d1f0ba32e06b140009f94596a6a8eed919c436e9016d6da09f;
    endcase
end

endmodule

module compressor_array_12_8_1033
(
    input  [11:0] col_in_0,
    input  [11:0] col_in_1,
    input  [11:0] col_in_2,
    input  [11:0] col_in_3,
    input  [11:0] col_in_4,
    input  [11:0] col_in_5,
    input  [11:0] col_in_6,
    input  [11:0] col_in_7,
    input  [11:0] col_in_8,
    input  [11:0] col_in_9,
    input  [11:0] col_in_10,
    input  [11:0] col_in_11,
    input  [11:0] col_in_12,
    input  [11:0] col_in_13,
    input  [11:0] col_in_14,
    input  [11:0] col_in_15,
    input  [11:0] col_in_16,
    input  [11:0] col_in_17,
    input  [11:0] col_in_18,
    input  [11:0] col_in_19,
    input  [11:0] col_in_20,
    input  [11:0] col_in_21,
    input  [11:0] col_in_22,
    input  [11:0] col_in_23,
    input  [11:0] col_in_24,
    input  [11:0] col_in_25,
    input  [11:0] col_in_26,
    input  [11:0] col_in_27,
    input  [11:0] col_in_28,
    input  [11:0] col_in_29,
    input  [11:0] col_in_30,
    input  [11:0] col_in_31,
    input  [11:0] col_in_32,
    input  [11:0] col_in_33,
    input  [11:0] col_in_34,
    input  [11:0] col_in_35,
    input  [11:0] col_in_36,
    input  [11:0] col_in_37,
    input  [11:0] col_in_38,
    input  [11:0] col_in_39,
    input  [11:0] col_in_40,
    input  [11:0] col_in_41,
    input  [11:0] col_in_42,
    input  [11:0] col_in_43,
    input  [11:0] col_in_44,
    input  [11:0] col_in_45,
    input  [11:0] col_in_46,
    input  [11:0] col_in_47,
    input  [11:0] col_in_48,
    input  [11:0] col_in_49,
    input  [11:0] col_in_50,
    input  [11:0] col_in_51,
    input  [11:0] col_in_52,
    input  [11:0] col_in_53,
    input  [11:0] col_in_54,
    input  [11:0] col_in_55,
    input  [11:0] col_in_56,
    input  [11:0] col_in_57,
    input  [11:0] col_in_58,
    input  [11:0] col_in_59,
    input  [11:0] col_in_60,
    input  [11:0] col_in_61,
    input  [11:0] col_in_62,
    input  [11:0] col_in_63,
    input  [11:0] col_in_64,
    input  [11:0] col_in_65,
    input  [11:0] col_in_66,
    input  [11:0] col_in_67,
    input  [11:0] col_in_68,
    input  [11:0] col_in_69,
    input  [11:0] col_in_70,
    input  [11:0] col_in_71,
    input  [11:0] col_in_72,
    input  [11:0] col_in_73,
    input  [11:0] col_in_74,
    input  [11:0] col_in_75,
    input  [11:0] col_in_76,
    input  [11:0] col_in_77,
    input  [11:0] col_in_78,
    input  [11:0] col_in_79,
    input  [11:0] col_in_80,
    input  [11:0] col_in_81,
    input  [11:0] col_in_82,
    input  [11:0] col_in_83,
    input  [11:0] col_in_84,
    input  [11:0] col_in_85,
    input  [11:0] col_in_86,
    input  [11:0] col_in_87,
    input  [11:0] col_in_88,
    input  [11:0] col_in_89,
    input  [11:0] col_in_90,
    input  [11:0] col_in_91,
    input  [11:0] col_in_92,
    input  [11:0] col_in_93,
    input  [11:0] col_in_94,
    input  [11:0] col_in_95,
    input  [11:0] col_in_96,
    input  [11:0] col_in_97,
    input  [11:0] col_in_98,
    input  [11:0] col_in_99,
    input  [11:0] col_in_100,
    input  [11:0] col_in_101,
    input  [11:0] col_in_102,
    input  [11:0] col_in_103,
    input  [11:0] col_in_104,
    input  [11:0] col_in_105,
    input  [11:0] col_in_106,
    input  [11:0] col_in_107,
    input  [11:0] col_in_108,
    input  [11:0] col_in_109,
    input  [11:0] col_in_110,
    input  [11:0] col_in_111,
    input  [11:0] col_in_112,
    input  [11:0] col_in_113,
    input  [11:0] col_in_114,
    input  [11:0] col_in_115,
    input  [11:0] col_in_116,
    input  [11:0] col_in_117,
    input  [11:0] col_in_118,
    input  [11:0] col_in_119,
    input  [11:0] col_in_120,
    input  [11:0] col_in_121,
    input  [11:0] col_in_122,
    input  [11:0] col_in_123,
    input  [11:0] col_in_124,
    input  [11:0] col_in_125,
    input  [11:0] col_in_126,
    input  [11:0] col_in_127,
    input  [11:0] col_in_128,
    input  [11:0] col_in_129,
    input  [11:0] col_in_130,
    input  [11:0] col_in_131,
    input  [11:0] col_in_132,
    input  [11:0] col_in_133,
    input  [11:0] col_in_134,
    input  [11:0] col_in_135,
    input  [11:0] col_in_136,
    input  [11:0] col_in_137,
    input  [11:0] col_in_138,
    input  [11:0] col_in_139,
    input  [11:0] col_in_140,
    input  [11:0] col_in_141,
    input  [11:0] col_in_142,
    input  [11:0] col_in_143,
    input  [11:0] col_in_144,
    input  [11:0] col_in_145,
    input  [11:0] col_in_146,
    input  [11:0] col_in_147,
    input  [11:0] col_in_148,
    input  [11:0] col_in_149,
    input  [11:0] col_in_150,
    input  [11:0] col_in_151,
    input  [11:0] col_in_152,
    input  [11:0] col_in_153,
    input  [11:0] col_in_154,
    input  [11:0] col_in_155,
    input  [11:0] col_in_156,
    input  [11:0] col_in_157,
    input  [11:0] col_in_158,
    input  [11:0] col_in_159,
    input  [11:0] col_in_160,
    input  [11:0] col_in_161,
    input  [11:0] col_in_162,
    input  [11:0] col_in_163,
    input  [11:0] col_in_164,
    input  [11:0] col_in_165,
    input  [11:0] col_in_166,
    input  [11:0] col_in_167,
    input  [11:0] col_in_168,
    input  [11:0] col_in_169,
    input  [11:0] col_in_170,
    input  [11:0] col_in_171,
    input  [11:0] col_in_172,
    input  [11:0] col_in_173,
    input  [11:0] col_in_174,
    input  [11:0] col_in_175,
    input  [11:0] col_in_176,
    input  [11:0] col_in_177,
    input  [11:0] col_in_178,
    input  [11:0] col_in_179,
    input  [11:0] col_in_180,
    input  [11:0] col_in_181,
    input  [11:0] col_in_182,
    input  [11:0] col_in_183,
    input  [11:0] col_in_184,
    input  [11:0] col_in_185,
    input  [11:0] col_in_186,
    input  [11:0] col_in_187,
    input  [11:0] col_in_188,
    input  [11:0] col_in_189,
    input  [11:0] col_in_190,
    input  [11:0] col_in_191,
    input  [11:0] col_in_192,
    input  [11:0] col_in_193,
    input  [11:0] col_in_194,
    input  [11:0] col_in_195,
    input  [11:0] col_in_196,
    input  [11:0] col_in_197,
    input  [11:0] col_in_198,
    input  [11:0] col_in_199,
    input  [11:0] col_in_200,
    input  [11:0] col_in_201,
    input  [11:0] col_in_202,
    input  [11:0] col_in_203,
    input  [11:0] col_in_204,
    input  [11:0] col_in_205,
    input  [11:0] col_in_206,
    input  [11:0] col_in_207,
    input  [11:0] col_in_208,
    input  [11:0] col_in_209,
    input  [11:0] col_in_210,
    input  [11:0] col_in_211,
    input  [11:0] col_in_212,
    input  [11:0] col_in_213,
    input  [11:0] col_in_214,
    input  [11:0] col_in_215,
    input  [11:0] col_in_216,
    input  [11:0] col_in_217,
    input  [11:0] col_in_218,
    input  [11:0] col_in_219,
    input  [11:0] col_in_220,
    input  [11:0] col_in_221,
    input  [11:0] col_in_222,
    input  [11:0] col_in_223,
    input  [11:0] col_in_224,
    input  [11:0] col_in_225,
    input  [11:0] col_in_226,
    input  [11:0] col_in_227,
    input  [11:0] col_in_228,
    input  [11:0] col_in_229,
    input  [11:0] col_in_230,
    input  [11:0] col_in_231,
    input  [11:0] col_in_232,
    input  [11:0] col_in_233,
    input  [11:0] col_in_234,
    input  [11:0] col_in_235,
    input  [11:0] col_in_236,
    input  [11:0] col_in_237,
    input  [11:0] col_in_238,
    input  [11:0] col_in_239,
    input  [11:0] col_in_240,
    input  [11:0] col_in_241,
    input  [11:0] col_in_242,
    input  [11:0] col_in_243,
    input  [11:0] col_in_244,
    input  [11:0] col_in_245,
    input  [11:0] col_in_246,
    input  [11:0] col_in_247,
    input  [11:0] col_in_248,
    input  [11:0] col_in_249,
    input  [11:0] col_in_250,
    input  [11:0] col_in_251,
    input  [11:0] col_in_252,
    input  [11:0] col_in_253,
    input  [11:0] col_in_254,
    input  [11:0] col_in_255,
    input  [11:0] col_in_256,
    input  [11:0] col_in_257,
    input  [11:0] col_in_258,
    input  [11:0] col_in_259,
    input  [11:0] col_in_260,
    input  [11:0] col_in_261,
    input  [11:0] col_in_262,
    input  [11:0] col_in_263,
    input  [11:0] col_in_264,
    input  [11:0] col_in_265,
    input  [11:0] col_in_266,
    input  [11:0] col_in_267,
    input  [11:0] col_in_268,
    input  [11:0] col_in_269,
    input  [11:0] col_in_270,
    input  [11:0] col_in_271,
    input  [11:0] col_in_272,
    input  [11:0] col_in_273,
    input  [11:0] col_in_274,
    input  [11:0] col_in_275,
    input  [11:0] col_in_276,
    input  [11:0] col_in_277,
    input  [11:0] col_in_278,
    input  [11:0] col_in_279,
    input  [11:0] col_in_280,
    input  [11:0] col_in_281,
    input  [11:0] col_in_282,
    input  [11:0] col_in_283,
    input  [11:0] col_in_284,
    input  [11:0] col_in_285,
    input  [11:0] col_in_286,
    input  [11:0] col_in_287,
    input  [11:0] col_in_288,
    input  [11:0] col_in_289,
    input  [11:0] col_in_290,
    input  [11:0] col_in_291,
    input  [11:0] col_in_292,
    input  [11:0] col_in_293,
    input  [11:0] col_in_294,
    input  [11:0] col_in_295,
    input  [11:0] col_in_296,
    input  [11:0] col_in_297,
    input  [11:0] col_in_298,
    input  [11:0] col_in_299,
    input  [11:0] col_in_300,
    input  [11:0] col_in_301,
    input  [11:0] col_in_302,
    input  [11:0] col_in_303,
    input  [11:0] col_in_304,
    input  [11:0] col_in_305,
    input  [11:0] col_in_306,
    input  [11:0] col_in_307,
    input  [11:0] col_in_308,
    input  [11:0] col_in_309,
    input  [11:0] col_in_310,
    input  [11:0] col_in_311,
    input  [11:0] col_in_312,
    input  [11:0] col_in_313,
    input  [11:0] col_in_314,
    input  [11:0] col_in_315,
    input  [11:0] col_in_316,
    input  [11:0] col_in_317,
    input  [11:0] col_in_318,
    input  [11:0] col_in_319,
    input  [11:0] col_in_320,
    input  [11:0] col_in_321,
    input  [11:0] col_in_322,
    input  [11:0] col_in_323,
    input  [11:0] col_in_324,
    input  [11:0] col_in_325,
    input  [11:0] col_in_326,
    input  [11:0] col_in_327,
    input  [11:0] col_in_328,
    input  [11:0] col_in_329,
    input  [11:0] col_in_330,
    input  [11:0] col_in_331,
    input  [11:0] col_in_332,
    input  [11:0] col_in_333,
    input  [11:0] col_in_334,
    input  [11:0] col_in_335,
    input  [11:0] col_in_336,
    input  [11:0] col_in_337,
    input  [11:0] col_in_338,
    input  [11:0] col_in_339,
    input  [11:0] col_in_340,
    input  [11:0] col_in_341,
    input  [11:0] col_in_342,
    input  [11:0] col_in_343,
    input  [11:0] col_in_344,
    input  [11:0] col_in_345,
    input  [11:0] col_in_346,
    input  [11:0] col_in_347,
    input  [11:0] col_in_348,
    input  [11:0] col_in_349,
    input  [11:0] col_in_350,
    input  [11:0] col_in_351,
    input  [11:0] col_in_352,
    input  [11:0] col_in_353,
    input  [11:0] col_in_354,
    input  [11:0] col_in_355,
    input  [11:0] col_in_356,
    input  [11:0] col_in_357,
    input  [11:0] col_in_358,
    input  [11:0] col_in_359,
    input  [11:0] col_in_360,
    input  [11:0] col_in_361,
    input  [11:0] col_in_362,
    input  [11:0] col_in_363,
    input  [11:0] col_in_364,
    input  [11:0] col_in_365,
    input  [11:0] col_in_366,
    input  [11:0] col_in_367,
    input  [11:0] col_in_368,
    input  [11:0] col_in_369,
    input  [11:0] col_in_370,
    input  [11:0] col_in_371,
    input  [11:0] col_in_372,
    input  [11:0] col_in_373,
    input  [11:0] col_in_374,
    input  [11:0] col_in_375,
    input  [11:0] col_in_376,
    input  [11:0] col_in_377,
    input  [11:0] col_in_378,
    input  [11:0] col_in_379,
    input  [11:0] col_in_380,
    input  [11:0] col_in_381,
    input  [11:0] col_in_382,
    input  [11:0] col_in_383,
    input  [11:0] col_in_384,
    input  [11:0] col_in_385,
    input  [11:0] col_in_386,
    input  [11:0] col_in_387,
    input  [11:0] col_in_388,
    input  [11:0] col_in_389,
    input  [11:0] col_in_390,
    input  [11:0] col_in_391,
    input  [11:0] col_in_392,
    input  [11:0] col_in_393,
    input  [11:0] col_in_394,
    input  [11:0] col_in_395,
    input  [11:0] col_in_396,
    input  [11:0] col_in_397,
    input  [11:0] col_in_398,
    input  [11:0] col_in_399,
    input  [11:0] col_in_400,
    input  [11:0] col_in_401,
    input  [11:0] col_in_402,
    input  [11:0] col_in_403,
    input  [11:0] col_in_404,
    input  [11:0] col_in_405,
    input  [11:0] col_in_406,
    input  [11:0] col_in_407,
    input  [11:0] col_in_408,
    input  [11:0] col_in_409,
    input  [11:0] col_in_410,
    input  [11:0] col_in_411,
    input  [11:0] col_in_412,
    input  [11:0] col_in_413,
    input  [11:0] col_in_414,
    input  [11:0] col_in_415,
    input  [11:0] col_in_416,
    input  [11:0] col_in_417,
    input  [11:0] col_in_418,
    input  [11:0] col_in_419,
    input  [11:0] col_in_420,
    input  [11:0] col_in_421,
    input  [11:0] col_in_422,
    input  [11:0] col_in_423,
    input  [11:0] col_in_424,
    input  [11:0] col_in_425,
    input  [11:0] col_in_426,
    input  [11:0] col_in_427,
    input  [11:0] col_in_428,
    input  [11:0] col_in_429,
    input  [11:0] col_in_430,
    input  [11:0] col_in_431,
    input  [11:0] col_in_432,
    input  [11:0] col_in_433,
    input  [11:0] col_in_434,
    input  [11:0] col_in_435,
    input  [11:0] col_in_436,
    input  [11:0] col_in_437,
    input  [11:0] col_in_438,
    input  [11:0] col_in_439,
    input  [11:0] col_in_440,
    input  [11:0] col_in_441,
    input  [11:0] col_in_442,
    input  [11:0] col_in_443,
    input  [11:0] col_in_444,
    input  [11:0] col_in_445,
    input  [11:0] col_in_446,
    input  [11:0] col_in_447,
    input  [11:0] col_in_448,
    input  [11:0] col_in_449,
    input  [11:0] col_in_450,
    input  [11:0] col_in_451,
    input  [11:0] col_in_452,
    input  [11:0] col_in_453,
    input  [11:0] col_in_454,
    input  [11:0] col_in_455,
    input  [11:0] col_in_456,
    input  [11:0] col_in_457,
    input  [11:0] col_in_458,
    input  [11:0] col_in_459,
    input  [11:0] col_in_460,
    input  [11:0] col_in_461,
    input  [11:0] col_in_462,
    input  [11:0] col_in_463,
    input  [11:0] col_in_464,
    input  [11:0] col_in_465,
    input  [11:0] col_in_466,
    input  [11:0] col_in_467,
    input  [11:0] col_in_468,
    input  [11:0] col_in_469,
    input  [11:0] col_in_470,
    input  [11:0] col_in_471,
    input  [11:0] col_in_472,
    input  [11:0] col_in_473,
    input  [11:0] col_in_474,
    input  [11:0] col_in_475,
    input  [11:0] col_in_476,
    input  [11:0] col_in_477,
    input  [11:0] col_in_478,
    input  [11:0] col_in_479,
    input  [11:0] col_in_480,
    input  [11:0] col_in_481,
    input  [11:0] col_in_482,
    input  [11:0] col_in_483,
    input  [11:0] col_in_484,
    input  [11:0] col_in_485,
    input  [11:0] col_in_486,
    input  [11:0] col_in_487,
    input  [11:0] col_in_488,
    input  [11:0] col_in_489,
    input  [11:0] col_in_490,
    input  [11:0] col_in_491,
    input  [11:0] col_in_492,
    input  [11:0] col_in_493,
    input  [11:0] col_in_494,
    input  [11:0] col_in_495,
    input  [11:0] col_in_496,
    input  [11:0] col_in_497,
    input  [11:0] col_in_498,
    input  [11:0] col_in_499,
    input  [11:0] col_in_500,
    input  [11:0] col_in_501,
    input  [11:0] col_in_502,
    input  [11:0] col_in_503,
    input  [11:0] col_in_504,
    input  [11:0] col_in_505,
    input  [11:0] col_in_506,
    input  [11:0] col_in_507,
    input  [11:0] col_in_508,
    input  [11:0] col_in_509,
    input  [11:0] col_in_510,
    input  [11:0] col_in_511,
    input  [11:0] col_in_512,
    input  [11:0] col_in_513,
    input  [11:0] col_in_514,
    input  [11:0] col_in_515,
    input  [11:0] col_in_516,
    input  [11:0] col_in_517,
    input  [11:0] col_in_518,
    input  [11:0] col_in_519,
    input  [11:0] col_in_520,
    input  [11:0] col_in_521,
    input  [11:0] col_in_522,
    input  [11:0] col_in_523,
    input  [11:0] col_in_524,
    input  [11:0] col_in_525,
    input  [11:0] col_in_526,
    input  [11:0] col_in_527,
    input  [11:0] col_in_528,
    input  [11:0] col_in_529,
    input  [11:0] col_in_530,
    input  [11:0] col_in_531,
    input  [11:0] col_in_532,
    input  [11:0] col_in_533,
    input  [11:0] col_in_534,
    input  [11:0] col_in_535,
    input  [11:0] col_in_536,
    input  [11:0] col_in_537,
    input  [11:0] col_in_538,
    input  [11:0] col_in_539,
    input  [11:0] col_in_540,
    input  [11:0] col_in_541,
    input  [11:0] col_in_542,
    input  [11:0] col_in_543,
    input  [11:0] col_in_544,
    input  [11:0] col_in_545,
    input  [11:0] col_in_546,
    input  [11:0] col_in_547,
    input  [11:0] col_in_548,
    input  [11:0] col_in_549,
    input  [11:0] col_in_550,
    input  [11:0] col_in_551,
    input  [11:0] col_in_552,
    input  [11:0] col_in_553,
    input  [11:0] col_in_554,
    input  [11:0] col_in_555,
    input  [11:0] col_in_556,
    input  [11:0] col_in_557,
    input  [11:0] col_in_558,
    input  [11:0] col_in_559,
    input  [11:0] col_in_560,
    input  [11:0] col_in_561,
    input  [11:0] col_in_562,
    input  [11:0] col_in_563,
    input  [11:0] col_in_564,
    input  [11:0] col_in_565,
    input  [11:0] col_in_566,
    input  [11:0] col_in_567,
    input  [11:0] col_in_568,
    input  [11:0] col_in_569,
    input  [11:0] col_in_570,
    input  [11:0] col_in_571,
    input  [11:0] col_in_572,
    input  [11:0] col_in_573,
    input  [11:0] col_in_574,
    input  [11:0] col_in_575,
    input  [11:0] col_in_576,
    input  [11:0] col_in_577,
    input  [11:0] col_in_578,
    input  [11:0] col_in_579,
    input  [11:0] col_in_580,
    input  [11:0] col_in_581,
    input  [11:0] col_in_582,
    input  [11:0] col_in_583,
    input  [11:0] col_in_584,
    input  [11:0] col_in_585,
    input  [11:0] col_in_586,
    input  [11:0] col_in_587,
    input  [11:0] col_in_588,
    input  [11:0] col_in_589,
    input  [11:0] col_in_590,
    input  [11:0] col_in_591,
    input  [11:0] col_in_592,
    input  [11:0] col_in_593,
    input  [11:0] col_in_594,
    input  [11:0] col_in_595,
    input  [11:0] col_in_596,
    input  [11:0] col_in_597,
    input  [11:0] col_in_598,
    input  [11:0] col_in_599,
    input  [11:0] col_in_600,
    input  [11:0] col_in_601,
    input  [11:0] col_in_602,
    input  [11:0] col_in_603,
    input  [11:0] col_in_604,
    input  [11:0] col_in_605,
    input  [11:0] col_in_606,
    input  [11:0] col_in_607,
    input  [11:0] col_in_608,
    input  [11:0] col_in_609,
    input  [11:0] col_in_610,
    input  [11:0] col_in_611,
    input  [11:0] col_in_612,
    input  [11:0] col_in_613,
    input  [11:0] col_in_614,
    input  [11:0] col_in_615,
    input  [11:0] col_in_616,
    input  [11:0] col_in_617,
    input  [11:0] col_in_618,
    input  [11:0] col_in_619,
    input  [11:0] col_in_620,
    input  [11:0] col_in_621,
    input  [11:0] col_in_622,
    input  [11:0] col_in_623,
    input  [11:0] col_in_624,
    input  [11:0] col_in_625,
    input  [11:0] col_in_626,
    input  [11:0] col_in_627,
    input  [11:0] col_in_628,
    input  [11:0] col_in_629,
    input  [11:0] col_in_630,
    input  [11:0] col_in_631,
    input  [11:0] col_in_632,
    input  [11:0] col_in_633,
    input  [11:0] col_in_634,
    input  [11:0] col_in_635,
    input  [11:0] col_in_636,
    input  [11:0] col_in_637,
    input  [11:0] col_in_638,
    input  [11:0] col_in_639,
    input  [11:0] col_in_640,
    input  [11:0] col_in_641,
    input  [11:0] col_in_642,
    input  [11:0] col_in_643,
    input  [11:0] col_in_644,
    input  [11:0] col_in_645,
    input  [11:0] col_in_646,
    input  [11:0] col_in_647,
    input  [11:0] col_in_648,
    input  [11:0] col_in_649,
    input  [11:0] col_in_650,
    input  [11:0] col_in_651,
    input  [11:0] col_in_652,
    input  [11:0] col_in_653,
    input  [11:0] col_in_654,
    input  [11:0] col_in_655,
    input  [11:0] col_in_656,
    input  [11:0] col_in_657,
    input  [11:0] col_in_658,
    input  [11:0] col_in_659,
    input  [11:0] col_in_660,
    input  [11:0] col_in_661,
    input  [11:0] col_in_662,
    input  [11:0] col_in_663,
    input  [11:0] col_in_664,
    input  [11:0] col_in_665,
    input  [11:0] col_in_666,
    input  [11:0] col_in_667,
    input  [11:0] col_in_668,
    input  [11:0] col_in_669,
    input  [11:0] col_in_670,
    input  [11:0] col_in_671,
    input  [11:0] col_in_672,
    input  [11:0] col_in_673,
    input  [11:0] col_in_674,
    input  [11:0] col_in_675,
    input  [11:0] col_in_676,
    input  [11:0] col_in_677,
    input  [11:0] col_in_678,
    input  [11:0] col_in_679,
    input  [11:0] col_in_680,
    input  [11:0] col_in_681,
    input  [11:0] col_in_682,
    input  [11:0] col_in_683,
    input  [11:0] col_in_684,
    input  [11:0] col_in_685,
    input  [11:0] col_in_686,
    input  [11:0] col_in_687,
    input  [11:0] col_in_688,
    input  [11:0] col_in_689,
    input  [11:0] col_in_690,
    input  [11:0] col_in_691,
    input  [11:0] col_in_692,
    input  [11:0] col_in_693,
    input  [11:0] col_in_694,
    input  [11:0] col_in_695,
    input  [11:0] col_in_696,
    input  [11:0] col_in_697,
    input  [11:0] col_in_698,
    input  [11:0] col_in_699,
    input  [11:0] col_in_700,
    input  [11:0] col_in_701,
    input  [11:0] col_in_702,
    input  [11:0] col_in_703,
    input  [11:0] col_in_704,
    input  [11:0] col_in_705,
    input  [11:0] col_in_706,
    input  [11:0] col_in_707,
    input  [11:0] col_in_708,
    input  [11:0] col_in_709,
    input  [11:0] col_in_710,
    input  [11:0] col_in_711,
    input  [11:0] col_in_712,
    input  [11:0] col_in_713,
    input  [11:0] col_in_714,
    input  [11:0] col_in_715,
    input  [11:0] col_in_716,
    input  [11:0] col_in_717,
    input  [11:0] col_in_718,
    input  [11:0] col_in_719,
    input  [11:0] col_in_720,
    input  [11:0] col_in_721,
    input  [11:0] col_in_722,
    input  [11:0] col_in_723,
    input  [11:0] col_in_724,
    input  [11:0] col_in_725,
    input  [11:0] col_in_726,
    input  [11:0] col_in_727,
    input  [11:0] col_in_728,
    input  [11:0] col_in_729,
    input  [11:0] col_in_730,
    input  [11:0] col_in_731,
    input  [11:0] col_in_732,
    input  [11:0] col_in_733,
    input  [11:0] col_in_734,
    input  [11:0] col_in_735,
    input  [11:0] col_in_736,
    input  [11:0] col_in_737,
    input  [11:0] col_in_738,
    input  [11:0] col_in_739,
    input  [11:0] col_in_740,
    input  [11:0] col_in_741,
    input  [11:0] col_in_742,
    input  [11:0] col_in_743,
    input  [11:0] col_in_744,
    input  [11:0] col_in_745,
    input  [11:0] col_in_746,
    input  [11:0] col_in_747,
    input  [11:0] col_in_748,
    input  [11:0] col_in_749,
    input  [11:0] col_in_750,
    input  [11:0] col_in_751,
    input  [11:0] col_in_752,
    input  [11:0] col_in_753,
    input  [11:0] col_in_754,
    input  [11:0] col_in_755,
    input  [11:0] col_in_756,
    input  [11:0] col_in_757,
    input  [11:0] col_in_758,
    input  [11:0] col_in_759,
    input  [11:0] col_in_760,
    input  [11:0] col_in_761,
    input  [11:0] col_in_762,
    input  [11:0] col_in_763,
    input  [11:0] col_in_764,
    input  [11:0] col_in_765,
    input  [11:0] col_in_766,
    input  [11:0] col_in_767,
    input  [11:0] col_in_768,
    input  [11:0] col_in_769,
    input  [11:0] col_in_770,
    input  [11:0] col_in_771,
    input  [11:0] col_in_772,
    input  [11:0] col_in_773,
    input  [11:0] col_in_774,
    input  [11:0] col_in_775,
    input  [11:0] col_in_776,
    input  [11:0] col_in_777,
    input  [11:0] col_in_778,
    input  [11:0] col_in_779,
    input  [11:0] col_in_780,
    input  [11:0] col_in_781,
    input  [11:0] col_in_782,
    input  [11:0] col_in_783,
    input  [11:0] col_in_784,
    input  [11:0] col_in_785,
    input  [11:0] col_in_786,
    input  [11:0] col_in_787,
    input  [11:0] col_in_788,
    input  [11:0] col_in_789,
    input  [11:0] col_in_790,
    input  [11:0] col_in_791,
    input  [11:0] col_in_792,
    input  [11:0] col_in_793,
    input  [11:0] col_in_794,
    input  [11:0] col_in_795,
    input  [11:0] col_in_796,
    input  [11:0] col_in_797,
    input  [11:0] col_in_798,
    input  [11:0] col_in_799,
    input  [11:0] col_in_800,
    input  [11:0] col_in_801,
    input  [11:0] col_in_802,
    input  [11:0] col_in_803,
    input  [11:0] col_in_804,
    input  [11:0] col_in_805,
    input  [11:0] col_in_806,
    input  [11:0] col_in_807,
    input  [11:0] col_in_808,
    input  [11:0] col_in_809,
    input  [11:0] col_in_810,
    input  [11:0] col_in_811,
    input  [11:0] col_in_812,
    input  [11:0] col_in_813,
    input  [11:0] col_in_814,
    input  [11:0] col_in_815,
    input  [11:0] col_in_816,
    input  [11:0] col_in_817,
    input  [11:0] col_in_818,
    input  [11:0] col_in_819,
    input  [11:0] col_in_820,
    input  [11:0] col_in_821,
    input  [11:0] col_in_822,
    input  [11:0] col_in_823,
    input  [11:0] col_in_824,
    input  [11:0] col_in_825,
    input  [11:0] col_in_826,
    input  [11:0] col_in_827,
    input  [11:0] col_in_828,
    input  [11:0] col_in_829,
    input  [11:0] col_in_830,
    input  [11:0] col_in_831,
    input  [11:0] col_in_832,
    input  [11:0] col_in_833,
    input  [11:0] col_in_834,
    input  [11:0] col_in_835,
    input  [11:0] col_in_836,
    input  [11:0] col_in_837,
    input  [11:0] col_in_838,
    input  [11:0] col_in_839,
    input  [11:0] col_in_840,
    input  [11:0] col_in_841,
    input  [11:0] col_in_842,
    input  [11:0] col_in_843,
    input  [11:0] col_in_844,
    input  [11:0] col_in_845,
    input  [11:0] col_in_846,
    input  [11:0] col_in_847,
    input  [11:0] col_in_848,
    input  [11:0] col_in_849,
    input  [11:0] col_in_850,
    input  [11:0] col_in_851,
    input  [11:0] col_in_852,
    input  [11:0] col_in_853,
    input  [11:0] col_in_854,
    input  [11:0] col_in_855,
    input  [11:0] col_in_856,
    input  [11:0] col_in_857,
    input  [11:0] col_in_858,
    input  [11:0] col_in_859,
    input  [11:0] col_in_860,
    input  [11:0] col_in_861,
    input  [11:0] col_in_862,
    input  [11:0] col_in_863,
    input  [11:0] col_in_864,
    input  [11:0] col_in_865,
    input  [11:0] col_in_866,
    input  [11:0] col_in_867,
    input  [11:0] col_in_868,
    input  [11:0] col_in_869,
    input  [11:0] col_in_870,
    input  [11:0] col_in_871,
    input  [11:0] col_in_872,
    input  [11:0] col_in_873,
    input  [11:0] col_in_874,
    input  [11:0] col_in_875,
    input  [11:0] col_in_876,
    input  [11:0] col_in_877,
    input  [11:0] col_in_878,
    input  [11:0] col_in_879,
    input  [11:0] col_in_880,
    input  [11:0] col_in_881,
    input  [11:0] col_in_882,
    input  [11:0] col_in_883,
    input  [11:0] col_in_884,
    input  [11:0] col_in_885,
    input  [11:0] col_in_886,
    input  [11:0] col_in_887,
    input  [11:0] col_in_888,
    input  [11:0] col_in_889,
    input  [11:0] col_in_890,
    input  [11:0] col_in_891,
    input  [11:0] col_in_892,
    input  [11:0] col_in_893,
    input  [11:0] col_in_894,
    input  [11:0] col_in_895,
    input  [11:0] col_in_896,
    input  [11:0] col_in_897,
    input  [11:0] col_in_898,
    input  [11:0] col_in_899,
    input  [11:0] col_in_900,
    input  [11:0] col_in_901,
    input  [11:0] col_in_902,
    input  [11:0] col_in_903,
    input  [11:0] col_in_904,
    input  [11:0] col_in_905,
    input  [11:0] col_in_906,
    input  [11:0] col_in_907,
    input  [11:0] col_in_908,
    input  [11:0] col_in_909,
    input  [11:0] col_in_910,
    input  [11:0] col_in_911,
    input  [11:0] col_in_912,
    input  [11:0] col_in_913,
    input  [11:0] col_in_914,
    input  [11:0] col_in_915,
    input  [11:0] col_in_916,
    input  [11:0] col_in_917,
    input  [11:0] col_in_918,
    input  [11:0] col_in_919,
    input  [11:0] col_in_920,
    input  [11:0] col_in_921,
    input  [11:0] col_in_922,
    input  [11:0] col_in_923,
    input  [11:0] col_in_924,
    input  [11:0] col_in_925,
    input  [11:0] col_in_926,
    input  [11:0] col_in_927,
    input  [11:0] col_in_928,
    input  [11:0] col_in_929,
    input  [11:0] col_in_930,
    input  [11:0] col_in_931,
    input  [11:0] col_in_932,
    input  [11:0] col_in_933,
    input  [11:0] col_in_934,
    input  [11:0] col_in_935,
    input  [11:0] col_in_936,
    input  [11:0] col_in_937,
    input  [11:0] col_in_938,
    input  [11:0] col_in_939,
    input  [11:0] col_in_940,
    input  [11:0] col_in_941,
    input  [11:0] col_in_942,
    input  [11:0] col_in_943,
    input  [11:0] col_in_944,
    input  [11:0] col_in_945,
    input  [11:0] col_in_946,
    input  [11:0] col_in_947,
    input  [11:0] col_in_948,
    input  [11:0] col_in_949,
    input  [11:0] col_in_950,
    input  [11:0] col_in_951,
    input  [11:0] col_in_952,
    input  [11:0] col_in_953,
    input  [11:0] col_in_954,
    input  [11:0] col_in_955,
    input  [11:0] col_in_956,
    input  [11:0] col_in_957,
    input  [11:0] col_in_958,
    input  [11:0] col_in_959,
    input  [11:0] col_in_960,
    input  [11:0] col_in_961,
    input  [11:0] col_in_962,
    input  [11:0] col_in_963,
    input  [11:0] col_in_964,
    input  [11:0] col_in_965,
    input  [11:0] col_in_966,
    input  [11:0] col_in_967,
    input  [11:0] col_in_968,
    input  [11:0] col_in_969,
    input  [11:0] col_in_970,
    input  [11:0] col_in_971,
    input  [11:0] col_in_972,
    input  [11:0] col_in_973,
    input  [11:0] col_in_974,
    input  [11:0] col_in_975,
    input  [11:0] col_in_976,
    input  [11:0] col_in_977,
    input  [11:0] col_in_978,
    input  [11:0] col_in_979,
    input  [11:0] col_in_980,
    input  [11:0] col_in_981,
    input  [11:0] col_in_982,
    input  [11:0] col_in_983,
    input  [11:0] col_in_984,
    input  [11:0] col_in_985,
    input  [11:0] col_in_986,
    input  [11:0] col_in_987,
    input  [11:0] col_in_988,
    input  [11:0] col_in_989,
    input  [11:0] col_in_990,
    input  [11:0] col_in_991,
    input  [11:0] col_in_992,
    input  [11:0] col_in_993,
    input  [11:0] col_in_994,
    input  [11:0] col_in_995,
    input  [11:0] col_in_996,
    input  [11:0] col_in_997,
    input  [11:0] col_in_998,
    input  [11:0] col_in_999,
    input  [11:0] col_in_1000,
    input  [11:0] col_in_1001,
    input  [11:0] col_in_1002,
    input  [11:0] col_in_1003,
    input  [11:0] col_in_1004,
    input  [11:0] col_in_1005,
    input  [11:0] col_in_1006,
    input  [11:0] col_in_1007,
    input  [11:0] col_in_1008,
    input  [11:0] col_in_1009,
    input  [11:0] col_in_1010,
    input  [11:0] col_in_1011,
    input  [11:0] col_in_1012,
    input  [11:0] col_in_1013,
    input  [11:0] col_in_1014,
    input  [11:0] col_in_1015,
    input  [11:0] col_in_1016,
    input  [11:0] col_in_1017,
    input  [11:0] col_in_1018,
    input  [11:0] col_in_1019,
    input  [11:0] col_in_1020,
    input  [11:0] col_in_1021,
    input  [11:0] col_in_1022,
    input  [11:0] col_in_1023,
    input  [11:0] col_in_1024,
    input  [11:0] col_in_1025,
    input  [11:0] col_in_1026,
    input  [11:0] col_in_1027,
    input  [11:0] col_in_1028,
    input  [11:0] col_in_1029,
    input  [11:0] col_in_1030,
    input  [11:0] col_in_1031,
    input  [11:0] col_in_1032,

    output [7:0] col_out_0,
    output [7:0] col_out_1,
    output [7:0] col_out_2,
    output [7:0] col_out_3,
    output [7:0] col_out_4,
    output [7:0] col_out_5,
    output [7:0] col_out_6,
    output [7:0] col_out_7,
    output [7:0] col_out_8,
    output [7:0] col_out_9,
    output [7:0] col_out_10,
    output [7:0] col_out_11,
    output [7:0] col_out_12,
    output [7:0] col_out_13,
    output [7:0] col_out_14,
    output [7:0] col_out_15,
    output [7:0] col_out_16,
    output [7:0] col_out_17,
    output [7:0] col_out_18,
    output [7:0] col_out_19,
    output [7:0] col_out_20,
    output [7:0] col_out_21,
    output [7:0] col_out_22,
    output [7:0] col_out_23,
    output [7:0] col_out_24,
    output [7:0] col_out_25,
    output [7:0] col_out_26,
    output [7:0] col_out_27,
    output [7:0] col_out_28,
    output [7:0] col_out_29,
    output [7:0] col_out_30,
    output [7:0] col_out_31,
    output [7:0] col_out_32,
    output [7:0] col_out_33,
    output [7:0] col_out_34,
    output [7:0] col_out_35,
    output [7:0] col_out_36,
    output [7:0] col_out_37,
    output [7:0] col_out_38,
    output [7:0] col_out_39,
    output [7:0] col_out_40,
    output [7:0] col_out_41,
    output [7:0] col_out_42,
    output [7:0] col_out_43,
    output [7:0] col_out_44,
    output [7:0] col_out_45,
    output [7:0] col_out_46,
    output [7:0] col_out_47,
    output [7:0] col_out_48,
    output [7:0] col_out_49,
    output [7:0] col_out_50,
    output [7:0] col_out_51,
    output [7:0] col_out_52,
    output [7:0] col_out_53,
    output [7:0] col_out_54,
    output [7:0] col_out_55,
    output [7:0] col_out_56,
    output [7:0] col_out_57,
    output [7:0] col_out_58,
    output [7:0] col_out_59,
    output [7:0] col_out_60,
    output [7:0] col_out_61,
    output [7:0] col_out_62,
    output [7:0] col_out_63,
    output [7:0] col_out_64,
    output [7:0] col_out_65,
    output [7:0] col_out_66,
    output [7:0] col_out_67,
    output [7:0] col_out_68,
    output [7:0] col_out_69,
    output [7:0] col_out_70,
    output [7:0] col_out_71,
    output [7:0] col_out_72,
    output [7:0] col_out_73,
    output [7:0] col_out_74,
    output [7:0] col_out_75,
    output [7:0] col_out_76,
    output [7:0] col_out_77,
    output [7:0] col_out_78,
    output [7:0] col_out_79,
    output [7:0] col_out_80,
    output [7:0] col_out_81,
    output [7:0] col_out_82,
    output [7:0] col_out_83,
    output [7:0] col_out_84,
    output [7:0] col_out_85,
    output [7:0] col_out_86,
    output [7:0] col_out_87,
    output [7:0] col_out_88,
    output [7:0] col_out_89,
    output [7:0] col_out_90,
    output [7:0] col_out_91,
    output [7:0] col_out_92,
    output [7:0] col_out_93,
    output [7:0] col_out_94,
    output [7:0] col_out_95,
    output [7:0] col_out_96,
    output [7:0] col_out_97,
    output [7:0] col_out_98,
    output [7:0] col_out_99,
    output [7:0] col_out_100,
    output [7:0] col_out_101,
    output [7:0] col_out_102,
    output [7:0] col_out_103,
    output [7:0] col_out_104,
    output [7:0] col_out_105,
    output [7:0] col_out_106,
    output [7:0] col_out_107,
    output [7:0] col_out_108,
    output [7:0] col_out_109,
    output [7:0] col_out_110,
    output [7:0] col_out_111,
    output [7:0] col_out_112,
    output [7:0] col_out_113,
    output [7:0] col_out_114,
    output [7:0] col_out_115,
    output [7:0] col_out_116,
    output [7:0] col_out_117,
    output [7:0] col_out_118,
    output [7:0] col_out_119,
    output [7:0] col_out_120,
    output [7:0] col_out_121,
    output [7:0] col_out_122,
    output [7:0] col_out_123,
    output [7:0] col_out_124,
    output [7:0] col_out_125,
    output [7:0] col_out_126,
    output [7:0] col_out_127,
    output [7:0] col_out_128,
    output [7:0] col_out_129,
    output [7:0] col_out_130,
    output [7:0] col_out_131,
    output [7:0] col_out_132,
    output [7:0] col_out_133,
    output [7:0] col_out_134,
    output [7:0] col_out_135,
    output [7:0] col_out_136,
    output [7:0] col_out_137,
    output [7:0] col_out_138,
    output [7:0] col_out_139,
    output [7:0] col_out_140,
    output [7:0] col_out_141,
    output [7:0] col_out_142,
    output [7:0] col_out_143,
    output [7:0] col_out_144,
    output [7:0] col_out_145,
    output [7:0] col_out_146,
    output [7:0] col_out_147,
    output [7:0] col_out_148,
    output [7:0] col_out_149,
    output [7:0] col_out_150,
    output [7:0] col_out_151,
    output [7:0] col_out_152,
    output [7:0] col_out_153,
    output [7:0] col_out_154,
    output [7:0] col_out_155,
    output [7:0] col_out_156,
    output [7:0] col_out_157,
    output [7:0] col_out_158,
    output [7:0] col_out_159,
    output [7:0] col_out_160,
    output [7:0] col_out_161,
    output [7:0] col_out_162,
    output [7:0] col_out_163,
    output [7:0] col_out_164,
    output [7:0] col_out_165,
    output [7:0] col_out_166,
    output [7:0] col_out_167,
    output [7:0] col_out_168,
    output [7:0] col_out_169,
    output [7:0] col_out_170,
    output [7:0] col_out_171,
    output [7:0] col_out_172,
    output [7:0] col_out_173,
    output [7:0] col_out_174,
    output [7:0] col_out_175,
    output [7:0] col_out_176,
    output [7:0] col_out_177,
    output [7:0] col_out_178,
    output [7:0] col_out_179,
    output [7:0] col_out_180,
    output [7:0] col_out_181,
    output [7:0] col_out_182,
    output [7:0] col_out_183,
    output [7:0] col_out_184,
    output [7:0] col_out_185,
    output [7:0] col_out_186,
    output [7:0] col_out_187,
    output [7:0] col_out_188,
    output [7:0] col_out_189,
    output [7:0] col_out_190,
    output [7:0] col_out_191,
    output [7:0] col_out_192,
    output [7:0] col_out_193,
    output [7:0] col_out_194,
    output [7:0] col_out_195,
    output [7:0] col_out_196,
    output [7:0] col_out_197,
    output [7:0] col_out_198,
    output [7:0] col_out_199,
    output [7:0] col_out_200,
    output [7:0] col_out_201,
    output [7:0] col_out_202,
    output [7:0] col_out_203,
    output [7:0] col_out_204,
    output [7:0] col_out_205,
    output [7:0] col_out_206,
    output [7:0] col_out_207,
    output [7:0] col_out_208,
    output [7:0] col_out_209,
    output [7:0] col_out_210,
    output [7:0] col_out_211,
    output [7:0] col_out_212,
    output [7:0] col_out_213,
    output [7:0] col_out_214,
    output [7:0] col_out_215,
    output [7:0] col_out_216,
    output [7:0] col_out_217,
    output [7:0] col_out_218,
    output [7:0] col_out_219,
    output [7:0] col_out_220,
    output [7:0] col_out_221,
    output [7:0] col_out_222,
    output [7:0] col_out_223,
    output [7:0] col_out_224,
    output [7:0] col_out_225,
    output [7:0] col_out_226,
    output [7:0] col_out_227,
    output [7:0] col_out_228,
    output [7:0] col_out_229,
    output [7:0] col_out_230,
    output [7:0] col_out_231,
    output [7:0] col_out_232,
    output [7:0] col_out_233,
    output [7:0] col_out_234,
    output [7:0] col_out_235,
    output [7:0] col_out_236,
    output [7:0] col_out_237,
    output [7:0] col_out_238,
    output [7:0] col_out_239,
    output [7:0] col_out_240,
    output [7:0] col_out_241,
    output [7:0] col_out_242,
    output [7:0] col_out_243,
    output [7:0] col_out_244,
    output [7:0] col_out_245,
    output [7:0] col_out_246,
    output [7:0] col_out_247,
    output [7:0] col_out_248,
    output [7:0] col_out_249,
    output [7:0] col_out_250,
    output [7:0] col_out_251,
    output [7:0] col_out_252,
    output [7:0] col_out_253,
    output [7:0] col_out_254,
    output [7:0] col_out_255,
    output [7:0] col_out_256,
    output [7:0] col_out_257,
    output [7:0] col_out_258,
    output [7:0] col_out_259,
    output [7:0] col_out_260,
    output [7:0] col_out_261,
    output [7:0] col_out_262,
    output [7:0] col_out_263,
    output [7:0] col_out_264,
    output [7:0] col_out_265,
    output [7:0] col_out_266,
    output [7:0] col_out_267,
    output [7:0] col_out_268,
    output [7:0] col_out_269,
    output [7:0] col_out_270,
    output [7:0] col_out_271,
    output [7:0] col_out_272,
    output [7:0] col_out_273,
    output [7:0] col_out_274,
    output [7:0] col_out_275,
    output [7:0] col_out_276,
    output [7:0] col_out_277,
    output [7:0] col_out_278,
    output [7:0] col_out_279,
    output [7:0] col_out_280,
    output [7:0] col_out_281,
    output [7:0] col_out_282,
    output [7:0] col_out_283,
    output [7:0] col_out_284,
    output [7:0] col_out_285,
    output [7:0] col_out_286,
    output [7:0] col_out_287,
    output [7:0] col_out_288,
    output [7:0] col_out_289,
    output [7:0] col_out_290,
    output [7:0] col_out_291,
    output [7:0] col_out_292,
    output [7:0] col_out_293,
    output [7:0] col_out_294,
    output [7:0] col_out_295,
    output [7:0] col_out_296,
    output [7:0] col_out_297,
    output [7:0] col_out_298,
    output [7:0] col_out_299,
    output [7:0] col_out_300,
    output [7:0] col_out_301,
    output [7:0] col_out_302,
    output [7:0] col_out_303,
    output [7:0] col_out_304,
    output [7:0] col_out_305,
    output [7:0] col_out_306,
    output [7:0] col_out_307,
    output [7:0] col_out_308,
    output [7:0] col_out_309,
    output [7:0] col_out_310,
    output [7:0] col_out_311,
    output [7:0] col_out_312,
    output [7:0] col_out_313,
    output [7:0] col_out_314,
    output [7:0] col_out_315,
    output [7:0] col_out_316,
    output [7:0] col_out_317,
    output [7:0] col_out_318,
    output [7:0] col_out_319,
    output [7:0] col_out_320,
    output [7:0] col_out_321,
    output [7:0] col_out_322,
    output [7:0] col_out_323,
    output [7:0] col_out_324,
    output [7:0] col_out_325,
    output [7:0] col_out_326,
    output [7:0] col_out_327,
    output [7:0] col_out_328,
    output [7:0] col_out_329,
    output [7:0] col_out_330,
    output [7:0] col_out_331,
    output [7:0] col_out_332,
    output [7:0] col_out_333,
    output [7:0] col_out_334,
    output [7:0] col_out_335,
    output [7:0] col_out_336,
    output [7:0] col_out_337,
    output [7:0] col_out_338,
    output [7:0] col_out_339,
    output [7:0] col_out_340,
    output [7:0] col_out_341,
    output [7:0] col_out_342,
    output [7:0] col_out_343,
    output [7:0] col_out_344,
    output [7:0] col_out_345,
    output [7:0] col_out_346,
    output [7:0] col_out_347,
    output [7:0] col_out_348,
    output [7:0] col_out_349,
    output [7:0] col_out_350,
    output [7:0] col_out_351,
    output [7:0] col_out_352,
    output [7:0] col_out_353,
    output [7:0] col_out_354,
    output [7:0] col_out_355,
    output [7:0] col_out_356,
    output [7:0] col_out_357,
    output [7:0] col_out_358,
    output [7:0] col_out_359,
    output [7:0] col_out_360,
    output [7:0] col_out_361,
    output [7:0] col_out_362,
    output [7:0] col_out_363,
    output [7:0] col_out_364,
    output [7:0] col_out_365,
    output [7:0] col_out_366,
    output [7:0] col_out_367,
    output [7:0] col_out_368,
    output [7:0] col_out_369,
    output [7:0] col_out_370,
    output [7:0] col_out_371,
    output [7:0] col_out_372,
    output [7:0] col_out_373,
    output [7:0] col_out_374,
    output [7:0] col_out_375,
    output [7:0] col_out_376,
    output [7:0] col_out_377,
    output [7:0] col_out_378,
    output [7:0] col_out_379,
    output [7:0] col_out_380,
    output [7:0] col_out_381,
    output [7:0] col_out_382,
    output [7:0] col_out_383,
    output [7:0] col_out_384,
    output [7:0] col_out_385,
    output [7:0] col_out_386,
    output [7:0] col_out_387,
    output [7:0] col_out_388,
    output [7:0] col_out_389,
    output [7:0] col_out_390,
    output [7:0] col_out_391,
    output [7:0] col_out_392,
    output [7:0] col_out_393,
    output [7:0] col_out_394,
    output [7:0] col_out_395,
    output [7:0] col_out_396,
    output [7:0] col_out_397,
    output [7:0] col_out_398,
    output [7:0] col_out_399,
    output [7:0] col_out_400,
    output [7:0] col_out_401,
    output [7:0] col_out_402,
    output [7:0] col_out_403,
    output [7:0] col_out_404,
    output [7:0] col_out_405,
    output [7:0] col_out_406,
    output [7:0] col_out_407,
    output [7:0] col_out_408,
    output [7:0] col_out_409,
    output [7:0] col_out_410,
    output [7:0] col_out_411,
    output [7:0] col_out_412,
    output [7:0] col_out_413,
    output [7:0] col_out_414,
    output [7:0] col_out_415,
    output [7:0] col_out_416,
    output [7:0] col_out_417,
    output [7:0] col_out_418,
    output [7:0] col_out_419,
    output [7:0] col_out_420,
    output [7:0] col_out_421,
    output [7:0] col_out_422,
    output [7:0] col_out_423,
    output [7:0] col_out_424,
    output [7:0] col_out_425,
    output [7:0] col_out_426,
    output [7:0] col_out_427,
    output [7:0] col_out_428,
    output [7:0] col_out_429,
    output [7:0] col_out_430,
    output [7:0] col_out_431,
    output [7:0] col_out_432,
    output [7:0] col_out_433,
    output [7:0] col_out_434,
    output [7:0] col_out_435,
    output [7:0] col_out_436,
    output [7:0] col_out_437,
    output [7:0] col_out_438,
    output [7:0] col_out_439,
    output [7:0] col_out_440,
    output [7:0] col_out_441,
    output [7:0] col_out_442,
    output [7:0] col_out_443,
    output [7:0] col_out_444,
    output [7:0] col_out_445,
    output [7:0] col_out_446,
    output [7:0] col_out_447,
    output [7:0] col_out_448,
    output [7:0] col_out_449,
    output [7:0] col_out_450,
    output [7:0] col_out_451,
    output [7:0] col_out_452,
    output [7:0] col_out_453,
    output [7:0] col_out_454,
    output [7:0] col_out_455,
    output [7:0] col_out_456,
    output [7:0] col_out_457,
    output [7:0] col_out_458,
    output [7:0] col_out_459,
    output [7:0] col_out_460,
    output [7:0] col_out_461,
    output [7:0] col_out_462,
    output [7:0] col_out_463,
    output [7:0] col_out_464,
    output [7:0] col_out_465,
    output [7:0] col_out_466,
    output [7:0] col_out_467,
    output [7:0] col_out_468,
    output [7:0] col_out_469,
    output [7:0] col_out_470,
    output [7:0] col_out_471,
    output [7:0] col_out_472,
    output [7:0] col_out_473,
    output [7:0] col_out_474,
    output [7:0] col_out_475,
    output [7:0] col_out_476,
    output [7:0] col_out_477,
    output [7:0] col_out_478,
    output [7:0] col_out_479,
    output [7:0] col_out_480,
    output [7:0] col_out_481,
    output [7:0] col_out_482,
    output [7:0] col_out_483,
    output [7:0] col_out_484,
    output [7:0] col_out_485,
    output [7:0] col_out_486,
    output [7:0] col_out_487,
    output [7:0] col_out_488,
    output [7:0] col_out_489,
    output [7:0] col_out_490,
    output [7:0] col_out_491,
    output [7:0] col_out_492,
    output [7:0] col_out_493,
    output [7:0] col_out_494,
    output [7:0] col_out_495,
    output [7:0] col_out_496,
    output [7:0] col_out_497,
    output [7:0] col_out_498,
    output [7:0] col_out_499,
    output [7:0] col_out_500,
    output [7:0] col_out_501,
    output [7:0] col_out_502,
    output [7:0] col_out_503,
    output [7:0] col_out_504,
    output [7:0] col_out_505,
    output [7:0] col_out_506,
    output [7:0] col_out_507,
    output [7:0] col_out_508,
    output [7:0] col_out_509,
    output [7:0] col_out_510,
    output [7:0] col_out_511,
    output [7:0] col_out_512,
    output [7:0] col_out_513,
    output [7:0] col_out_514,
    output [7:0] col_out_515,
    output [7:0] col_out_516,
    output [7:0] col_out_517,
    output [7:0] col_out_518,
    output [7:0] col_out_519,
    output [7:0] col_out_520,
    output [7:0] col_out_521,
    output [7:0] col_out_522,
    output [7:0] col_out_523,
    output [7:0] col_out_524,
    output [7:0] col_out_525,
    output [7:0] col_out_526,
    output [7:0] col_out_527,
    output [7:0] col_out_528,
    output [7:0] col_out_529,
    output [7:0] col_out_530,
    output [7:0] col_out_531,
    output [7:0] col_out_532,
    output [7:0] col_out_533,
    output [7:0] col_out_534,
    output [7:0] col_out_535,
    output [7:0] col_out_536,
    output [7:0] col_out_537,
    output [7:0] col_out_538,
    output [7:0] col_out_539,
    output [7:0] col_out_540,
    output [7:0] col_out_541,
    output [7:0] col_out_542,
    output [7:0] col_out_543,
    output [7:0] col_out_544,
    output [7:0] col_out_545,
    output [7:0] col_out_546,
    output [7:0] col_out_547,
    output [7:0] col_out_548,
    output [7:0] col_out_549,
    output [7:0] col_out_550,
    output [7:0] col_out_551,
    output [7:0] col_out_552,
    output [7:0] col_out_553,
    output [7:0] col_out_554,
    output [7:0] col_out_555,
    output [7:0] col_out_556,
    output [7:0] col_out_557,
    output [7:0] col_out_558,
    output [7:0] col_out_559,
    output [7:0] col_out_560,
    output [7:0] col_out_561,
    output [7:0] col_out_562,
    output [7:0] col_out_563,
    output [7:0] col_out_564,
    output [7:0] col_out_565,
    output [7:0] col_out_566,
    output [7:0] col_out_567,
    output [7:0] col_out_568,
    output [7:0] col_out_569,
    output [7:0] col_out_570,
    output [7:0] col_out_571,
    output [7:0] col_out_572,
    output [7:0] col_out_573,
    output [7:0] col_out_574,
    output [7:0] col_out_575,
    output [7:0] col_out_576,
    output [7:0] col_out_577,
    output [7:0] col_out_578,
    output [7:0] col_out_579,
    output [7:0] col_out_580,
    output [7:0] col_out_581,
    output [7:0] col_out_582,
    output [7:0] col_out_583,
    output [7:0] col_out_584,
    output [7:0] col_out_585,
    output [7:0] col_out_586,
    output [7:0] col_out_587,
    output [7:0] col_out_588,
    output [7:0] col_out_589,
    output [7:0] col_out_590,
    output [7:0] col_out_591,
    output [7:0] col_out_592,
    output [7:0] col_out_593,
    output [7:0] col_out_594,
    output [7:0] col_out_595,
    output [7:0] col_out_596,
    output [7:0] col_out_597,
    output [7:0] col_out_598,
    output [7:0] col_out_599,
    output [7:0] col_out_600,
    output [7:0] col_out_601,
    output [7:0] col_out_602,
    output [7:0] col_out_603,
    output [7:0] col_out_604,
    output [7:0] col_out_605,
    output [7:0] col_out_606,
    output [7:0] col_out_607,
    output [7:0] col_out_608,
    output [7:0] col_out_609,
    output [7:0] col_out_610,
    output [7:0] col_out_611,
    output [7:0] col_out_612,
    output [7:0] col_out_613,
    output [7:0] col_out_614,
    output [7:0] col_out_615,
    output [7:0] col_out_616,
    output [7:0] col_out_617,
    output [7:0] col_out_618,
    output [7:0] col_out_619,
    output [7:0] col_out_620,
    output [7:0] col_out_621,
    output [7:0] col_out_622,
    output [7:0] col_out_623,
    output [7:0] col_out_624,
    output [7:0] col_out_625,
    output [7:0] col_out_626,
    output [7:0] col_out_627,
    output [7:0] col_out_628,
    output [7:0] col_out_629,
    output [7:0] col_out_630,
    output [7:0] col_out_631,
    output [7:0] col_out_632,
    output [7:0] col_out_633,
    output [7:0] col_out_634,
    output [7:0] col_out_635,
    output [7:0] col_out_636,
    output [7:0] col_out_637,
    output [7:0] col_out_638,
    output [7:0] col_out_639,
    output [7:0] col_out_640,
    output [7:0] col_out_641,
    output [7:0] col_out_642,
    output [7:0] col_out_643,
    output [7:0] col_out_644,
    output [7:0] col_out_645,
    output [7:0] col_out_646,
    output [7:0] col_out_647,
    output [7:0] col_out_648,
    output [7:0] col_out_649,
    output [7:0] col_out_650,
    output [7:0] col_out_651,
    output [7:0] col_out_652,
    output [7:0] col_out_653,
    output [7:0] col_out_654,
    output [7:0] col_out_655,
    output [7:0] col_out_656,
    output [7:0] col_out_657,
    output [7:0] col_out_658,
    output [7:0] col_out_659,
    output [7:0] col_out_660,
    output [7:0] col_out_661,
    output [7:0] col_out_662,
    output [7:0] col_out_663,
    output [7:0] col_out_664,
    output [7:0] col_out_665,
    output [7:0] col_out_666,
    output [7:0] col_out_667,
    output [7:0] col_out_668,
    output [7:0] col_out_669,
    output [7:0] col_out_670,
    output [7:0] col_out_671,
    output [7:0] col_out_672,
    output [7:0] col_out_673,
    output [7:0] col_out_674,
    output [7:0] col_out_675,
    output [7:0] col_out_676,
    output [7:0] col_out_677,
    output [7:0] col_out_678,
    output [7:0] col_out_679,
    output [7:0] col_out_680,
    output [7:0] col_out_681,
    output [7:0] col_out_682,
    output [7:0] col_out_683,
    output [7:0] col_out_684,
    output [7:0] col_out_685,
    output [7:0] col_out_686,
    output [7:0] col_out_687,
    output [7:0] col_out_688,
    output [7:0] col_out_689,
    output [7:0] col_out_690,
    output [7:0] col_out_691,
    output [7:0] col_out_692,
    output [7:0] col_out_693,
    output [7:0] col_out_694,
    output [7:0] col_out_695,
    output [7:0] col_out_696,
    output [7:0] col_out_697,
    output [7:0] col_out_698,
    output [7:0] col_out_699,
    output [7:0] col_out_700,
    output [7:0] col_out_701,
    output [7:0] col_out_702,
    output [7:0] col_out_703,
    output [7:0] col_out_704,
    output [7:0] col_out_705,
    output [7:0] col_out_706,
    output [7:0] col_out_707,
    output [7:0] col_out_708,
    output [7:0] col_out_709,
    output [7:0] col_out_710,
    output [7:0] col_out_711,
    output [7:0] col_out_712,
    output [7:0] col_out_713,
    output [7:0] col_out_714,
    output [7:0] col_out_715,
    output [7:0] col_out_716,
    output [7:0] col_out_717,
    output [7:0] col_out_718,
    output [7:0] col_out_719,
    output [7:0] col_out_720,
    output [7:0] col_out_721,
    output [7:0] col_out_722,
    output [7:0] col_out_723,
    output [7:0] col_out_724,
    output [7:0] col_out_725,
    output [7:0] col_out_726,
    output [7:0] col_out_727,
    output [7:0] col_out_728,
    output [7:0] col_out_729,
    output [7:0] col_out_730,
    output [7:0] col_out_731,
    output [7:0] col_out_732,
    output [7:0] col_out_733,
    output [7:0] col_out_734,
    output [7:0] col_out_735,
    output [7:0] col_out_736,
    output [7:0] col_out_737,
    output [7:0] col_out_738,
    output [7:0] col_out_739,
    output [7:0] col_out_740,
    output [7:0] col_out_741,
    output [7:0] col_out_742,
    output [7:0] col_out_743,
    output [7:0] col_out_744,
    output [7:0] col_out_745,
    output [7:0] col_out_746,
    output [7:0] col_out_747,
    output [7:0] col_out_748,
    output [7:0] col_out_749,
    output [7:0] col_out_750,
    output [7:0] col_out_751,
    output [7:0] col_out_752,
    output [7:0] col_out_753,
    output [7:0] col_out_754,
    output [7:0] col_out_755,
    output [7:0] col_out_756,
    output [7:0] col_out_757,
    output [7:0] col_out_758,
    output [7:0] col_out_759,
    output [7:0] col_out_760,
    output [7:0] col_out_761,
    output [7:0] col_out_762,
    output [7:0] col_out_763,
    output [7:0] col_out_764,
    output [7:0] col_out_765,
    output [7:0] col_out_766,
    output [7:0] col_out_767,
    output [7:0] col_out_768,
    output [7:0] col_out_769,
    output [7:0] col_out_770,
    output [7:0] col_out_771,
    output [7:0] col_out_772,
    output [7:0] col_out_773,
    output [7:0] col_out_774,
    output [7:0] col_out_775,
    output [7:0] col_out_776,
    output [7:0] col_out_777,
    output [7:0] col_out_778,
    output [7:0] col_out_779,
    output [7:0] col_out_780,
    output [7:0] col_out_781,
    output [7:0] col_out_782,
    output [7:0] col_out_783,
    output [7:0] col_out_784,
    output [7:0] col_out_785,
    output [7:0] col_out_786,
    output [7:0] col_out_787,
    output [7:0] col_out_788,
    output [7:0] col_out_789,
    output [7:0] col_out_790,
    output [7:0] col_out_791,
    output [7:0] col_out_792,
    output [7:0] col_out_793,
    output [7:0] col_out_794,
    output [7:0] col_out_795,
    output [7:0] col_out_796,
    output [7:0] col_out_797,
    output [7:0] col_out_798,
    output [7:0] col_out_799,
    output [7:0] col_out_800,
    output [7:0] col_out_801,
    output [7:0] col_out_802,
    output [7:0] col_out_803,
    output [7:0] col_out_804,
    output [7:0] col_out_805,
    output [7:0] col_out_806,
    output [7:0] col_out_807,
    output [7:0] col_out_808,
    output [7:0] col_out_809,
    output [7:0] col_out_810,
    output [7:0] col_out_811,
    output [7:0] col_out_812,
    output [7:0] col_out_813,
    output [7:0] col_out_814,
    output [7:0] col_out_815,
    output [7:0] col_out_816,
    output [7:0] col_out_817,
    output [7:0] col_out_818,
    output [7:0] col_out_819,
    output [7:0] col_out_820,
    output [7:0] col_out_821,
    output [7:0] col_out_822,
    output [7:0] col_out_823,
    output [7:0] col_out_824,
    output [7:0] col_out_825,
    output [7:0] col_out_826,
    output [7:0] col_out_827,
    output [7:0] col_out_828,
    output [7:0] col_out_829,
    output [7:0] col_out_830,
    output [7:0] col_out_831,
    output [7:0] col_out_832,
    output [7:0] col_out_833,
    output [7:0] col_out_834,
    output [7:0] col_out_835,
    output [7:0] col_out_836,
    output [7:0] col_out_837,
    output [7:0] col_out_838,
    output [7:0] col_out_839,
    output [7:0] col_out_840,
    output [7:0] col_out_841,
    output [7:0] col_out_842,
    output [7:0] col_out_843,
    output [7:0] col_out_844,
    output [7:0] col_out_845,
    output [7:0] col_out_846,
    output [7:0] col_out_847,
    output [7:0] col_out_848,
    output [7:0] col_out_849,
    output [7:0] col_out_850,
    output [7:0] col_out_851,
    output [7:0] col_out_852,
    output [7:0] col_out_853,
    output [7:0] col_out_854,
    output [7:0] col_out_855,
    output [7:0] col_out_856,
    output [7:0] col_out_857,
    output [7:0] col_out_858,
    output [7:0] col_out_859,
    output [7:0] col_out_860,
    output [7:0] col_out_861,
    output [7:0] col_out_862,
    output [7:0] col_out_863,
    output [7:0] col_out_864,
    output [7:0] col_out_865,
    output [7:0] col_out_866,
    output [7:0] col_out_867,
    output [7:0] col_out_868,
    output [7:0] col_out_869,
    output [7:0] col_out_870,
    output [7:0] col_out_871,
    output [7:0] col_out_872,
    output [7:0] col_out_873,
    output [7:0] col_out_874,
    output [7:0] col_out_875,
    output [7:0] col_out_876,
    output [7:0] col_out_877,
    output [7:0] col_out_878,
    output [7:0] col_out_879,
    output [7:0] col_out_880,
    output [7:0] col_out_881,
    output [7:0] col_out_882,
    output [7:0] col_out_883,
    output [7:0] col_out_884,
    output [7:0] col_out_885,
    output [7:0] col_out_886,
    output [7:0] col_out_887,
    output [7:0] col_out_888,
    output [7:0] col_out_889,
    output [7:0] col_out_890,
    output [7:0] col_out_891,
    output [7:0] col_out_892,
    output [7:0] col_out_893,
    output [7:0] col_out_894,
    output [7:0] col_out_895,
    output [7:0] col_out_896,
    output [7:0] col_out_897,
    output [7:0] col_out_898,
    output [7:0] col_out_899,
    output [7:0] col_out_900,
    output [7:0] col_out_901,
    output [7:0] col_out_902,
    output [7:0] col_out_903,
    output [7:0] col_out_904,
    output [7:0] col_out_905,
    output [7:0] col_out_906,
    output [7:0] col_out_907,
    output [7:0] col_out_908,
    output [7:0] col_out_909,
    output [7:0] col_out_910,
    output [7:0] col_out_911,
    output [7:0] col_out_912,
    output [7:0] col_out_913,
    output [7:0] col_out_914,
    output [7:0] col_out_915,
    output [7:0] col_out_916,
    output [7:0] col_out_917,
    output [7:0] col_out_918,
    output [7:0] col_out_919,
    output [7:0] col_out_920,
    output [7:0] col_out_921,
    output [7:0] col_out_922,
    output [7:0] col_out_923,
    output [7:0] col_out_924,
    output [7:0] col_out_925,
    output [7:0] col_out_926,
    output [7:0] col_out_927,
    output [7:0] col_out_928,
    output [7:0] col_out_929,
    output [7:0] col_out_930,
    output [7:0] col_out_931,
    output [7:0] col_out_932,
    output [7:0] col_out_933,
    output [7:0] col_out_934,
    output [7:0] col_out_935,
    output [7:0] col_out_936,
    output [7:0] col_out_937,
    output [7:0] col_out_938,
    output [7:0] col_out_939,
    output [7:0] col_out_940,
    output [7:0] col_out_941,
    output [7:0] col_out_942,
    output [7:0] col_out_943,
    output [7:0] col_out_944,
    output [7:0] col_out_945,
    output [7:0] col_out_946,
    output [7:0] col_out_947,
    output [7:0] col_out_948,
    output [7:0] col_out_949,
    output [7:0] col_out_950,
    output [7:0] col_out_951,
    output [7:0] col_out_952,
    output [7:0] col_out_953,
    output [7:0] col_out_954,
    output [7:0] col_out_955,
    output [7:0] col_out_956,
    output [7:0] col_out_957,
    output [7:0] col_out_958,
    output [7:0] col_out_959,
    output [7:0] col_out_960,
    output [7:0] col_out_961,
    output [7:0] col_out_962,
    output [7:0] col_out_963,
    output [7:0] col_out_964,
    output [7:0] col_out_965,
    output [7:0] col_out_966,
    output [7:0] col_out_967,
    output [7:0] col_out_968,
    output [7:0] col_out_969,
    output [7:0] col_out_970,
    output [7:0] col_out_971,
    output [7:0] col_out_972,
    output [7:0] col_out_973,
    output [7:0] col_out_974,
    output [7:0] col_out_975,
    output [7:0] col_out_976,
    output [7:0] col_out_977,
    output [7:0] col_out_978,
    output [7:0] col_out_979,
    output [7:0] col_out_980,
    output [7:0] col_out_981,
    output [7:0] col_out_982,
    output [7:0] col_out_983,
    output [7:0] col_out_984,
    output [7:0] col_out_985,
    output [7:0] col_out_986,
    output [7:0] col_out_987,
    output [7:0] col_out_988,
    output [7:0] col_out_989,
    output [7:0] col_out_990,
    output [7:0] col_out_991,
    output [7:0] col_out_992,
    output [7:0] col_out_993,
    output [7:0] col_out_994,
    output [7:0] col_out_995,
    output [7:0] col_out_996,
    output [7:0] col_out_997,
    output [7:0] col_out_998,
    output [7:0] col_out_999,
    output [7:0] col_out_1000,
    output [7:0] col_out_1001,
    output [7:0] col_out_1002,
    output [7:0] col_out_1003,
    output [7:0] col_out_1004,
    output [7:0] col_out_1005,
    output [7:0] col_out_1006,
    output [7:0] col_out_1007,
    output [7:0] col_out_1008,
    output [7:0] col_out_1009,
    output [7:0] col_out_1010,
    output [7:0] col_out_1011,
    output [7:0] col_out_1012,
    output [7:0] col_out_1013,
    output [7:0] col_out_1014,
    output [7:0] col_out_1015,
    output [7:0] col_out_1016,
    output [7:0] col_out_1017,
    output [7:0] col_out_1018,
    output [7:0] col_out_1019,
    output [7:0] col_out_1020,
    output [7:0] col_out_1021,
    output [7:0] col_out_1022,
    output [7:0] col_out_1023,
    output [7:0] col_out_1024,
    output [7:0] col_out_1025,
    output [7:0] col_out_1026,
    output [7:0] col_out_1027,
    output [7:0] col_out_1028,
    output [7:0] col_out_1029,
    output [7:0] col_out_1030,
    output [7:0] col_out_1031,
    output [7:0] col_out_1032,
    output [7:0] col_out_1033
);



//--compressor_array input and output----------------------

wire [11:0] u_ca_in_0;
wire [11:0] u_ca_in_1;
wire [11:0] u_ca_in_2;
wire [11:0] u_ca_in_3;
wire [11:0] u_ca_in_4;
wire [11:0] u_ca_in_5;
wire [11:0] u_ca_in_6;
wire [11:0] u_ca_in_7;
wire [11:0] u_ca_in_8;
wire [11:0] u_ca_in_9;
wire [11:0] u_ca_in_10;
wire [11:0] u_ca_in_11;
wire [11:0] u_ca_in_12;
wire [11:0] u_ca_in_13;
wire [11:0] u_ca_in_14;
wire [11:0] u_ca_in_15;
wire [11:0] u_ca_in_16;
wire [11:0] u_ca_in_17;
wire [11:0] u_ca_in_18;
wire [11:0] u_ca_in_19;
wire [11:0] u_ca_in_20;
wire [11:0] u_ca_in_21;
wire [11:0] u_ca_in_22;
wire [11:0] u_ca_in_23;
wire [11:0] u_ca_in_24;
wire [11:0] u_ca_in_25;
wire [11:0] u_ca_in_26;
wire [11:0] u_ca_in_27;
wire [11:0] u_ca_in_28;
wire [11:0] u_ca_in_29;
wire [11:0] u_ca_in_30;
wire [11:0] u_ca_in_31;
wire [11:0] u_ca_in_32;
wire [11:0] u_ca_in_33;
wire [11:0] u_ca_in_34;
wire [11:0] u_ca_in_35;
wire [11:0] u_ca_in_36;
wire [11:0] u_ca_in_37;
wire [11:0] u_ca_in_38;
wire [11:0] u_ca_in_39;
wire [11:0] u_ca_in_40;
wire [11:0] u_ca_in_41;
wire [11:0] u_ca_in_42;
wire [11:0] u_ca_in_43;
wire [11:0] u_ca_in_44;
wire [11:0] u_ca_in_45;
wire [11:0] u_ca_in_46;
wire [11:0] u_ca_in_47;
wire [11:0] u_ca_in_48;
wire [11:0] u_ca_in_49;
wire [11:0] u_ca_in_50;
wire [11:0] u_ca_in_51;
wire [11:0] u_ca_in_52;
wire [11:0] u_ca_in_53;
wire [11:0] u_ca_in_54;
wire [11:0] u_ca_in_55;
wire [11:0] u_ca_in_56;
wire [11:0] u_ca_in_57;
wire [11:0] u_ca_in_58;
wire [11:0] u_ca_in_59;
wire [11:0] u_ca_in_60;
wire [11:0] u_ca_in_61;
wire [11:0] u_ca_in_62;
wire [11:0] u_ca_in_63;
wire [11:0] u_ca_in_64;
wire [11:0] u_ca_in_65;
wire [11:0] u_ca_in_66;
wire [11:0] u_ca_in_67;
wire [11:0] u_ca_in_68;
wire [11:0] u_ca_in_69;
wire [11:0] u_ca_in_70;
wire [11:0] u_ca_in_71;
wire [11:0] u_ca_in_72;
wire [11:0] u_ca_in_73;
wire [11:0] u_ca_in_74;
wire [11:0] u_ca_in_75;
wire [11:0] u_ca_in_76;
wire [11:0] u_ca_in_77;
wire [11:0] u_ca_in_78;
wire [11:0] u_ca_in_79;
wire [11:0] u_ca_in_80;
wire [11:0] u_ca_in_81;
wire [11:0] u_ca_in_82;
wire [11:0] u_ca_in_83;
wire [11:0] u_ca_in_84;
wire [11:0] u_ca_in_85;
wire [11:0] u_ca_in_86;
wire [11:0] u_ca_in_87;
wire [11:0] u_ca_in_88;
wire [11:0] u_ca_in_89;
wire [11:0] u_ca_in_90;
wire [11:0] u_ca_in_91;
wire [11:0] u_ca_in_92;
wire [11:0] u_ca_in_93;
wire [11:0] u_ca_in_94;
wire [11:0] u_ca_in_95;
wire [11:0] u_ca_in_96;
wire [11:0] u_ca_in_97;
wire [11:0] u_ca_in_98;
wire [11:0] u_ca_in_99;
wire [11:0] u_ca_in_100;
wire [11:0] u_ca_in_101;
wire [11:0] u_ca_in_102;
wire [11:0] u_ca_in_103;
wire [11:0] u_ca_in_104;
wire [11:0] u_ca_in_105;
wire [11:0] u_ca_in_106;
wire [11:0] u_ca_in_107;
wire [11:0] u_ca_in_108;
wire [11:0] u_ca_in_109;
wire [11:0] u_ca_in_110;
wire [11:0] u_ca_in_111;
wire [11:0] u_ca_in_112;
wire [11:0] u_ca_in_113;
wire [11:0] u_ca_in_114;
wire [11:0] u_ca_in_115;
wire [11:0] u_ca_in_116;
wire [11:0] u_ca_in_117;
wire [11:0] u_ca_in_118;
wire [11:0] u_ca_in_119;
wire [11:0] u_ca_in_120;
wire [11:0] u_ca_in_121;
wire [11:0] u_ca_in_122;
wire [11:0] u_ca_in_123;
wire [11:0] u_ca_in_124;
wire [11:0] u_ca_in_125;
wire [11:0] u_ca_in_126;
wire [11:0] u_ca_in_127;
wire [11:0] u_ca_in_128;
wire [11:0] u_ca_in_129;
wire [11:0] u_ca_in_130;
wire [11:0] u_ca_in_131;
wire [11:0] u_ca_in_132;
wire [11:0] u_ca_in_133;
wire [11:0] u_ca_in_134;
wire [11:0] u_ca_in_135;
wire [11:0] u_ca_in_136;
wire [11:0] u_ca_in_137;
wire [11:0] u_ca_in_138;
wire [11:0] u_ca_in_139;
wire [11:0] u_ca_in_140;
wire [11:0] u_ca_in_141;
wire [11:0] u_ca_in_142;
wire [11:0] u_ca_in_143;
wire [11:0] u_ca_in_144;
wire [11:0] u_ca_in_145;
wire [11:0] u_ca_in_146;
wire [11:0] u_ca_in_147;
wire [11:0] u_ca_in_148;
wire [11:0] u_ca_in_149;
wire [11:0] u_ca_in_150;
wire [11:0] u_ca_in_151;
wire [11:0] u_ca_in_152;
wire [11:0] u_ca_in_153;
wire [11:0] u_ca_in_154;
wire [11:0] u_ca_in_155;
wire [11:0] u_ca_in_156;
wire [11:0] u_ca_in_157;
wire [11:0] u_ca_in_158;
wire [11:0] u_ca_in_159;
wire [11:0] u_ca_in_160;
wire [11:0] u_ca_in_161;
wire [11:0] u_ca_in_162;
wire [11:0] u_ca_in_163;
wire [11:0] u_ca_in_164;
wire [11:0] u_ca_in_165;
wire [11:0] u_ca_in_166;
wire [11:0] u_ca_in_167;
wire [11:0] u_ca_in_168;
wire [11:0] u_ca_in_169;
wire [11:0] u_ca_in_170;
wire [11:0] u_ca_in_171;
wire [11:0] u_ca_in_172;
wire [11:0] u_ca_in_173;
wire [11:0] u_ca_in_174;
wire [11:0] u_ca_in_175;
wire [11:0] u_ca_in_176;
wire [11:0] u_ca_in_177;
wire [11:0] u_ca_in_178;
wire [11:0] u_ca_in_179;
wire [11:0] u_ca_in_180;
wire [11:0] u_ca_in_181;
wire [11:0] u_ca_in_182;
wire [11:0] u_ca_in_183;
wire [11:0] u_ca_in_184;
wire [11:0] u_ca_in_185;
wire [11:0] u_ca_in_186;
wire [11:0] u_ca_in_187;
wire [11:0] u_ca_in_188;
wire [11:0] u_ca_in_189;
wire [11:0] u_ca_in_190;
wire [11:0] u_ca_in_191;
wire [11:0] u_ca_in_192;
wire [11:0] u_ca_in_193;
wire [11:0] u_ca_in_194;
wire [11:0] u_ca_in_195;
wire [11:0] u_ca_in_196;
wire [11:0] u_ca_in_197;
wire [11:0] u_ca_in_198;
wire [11:0] u_ca_in_199;
wire [11:0] u_ca_in_200;
wire [11:0] u_ca_in_201;
wire [11:0] u_ca_in_202;
wire [11:0] u_ca_in_203;
wire [11:0] u_ca_in_204;
wire [11:0] u_ca_in_205;
wire [11:0] u_ca_in_206;
wire [11:0] u_ca_in_207;
wire [11:0] u_ca_in_208;
wire [11:0] u_ca_in_209;
wire [11:0] u_ca_in_210;
wire [11:0] u_ca_in_211;
wire [11:0] u_ca_in_212;
wire [11:0] u_ca_in_213;
wire [11:0] u_ca_in_214;
wire [11:0] u_ca_in_215;
wire [11:0] u_ca_in_216;
wire [11:0] u_ca_in_217;
wire [11:0] u_ca_in_218;
wire [11:0] u_ca_in_219;
wire [11:0] u_ca_in_220;
wire [11:0] u_ca_in_221;
wire [11:0] u_ca_in_222;
wire [11:0] u_ca_in_223;
wire [11:0] u_ca_in_224;
wire [11:0] u_ca_in_225;
wire [11:0] u_ca_in_226;
wire [11:0] u_ca_in_227;
wire [11:0] u_ca_in_228;
wire [11:0] u_ca_in_229;
wire [11:0] u_ca_in_230;
wire [11:0] u_ca_in_231;
wire [11:0] u_ca_in_232;
wire [11:0] u_ca_in_233;
wire [11:0] u_ca_in_234;
wire [11:0] u_ca_in_235;
wire [11:0] u_ca_in_236;
wire [11:0] u_ca_in_237;
wire [11:0] u_ca_in_238;
wire [11:0] u_ca_in_239;
wire [11:0] u_ca_in_240;
wire [11:0] u_ca_in_241;
wire [11:0] u_ca_in_242;
wire [11:0] u_ca_in_243;
wire [11:0] u_ca_in_244;
wire [11:0] u_ca_in_245;
wire [11:0] u_ca_in_246;
wire [11:0] u_ca_in_247;
wire [11:0] u_ca_in_248;
wire [11:0] u_ca_in_249;
wire [11:0] u_ca_in_250;
wire [11:0] u_ca_in_251;
wire [11:0] u_ca_in_252;
wire [11:0] u_ca_in_253;
wire [11:0] u_ca_in_254;
wire [11:0] u_ca_in_255;
wire [11:0] u_ca_in_256;
wire [11:0] u_ca_in_257;
wire [11:0] u_ca_in_258;
wire [11:0] u_ca_in_259;
wire [11:0] u_ca_in_260;
wire [11:0] u_ca_in_261;
wire [11:0] u_ca_in_262;
wire [11:0] u_ca_in_263;
wire [11:0] u_ca_in_264;
wire [11:0] u_ca_in_265;
wire [11:0] u_ca_in_266;
wire [11:0] u_ca_in_267;
wire [11:0] u_ca_in_268;
wire [11:0] u_ca_in_269;
wire [11:0] u_ca_in_270;
wire [11:0] u_ca_in_271;
wire [11:0] u_ca_in_272;
wire [11:0] u_ca_in_273;
wire [11:0] u_ca_in_274;
wire [11:0] u_ca_in_275;
wire [11:0] u_ca_in_276;
wire [11:0] u_ca_in_277;
wire [11:0] u_ca_in_278;
wire [11:0] u_ca_in_279;
wire [11:0] u_ca_in_280;
wire [11:0] u_ca_in_281;
wire [11:0] u_ca_in_282;
wire [11:0] u_ca_in_283;
wire [11:0] u_ca_in_284;
wire [11:0] u_ca_in_285;
wire [11:0] u_ca_in_286;
wire [11:0] u_ca_in_287;
wire [11:0] u_ca_in_288;
wire [11:0] u_ca_in_289;
wire [11:0] u_ca_in_290;
wire [11:0] u_ca_in_291;
wire [11:0] u_ca_in_292;
wire [11:0] u_ca_in_293;
wire [11:0] u_ca_in_294;
wire [11:0] u_ca_in_295;
wire [11:0] u_ca_in_296;
wire [11:0] u_ca_in_297;
wire [11:0] u_ca_in_298;
wire [11:0] u_ca_in_299;
wire [11:0] u_ca_in_300;
wire [11:0] u_ca_in_301;
wire [11:0] u_ca_in_302;
wire [11:0] u_ca_in_303;
wire [11:0] u_ca_in_304;
wire [11:0] u_ca_in_305;
wire [11:0] u_ca_in_306;
wire [11:0] u_ca_in_307;
wire [11:0] u_ca_in_308;
wire [11:0] u_ca_in_309;
wire [11:0] u_ca_in_310;
wire [11:0] u_ca_in_311;
wire [11:0] u_ca_in_312;
wire [11:0] u_ca_in_313;
wire [11:0] u_ca_in_314;
wire [11:0] u_ca_in_315;
wire [11:0] u_ca_in_316;
wire [11:0] u_ca_in_317;
wire [11:0] u_ca_in_318;
wire [11:0] u_ca_in_319;
wire [11:0] u_ca_in_320;
wire [11:0] u_ca_in_321;
wire [11:0] u_ca_in_322;
wire [11:0] u_ca_in_323;
wire [11:0] u_ca_in_324;
wire [11:0] u_ca_in_325;
wire [11:0] u_ca_in_326;
wire [11:0] u_ca_in_327;
wire [11:0] u_ca_in_328;
wire [11:0] u_ca_in_329;
wire [11:0] u_ca_in_330;
wire [11:0] u_ca_in_331;
wire [11:0] u_ca_in_332;
wire [11:0] u_ca_in_333;
wire [11:0] u_ca_in_334;
wire [11:0] u_ca_in_335;
wire [11:0] u_ca_in_336;
wire [11:0] u_ca_in_337;
wire [11:0] u_ca_in_338;
wire [11:0] u_ca_in_339;
wire [11:0] u_ca_in_340;
wire [11:0] u_ca_in_341;
wire [11:0] u_ca_in_342;
wire [11:0] u_ca_in_343;
wire [11:0] u_ca_in_344;
wire [11:0] u_ca_in_345;
wire [11:0] u_ca_in_346;
wire [11:0] u_ca_in_347;
wire [11:0] u_ca_in_348;
wire [11:0] u_ca_in_349;
wire [11:0] u_ca_in_350;
wire [11:0] u_ca_in_351;
wire [11:0] u_ca_in_352;
wire [11:0] u_ca_in_353;
wire [11:0] u_ca_in_354;
wire [11:0] u_ca_in_355;
wire [11:0] u_ca_in_356;
wire [11:0] u_ca_in_357;
wire [11:0] u_ca_in_358;
wire [11:0] u_ca_in_359;
wire [11:0] u_ca_in_360;
wire [11:0] u_ca_in_361;
wire [11:0] u_ca_in_362;
wire [11:0] u_ca_in_363;
wire [11:0] u_ca_in_364;
wire [11:0] u_ca_in_365;
wire [11:0] u_ca_in_366;
wire [11:0] u_ca_in_367;
wire [11:0] u_ca_in_368;
wire [11:0] u_ca_in_369;
wire [11:0] u_ca_in_370;
wire [11:0] u_ca_in_371;
wire [11:0] u_ca_in_372;
wire [11:0] u_ca_in_373;
wire [11:0] u_ca_in_374;
wire [11:0] u_ca_in_375;
wire [11:0] u_ca_in_376;
wire [11:0] u_ca_in_377;
wire [11:0] u_ca_in_378;
wire [11:0] u_ca_in_379;
wire [11:0] u_ca_in_380;
wire [11:0] u_ca_in_381;
wire [11:0] u_ca_in_382;
wire [11:0] u_ca_in_383;
wire [11:0] u_ca_in_384;
wire [11:0] u_ca_in_385;
wire [11:0] u_ca_in_386;
wire [11:0] u_ca_in_387;
wire [11:0] u_ca_in_388;
wire [11:0] u_ca_in_389;
wire [11:0] u_ca_in_390;
wire [11:0] u_ca_in_391;
wire [11:0] u_ca_in_392;
wire [11:0] u_ca_in_393;
wire [11:0] u_ca_in_394;
wire [11:0] u_ca_in_395;
wire [11:0] u_ca_in_396;
wire [11:0] u_ca_in_397;
wire [11:0] u_ca_in_398;
wire [11:0] u_ca_in_399;
wire [11:0] u_ca_in_400;
wire [11:0] u_ca_in_401;
wire [11:0] u_ca_in_402;
wire [11:0] u_ca_in_403;
wire [11:0] u_ca_in_404;
wire [11:0] u_ca_in_405;
wire [11:0] u_ca_in_406;
wire [11:0] u_ca_in_407;
wire [11:0] u_ca_in_408;
wire [11:0] u_ca_in_409;
wire [11:0] u_ca_in_410;
wire [11:0] u_ca_in_411;
wire [11:0] u_ca_in_412;
wire [11:0] u_ca_in_413;
wire [11:0] u_ca_in_414;
wire [11:0] u_ca_in_415;
wire [11:0] u_ca_in_416;
wire [11:0] u_ca_in_417;
wire [11:0] u_ca_in_418;
wire [11:0] u_ca_in_419;
wire [11:0] u_ca_in_420;
wire [11:0] u_ca_in_421;
wire [11:0] u_ca_in_422;
wire [11:0] u_ca_in_423;
wire [11:0] u_ca_in_424;
wire [11:0] u_ca_in_425;
wire [11:0] u_ca_in_426;
wire [11:0] u_ca_in_427;
wire [11:0] u_ca_in_428;
wire [11:0] u_ca_in_429;
wire [11:0] u_ca_in_430;
wire [11:0] u_ca_in_431;
wire [11:0] u_ca_in_432;
wire [11:0] u_ca_in_433;
wire [11:0] u_ca_in_434;
wire [11:0] u_ca_in_435;
wire [11:0] u_ca_in_436;
wire [11:0] u_ca_in_437;
wire [11:0] u_ca_in_438;
wire [11:0] u_ca_in_439;
wire [11:0] u_ca_in_440;
wire [11:0] u_ca_in_441;
wire [11:0] u_ca_in_442;
wire [11:0] u_ca_in_443;
wire [11:0] u_ca_in_444;
wire [11:0] u_ca_in_445;
wire [11:0] u_ca_in_446;
wire [11:0] u_ca_in_447;
wire [11:0] u_ca_in_448;
wire [11:0] u_ca_in_449;
wire [11:0] u_ca_in_450;
wire [11:0] u_ca_in_451;
wire [11:0] u_ca_in_452;
wire [11:0] u_ca_in_453;
wire [11:0] u_ca_in_454;
wire [11:0] u_ca_in_455;
wire [11:0] u_ca_in_456;
wire [11:0] u_ca_in_457;
wire [11:0] u_ca_in_458;
wire [11:0] u_ca_in_459;
wire [11:0] u_ca_in_460;
wire [11:0] u_ca_in_461;
wire [11:0] u_ca_in_462;
wire [11:0] u_ca_in_463;
wire [11:0] u_ca_in_464;
wire [11:0] u_ca_in_465;
wire [11:0] u_ca_in_466;
wire [11:0] u_ca_in_467;
wire [11:0] u_ca_in_468;
wire [11:0] u_ca_in_469;
wire [11:0] u_ca_in_470;
wire [11:0] u_ca_in_471;
wire [11:0] u_ca_in_472;
wire [11:0] u_ca_in_473;
wire [11:0] u_ca_in_474;
wire [11:0] u_ca_in_475;
wire [11:0] u_ca_in_476;
wire [11:0] u_ca_in_477;
wire [11:0] u_ca_in_478;
wire [11:0] u_ca_in_479;
wire [11:0] u_ca_in_480;
wire [11:0] u_ca_in_481;
wire [11:0] u_ca_in_482;
wire [11:0] u_ca_in_483;
wire [11:0] u_ca_in_484;
wire [11:0] u_ca_in_485;
wire [11:0] u_ca_in_486;
wire [11:0] u_ca_in_487;
wire [11:0] u_ca_in_488;
wire [11:0] u_ca_in_489;
wire [11:0] u_ca_in_490;
wire [11:0] u_ca_in_491;
wire [11:0] u_ca_in_492;
wire [11:0] u_ca_in_493;
wire [11:0] u_ca_in_494;
wire [11:0] u_ca_in_495;
wire [11:0] u_ca_in_496;
wire [11:0] u_ca_in_497;
wire [11:0] u_ca_in_498;
wire [11:0] u_ca_in_499;
wire [11:0] u_ca_in_500;
wire [11:0] u_ca_in_501;
wire [11:0] u_ca_in_502;
wire [11:0] u_ca_in_503;
wire [11:0] u_ca_in_504;
wire [11:0] u_ca_in_505;
wire [11:0] u_ca_in_506;
wire [11:0] u_ca_in_507;
wire [11:0] u_ca_in_508;
wire [11:0] u_ca_in_509;
wire [11:0] u_ca_in_510;
wire [11:0] u_ca_in_511;
wire [11:0] u_ca_in_512;
wire [11:0] u_ca_in_513;
wire [11:0] u_ca_in_514;
wire [11:0] u_ca_in_515;
wire [11:0] u_ca_in_516;
wire [11:0] u_ca_in_517;
wire [11:0] u_ca_in_518;
wire [11:0] u_ca_in_519;
wire [11:0] u_ca_in_520;
wire [11:0] u_ca_in_521;
wire [11:0] u_ca_in_522;
wire [11:0] u_ca_in_523;
wire [11:0] u_ca_in_524;
wire [11:0] u_ca_in_525;
wire [11:0] u_ca_in_526;
wire [11:0] u_ca_in_527;
wire [11:0] u_ca_in_528;
wire [11:0] u_ca_in_529;
wire [11:0] u_ca_in_530;
wire [11:0] u_ca_in_531;
wire [11:0] u_ca_in_532;
wire [11:0] u_ca_in_533;
wire [11:0] u_ca_in_534;
wire [11:0] u_ca_in_535;
wire [11:0] u_ca_in_536;
wire [11:0] u_ca_in_537;
wire [11:0] u_ca_in_538;
wire [11:0] u_ca_in_539;
wire [11:0] u_ca_in_540;
wire [11:0] u_ca_in_541;
wire [11:0] u_ca_in_542;
wire [11:0] u_ca_in_543;
wire [11:0] u_ca_in_544;
wire [11:0] u_ca_in_545;
wire [11:0] u_ca_in_546;
wire [11:0] u_ca_in_547;
wire [11:0] u_ca_in_548;
wire [11:0] u_ca_in_549;
wire [11:0] u_ca_in_550;
wire [11:0] u_ca_in_551;
wire [11:0] u_ca_in_552;
wire [11:0] u_ca_in_553;
wire [11:0] u_ca_in_554;
wire [11:0] u_ca_in_555;
wire [11:0] u_ca_in_556;
wire [11:0] u_ca_in_557;
wire [11:0] u_ca_in_558;
wire [11:0] u_ca_in_559;
wire [11:0] u_ca_in_560;
wire [11:0] u_ca_in_561;
wire [11:0] u_ca_in_562;
wire [11:0] u_ca_in_563;
wire [11:0] u_ca_in_564;
wire [11:0] u_ca_in_565;
wire [11:0] u_ca_in_566;
wire [11:0] u_ca_in_567;
wire [11:0] u_ca_in_568;
wire [11:0] u_ca_in_569;
wire [11:0] u_ca_in_570;
wire [11:0] u_ca_in_571;
wire [11:0] u_ca_in_572;
wire [11:0] u_ca_in_573;
wire [11:0] u_ca_in_574;
wire [11:0] u_ca_in_575;
wire [11:0] u_ca_in_576;
wire [11:0] u_ca_in_577;
wire [11:0] u_ca_in_578;
wire [11:0] u_ca_in_579;
wire [11:0] u_ca_in_580;
wire [11:0] u_ca_in_581;
wire [11:0] u_ca_in_582;
wire [11:0] u_ca_in_583;
wire [11:0] u_ca_in_584;
wire [11:0] u_ca_in_585;
wire [11:0] u_ca_in_586;
wire [11:0] u_ca_in_587;
wire [11:0] u_ca_in_588;
wire [11:0] u_ca_in_589;
wire [11:0] u_ca_in_590;
wire [11:0] u_ca_in_591;
wire [11:0] u_ca_in_592;
wire [11:0] u_ca_in_593;
wire [11:0] u_ca_in_594;
wire [11:0] u_ca_in_595;
wire [11:0] u_ca_in_596;
wire [11:0] u_ca_in_597;
wire [11:0] u_ca_in_598;
wire [11:0] u_ca_in_599;
wire [11:0] u_ca_in_600;
wire [11:0] u_ca_in_601;
wire [11:0] u_ca_in_602;
wire [11:0] u_ca_in_603;
wire [11:0] u_ca_in_604;
wire [11:0] u_ca_in_605;
wire [11:0] u_ca_in_606;
wire [11:0] u_ca_in_607;
wire [11:0] u_ca_in_608;
wire [11:0] u_ca_in_609;
wire [11:0] u_ca_in_610;
wire [11:0] u_ca_in_611;
wire [11:0] u_ca_in_612;
wire [11:0] u_ca_in_613;
wire [11:0] u_ca_in_614;
wire [11:0] u_ca_in_615;
wire [11:0] u_ca_in_616;
wire [11:0] u_ca_in_617;
wire [11:0] u_ca_in_618;
wire [11:0] u_ca_in_619;
wire [11:0] u_ca_in_620;
wire [11:0] u_ca_in_621;
wire [11:0] u_ca_in_622;
wire [11:0] u_ca_in_623;
wire [11:0] u_ca_in_624;
wire [11:0] u_ca_in_625;
wire [11:0] u_ca_in_626;
wire [11:0] u_ca_in_627;
wire [11:0] u_ca_in_628;
wire [11:0] u_ca_in_629;
wire [11:0] u_ca_in_630;
wire [11:0] u_ca_in_631;
wire [11:0] u_ca_in_632;
wire [11:0] u_ca_in_633;
wire [11:0] u_ca_in_634;
wire [11:0] u_ca_in_635;
wire [11:0] u_ca_in_636;
wire [11:0] u_ca_in_637;
wire [11:0] u_ca_in_638;
wire [11:0] u_ca_in_639;
wire [11:0] u_ca_in_640;
wire [11:0] u_ca_in_641;
wire [11:0] u_ca_in_642;
wire [11:0] u_ca_in_643;
wire [11:0] u_ca_in_644;
wire [11:0] u_ca_in_645;
wire [11:0] u_ca_in_646;
wire [11:0] u_ca_in_647;
wire [11:0] u_ca_in_648;
wire [11:0] u_ca_in_649;
wire [11:0] u_ca_in_650;
wire [11:0] u_ca_in_651;
wire [11:0] u_ca_in_652;
wire [11:0] u_ca_in_653;
wire [11:0] u_ca_in_654;
wire [11:0] u_ca_in_655;
wire [11:0] u_ca_in_656;
wire [11:0] u_ca_in_657;
wire [11:0] u_ca_in_658;
wire [11:0] u_ca_in_659;
wire [11:0] u_ca_in_660;
wire [11:0] u_ca_in_661;
wire [11:0] u_ca_in_662;
wire [11:0] u_ca_in_663;
wire [11:0] u_ca_in_664;
wire [11:0] u_ca_in_665;
wire [11:0] u_ca_in_666;
wire [11:0] u_ca_in_667;
wire [11:0] u_ca_in_668;
wire [11:0] u_ca_in_669;
wire [11:0] u_ca_in_670;
wire [11:0] u_ca_in_671;
wire [11:0] u_ca_in_672;
wire [11:0] u_ca_in_673;
wire [11:0] u_ca_in_674;
wire [11:0] u_ca_in_675;
wire [11:0] u_ca_in_676;
wire [11:0] u_ca_in_677;
wire [11:0] u_ca_in_678;
wire [11:0] u_ca_in_679;
wire [11:0] u_ca_in_680;
wire [11:0] u_ca_in_681;
wire [11:0] u_ca_in_682;
wire [11:0] u_ca_in_683;
wire [11:0] u_ca_in_684;
wire [11:0] u_ca_in_685;
wire [11:0] u_ca_in_686;
wire [11:0] u_ca_in_687;
wire [11:0] u_ca_in_688;
wire [11:0] u_ca_in_689;
wire [11:0] u_ca_in_690;
wire [11:0] u_ca_in_691;
wire [11:0] u_ca_in_692;
wire [11:0] u_ca_in_693;
wire [11:0] u_ca_in_694;
wire [11:0] u_ca_in_695;
wire [11:0] u_ca_in_696;
wire [11:0] u_ca_in_697;
wire [11:0] u_ca_in_698;
wire [11:0] u_ca_in_699;
wire [11:0] u_ca_in_700;
wire [11:0] u_ca_in_701;
wire [11:0] u_ca_in_702;
wire [11:0] u_ca_in_703;
wire [11:0] u_ca_in_704;
wire [11:0] u_ca_in_705;
wire [11:0] u_ca_in_706;
wire [11:0] u_ca_in_707;
wire [11:0] u_ca_in_708;
wire [11:0] u_ca_in_709;
wire [11:0] u_ca_in_710;
wire [11:0] u_ca_in_711;
wire [11:0] u_ca_in_712;
wire [11:0] u_ca_in_713;
wire [11:0] u_ca_in_714;
wire [11:0] u_ca_in_715;
wire [11:0] u_ca_in_716;
wire [11:0] u_ca_in_717;
wire [11:0] u_ca_in_718;
wire [11:0] u_ca_in_719;
wire [11:0] u_ca_in_720;
wire [11:0] u_ca_in_721;
wire [11:0] u_ca_in_722;
wire [11:0] u_ca_in_723;
wire [11:0] u_ca_in_724;
wire [11:0] u_ca_in_725;
wire [11:0] u_ca_in_726;
wire [11:0] u_ca_in_727;
wire [11:0] u_ca_in_728;
wire [11:0] u_ca_in_729;
wire [11:0] u_ca_in_730;
wire [11:0] u_ca_in_731;
wire [11:0] u_ca_in_732;
wire [11:0] u_ca_in_733;
wire [11:0] u_ca_in_734;
wire [11:0] u_ca_in_735;
wire [11:0] u_ca_in_736;
wire [11:0] u_ca_in_737;
wire [11:0] u_ca_in_738;
wire [11:0] u_ca_in_739;
wire [11:0] u_ca_in_740;
wire [11:0] u_ca_in_741;
wire [11:0] u_ca_in_742;
wire [11:0] u_ca_in_743;
wire [11:0] u_ca_in_744;
wire [11:0] u_ca_in_745;
wire [11:0] u_ca_in_746;
wire [11:0] u_ca_in_747;
wire [11:0] u_ca_in_748;
wire [11:0] u_ca_in_749;
wire [11:0] u_ca_in_750;
wire [11:0] u_ca_in_751;
wire [11:0] u_ca_in_752;
wire [11:0] u_ca_in_753;
wire [11:0] u_ca_in_754;
wire [11:0] u_ca_in_755;
wire [11:0] u_ca_in_756;
wire [11:0] u_ca_in_757;
wire [11:0] u_ca_in_758;
wire [11:0] u_ca_in_759;
wire [11:0] u_ca_in_760;
wire [11:0] u_ca_in_761;
wire [11:0] u_ca_in_762;
wire [11:0] u_ca_in_763;
wire [11:0] u_ca_in_764;
wire [11:0] u_ca_in_765;
wire [11:0] u_ca_in_766;
wire [11:0] u_ca_in_767;
wire [11:0] u_ca_in_768;
wire [11:0] u_ca_in_769;
wire [11:0] u_ca_in_770;
wire [11:0] u_ca_in_771;
wire [11:0] u_ca_in_772;
wire [11:0] u_ca_in_773;
wire [11:0] u_ca_in_774;
wire [11:0] u_ca_in_775;
wire [11:0] u_ca_in_776;
wire [11:0] u_ca_in_777;
wire [11:0] u_ca_in_778;
wire [11:0] u_ca_in_779;
wire [11:0] u_ca_in_780;
wire [11:0] u_ca_in_781;
wire [11:0] u_ca_in_782;
wire [11:0] u_ca_in_783;
wire [11:0] u_ca_in_784;
wire [11:0] u_ca_in_785;
wire [11:0] u_ca_in_786;
wire [11:0] u_ca_in_787;
wire [11:0] u_ca_in_788;
wire [11:0] u_ca_in_789;
wire [11:0] u_ca_in_790;
wire [11:0] u_ca_in_791;
wire [11:0] u_ca_in_792;
wire [11:0] u_ca_in_793;
wire [11:0] u_ca_in_794;
wire [11:0] u_ca_in_795;
wire [11:0] u_ca_in_796;
wire [11:0] u_ca_in_797;
wire [11:0] u_ca_in_798;
wire [11:0] u_ca_in_799;
wire [11:0] u_ca_in_800;
wire [11:0] u_ca_in_801;
wire [11:0] u_ca_in_802;
wire [11:0] u_ca_in_803;
wire [11:0] u_ca_in_804;
wire [11:0] u_ca_in_805;
wire [11:0] u_ca_in_806;
wire [11:0] u_ca_in_807;
wire [11:0] u_ca_in_808;
wire [11:0] u_ca_in_809;
wire [11:0] u_ca_in_810;
wire [11:0] u_ca_in_811;
wire [11:0] u_ca_in_812;
wire [11:0] u_ca_in_813;
wire [11:0] u_ca_in_814;
wire [11:0] u_ca_in_815;
wire [11:0] u_ca_in_816;
wire [11:0] u_ca_in_817;
wire [11:0] u_ca_in_818;
wire [11:0] u_ca_in_819;
wire [11:0] u_ca_in_820;
wire [11:0] u_ca_in_821;
wire [11:0] u_ca_in_822;
wire [11:0] u_ca_in_823;
wire [11:0] u_ca_in_824;
wire [11:0] u_ca_in_825;
wire [11:0] u_ca_in_826;
wire [11:0] u_ca_in_827;
wire [11:0] u_ca_in_828;
wire [11:0] u_ca_in_829;
wire [11:0] u_ca_in_830;
wire [11:0] u_ca_in_831;
wire [11:0] u_ca_in_832;
wire [11:0] u_ca_in_833;
wire [11:0] u_ca_in_834;
wire [11:0] u_ca_in_835;
wire [11:0] u_ca_in_836;
wire [11:0] u_ca_in_837;
wire [11:0] u_ca_in_838;
wire [11:0] u_ca_in_839;
wire [11:0] u_ca_in_840;
wire [11:0] u_ca_in_841;
wire [11:0] u_ca_in_842;
wire [11:0] u_ca_in_843;
wire [11:0] u_ca_in_844;
wire [11:0] u_ca_in_845;
wire [11:0] u_ca_in_846;
wire [11:0] u_ca_in_847;
wire [11:0] u_ca_in_848;
wire [11:0] u_ca_in_849;
wire [11:0] u_ca_in_850;
wire [11:0] u_ca_in_851;
wire [11:0] u_ca_in_852;
wire [11:0] u_ca_in_853;
wire [11:0] u_ca_in_854;
wire [11:0] u_ca_in_855;
wire [11:0] u_ca_in_856;
wire [11:0] u_ca_in_857;
wire [11:0] u_ca_in_858;
wire [11:0] u_ca_in_859;
wire [11:0] u_ca_in_860;
wire [11:0] u_ca_in_861;
wire [11:0] u_ca_in_862;
wire [11:0] u_ca_in_863;
wire [11:0] u_ca_in_864;
wire [11:0] u_ca_in_865;
wire [11:0] u_ca_in_866;
wire [11:0] u_ca_in_867;
wire [11:0] u_ca_in_868;
wire [11:0] u_ca_in_869;
wire [11:0] u_ca_in_870;
wire [11:0] u_ca_in_871;
wire [11:0] u_ca_in_872;
wire [11:0] u_ca_in_873;
wire [11:0] u_ca_in_874;
wire [11:0] u_ca_in_875;
wire [11:0] u_ca_in_876;
wire [11:0] u_ca_in_877;
wire [11:0] u_ca_in_878;
wire [11:0] u_ca_in_879;
wire [11:0] u_ca_in_880;
wire [11:0] u_ca_in_881;
wire [11:0] u_ca_in_882;
wire [11:0] u_ca_in_883;
wire [11:0] u_ca_in_884;
wire [11:0] u_ca_in_885;
wire [11:0] u_ca_in_886;
wire [11:0] u_ca_in_887;
wire [11:0] u_ca_in_888;
wire [11:0] u_ca_in_889;
wire [11:0] u_ca_in_890;
wire [11:0] u_ca_in_891;
wire [11:0] u_ca_in_892;
wire [11:0] u_ca_in_893;
wire [11:0] u_ca_in_894;
wire [11:0] u_ca_in_895;
wire [11:0] u_ca_in_896;
wire [11:0] u_ca_in_897;
wire [11:0] u_ca_in_898;
wire [11:0] u_ca_in_899;
wire [11:0] u_ca_in_900;
wire [11:0] u_ca_in_901;
wire [11:0] u_ca_in_902;
wire [11:0] u_ca_in_903;
wire [11:0] u_ca_in_904;
wire [11:0] u_ca_in_905;
wire [11:0] u_ca_in_906;
wire [11:0] u_ca_in_907;
wire [11:0] u_ca_in_908;
wire [11:0] u_ca_in_909;
wire [11:0] u_ca_in_910;
wire [11:0] u_ca_in_911;
wire [11:0] u_ca_in_912;
wire [11:0] u_ca_in_913;
wire [11:0] u_ca_in_914;
wire [11:0] u_ca_in_915;
wire [11:0] u_ca_in_916;
wire [11:0] u_ca_in_917;
wire [11:0] u_ca_in_918;
wire [11:0] u_ca_in_919;
wire [11:0] u_ca_in_920;
wire [11:0] u_ca_in_921;
wire [11:0] u_ca_in_922;
wire [11:0] u_ca_in_923;
wire [11:0] u_ca_in_924;
wire [11:0] u_ca_in_925;
wire [11:0] u_ca_in_926;
wire [11:0] u_ca_in_927;
wire [11:0] u_ca_in_928;
wire [11:0] u_ca_in_929;
wire [11:0] u_ca_in_930;
wire [11:0] u_ca_in_931;
wire [11:0] u_ca_in_932;
wire [11:0] u_ca_in_933;
wire [11:0] u_ca_in_934;
wire [11:0] u_ca_in_935;
wire [11:0] u_ca_in_936;
wire [11:0] u_ca_in_937;
wire [11:0] u_ca_in_938;
wire [11:0] u_ca_in_939;
wire [11:0] u_ca_in_940;
wire [11:0] u_ca_in_941;
wire [11:0] u_ca_in_942;
wire [11:0] u_ca_in_943;
wire [11:0] u_ca_in_944;
wire [11:0] u_ca_in_945;
wire [11:0] u_ca_in_946;
wire [11:0] u_ca_in_947;
wire [11:0] u_ca_in_948;
wire [11:0] u_ca_in_949;
wire [11:0] u_ca_in_950;
wire [11:0] u_ca_in_951;
wire [11:0] u_ca_in_952;
wire [11:0] u_ca_in_953;
wire [11:0] u_ca_in_954;
wire [11:0] u_ca_in_955;
wire [11:0] u_ca_in_956;
wire [11:0] u_ca_in_957;
wire [11:0] u_ca_in_958;
wire [11:0] u_ca_in_959;
wire [11:0] u_ca_in_960;
wire [11:0] u_ca_in_961;
wire [11:0] u_ca_in_962;
wire [11:0] u_ca_in_963;
wire [11:0] u_ca_in_964;
wire [11:0] u_ca_in_965;
wire [11:0] u_ca_in_966;
wire [11:0] u_ca_in_967;
wire [11:0] u_ca_in_968;
wire [11:0] u_ca_in_969;
wire [11:0] u_ca_in_970;
wire [11:0] u_ca_in_971;
wire [11:0] u_ca_in_972;
wire [11:0] u_ca_in_973;
wire [11:0] u_ca_in_974;
wire [11:0] u_ca_in_975;
wire [11:0] u_ca_in_976;
wire [11:0] u_ca_in_977;
wire [11:0] u_ca_in_978;
wire [11:0] u_ca_in_979;
wire [11:0] u_ca_in_980;
wire [11:0] u_ca_in_981;
wire [11:0] u_ca_in_982;
wire [11:0] u_ca_in_983;
wire [11:0] u_ca_in_984;
wire [11:0] u_ca_in_985;
wire [11:0] u_ca_in_986;
wire [11:0] u_ca_in_987;
wire [11:0] u_ca_in_988;
wire [11:0] u_ca_in_989;
wire [11:0] u_ca_in_990;
wire [11:0] u_ca_in_991;
wire [11:0] u_ca_in_992;
wire [11:0] u_ca_in_993;
wire [11:0] u_ca_in_994;
wire [11:0] u_ca_in_995;
wire [11:0] u_ca_in_996;
wire [11:0] u_ca_in_997;
wire [11:0] u_ca_in_998;
wire [11:0] u_ca_in_999;
wire [11:0] u_ca_in_1000;
wire [11:0] u_ca_in_1001;
wire [11:0] u_ca_in_1002;
wire [11:0] u_ca_in_1003;
wire [11:0] u_ca_in_1004;
wire [11:0] u_ca_in_1005;
wire [11:0] u_ca_in_1006;
wire [11:0] u_ca_in_1007;
wire [11:0] u_ca_in_1008;
wire [11:0] u_ca_in_1009;
wire [11:0] u_ca_in_1010;
wire [11:0] u_ca_in_1011;
wire [11:0] u_ca_in_1012;
wire [11:0] u_ca_in_1013;
wire [11:0] u_ca_in_1014;
wire [11:0] u_ca_in_1015;
wire [11:0] u_ca_in_1016;
wire [11:0] u_ca_in_1017;
wire [11:0] u_ca_in_1018;
wire [11:0] u_ca_in_1019;
wire [11:0] u_ca_in_1020;
wire [11:0] u_ca_in_1021;
wire [11:0] u_ca_in_1022;
wire [11:0] u_ca_in_1023;
wire [11:0] u_ca_in_1024;
wire [11:0] u_ca_in_1025;
wire [11:0] u_ca_in_1026;
wire [11:0] u_ca_in_1027;
wire [11:0] u_ca_in_1028;
wire [11:0] u_ca_in_1029;
wire [11:0] u_ca_in_1030;
wire [11:0] u_ca_in_1031;
wire [11:0] u_ca_in_1032;

wire [7:0] u_ca_out_0;
wire [7:0] u_ca_out_1;
wire [7:0] u_ca_out_2;
wire [7:0] u_ca_out_3;
wire [7:0] u_ca_out_4;
wire [7:0] u_ca_out_5;
wire [7:0] u_ca_out_6;
wire [7:0] u_ca_out_7;
wire [7:0] u_ca_out_8;
wire [7:0] u_ca_out_9;
wire [7:0] u_ca_out_10;
wire [7:0] u_ca_out_11;
wire [7:0] u_ca_out_12;
wire [7:0] u_ca_out_13;
wire [7:0] u_ca_out_14;
wire [7:0] u_ca_out_15;
wire [7:0] u_ca_out_16;
wire [7:0] u_ca_out_17;
wire [7:0] u_ca_out_18;
wire [7:0] u_ca_out_19;
wire [7:0] u_ca_out_20;
wire [7:0] u_ca_out_21;
wire [7:0] u_ca_out_22;
wire [7:0] u_ca_out_23;
wire [7:0] u_ca_out_24;
wire [7:0] u_ca_out_25;
wire [7:0] u_ca_out_26;
wire [7:0] u_ca_out_27;
wire [7:0] u_ca_out_28;
wire [7:0] u_ca_out_29;
wire [7:0] u_ca_out_30;
wire [7:0] u_ca_out_31;
wire [7:0] u_ca_out_32;
wire [7:0] u_ca_out_33;
wire [7:0] u_ca_out_34;
wire [7:0] u_ca_out_35;
wire [7:0] u_ca_out_36;
wire [7:0] u_ca_out_37;
wire [7:0] u_ca_out_38;
wire [7:0] u_ca_out_39;
wire [7:0] u_ca_out_40;
wire [7:0] u_ca_out_41;
wire [7:0] u_ca_out_42;
wire [7:0] u_ca_out_43;
wire [7:0] u_ca_out_44;
wire [7:0] u_ca_out_45;
wire [7:0] u_ca_out_46;
wire [7:0] u_ca_out_47;
wire [7:0] u_ca_out_48;
wire [7:0] u_ca_out_49;
wire [7:0] u_ca_out_50;
wire [7:0] u_ca_out_51;
wire [7:0] u_ca_out_52;
wire [7:0] u_ca_out_53;
wire [7:0] u_ca_out_54;
wire [7:0] u_ca_out_55;
wire [7:0] u_ca_out_56;
wire [7:0] u_ca_out_57;
wire [7:0] u_ca_out_58;
wire [7:0] u_ca_out_59;
wire [7:0] u_ca_out_60;
wire [7:0] u_ca_out_61;
wire [7:0] u_ca_out_62;
wire [7:0] u_ca_out_63;
wire [7:0] u_ca_out_64;
wire [7:0] u_ca_out_65;
wire [7:0] u_ca_out_66;
wire [7:0] u_ca_out_67;
wire [7:0] u_ca_out_68;
wire [7:0] u_ca_out_69;
wire [7:0] u_ca_out_70;
wire [7:0] u_ca_out_71;
wire [7:0] u_ca_out_72;
wire [7:0] u_ca_out_73;
wire [7:0] u_ca_out_74;
wire [7:0] u_ca_out_75;
wire [7:0] u_ca_out_76;
wire [7:0] u_ca_out_77;
wire [7:0] u_ca_out_78;
wire [7:0] u_ca_out_79;
wire [7:0] u_ca_out_80;
wire [7:0] u_ca_out_81;
wire [7:0] u_ca_out_82;
wire [7:0] u_ca_out_83;
wire [7:0] u_ca_out_84;
wire [7:0] u_ca_out_85;
wire [7:0] u_ca_out_86;
wire [7:0] u_ca_out_87;
wire [7:0] u_ca_out_88;
wire [7:0] u_ca_out_89;
wire [7:0] u_ca_out_90;
wire [7:0] u_ca_out_91;
wire [7:0] u_ca_out_92;
wire [7:0] u_ca_out_93;
wire [7:0] u_ca_out_94;
wire [7:0] u_ca_out_95;
wire [7:0] u_ca_out_96;
wire [7:0] u_ca_out_97;
wire [7:0] u_ca_out_98;
wire [7:0] u_ca_out_99;
wire [7:0] u_ca_out_100;
wire [7:0] u_ca_out_101;
wire [7:0] u_ca_out_102;
wire [7:0] u_ca_out_103;
wire [7:0] u_ca_out_104;
wire [7:0] u_ca_out_105;
wire [7:0] u_ca_out_106;
wire [7:0] u_ca_out_107;
wire [7:0] u_ca_out_108;
wire [7:0] u_ca_out_109;
wire [7:0] u_ca_out_110;
wire [7:0] u_ca_out_111;
wire [7:0] u_ca_out_112;
wire [7:0] u_ca_out_113;
wire [7:0] u_ca_out_114;
wire [7:0] u_ca_out_115;
wire [7:0] u_ca_out_116;
wire [7:0] u_ca_out_117;
wire [7:0] u_ca_out_118;
wire [7:0] u_ca_out_119;
wire [7:0] u_ca_out_120;
wire [7:0] u_ca_out_121;
wire [7:0] u_ca_out_122;
wire [7:0] u_ca_out_123;
wire [7:0] u_ca_out_124;
wire [7:0] u_ca_out_125;
wire [7:0] u_ca_out_126;
wire [7:0] u_ca_out_127;
wire [7:0] u_ca_out_128;
wire [7:0] u_ca_out_129;
wire [7:0] u_ca_out_130;
wire [7:0] u_ca_out_131;
wire [7:0] u_ca_out_132;
wire [7:0] u_ca_out_133;
wire [7:0] u_ca_out_134;
wire [7:0] u_ca_out_135;
wire [7:0] u_ca_out_136;
wire [7:0] u_ca_out_137;
wire [7:0] u_ca_out_138;
wire [7:0] u_ca_out_139;
wire [7:0] u_ca_out_140;
wire [7:0] u_ca_out_141;
wire [7:0] u_ca_out_142;
wire [7:0] u_ca_out_143;
wire [7:0] u_ca_out_144;
wire [7:0] u_ca_out_145;
wire [7:0] u_ca_out_146;
wire [7:0] u_ca_out_147;
wire [7:0] u_ca_out_148;
wire [7:0] u_ca_out_149;
wire [7:0] u_ca_out_150;
wire [7:0] u_ca_out_151;
wire [7:0] u_ca_out_152;
wire [7:0] u_ca_out_153;
wire [7:0] u_ca_out_154;
wire [7:0] u_ca_out_155;
wire [7:0] u_ca_out_156;
wire [7:0] u_ca_out_157;
wire [7:0] u_ca_out_158;
wire [7:0] u_ca_out_159;
wire [7:0] u_ca_out_160;
wire [7:0] u_ca_out_161;
wire [7:0] u_ca_out_162;
wire [7:0] u_ca_out_163;
wire [7:0] u_ca_out_164;
wire [7:0] u_ca_out_165;
wire [7:0] u_ca_out_166;
wire [7:0] u_ca_out_167;
wire [7:0] u_ca_out_168;
wire [7:0] u_ca_out_169;
wire [7:0] u_ca_out_170;
wire [7:0] u_ca_out_171;
wire [7:0] u_ca_out_172;
wire [7:0] u_ca_out_173;
wire [7:0] u_ca_out_174;
wire [7:0] u_ca_out_175;
wire [7:0] u_ca_out_176;
wire [7:0] u_ca_out_177;
wire [7:0] u_ca_out_178;
wire [7:0] u_ca_out_179;
wire [7:0] u_ca_out_180;
wire [7:0] u_ca_out_181;
wire [7:0] u_ca_out_182;
wire [7:0] u_ca_out_183;
wire [7:0] u_ca_out_184;
wire [7:0] u_ca_out_185;
wire [7:0] u_ca_out_186;
wire [7:0] u_ca_out_187;
wire [7:0] u_ca_out_188;
wire [7:0] u_ca_out_189;
wire [7:0] u_ca_out_190;
wire [7:0] u_ca_out_191;
wire [7:0] u_ca_out_192;
wire [7:0] u_ca_out_193;
wire [7:0] u_ca_out_194;
wire [7:0] u_ca_out_195;
wire [7:0] u_ca_out_196;
wire [7:0] u_ca_out_197;
wire [7:0] u_ca_out_198;
wire [7:0] u_ca_out_199;
wire [7:0] u_ca_out_200;
wire [7:0] u_ca_out_201;
wire [7:0] u_ca_out_202;
wire [7:0] u_ca_out_203;
wire [7:0] u_ca_out_204;
wire [7:0] u_ca_out_205;
wire [7:0] u_ca_out_206;
wire [7:0] u_ca_out_207;
wire [7:0] u_ca_out_208;
wire [7:0] u_ca_out_209;
wire [7:0] u_ca_out_210;
wire [7:0] u_ca_out_211;
wire [7:0] u_ca_out_212;
wire [7:0] u_ca_out_213;
wire [7:0] u_ca_out_214;
wire [7:0] u_ca_out_215;
wire [7:0] u_ca_out_216;
wire [7:0] u_ca_out_217;
wire [7:0] u_ca_out_218;
wire [7:0] u_ca_out_219;
wire [7:0] u_ca_out_220;
wire [7:0] u_ca_out_221;
wire [7:0] u_ca_out_222;
wire [7:0] u_ca_out_223;
wire [7:0] u_ca_out_224;
wire [7:0] u_ca_out_225;
wire [7:0] u_ca_out_226;
wire [7:0] u_ca_out_227;
wire [7:0] u_ca_out_228;
wire [7:0] u_ca_out_229;
wire [7:0] u_ca_out_230;
wire [7:0] u_ca_out_231;
wire [7:0] u_ca_out_232;
wire [7:0] u_ca_out_233;
wire [7:0] u_ca_out_234;
wire [7:0] u_ca_out_235;
wire [7:0] u_ca_out_236;
wire [7:0] u_ca_out_237;
wire [7:0] u_ca_out_238;
wire [7:0] u_ca_out_239;
wire [7:0] u_ca_out_240;
wire [7:0] u_ca_out_241;
wire [7:0] u_ca_out_242;
wire [7:0] u_ca_out_243;
wire [7:0] u_ca_out_244;
wire [7:0] u_ca_out_245;
wire [7:0] u_ca_out_246;
wire [7:0] u_ca_out_247;
wire [7:0] u_ca_out_248;
wire [7:0] u_ca_out_249;
wire [7:0] u_ca_out_250;
wire [7:0] u_ca_out_251;
wire [7:0] u_ca_out_252;
wire [7:0] u_ca_out_253;
wire [7:0] u_ca_out_254;
wire [7:0] u_ca_out_255;
wire [7:0] u_ca_out_256;
wire [7:0] u_ca_out_257;
wire [7:0] u_ca_out_258;
wire [7:0] u_ca_out_259;
wire [7:0] u_ca_out_260;
wire [7:0] u_ca_out_261;
wire [7:0] u_ca_out_262;
wire [7:0] u_ca_out_263;
wire [7:0] u_ca_out_264;
wire [7:0] u_ca_out_265;
wire [7:0] u_ca_out_266;
wire [7:0] u_ca_out_267;
wire [7:0] u_ca_out_268;
wire [7:0] u_ca_out_269;
wire [7:0] u_ca_out_270;
wire [7:0] u_ca_out_271;
wire [7:0] u_ca_out_272;
wire [7:0] u_ca_out_273;
wire [7:0] u_ca_out_274;
wire [7:0] u_ca_out_275;
wire [7:0] u_ca_out_276;
wire [7:0] u_ca_out_277;
wire [7:0] u_ca_out_278;
wire [7:0] u_ca_out_279;
wire [7:0] u_ca_out_280;
wire [7:0] u_ca_out_281;
wire [7:0] u_ca_out_282;
wire [7:0] u_ca_out_283;
wire [7:0] u_ca_out_284;
wire [7:0] u_ca_out_285;
wire [7:0] u_ca_out_286;
wire [7:0] u_ca_out_287;
wire [7:0] u_ca_out_288;
wire [7:0] u_ca_out_289;
wire [7:0] u_ca_out_290;
wire [7:0] u_ca_out_291;
wire [7:0] u_ca_out_292;
wire [7:0] u_ca_out_293;
wire [7:0] u_ca_out_294;
wire [7:0] u_ca_out_295;
wire [7:0] u_ca_out_296;
wire [7:0] u_ca_out_297;
wire [7:0] u_ca_out_298;
wire [7:0] u_ca_out_299;
wire [7:0] u_ca_out_300;
wire [7:0] u_ca_out_301;
wire [7:0] u_ca_out_302;
wire [7:0] u_ca_out_303;
wire [7:0] u_ca_out_304;
wire [7:0] u_ca_out_305;
wire [7:0] u_ca_out_306;
wire [7:0] u_ca_out_307;
wire [7:0] u_ca_out_308;
wire [7:0] u_ca_out_309;
wire [7:0] u_ca_out_310;
wire [7:0] u_ca_out_311;
wire [7:0] u_ca_out_312;
wire [7:0] u_ca_out_313;
wire [7:0] u_ca_out_314;
wire [7:0] u_ca_out_315;
wire [7:0] u_ca_out_316;
wire [7:0] u_ca_out_317;
wire [7:0] u_ca_out_318;
wire [7:0] u_ca_out_319;
wire [7:0] u_ca_out_320;
wire [7:0] u_ca_out_321;
wire [7:0] u_ca_out_322;
wire [7:0] u_ca_out_323;
wire [7:0] u_ca_out_324;
wire [7:0] u_ca_out_325;
wire [7:0] u_ca_out_326;
wire [7:0] u_ca_out_327;
wire [7:0] u_ca_out_328;
wire [7:0] u_ca_out_329;
wire [7:0] u_ca_out_330;
wire [7:0] u_ca_out_331;
wire [7:0] u_ca_out_332;
wire [7:0] u_ca_out_333;
wire [7:0] u_ca_out_334;
wire [7:0] u_ca_out_335;
wire [7:0] u_ca_out_336;
wire [7:0] u_ca_out_337;
wire [7:0] u_ca_out_338;
wire [7:0] u_ca_out_339;
wire [7:0] u_ca_out_340;
wire [7:0] u_ca_out_341;
wire [7:0] u_ca_out_342;
wire [7:0] u_ca_out_343;
wire [7:0] u_ca_out_344;
wire [7:0] u_ca_out_345;
wire [7:0] u_ca_out_346;
wire [7:0] u_ca_out_347;
wire [7:0] u_ca_out_348;
wire [7:0] u_ca_out_349;
wire [7:0] u_ca_out_350;
wire [7:0] u_ca_out_351;
wire [7:0] u_ca_out_352;
wire [7:0] u_ca_out_353;
wire [7:0] u_ca_out_354;
wire [7:0] u_ca_out_355;
wire [7:0] u_ca_out_356;
wire [7:0] u_ca_out_357;
wire [7:0] u_ca_out_358;
wire [7:0] u_ca_out_359;
wire [7:0] u_ca_out_360;
wire [7:0] u_ca_out_361;
wire [7:0] u_ca_out_362;
wire [7:0] u_ca_out_363;
wire [7:0] u_ca_out_364;
wire [7:0] u_ca_out_365;
wire [7:0] u_ca_out_366;
wire [7:0] u_ca_out_367;
wire [7:0] u_ca_out_368;
wire [7:0] u_ca_out_369;
wire [7:0] u_ca_out_370;
wire [7:0] u_ca_out_371;
wire [7:0] u_ca_out_372;
wire [7:0] u_ca_out_373;
wire [7:0] u_ca_out_374;
wire [7:0] u_ca_out_375;
wire [7:0] u_ca_out_376;
wire [7:0] u_ca_out_377;
wire [7:0] u_ca_out_378;
wire [7:0] u_ca_out_379;
wire [7:0] u_ca_out_380;
wire [7:0] u_ca_out_381;
wire [7:0] u_ca_out_382;
wire [7:0] u_ca_out_383;
wire [7:0] u_ca_out_384;
wire [7:0] u_ca_out_385;
wire [7:0] u_ca_out_386;
wire [7:0] u_ca_out_387;
wire [7:0] u_ca_out_388;
wire [7:0] u_ca_out_389;
wire [7:0] u_ca_out_390;
wire [7:0] u_ca_out_391;
wire [7:0] u_ca_out_392;
wire [7:0] u_ca_out_393;
wire [7:0] u_ca_out_394;
wire [7:0] u_ca_out_395;
wire [7:0] u_ca_out_396;
wire [7:0] u_ca_out_397;
wire [7:0] u_ca_out_398;
wire [7:0] u_ca_out_399;
wire [7:0] u_ca_out_400;
wire [7:0] u_ca_out_401;
wire [7:0] u_ca_out_402;
wire [7:0] u_ca_out_403;
wire [7:0] u_ca_out_404;
wire [7:0] u_ca_out_405;
wire [7:0] u_ca_out_406;
wire [7:0] u_ca_out_407;
wire [7:0] u_ca_out_408;
wire [7:0] u_ca_out_409;
wire [7:0] u_ca_out_410;
wire [7:0] u_ca_out_411;
wire [7:0] u_ca_out_412;
wire [7:0] u_ca_out_413;
wire [7:0] u_ca_out_414;
wire [7:0] u_ca_out_415;
wire [7:0] u_ca_out_416;
wire [7:0] u_ca_out_417;
wire [7:0] u_ca_out_418;
wire [7:0] u_ca_out_419;
wire [7:0] u_ca_out_420;
wire [7:0] u_ca_out_421;
wire [7:0] u_ca_out_422;
wire [7:0] u_ca_out_423;
wire [7:0] u_ca_out_424;
wire [7:0] u_ca_out_425;
wire [7:0] u_ca_out_426;
wire [7:0] u_ca_out_427;
wire [7:0] u_ca_out_428;
wire [7:0] u_ca_out_429;
wire [7:0] u_ca_out_430;
wire [7:0] u_ca_out_431;
wire [7:0] u_ca_out_432;
wire [7:0] u_ca_out_433;
wire [7:0] u_ca_out_434;
wire [7:0] u_ca_out_435;
wire [7:0] u_ca_out_436;
wire [7:0] u_ca_out_437;
wire [7:0] u_ca_out_438;
wire [7:0] u_ca_out_439;
wire [7:0] u_ca_out_440;
wire [7:0] u_ca_out_441;
wire [7:0] u_ca_out_442;
wire [7:0] u_ca_out_443;
wire [7:0] u_ca_out_444;
wire [7:0] u_ca_out_445;
wire [7:0] u_ca_out_446;
wire [7:0] u_ca_out_447;
wire [7:0] u_ca_out_448;
wire [7:0] u_ca_out_449;
wire [7:0] u_ca_out_450;
wire [7:0] u_ca_out_451;
wire [7:0] u_ca_out_452;
wire [7:0] u_ca_out_453;
wire [7:0] u_ca_out_454;
wire [7:0] u_ca_out_455;
wire [7:0] u_ca_out_456;
wire [7:0] u_ca_out_457;
wire [7:0] u_ca_out_458;
wire [7:0] u_ca_out_459;
wire [7:0] u_ca_out_460;
wire [7:0] u_ca_out_461;
wire [7:0] u_ca_out_462;
wire [7:0] u_ca_out_463;
wire [7:0] u_ca_out_464;
wire [7:0] u_ca_out_465;
wire [7:0] u_ca_out_466;
wire [7:0] u_ca_out_467;
wire [7:0] u_ca_out_468;
wire [7:0] u_ca_out_469;
wire [7:0] u_ca_out_470;
wire [7:0] u_ca_out_471;
wire [7:0] u_ca_out_472;
wire [7:0] u_ca_out_473;
wire [7:0] u_ca_out_474;
wire [7:0] u_ca_out_475;
wire [7:0] u_ca_out_476;
wire [7:0] u_ca_out_477;
wire [7:0] u_ca_out_478;
wire [7:0] u_ca_out_479;
wire [7:0] u_ca_out_480;
wire [7:0] u_ca_out_481;
wire [7:0] u_ca_out_482;
wire [7:0] u_ca_out_483;
wire [7:0] u_ca_out_484;
wire [7:0] u_ca_out_485;
wire [7:0] u_ca_out_486;
wire [7:0] u_ca_out_487;
wire [7:0] u_ca_out_488;
wire [7:0] u_ca_out_489;
wire [7:0] u_ca_out_490;
wire [7:0] u_ca_out_491;
wire [7:0] u_ca_out_492;
wire [7:0] u_ca_out_493;
wire [7:0] u_ca_out_494;
wire [7:0] u_ca_out_495;
wire [7:0] u_ca_out_496;
wire [7:0] u_ca_out_497;
wire [7:0] u_ca_out_498;
wire [7:0] u_ca_out_499;
wire [7:0] u_ca_out_500;
wire [7:0] u_ca_out_501;
wire [7:0] u_ca_out_502;
wire [7:0] u_ca_out_503;
wire [7:0] u_ca_out_504;
wire [7:0] u_ca_out_505;
wire [7:0] u_ca_out_506;
wire [7:0] u_ca_out_507;
wire [7:0] u_ca_out_508;
wire [7:0] u_ca_out_509;
wire [7:0] u_ca_out_510;
wire [7:0] u_ca_out_511;
wire [7:0] u_ca_out_512;
wire [7:0] u_ca_out_513;
wire [7:0] u_ca_out_514;
wire [7:0] u_ca_out_515;
wire [7:0] u_ca_out_516;
wire [7:0] u_ca_out_517;
wire [7:0] u_ca_out_518;
wire [7:0] u_ca_out_519;
wire [7:0] u_ca_out_520;
wire [7:0] u_ca_out_521;
wire [7:0] u_ca_out_522;
wire [7:0] u_ca_out_523;
wire [7:0] u_ca_out_524;
wire [7:0] u_ca_out_525;
wire [7:0] u_ca_out_526;
wire [7:0] u_ca_out_527;
wire [7:0] u_ca_out_528;
wire [7:0] u_ca_out_529;
wire [7:0] u_ca_out_530;
wire [7:0] u_ca_out_531;
wire [7:0] u_ca_out_532;
wire [7:0] u_ca_out_533;
wire [7:0] u_ca_out_534;
wire [7:0] u_ca_out_535;
wire [7:0] u_ca_out_536;
wire [7:0] u_ca_out_537;
wire [7:0] u_ca_out_538;
wire [7:0] u_ca_out_539;
wire [7:0] u_ca_out_540;
wire [7:0] u_ca_out_541;
wire [7:0] u_ca_out_542;
wire [7:0] u_ca_out_543;
wire [7:0] u_ca_out_544;
wire [7:0] u_ca_out_545;
wire [7:0] u_ca_out_546;
wire [7:0] u_ca_out_547;
wire [7:0] u_ca_out_548;
wire [7:0] u_ca_out_549;
wire [7:0] u_ca_out_550;
wire [7:0] u_ca_out_551;
wire [7:0] u_ca_out_552;
wire [7:0] u_ca_out_553;
wire [7:0] u_ca_out_554;
wire [7:0] u_ca_out_555;
wire [7:0] u_ca_out_556;
wire [7:0] u_ca_out_557;
wire [7:0] u_ca_out_558;
wire [7:0] u_ca_out_559;
wire [7:0] u_ca_out_560;
wire [7:0] u_ca_out_561;
wire [7:0] u_ca_out_562;
wire [7:0] u_ca_out_563;
wire [7:0] u_ca_out_564;
wire [7:0] u_ca_out_565;
wire [7:0] u_ca_out_566;
wire [7:0] u_ca_out_567;
wire [7:0] u_ca_out_568;
wire [7:0] u_ca_out_569;
wire [7:0] u_ca_out_570;
wire [7:0] u_ca_out_571;
wire [7:0] u_ca_out_572;
wire [7:0] u_ca_out_573;
wire [7:0] u_ca_out_574;
wire [7:0] u_ca_out_575;
wire [7:0] u_ca_out_576;
wire [7:0] u_ca_out_577;
wire [7:0] u_ca_out_578;
wire [7:0] u_ca_out_579;
wire [7:0] u_ca_out_580;
wire [7:0] u_ca_out_581;
wire [7:0] u_ca_out_582;
wire [7:0] u_ca_out_583;
wire [7:0] u_ca_out_584;
wire [7:0] u_ca_out_585;
wire [7:0] u_ca_out_586;
wire [7:0] u_ca_out_587;
wire [7:0] u_ca_out_588;
wire [7:0] u_ca_out_589;
wire [7:0] u_ca_out_590;
wire [7:0] u_ca_out_591;
wire [7:0] u_ca_out_592;
wire [7:0] u_ca_out_593;
wire [7:0] u_ca_out_594;
wire [7:0] u_ca_out_595;
wire [7:0] u_ca_out_596;
wire [7:0] u_ca_out_597;
wire [7:0] u_ca_out_598;
wire [7:0] u_ca_out_599;
wire [7:0] u_ca_out_600;
wire [7:0] u_ca_out_601;
wire [7:0] u_ca_out_602;
wire [7:0] u_ca_out_603;
wire [7:0] u_ca_out_604;
wire [7:0] u_ca_out_605;
wire [7:0] u_ca_out_606;
wire [7:0] u_ca_out_607;
wire [7:0] u_ca_out_608;
wire [7:0] u_ca_out_609;
wire [7:0] u_ca_out_610;
wire [7:0] u_ca_out_611;
wire [7:0] u_ca_out_612;
wire [7:0] u_ca_out_613;
wire [7:0] u_ca_out_614;
wire [7:0] u_ca_out_615;
wire [7:0] u_ca_out_616;
wire [7:0] u_ca_out_617;
wire [7:0] u_ca_out_618;
wire [7:0] u_ca_out_619;
wire [7:0] u_ca_out_620;
wire [7:0] u_ca_out_621;
wire [7:0] u_ca_out_622;
wire [7:0] u_ca_out_623;
wire [7:0] u_ca_out_624;
wire [7:0] u_ca_out_625;
wire [7:0] u_ca_out_626;
wire [7:0] u_ca_out_627;
wire [7:0] u_ca_out_628;
wire [7:0] u_ca_out_629;
wire [7:0] u_ca_out_630;
wire [7:0] u_ca_out_631;
wire [7:0] u_ca_out_632;
wire [7:0] u_ca_out_633;
wire [7:0] u_ca_out_634;
wire [7:0] u_ca_out_635;
wire [7:0] u_ca_out_636;
wire [7:0] u_ca_out_637;
wire [7:0] u_ca_out_638;
wire [7:0] u_ca_out_639;
wire [7:0] u_ca_out_640;
wire [7:0] u_ca_out_641;
wire [7:0] u_ca_out_642;
wire [7:0] u_ca_out_643;
wire [7:0] u_ca_out_644;
wire [7:0] u_ca_out_645;
wire [7:0] u_ca_out_646;
wire [7:0] u_ca_out_647;
wire [7:0] u_ca_out_648;
wire [7:0] u_ca_out_649;
wire [7:0] u_ca_out_650;
wire [7:0] u_ca_out_651;
wire [7:0] u_ca_out_652;
wire [7:0] u_ca_out_653;
wire [7:0] u_ca_out_654;
wire [7:0] u_ca_out_655;
wire [7:0] u_ca_out_656;
wire [7:0] u_ca_out_657;
wire [7:0] u_ca_out_658;
wire [7:0] u_ca_out_659;
wire [7:0] u_ca_out_660;
wire [7:0] u_ca_out_661;
wire [7:0] u_ca_out_662;
wire [7:0] u_ca_out_663;
wire [7:0] u_ca_out_664;
wire [7:0] u_ca_out_665;
wire [7:0] u_ca_out_666;
wire [7:0] u_ca_out_667;
wire [7:0] u_ca_out_668;
wire [7:0] u_ca_out_669;
wire [7:0] u_ca_out_670;
wire [7:0] u_ca_out_671;
wire [7:0] u_ca_out_672;
wire [7:0] u_ca_out_673;
wire [7:0] u_ca_out_674;
wire [7:0] u_ca_out_675;
wire [7:0] u_ca_out_676;
wire [7:0] u_ca_out_677;
wire [7:0] u_ca_out_678;
wire [7:0] u_ca_out_679;
wire [7:0] u_ca_out_680;
wire [7:0] u_ca_out_681;
wire [7:0] u_ca_out_682;
wire [7:0] u_ca_out_683;
wire [7:0] u_ca_out_684;
wire [7:0] u_ca_out_685;
wire [7:0] u_ca_out_686;
wire [7:0] u_ca_out_687;
wire [7:0] u_ca_out_688;
wire [7:0] u_ca_out_689;
wire [7:0] u_ca_out_690;
wire [7:0] u_ca_out_691;
wire [7:0] u_ca_out_692;
wire [7:0] u_ca_out_693;
wire [7:0] u_ca_out_694;
wire [7:0] u_ca_out_695;
wire [7:0] u_ca_out_696;
wire [7:0] u_ca_out_697;
wire [7:0] u_ca_out_698;
wire [7:0] u_ca_out_699;
wire [7:0] u_ca_out_700;
wire [7:0] u_ca_out_701;
wire [7:0] u_ca_out_702;
wire [7:0] u_ca_out_703;
wire [7:0] u_ca_out_704;
wire [7:0] u_ca_out_705;
wire [7:0] u_ca_out_706;
wire [7:0] u_ca_out_707;
wire [7:0] u_ca_out_708;
wire [7:0] u_ca_out_709;
wire [7:0] u_ca_out_710;
wire [7:0] u_ca_out_711;
wire [7:0] u_ca_out_712;
wire [7:0] u_ca_out_713;
wire [7:0] u_ca_out_714;
wire [7:0] u_ca_out_715;
wire [7:0] u_ca_out_716;
wire [7:0] u_ca_out_717;
wire [7:0] u_ca_out_718;
wire [7:0] u_ca_out_719;
wire [7:0] u_ca_out_720;
wire [7:0] u_ca_out_721;
wire [7:0] u_ca_out_722;
wire [7:0] u_ca_out_723;
wire [7:0] u_ca_out_724;
wire [7:0] u_ca_out_725;
wire [7:0] u_ca_out_726;
wire [7:0] u_ca_out_727;
wire [7:0] u_ca_out_728;
wire [7:0] u_ca_out_729;
wire [7:0] u_ca_out_730;
wire [7:0] u_ca_out_731;
wire [7:0] u_ca_out_732;
wire [7:0] u_ca_out_733;
wire [7:0] u_ca_out_734;
wire [7:0] u_ca_out_735;
wire [7:0] u_ca_out_736;
wire [7:0] u_ca_out_737;
wire [7:0] u_ca_out_738;
wire [7:0] u_ca_out_739;
wire [7:0] u_ca_out_740;
wire [7:0] u_ca_out_741;
wire [7:0] u_ca_out_742;
wire [7:0] u_ca_out_743;
wire [7:0] u_ca_out_744;
wire [7:0] u_ca_out_745;
wire [7:0] u_ca_out_746;
wire [7:0] u_ca_out_747;
wire [7:0] u_ca_out_748;
wire [7:0] u_ca_out_749;
wire [7:0] u_ca_out_750;
wire [7:0] u_ca_out_751;
wire [7:0] u_ca_out_752;
wire [7:0] u_ca_out_753;
wire [7:0] u_ca_out_754;
wire [7:0] u_ca_out_755;
wire [7:0] u_ca_out_756;
wire [7:0] u_ca_out_757;
wire [7:0] u_ca_out_758;
wire [7:0] u_ca_out_759;
wire [7:0] u_ca_out_760;
wire [7:0] u_ca_out_761;
wire [7:0] u_ca_out_762;
wire [7:0] u_ca_out_763;
wire [7:0] u_ca_out_764;
wire [7:0] u_ca_out_765;
wire [7:0] u_ca_out_766;
wire [7:0] u_ca_out_767;
wire [7:0] u_ca_out_768;
wire [7:0] u_ca_out_769;
wire [7:0] u_ca_out_770;
wire [7:0] u_ca_out_771;
wire [7:0] u_ca_out_772;
wire [7:0] u_ca_out_773;
wire [7:0] u_ca_out_774;
wire [7:0] u_ca_out_775;
wire [7:0] u_ca_out_776;
wire [7:0] u_ca_out_777;
wire [7:0] u_ca_out_778;
wire [7:0] u_ca_out_779;
wire [7:0] u_ca_out_780;
wire [7:0] u_ca_out_781;
wire [7:0] u_ca_out_782;
wire [7:0] u_ca_out_783;
wire [7:0] u_ca_out_784;
wire [7:0] u_ca_out_785;
wire [7:0] u_ca_out_786;
wire [7:0] u_ca_out_787;
wire [7:0] u_ca_out_788;
wire [7:0] u_ca_out_789;
wire [7:0] u_ca_out_790;
wire [7:0] u_ca_out_791;
wire [7:0] u_ca_out_792;
wire [7:0] u_ca_out_793;
wire [7:0] u_ca_out_794;
wire [7:0] u_ca_out_795;
wire [7:0] u_ca_out_796;
wire [7:0] u_ca_out_797;
wire [7:0] u_ca_out_798;
wire [7:0] u_ca_out_799;
wire [7:0] u_ca_out_800;
wire [7:0] u_ca_out_801;
wire [7:0] u_ca_out_802;
wire [7:0] u_ca_out_803;
wire [7:0] u_ca_out_804;
wire [7:0] u_ca_out_805;
wire [7:0] u_ca_out_806;
wire [7:0] u_ca_out_807;
wire [7:0] u_ca_out_808;
wire [7:0] u_ca_out_809;
wire [7:0] u_ca_out_810;
wire [7:0] u_ca_out_811;
wire [7:0] u_ca_out_812;
wire [7:0] u_ca_out_813;
wire [7:0] u_ca_out_814;
wire [7:0] u_ca_out_815;
wire [7:0] u_ca_out_816;
wire [7:0] u_ca_out_817;
wire [7:0] u_ca_out_818;
wire [7:0] u_ca_out_819;
wire [7:0] u_ca_out_820;
wire [7:0] u_ca_out_821;
wire [7:0] u_ca_out_822;
wire [7:0] u_ca_out_823;
wire [7:0] u_ca_out_824;
wire [7:0] u_ca_out_825;
wire [7:0] u_ca_out_826;
wire [7:0] u_ca_out_827;
wire [7:0] u_ca_out_828;
wire [7:0] u_ca_out_829;
wire [7:0] u_ca_out_830;
wire [7:0] u_ca_out_831;
wire [7:0] u_ca_out_832;
wire [7:0] u_ca_out_833;
wire [7:0] u_ca_out_834;
wire [7:0] u_ca_out_835;
wire [7:0] u_ca_out_836;
wire [7:0] u_ca_out_837;
wire [7:0] u_ca_out_838;
wire [7:0] u_ca_out_839;
wire [7:0] u_ca_out_840;
wire [7:0] u_ca_out_841;
wire [7:0] u_ca_out_842;
wire [7:0] u_ca_out_843;
wire [7:0] u_ca_out_844;
wire [7:0] u_ca_out_845;
wire [7:0] u_ca_out_846;
wire [7:0] u_ca_out_847;
wire [7:0] u_ca_out_848;
wire [7:0] u_ca_out_849;
wire [7:0] u_ca_out_850;
wire [7:0] u_ca_out_851;
wire [7:0] u_ca_out_852;
wire [7:0] u_ca_out_853;
wire [7:0] u_ca_out_854;
wire [7:0] u_ca_out_855;
wire [7:0] u_ca_out_856;
wire [7:0] u_ca_out_857;
wire [7:0] u_ca_out_858;
wire [7:0] u_ca_out_859;
wire [7:0] u_ca_out_860;
wire [7:0] u_ca_out_861;
wire [7:0] u_ca_out_862;
wire [7:0] u_ca_out_863;
wire [7:0] u_ca_out_864;
wire [7:0] u_ca_out_865;
wire [7:0] u_ca_out_866;
wire [7:0] u_ca_out_867;
wire [7:0] u_ca_out_868;
wire [7:0] u_ca_out_869;
wire [7:0] u_ca_out_870;
wire [7:0] u_ca_out_871;
wire [7:0] u_ca_out_872;
wire [7:0] u_ca_out_873;
wire [7:0] u_ca_out_874;
wire [7:0] u_ca_out_875;
wire [7:0] u_ca_out_876;
wire [7:0] u_ca_out_877;
wire [7:0] u_ca_out_878;
wire [7:0] u_ca_out_879;
wire [7:0] u_ca_out_880;
wire [7:0] u_ca_out_881;
wire [7:0] u_ca_out_882;
wire [7:0] u_ca_out_883;
wire [7:0] u_ca_out_884;
wire [7:0] u_ca_out_885;
wire [7:0] u_ca_out_886;
wire [7:0] u_ca_out_887;
wire [7:0] u_ca_out_888;
wire [7:0] u_ca_out_889;
wire [7:0] u_ca_out_890;
wire [7:0] u_ca_out_891;
wire [7:0] u_ca_out_892;
wire [7:0] u_ca_out_893;
wire [7:0] u_ca_out_894;
wire [7:0] u_ca_out_895;
wire [7:0] u_ca_out_896;
wire [7:0] u_ca_out_897;
wire [7:0] u_ca_out_898;
wire [7:0] u_ca_out_899;
wire [7:0] u_ca_out_900;
wire [7:0] u_ca_out_901;
wire [7:0] u_ca_out_902;
wire [7:0] u_ca_out_903;
wire [7:0] u_ca_out_904;
wire [7:0] u_ca_out_905;
wire [7:0] u_ca_out_906;
wire [7:0] u_ca_out_907;
wire [7:0] u_ca_out_908;
wire [7:0] u_ca_out_909;
wire [7:0] u_ca_out_910;
wire [7:0] u_ca_out_911;
wire [7:0] u_ca_out_912;
wire [7:0] u_ca_out_913;
wire [7:0] u_ca_out_914;
wire [7:0] u_ca_out_915;
wire [7:0] u_ca_out_916;
wire [7:0] u_ca_out_917;
wire [7:0] u_ca_out_918;
wire [7:0] u_ca_out_919;
wire [7:0] u_ca_out_920;
wire [7:0] u_ca_out_921;
wire [7:0] u_ca_out_922;
wire [7:0] u_ca_out_923;
wire [7:0] u_ca_out_924;
wire [7:0] u_ca_out_925;
wire [7:0] u_ca_out_926;
wire [7:0] u_ca_out_927;
wire [7:0] u_ca_out_928;
wire [7:0] u_ca_out_929;
wire [7:0] u_ca_out_930;
wire [7:0] u_ca_out_931;
wire [7:0] u_ca_out_932;
wire [7:0] u_ca_out_933;
wire [7:0] u_ca_out_934;
wire [7:0] u_ca_out_935;
wire [7:0] u_ca_out_936;
wire [7:0] u_ca_out_937;
wire [7:0] u_ca_out_938;
wire [7:0] u_ca_out_939;
wire [7:0] u_ca_out_940;
wire [7:0] u_ca_out_941;
wire [7:0] u_ca_out_942;
wire [7:0] u_ca_out_943;
wire [7:0] u_ca_out_944;
wire [7:0] u_ca_out_945;
wire [7:0] u_ca_out_946;
wire [7:0] u_ca_out_947;
wire [7:0] u_ca_out_948;
wire [7:0] u_ca_out_949;
wire [7:0] u_ca_out_950;
wire [7:0] u_ca_out_951;
wire [7:0] u_ca_out_952;
wire [7:0] u_ca_out_953;
wire [7:0] u_ca_out_954;
wire [7:0] u_ca_out_955;
wire [7:0] u_ca_out_956;
wire [7:0] u_ca_out_957;
wire [7:0] u_ca_out_958;
wire [7:0] u_ca_out_959;
wire [7:0] u_ca_out_960;
wire [7:0] u_ca_out_961;
wire [7:0] u_ca_out_962;
wire [7:0] u_ca_out_963;
wire [7:0] u_ca_out_964;
wire [7:0] u_ca_out_965;
wire [7:0] u_ca_out_966;
wire [7:0] u_ca_out_967;
wire [7:0] u_ca_out_968;
wire [7:0] u_ca_out_969;
wire [7:0] u_ca_out_970;
wire [7:0] u_ca_out_971;
wire [7:0] u_ca_out_972;
wire [7:0] u_ca_out_973;
wire [7:0] u_ca_out_974;
wire [7:0] u_ca_out_975;
wire [7:0] u_ca_out_976;
wire [7:0] u_ca_out_977;
wire [7:0] u_ca_out_978;
wire [7:0] u_ca_out_979;
wire [7:0] u_ca_out_980;
wire [7:0] u_ca_out_981;
wire [7:0] u_ca_out_982;
wire [7:0] u_ca_out_983;
wire [7:0] u_ca_out_984;
wire [7:0] u_ca_out_985;
wire [7:0] u_ca_out_986;
wire [7:0] u_ca_out_987;
wire [7:0] u_ca_out_988;
wire [7:0] u_ca_out_989;
wire [7:0] u_ca_out_990;
wire [7:0] u_ca_out_991;
wire [7:0] u_ca_out_992;
wire [7:0] u_ca_out_993;
wire [7:0] u_ca_out_994;
wire [7:0] u_ca_out_995;
wire [7:0] u_ca_out_996;
wire [7:0] u_ca_out_997;
wire [7:0] u_ca_out_998;
wire [7:0] u_ca_out_999;
wire [7:0] u_ca_out_1000;
wire [7:0] u_ca_out_1001;
wire [7:0] u_ca_out_1002;
wire [7:0] u_ca_out_1003;
wire [7:0] u_ca_out_1004;
wire [7:0] u_ca_out_1005;
wire [7:0] u_ca_out_1006;
wire [7:0] u_ca_out_1007;
wire [7:0] u_ca_out_1008;
wire [7:0] u_ca_out_1009;
wire [7:0] u_ca_out_1010;
wire [7:0] u_ca_out_1011;
wire [7:0] u_ca_out_1012;
wire [7:0] u_ca_out_1013;
wire [7:0] u_ca_out_1014;
wire [7:0] u_ca_out_1015;
wire [7:0] u_ca_out_1016;
wire [7:0] u_ca_out_1017;
wire [7:0] u_ca_out_1018;
wire [7:0] u_ca_out_1019;
wire [7:0] u_ca_out_1020;
wire [7:0] u_ca_out_1021;
wire [7:0] u_ca_out_1022;
wire [7:0] u_ca_out_1023;
wire [7:0] u_ca_out_1024;
wire [7:0] u_ca_out_1025;
wire [7:0] u_ca_out_1026;
wire [7:0] u_ca_out_1027;
wire [7:0] u_ca_out_1028;
wire [7:0] u_ca_out_1029;
wire [7:0] u_ca_out_1030;
wire [7:0] u_ca_out_1031;
wire [7:0] u_ca_out_1032;
wire [7:0] u_ca_out_1033;

assign u_ca_in_0 = col_in_0;
assign u_ca_in_1 = col_in_1;
assign u_ca_in_2 = col_in_2;
assign u_ca_in_3 = col_in_3;
assign u_ca_in_4 = col_in_4;
assign u_ca_in_5 = col_in_5;
assign u_ca_in_6 = col_in_6;
assign u_ca_in_7 = col_in_7;
assign u_ca_in_8 = col_in_8;
assign u_ca_in_9 = col_in_9;
assign u_ca_in_10 = col_in_10;
assign u_ca_in_11 = col_in_11;
assign u_ca_in_12 = col_in_12;
assign u_ca_in_13 = col_in_13;
assign u_ca_in_14 = col_in_14;
assign u_ca_in_15 = col_in_15;
assign u_ca_in_16 = col_in_16;
assign u_ca_in_17 = col_in_17;
assign u_ca_in_18 = col_in_18;
assign u_ca_in_19 = col_in_19;
assign u_ca_in_20 = col_in_20;
assign u_ca_in_21 = col_in_21;
assign u_ca_in_22 = col_in_22;
assign u_ca_in_23 = col_in_23;
assign u_ca_in_24 = col_in_24;
assign u_ca_in_25 = col_in_25;
assign u_ca_in_26 = col_in_26;
assign u_ca_in_27 = col_in_27;
assign u_ca_in_28 = col_in_28;
assign u_ca_in_29 = col_in_29;
assign u_ca_in_30 = col_in_30;
assign u_ca_in_31 = col_in_31;
assign u_ca_in_32 = col_in_32;
assign u_ca_in_33 = col_in_33;
assign u_ca_in_34 = col_in_34;
assign u_ca_in_35 = col_in_35;
assign u_ca_in_36 = col_in_36;
assign u_ca_in_37 = col_in_37;
assign u_ca_in_38 = col_in_38;
assign u_ca_in_39 = col_in_39;
assign u_ca_in_40 = col_in_40;
assign u_ca_in_41 = col_in_41;
assign u_ca_in_42 = col_in_42;
assign u_ca_in_43 = col_in_43;
assign u_ca_in_44 = col_in_44;
assign u_ca_in_45 = col_in_45;
assign u_ca_in_46 = col_in_46;
assign u_ca_in_47 = col_in_47;
assign u_ca_in_48 = col_in_48;
assign u_ca_in_49 = col_in_49;
assign u_ca_in_50 = col_in_50;
assign u_ca_in_51 = col_in_51;
assign u_ca_in_52 = col_in_52;
assign u_ca_in_53 = col_in_53;
assign u_ca_in_54 = col_in_54;
assign u_ca_in_55 = col_in_55;
assign u_ca_in_56 = col_in_56;
assign u_ca_in_57 = col_in_57;
assign u_ca_in_58 = col_in_58;
assign u_ca_in_59 = col_in_59;
assign u_ca_in_60 = col_in_60;
assign u_ca_in_61 = col_in_61;
assign u_ca_in_62 = col_in_62;
assign u_ca_in_63 = col_in_63;
assign u_ca_in_64 = col_in_64;
assign u_ca_in_65 = col_in_65;
assign u_ca_in_66 = col_in_66;
assign u_ca_in_67 = col_in_67;
assign u_ca_in_68 = col_in_68;
assign u_ca_in_69 = col_in_69;
assign u_ca_in_70 = col_in_70;
assign u_ca_in_71 = col_in_71;
assign u_ca_in_72 = col_in_72;
assign u_ca_in_73 = col_in_73;
assign u_ca_in_74 = col_in_74;
assign u_ca_in_75 = col_in_75;
assign u_ca_in_76 = col_in_76;
assign u_ca_in_77 = col_in_77;
assign u_ca_in_78 = col_in_78;
assign u_ca_in_79 = col_in_79;
assign u_ca_in_80 = col_in_80;
assign u_ca_in_81 = col_in_81;
assign u_ca_in_82 = col_in_82;
assign u_ca_in_83 = col_in_83;
assign u_ca_in_84 = col_in_84;
assign u_ca_in_85 = col_in_85;
assign u_ca_in_86 = col_in_86;
assign u_ca_in_87 = col_in_87;
assign u_ca_in_88 = col_in_88;
assign u_ca_in_89 = col_in_89;
assign u_ca_in_90 = col_in_90;
assign u_ca_in_91 = col_in_91;
assign u_ca_in_92 = col_in_92;
assign u_ca_in_93 = col_in_93;
assign u_ca_in_94 = col_in_94;
assign u_ca_in_95 = col_in_95;
assign u_ca_in_96 = col_in_96;
assign u_ca_in_97 = col_in_97;
assign u_ca_in_98 = col_in_98;
assign u_ca_in_99 = col_in_99;
assign u_ca_in_100 = col_in_100;
assign u_ca_in_101 = col_in_101;
assign u_ca_in_102 = col_in_102;
assign u_ca_in_103 = col_in_103;
assign u_ca_in_104 = col_in_104;
assign u_ca_in_105 = col_in_105;
assign u_ca_in_106 = col_in_106;
assign u_ca_in_107 = col_in_107;
assign u_ca_in_108 = col_in_108;
assign u_ca_in_109 = col_in_109;
assign u_ca_in_110 = col_in_110;
assign u_ca_in_111 = col_in_111;
assign u_ca_in_112 = col_in_112;
assign u_ca_in_113 = col_in_113;
assign u_ca_in_114 = col_in_114;
assign u_ca_in_115 = col_in_115;
assign u_ca_in_116 = col_in_116;
assign u_ca_in_117 = col_in_117;
assign u_ca_in_118 = col_in_118;
assign u_ca_in_119 = col_in_119;
assign u_ca_in_120 = col_in_120;
assign u_ca_in_121 = col_in_121;
assign u_ca_in_122 = col_in_122;
assign u_ca_in_123 = col_in_123;
assign u_ca_in_124 = col_in_124;
assign u_ca_in_125 = col_in_125;
assign u_ca_in_126 = col_in_126;
assign u_ca_in_127 = col_in_127;
assign u_ca_in_128 = col_in_128;
assign u_ca_in_129 = col_in_129;
assign u_ca_in_130 = col_in_130;
assign u_ca_in_131 = col_in_131;
assign u_ca_in_132 = col_in_132;
assign u_ca_in_133 = col_in_133;
assign u_ca_in_134 = col_in_134;
assign u_ca_in_135 = col_in_135;
assign u_ca_in_136 = col_in_136;
assign u_ca_in_137 = col_in_137;
assign u_ca_in_138 = col_in_138;
assign u_ca_in_139 = col_in_139;
assign u_ca_in_140 = col_in_140;
assign u_ca_in_141 = col_in_141;
assign u_ca_in_142 = col_in_142;
assign u_ca_in_143 = col_in_143;
assign u_ca_in_144 = col_in_144;
assign u_ca_in_145 = col_in_145;
assign u_ca_in_146 = col_in_146;
assign u_ca_in_147 = col_in_147;
assign u_ca_in_148 = col_in_148;
assign u_ca_in_149 = col_in_149;
assign u_ca_in_150 = col_in_150;
assign u_ca_in_151 = col_in_151;
assign u_ca_in_152 = col_in_152;
assign u_ca_in_153 = col_in_153;
assign u_ca_in_154 = col_in_154;
assign u_ca_in_155 = col_in_155;
assign u_ca_in_156 = col_in_156;
assign u_ca_in_157 = col_in_157;
assign u_ca_in_158 = col_in_158;
assign u_ca_in_159 = col_in_159;
assign u_ca_in_160 = col_in_160;
assign u_ca_in_161 = col_in_161;
assign u_ca_in_162 = col_in_162;
assign u_ca_in_163 = col_in_163;
assign u_ca_in_164 = col_in_164;
assign u_ca_in_165 = col_in_165;
assign u_ca_in_166 = col_in_166;
assign u_ca_in_167 = col_in_167;
assign u_ca_in_168 = col_in_168;
assign u_ca_in_169 = col_in_169;
assign u_ca_in_170 = col_in_170;
assign u_ca_in_171 = col_in_171;
assign u_ca_in_172 = col_in_172;
assign u_ca_in_173 = col_in_173;
assign u_ca_in_174 = col_in_174;
assign u_ca_in_175 = col_in_175;
assign u_ca_in_176 = col_in_176;
assign u_ca_in_177 = col_in_177;
assign u_ca_in_178 = col_in_178;
assign u_ca_in_179 = col_in_179;
assign u_ca_in_180 = col_in_180;
assign u_ca_in_181 = col_in_181;
assign u_ca_in_182 = col_in_182;
assign u_ca_in_183 = col_in_183;
assign u_ca_in_184 = col_in_184;
assign u_ca_in_185 = col_in_185;
assign u_ca_in_186 = col_in_186;
assign u_ca_in_187 = col_in_187;
assign u_ca_in_188 = col_in_188;
assign u_ca_in_189 = col_in_189;
assign u_ca_in_190 = col_in_190;
assign u_ca_in_191 = col_in_191;
assign u_ca_in_192 = col_in_192;
assign u_ca_in_193 = col_in_193;
assign u_ca_in_194 = col_in_194;
assign u_ca_in_195 = col_in_195;
assign u_ca_in_196 = col_in_196;
assign u_ca_in_197 = col_in_197;
assign u_ca_in_198 = col_in_198;
assign u_ca_in_199 = col_in_199;
assign u_ca_in_200 = col_in_200;
assign u_ca_in_201 = col_in_201;
assign u_ca_in_202 = col_in_202;
assign u_ca_in_203 = col_in_203;
assign u_ca_in_204 = col_in_204;
assign u_ca_in_205 = col_in_205;
assign u_ca_in_206 = col_in_206;
assign u_ca_in_207 = col_in_207;
assign u_ca_in_208 = col_in_208;
assign u_ca_in_209 = col_in_209;
assign u_ca_in_210 = col_in_210;
assign u_ca_in_211 = col_in_211;
assign u_ca_in_212 = col_in_212;
assign u_ca_in_213 = col_in_213;
assign u_ca_in_214 = col_in_214;
assign u_ca_in_215 = col_in_215;
assign u_ca_in_216 = col_in_216;
assign u_ca_in_217 = col_in_217;
assign u_ca_in_218 = col_in_218;
assign u_ca_in_219 = col_in_219;
assign u_ca_in_220 = col_in_220;
assign u_ca_in_221 = col_in_221;
assign u_ca_in_222 = col_in_222;
assign u_ca_in_223 = col_in_223;
assign u_ca_in_224 = col_in_224;
assign u_ca_in_225 = col_in_225;
assign u_ca_in_226 = col_in_226;
assign u_ca_in_227 = col_in_227;
assign u_ca_in_228 = col_in_228;
assign u_ca_in_229 = col_in_229;
assign u_ca_in_230 = col_in_230;
assign u_ca_in_231 = col_in_231;
assign u_ca_in_232 = col_in_232;
assign u_ca_in_233 = col_in_233;
assign u_ca_in_234 = col_in_234;
assign u_ca_in_235 = col_in_235;
assign u_ca_in_236 = col_in_236;
assign u_ca_in_237 = col_in_237;
assign u_ca_in_238 = col_in_238;
assign u_ca_in_239 = col_in_239;
assign u_ca_in_240 = col_in_240;
assign u_ca_in_241 = col_in_241;
assign u_ca_in_242 = col_in_242;
assign u_ca_in_243 = col_in_243;
assign u_ca_in_244 = col_in_244;
assign u_ca_in_245 = col_in_245;
assign u_ca_in_246 = col_in_246;
assign u_ca_in_247 = col_in_247;
assign u_ca_in_248 = col_in_248;
assign u_ca_in_249 = col_in_249;
assign u_ca_in_250 = col_in_250;
assign u_ca_in_251 = col_in_251;
assign u_ca_in_252 = col_in_252;
assign u_ca_in_253 = col_in_253;
assign u_ca_in_254 = col_in_254;
assign u_ca_in_255 = col_in_255;
assign u_ca_in_256 = col_in_256;
assign u_ca_in_257 = col_in_257;
assign u_ca_in_258 = col_in_258;
assign u_ca_in_259 = col_in_259;
assign u_ca_in_260 = col_in_260;
assign u_ca_in_261 = col_in_261;
assign u_ca_in_262 = col_in_262;
assign u_ca_in_263 = col_in_263;
assign u_ca_in_264 = col_in_264;
assign u_ca_in_265 = col_in_265;
assign u_ca_in_266 = col_in_266;
assign u_ca_in_267 = col_in_267;
assign u_ca_in_268 = col_in_268;
assign u_ca_in_269 = col_in_269;
assign u_ca_in_270 = col_in_270;
assign u_ca_in_271 = col_in_271;
assign u_ca_in_272 = col_in_272;
assign u_ca_in_273 = col_in_273;
assign u_ca_in_274 = col_in_274;
assign u_ca_in_275 = col_in_275;
assign u_ca_in_276 = col_in_276;
assign u_ca_in_277 = col_in_277;
assign u_ca_in_278 = col_in_278;
assign u_ca_in_279 = col_in_279;
assign u_ca_in_280 = col_in_280;
assign u_ca_in_281 = col_in_281;
assign u_ca_in_282 = col_in_282;
assign u_ca_in_283 = col_in_283;
assign u_ca_in_284 = col_in_284;
assign u_ca_in_285 = col_in_285;
assign u_ca_in_286 = col_in_286;
assign u_ca_in_287 = col_in_287;
assign u_ca_in_288 = col_in_288;
assign u_ca_in_289 = col_in_289;
assign u_ca_in_290 = col_in_290;
assign u_ca_in_291 = col_in_291;
assign u_ca_in_292 = col_in_292;
assign u_ca_in_293 = col_in_293;
assign u_ca_in_294 = col_in_294;
assign u_ca_in_295 = col_in_295;
assign u_ca_in_296 = col_in_296;
assign u_ca_in_297 = col_in_297;
assign u_ca_in_298 = col_in_298;
assign u_ca_in_299 = col_in_299;
assign u_ca_in_300 = col_in_300;
assign u_ca_in_301 = col_in_301;
assign u_ca_in_302 = col_in_302;
assign u_ca_in_303 = col_in_303;
assign u_ca_in_304 = col_in_304;
assign u_ca_in_305 = col_in_305;
assign u_ca_in_306 = col_in_306;
assign u_ca_in_307 = col_in_307;
assign u_ca_in_308 = col_in_308;
assign u_ca_in_309 = col_in_309;
assign u_ca_in_310 = col_in_310;
assign u_ca_in_311 = col_in_311;
assign u_ca_in_312 = col_in_312;
assign u_ca_in_313 = col_in_313;
assign u_ca_in_314 = col_in_314;
assign u_ca_in_315 = col_in_315;
assign u_ca_in_316 = col_in_316;
assign u_ca_in_317 = col_in_317;
assign u_ca_in_318 = col_in_318;
assign u_ca_in_319 = col_in_319;
assign u_ca_in_320 = col_in_320;
assign u_ca_in_321 = col_in_321;
assign u_ca_in_322 = col_in_322;
assign u_ca_in_323 = col_in_323;
assign u_ca_in_324 = col_in_324;
assign u_ca_in_325 = col_in_325;
assign u_ca_in_326 = col_in_326;
assign u_ca_in_327 = col_in_327;
assign u_ca_in_328 = col_in_328;
assign u_ca_in_329 = col_in_329;
assign u_ca_in_330 = col_in_330;
assign u_ca_in_331 = col_in_331;
assign u_ca_in_332 = col_in_332;
assign u_ca_in_333 = col_in_333;
assign u_ca_in_334 = col_in_334;
assign u_ca_in_335 = col_in_335;
assign u_ca_in_336 = col_in_336;
assign u_ca_in_337 = col_in_337;
assign u_ca_in_338 = col_in_338;
assign u_ca_in_339 = col_in_339;
assign u_ca_in_340 = col_in_340;
assign u_ca_in_341 = col_in_341;
assign u_ca_in_342 = col_in_342;
assign u_ca_in_343 = col_in_343;
assign u_ca_in_344 = col_in_344;
assign u_ca_in_345 = col_in_345;
assign u_ca_in_346 = col_in_346;
assign u_ca_in_347 = col_in_347;
assign u_ca_in_348 = col_in_348;
assign u_ca_in_349 = col_in_349;
assign u_ca_in_350 = col_in_350;
assign u_ca_in_351 = col_in_351;
assign u_ca_in_352 = col_in_352;
assign u_ca_in_353 = col_in_353;
assign u_ca_in_354 = col_in_354;
assign u_ca_in_355 = col_in_355;
assign u_ca_in_356 = col_in_356;
assign u_ca_in_357 = col_in_357;
assign u_ca_in_358 = col_in_358;
assign u_ca_in_359 = col_in_359;
assign u_ca_in_360 = col_in_360;
assign u_ca_in_361 = col_in_361;
assign u_ca_in_362 = col_in_362;
assign u_ca_in_363 = col_in_363;
assign u_ca_in_364 = col_in_364;
assign u_ca_in_365 = col_in_365;
assign u_ca_in_366 = col_in_366;
assign u_ca_in_367 = col_in_367;
assign u_ca_in_368 = col_in_368;
assign u_ca_in_369 = col_in_369;
assign u_ca_in_370 = col_in_370;
assign u_ca_in_371 = col_in_371;
assign u_ca_in_372 = col_in_372;
assign u_ca_in_373 = col_in_373;
assign u_ca_in_374 = col_in_374;
assign u_ca_in_375 = col_in_375;
assign u_ca_in_376 = col_in_376;
assign u_ca_in_377 = col_in_377;
assign u_ca_in_378 = col_in_378;
assign u_ca_in_379 = col_in_379;
assign u_ca_in_380 = col_in_380;
assign u_ca_in_381 = col_in_381;
assign u_ca_in_382 = col_in_382;
assign u_ca_in_383 = col_in_383;
assign u_ca_in_384 = col_in_384;
assign u_ca_in_385 = col_in_385;
assign u_ca_in_386 = col_in_386;
assign u_ca_in_387 = col_in_387;
assign u_ca_in_388 = col_in_388;
assign u_ca_in_389 = col_in_389;
assign u_ca_in_390 = col_in_390;
assign u_ca_in_391 = col_in_391;
assign u_ca_in_392 = col_in_392;
assign u_ca_in_393 = col_in_393;
assign u_ca_in_394 = col_in_394;
assign u_ca_in_395 = col_in_395;
assign u_ca_in_396 = col_in_396;
assign u_ca_in_397 = col_in_397;
assign u_ca_in_398 = col_in_398;
assign u_ca_in_399 = col_in_399;
assign u_ca_in_400 = col_in_400;
assign u_ca_in_401 = col_in_401;
assign u_ca_in_402 = col_in_402;
assign u_ca_in_403 = col_in_403;
assign u_ca_in_404 = col_in_404;
assign u_ca_in_405 = col_in_405;
assign u_ca_in_406 = col_in_406;
assign u_ca_in_407 = col_in_407;
assign u_ca_in_408 = col_in_408;
assign u_ca_in_409 = col_in_409;
assign u_ca_in_410 = col_in_410;
assign u_ca_in_411 = col_in_411;
assign u_ca_in_412 = col_in_412;
assign u_ca_in_413 = col_in_413;
assign u_ca_in_414 = col_in_414;
assign u_ca_in_415 = col_in_415;
assign u_ca_in_416 = col_in_416;
assign u_ca_in_417 = col_in_417;
assign u_ca_in_418 = col_in_418;
assign u_ca_in_419 = col_in_419;
assign u_ca_in_420 = col_in_420;
assign u_ca_in_421 = col_in_421;
assign u_ca_in_422 = col_in_422;
assign u_ca_in_423 = col_in_423;
assign u_ca_in_424 = col_in_424;
assign u_ca_in_425 = col_in_425;
assign u_ca_in_426 = col_in_426;
assign u_ca_in_427 = col_in_427;
assign u_ca_in_428 = col_in_428;
assign u_ca_in_429 = col_in_429;
assign u_ca_in_430 = col_in_430;
assign u_ca_in_431 = col_in_431;
assign u_ca_in_432 = col_in_432;
assign u_ca_in_433 = col_in_433;
assign u_ca_in_434 = col_in_434;
assign u_ca_in_435 = col_in_435;
assign u_ca_in_436 = col_in_436;
assign u_ca_in_437 = col_in_437;
assign u_ca_in_438 = col_in_438;
assign u_ca_in_439 = col_in_439;
assign u_ca_in_440 = col_in_440;
assign u_ca_in_441 = col_in_441;
assign u_ca_in_442 = col_in_442;
assign u_ca_in_443 = col_in_443;
assign u_ca_in_444 = col_in_444;
assign u_ca_in_445 = col_in_445;
assign u_ca_in_446 = col_in_446;
assign u_ca_in_447 = col_in_447;
assign u_ca_in_448 = col_in_448;
assign u_ca_in_449 = col_in_449;
assign u_ca_in_450 = col_in_450;
assign u_ca_in_451 = col_in_451;
assign u_ca_in_452 = col_in_452;
assign u_ca_in_453 = col_in_453;
assign u_ca_in_454 = col_in_454;
assign u_ca_in_455 = col_in_455;
assign u_ca_in_456 = col_in_456;
assign u_ca_in_457 = col_in_457;
assign u_ca_in_458 = col_in_458;
assign u_ca_in_459 = col_in_459;
assign u_ca_in_460 = col_in_460;
assign u_ca_in_461 = col_in_461;
assign u_ca_in_462 = col_in_462;
assign u_ca_in_463 = col_in_463;
assign u_ca_in_464 = col_in_464;
assign u_ca_in_465 = col_in_465;
assign u_ca_in_466 = col_in_466;
assign u_ca_in_467 = col_in_467;
assign u_ca_in_468 = col_in_468;
assign u_ca_in_469 = col_in_469;
assign u_ca_in_470 = col_in_470;
assign u_ca_in_471 = col_in_471;
assign u_ca_in_472 = col_in_472;
assign u_ca_in_473 = col_in_473;
assign u_ca_in_474 = col_in_474;
assign u_ca_in_475 = col_in_475;
assign u_ca_in_476 = col_in_476;
assign u_ca_in_477 = col_in_477;
assign u_ca_in_478 = col_in_478;
assign u_ca_in_479 = col_in_479;
assign u_ca_in_480 = col_in_480;
assign u_ca_in_481 = col_in_481;
assign u_ca_in_482 = col_in_482;
assign u_ca_in_483 = col_in_483;
assign u_ca_in_484 = col_in_484;
assign u_ca_in_485 = col_in_485;
assign u_ca_in_486 = col_in_486;
assign u_ca_in_487 = col_in_487;
assign u_ca_in_488 = col_in_488;
assign u_ca_in_489 = col_in_489;
assign u_ca_in_490 = col_in_490;
assign u_ca_in_491 = col_in_491;
assign u_ca_in_492 = col_in_492;
assign u_ca_in_493 = col_in_493;
assign u_ca_in_494 = col_in_494;
assign u_ca_in_495 = col_in_495;
assign u_ca_in_496 = col_in_496;
assign u_ca_in_497 = col_in_497;
assign u_ca_in_498 = col_in_498;
assign u_ca_in_499 = col_in_499;
assign u_ca_in_500 = col_in_500;
assign u_ca_in_501 = col_in_501;
assign u_ca_in_502 = col_in_502;
assign u_ca_in_503 = col_in_503;
assign u_ca_in_504 = col_in_504;
assign u_ca_in_505 = col_in_505;
assign u_ca_in_506 = col_in_506;
assign u_ca_in_507 = col_in_507;
assign u_ca_in_508 = col_in_508;
assign u_ca_in_509 = col_in_509;
assign u_ca_in_510 = col_in_510;
assign u_ca_in_511 = col_in_511;
assign u_ca_in_512 = col_in_512;
assign u_ca_in_513 = col_in_513;
assign u_ca_in_514 = col_in_514;
assign u_ca_in_515 = col_in_515;
assign u_ca_in_516 = col_in_516;
assign u_ca_in_517 = col_in_517;
assign u_ca_in_518 = col_in_518;
assign u_ca_in_519 = col_in_519;
assign u_ca_in_520 = col_in_520;
assign u_ca_in_521 = col_in_521;
assign u_ca_in_522 = col_in_522;
assign u_ca_in_523 = col_in_523;
assign u_ca_in_524 = col_in_524;
assign u_ca_in_525 = col_in_525;
assign u_ca_in_526 = col_in_526;
assign u_ca_in_527 = col_in_527;
assign u_ca_in_528 = col_in_528;
assign u_ca_in_529 = col_in_529;
assign u_ca_in_530 = col_in_530;
assign u_ca_in_531 = col_in_531;
assign u_ca_in_532 = col_in_532;
assign u_ca_in_533 = col_in_533;
assign u_ca_in_534 = col_in_534;
assign u_ca_in_535 = col_in_535;
assign u_ca_in_536 = col_in_536;
assign u_ca_in_537 = col_in_537;
assign u_ca_in_538 = col_in_538;
assign u_ca_in_539 = col_in_539;
assign u_ca_in_540 = col_in_540;
assign u_ca_in_541 = col_in_541;
assign u_ca_in_542 = col_in_542;
assign u_ca_in_543 = col_in_543;
assign u_ca_in_544 = col_in_544;
assign u_ca_in_545 = col_in_545;
assign u_ca_in_546 = col_in_546;
assign u_ca_in_547 = col_in_547;
assign u_ca_in_548 = col_in_548;
assign u_ca_in_549 = col_in_549;
assign u_ca_in_550 = col_in_550;
assign u_ca_in_551 = col_in_551;
assign u_ca_in_552 = col_in_552;
assign u_ca_in_553 = col_in_553;
assign u_ca_in_554 = col_in_554;
assign u_ca_in_555 = col_in_555;
assign u_ca_in_556 = col_in_556;
assign u_ca_in_557 = col_in_557;
assign u_ca_in_558 = col_in_558;
assign u_ca_in_559 = col_in_559;
assign u_ca_in_560 = col_in_560;
assign u_ca_in_561 = col_in_561;
assign u_ca_in_562 = col_in_562;
assign u_ca_in_563 = col_in_563;
assign u_ca_in_564 = col_in_564;
assign u_ca_in_565 = col_in_565;
assign u_ca_in_566 = col_in_566;
assign u_ca_in_567 = col_in_567;
assign u_ca_in_568 = col_in_568;
assign u_ca_in_569 = col_in_569;
assign u_ca_in_570 = col_in_570;
assign u_ca_in_571 = col_in_571;
assign u_ca_in_572 = col_in_572;
assign u_ca_in_573 = col_in_573;
assign u_ca_in_574 = col_in_574;
assign u_ca_in_575 = col_in_575;
assign u_ca_in_576 = col_in_576;
assign u_ca_in_577 = col_in_577;
assign u_ca_in_578 = col_in_578;
assign u_ca_in_579 = col_in_579;
assign u_ca_in_580 = col_in_580;
assign u_ca_in_581 = col_in_581;
assign u_ca_in_582 = col_in_582;
assign u_ca_in_583 = col_in_583;
assign u_ca_in_584 = col_in_584;
assign u_ca_in_585 = col_in_585;
assign u_ca_in_586 = col_in_586;
assign u_ca_in_587 = col_in_587;
assign u_ca_in_588 = col_in_588;
assign u_ca_in_589 = col_in_589;
assign u_ca_in_590 = col_in_590;
assign u_ca_in_591 = col_in_591;
assign u_ca_in_592 = col_in_592;
assign u_ca_in_593 = col_in_593;
assign u_ca_in_594 = col_in_594;
assign u_ca_in_595 = col_in_595;
assign u_ca_in_596 = col_in_596;
assign u_ca_in_597 = col_in_597;
assign u_ca_in_598 = col_in_598;
assign u_ca_in_599 = col_in_599;
assign u_ca_in_600 = col_in_600;
assign u_ca_in_601 = col_in_601;
assign u_ca_in_602 = col_in_602;
assign u_ca_in_603 = col_in_603;
assign u_ca_in_604 = col_in_604;
assign u_ca_in_605 = col_in_605;
assign u_ca_in_606 = col_in_606;
assign u_ca_in_607 = col_in_607;
assign u_ca_in_608 = col_in_608;
assign u_ca_in_609 = col_in_609;
assign u_ca_in_610 = col_in_610;
assign u_ca_in_611 = col_in_611;
assign u_ca_in_612 = col_in_612;
assign u_ca_in_613 = col_in_613;
assign u_ca_in_614 = col_in_614;
assign u_ca_in_615 = col_in_615;
assign u_ca_in_616 = col_in_616;
assign u_ca_in_617 = col_in_617;
assign u_ca_in_618 = col_in_618;
assign u_ca_in_619 = col_in_619;
assign u_ca_in_620 = col_in_620;
assign u_ca_in_621 = col_in_621;
assign u_ca_in_622 = col_in_622;
assign u_ca_in_623 = col_in_623;
assign u_ca_in_624 = col_in_624;
assign u_ca_in_625 = col_in_625;
assign u_ca_in_626 = col_in_626;
assign u_ca_in_627 = col_in_627;
assign u_ca_in_628 = col_in_628;
assign u_ca_in_629 = col_in_629;
assign u_ca_in_630 = col_in_630;
assign u_ca_in_631 = col_in_631;
assign u_ca_in_632 = col_in_632;
assign u_ca_in_633 = col_in_633;
assign u_ca_in_634 = col_in_634;
assign u_ca_in_635 = col_in_635;
assign u_ca_in_636 = col_in_636;
assign u_ca_in_637 = col_in_637;
assign u_ca_in_638 = col_in_638;
assign u_ca_in_639 = col_in_639;
assign u_ca_in_640 = col_in_640;
assign u_ca_in_641 = col_in_641;
assign u_ca_in_642 = col_in_642;
assign u_ca_in_643 = col_in_643;
assign u_ca_in_644 = col_in_644;
assign u_ca_in_645 = col_in_645;
assign u_ca_in_646 = col_in_646;
assign u_ca_in_647 = col_in_647;
assign u_ca_in_648 = col_in_648;
assign u_ca_in_649 = col_in_649;
assign u_ca_in_650 = col_in_650;
assign u_ca_in_651 = col_in_651;
assign u_ca_in_652 = col_in_652;
assign u_ca_in_653 = col_in_653;
assign u_ca_in_654 = col_in_654;
assign u_ca_in_655 = col_in_655;
assign u_ca_in_656 = col_in_656;
assign u_ca_in_657 = col_in_657;
assign u_ca_in_658 = col_in_658;
assign u_ca_in_659 = col_in_659;
assign u_ca_in_660 = col_in_660;
assign u_ca_in_661 = col_in_661;
assign u_ca_in_662 = col_in_662;
assign u_ca_in_663 = col_in_663;
assign u_ca_in_664 = col_in_664;
assign u_ca_in_665 = col_in_665;
assign u_ca_in_666 = col_in_666;
assign u_ca_in_667 = col_in_667;
assign u_ca_in_668 = col_in_668;
assign u_ca_in_669 = col_in_669;
assign u_ca_in_670 = col_in_670;
assign u_ca_in_671 = col_in_671;
assign u_ca_in_672 = col_in_672;
assign u_ca_in_673 = col_in_673;
assign u_ca_in_674 = col_in_674;
assign u_ca_in_675 = col_in_675;
assign u_ca_in_676 = col_in_676;
assign u_ca_in_677 = col_in_677;
assign u_ca_in_678 = col_in_678;
assign u_ca_in_679 = col_in_679;
assign u_ca_in_680 = col_in_680;
assign u_ca_in_681 = col_in_681;
assign u_ca_in_682 = col_in_682;
assign u_ca_in_683 = col_in_683;
assign u_ca_in_684 = col_in_684;
assign u_ca_in_685 = col_in_685;
assign u_ca_in_686 = col_in_686;
assign u_ca_in_687 = col_in_687;
assign u_ca_in_688 = col_in_688;
assign u_ca_in_689 = col_in_689;
assign u_ca_in_690 = col_in_690;
assign u_ca_in_691 = col_in_691;
assign u_ca_in_692 = col_in_692;
assign u_ca_in_693 = col_in_693;
assign u_ca_in_694 = col_in_694;
assign u_ca_in_695 = col_in_695;
assign u_ca_in_696 = col_in_696;
assign u_ca_in_697 = col_in_697;
assign u_ca_in_698 = col_in_698;
assign u_ca_in_699 = col_in_699;
assign u_ca_in_700 = col_in_700;
assign u_ca_in_701 = col_in_701;
assign u_ca_in_702 = col_in_702;
assign u_ca_in_703 = col_in_703;
assign u_ca_in_704 = col_in_704;
assign u_ca_in_705 = col_in_705;
assign u_ca_in_706 = col_in_706;
assign u_ca_in_707 = col_in_707;
assign u_ca_in_708 = col_in_708;
assign u_ca_in_709 = col_in_709;
assign u_ca_in_710 = col_in_710;
assign u_ca_in_711 = col_in_711;
assign u_ca_in_712 = col_in_712;
assign u_ca_in_713 = col_in_713;
assign u_ca_in_714 = col_in_714;
assign u_ca_in_715 = col_in_715;
assign u_ca_in_716 = col_in_716;
assign u_ca_in_717 = col_in_717;
assign u_ca_in_718 = col_in_718;
assign u_ca_in_719 = col_in_719;
assign u_ca_in_720 = col_in_720;
assign u_ca_in_721 = col_in_721;
assign u_ca_in_722 = col_in_722;
assign u_ca_in_723 = col_in_723;
assign u_ca_in_724 = col_in_724;
assign u_ca_in_725 = col_in_725;
assign u_ca_in_726 = col_in_726;
assign u_ca_in_727 = col_in_727;
assign u_ca_in_728 = col_in_728;
assign u_ca_in_729 = col_in_729;
assign u_ca_in_730 = col_in_730;
assign u_ca_in_731 = col_in_731;
assign u_ca_in_732 = col_in_732;
assign u_ca_in_733 = col_in_733;
assign u_ca_in_734 = col_in_734;
assign u_ca_in_735 = col_in_735;
assign u_ca_in_736 = col_in_736;
assign u_ca_in_737 = col_in_737;
assign u_ca_in_738 = col_in_738;
assign u_ca_in_739 = col_in_739;
assign u_ca_in_740 = col_in_740;
assign u_ca_in_741 = col_in_741;
assign u_ca_in_742 = col_in_742;
assign u_ca_in_743 = col_in_743;
assign u_ca_in_744 = col_in_744;
assign u_ca_in_745 = col_in_745;
assign u_ca_in_746 = col_in_746;
assign u_ca_in_747 = col_in_747;
assign u_ca_in_748 = col_in_748;
assign u_ca_in_749 = col_in_749;
assign u_ca_in_750 = col_in_750;
assign u_ca_in_751 = col_in_751;
assign u_ca_in_752 = col_in_752;
assign u_ca_in_753 = col_in_753;
assign u_ca_in_754 = col_in_754;
assign u_ca_in_755 = col_in_755;
assign u_ca_in_756 = col_in_756;
assign u_ca_in_757 = col_in_757;
assign u_ca_in_758 = col_in_758;
assign u_ca_in_759 = col_in_759;
assign u_ca_in_760 = col_in_760;
assign u_ca_in_761 = col_in_761;
assign u_ca_in_762 = col_in_762;
assign u_ca_in_763 = col_in_763;
assign u_ca_in_764 = col_in_764;
assign u_ca_in_765 = col_in_765;
assign u_ca_in_766 = col_in_766;
assign u_ca_in_767 = col_in_767;
assign u_ca_in_768 = col_in_768;
assign u_ca_in_769 = col_in_769;
assign u_ca_in_770 = col_in_770;
assign u_ca_in_771 = col_in_771;
assign u_ca_in_772 = col_in_772;
assign u_ca_in_773 = col_in_773;
assign u_ca_in_774 = col_in_774;
assign u_ca_in_775 = col_in_775;
assign u_ca_in_776 = col_in_776;
assign u_ca_in_777 = col_in_777;
assign u_ca_in_778 = col_in_778;
assign u_ca_in_779 = col_in_779;
assign u_ca_in_780 = col_in_780;
assign u_ca_in_781 = col_in_781;
assign u_ca_in_782 = col_in_782;
assign u_ca_in_783 = col_in_783;
assign u_ca_in_784 = col_in_784;
assign u_ca_in_785 = col_in_785;
assign u_ca_in_786 = col_in_786;
assign u_ca_in_787 = col_in_787;
assign u_ca_in_788 = col_in_788;
assign u_ca_in_789 = col_in_789;
assign u_ca_in_790 = col_in_790;
assign u_ca_in_791 = col_in_791;
assign u_ca_in_792 = col_in_792;
assign u_ca_in_793 = col_in_793;
assign u_ca_in_794 = col_in_794;
assign u_ca_in_795 = col_in_795;
assign u_ca_in_796 = col_in_796;
assign u_ca_in_797 = col_in_797;
assign u_ca_in_798 = col_in_798;
assign u_ca_in_799 = col_in_799;
assign u_ca_in_800 = col_in_800;
assign u_ca_in_801 = col_in_801;
assign u_ca_in_802 = col_in_802;
assign u_ca_in_803 = col_in_803;
assign u_ca_in_804 = col_in_804;
assign u_ca_in_805 = col_in_805;
assign u_ca_in_806 = col_in_806;
assign u_ca_in_807 = col_in_807;
assign u_ca_in_808 = col_in_808;
assign u_ca_in_809 = col_in_809;
assign u_ca_in_810 = col_in_810;
assign u_ca_in_811 = col_in_811;
assign u_ca_in_812 = col_in_812;
assign u_ca_in_813 = col_in_813;
assign u_ca_in_814 = col_in_814;
assign u_ca_in_815 = col_in_815;
assign u_ca_in_816 = col_in_816;
assign u_ca_in_817 = col_in_817;
assign u_ca_in_818 = col_in_818;
assign u_ca_in_819 = col_in_819;
assign u_ca_in_820 = col_in_820;
assign u_ca_in_821 = col_in_821;
assign u_ca_in_822 = col_in_822;
assign u_ca_in_823 = col_in_823;
assign u_ca_in_824 = col_in_824;
assign u_ca_in_825 = col_in_825;
assign u_ca_in_826 = col_in_826;
assign u_ca_in_827 = col_in_827;
assign u_ca_in_828 = col_in_828;
assign u_ca_in_829 = col_in_829;
assign u_ca_in_830 = col_in_830;
assign u_ca_in_831 = col_in_831;
assign u_ca_in_832 = col_in_832;
assign u_ca_in_833 = col_in_833;
assign u_ca_in_834 = col_in_834;
assign u_ca_in_835 = col_in_835;
assign u_ca_in_836 = col_in_836;
assign u_ca_in_837 = col_in_837;
assign u_ca_in_838 = col_in_838;
assign u_ca_in_839 = col_in_839;
assign u_ca_in_840 = col_in_840;
assign u_ca_in_841 = col_in_841;
assign u_ca_in_842 = col_in_842;
assign u_ca_in_843 = col_in_843;
assign u_ca_in_844 = col_in_844;
assign u_ca_in_845 = col_in_845;
assign u_ca_in_846 = col_in_846;
assign u_ca_in_847 = col_in_847;
assign u_ca_in_848 = col_in_848;
assign u_ca_in_849 = col_in_849;
assign u_ca_in_850 = col_in_850;
assign u_ca_in_851 = col_in_851;
assign u_ca_in_852 = col_in_852;
assign u_ca_in_853 = col_in_853;
assign u_ca_in_854 = col_in_854;
assign u_ca_in_855 = col_in_855;
assign u_ca_in_856 = col_in_856;
assign u_ca_in_857 = col_in_857;
assign u_ca_in_858 = col_in_858;
assign u_ca_in_859 = col_in_859;
assign u_ca_in_860 = col_in_860;
assign u_ca_in_861 = col_in_861;
assign u_ca_in_862 = col_in_862;
assign u_ca_in_863 = col_in_863;
assign u_ca_in_864 = col_in_864;
assign u_ca_in_865 = col_in_865;
assign u_ca_in_866 = col_in_866;
assign u_ca_in_867 = col_in_867;
assign u_ca_in_868 = col_in_868;
assign u_ca_in_869 = col_in_869;
assign u_ca_in_870 = col_in_870;
assign u_ca_in_871 = col_in_871;
assign u_ca_in_872 = col_in_872;
assign u_ca_in_873 = col_in_873;
assign u_ca_in_874 = col_in_874;
assign u_ca_in_875 = col_in_875;
assign u_ca_in_876 = col_in_876;
assign u_ca_in_877 = col_in_877;
assign u_ca_in_878 = col_in_878;
assign u_ca_in_879 = col_in_879;
assign u_ca_in_880 = col_in_880;
assign u_ca_in_881 = col_in_881;
assign u_ca_in_882 = col_in_882;
assign u_ca_in_883 = col_in_883;
assign u_ca_in_884 = col_in_884;
assign u_ca_in_885 = col_in_885;
assign u_ca_in_886 = col_in_886;
assign u_ca_in_887 = col_in_887;
assign u_ca_in_888 = col_in_888;
assign u_ca_in_889 = col_in_889;
assign u_ca_in_890 = col_in_890;
assign u_ca_in_891 = col_in_891;
assign u_ca_in_892 = col_in_892;
assign u_ca_in_893 = col_in_893;
assign u_ca_in_894 = col_in_894;
assign u_ca_in_895 = col_in_895;
assign u_ca_in_896 = col_in_896;
assign u_ca_in_897 = col_in_897;
assign u_ca_in_898 = col_in_898;
assign u_ca_in_899 = col_in_899;
assign u_ca_in_900 = col_in_900;
assign u_ca_in_901 = col_in_901;
assign u_ca_in_902 = col_in_902;
assign u_ca_in_903 = col_in_903;
assign u_ca_in_904 = col_in_904;
assign u_ca_in_905 = col_in_905;
assign u_ca_in_906 = col_in_906;
assign u_ca_in_907 = col_in_907;
assign u_ca_in_908 = col_in_908;
assign u_ca_in_909 = col_in_909;
assign u_ca_in_910 = col_in_910;
assign u_ca_in_911 = col_in_911;
assign u_ca_in_912 = col_in_912;
assign u_ca_in_913 = col_in_913;
assign u_ca_in_914 = col_in_914;
assign u_ca_in_915 = col_in_915;
assign u_ca_in_916 = col_in_916;
assign u_ca_in_917 = col_in_917;
assign u_ca_in_918 = col_in_918;
assign u_ca_in_919 = col_in_919;
assign u_ca_in_920 = col_in_920;
assign u_ca_in_921 = col_in_921;
assign u_ca_in_922 = col_in_922;
assign u_ca_in_923 = col_in_923;
assign u_ca_in_924 = col_in_924;
assign u_ca_in_925 = col_in_925;
assign u_ca_in_926 = col_in_926;
assign u_ca_in_927 = col_in_927;
assign u_ca_in_928 = col_in_928;
assign u_ca_in_929 = col_in_929;
assign u_ca_in_930 = col_in_930;
assign u_ca_in_931 = col_in_931;
assign u_ca_in_932 = col_in_932;
assign u_ca_in_933 = col_in_933;
assign u_ca_in_934 = col_in_934;
assign u_ca_in_935 = col_in_935;
assign u_ca_in_936 = col_in_936;
assign u_ca_in_937 = col_in_937;
assign u_ca_in_938 = col_in_938;
assign u_ca_in_939 = col_in_939;
assign u_ca_in_940 = col_in_940;
assign u_ca_in_941 = col_in_941;
assign u_ca_in_942 = col_in_942;
assign u_ca_in_943 = col_in_943;
assign u_ca_in_944 = col_in_944;
assign u_ca_in_945 = col_in_945;
assign u_ca_in_946 = col_in_946;
assign u_ca_in_947 = col_in_947;
assign u_ca_in_948 = col_in_948;
assign u_ca_in_949 = col_in_949;
assign u_ca_in_950 = col_in_950;
assign u_ca_in_951 = col_in_951;
assign u_ca_in_952 = col_in_952;
assign u_ca_in_953 = col_in_953;
assign u_ca_in_954 = col_in_954;
assign u_ca_in_955 = col_in_955;
assign u_ca_in_956 = col_in_956;
assign u_ca_in_957 = col_in_957;
assign u_ca_in_958 = col_in_958;
assign u_ca_in_959 = col_in_959;
assign u_ca_in_960 = col_in_960;
assign u_ca_in_961 = col_in_961;
assign u_ca_in_962 = col_in_962;
assign u_ca_in_963 = col_in_963;
assign u_ca_in_964 = col_in_964;
assign u_ca_in_965 = col_in_965;
assign u_ca_in_966 = col_in_966;
assign u_ca_in_967 = col_in_967;
assign u_ca_in_968 = col_in_968;
assign u_ca_in_969 = col_in_969;
assign u_ca_in_970 = col_in_970;
assign u_ca_in_971 = col_in_971;
assign u_ca_in_972 = col_in_972;
assign u_ca_in_973 = col_in_973;
assign u_ca_in_974 = col_in_974;
assign u_ca_in_975 = col_in_975;
assign u_ca_in_976 = col_in_976;
assign u_ca_in_977 = col_in_977;
assign u_ca_in_978 = col_in_978;
assign u_ca_in_979 = col_in_979;
assign u_ca_in_980 = col_in_980;
assign u_ca_in_981 = col_in_981;
assign u_ca_in_982 = col_in_982;
assign u_ca_in_983 = col_in_983;
assign u_ca_in_984 = col_in_984;
assign u_ca_in_985 = col_in_985;
assign u_ca_in_986 = col_in_986;
assign u_ca_in_987 = col_in_987;
assign u_ca_in_988 = col_in_988;
assign u_ca_in_989 = col_in_989;
assign u_ca_in_990 = col_in_990;
assign u_ca_in_991 = col_in_991;
assign u_ca_in_992 = col_in_992;
assign u_ca_in_993 = col_in_993;
assign u_ca_in_994 = col_in_994;
assign u_ca_in_995 = col_in_995;
assign u_ca_in_996 = col_in_996;
assign u_ca_in_997 = col_in_997;
assign u_ca_in_998 = col_in_998;
assign u_ca_in_999 = col_in_999;
assign u_ca_in_1000 = col_in_1000;
assign u_ca_in_1001 = col_in_1001;
assign u_ca_in_1002 = col_in_1002;
assign u_ca_in_1003 = col_in_1003;
assign u_ca_in_1004 = col_in_1004;
assign u_ca_in_1005 = col_in_1005;
assign u_ca_in_1006 = col_in_1006;
assign u_ca_in_1007 = col_in_1007;
assign u_ca_in_1008 = col_in_1008;
assign u_ca_in_1009 = col_in_1009;
assign u_ca_in_1010 = col_in_1010;
assign u_ca_in_1011 = col_in_1011;
assign u_ca_in_1012 = col_in_1012;
assign u_ca_in_1013 = col_in_1013;
assign u_ca_in_1014 = col_in_1014;
assign u_ca_in_1015 = col_in_1015;
assign u_ca_in_1016 = col_in_1016;
assign u_ca_in_1017 = col_in_1017;
assign u_ca_in_1018 = col_in_1018;
assign u_ca_in_1019 = col_in_1019;
assign u_ca_in_1020 = col_in_1020;
assign u_ca_in_1021 = col_in_1021;
assign u_ca_in_1022 = col_in_1022;
assign u_ca_in_1023 = col_in_1023;
assign u_ca_in_1024 = col_in_1024;
assign u_ca_in_1025 = col_in_1025;
assign u_ca_in_1026 = col_in_1026;
assign u_ca_in_1027 = col_in_1027;
assign u_ca_in_1028 = col_in_1028;
assign u_ca_in_1029 = col_in_1029;
assign u_ca_in_1030 = col_in_1030;
assign u_ca_in_1031 = col_in_1031;
assign u_ca_in_1032 = col_in_1032;


//---------------------------------------------------------



//--compressor_array---------------------------------------
compressor_12_8 u_ca_12_8_0(.d_in(u_ca_in_0), .d_out(u_ca_out_0));
compressor_12_8 u_ca_12_8_1(.d_in(u_ca_in_1), .d_out(u_ca_out_1));
compressor_12_8 u_ca_12_8_2(.d_in(u_ca_in_2), .d_out(u_ca_out_2));
compressor_12_8 u_ca_12_8_3(.d_in(u_ca_in_3), .d_out(u_ca_out_3));
compressor_12_8 u_ca_12_8_4(.d_in(u_ca_in_4), .d_out(u_ca_out_4));
compressor_12_8 u_ca_12_8_5(.d_in(u_ca_in_5), .d_out(u_ca_out_5));
compressor_12_8 u_ca_12_8_6(.d_in(u_ca_in_6), .d_out(u_ca_out_6));
compressor_12_8 u_ca_12_8_7(.d_in(u_ca_in_7), .d_out(u_ca_out_7));
compressor_12_8 u_ca_12_8_8(.d_in(u_ca_in_8), .d_out(u_ca_out_8));
compressor_12_8 u_ca_12_8_9(.d_in(u_ca_in_9), .d_out(u_ca_out_9));
compressor_12_8 u_ca_12_8_10(.d_in(u_ca_in_10), .d_out(u_ca_out_10));
compressor_12_8 u_ca_12_8_11(.d_in(u_ca_in_11), .d_out(u_ca_out_11));
compressor_12_8 u_ca_12_8_12(.d_in(u_ca_in_12), .d_out(u_ca_out_12));
compressor_12_8 u_ca_12_8_13(.d_in(u_ca_in_13), .d_out(u_ca_out_13));
compressor_12_8 u_ca_12_8_14(.d_in(u_ca_in_14), .d_out(u_ca_out_14));
compressor_12_8 u_ca_12_8_15(.d_in(u_ca_in_15), .d_out(u_ca_out_15));
compressor_12_8 u_ca_12_8_16(.d_in(u_ca_in_16), .d_out(u_ca_out_16));
compressor_12_8 u_ca_12_8_17(.d_in(u_ca_in_17), .d_out(u_ca_out_17));
compressor_12_8 u_ca_12_8_18(.d_in(u_ca_in_18), .d_out(u_ca_out_18));
compressor_12_8 u_ca_12_8_19(.d_in(u_ca_in_19), .d_out(u_ca_out_19));
compressor_12_8 u_ca_12_8_20(.d_in(u_ca_in_20), .d_out(u_ca_out_20));
compressor_12_8 u_ca_12_8_21(.d_in(u_ca_in_21), .d_out(u_ca_out_21));
compressor_12_8 u_ca_12_8_22(.d_in(u_ca_in_22), .d_out(u_ca_out_22));
compressor_12_8 u_ca_12_8_23(.d_in(u_ca_in_23), .d_out(u_ca_out_23));
compressor_12_8 u_ca_12_8_24(.d_in(u_ca_in_24), .d_out(u_ca_out_24));
compressor_12_8 u_ca_12_8_25(.d_in(u_ca_in_25), .d_out(u_ca_out_25));
compressor_12_8 u_ca_12_8_26(.d_in(u_ca_in_26), .d_out(u_ca_out_26));
compressor_12_8 u_ca_12_8_27(.d_in(u_ca_in_27), .d_out(u_ca_out_27));
compressor_12_8 u_ca_12_8_28(.d_in(u_ca_in_28), .d_out(u_ca_out_28));
compressor_12_8 u_ca_12_8_29(.d_in(u_ca_in_29), .d_out(u_ca_out_29));
compressor_12_8 u_ca_12_8_30(.d_in(u_ca_in_30), .d_out(u_ca_out_30));
compressor_12_8 u_ca_12_8_31(.d_in(u_ca_in_31), .d_out(u_ca_out_31));
compressor_12_8 u_ca_12_8_32(.d_in(u_ca_in_32), .d_out(u_ca_out_32));
compressor_12_8 u_ca_12_8_33(.d_in(u_ca_in_33), .d_out(u_ca_out_33));
compressor_12_8 u_ca_12_8_34(.d_in(u_ca_in_34), .d_out(u_ca_out_34));
compressor_12_8 u_ca_12_8_35(.d_in(u_ca_in_35), .d_out(u_ca_out_35));
compressor_12_8 u_ca_12_8_36(.d_in(u_ca_in_36), .d_out(u_ca_out_36));
compressor_12_8 u_ca_12_8_37(.d_in(u_ca_in_37), .d_out(u_ca_out_37));
compressor_12_8 u_ca_12_8_38(.d_in(u_ca_in_38), .d_out(u_ca_out_38));
compressor_12_8 u_ca_12_8_39(.d_in(u_ca_in_39), .d_out(u_ca_out_39));
compressor_12_8 u_ca_12_8_40(.d_in(u_ca_in_40), .d_out(u_ca_out_40));
compressor_12_8 u_ca_12_8_41(.d_in(u_ca_in_41), .d_out(u_ca_out_41));
compressor_12_8 u_ca_12_8_42(.d_in(u_ca_in_42), .d_out(u_ca_out_42));
compressor_12_8 u_ca_12_8_43(.d_in(u_ca_in_43), .d_out(u_ca_out_43));
compressor_12_8 u_ca_12_8_44(.d_in(u_ca_in_44), .d_out(u_ca_out_44));
compressor_12_8 u_ca_12_8_45(.d_in(u_ca_in_45), .d_out(u_ca_out_45));
compressor_12_8 u_ca_12_8_46(.d_in(u_ca_in_46), .d_out(u_ca_out_46));
compressor_12_8 u_ca_12_8_47(.d_in(u_ca_in_47), .d_out(u_ca_out_47));
compressor_12_8 u_ca_12_8_48(.d_in(u_ca_in_48), .d_out(u_ca_out_48));
compressor_12_8 u_ca_12_8_49(.d_in(u_ca_in_49), .d_out(u_ca_out_49));
compressor_12_8 u_ca_12_8_50(.d_in(u_ca_in_50), .d_out(u_ca_out_50));
compressor_12_8 u_ca_12_8_51(.d_in(u_ca_in_51), .d_out(u_ca_out_51));
compressor_12_8 u_ca_12_8_52(.d_in(u_ca_in_52), .d_out(u_ca_out_52));
compressor_12_8 u_ca_12_8_53(.d_in(u_ca_in_53), .d_out(u_ca_out_53));
compressor_12_8 u_ca_12_8_54(.d_in(u_ca_in_54), .d_out(u_ca_out_54));
compressor_12_8 u_ca_12_8_55(.d_in(u_ca_in_55), .d_out(u_ca_out_55));
compressor_12_8 u_ca_12_8_56(.d_in(u_ca_in_56), .d_out(u_ca_out_56));
compressor_12_8 u_ca_12_8_57(.d_in(u_ca_in_57), .d_out(u_ca_out_57));
compressor_12_8 u_ca_12_8_58(.d_in(u_ca_in_58), .d_out(u_ca_out_58));
compressor_12_8 u_ca_12_8_59(.d_in(u_ca_in_59), .d_out(u_ca_out_59));
compressor_12_8 u_ca_12_8_60(.d_in(u_ca_in_60), .d_out(u_ca_out_60));
compressor_12_8 u_ca_12_8_61(.d_in(u_ca_in_61), .d_out(u_ca_out_61));
compressor_12_8 u_ca_12_8_62(.d_in(u_ca_in_62), .d_out(u_ca_out_62));
compressor_12_8 u_ca_12_8_63(.d_in(u_ca_in_63), .d_out(u_ca_out_63));
compressor_12_8 u_ca_12_8_64(.d_in(u_ca_in_64), .d_out(u_ca_out_64));
compressor_12_8 u_ca_12_8_65(.d_in(u_ca_in_65), .d_out(u_ca_out_65));
compressor_12_8 u_ca_12_8_66(.d_in(u_ca_in_66), .d_out(u_ca_out_66));
compressor_12_8 u_ca_12_8_67(.d_in(u_ca_in_67), .d_out(u_ca_out_67));
compressor_12_8 u_ca_12_8_68(.d_in(u_ca_in_68), .d_out(u_ca_out_68));
compressor_12_8 u_ca_12_8_69(.d_in(u_ca_in_69), .d_out(u_ca_out_69));
compressor_12_8 u_ca_12_8_70(.d_in(u_ca_in_70), .d_out(u_ca_out_70));
compressor_12_8 u_ca_12_8_71(.d_in(u_ca_in_71), .d_out(u_ca_out_71));
compressor_12_8 u_ca_12_8_72(.d_in(u_ca_in_72), .d_out(u_ca_out_72));
compressor_12_8 u_ca_12_8_73(.d_in(u_ca_in_73), .d_out(u_ca_out_73));
compressor_12_8 u_ca_12_8_74(.d_in(u_ca_in_74), .d_out(u_ca_out_74));
compressor_12_8 u_ca_12_8_75(.d_in(u_ca_in_75), .d_out(u_ca_out_75));
compressor_12_8 u_ca_12_8_76(.d_in(u_ca_in_76), .d_out(u_ca_out_76));
compressor_12_8 u_ca_12_8_77(.d_in(u_ca_in_77), .d_out(u_ca_out_77));
compressor_12_8 u_ca_12_8_78(.d_in(u_ca_in_78), .d_out(u_ca_out_78));
compressor_12_8 u_ca_12_8_79(.d_in(u_ca_in_79), .d_out(u_ca_out_79));
compressor_12_8 u_ca_12_8_80(.d_in(u_ca_in_80), .d_out(u_ca_out_80));
compressor_12_8 u_ca_12_8_81(.d_in(u_ca_in_81), .d_out(u_ca_out_81));
compressor_12_8 u_ca_12_8_82(.d_in(u_ca_in_82), .d_out(u_ca_out_82));
compressor_12_8 u_ca_12_8_83(.d_in(u_ca_in_83), .d_out(u_ca_out_83));
compressor_12_8 u_ca_12_8_84(.d_in(u_ca_in_84), .d_out(u_ca_out_84));
compressor_12_8 u_ca_12_8_85(.d_in(u_ca_in_85), .d_out(u_ca_out_85));
compressor_12_8 u_ca_12_8_86(.d_in(u_ca_in_86), .d_out(u_ca_out_86));
compressor_12_8 u_ca_12_8_87(.d_in(u_ca_in_87), .d_out(u_ca_out_87));
compressor_12_8 u_ca_12_8_88(.d_in(u_ca_in_88), .d_out(u_ca_out_88));
compressor_12_8 u_ca_12_8_89(.d_in(u_ca_in_89), .d_out(u_ca_out_89));
compressor_12_8 u_ca_12_8_90(.d_in(u_ca_in_90), .d_out(u_ca_out_90));
compressor_12_8 u_ca_12_8_91(.d_in(u_ca_in_91), .d_out(u_ca_out_91));
compressor_12_8 u_ca_12_8_92(.d_in(u_ca_in_92), .d_out(u_ca_out_92));
compressor_12_8 u_ca_12_8_93(.d_in(u_ca_in_93), .d_out(u_ca_out_93));
compressor_12_8 u_ca_12_8_94(.d_in(u_ca_in_94), .d_out(u_ca_out_94));
compressor_12_8 u_ca_12_8_95(.d_in(u_ca_in_95), .d_out(u_ca_out_95));
compressor_12_8 u_ca_12_8_96(.d_in(u_ca_in_96), .d_out(u_ca_out_96));
compressor_12_8 u_ca_12_8_97(.d_in(u_ca_in_97), .d_out(u_ca_out_97));
compressor_12_8 u_ca_12_8_98(.d_in(u_ca_in_98), .d_out(u_ca_out_98));
compressor_12_8 u_ca_12_8_99(.d_in(u_ca_in_99), .d_out(u_ca_out_99));
compressor_12_8 u_ca_12_8_100(.d_in(u_ca_in_100), .d_out(u_ca_out_100));
compressor_12_8 u_ca_12_8_101(.d_in(u_ca_in_101), .d_out(u_ca_out_101));
compressor_12_8 u_ca_12_8_102(.d_in(u_ca_in_102), .d_out(u_ca_out_102));
compressor_12_8 u_ca_12_8_103(.d_in(u_ca_in_103), .d_out(u_ca_out_103));
compressor_12_8 u_ca_12_8_104(.d_in(u_ca_in_104), .d_out(u_ca_out_104));
compressor_12_8 u_ca_12_8_105(.d_in(u_ca_in_105), .d_out(u_ca_out_105));
compressor_12_8 u_ca_12_8_106(.d_in(u_ca_in_106), .d_out(u_ca_out_106));
compressor_12_8 u_ca_12_8_107(.d_in(u_ca_in_107), .d_out(u_ca_out_107));
compressor_12_8 u_ca_12_8_108(.d_in(u_ca_in_108), .d_out(u_ca_out_108));
compressor_12_8 u_ca_12_8_109(.d_in(u_ca_in_109), .d_out(u_ca_out_109));
compressor_12_8 u_ca_12_8_110(.d_in(u_ca_in_110), .d_out(u_ca_out_110));
compressor_12_8 u_ca_12_8_111(.d_in(u_ca_in_111), .d_out(u_ca_out_111));
compressor_12_8 u_ca_12_8_112(.d_in(u_ca_in_112), .d_out(u_ca_out_112));
compressor_12_8 u_ca_12_8_113(.d_in(u_ca_in_113), .d_out(u_ca_out_113));
compressor_12_8 u_ca_12_8_114(.d_in(u_ca_in_114), .d_out(u_ca_out_114));
compressor_12_8 u_ca_12_8_115(.d_in(u_ca_in_115), .d_out(u_ca_out_115));
compressor_12_8 u_ca_12_8_116(.d_in(u_ca_in_116), .d_out(u_ca_out_116));
compressor_12_8 u_ca_12_8_117(.d_in(u_ca_in_117), .d_out(u_ca_out_117));
compressor_12_8 u_ca_12_8_118(.d_in(u_ca_in_118), .d_out(u_ca_out_118));
compressor_12_8 u_ca_12_8_119(.d_in(u_ca_in_119), .d_out(u_ca_out_119));
compressor_12_8 u_ca_12_8_120(.d_in(u_ca_in_120), .d_out(u_ca_out_120));
compressor_12_8 u_ca_12_8_121(.d_in(u_ca_in_121), .d_out(u_ca_out_121));
compressor_12_8 u_ca_12_8_122(.d_in(u_ca_in_122), .d_out(u_ca_out_122));
compressor_12_8 u_ca_12_8_123(.d_in(u_ca_in_123), .d_out(u_ca_out_123));
compressor_12_8 u_ca_12_8_124(.d_in(u_ca_in_124), .d_out(u_ca_out_124));
compressor_12_8 u_ca_12_8_125(.d_in(u_ca_in_125), .d_out(u_ca_out_125));
compressor_12_8 u_ca_12_8_126(.d_in(u_ca_in_126), .d_out(u_ca_out_126));
compressor_12_8 u_ca_12_8_127(.d_in(u_ca_in_127), .d_out(u_ca_out_127));
compressor_12_8 u_ca_12_8_128(.d_in(u_ca_in_128), .d_out(u_ca_out_128));
compressor_12_8 u_ca_12_8_129(.d_in(u_ca_in_129), .d_out(u_ca_out_129));
compressor_12_8 u_ca_12_8_130(.d_in(u_ca_in_130), .d_out(u_ca_out_130));
compressor_12_8 u_ca_12_8_131(.d_in(u_ca_in_131), .d_out(u_ca_out_131));
compressor_12_8 u_ca_12_8_132(.d_in(u_ca_in_132), .d_out(u_ca_out_132));
compressor_12_8 u_ca_12_8_133(.d_in(u_ca_in_133), .d_out(u_ca_out_133));
compressor_12_8 u_ca_12_8_134(.d_in(u_ca_in_134), .d_out(u_ca_out_134));
compressor_12_8 u_ca_12_8_135(.d_in(u_ca_in_135), .d_out(u_ca_out_135));
compressor_12_8 u_ca_12_8_136(.d_in(u_ca_in_136), .d_out(u_ca_out_136));
compressor_12_8 u_ca_12_8_137(.d_in(u_ca_in_137), .d_out(u_ca_out_137));
compressor_12_8 u_ca_12_8_138(.d_in(u_ca_in_138), .d_out(u_ca_out_138));
compressor_12_8 u_ca_12_8_139(.d_in(u_ca_in_139), .d_out(u_ca_out_139));
compressor_12_8 u_ca_12_8_140(.d_in(u_ca_in_140), .d_out(u_ca_out_140));
compressor_12_8 u_ca_12_8_141(.d_in(u_ca_in_141), .d_out(u_ca_out_141));
compressor_12_8 u_ca_12_8_142(.d_in(u_ca_in_142), .d_out(u_ca_out_142));
compressor_12_8 u_ca_12_8_143(.d_in(u_ca_in_143), .d_out(u_ca_out_143));
compressor_12_8 u_ca_12_8_144(.d_in(u_ca_in_144), .d_out(u_ca_out_144));
compressor_12_8 u_ca_12_8_145(.d_in(u_ca_in_145), .d_out(u_ca_out_145));
compressor_12_8 u_ca_12_8_146(.d_in(u_ca_in_146), .d_out(u_ca_out_146));
compressor_12_8 u_ca_12_8_147(.d_in(u_ca_in_147), .d_out(u_ca_out_147));
compressor_12_8 u_ca_12_8_148(.d_in(u_ca_in_148), .d_out(u_ca_out_148));
compressor_12_8 u_ca_12_8_149(.d_in(u_ca_in_149), .d_out(u_ca_out_149));
compressor_12_8 u_ca_12_8_150(.d_in(u_ca_in_150), .d_out(u_ca_out_150));
compressor_12_8 u_ca_12_8_151(.d_in(u_ca_in_151), .d_out(u_ca_out_151));
compressor_12_8 u_ca_12_8_152(.d_in(u_ca_in_152), .d_out(u_ca_out_152));
compressor_12_8 u_ca_12_8_153(.d_in(u_ca_in_153), .d_out(u_ca_out_153));
compressor_12_8 u_ca_12_8_154(.d_in(u_ca_in_154), .d_out(u_ca_out_154));
compressor_12_8 u_ca_12_8_155(.d_in(u_ca_in_155), .d_out(u_ca_out_155));
compressor_12_8 u_ca_12_8_156(.d_in(u_ca_in_156), .d_out(u_ca_out_156));
compressor_12_8 u_ca_12_8_157(.d_in(u_ca_in_157), .d_out(u_ca_out_157));
compressor_12_8 u_ca_12_8_158(.d_in(u_ca_in_158), .d_out(u_ca_out_158));
compressor_12_8 u_ca_12_8_159(.d_in(u_ca_in_159), .d_out(u_ca_out_159));
compressor_12_8 u_ca_12_8_160(.d_in(u_ca_in_160), .d_out(u_ca_out_160));
compressor_12_8 u_ca_12_8_161(.d_in(u_ca_in_161), .d_out(u_ca_out_161));
compressor_12_8 u_ca_12_8_162(.d_in(u_ca_in_162), .d_out(u_ca_out_162));
compressor_12_8 u_ca_12_8_163(.d_in(u_ca_in_163), .d_out(u_ca_out_163));
compressor_12_8 u_ca_12_8_164(.d_in(u_ca_in_164), .d_out(u_ca_out_164));
compressor_12_8 u_ca_12_8_165(.d_in(u_ca_in_165), .d_out(u_ca_out_165));
compressor_12_8 u_ca_12_8_166(.d_in(u_ca_in_166), .d_out(u_ca_out_166));
compressor_12_8 u_ca_12_8_167(.d_in(u_ca_in_167), .d_out(u_ca_out_167));
compressor_12_8 u_ca_12_8_168(.d_in(u_ca_in_168), .d_out(u_ca_out_168));
compressor_12_8 u_ca_12_8_169(.d_in(u_ca_in_169), .d_out(u_ca_out_169));
compressor_12_8 u_ca_12_8_170(.d_in(u_ca_in_170), .d_out(u_ca_out_170));
compressor_12_8 u_ca_12_8_171(.d_in(u_ca_in_171), .d_out(u_ca_out_171));
compressor_12_8 u_ca_12_8_172(.d_in(u_ca_in_172), .d_out(u_ca_out_172));
compressor_12_8 u_ca_12_8_173(.d_in(u_ca_in_173), .d_out(u_ca_out_173));
compressor_12_8 u_ca_12_8_174(.d_in(u_ca_in_174), .d_out(u_ca_out_174));
compressor_12_8 u_ca_12_8_175(.d_in(u_ca_in_175), .d_out(u_ca_out_175));
compressor_12_8 u_ca_12_8_176(.d_in(u_ca_in_176), .d_out(u_ca_out_176));
compressor_12_8 u_ca_12_8_177(.d_in(u_ca_in_177), .d_out(u_ca_out_177));
compressor_12_8 u_ca_12_8_178(.d_in(u_ca_in_178), .d_out(u_ca_out_178));
compressor_12_8 u_ca_12_8_179(.d_in(u_ca_in_179), .d_out(u_ca_out_179));
compressor_12_8 u_ca_12_8_180(.d_in(u_ca_in_180), .d_out(u_ca_out_180));
compressor_12_8 u_ca_12_8_181(.d_in(u_ca_in_181), .d_out(u_ca_out_181));
compressor_12_8 u_ca_12_8_182(.d_in(u_ca_in_182), .d_out(u_ca_out_182));
compressor_12_8 u_ca_12_8_183(.d_in(u_ca_in_183), .d_out(u_ca_out_183));
compressor_12_8 u_ca_12_8_184(.d_in(u_ca_in_184), .d_out(u_ca_out_184));
compressor_12_8 u_ca_12_8_185(.d_in(u_ca_in_185), .d_out(u_ca_out_185));
compressor_12_8 u_ca_12_8_186(.d_in(u_ca_in_186), .d_out(u_ca_out_186));
compressor_12_8 u_ca_12_8_187(.d_in(u_ca_in_187), .d_out(u_ca_out_187));
compressor_12_8 u_ca_12_8_188(.d_in(u_ca_in_188), .d_out(u_ca_out_188));
compressor_12_8 u_ca_12_8_189(.d_in(u_ca_in_189), .d_out(u_ca_out_189));
compressor_12_8 u_ca_12_8_190(.d_in(u_ca_in_190), .d_out(u_ca_out_190));
compressor_12_8 u_ca_12_8_191(.d_in(u_ca_in_191), .d_out(u_ca_out_191));
compressor_12_8 u_ca_12_8_192(.d_in(u_ca_in_192), .d_out(u_ca_out_192));
compressor_12_8 u_ca_12_8_193(.d_in(u_ca_in_193), .d_out(u_ca_out_193));
compressor_12_8 u_ca_12_8_194(.d_in(u_ca_in_194), .d_out(u_ca_out_194));
compressor_12_8 u_ca_12_8_195(.d_in(u_ca_in_195), .d_out(u_ca_out_195));
compressor_12_8 u_ca_12_8_196(.d_in(u_ca_in_196), .d_out(u_ca_out_196));
compressor_12_8 u_ca_12_8_197(.d_in(u_ca_in_197), .d_out(u_ca_out_197));
compressor_12_8 u_ca_12_8_198(.d_in(u_ca_in_198), .d_out(u_ca_out_198));
compressor_12_8 u_ca_12_8_199(.d_in(u_ca_in_199), .d_out(u_ca_out_199));
compressor_12_8 u_ca_12_8_200(.d_in(u_ca_in_200), .d_out(u_ca_out_200));
compressor_12_8 u_ca_12_8_201(.d_in(u_ca_in_201), .d_out(u_ca_out_201));
compressor_12_8 u_ca_12_8_202(.d_in(u_ca_in_202), .d_out(u_ca_out_202));
compressor_12_8 u_ca_12_8_203(.d_in(u_ca_in_203), .d_out(u_ca_out_203));
compressor_12_8 u_ca_12_8_204(.d_in(u_ca_in_204), .d_out(u_ca_out_204));
compressor_12_8 u_ca_12_8_205(.d_in(u_ca_in_205), .d_out(u_ca_out_205));
compressor_12_8 u_ca_12_8_206(.d_in(u_ca_in_206), .d_out(u_ca_out_206));
compressor_12_8 u_ca_12_8_207(.d_in(u_ca_in_207), .d_out(u_ca_out_207));
compressor_12_8 u_ca_12_8_208(.d_in(u_ca_in_208), .d_out(u_ca_out_208));
compressor_12_8 u_ca_12_8_209(.d_in(u_ca_in_209), .d_out(u_ca_out_209));
compressor_12_8 u_ca_12_8_210(.d_in(u_ca_in_210), .d_out(u_ca_out_210));
compressor_12_8 u_ca_12_8_211(.d_in(u_ca_in_211), .d_out(u_ca_out_211));
compressor_12_8 u_ca_12_8_212(.d_in(u_ca_in_212), .d_out(u_ca_out_212));
compressor_12_8 u_ca_12_8_213(.d_in(u_ca_in_213), .d_out(u_ca_out_213));
compressor_12_8 u_ca_12_8_214(.d_in(u_ca_in_214), .d_out(u_ca_out_214));
compressor_12_8 u_ca_12_8_215(.d_in(u_ca_in_215), .d_out(u_ca_out_215));
compressor_12_8 u_ca_12_8_216(.d_in(u_ca_in_216), .d_out(u_ca_out_216));
compressor_12_8 u_ca_12_8_217(.d_in(u_ca_in_217), .d_out(u_ca_out_217));
compressor_12_8 u_ca_12_8_218(.d_in(u_ca_in_218), .d_out(u_ca_out_218));
compressor_12_8 u_ca_12_8_219(.d_in(u_ca_in_219), .d_out(u_ca_out_219));
compressor_12_8 u_ca_12_8_220(.d_in(u_ca_in_220), .d_out(u_ca_out_220));
compressor_12_8 u_ca_12_8_221(.d_in(u_ca_in_221), .d_out(u_ca_out_221));
compressor_12_8 u_ca_12_8_222(.d_in(u_ca_in_222), .d_out(u_ca_out_222));
compressor_12_8 u_ca_12_8_223(.d_in(u_ca_in_223), .d_out(u_ca_out_223));
compressor_12_8 u_ca_12_8_224(.d_in(u_ca_in_224), .d_out(u_ca_out_224));
compressor_12_8 u_ca_12_8_225(.d_in(u_ca_in_225), .d_out(u_ca_out_225));
compressor_12_8 u_ca_12_8_226(.d_in(u_ca_in_226), .d_out(u_ca_out_226));
compressor_12_8 u_ca_12_8_227(.d_in(u_ca_in_227), .d_out(u_ca_out_227));
compressor_12_8 u_ca_12_8_228(.d_in(u_ca_in_228), .d_out(u_ca_out_228));
compressor_12_8 u_ca_12_8_229(.d_in(u_ca_in_229), .d_out(u_ca_out_229));
compressor_12_8 u_ca_12_8_230(.d_in(u_ca_in_230), .d_out(u_ca_out_230));
compressor_12_8 u_ca_12_8_231(.d_in(u_ca_in_231), .d_out(u_ca_out_231));
compressor_12_8 u_ca_12_8_232(.d_in(u_ca_in_232), .d_out(u_ca_out_232));
compressor_12_8 u_ca_12_8_233(.d_in(u_ca_in_233), .d_out(u_ca_out_233));
compressor_12_8 u_ca_12_8_234(.d_in(u_ca_in_234), .d_out(u_ca_out_234));
compressor_12_8 u_ca_12_8_235(.d_in(u_ca_in_235), .d_out(u_ca_out_235));
compressor_12_8 u_ca_12_8_236(.d_in(u_ca_in_236), .d_out(u_ca_out_236));
compressor_12_8 u_ca_12_8_237(.d_in(u_ca_in_237), .d_out(u_ca_out_237));
compressor_12_8 u_ca_12_8_238(.d_in(u_ca_in_238), .d_out(u_ca_out_238));
compressor_12_8 u_ca_12_8_239(.d_in(u_ca_in_239), .d_out(u_ca_out_239));
compressor_12_8 u_ca_12_8_240(.d_in(u_ca_in_240), .d_out(u_ca_out_240));
compressor_12_8 u_ca_12_8_241(.d_in(u_ca_in_241), .d_out(u_ca_out_241));
compressor_12_8 u_ca_12_8_242(.d_in(u_ca_in_242), .d_out(u_ca_out_242));
compressor_12_8 u_ca_12_8_243(.d_in(u_ca_in_243), .d_out(u_ca_out_243));
compressor_12_8 u_ca_12_8_244(.d_in(u_ca_in_244), .d_out(u_ca_out_244));
compressor_12_8 u_ca_12_8_245(.d_in(u_ca_in_245), .d_out(u_ca_out_245));
compressor_12_8 u_ca_12_8_246(.d_in(u_ca_in_246), .d_out(u_ca_out_246));
compressor_12_8 u_ca_12_8_247(.d_in(u_ca_in_247), .d_out(u_ca_out_247));
compressor_12_8 u_ca_12_8_248(.d_in(u_ca_in_248), .d_out(u_ca_out_248));
compressor_12_8 u_ca_12_8_249(.d_in(u_ca_in_249), .d_out(u_ca_out_249));
compressor_12_8 u_ca_12_8_250(.d_in(u_ca_in_250), .d_out(u_ca_out_250));
compressor_12_8 u_ca_12_8_251(.d_in(u_ca_in_251), .d_out(u_ca_out_251));
compressor_12_8 u_ca_12_8_252(.d_in(u_ca_in_252), .d_out(u_ca_out_252));
compressor_12_8 u_ca_12_8_253(.d_in(u_ca_in_253), .d_out(u_ca_out_253));
compressor_12_8 u_ca_12_8_254(.d_in(u_ca_in_254), .d_out(u_ca_out_254));
compressor_12_8 u_ca_12_8_255(.d_in(u_ca_in_255), .d_out(u_ca_out_255));
compressor_12_8 u_ca_12_8_256(.d_in(u_ca_in_256), .d_out(u_ca_out_256));
compressor_12_8 u_ca_12_8_257(.d_in(u_ca_in_257), .d_out(u_ca_out_257));
compressor_12_8 u_ca_12_8_258(.d_in(u_ca_in_258), .d_out(u_ca_out_258));
compressor_12_8 u_ca_12_8_259(.d_in(u_ca_in_259), .d_out(u_ca_out_259));
compressor_12_8 u_ca_12_8_260(.d_in(u_ca_in_260), .d_out(u_ca_out_260));
compressor_12_8 u_ca_12_8_261(.d_in(u_ca_in_261), .d_out(u_ca_out_261));
compressor_12_8 u_ca_12_8_262(.d_in(u_ca_in_262), .d_out(u_ca_out_262));
compressor_12_8 u_ca_12_8_263(.d_in(u_ca_in_263), .d_out(u_ca_out_263));
compressor_12_8 u_ca_12_8_264(.d_in(u_ca_in_264), .d_out(u_ca_out_264));
compressor_12_8 u_ca_12_8_265(.d_in(u_ca_in_265), .d_out(u_ca_out_265));
compressor_12_8 u_ca_12_8_266(.d_in(u_ca_in_266), .d_out(u_ca_out_266));
compressor_12_8 u_ca_12_8_267(.d_in(u_ca_in_267), .d_out(u_ca_out_267));
compressor_12_8 u_ca_12_8_268(.d_in(u_ca_in_268), .d_out(u_ca_out_268));
compressor_12_8 u_ca_12_8_269(.d_in(u_ca_in_269), .d_out(u_ca_out_269));
compressor_12_8 u_ca_12_8_270(.d_in(u_ca_in_270), .d_out(u_ca_out_270));
compressor_12_8 u_ca_12_8_271(.d_in(u_ca_in_271), .d_out(u_ca_out_271));
compressor_12_8 u_ca_12_8_272(.d_in(u_ca_in_272), .d_out(u_ca_out_272));
compressor_12_8 u_ca_12_8_273(.d_in(u_ca_in_273), .d_out(u_ca_out_273));
compressor_12_8 u_ca_12_8_274(.d_in(u_ca_in_274), .d_out(u_ca_out_274));
compressor_12_8 u_ca_12_8_275(.d_in(u_ca_in_275), .d_out(u_ca_out_275));
compressor_12_8 u_ca_12_8_276(.d_in(u_ca_in_276), .d_out(u_ca_out_276));
compressor_12_8 u_ca_12_8_277(.d_in(u_ca_in_277), .d_out(u_ca_out_277));
compressor_12_8 u_ca_12_8_278(.d_in(u_ca_in_278), .d_out(u_ca_out_278));
compressor_12_8 u_ca_12_8_279(.d_in(u_ca_in_279), .d_out(u_ca_out_279));
compressor_12_8 u_ca_12_8_280(.d_in(u_ca_in_280), .d_out(u_ca_out_280));
compressor_12_8 u_ca_12_8_281(.d_in(u_ca_in_281), .d_out(u_ca_out_281));
compressor_12_8 u_ca_12_8_282(.d_in(u_ca_in_282), .d_out(u_ca_out_282));
compressor_12_8 u_ca_12_8_283(.d_in(u_ca_in_283), .d_out(u_ca_out_283));
compressor_12_8 u_ca_12_8_284(.d_in(u_ca_in_284), .d_out(u_ca_out_284));
compressor_12_8 u_ca_12_8_285(.d_in(u_ca_in_285), .d_out(u_ca_out_285));
compressor_12_8 u_ca_12_8_286(.d_in(u_ca_in_286), .d_out(u_ca_out_286));
compressor_12_8 u_ca_12_8_287(.d_in(u_ca_in_287), .d_out(u_ca_out_287));
compressor_12_8 u_ca_12_8_288(.d_in(u_ca_in_288), .d_out(u_ca_out_288));
compressor_12_8 u_ca_12_8_289(.d_in(u_ca_in_289), .d_out(u_ca_out_289));
compressor_12_8 u_ca_12_8_290(.d_in(u_ca_in_290), .d_out(u_ca_out_290));
compressor_12_8 u_ca_12_8_291(.d_in(u_ca_in_291), .d_out(u_ca_out_291));
compressor_12_8 u_ca_12_8_292(.d_in(u_ca_in_292), .d_out(u_ca_out_292));
compressor_12_8 u_ca_12_8_293(.d_in(u_ca_in_293), .d_out(u_ca_out_293));
compressor_12_8 u_ca_12_8_294(.d_in(u_ca_in_294), .d_out(u_ca_out_294));
compressor_12_8 u_ca_12_8_295(.d_in(u_ca_in_295), .d_out(u_ca_out_295));
compressor_12_8 u_ca_12_8_296(.d_in(u_ca_in_296), .d_out(u_ca_out_296));
compressor_12_8 u_ca_12_8_297(.d_in(u_ca_in_297), .d_out(u_ca_out_297));
compressor_12_8 u_ca_12_8_298(.d_in(u_ca_in_298), .d_out(u_ca_out_298));
compressor_12_8 u_ca_12_8_299(.d_in(u_ca_in_299), .d_out(u_ca_out_299));
compressor_12_8 u_ca_12_8_300(.d_in(u_ca_in_300), .d_out(u_ca_out_300));
compressor_12_8 u_ca_12_8_301(.d_in(u_ca_in_301), .d_out(u_ca_out_301));
compressor_12_8 u_ca_12_8_302(.d_in(u_ca_in_302), .d_out(u_ca_out_302));
compressor_12_8 u_ca_12_8_303(.d_in(u_ca_in_303), .d_out(u_ca_out_303));
compressor_12_8 u_ca_12_8_304(.d_in(u_ca_in_304), .d_out(u_ca_out_304));
compressor_12_8 u_ca_12_8_305(.d_in(u_ca_in_305), .d_out(u_ca_out_305));
compressor_12_8 u_ca_12_8_306(.d_in(u_ca_in_306), .d_out(u_ca_out_306));
compressor_12_8 u_ca_12_8_307(.d_in(u_ca_in_307), .d_out(u_ca_out_307));
compressor_12_8 u_ca_12_8_308(.d_in(u_ca_in_308), .d_out(u_ca_out_308));
compressor_12_8 u_ca_12_8_309(.d_in(u_ca_in_309), .d_out(u_ca_out_309));
compressor_12_8 u_ca_12_8_310(.d_in(u_ca_in_310), .d_out(u_ca_out_310));
compressor_12_8 u_ca_12_8_311(.d_in(u_ca_in_311), .d_out(u_ca_out_311));
compressor_12_8 u_ca_12_8_312(.d_in(u_ca_in_312), .d_out(u_ca_out_312));
compressor_12_8 u_ca_12_8_313(.d_in(u_ca_in_313), .d_out(u_ca_out_313));
compressor_12_8 u_ca_12_8_314(.d_in(u_ca_in_314), .d_out(u_ca_out_314));
compressor_12_8 u_ca_12_8_315(.d_in(u_ca_in_315), .d_out(u_ca_out_315));
compressor_12_8 u_ca_12_8_316(.d_in(u_ca_in_316), .d_out(u_ca_out_316));
compressor_12_8 u_ca_12_8_317(.d_in(u_ca_in_317), .d_out(u_ca_out_317));
compressor_12_8 u_ca_12_8_318(.d_in(u_ca_in_318), .d_out(u_ca_out_318));
compressor_12_8 u_ca_12_8_319(.d_in(u_ca_in_319), .d_out(u_ca_out_319));
compressor_12_8 u_ca_12_8_320(.d_in(u_ca_in_320), .d_out(u_ca_out_320));
compressor_12_8 u_ca_12_8_321(.d_in(u_ca_in_321), .d_out(u_ca_out_321));
compressor_12_8 u_ca_12_8_322(.d_in(u_ca_in_322), .d_out(u_ca_out_322));
compressor_12_8 u_ca_12_8_323(.d_in(u_ca_in_323), .d_out(u_ca_out_323));
compressor_12_8 u_ca_12_8_324(.d_in(u_ca_in_324), .d_out(u_ca_out_324));
compressor_12_8 u_ca_12_8_325(.d_in(u_ca_in_325), .d_out(u_ca_out_325));
compressor_12_8 u_ca_12_8_326(.d_in(u_ca_in_326), .d_out(u_ca_out_326));
compressor_12_8 u_ca_12_8_327(.d_in(u_ca_in_327), .d_out(u_ca_out_327));
compressor_12_8 u_ca_12_8_328(.d_in(u_ca_in_328), .d_out(u_ca_out_328));
compressor_12_8 u_ca_12_8_329(.d_in(u_ca_in_329), .d_out(u_ca_out_329));
compressor_12_8 u_ca_12_8_330(.d_in(u_ca_in_330), .d_out(u_ca_out_330));
compressor_12_8 u_ca_12_8_331(.d_in(u_ca_in_331), .d_out(u_ca_out_331));
compressor_12_8 u_ca_12_8_332(.d_in(u_ca_in_332), .d_out(u_ca_out_332));
compressor_12_8 u_ca_12_8_333(.d_in(u_ca_in_333), .d_out(u_ca_out_333));
compressor_12_8 u_ca_12_8_334(.d_in(u_ca_in_334), .d_out(u_ca_out_334));
compressor_12_8 u_ca_12_8_335(.d_in(u_ca_in_335), .d_out(u_ca_out_335));
compressor_12_8 u_ca_12_8_336(.d_in(u_ca_in_336), .d_out(u_ca_out_336));
compressor_12_8 u_ca_12_8_337(.d_in(u_ca_in_337), .d_out(u_ca_out_337));
compressor_12_8 u_ca_12_8_338(.d_in(u_ca_in_338), .d_out(u_ca_out_338));
compressor_12_8 u_ca_12_8_339(.d_in(u_ca_in_339), .d_out(u_ca_out_339));
compressor_12_8 u_ca_12_8_340(.d_in(u_ca_in_340), .d_out(u_ca_out_340));
compressor_12_8 u_ca_12_8_341(.d_in(u_ca_in_341), .d_out(u_ca_out_341));
compressor_12_8 u_ca_12_8_342(.d_in(u_ca_in_342), .d_out(u_ca_out_342));
compressor_12_8 u_ca_12_8_343(.d_in(u_ca_in_343), .d_out(u_ca_out_343));
compressor_12_8 u_ca_12_8_344(.d_in(u_ca_in_344), .d_out(u_ca_out_344));
compressor_12_8 u_ca_12_8_345(.d_in(u_ca_in_345), .d_out(u_ca_out_345));
compressor_12_8 u_ca_12_8_346(.d_in(u_ca_in_346), .d_out(u_ca_out_346));
compressor_12_8 u_ca_12_8_347(.d_in(u_ca_in_347), .d_out(u_ca_out_347));
compressor_12_8 u_ca_12_8_348(.d_in(u_ca_in_348), .d_out(u_ca_out_348));
compressor_12_8 u_ca_12_8_349(.d_in(u_ca_in_349), .d_out(u_ca_out_349));
compressor_12_8 u_ca_12_8_350(.d_in(u_ca_in_350), .d_out(u_ca_out_350));
compressor_12_8 u_ca_12_8_351(.d_in(u_ca_in_351), .d_out(u_ca_out_351));
compressor_12_8 u_ca_12_8_352(.d_in(u_ca_in_352), .d_out(u_ca_out_352));
compressor_12_8 u_ca_12_8_353(.d_in(u_ca_in_353), .d_out(u_ca_out_353));
compressor_12_8 u_ca_12_8_354(.d_in(u_ca_in_354), .d_out(u_ca_out_354));
compressor_12_8 u_ca_12_8_355(.d_in(u_ca_in_355), .d_out(u_ca_out_355));
compressor_12_8 u_ca_12_8_356(.d_in(u_ca_in_356), .d_out(u_ca_out_356));
compressor_12_8 u_ca_12_8_357(.d_in(u_ca_in_357), .d_out(u_ca_out_357));
compressor_12_8 u_ca_12_8_358(.d_in(u_ca_in_358), .d_out(u_ca_out_358));
compressor_12_8 u_ca_12_8_359(.d_in(u_ca_in_359), .d_out(u_ca_out_359));
compressor_12_8 u_ca_12_8_360(.d_in(u_ca_in_360), .d_out(u_ca_out_360));
compressor_12_8 u_ca_12_8_361(.d_in(u_ca_in_361), .d_out(u_ca_out_361));
compressor_12_8 u_ca_12_8_362(.d_in(u_ca_in_362), .d_out(u_ca_out_362));
compressor_12_8 u_ca_12_8_363(.d_in(u_ca_in_363), .d_out(u_ca_out_363));
compressor_12_8 u_ca_12_8_364(.d_in(u_ca_in_364), .d_out(u_ca_out_364));
compressor_12_8 u_ca_12_8_365(.d_in(u_ca_in_365), .d_out(u_ca_out_365));
compressor_12_8 u_ca_12_8_366(.d_in(u_ca_in_366), .d_out(u_ca_out_366));
compressor_12_8 u_ca_12_8_367(.d_in(u_ca_in_367), .d_out(u_ca_out_367));
compressor_12_8 u_ca_12_8_368(.d_in(u_ca_in_368), .d_out(u_ca_out_368));
compressor_12_8 u_ca_12_8_369(.d_in(u_ca_in_369), .d_out(u_ca_out_369));
compressor_12_8 u_ca_12_8_370(.d_in(u_ca_in_370), .d_out(u_ca_out_370));
compressor_12_8 u_ca_12_8_371(.d_in(u_ca_in_371), .d_out(u_ca_out_371));
compressor_12_8 u_ca_12_8_372(.d_in(u_ca_in_372), .d_out(u_ca_out_372));
compressor_12_8 u_ca_12_8_373(.d_in(u_ca_in_373), .d_out(u_ca_out_373));
compressor_12_8 u_ca_12_8_374(.d_in(u_ca_in_374), .d_out(u_ca_out_374));
compressor_12_8 u_ca_12_8_375(.d_in(u_ca_in_375), .d_out(u_ca_out_375));
compressor_12_8 u_ca_12_8_376(.d_in(u_ca_in_376), .d_out(u_ca_out_376));
compressor_12_8 u_ca_12_8_377(.d_in(u_ca_in_377), .d_out(u_ca_out_377));
compressor_12_8 u_ca_12_8_378(.d_in(u_ca_in_378), .d_out(u_ca_out_378));
compressor_12_8 u_ca_12_8_379(.d_in(u_ca_in_379), .d_out(u_ca_out_379));
compressor_12_8 u_ca_12_8_380(.d_in(u_ca_in_380), .d_out(u_ca_out_380));
compressor_12_8 u_ca_12_8_381(.d_in(u_ca_in_381), .d_out(u_ca_out_381));
compressor_12_8 u_ca_12_8_382(.d_in(u_ca_in_382), .d_out(u_ca_out_382));
compressor_12_8 u_ca_12_8_383(.d_in(u_ca_in_383), .d_out(u_ca_out_383));
compressor_12_8 u_ca_12_8_384(.d_in(u_ca_in_384), .d_out(u_ca_out_384));
compressor_12_8 u_ca_12_8_385(.d_in(u_ca_in_385), .d_out(u_ca_out_385));
compressor_12_8 u_ca_12_8_386(.d_in(u_ca_in_386), .d_out(u_ca_out_386));
compressor_12_8 u_ca_12_8_387(.d_in(u_ca_in_387), .d_out(u_ca_out_387));
compressor_12_8 u_ca_12_8_388(.d_in(u_ca_in_388), .d_out(u_ca_out_388));
compressor_12_8 u_ca_12_8_389(.d_in(u_ca_in_389), .d_out(u_ca_out_389));
compressor_12_8 u_ca_12_8_390(.d_in(u_ca_in_390), .d_out(u_ca_out_390));
compressor_12_8 u_ca_12_8_391(.d_in(u_ca_in_391), .d_out(u_ca_out_391));
compressor_12_8 u_ca_12_8_392(.d_in(u_ca_in_392), .d_out(u_ca_out_392));
compressor_12_8 u_ca_12_8_393(.d_in(u_ca_in_393), .d_out(u_ca_out_393));
compressor_12_8 u_ca_12_8_394(.d_in(u_ca_in_394), .d_out(u_ca_out_394));
compressor_12_8 u_ca_12_8_395(.d_in(u_ca_in_395), .d_out(u_ca_out_395));
compressor_12_8 u_ca_12_8_396(.d_in(u_ca_in_396), .d_out(u_ca_out_396));
compressor_12_8 u_ca_12_8_397(.d_in(u_ca_in_397), .d_out(u_ca_out_397));
compressor_12_8 u_ca_12_8_398(.d_in(u_ca_in_398), .d_out(u_ca_out_398));
compressor_12_8 u_ca_12_8_399(.d_in(u_ca_in_399), .d_out(u_ca_out_399));
compressor_12_8 u_ca_12_8_400(.d_in(u_ca_in_400), .d_out(u_ca_out_400));
compressor_12_8 u_ca_12_8_401(.d_in(u_ca_in_401), .d_out(u_ca_out_401));
compressor_12_8 u_ca_12_8_402(.d_in(u_ca_in_402), .d_out(u_ca_out_402));
compressor_12_8 u_ca_12_8_403(.d_in(u_ca_in_403), .d_out(u_ca_out_403));
compressor_12_8 u_ca_12_8_404(.d_in(u_ca_in_404), .d_out(u_ca_out_404));
compressor_12_8 u_ca_12_8_405(.d_in(u_ca_in_405), .d_out(u_ca_out_405));
compressor_12_8 u_ca_12_8_406(.d_in(u_ca_in_406), .d_out(u_ca_out_406));
compressor_12_8 u_ca_12_8_407(.d_in(u_ca_in_407), .d_out(u_ca_out_407));
compressor_12_8 u_ca_12_8_408(.d_in(u_ca_in_408), .d_out(u_ca_out_408));
compressor_12_8 u_ca_12_8_409(.d_in(u_ca_in_409), .d_out(u_ca_out_409));
compressor_12_8 u_ca_12_8_410(.d_in(u_ca_in_410), .d_out(u_ca_out_410));
compressor_12_8 u_ca_12_8_411(.d_in(u_ca_in_411), .d_out(u_ca_out_411));
compressor_12_8 u_ca_12_8_412(.d_in(u_ca_in_412), .d_out(u_ca_out_412));
compressor_12_8 u_ca_12_8_413(.d_in(u_ca_in_413), .d_out(u_ca_out_413));
compressor_12_8 u_ca_12_8_414(.d_in(u_ca_in_414), .d_out(u_ca_out_414));
compressor_12_8 u_ca_12_8_415(.d_in(u_ca_in_415), .d_out(u_ca_out_415));
compressor_12_8 u_ca_12_8_416(.d_in(u_ca_in_416), .d_out(u_ca_out_416));
compressor_12_8 u_ca_12_8_417(.d_in(u_ca_in_417), .d_out(u_ca_out_417));
compressor_12_8 u_ca_12_8_418(.d_in(u_ca_in_418), .d_out(u_ca_out_418));
compressor_12_8 u_ca_12_8_419(.d_in(u_ca_in_419), .d_out(u_ca_out_419));
compressor_12_8 u_ca_12_8_420(.d_in(u_ca_in_420), .d_out(u_ca_out_420));
compressor_12_8 u_ca_12_8_421(.d_in(u_ca_in_421), .d_out(u_ca_out_421));
compressor_12_8 u_ca_12_8_422(.d_in(u_ca_in_422), .d_out(u_ca_out_422));
compressor_12_8 u_ca_12_8_423(.d_in(u_ca_in_423), .d_out(u_ca_out_423));
compressor_12_8 u_ca_12_8_424(.d_in(u_ca_in_424), .d_out(u_ca_out_424));
compressor_12_8 u_ca_12_8_425(.d_in(u_ca_in_425), .d_out(u_ca_out_425));
compressor_12_8 u_ca_12_8_426(.d_in(u_ca_in_426), .d_out(u_ca_out_426));
compressor_12_8 u_ca_12_8_427(.d_in(u_ca_in_427), .d_out(u_ca_out_427));
compressor_12_8 u_ca_12_8_428(.d_in(u_ca_in_428), .d_out(u_ca_out_428));
compressor_12_8 u_ca_12_8_429(.d_in(u_ca_in_429), .d_out(u_ca_out_429));
compressor_12_8 u_ca_12_8_430(.d_in(u_ca_in_430), .d_out(u_ca_out_430));
compressor_12_8 u_ca_12_8_431(.d_in(u_ca_in_431), .d_out(u_ca_out_431));
compressor_12_8 u_ca_12_8_432(.d_in(u_ca_in_432), .d_out(u_ca_out_432));
compressor_12_8 u_ca_12_8_433(.d_in(u_ca_in_433), .d_out(u_ca_out_433));
compressor_12_8 u_ca_12_8_434(.d_in(u_ca_in_434), .d_out(u_ca_out_434));
compressor_12_8 u_ca_12_8_435(.d_in(u_ca_in_435), .d_out(u_ca_out_435));
compressor_12_8 u_ca_12_8_436(.d_in(u_ca_in_436), .d_out(u_ca_out_436));
compressor_12_8 u_ca_12_8_437(.d_in(u_ca_in_437), .d_out(u_ca_out_437));
compressor_12_8 u_ca_12_8_438(.d_in(u_ca_in_438), .d_out(u_ca_out_438));
compressor_12_8 u_ca_12_8_439(.d_in(u_ca_in_439), .d_out(u_ca_out_439));
compressor_12_8 u_ca_12_8_440(.d_in(u_ca_in_440), .d_out(u_ca_out_440));
compressor_12_8 u_ca_12_8_441(.d_in(u_ca_in_441), .d_out(u_ca_out_441));
compressor_12_8 u_ca_12_8_442(.d_in(u_ca_in_442), .d_out(u_ca_out_442));
compressor_12_8 u_ca_12_8_443(.d_in(u_ca_in_443), .d_out(u_ca_out_443));
compressor_12_8 u_ca_12_8_444(.d_in(u_ca_in_444), .d_out(u_ca_out_444));
compressor_12_8 u_ca_12_8_445(.d_in(u_ca_in_445), .d_out(u_ca_out_445));
compressor_12_8 u_ca_12_8_446(.d_in(u_ca_in_446), .d_out(u_ca_out_446));
compressor_12_8 u_ca_12_8_447(.d_in(u_ca_in_447), .d_out(u_ca_out_447));
compressor_12_8 u_ca_12_8_448(.d_in(u_ca_in_448), .d_out(u_ca_out_448));
compressor_12_8 u_ca_12_8_449(.d_in(u_ca_in_449), .d_out(u_ca_out_449));
compressor_12_8 u_ca_12_8_450(.d_in(u_ca_in_450), .d_out(u_ca_out_450));
compressor_12_8 u_ca_12_8_451(.d_in(u_ca_in_451), .d_out(u_ca_out_451));
compressor_12_8 u_ca_12_8_452(.d_in(u_ca_in_452), .d_out(u_ca_out_452));
compressor_12_8 u_ca_12_8_453(.d_in(u_ca_in_453), .d_out(u_ca_out_453));
compressor_12_8 u_ca_12_8_454(.d_in(u_ca_in_454), .d_out(u_ca_out_454));
compressor_12_8 u_ca_12_8_455(.d_in(u_ca_in_455), .d_out(u_ca_out_455));
compressor_12_8 u_ca_12_8_456(.d_in(u_ca_in_456), .d_out(u_ca_out_456));
compressor_12_8 u_ca_12_8_457(.d_in(u_ca_in_457), .d_out(u_ca_out_457));
compressor_12_8 u_ca_12_8_458(.d_in(u_ca_in_458), .d_out(u_ca_out_458));
compressor_12_8 u_ca_12_8_459(.d_in(u_ca_in_459), .d_out(u_ca_out_459));
compressor_12_8 u_ca_12_8_460(.d_in(u_ca_in_460), .d_out(u_ca_out_460));
compressor_12_8 u_ca_12_8_461(.d_in(u_ca_in_461), .d_out(u_ca_out_461));
compressor_12_8 u_ca_12_8_462(.d_in(u_ca_in_462), .d_out(u_ca_out_462));
compressor_12_8 u_ca_12_8_463(.d_in(u_ca_in_463), .d_out(u_ca_out_463));
compressor_12_8 u_ca_12_8_464(.d_in(u_ca_in_464), .d_out(u_ca_out_464));
compressor_12_8 u_ca_12_8_465(.d_in(u_ca_in_465), .d_out(u_ca_out_465));
compressor_12_8 u_ca_12_8_466(.d_in(u_ca_in_466), .d_out(u_ca_out_466));
compressor_12_8 u_ca_12_8_467(.d_in(u_ca_in_467), .d_out(u_ca_out_467));
compressor_12_8 u_ca_12_8_468(.d_in(u_ca_in_468), .d_out(u_ca_out_468));
compressor_12_8 u_ca_12_8_469(.d_in(u_ca_in_469), .d_out(u_ca_out_469));
compressor_12_8 u_ca_12_8_470(.d_in(u_ca_in_470), .d_out(u_ca_out_470));
compressor_12_8 u_ca_12_8_471(.d_in(u_ca_in_471), .d_out(u_ca_out_471));
compressor_12_8 u_ca_12_8_472(.d_in(u_ca_in_472), .d_out(u_ca_out_472));
compressor_12_8 u_ca_12_8_473(.d_in(u_ca_in_473), .d_out(u_ca_out_473));
compressor_12_8 u_ca_12_8_474(.d_in(u_ca_in_474), .d_out(u_ca_out_474));
compressor_12_8 u_ca_12_8_475(.d_in(u_ca_in_475), .d_out(u_ca_out_475));
compressor_12_8 u_ca_12_8_476(.d_in(u_ca_in_476), .d_out(u_ca_out_476));
compressor_12_8 u_ca_12_8_477(.d_in(u_ca_in_477), .d_out(u_ca_out_477));
compressor_12_8 u_ca_12_8_478(.d_in(u_ca_in_478), .d_out(u_ca_out_478));
compressor_12_8 u_ca_12_8_479(.d_in(u_ca_in_479), .d_out(u_ca_out_479));
compressor_12_8 u_ca_12_8_480(.d_in(u_ca_in_480), .d_out(u_ca_out_480));
compressor_12_8 u_ca_12_8_481(.d_in(u_ca_in_481), .d_out(u_ca_out_481));
compressor_12_8 u_ca_12_8_482(.d_in(u_ca_in_482), .d_out(u_ca_out_482));
compressor_12_8 u_ca_12_8_483(.d_in(u_ca_in_483), .d_out(u_ca_out_483));
compressor_12_8 u_ca_12_8_484(.d_in(u_ca_in_484), .d_out(u_ca_out_484));
compressor_12_8 u_ca_12_8_485(.d_in(u_ca_in_485), .d_out(u_ca_out_485));
compressor_12_8 u_ca_12_8_486(.d_in(u_ca_in_486), .d_out(u_ca_out_486));
compressor_12_8 u_ca_12_8_487(.d_in(u_ca_in_487), .d_out(u_ca_out_487));
compressor_12_8 u_ca_12_8_488(.d_in(u_ca_in_488), .d_out(u_ca_out_488));
compressor_12_8 u_ca_12_8_489(.d_in(u_ca_in_489), .d_out(u_ca_out_489));
compressor_12_8 u_ca_12_8_490(.d_in(u_ca_in_490), .d_out(u_ca_out_490));
compressor_12_8 u_ca_12_8_491(.d_in(u_ca_in_491), .d_out(u_ca_out_491));
compressor_12_8 u_ca_12_8_492(.d_in(u_ca_in_492), .d_out(u_ca_out_492));
compressor_12_8 u_ca_12_8_493(.d_in(u_ca_in_493), .d_out(u_ca_out_493));
compressor_12_8 u_ca_12_8_494(.d_in(u_ca_in_494), .d_out(u_ca_out_494));
compressor_12_8 u_ca_12_8_495(.d_in(u_ca_in_495), .d_out(u_ca_out_495));
compressor_12_8 u_ca_12_8_496(.d_in(u_ca_in_496), .d_out(u_ca_out_496));
compressor_12_8 u_ca_12_8_497(.d_in(u_ca_in_497), .d_out(u_ca_out_497));
compressor_12_8 u_ca_12_8_498(.d_in(u_ca_in_498), .d_out(u_ca_out_498));
compressor_12_8 u_ca_12_8_499(.d_in(u_ca_in_499), .d_out(u_ca_out_499));
compressor_12_8 u_ca_12_8_500(.d_in(u_ca_in_500), .d_out(u_ca_out_500));
compressor_12_8 u_ca_12_8_501(.d_in(u_ca_in_501), .d_out(u_ca_out_501));
compressor_12_8 u_ca_12_8_502(.d_in(u_ca_in_502), .d_out(u_ca_out_502));
compressor_12_8 u_ca_12_8_503(.d_in(u_ca_in_503), .d_out(u_ca_out_503));
compressor_12_8 u_ca_12_8_504(.d_in(u_ca_in_504), .d_out(u_ca_out_504));
compressor_12_8 u_ca_12_8_505(.d_in(u_ca_in_505), .d_out(u_ca_out_505));
compressor_12_8 u_ca_12_8_506(.d_in(u_ca_in_506), .d_out(u_ca_out_506));
compressor_12_8 u_ca_12_8_507(.d_in(u_ca_in_507), .d_out(u_ca_out_507));
compressor_12_8 u_ca_12_8_508(.d_in(u_ca_in_508), .d_out(u_ca_out_508));
compressor_12_8 u_ca_12_8_509(.d_in(u_ca_in_509), .d_out(u_ca_out_509));
compressor_12_8 u_ca_12_8_510(.d_in(u_ca_in_510), .d_out(u_ca_out_510));
compressor_12_8 u_ca_12_8_511(.d_in(u_ca_in_511), .d_out(u_ca_out_511));
compressor_12_8 u_ca_12_8_512(.d_in(u_ca_in_512), .d_out(u_ca_out_512));
compressor_12_8 u_ca_12_8_513(.d_in(u_ca_in_513), .d_out(u_ca_out_513));
compressor_12_8 u_ca_12_8_514(.d_in(u_ca_in_514), .d_out(u_ca_out_514));
compressor_12_8 u_ca_12_8_515(.d_in(u_ca_in_515), .d_out(u_ca_out_515));
compressor_12_8 u_ca_12_8_516(.d_in(u_ca_in_516), .d_out(u_ca_out_516));
compressor_12_8 u_ca_12_8_517(.d_in(u_ca_in_517), .d_out(u_ca_out_517));
compressor_12_8 u_ca_12_8_518(.d_in(u_ca_in_518), .d_out(u_ca_out_518));
compressor_12_8 u_ca_12_8_519(.d_in(u_ca_in_519), .d_out(u_ca_out_519));
compressor_12_8 u_ca_12_8_520(.d_in(u_ca_in_520), .d_out(u_ca_out_520));
compressor_12_8 u_ca_12_8_521(.d_in(u_ca_in_521), .d_out(u_ca_out_521));
compressor_12_8 u_ca_12_8_522(.d_in(u_ca_in_522), .d_out(u_ca_out_522));
compressor_12_8 u_ca_12_8_523(.d_in(u_ca_in_523), .d_out(u_ca_out_523));
compressor_12_8 u_ca_12_8_524(.d_in(u_ca_in_524), .d_out(u_ca_out_524));
compressor_12_8 u_ca_12_8_525(.d_in(u_ca_in_525), .d_out(u_ca_out_525));
compressor_12_8 u_ca_12_8_526(.d_in(u_ca_in_526), .d_out(u_ca_out_526));
compressor_12_8 u_ca_12_8_527(.d_in(u_ca_in_527), .d_out(u_ca_out_527));
compressor_12_8 u_ca_12_8_528(.d_in(u_ca_in_528), .d_out(u_ca_out_528));
compressor_12_8 u_ca_12_8_529(.d_in(u_ca_in_529), .d_out(u_ca_out_529));
compressor_12_8 u_ca_12_8_530(.d_in(u_ca_in_530), .d_out(u_ca_out_530));
compressor_12_8 u_ca_12_8_531(.d_in(u_ca_in_531), .d_out(u_ca_out_531));
compressor_12_8 u_ca_12_8_532(.d_in(u_ca_in_532), .d_out(u_ca_out_532));
compressor_12_8 u_ca_12_8_533(.d_in(u_ca_in_533), .d_out(u_ca_out_533));
compressor_12_8 u_ca_12_8_534(.d_in(u_ca_in_534), .d_out(u_ca_out_534));
compressor_12_8 u_ca_12_8_535(.d_in(u_ca_in_535), .d_out(u_ca_out_535));
compressor_12_8 u_ca_12_8_536(.d_in(u_ca_in_536), .d_out(u_ca_out_536));
compressor_12_8 u_ca_12_8_537(.d_in(u_ca_in_537), .d_out(u_ca_out_537));
compressor_12_8 u_ca_12_8_538(.d_in(u_ca_in_538), .d_out(u_ca_out_538));
compressor_12_8 u_ca_12_8_539(.d_in(u_ca_in_539), .d_out(u_ca_out_539));
compressor_12_8 u_ca_12_8_540(.d_in(u_ca_in_540), .d_out(u_ca_out_540));
compressor_12_8 u_ca_12_8_541(.d_in(u_ca_in_541), .d_out(u_ca_out_541));
compressor_12_8 u_ca_12_8_542(.d_in(u_ca_in_542), .d_out(u_ca_out_542));
compressor_12_8 u_ca_12_8_543(.d_in(u_ca_in_543), .d_out(u_ca_out_543));
compressor_12_8 u_ca_12_8_544(.d_in(u_ca_in_544), .d_out(u_ca_out_544));
compressor_12_8 u_ca_12_8_545(.d_in(u_ca_in_545), .d_out(u_ca_out_545));
compressor_12_8 u_ca_12_8_546(.d_in(u_ca_in_546), .d_out(u_ca_out_546));
compressor_12_8 u_ca_12_8_547(.d_in(u_ca_in_547), .d_out(u_ca_out_547));
compressor_12_8 u_ca_12_8_548(.d_in(u_ca_in_548), .d_out(u_ca_out_548));
compressor_12_8 u_ca_12_8_549(.d_in(u_ca_in_549), .d_out(u_ca_out_549));
compressor_12_8 u_ca_12_8_550(.d_in(u_ca_in_550), .d_out(u_ca_out_550));
compressor_12_8 u_ca_12_8_551(.d_in(u_ca_in_551), .d_out(u_ca_out_551));
compressor_12_8 u_ca_12_8_552(.d_in(u_ca_in_552), .d_out(u_ca_out_552));
compressor_12_8 u_ca_12_8_553(.d_in(u_ca_in_553), .d_out(u_ca_out_553));
compressor_12_8 u_ca_12_8_554(.d_in(u_ca_in_554), .d_out(u_ca_out_554));
compressor_12_8 u_ca_12_8_555(.d_in(u_ca_in_555), .d_out(u_ca_out_555));
compressor_12_8 u_ca_12_8_556(.d_in(u_ca_in_556), .d_out(u_ca_out_556));
compressor_12_8 u_ca_12_8_557(.d_in(u_ca_in_557), .d_out(u_ca_out_557));
compressor_12_8 u_ca_12_8_558(.d_in(u_ca_in_558), .d_out(u_ca_out_558));
compressor_12_8 u_ca_12_8_559(.d_in(u_ca_in_559), .d_out(u_ca_out_559));
compressor_12_8 u_ca_12_8_560(.d_in(u_ca_in_560), .d_out(u_ca_out_560));
compressor_12_8 u_ca_12_8_561(.d_in(u_ca_in_561), .d_out(u_ca_out_561));
compressor_12_8 u_ca_12_8_562(.d_in(u_ca_in_562), .d_out(u_ca_out_562));
compressor_12_8 u_ca_12_8_563(.d_in(u_ca_in_563), .d_out(u_ca_out_563));
compressor_12_8 u_ca_12_8_564(.d_in(u_ca_in_564), .d_out(u_ca_out_564));
compressor_12_8 u_ca_12_8_565(.d_in(u_ca_in_565), .d_out(u_ca_out_565));
compressor_12_8 u_ca_12_8_566(.d_in(u_ca_in_566), .d_out(u_ca_out_566));
compressor_12_8 u_ca_12_8_567(.d_in(u_ca_in_567), .d_out(u_ca_out_567));
compressor_12_8 u_ca_12_8_568(.d_in(u_ca_in_568), .d_out(u_ca_out_568));
compressor_12_8 u_ca_12_8_569(.d_in(u_ca_in_569), .d_out(u_ca_out_569));
compressor_12_8 u_ca_12_8_570(.d_in(u_ca_in_570), .d_out(u_ca_out_570));
compressor_12_8 u_ca_12_8_571(.d_in(u_ca_in_571), .d_out(u_ca_out_571));
compressor_12_8 u_ca_12_8_572(.d_in(u_ca_in_572), .d_out(u_ca_out_572));
compressor_12_8 u_ca_12_8_573(.d_in(u_ca_in_573), .d_out(u_ca_out_573));
compressor_12_8 u_ca_12_8_574(.d_in(u_ca_in_574), .d_out(u_ca_out_574));
compressor_12_8 u_ca_12_8_575(.d_in(u_ca_in_575), .d_out(u_ca_out_575));
compressor_12_8 u_ca_12_8_576(.d_in(u_ca_in_576), .d_out(u_ca_out_576));
compressor_12_8 u_ca_12_8_577(.d_in(u_ca_in_577), .d_out(u_ca_out_577));
compressor_12_8 u_ca_12_8_578(.d_in(u_ca_in_578), .d_out(u_ca_out_578));
compressor_12_8 u_ca_12_8_579(.d_in(u_ca_in_579), .d_out(u_ca_out_579));
compressor_12_8 u_ca_12_8_580(.d_in(u_ca_in_580), .d_out(u_ca_out_580));
compressor_12_8 u_ca_12_8_581(.d_in(u_ca_in_581), .d_out(u_ca_out_581));
compressor_12_8 u_ca_12_8_582(.d_in(u_ca_in_582), .d_out(u_ca_out_582));
compressor_12_8 u_ca_12_8_583(.d_in(u_ca_in_583), .d_out(u_ca_out_583));
compressor_12_8 u_ca_12_8_584(.d_in(u_ca_in_584), .d_out(u_ca_out_584));
compressor_12_8 u_ca_12_8_585(.d_in(u_ca_in_585), .d_out(u_ca_out_585));
compressor_12_8 u_ca_12_8_586(.d_in(u_ca_in_586), .d_out(u_ca_out_586));
compressor_12_8 u_ca_12_8_587(.d_in(u_ca_in_587), .d_out(u_ca_out_587));
compressor_12_8 u_ca_12_8_588(.d_in(u_ca_in_588), .d_out(u_ca_out_588));
compressor_12_8 u_ca_12_8_589(.d_in(u_ca_in_589), .d_out(u_ca_out_589));
compressor_12_8 u_ca_12_8_590(.d_in(u_ca_in_590), .d_out(u_ca_out_590));
compressor_12_8 u_ca_12_8_591(.d_in(u_ca_in_591), .d_out(u_ca_out_591));
compressor_12_8 u_ca_12_8_592(.d_in(u_ca_in_592), .d_out(u_ca_out_592));
compressor_12_8 u_ca_12_8_593(.d_in(u_ca_in_593), .d_out(u_ca_out_593));
compressor_12_8 u_ca_12_8_594(.d_in(u_ca_in_594), .d_out(u_ca_out_594));
compressor_12_8 u_ca_12_8_595(.d_in(u_ca_in_595), .d_out(u_ca_out_595));
compressor_12_8 u_ca_12_8_596(.d_in(u_ca_in_596), .d_out(u_ca_out_596));
compressor_12_8 u_ca_12_8_597(.d_in(u_ca_in_597), .d_out(u_ca_out_597));
compressor_12_8 u_ca_12_8_598(.d_in(u_ca_in_598), .d_out(u_ca_out_598));
compressor_12_8 u_ca_12_8_599(.d_in(u_ca_in_599), .d_out(u_ca_out_599));
compressor_12_8 u_ca_12_8_600(.d_in(u_ca_in_600), .d_out(u_ca_out_600));
compressor_12_8 u_ca_12_8_601(.d_in(u_ca_in_601), .d_out(u_ca_out_601));
compressor_12_8 u_ca_12_8_602(.d_in(u_ca_in_602), .d_out(u_ca_out_602));
compressor_12_8 u_ca_12_8_603(.d_in(u_ca_in_603), .d_out(u_ca_out_603));
compressor_12_8 u_ca_12_8_604(.d_in(u_ca_in_604), .d_out(u_ca_out_604));
compressor_12_8 u_ca_12_8_605(.d_in(u_ca_in_605), .d_out(u_ca_out_605));
compressor_12_8 u_ca_12_8_606(.d_in(u_ca_in_606), .d_out(u_ca_out_606));
compressor_12_8 u_ca_12_8_607(.d_in(u_ca_in_607), .d_out(u_ca_out_607));
compressor_12_8 u_ca_12_8_608(.d_in(u_ca_in_608), .d_out(u_ca_out_608));
compressor_12_8 u_ca_12_8_609(.d_in(u_ca_in_609), .d_out(u_ca_out_609));
compressor_12_8 u_ca_12_8_610(.d_in(u_ca_in_610), .d_out(u_ca_out_610));
compressor_12_8 u_ca_12_8_611(.d_in(u_ca_in_611), .d_out(u_ca_out_611));
compressor_12_8 u_ca_12_8_612(.d_in(u_ca_in_612), .d_out(u_ca_out_612));
compressor_12_8 u_ca_12_8_613(.d_in(u_ca_in_613), .d_out(u_ca_out_613));
compressor_12_8 u_ca_12_8_614(.d_in(u_ca_in_614), .d_out(u_ca_out_614));
compressor_12_8 u_ca_12_8_615(.d_in(u_ca_in_615), .d_out(u_ca_out_615));
compressor_12_8 u_ca_12_8_616(.d_in(u_ca_in_616), .d_out(u_ca_out_616));
compressor_12_8 u_ca_12_8_617(.d_in(u_ca_in_617), .d_out(u_ca_out_617));
compressor_12_8 u_ca_12_8_618(.d_in(u_ca_in_618), .d_out(u_ca_out_618));
compressor_12_8 u_ca_12_8_619(.d_in(u_ca_in_619), .d_out(u_ca_out_619));
compressor_12_8 u_ca_12_8_620(.d_in(u_ca_in_620), .d_out(u_ca_out_620));
compressor_12_8 u_ca_12_8_621(.d_in(u_ca_in_621), .d_out(u_ca_out_621));
compressor_12_8 u_ca_12_8_622(.d_in(u_ca_in_622), .d_out(u_ca_out_622));
compressor_12_8 u_ca_12_8_623(.d_in(u_ca_in_623), .d_out(u_ca_out_623));
compressor_12_8 u_ca_12_8_624(.d_in(u_ca_in_624), .d_out(u_ca_out_624));
compressor_12_8 u_ca_12_8_625(.d_in(u_ca_in_625), .d_out(u_ca_out_625));
compressor_12_8 u_ca_12_8_626(.d_in(u_ca_in_626), .d_out(u_ca_out_626));
compressor_12_8 u_ca_12_8_627(.d_in(u_ca_in_627), .d_out(u_ca_out_627));
compressor_12_8 u_ca_12_8_628(.d_in(u_ca_in_628), .d_out(u_ca_out_628));
compressor_12_8 u_ca_12_8_629(.d_in(u_ca_in_629), .d_out(u_ca_out_629));
compressor_12_8 u_ca_12_8_630(.d_in(u_ca_in_630), .d_out(u_ca_out_630));
compressor_12_8 u_ca_12_8_631(.d_in(u_ca_in_631), .d_out(u_ca_out_631));
compressor_12_8 u_ca_12_8_632(.d_in(u_ca_in_632), .d_out(u_ca_out_632));
compressor_12_8 u_ca_12_8_633(.d_in(u_ca_in_633), .d_out(u_ca_out_633));
compressor_12_8 u_ca_12_8_634(.d_in(u_ca_in_634), .d_out(u_ca_out_634));
compressor_12_8 u_ca_12_8_635(.d_in(u_ca_in_635), .d_out(u_ca_out_635));
compressor_12_8 u_ca_12_8_636(.d_in(u_ca_in_636), .d_out(u_ca_out_636));
compressor_12_8 u_ca_12_8_637(.d_in(u_ca_in_637), .d_out(u_ca_out_637));
compressor_12_8 u_ca_12_8_638(.d_in(u_ca_in_638), .d_out(u_ca_out_638));
compressor_12_8 u_ca_12_8_639(.d_in(u_ca_in_639), .d_out(u_ca_out_639));
compressor_12_8 u_ca_12_8_640(.d_in(u_ca_in_640), .d_out(u_ca_out_640));
compressor_12_8 u_ca_12_8_641(.d_in(u_ca_in_641), .d_out(u_ca_out_641));
compressor_12_8 u_ca_12_8_642(.d_in(u_ca_in_642), .d_out(u_ca_out_642));
compressor_12_8 u_ca_12_8_643(.d_in(u_ca_in_643), .d_out(u_ca_out_643));
compressor_12_8 u_ca_12_8_644(.d_in(u_ca_in_644), .d_out(u_ca_out_644));
compressor_12_8 u_ca_12_8_645(.d_in(u_ca_in_645), .d_out(u_ca_out_645));
compressor_12_8 u_ca_12_8_646(.d_in(u_ca_in_646), .d_out(u_ca_out_646));
compressor_12_8 u_ca_12_8_647(.d_in(u_ca_in_647), .d_out(u_ca_out_647));
compressor_12_8 u_ca_12_8_648(.d_in(u_ca_in_648), .d_out(u_ca_out_648));
compressor_12_8 u_ca_12_8_649(.d_in(u_ca_in_649), .d_out(u_ca_out_649));
compressor_12_8 u_ca_12_8_650(.d_in(u_ca_in_650), .d_out(u_ca_out_650));
compressor_12_8 u_ca_12_8_651(.d_in(u_ca_in_651), .d_out(u_ca_out_651));
compressor_12_8 u_ca_12_8_652(.d_in(u_ca_in_652), .d_out(u_ca_out_652));
compressor_12_8 u_ca_12_8_653(.d_in(u_ca_in_653), .d_out(u_ca_out_653));
compressor_12_8 u_ca_12_8_654(.d_in(u_ca_in_654), .d_out(u_ca_out_654));
compressor_12_8 u_ca_12_8_655(.d_in(u_ca_in_655), .d_out(u_ca_out_655));
compressor_12_8 u_ca_12_8_656(.d_in(u_ca_in_656), .d_out(u_ca_out_656));
compressor_12_8 u_ca_12_8_657(.d_in(u_ca_in_657), .d_out(u_ca_out_657));
compressor_12_8 u_ca_12_8_658(.d_in(u_ca_in_658), .d_out(u_ca_out_658));
compressor_12_8 u_ca_12_8_659(.d_in(u_ca_in_659), .d_out(u_ca_out_659));
compressor_12_8 u_ca_12_8_660(.d_in(u_ca_in_660), .d_out(u_ca_out_660));
compressor_12_8 u_ca_12_8_661(.d_in(u_ca_in_661), .d_out(u_ca_out_661));
compressor_12_8 u_ca_12_8_662(.d_in(u_ca_in_662), .d_out(u_ca_out_662));
compressor_12_8 u_ca_12_8_663(.d_in(u_ca_in_663), .d_out(u_ca_out_663));
compressor_12_8 u_ca_12_8_664(.d_in(u_ca_in_664), .d_out(u_ca_out_664));
compressor_12_8 u_ca_12_8_665(.d_in(u_ca_in_665), .d_out(u_ca_out_665));
compressor_12_8 u_ca_12_8_666(.d_in(u_ca_in_666), .d_out(u_ca_out_666));
compressor_12_8 u_ca_12_8_667(.d_in(u_ca_in_667), .d_out(u_ca_out_667));
compressor_12_8 u_ca_12_8_668(.d_in(u_ca_in_668), .d_out(u_ca_out_668));
compressor_12_8 u_ca_12_8_669(.d_in(u_ca_in_669), .d_out(u_ca_out_669));
compressor_12_8 u_ca_12_8_670(.d_in(u_ca_in_670), .d_out(u_ca_out_670));
compressor_12_8 u_ca_12_8_671(.d_in(u_ca_in_671), .d_out(u_ca_out_671));
compressor_12_8 u_ca_12_8_672(.d_in(u_ca_in_672), .d_out(u_ca_out_672));
compressor_12_8 u_ca_12_8_673(.d_in(u_ca_in_673), .d_out(u_ca_out_673));
compressor_12_8 u_ca_12_8_674(.d_in(u_ca_in_674), .d_out(u_ca_out_674));
compressor_12_8 u_ca_12_8_675(.d_in(u_ca_in_675), .d_out(u_ca_out_675));
compressor_12_8 u_ca_12_8_676(.d_in(u_ca_in_676), .d_out(u_ca_out_676));
compressor_12_8 u_ca_12_8_677(.d_in(u_ca_in_677), .d_out(u_ca_out_677));
compressor_12_8 u_ca_12_8_678(.d_in(u_ca_in_678), .d_out(u_ca_out_678));
compressor_12_8 u_ca_12_8_679(.d_in(u_ca_in_679), .d_out(u_ca_out_679));
compressor_12_8 u_ca_12_8_680(.d_in(u_ca_in_680), .d_out(u_ca_out_680));
compressor_12_8 u_ca_12_8_681(.d_in(u_ca_in_681), .d_out(u_ca_out_681));
compressor_12_8 u_ca_12_8_682(.d_in(u_ca_in_682), .d_out(u_ca_out_682));
compressor_12_8 u_ca_12_8_683(.d_in(u_ca_in_683), .d_out(u_ca_out_683));
compressor_12_8 u_ca_12_8_684(.d_in(u_ca_in_684), .d_out(u_ca_out_684));
compressor_12_8 u_ca_12_8_685(.d_in(u_ca_in_685), .d_out(u_ca_out_685));
compressor_12_8 u_ca_12_8_686(.d_in(u_ca_in_686), .d_out(u_ca_out_686));
compressor_12_8 u_ca_12_8_687(.d_in(u_ca_in_687), .d_out(u_ca_out_687));
compressor_12_8 u_ca_12_8_688(.d_in(u_ca_in_688), .d_out(u_ca_out_688));
compressor_12_8 u_ca_12_8_689(.d_in(u_ca_in_689), .d_out(u_ca_out_689));
compressor_12_8 u_ca_12_8_690(.d_in(u_ca_in_690), .d_out(u_ca_out_690));
compressor_12_8 u_ca_12_8_691(.d_in(u_ca_in_691), .d_out(u_ca_out_691));
compressor_12_8 u_ca_12_8_692(.d_in(u_ca_in_692), .d_out(u_ca_out_692));
compressor_12_8 u_ca_12_8_693(.d_in(u_ca_in_693), .d_out(u_ca_out_693));
compressor_12_8 u_ca_12_8_694(.d_in(u_ca_in_694), .d_out(u_ca_out_694));
compressor_12_8 u_ca_12_8_695(.d_in(u_ca_in_695), .d_out(u_ca_out_695));
compressor_12_8 u_ca_12_8_696(.d_in(u_ca_in_696), .d_out(u_ca_out_696));
compressor_12_8 u_ca_12_8_697(.d_in(u_ca_in_697), .d_out(u_ca_out_697));
compressor_12_8 u_ca_12_8_698(.d_in(u_ca_in_698), .d_out(u_ca_out_698));
compressor_12_8 u_ca_12_8_699(.d_in(u_ca_in_699), .d_out(u_ca_out_699));
compressor_12_8 u_ca_12_8_700(.d_in(u_ca_in_700), .d_out(u_ca_out_700));
compressor_12_8 u_ca_12_8_701(.d_in(u_ca_in_701), .d_out(u_ca_out_701));
compressor_12_8 u_ca_12_8_702(.d_in(u_ca_in_702), .d_out(u_ca_out_702));
compressor_12_8 u_ca_12_8_703(.d_in(u_ca_in_703), .d_out(u_ca_out_703));
compressor_12_8 u_ca_12_8_704(.d_in(u_ca_in_704), .d_out(u_ca_out_704));
compressor_12_8 u_ca_12_8_705(.d_in(u_ca_in_705), .d_out(u_ca_out_705));
compressor_12_8 u_ca_12_8_706(.d_in(u_ca_in_706), .d_out(u_ca_out_706));
compressor_12_8 u_ca_12_8_707(.d_in(u_ca_in_707), .d_out(u_ca_out_707));
compressor_12_8 u_ca_12_8_708(.d_in(u_ca_in_708), .d_out(u_ca_out_708));
compressor_12_8 u_ca_12_8_709(.d_in(u_ca_in_709), .d_out(u_ca_out_709));
compressor_12_8 u_ca_12_8_710(.d_in(u_ca_in_710), .d_out(u_ca_out_710));
compressor_12_8 u_ca_12_8_711(.d_in(u_ca_in_711), .d_out(u_ca_out_711));
compressor_12_8 u_ca_12_8_712(.d_in(u_ca_in_712), .d_out(u_ca_out_712));
compressor_12_8 u_ca_12_8_713(.d_in(u_ca_in_713), .d_out(u_ca_out_713));
compressor_12_8 u_ca_12_8_714(.d_in(u_ca_in_714), .d_out(u_ca_out_714));
compressor_12_8 u_ca_12_8_715(.d_in(u_ca_in_715), .d_out(u_ca_out_715));
compressor_12_8 u_ca_12_8_716(.d_in(u_ca_in_716), .d_out(u_ca_out_716));
compressor_12_8 u_ca_12_8_717(.d_in(u_ca_in_717), .d_out(u_ca_out_717));
compressor_12_8 u_ca_12_8_718(.d_in(u_ca_in_718), .d_out(u_ca_out_718));
compressor_12_8 u_ca_12_8_719(.d_in(u_ca_in_719), .d_out(u_ca_out_719));
compressor_12_8 u_ca_12_8_720(.d_in(u_ca_in_720), .d_out(u_ca_out_720));
compressor_12_8 u_ca_12_8_721(.d_in(u_ca_in_721), .d_out(u_ca_out_721));
compressor_12_8 u_ca_12_8_722(.d_in(u_ca_in_722), .d_out(u_ca_out_722));
compressor_12_8 u_ca_12_8_723(.d_in(u_ca_in_723), .d_out(u_ca_out_723));
compressor_12_8 u_ca_12_8_724(.d_in(u_ca_in_724), .d_out(u_ca_out_724));
compressor_12_8 u_ca_12_8_725(.d_in(u_ca_in_725), .d_out(u_ca_out_725));
compressor_12_8 u_ca_12_8_726(.d_in(u_ca_in_726), .d_out(u_ca_out_726));
compressor_12_8 u_ca_12_8_727(.d_in(u_ca_in_727), .d_out(u_ca_out_727));
compressor_12_8 u_ca_12_8_728(.d_in(u_ca_in_728), .d_out(u_ca_out_728));
compressor_12_8 u_ca_12_8_729(.d_in(u_ca_in_729), .d_out(u_ca_out_729));
compressor_12_8 u_ca_12_8_730(.d_in(u_ca_in_730), .d_out(u_ca_out_730));
compressor_12_8 u_ca_12_8_731(.d_in(u_ca_in_731), .d_out(u_ca_out_731));
compressor_12_8 u_ca_12_8_732(.d_in(u_ca_in_732), .d_out(u_ca_out_732));
compressor_12_8 u_ca_12_8_733(.d_in(u_ca_in_733), .d_out(u_ca_out_733));
compressor_12_8 u_ca_12_8_734(.d_in(u_ca_in_734), .d_out(u_ca_out_734));
compressor_12_8 u_ca_12_8_735(.d_in(u_ca_in_735), .d_out(u_ca_out_735));
compressor_12_8 u_ca_12_8_736(.d_in(u_ca_in_736), .d_out(u_ca_out_736));
compressor_12_8 u_ca_12_8_737(.d_in(u_ca_in_737), .d_out(u_ca_out_737));
compressor_12_8 u_ca_12_8_738(.d_in(u_ca_in_738), .d_out(u_ca_out_738));
compressor_12_8 u_ca_12_8_739(.d_in(u_ca_in_739), .d_out(u_ca_out_739));
compressor_12_8 u_ca_12_8_740(.d_in(u_ca_in_740), .d_out(u_ca_out_740));
compressor_12_8 u_ca_12_8_741(.d_in(u_ca_in_741), .d_out(u_ca_out_741));
compressor_12_8 u_ca_12_8_742(.d_in(u_ca_in_742), .d_out(u_ca_out_742));
compressor_12_8 u_ca_12_8_743(.d_in(u_ca_in_743), .d_out(u_ca_out_743));
compressor_12_8 u_ca_12_8_744(.d_in(u_ca_in_744), .d_out(u_ca_out_744));
compressor_12_8 u_ca_12_8_745(.d_in(u_ca_in_745), .d_out(u_ca_out_745));
compressor_12_8 u_ca_12_8_746(.d_in(u_ca_in_746), .d_out(u_ca_out_746));
compressor_12_8 u_ca_12_8_747(.d_in(u_ca_in_747), .d_out(u_ca_out_747));
compressor_12_8 u_ca_12_8_748(.d_in(u_ca_in_748), .d_out(u_ca_out_748));
compressor_12_8 u_ca_12_8_749(.d_in(u_ca_in_749), .d_out(u_ca_out_749));
compressor_12_8 u_ca_12_8_750(.d_in(u_ca_in_750), .d_out(u_ca_out_750));
compressor_12_8 u_ca_12_8_751(.d_in(u_ca_in_751), .d_out(u_ca_out_751));
compressor_12_8 u_ca_12_8_752(.d_in(u_ca_in_752), .d_out(u_ca_out_752));
compressor_12_8 u_ca_12_8_753(.d_in(u_ca_in_753), .d_out(u_ca_out_753));
compressor_12_8 u_ca_12_8_754(.d_in(u_ca_in_754), .d_out(u_ca_out_754));
compressor_12_8 u_ca_12_8_755(.d_in(u_ca_in_755), .d_out(u_ca_out_755));
compressor_12_8 u_ca_12_8_756(.d_in(u_ca_in_756), .d_out(u_ca_out_756));
compressor_12_8 u_ca_12_8_757(.d_in(u_ca_in_757), .d_out(u_ca_out_757));
compressor_12_8 u_ca_12_8_758(.d_in(u_ca_in_758), .d_out(u_ca_out_758));
compressor_12_8 u_ca_12_8_759(.d_in(u_ca_in_759), .d_out(u_ca_out_759));
compressor_12_8 u_ca_12_8_760(.d_in(u_ca_in_760), .d_out(u_ca_out_760));
compressor_12_8 u_ca_12_8_761(.d_in(u_ca_in_761), .d_out(u_ca_out_761));
compressor_12_8 u_ca_12_8_762(.d_in(u_ca_in_762), .d_out(u_ca_out_762));
compressor_12_8 u_ca_12_8_763(.d_in(u_ca_in_763), .d_out(u_ca_out_763));
compressor_12_8 u_ca_12_8_764(.d_in(u_ca_in_764), .d_out(u_ca_out_764));
compressor_12_8 u_ca_12_8_765(.d_in(u_ca_in_765), .d_out(u_ca_out_765));
compressor_12_8 u_ca_12_8_766(.d_in(u_ca_in_766), .d_out(u_ca_out_766));
compressor_12_8 u_ca_12_8_767(.d_in(u_ca_in_767), .d_out(u_ca_out_767));
compressor_12_8 u_ca_12_8_768(.d_in(u_ca_in_768), .d_out(u_ca_out_768));
compressor_12_8 u_ca_12_8_769(.d_in(u_ca_in_769), .d_out(u_ca_out_769));
compressor_12_8 u_ca_12_8_770(.d_in(u_ca_in_770), .d_out(u_ca_out_770));
compressor_12_8 u_ca_12_8_771(.d_in(u_ca_in_771), .d_out(u_ca_out_771));
compressor_12_8 u_ca_12_8_772(.d_in(u_ca_in_772), .d_out(u_ca_out_772));
compressor_12_8 u_ca_12_8_773(.d_in(u_ca_in_773), .d_out(u_ca_out_773));
compressor_12_8 u_ca_12_8_774(.d_in(u_ca_in_774), .d_out(u_ca_out_774));
compressor_12_8 u_ca_12_8_775(.d_in(u_ca_in_775), .d_out(u_ca_out_775));
compressor_12_8 u_ca_12_8_776(.d_in(u_ca_in_776), .d_out(u_ca_out_776));
compressor_12_8 u_ca_12_8_777(.d_in(u_ca_in_777), .d_out(u_ca_out_777));
compressor_12_8 u_ca_12_8_778(.d_in(u_ca_in_778), .d_out(u_ca_out_778));
compressor_12_8 u_ca_12_8_779(.d_in(u_ca_in_779), .d_out(u_ca_out_779));
compressor_12_8 u_ca_12_8_780(.d_in(u_ca_in_780), .d_out(u_ca_out_780));
compressor_12_8 u_ca_12_8_781(.d_in(u_ca_in_781), .d_out(u_ca_out_781));
compressor_12_8 u_ca_12_8_782(.d_in(u_ca_in_782), .d_out(u_ca_out_782));
compressor_12_8 u_ca_12_8_783(.d_in(u_ca_in_783), .d_out(u_ca_out_783));
compressor_12_8 u_ca_12_8_784(.d_in(u_ca_in_784), .d_out(u_ca_out_784));
compressor_12_8 u_ca_12_8_785(.d_in(u_ca_in_785), .d_out(u_ca_out_785));
compressor_12_8 u_ca_12_8_786(.d_in(u_ca_in_786), .d_out(u_ca_out_786));
compressor_12_8 u_ca_12_8_787(.d_in(u_ca_in_787), .d_out(u_ca_out_787));
compressor_12_8 u_ca_12_8_788(.d_in(u_ca_in_788), .d_out(u_ca_out_788));
compressor_12_8 u_ca_12_8_789(.d_in(u_ca_in_789), .d_out(u_ca_out_789));
compressor_12_8 u_ca_12_8_790(.d_in(u_ca_in_790), .d_out(u_ca_out_790));
compressor_12_8 u_ca_12_8_791(.d_in(u_ca_in_791), .d_out(u_ca_out_791));
compressor_12_8 u_ca_12_8_792(.d_in(u_ca_in_792), .d_out(u_ca_out_792));
compressor_12_8 u_ca_12_8_793(.d_in(u_ca_in_793), .d_out(u_ca_out_793));
compressor_12_8 u_ca_12_8_794(.d_in(u_ca_in_794), .d_out(u_ca_out_794));
compressor_12_8 u_ca_12_8_795(.d_in(u_ca_in_795), .d_out(u_ca_out_795));
compressor_12_8 u_ca_12_8_796(.d_in(u_ca_in_796), .d_out(u_ca_out_796));
compressor_12_8 u_ca_12_8_797(.d_in(u_ca_in_797), .d_out(u_ca_out_797));
compressor_12_8 u_ca_12_8_798(.d_in(u_ca_in_798), .d_out(u_ca_out_798));
compressor_12_8 u_ca_12_8_799(.d_in(u_ca_in_799), .d_out(u_ca_out_799));
compressor_12_8 u_ca_12_8_800(.d_in(u_ca_in_800), .d_out(u_ca_out_800));
compressor_12_8 u_ca_12_8_801(.d_in(u_ca_in_801), .d_out(u_ca_out_801));
compressor_12_8 u_ca_12_8_802(.d_in(u_ca_in_802), .d_out(u_ca_out_802));
compressor_12_8 u_ca_12_8_803(.d_in(u_ca_in_803), .d_out(u_ca_out_803));
compressor_12_8 u_ca_12_8_804(.d_in(u_ca_in_804), .d_out(u_ca_out_804));
compressor_12_8 u_ca_12_8_805(.d_in(u_ca_in_805), .d_out(u_ca_out_805));
compressor_12_8 u_ca_12_8_806(.d_in(u_ca_in_806), .d_out(u_ca_out_806));
compressor_12_8 u_ca_12_8_807(.d_in(u_ca_in_807), .d_out(u_ca_out_807));
compressor_12_8 u_ca_12_8_808(.d_in(u_ca_in_808), .d_out(u_ca_out_808));
compressor_12_8 u_ca_12_8_809(.d_in(u_ca_in_809), .d_out(u_ca_out_809));
compressor_12_8 u_ca_12_8_810(.d_in(u_ca_in_810), .d_out(u_ca_out_810));
compressor_12_8 u_ca_12_8_811(.d_in(u_ca_in_811), .d_out(u_ca_out_811));
compressor_12_8 u_ca_12_8_812(.d_in(u_ca_in_812), .d_out(u_ca_out_812));
compressor_12_8 u_ca_12_8_813(.d_in(u_ca_in_813), .d_out(u_ca_out_813));
compressor_12_8 u_ca_12_8_814(.d_in(u_ca_in_814), .d_out(u_ca_out_814));
compressor_12_8 u_ca_12_8_815(.d_in(u_ca_in_815), .d_out(u_ca_out_815));
compressor_12_8 u_ca_12_8_816(.d_in(u_ca_in_816), .d_out(u_ca_out_816));
compressor_12_8 u_ca_12_8_817(.d_in(u_ca_in_817), .d_out(u_ca_out_817));
compressor_12_8 u_ca_12_8_818(.d_in(u_ca_in_818), .d_out(u_ca_out_818));
compressor_12_8 u_ca_12_8_819(.d_in(u_ca_in_819), .d_out(u_ca_out_819));
compressor_12_8 u_ca_12_8_820(.d_in(u_ca_in_820), .d_out(u_ca_out_820));
compressor_12_8 u_ca_12_8_821(.d_in(u_ca_in_821), .d_out(u_ca_out_821));
compressor_12_8 u_ca_12_8_822(.d_in(u_ca_in_822), .d_out(u_ca_out_822));
compressor_12_8 u_ca_12_8_823(.d_in(u_ca_in_823), .d_out(u_ca_out_823));
compressor_12_8 u_ca_12_8_824(.d_in(u_ca_in_824), .d_out(u_ca_out_824));
compressor_12_8 u_ca_12_8_825(.d_in(u_ca_in_825), .d_out(u_ca_out_825));
compressor_12_8 u_ca_12_8_826(.d_in(u_ca_in_826), .d_out(u_ca_out_826));
compressor_12_8 u_ca_12_8_827(.d_in(u_ca_in_827), .d_out(u_ca_out_827));
compressor_12_8 u_ca_12_8_828(.d_in(u_ca_in_828), .d_out(u_ca_out_828));
compressor_12_8 u_ca_12_8_829(.d_in(u_ca_in_829), .d_out(u_ca_out_829));
compressor_12_8 u_ca_12_8_830(.d_in(u_ca_in_830), .d_out(u_ca_out_830));
compressor_12_8 u_ca_12_8_831(.d_in(u_ca_in_831), .d_out(u_ca_out_831));
compressor_12_8 u_ca_12_8_832(.d_in(u_ca_in_832), .d_out(u_ca_out_832));
compressor_12_8 u_ca_12_8_833(.d_in(u_ca_in_833), .d_out(u_ca_out_833));
compressor_12_8 u_ca_12_8_834(.d_in(u_ca_in_834), .d_out(u_ca_out_834));
compressor_12_8 u_ca_12_8_835(.d_in(u_ca_in_835), .d_out(u_ca_out_835));
compressor_12_8 u_ca_12_8_836(.d_in(u_ca_in_836), .d_out(u_ca_out_836));
compressor_12_8 u_ca_12_8_837(.d_in(u_ca_in_837), .d_out(u_ca_out_837));
compressor_12_8 u_ca_12_8_838(.d_in(u_ca_in_838), .d_out(u_ca_out_838));
compressor_12_8 u_ca_12_8_839(.d_in(u_ca_in_839), .d_out(u_ca_out_839));
compressor_12_8 u_ca_12_8_840(.d_in(u_ca_in_840), .d_out(u_ca_out_840));
compressor_12_8 u_ca_12_8_841(.d_in(u_ca_in_841), .d_out(u_ca_out_841));
compressor_12_8 u_ca_12_8_842(.d_in(u_ca_in_842), .d_out(u_ca_out_842));
compressor_12_8 u_ca_12_8_843(.d_in(u_ca_in_843), .d_out(u_ca_out_843));
compressor_12_8 u_ca_12_8_844(.d_in(u_ca_in_844), .d_out(u_ca_out_844));
compressor_12_8 u_ca_12_8_845(.d_in(u_ca_in_845), .d_out(u_ca_out_845));
compressor_12_8 u_ca_12_8_846(.d_in(u_ca_in_846), .d_out(u_ca_out_846));
compressor_12_8 u_ca_12_8_847(.d_in(u_ca_in_847), .d_out(u_ca_out_847));
compressor_12_8 u_ca_12_8_848(.d_in(u_ca_in_848), .d_out(u_ca_out_848));
compressor_12_8 u_ca_12_8_849(.d_in(u_ca_in_849), .d_out(u_ca_out_849));
compressor_12_8 u_ca_12_8_850(.d_in(u_ca_in_850), .d_out(u_ca_out_850));
compressor_12_8 u_ca_12_8_851(.d_in(u_ca_in_851), .d_out(u_ca_out_851));
compressor_12_8 u_ca_12_8_852(.d_in(u_ca_in_852), .d_out(u_ca_out_852));
compressor_12_8 u_ca_12_8_853(.d_in(u_ca_in_853), .d_out(u_ca_out_853));
compressor_12_8 u_ca_12_8_854(.d_in(u_ca_in_854), .d_out(u_ca_out_854));
compressor_12_8 u_ca_12_8_855(.d_in(u_ca_in_855), .d_out(u_ca_out_855));
compressor_12_8 u_ca_12_8_856(.d_in(u_ca_in_856), .d_out(u_ca_out_856));
compressor_12_8 u_ca_12_8_857(.d_in(u_ca_in_857), .d_out(u_ca_out_857));
compressor_12_8 u_ca_12_8_858(.d_in(u_ca_in_858), .d_out(u_ca_out_858));
compressor_12_8 u_ca_12_8_859(.d_in(u_ca_in_859), .d_out(u_ca_out_859));
compressor_12_8 u_ca_12_8_860(.d_in(u_ca_in_860), .d_out(u_ca_out_860));
compressor_12_8 u_ca_12_8_861(.d_in(u_ca_in_861), .d_out(u_ca_out_861));
compressor_12_8 u_ca_12_8_862(.d_in(u_ca_in_862), .d_out(u_ca_out_862));
compressor_12_8 u_ca_12_8_863(.d_in(u_ca_in_863), .d_out(u_ca_out_863));
compressor_12_8 u_ca_12_8_864(.d_in(u_ca_in_864), .d_out(u_ca_out_864));
compressor_12_8 u_ca_12_8_865(.d_in(u_ca_in_865), .d_out(u_ca_out_865));
compressor_12_8 u_ca_12_8_866(.d_in(u_ca_in_866), .d_out(u_ca_out_866));
compressor_12_8 u_ca_12_8_867(.d_in(u_ca_in_867), .d_out(u_ca_out_867));
compressor_12_8 u_ca_12_8_868(.d_in(u_ca_in_868), .d_out(u_ca_out_868));
compressor_12_8 u_ca_12_8_869(.d_in(u_ca_in_869), .d_out(u_ca_out_869));
compressor_12_8 u_ca_12_8_870(.d_in(u_ca_in_870), .d_out(u_ca_out_870));
compressor_12_8 u_ca_12_8_871(.d_in(u_ca_in_871), .d_out(u_ca_out_871));
compressor_12_8 u_ca_12_8_872(.d_in(u_ca_in_872), .d_out(u_ca_out_872));
compressor_12_8 u_ca_12_8_873(.d_in(u_ca_in_873), .d_out(u_ca_out_873));
compressor_12_8 u_ca_12_8_874(.d_in(u_ca_in_874), .d_out(u_ca_out_874));
compressor_12_8 u_ca_12_8_875(.d_in(u_ca_in_875), .d_out(u_ca_out_875));
compressor_12_8 u_ca_12_8_876(.d_in(u_ca_in_876), .d_out(u_ca_out_876));
compressor_12_8 u_ca_12_8_877(.d_in(u_ca_in_877), .d_out(u_ca_out_877));
compressor_12_8 u_ca_12_8_878(.d_in(u_ca_in_878), .d_out(u_ca_out_878));
compressor_12_8 u_ca_12_8_879(.d_in(u_ca_in_879), .d_out(u_ca_out_879));
compressor_12_8 u_ca_12_8_880(.d_in(u_ca_in_880), .d_out(u_ca_out_880));
compressor_12_8 u_ca_12_8_881(.d_in(u_ca_in_881), .d_out(u_ca_out_881));
compressor_12_8 u_ca_12_8_882(.d_in(u_ca_in_882), .d_out(u_ca_out_882));
compressor_12_8 u_ca_12_8_883(.d_in(u_ca_in_883), .d_out(u_ca_out_883));
compressor_12_8 u_ca_12_8_884(.d_in(u_ca_in_884), .d_out(u_ca_out_884));
compressor_12_8 u_ca_12_8_885(.d_in(u_ca_in_885), .d_out(u_ca_out_885));
compressor_12_8 u_ca_12_8_886(.d_in(u_ca_in_886), .d_out(u_ca_out_886));
compressor_12_8 u_ca_12_8_887(.d_in(u_ca_in_887), .d_out(u_ca_out_887));
compressor_12_8 u_ca_12_8_888(.d_in(u_ca_in_888), .d_out(u_ca_out_888));
compressor_12_8 u_ca_12_8_889(.d_in(u_ca_in_889), .d_out(u_ca_out_889));
compressor_12_8 u_ca_12_8_890(.d_in(u_ca_in_890), .d_out(u_ca_out_890));
compressor_12_8 u_ca_12_8_891(.d_in(u_ca_in_891), .d_out(u_ca_out_891));
compressor_12_8 u_ca_12_8_892(.d_in(u_ca_in_892), .d_out(u_ca_out_892));
compressor_12_8 u_ca_12_8_893(.d_in(u_ca_in_893), .d_out(u_ca_out_893));
compressor_12_8 u_ca_12_8_894(.d_in(u_ca_in_894), .d_out(u_ca_out_894));
compressor_12_8 u_ca_12_8_895(.d_in(u_ca_in_895), .d_out(u_ca_out_895));
compressor_12_8 u_ca_12_8_896(.d_in(u_ca_in_896), .d_out(u_ca_out_896));
compressor_12_8 u_ca_12_8_897(.d_in(u_ca_in_897), .d_out(u_ca_out_897));
compressor_12_8 u_ca_12_8_898(.d_in(u_ca_in_898), .d_out(u_ca_out_898));
compressor_12_8 u_ca_12_8_899(.d_in(u_ca_in_899), .d_out(u_ca_out_899));
compressor_12_8 u_ca_12_8_900(.d_in(u_ca_in_900), .d_out(u_ca_out_900));
compressor_12_8 u_ca_12_8_901(.d_in(u_ca_in_901), .d_out(u_ca_out_901));
compressor_12_8 u_ca_12_8_902(.d_in(u_ca_in_902), .d_out(u_ca_out_902));
compressor_12_8 u_ca_12_8_903(.d_in(u_ca_in_903), .d_out(u_ca_out_903));
compressor_12_8 u_ca_12_8_904(.d_in(u_ca_in_904), .d_out(u_ca_out_904));
compressor_12_8 u_ca_12_8_905(.d_in(u_ca_in_905), .d_out(u_ca_out_905));
compressor_12_8 u_ca_12_8_906(.d_in(u_ca_in_906), .d_out(u_ca_out_906));
compressor_12_8 u_ca_12_8_907(.d_in(u_ca_in_907), .d_out(u_ca_out_907));
compressor_12_8 u_ca_12_8_908(.d_in(u_ca_in_908), .d_out(u_ca_out_908));
compressor_12_8 u_ca_12_8_909(.d_in(u_ca_in_909), .d_out(u_ca_out_909));
compressor_12_8 u_ca_12_8_910(.d_in(u_ca_in_910), .d_out(u_ca_out_910));
compressor_12_8 u_ca_12_8_911(.d_in(u_ca_in_911), .d_out(u_ca_out_911));
compressor_12_8 u_ca_12_8_912(.d_in(u_ca_in_912), .d_out(u_ca_out_912));
compressor_12_8 u_ca_12_8_913(.d_in(u_ca_in_913), .d_out(u_ca_out_913));
compressor_12_8 u_ca_12_8_914(.d_in(u_ca_in_914), .d_out(u_ca_out_914));
compressor_12_8 u_ca_12_8_915(.d_in(u_ca_in_915), .d_out(u_ca_out_915));
compressor_12_8 u_ca_12_8_916(.d_in(u_ca_in_916), .d_out(u_ca_out_916));
compressor_12_8 u_ca_12_8_917(.d_in(u_ca_in_917), .d_out(u_ca_out_917));
compressor_12_8 u_ca_12_8_918(.d_in(u_ca_in_918), .d_out(u_ca_out_918));
compressor_12_8 u_ca_12_8_919(.d_in(u_ca_in_919), .d_out(u_ca_out_919));
compressor_12_8 u_ca_12_8_920(.d_in(u_ca_in_920), .d_out(u_ca_out_920));
compressor_12_8 u_ca_12_8_921(.d_in(u_ca_in_921), .d_out(u_ca_out_921));
compressor_12_8 u_ca_12_8_922(.d_in(u_ca_in_922), .d_out(u_ca_out_922));
compressor_12_8 u_ca_12_8_923(.d_in(u_ca_in_923), .d_out(u_ca_out_923));
compressor_12_8 u_ca_12_8_924(.d_in(u_ca_in_924), .d_out(u_ca_out_924));
compressor_12_8 u_ca_12_8_925(.d_in(u_ca_in_925), .d_out(u_ca_out_925));
compressor_12_8 u_ca_12_8_926(.d_in(u_ca_in_926), .d_out(u_ca_out_926));
compressor_12_8 u_ca_12_8_927(.d_in(u_ca_in_927), .d_out(u_ca_out_927));
compressor_12_8 u_ca_12_8_928(.d_in(u_ca_in_928), .d_out(u_ca_out_928));
compressor_12_8 u_ca_12_8_929(.d_in(u_ca_in_929), .d_out(u_ca_out_929));
compressor_12_8 u_ca_12_8_930(.d_in(u_ca_in_930), .d_out(u_ca_out_930));
compressor_12_8 u_ca_12_8_931(.d_in(u_ca_in_931), .d_out(u_ca_out_931));
compressor_12_8 u_ca_12_8_932(.d_in(u_ca_in_932), .d_out(u_ca_out_932));
compressor_12_8 u_ca_12_8_933(.d_in(u_ca_in_933), .d_out(u_ca_out_933));
compressor_12_8 u_ca_12_8_934(.d_in(u_ca_in_934), .d_out(u_ca_out_934));
compressor_12_8 u_ca_12_8_935(.d_in(u_ca_in_935), .d_out(u_ca_out_935));
compressor_12_8 u_ca_12_8_936(.d_in(u_ca_in_936), .d_out(u_ca_out_936));
compressor_12_8 u_ca_12_8_937(.d_in(u_ca_in_937), .d_out(u_ca_out_937));
compressor_12_8 u_ca_12_8_938(.d_in(u_ca_in_938), .d_out(u_ca_out_938));
compressor_12_8 u_ca_12_8_939(.d_in(u_ca_in_939), .d_out(u_ca_out_939));
compressor_12_8 u_ca_12_8_940(.d_in(u_ca_in_940), .d_out(u_ca_out_940));
compressor_12_8 u_ca_12_8_941(.d_in(u_ca_in_941), .d_out(u_ca_out_941));
compressor_12_8 u_ca_12_8_942(.d_in(u_ca_in_942), .d_out(u_ca_out_942));
compressor_12_8 u_ca_12_8_943(.d_in(u_ca_in_943), .d_out(u_ca_out_943));
compressor_12_8 u_ca_12_8_944(.d_in(u_ca_in_944), .d_out(u_ca_out_944));
compressor_12_8 u_ca_12_8_945(.d_in(u_ca_in_945), .d_out(u_ca_out_945));
compressor_12_8 u_ca_12_8_946(.d_in(u_ca_in_946), .d_out(u_ca_out_946));
compressor_12_8 u_ca_12_8_947(.d_in(u_ca_in_947), .d_out(u_ca_out_947));
compressor_12_8 u_ca_12_8_948(.d_in(u_ca_in_948), .d_out(u_ca_out_948));
compressor_12_8 u_ca_12_8_949(.d_in(u_ca_in_949), .d_out(u_ca_out_949));
compressor_12_8 u_ca_12_8_950(.d_in(u_ca_in_950), .d_out(u_ca_out_950));
compressor_12_8 u_ca_12_8_951(.d_in(u_ca_in_951), .d_out(u_ca_out_951));
compressor_12_8 u_ca_12_8_952(.d_in(u_ca_in_952), .d_out(u_ca_out_952));
compressor_12_8 u_ca_12_8_953(.d_in(u_ca_in_953), .d_out(u_ca_out_953));
compressor_12_8 u_ca_12_8_954(.d_in(u_ca_in_954), .d_out(u_ca_out_954));
compressor_12_8 u_ca_12_8_955(.d_in(u_ca_in_955), .d_out(u_ca_out_955));
compressor_12_8 u_ca_12_8_956(.d_in(u_ca_in_956), .d_out(u_ca_out_956));
compressor_12_8 u_ca_12_8_957(.d_in(u_ca_in_957), .d_out(u_ca_out_957));
compressor_12_8 u_ca_12_8_958(.d_in(u_ca_in_958), .d_out(u_ca_out_958));
compressor_12_8 u_ca_12_8_959(.d_in(u_ca_in_959), .d_out(u_ca_out_959));
compressor_12_8 u_ca_12_8_960(.d_in(u_ca_in_960), .d_out(u_ca_out_960));
compressor_12_8 u_ca_12_8_961(.d_in(u_ca_in_961), .d_out(u_ca_out_961));
compressor_12_8 u_ca_12_8_962(.d_in(u_ca_in_962), .d_out(u_ca_out_962));
compressor_12_8 u_ca_12_8_963(.d_in(u_ca_in_963), .d_out(u_ca_out_963));
compressor_12_8 u_ca_12_8_964(.d_in(u_ca_in_964), .d_out(u_ca_out_964));
compressor_12_8 u_ca_12_8_965(.d_in(u_ca_in_965), .d_out(u_ca_out_965));
compressor_12_8 u_ca_12_8_966(.d_in(u_ca_in_966), .d_out(u_ca_out_966));
compressor_12_8 u_ca_12_8_967(.d_in(u_ca_in_967), .d_out(u_ca_out_967));
compressor_12_8 u_ca_12_8_968(.d_in(u_ca_in_968), .d_out(u_ca_out_968));
compressor_12_8 u_ca_12_8_969(.d_in(u_ca_in_969), .d_out(u_ca_out_969));
compressor_12_8 u_ca_12_8_970(.d_in(u_ca_in_970), .d_out(u_ca_out_970));
compressor_12_8 u_ca_12_8_971(.d_in(u_ca_in_971), .d_out(u_ca_out_971));
compressor_12_8 u_ca_12_8_972(.d_in(u_ca_in_972), .d_out(u_ca_out_972));
compressor_12_8 u_ca_12_8_973(.d_in(u_ca_in_973), .d_out(u_ca_out_973));
compressor_12_8 u_ca_12_8_974(.d_in(u_ca_in_974), .d_out(u_ca_out_974));
compressor_12_8 u_ca_12_8_975(.d_in(u_ca_in_975), .d_out(u_ca_out_975));
compressor_12_8 u_ca_12_8_976(.d_in(u_ca_in_976), .d_out(u_ca_out_976));
compressor_12_8 u_ca_12_8_977(.d_in(u_ca_in_977), .d_out(u_ca_out_977));
compressor_12_8 u_ca_12_8_978(.d_in(u_ca_in_978), .d_out(u_ca_out_978));
compressor_12_8 u_ca_12_8_979(.d_in(u_ca_in_979), .d_out(u_ca_out_979));
compressor_12_8 u_ca_12_8_980(.d_in(u_ca_in_980), .d_out(u_ca_out_980));
compressor_12_8 u_ca_12_8_981(.d_in(u_ca_in_981), .d_out(u_ca_out_981));
compressor_12_8 u_ca_12_8_982(.d_in(u_ca_in_982), .d_out(u_ca_out_982));
compressor_12_8 u_ca_12_8_983(.d_in(u_ca_in_983), .d_out(u_ca_out_983));
compressor_12_8 u_ca_12_8_984(.d_in(u_ca_in_984), .d_out(u_ca_out_984));
compressor_12_8 u_ca_12_8_985(.d_in(u_ca_in_985), .d_out(u_ca_out_985));
compressor_12_8 u_ca_12_8_986(.d_in(u_ca_in_986), .d_out(u_ca_out_986));
compressor_12_8 u_ca_12_8_987(.d_in(u_ca_in_987), .d_out(u_ca_out_987));
compressor_12_8 u_ca_12_8_988(.d_in(u_ca_in_988), .d_out(u_ca_out_988));
compressor_12_8 u_ca_12_8_989(.d_in(u_ca_in_989), .d_out(u_ca_out_989));
compressor_12_8 u_ca_12_8_990(.d_in(u_ca_in_990), .d_out(u_ca_out_990));
compressor_12_8 u_ca_12_8_991(.d_in(u_ca_in_991), .d_out(u_ca_out_991));
compressor_12_8 u_ca_12_8_992(.d_in(u_ca_in_992), .d_out(u_ca_out_992));
compressor_12_8 u_ca_12_8_993(.d_in(u_ca_in_993), .d_out(u_ca_out_993));
compressor_12_8 u_ca_12_8_994(.d_in(u_ca_in_994), .d_out(u_ca_out_994));
compressor_12_8 u_ca_12_8_995(.d_in(u_ca_in_995), .d_out(u_ca_out_995));
compressor_12_8 u_ca_12_8_996(.d_in(u_ca_in_996), .d_out(u_ca_out_996));
compressor_12_8 u_ca_12_8_997(.d_in(u_ca_in_997), .d_out(u_ca_out_997));
compressor_12_8 u_ca_12_8_998(.d_in(u_ca_in_998), .d_out(u_ca_out_998));
compressor_12_8 u_ca_12_8_999(.d_in(u_ca_in_999), .d_out(u_ca_out_999));
compressor_12_8 u_ca_12_8_1000(.d_in(u_ca_in_1000), .d_out(u_ca_out_1000));
compressor_12_8 u_ca_12_8_1001(.d_in(u_ca_in_1001), .d_out(u_ca_out_1001));
compressor_12_8 u_ca_12_8_1002(.d_in(u_ca_in_1002), .d_out(u_ca_out_1002));
compressor_12_8 u_ca_12_8_1003(.d_in(u_ca_in_1003), .d_out(u_ca_out_1003));
compressor_12_8 u_ca_12_8_1004(.d_in(u_ca_in_1004), .d_out(u_ca_out_1004));
compressor_12_8 u_ca_12_8_1005(.d_in(u_ca_in_1005), .d_out(u_ca_out_1005));
compressor_12_8 u_ca_12_8_1006(.d_in(u_ca_in_1006), .d_out(u_ca_out_1006));
compressor_12_8 u_ca_12_8_1007(.d_in(u_ca_in_1007), .d_out(u_ca_out_1007));
compressor_12_8 u_ca_12_8_1008(.d_in(u_ca_in_1008), .d_out(u_ca_out_1008));
compressor_12_8 u_ca_12_8_1009(.d_in(u_ca_in_1009), .d_out(u_ca_out_1009));
compressor_12_8 u_ca_12_8_1010(.d_in(u_ca_in_1010), .d_out(u_ca_out_1010));
compressor_12_8 u_ca_12_8_1011(.d_in(u_ca_in_1011), .d_out(u_ca_out_1011));
compressor_12_8 u_ca_12_8_1012(.d_in(u_ca_in_1012), .d_out(u_ca_out_1012));
compressor_12_8 u_ca_12_8_1013(.d_in(u_ca_in_1013), .d_out(u_ca_out_1013));
compressor_12_8 u_ca_12_8_1014(.d_in(u_ca_in_1014), .d_out(u_ca_out_1014));
compressor_12_8 u_ca_12_8_1015(.d_in(u_ca_in_1015), .d_out(u_ca_out_1015));
compressor_12_8 u_ca_12_8_1016(.d_in(u_ca_in_1016), .d_out(u_ca_out_1016));
compressor_12_8 u_ca_12_8_1017(.d_in(u_ca_in_1017), .d_out(u_ca_out_1017));
compressor_12_8 u_ca_12_8_1018(.d_in(u_ca_in_1018), .d_out(u_ca_out_1018));
compressor_12_8 u_ca_12_8_1019(.d_in(u_ca_in_1019), .d_out(u_ca_out_1019));
compressor_12_8 u_ca_12_8_1020(.d_in(u_ca_in_1020), .d_out(u_ca_out_1020));
compressor_12_8 u_ca_12_8_1021(.d_in(u_ca_in_1021), .d_out(u_ca_out_1021));
compressor_12_8 u_ca_12_8_1022(.d_in(u_ca_in_1022), .d_out(u_ca_out_1022));
compressor_12_8 u_ca_12_8_1023(.d_in(u_ca_in_1023), .d_out(u_ca_out_1023));
compressor_12_8 u_ca_12_8_1024(.d_in(u_ca_in_1024), .d_out(u_ca_out_1024));
compressor_12_8 u_ca_12_8_1025(.d_in(u_ca_in_1025), .d_out(u_ca_out_1025));
compressor_12_8 u_ca_12_8_1026(.d_in(u_ca_in_1026), .d_out(u_ca_out_1026));
compressor_12_8 u_ca_12_8_1027(.d_in(u_ca_in_1027), .d_out(u_ca_out_1027));
compressor_12_8 u_ca_12_8_1028(.d_in(u_ca_in_1028), .d_out(u_ca_out_1028));
compressor_12_8 u_ca_12_8_1029(.d_in(u_ca_in_1029), .d_out(u_ca_out_1029));
compressor_12_8 u_ca_12_8_1030(.d_in(u_ca_in_1030), .d_out(u_ca_out_1030));
compressor_12_8 u_ca_12_8_1031(.d_in(u_ca_in_1031), .d_out(u_ca_out_1031));
compressor_12_8 u_ca_12_8_1032(.d_in(u_ca_in_1032), .d_out(u_ca_out_1032));


//---------------------------------------------------------



//--output-------------------------------------------------

assign col_out_0 = {{4{1'b0}}, u_ca_out_0[3:0]};
assign col_out_1 = {u_ca_out_1[3:0], u_ca_out_0[7:4]};
assign col_out_2 = {u_ca_out_2[3:0], u_ca_out_1[7:4]};
assign col_out_3 = {u_ca_out_3[3:0], u_ca_out_2[7:4]};
assign col_out_4 = {u_ca_out_4[3:0], u_ca_out_3[7:4]};
assign col_out_5 = {u_ca_out_5[3:0], u_ca_out_4[7:4]};
assign col_out_6 = {u_ca_out_6[3:0], u_ca_out_5[7:4]};
assign col_out_7 = {u_ca_out_7[3:0], u_ca_out_6[7:4]};
assign col_out_8 = {u_ca_out_8[3:0], u_ca_out_7[7:4]};
assign col_out_9 = {u_ca_out_9[3:0], u_ca_out_8[7:4]};
assign col_out_10 = {u_ca_out_10[3:0], u_ca_out_9[7:4]};
assign col_out_11 = {u_ca_out_11[3:0], u_ca_out_10[7:4]};
assign col_out_12 = {u_ca_out_12[3:0], u_ca_out_11[7:4]};
assign col_out_13 = {u_ca_out_13[3:0], u_ca_out_12[7:4]};
assign col_out_14 = {u_ca_out_14[3:0], u_ca_out_13[7:4]};
assign col_out_15 = {u_ca_out_15[3:0], u_ca_out_14[7:4]};
assign col_out_16 = {u_ca_out_16[3:0], u_ca_out_15[7:4]};
assign col_out_17 = {u_ca_out_17[3:0], u_ca_out_16[7:4]};
assign col_out_18 = {u_ca_out_18[3:0], u_ca_out_17[7:4]};
assign col_out_19 = {u_ca_out_19[3:0], u_ca_out_18[7:4]};
assign col_out_20 = {u_ca_out_20[3:0], u_ca_out_19[7:4]};
assign col_out_21 = {u_ca_out_21[3:0], u_ca_out_20[7:4]};
assign col_out_22 = {u_ca_out_22[3:0], u_ca_out_21[7:4]};
assign col_out_23 = {u_ca_out_23[3:0], u_ca_out_22[7:4]};
assign col_out_24 = {u_ca_out_24[3:0], u_ca_out_23[7:4]};
assign col_out_25 = {u_ca_out_25[3:0], u_ca_out_24[7:4]};
assign col_out_26 = {u_ca_out_26[3:0], u_ca_out_25[7:4]};
assign col_out_27 = {u_ca_out_27[3:0], u_ca_out_26[7:4]};
assign col_out_28 = {u_ca_out_28[3:0], u_ca_out_27[7:4]};
assign col_out_29 = {u_ca_out_29[3:0], u_ca_out_28[7:4]};
assign col_out_30 = {u_ca_out_30[3:0], u_ca_out_29[7:4]};
assign col_out_31 = {u_ca_out_31[3:0], u_ca_out_30[7:4]};
assign col_out_32 = {u_ca_out_32[3:0], u_ca_out_31[7:4]};
assign col_out_33 = {u_ca_out_33[3:0], u_ca_out_32[7:4]};
assign col_out_34 = {u_ca_out_34[3:0], u_ca_out_33[7:4]};
assign col_out_35 = {u_ca_out_35[3:0], u_ca_out_34[7:4]};
assign col_out_36 = {u_ca_out_36[3:0], u_ca_out_35[7:4]};
assign col_out_37 = {u_ca_out_37[3:0], u_ca_out_36[7:4]};
assign col_out_38 = {u_ca_out_38[3:0], u_ca_out_37[7:4]};
assign col_out_39 = {u_ca_out_39[3:0], u_ca_out_38[7:4]};
assign col_out_40 = {u_ca_out_40[3:0], u_ca_out_39[7:4]};
assign col_out_41 = {u_ca_out_41[3:0], u_ca_out_40[7:4]};
assign col_out_42 = {u_ca_out_42[3:0], u_ca_out_41[7:4]};
assign col_out_43 = {u_ca_out_43[3:0], u_ca_out_42[7:4]};
assign col_out_44 = {u_ca_out_44[3:0], u_ca_out_43[7:4]};
assign col_out_45 = {u_ca_out_45[3:0], u_ca_out_44[7:4]};
assign col_out_46 = {u_ca_out_46[3:0], u_ca_out_45[7:4]};
assign col_out_47 = {u_ca_out_47[3:0], u_ca_out_46[7:4]};
assign col_out_48 = {u_ca_out_48[3:0], u_ca_out_47[7:4]};
assign col_out_49 = {u_ca_out_49[3:0], u_ca_out_48[7:4]};
assign col_out_50 = {u_ca_out_50[3:0], u_ca_out_49[7:4]};
assign col_out_51 = {u_ca_out_51[3:0], u_ca_out_50[7:4]};
assign col_out_52 = {u_ca_out_52[3:0], u_ca_out_51[7:4]};
assign col_out_53 = {u_ca_out_53[3:0], u_ca_out_52[7:4]};
assign col_out_54 = {u_ca_out_54[3:0], u_ca_out_53[7:4]};
assign col_out_55 = {u_ca_out_55[3:0], u_ca_out_54[7:4]};
assign col_out_56 = {u_ca_out_56[3:0], u_ca_out_55[7:4]};
assign col_out_57 = {u_ca_out_57[3:0], u_ca_out_56[7:4]};
assign col_out_58 = {u_ca_out_58[3:0], u_ca_out_57[7:4]};
assign col_out_59 = {u_ca_out_59[3:0], u_ca_out_58[7:4]};
assign col_out_60 = {u_ca_out_60[3:0], u_ca_out_59[7:4]};
assign col_out_61 = {u_ca_out_61[3:0], u_ca_out_60[7:4]};
assign col_out_62 = {u_ca_out_62[3:0], u_ca_out_61[7:4]};
assign col_out_63 = {u_ca_out_63[3:0], u_ca_out_62[7:4]};
assign col_out_64 = {u_ca_out_64[3:0], u_ca_out_63[7:4]};
assign col_out_65 = {u_ca_out_65[3:0], u_ca_out_64[7:4]};
assign col_out_66 = {u_ca_out_66[3:0], u_ca_out_65[7:4]};
assign col_out_67 = {u_ca_out_67[3:0], u_ca_out_66[7:4]};
assign col_out_68 = {u_ca_out_68[3:0], u_ca_out_67[7:4]};
assign col_out_69 = {u_ca_out_69[3:0], u_ca_out_68[7:4]};
assign col_out_70 = {u_ca_out_70[3:0], u_ca_out_69[7:4]};
assign col_out_71 = {u_ca_out_71[3:0], u_ca_out_70[7:4]};
assign col_out_72 = {u_ca_out_72[3:0], u_ca_out_71[7:4]};
assign col_out_73 = {u_ca_out_73[3:0], u_ca_out_72[7:4]};
assign col_out_74 = {u_ca_out_74[3:0], u_ca_out_73[7:4]};
assign col_out_75 = {u_ca_out_75[3:0], u_ca_out_74[7:4]};
assign col_out_76 = {u_ca_out_76[3:0], u_ca_out_75[7:4]};
assign col_out_77 = {u_ca_out_77[3:0], u_ca_out_76[7:4]};
assign col_out_78 = {u_ca_out_78[3:0], u_ca_out_77[7:4]};
assign col_out_79 = {u_ca_out_79[3:0], u_ca_out_78[7:4]};
assign col_out_80 = {u_ca_out_80[3:0], u_ca_out_79[7:4]};
assign col_out_81 = {u_ca_out_81[3:0], u_ca_out_80[7:4]};
assign col_out_82 = {u_ca_out_82[3:0], u_ca_out_81[7:4]};
assign col_out_83 = {u_ca_out_83[3:0], u_ca_out_82[7:4]};
assign col_out_84 = {u_ca_out_84[3:0], u_ca_out_83[7:4]};
assign col_out_85 = {u_ca_out_85[3:0], u_ca_out_84[7:4]};
assign col_out_86 = {u_ca_out_86[3:0], u_ca_out_85[7:4]};
assign col_out_87 = {u_ca_out_87[3:0], u_ca_out_86[7:4]};
assign col_out_88 = {u_ca_out_88[3:0], u_ca_out_87[7:4]};
assign col_out_89 = {u_ca_out_89[3:0], u_ca_out_88[7:4]};
assign col_out_90 = {u_ca_out_90[3:0], u_ca_out_89[7:4]};
assign col_out_91 = {u_ca_out_91[3:0], u_ca_out_90[7:4]};
assign col_out_92 = {u_ca_out_92[3:0], u_ca_out_91[7:4]};
assign col_out_93 = {u_ca_out_93[3:0], u_ca_out_92[7:4]};
assign col_out_94 = {u_ca_out_94[3:0], u_ca_out_93[7:4]};
assign col_out_95 = {u_ca_out_95[3:0], u_ca_out_94[7:4]};
assign col_out_96 = {u_ca_out_96[3:0], u_ca_out_95[7:4]};
assign col_out_97 = {u_ca_out_97[3:0], u_ca_out_96[7:4]};
assign col_out_98 = {u_ca_out_98[3:0], u_ca_out_97[7:4]};
assign col_out_99 = {u_ca_out_99[3:0], u_ca_out_98[7:4]};
assign col_out_100 = {u_ca_out_100[3:0], u_ca_out_99[7:4]};
assign col_out_101 = {u_ca_out_101[3:0], u_ca_out_100[7:4]};
assign col_out_102 = {u_ca_out_102[3:0], u_ca_out_101[7:4]};
assign col_out_103 = {u_ca_out_103[3:0], u_ca_out_102[7:4]};
assign col_out_104 = {u_ca_out_104[3:0], u_ca_out_103[7:4]};
assign col_out_105 = {u_ca_out_105[3:0], u_ca_out_104[7:4]};
assign col_out_106 = {u_ca_out_106[3:0], u_ca_out_105[7:4]};
assign col_out_107 = {u_ca_out_107[3:0], u_ca_out_106[7:4]};
assign col_out_108 = {u_ca_out_108[3:0], u_ca_out_107[7:4]};
assign col_out_109 = {u_ca_out_109[3:0], u_ca_out_108[7:4]};
assign col_out_110 = {u_ca_out_110[3:0], u_ca_out_109[7:4]};
assign col_out_111 = {u_ca_out_111[3:0], u_ca_out_110[7:4]};
assign col_out_112 = {u_ca_out_112[3:0], u_ca_out_111[7:4]};
assign col_out_113 = {u_ca_out_113[3:0], u_ca_out_112[7:4]};
assign col_out_114 = {u_ca_out_114[3:0], u_ca_out_113[7:4]};
assign col_out_115 = {u_ca_out_115[3:0], u_ca_out_114[7:4]};
assign col_out_116 = {u_ca_out_116[3:0], u_ca_out_115[7:4]};
assign col_out_117 = {u_ca_out_117[3:0], u_ca_out_116[7:4]};
assign col_out_118 = {u_ca_out_118[3:0], u_ca_out_117[7:4]};
assign col_out_119 = {u_ca_out_119[3:0], u_ca_out_118[7:4]};
assign col_out_120 = {u_ca_out_120[3:0], u_ca_out_119[7:4]};
assign col_out_121 = {u_ca_out_121[3:0], u_ca_out_120[7:4]};
assign col_out_122 = {u_ca_out_122[3:0], u_ca_out_121[7:4]};
assign col_out_123 = {u_ca_out_123[3:0], u_ca_out_122[7:4]};
assign col_out_124 = {u_ca_out_124[3:0], u_ca_out_123[7:4]};
assign col_out_125 = {u_ca_out_125[3:0], u_ca_out_124[7:4]};
assign col_out_126 = {u_ca_out_126[3:0], u_ca_out_125[7:4]};
assign col_out_127 = {u_ca_out_127[3:0], u_ca_out_126[7:4]};
assign col_out_128 = {u_ca_out_128[3:0], u_ca_out_127[7:4]};
assign col_out_129 = {u_ca_out_129[3:0], u_ca_out_128[7:4]};
assign col_out_130 = {u_ca_out_130[3:0], u_ca_out_129[7:4]};
assign col_out_131 = {u_ca_out_131[3:0], u_ca_out_130[7:4]};
assign col_out_132 = {u_ca_out_132[3:0], u_ca_out_131[7:4]};
assign col_out_133 = {u_ca_out_133[3:0], u_ca_out_132[7:4]};
assign col_out_134 = {u_ca_out_134[3:0], u_ca_out_133[7:4]};
assign col_out_135 = {u_ca_out_135[3:0], u_ca_out_134[7:4]};
assign col_out_136 = {u_ca_out_136[3:0], u_ca_out_135[7:4]};
assign col_out_137 = {u_ca_out_137[3:0], u_ca_out_136[7:4]};
assign col_out_138 = {u_ca_out_138[3:0], u_ca_out_137[7:4]};
assign col_out_139 = {u_ca_out_139[3:0], u_ca_out_138[7:4]};
assign col_out_140 = {u_ca_out_140[3:0], u_ca_out_139[7:4]};
assign col_out_141 = {u_ca_out_141[3:0], u_ca_out_140[7:4]};
assign col_out_142 = {u_ca_out_142[3:0], u_ca_out_141[7:4]};
assign col_out_143 = {u_ca_out_143[3:0], u_ca_out_142[7:4]};
assign col_out_144 = {u_ca_out_144[3:0], u_ca_out_143[7:4]};
assign col_out_145 = {u_ca_out_145[3:0], u_ca_out_144[7:4]};
assign col_out_146 = {u_ca_out_146[3:0], u_ca_out_145[7:4]};
assign col_out_147 = {u_ca_out_147[3:0], u_ca_out_146[7:4]};
assign col_out_148 = {u_ca_out_148[3:0], u_ca_out_147[7:4]};
assign col_out_149 = {u_ca_out_149[3:0], u_ca_out_148[7:4]};
assign col_out_150 = {u_ca_out_150[3:0], u_ca_out_149[7:4]};
assign col_out_151 = {u_ca_out_151[3:0], u_ca_out_150[7:4]};
assign col_out_152 = {u_ca_out_152[3:0], u_ca_out_151[7:4]};
assign col_out_153 = {u_ca_out_153[3:0], u_ca_out_152[7:4]};
assign col_out_154 = {u_ca_out_154[3:0], u_ca_out_153[7:4]};
assign col_out_155 = {u_ca_out_155[3:0], u_ca_out_154[7:4]};
assign col_out_156 = {u_ca_out_156[3:0], u_ca_out_155[7:4]};
assign col_out_157 = {u_ca_out_157[3:0], u_ca_out_156[7:4]};
assign col_out_158 = {u_ca_out_158[3:0], u_ca_out_157[7:4]};
assign col_out_159 = {u_ca_out_159[3:0], u_ca_out_158[7:4]};
assign col_out_160 = {u_ca_out_160[3:0], u_ca_out_159[7:4]};
assign col_out_161 = {u_ca_out_161[3:0], u_ca_out_160[7:4]};
assign col_out_162 = {u_ca_out_162[3:0], u_ca_out_161[7:4]};
assign col_out_163 = {u_ca_out_163[3:0], u_ca_out_162[7:4]};
assign col_out_164 = {u_ca_out_164[3:0], u_ca_out_163[7:4]};
assign col_out_165 = {u_ca_out_165[3:0], u_ca_out_164[7:4]};
assign col_out_166 = {u_ca_out_166[3:0], u_ca_out_165[7:4]};
assign col_out_167 = {u_ca_out_167[3:0], u_ca_out_166[7:4]};
assign col_out_168 = {u_ca_out_168[3:0], u_ca_out_167[7:4]};
assign col_out_169 = {u_ca_out_169[3:0], u_ca_out_168[7:4]};
assign col_out_170 = {u_ca_out_170[3:0], u_ca_out_169[7:4]};
assign col_out_171 = {u_ca_out_171[3:0], u_ca_out_170[7:4]};
assign col_out_172 = {u_ca_out_172[3:0], u_ca_out_171[7:4]};
assign col_out_173 = {u_ca_out_173[3:0], u_ca_out_172[7:4]};
assign col_out_174 = {u_ca_out_174[3:0], u_ca_out_173[7:4]};
assign col_out_175 = {u_ca_out_175[3:0], u_ca_out_174[7:4]};
assign col_out_176 = {u_ca_out_176[3:0], u_ca_out_175[7:4]};
assign col_out_177 = {u_ca_out_177[3:0], u_ca_out_176[7:4]};
assign col_out_178 = {u_ca_out_178[3:0], u_ca_out_177[7:4]};
assign col_out_179 = {u_ca_out_179[3:0], u_ca_out_178[7:4]};
assign col_out_180 = {u_ca_out_180[3:0], u_ca_out_179[7:4]};
assign col_out_181 = {u_ca_out_181[3:0], u_ca_out_180[7:4]};
assign col_out_182 = {u_ca_out_182[3:0], u_ca_out_181[7:4]};
assign col_out_183 = {u_ca_out_183[3:0], u_ca_out_182[7:4]};
assign col_out_184 = {u_ca_out_184[3:0], u_ca_out_183[7:4]};
assign col_out_185 = {u_ca_out_185[3:0], u_ca_out_184[7:4]};
assign col_out_186 = {u_ca_out_186[3:0], u_ca_out_185[7:4]};
assign col_out_187 = {u_ca_out_187[3:0], u_ca_out_186[7:4]};
assign col_out_188 = {u_ca_out_188[3:0], u_ca_out_187[7:4]};
assign col_out_189 = {u_ca_out_189[3:0], u_ca_out_188[7:4]};
assign col_out_190 = {u_ca_out_190[3:0], u_ca_out_189[7:4]};
assign col_out_191 = {u_ca_out_191[3:0], u_ca_out_190[7:4]};
assign col_out_192 = {u_ca_out_192[3:0], u_ca_out_191[7:4]};
assign col_out_193 = {u_ca_out_193[3:0], u_ca_out_192[7:4]};
assign col_out_194 = {u_ca_out_194[3:0], u_ca_out_193[7:4]};
assign col_out_195 = {u_ca_out_195[3:0], u_ca_out_194[7:4]};
assign col_out_196 = {u_ca_out_196[3:0], u_ca_out_195[7:4]};
assign col_out_197 = {u_ca_out_197[3:0], u_ca_out_196[7:4]};
assign col_out_198 = {u_ca_out_198[3:0], u_ca_out_197[7:4]};
assign col_out_199 = {u_ca_out_199[3:0], u_ca_out_198[7:4]};
assign col_out_200 = {u_ca_out_200[3:0], u_ca_out_199[7:4]};
assign col_out_201 = {u_ca_out_201[3:0], u_ca_out_200[7:4]};
assign col_out_202 = {u_ca_out_202[3:0], u_ca_out_201[7:4]};
assign col_out_203 = {u_ca_out_203[3:0], u_ca_out_202[7:4]};
assign col_out_204 = {u_ca_out_204[3:0], u_ca_out_203[7:4]};
assign col_out_205 = {u_ca_out_205[3:0], u_ca_out_204[7:4]};
assign col_out_206 = {u_ca_out_206[3:0], u_ca_out_205[7:4]};
assign col_out_207 = {u_ca_out_207[3:0], u_ca_out_206[7:4]};
assign col_out_208 = {u_ca_out_208[3:0], u_ca_out_207[7:4]};
assign col_out_209 = {u_ca_out_209[3:0], u_ca_out_208[7:4]};
assign col_out_210 = {u_ca_out_210[3:0], u_ca_out_209[7:4]};
assign col_out_211 = {u_ca_out_211[3:0], u_ca_out_210[7:4]};
assign col_out_212 = {u_ca_out_212[3:0], u_ca_out_211[7:4]};
assign col_out_213 = {u_ca_out_213[3:0], u_ca_out_212[7:4]};
assign col_out_214 = {u_ca_out_214[3:0], u_ca_out_213[7:4]};
assign col_out_215 = {u_ca_out_215[3:0], u_ca_out_214[7:4]};
assign col_out_216 = {u_ca_out_216[3:0], u_ca_out_215[7:4]};
assign col_out_217 = {u_ca_out_217[3:0], u_ca_out_216[7:4]};
assign col_out_218 = {u_ca_out_218[3:0], u_ca_out_217[7:4]};
assign col_out_219 = {u_ca_out_219[3:0], u_ca_out_218[7:4]};
assign col_out_220 = {u_ca_out_220[3:0], u_ca_out_219[7:4]};
assign col_out_221 = {u_ca_out_221[3:0], u_ca_out_220[7:4]};
assign col_out_222 = {u_ca_out_222[3:0], u_ca_out_221[7:4]};
assign col_out_223 = {u_ca_out_223[3:0], u_ca_out_222[7:4]};
assign col_out_224 = {u_ca_out_224[3:0], u_ca_out_223[7:4]};
assign col_out_225 = {u_ca_out_225[3:0], u_ca_out_224[7:4]};
assign col_out_226 = {u_ca_out_226[3:0], u_ca_out_225[7:4]};
assign col_out_227 = {u_ca_out_227[3:0], u_ca_out_226[7:4]};
assign col_out_228 = {u_ca_out_228[3:0], u_ca_out_227[7:4]};
assign col_out_229 = {u_ca_out_229[3:0], u_ca_out_228[7:4]};
assign col_out_230 = {u_ca_out_230[3:0], u_ca_out_229[7:4]};
assign col_out_231 = {u_ca_out_231[3:0], u_ca_out_230[7:4]};
assign col_out_232 = {u_ca_out_232[3:0], u_ca_out_231[7:4]};
assign col_out_233 = {u_ca_out_233[3:0], u_ca_out_232[7:4]};
assign col_out_234 = {u_ca_out_234[3:0], u_ca_out_233[7:4]};
assign col_out_235 = {u_ca_out_235[3:0], u_ca_out_234[7:4]};
assign col_out_236 = {u_ca_out_236[3:0], u_ca_out_235[7:4]};
assign col_out_237 = {u_ca_out_237[3:0], u_ca_out_236[7:4]};
assign col_out_238 = {u_ca_out_238[3:0], u_ca_out_237[7:4]};
assign col_out_239 = {u_ca_out_239[3:0], u_ca_out_238[7:4]};
assign col_out_240 = {u_ca_out_240[3:0], u_ca_out_239[7:4]};
assign col_out_241 = {u_ca_out_241[3:0], u_ca_out_240[7:4]};
assign col_out_242 = {u_ca_out_242[3:0], u_ca_out_241[7:4]};
assign col_out_243 = {u_ca_out_243[3:0], u_ca_out_242[7:4]};
assign col_out_244 = {u_ca_out_244[3:0], u_ca_out_243[7:4]};
assign col_out_245 = {u_ca_out_245[3:0], u_ca_out_244[7:4]};
assign col_out_246 = {u_ca_out_246[3:0], u_ca_out_245[7:4]};
assign col_out_247 = {u_ca_out_247[3:0], u_ca_out_246[7:4]};
assign col_out_248 = {u_ca_out_248[3:0], u_ca_out_247[7:4]};
assign col_out_249 = {u_ca_out_249[3:0], u_ca_out_248[7:4]};
assign col_out_250 = {u_ca_out_250[3:0], u_ca_out_249[7:4]};
assign col_out_251 = {u_ca_out_251[3:0], u_ca_out_250[7:4]};
assign col_out_252 = {u_ca_out_252[3:0], u_ca_out_251[7:4]};
assign col_out_253 = {u_ca_out_253[3:0], u_ca_out_252[7:4]};
assign col_out_254 = {u_ca_out_254[3:0], u_ca_out_253[7:4]};
assign col_out_255 = {u_ca_out_255[3:0], u_ca_out_254[7:4]};
assign col_out_256 = {u_ca_out_256[3:0], u_ca_out_255[7:4]};
assign col_out_257 = {u_ca_out_257[3:0], u_ca_out_256[7:4]};
assign col_out_258 = {u_ca_out_258[3:0], u_ca_out_257[7:4]};
assign col_out_259 = {u_ca_out_259[3:0], u_ca_out_258[7:4]};
assign col_out_260 = {u_ca_out_260[3:0], u_ca_out_259[7:4]};
assign col_out_261 = {u_ca_out_261[3:0], u_ca_out_260[7:4]};
assign col_out_262 = {u_ca_out_262[3:0], u_ca_out_261[7:4]};
assign col_out_263 = {u_ca_out_263[3:0], u_ca_out_262[7:4]};
assign col_out_264 = {u_ca_out_264[3:0], u_ca_out_263[7:4]};
assign col_out_265 = {u_ca_out_265[3:0], u_ca_out_264[7:4]};
assign col_out_266 = {u_ca_out_266[3:0], u_ca_out_265[7:4]};
assign col_out_267 = {u_ca_out_267[3:0], u_ca_out_266[7:4]};
assign col_out_268 = {u_ca_out_268[3:0], u_ca_out_267[7:4]};
assign col_out_269 = {u_ca_out_269[3:0], u_ca_out_268[7:4]};
assign col_out_270 = {u_ca_out_270[3:0], u_ca_out_269[7:4]};
assign col_out_271 = {u_ca_out_271[3:0], u_ca_out_270[7:4]};
assign col_out_272 = {u_ca_out_272[3:0], u_ca_out_271[7:4]};
assign col_out_273 = {u_ca_out_273[3:0], u_ca_out_272[7:4]};
assign col_out_274 = {u_ca_out_274[3:0], u_ca_out_273[7:4]};
assign col_out_275 = {u_ca_out_275[3:0], u_ca_out_274[7:4]};
assign col_out_276 = {u_ca_out_276[3:0], u_ca_out_275[7:4]};
assign col_out_277 = {u_ca_out_277[3:0], u_ca_out_276[7:4]};
assign col_out_278 = {u_ca_out_278[3:0], u_ca_out_277[7:4]};
assign col_out_279 = {u_ca_out_279[3:0], u_ca_out_278[7:4]};
assign col_out_280 = {u_ca_out_280[3:0], u_ca_out_279[7:4]};
assign col_out_281 = {u_ca_out_281[3:0], u_ca_out_280[7:4]};
assign col_out_282 = {u_ca_out_282[3:0], u_ca_out_281[7:4]};
assign col_out_283 = {u_ca_out_283[3:0], u_ca_out_282[7:4]};
assign col_out_284 = {u_ca_out_284[3:0], u_ca_out_283[7:4]};
assign col_out_285 = {u_ca_out_285[3:0], u_ca_out_284[7:4]};
assign col_out_286 = {u_ca_out_286[3:0], u_ca_out_285[7:4]};
assign col_out_287 = {u_ca_out_287[3:0], u_ca_out_286[7:4]};
assign col_out_288 = {u_ca_out_288[3:0], u_ca_out_287[7:4]};
assign col_out_289 = {u_ca_out_289[3:0], u_ca_out_288[7:4]};
assign col_out_290 = {u_ca_out_290[3:0], u_ca_out_289[7:4]};
assign col_out_291 = {u_ca_out_291[3:0], u_ca_out_290[7:4]};
assign col_out_292 = {u_ca_out_292[3:0], u_ca_out_291[7:4]};
assign col_out_293 = {u_ca_out_293[3:0], u_ca_out_292[7:4]};
assign col_out_294 = {u_ca_out_294[3:0], u_ca_out_293[7:4]};
assign col_out_295 = {u_ca_out_295[3:0], u_ca_out_294[7:4]};
assign col_out_296 = {u_ca_out_296[3:0], u_ca_out_295[7:4]};
assign col_out_297 = {u_ca_out_297[3:0], u_ca_out_296[7:4]};
assign col_out_298 = {u_ca_out_298[3:0], u_ca_out_297[7:4]};
assign col_out_299 = {u_ca_out_299[3:0], u_ca_out_298[7:4]};
assign col_out_300 = {u_ca_out_300[3:0], u_ca_out_299[7:4]};
assign col_out_301 = {u_ca_out_301[3:0], u_ca_out_300[7:4]};
assign col_out_302 = {u_ca_out_302[3:0], u_ca_out_301[7:4]};
assign col_out_303 = {u_ca_out_303[3:0], u_ca_out_302[7:4]};
assign col_out_304 = {u_ca_out_304[3:0], u_ca_out_303[7:4]};
assign col_out_305 = {u_ca_out_305[3:0], u_ca_out_304[7:4]};
assign col_out_306 = {u_ca_out_306[3:0], u_ca_out_305[7:4]};
assign col_out_307 = {u_ca_out_307[3:0], u_ca_out_306[7:4]};
assign col_out_308 = {u_ca_out_308[3:0], u_ca_out_307[7:4]};
assign col_out_309 = {u_ca_out_309[3:0], u_ca_out_308[7:4]};
assign col_out_310 = {u_ca_out_310[3:0], u_ca_out_309[7:4]};
assign col_out_311 = {u_ca_out_311[3:0], u_ca_out_310[7:4]};
assign col_out_312 = {u_ca_out_312[3:0], u_ca_out_311[7:4]};
assign col_out_313 = {u_ca_out_313[3:0], u_ca_out_312[7:4]};
assign col_out_314 = {u_ca_out_314[3:0], u_ca_out_313[7:4]};
assign col_out_315 = {u_ca_out_315[3:0], u_ca_out_314[7:4]};
assign col_out_316 = {u_ca_out_316[3:0], u_ca_out_315[7:4]};
assign col_out_317 = {u_ca_out_317[3:0], u_ca_out_316[7:4]};
assign col_out_318 = {u_ca_out_318[3:0], u_ca_out_317[7:4]};
assign col_out_319 = {u_ca_out_319[3:0], u_ca_out_318[7:4]};
assign col_out_320 = {u_ca_out_320[3:0], u_ca_out_319[7:4]};
assign col_out_321 = {u_ca_out_321[3:0], u_ca_out_320[7:4]};
assign col_out_322 = {u_ca_out_322[3:0], u_ca_out_321[7:4]};
assign col_out_323 = {u_ca_out_323[3:0], u_ca_out_322[7:4]};
assign col_out_324 = {u_ca_out_324[3:0], u_ca_out_323[7:4]};
assign col_out_325 = {u_ca_out_325[3:0], u_ca_out_324[7:4]};
assign col_out_326 = {u_ca_out_326[3:0], u_ca_out_325[7:4]};
assign col_out_327 = {u_ca_out_327[3:0], u_ca_out_326[7:4]};
assign col_out_328 = {u_ca_out_328[3:0], u_ca_out_327[7:4]};
assign col_out_329 = {u_ca_out_329[3:0], u_ca_out_328[7:4]};
assign col_out_330 = {u_ca_out_330[3:0], u_ca_out_329[7:4]};
assign col_out_331 = {u_ca_out_331[3:0], u_ca_out_330[7:4]};
assign col_out_332 = {u_ca_out_332[3:0], u_ca_out_331[7:4]};
assign col_out_333 = {u_ca_out_333[3:0], u_ca_out_332[7:4]};
assign col_out_334 = {u_ca_out_334[3:0], u_ca_out_333[7:4]};
assign col_out_335 = {u_ca_out_335[3:0], u_ca_out_334[7:4]};
assign col_out_336 = {u_ca_out_336[3:0], u_ca_out_335[7:4]};
assign col_out_337 = {u_ca_out_337[3:0], u_ca_out_336[7:4]};
assign col_out_338 = {u_ca_out_338[3:0], u_ca_out_337[7:4]};
assign col_out_339 = {u_ca_out_339[3:0], u_ca_out_338[7:4]};
assign col_out_340 = {u_ca_out_340[3:0], u_ca_out_339[7:4]};
assign col_out_341 = {u_ca_out_341[3:0], u_ca_out_340[7:4]};
assign col_out_342 = {u_ca_out_342[3:0], u_ca_out_341[7:4]};
assign col_out_343 = {u_ca_out_343[3:0], u_ca_out_342[7:4]};
assign col_out_344 = {u_ca_out_344[3:0], u_ca_out_343[7:4]};
assign col_out_345 = {u_ca_out_345[3:0], u_ca_out_344[7:4]};
assign col_out_346 = {u_ca_out_346[3:0], u_ca_out_345[7:4]};
assign col_out_347 = {u_ca_out_347[3:0], u_ca_out_346[7:4]};
assign col_out_348 = {u_ca_out_348[3:0], u_ca_out_347[7:4]};
assign col_out_349 = {u_ca_out_349[3:0], u_ca_out_348[7:4]};
assign col_out_350 = {u_ca_out_350[3:0], u_ca_out_349[7:4]};
assign col_out_351 = {u_ca_out_351[3:0], u_ca_out_350[7:4]};
assign col_out_352 = {u_ca_out_352[3:0], u_ca_out_351[7:4]};
assign col_out_353 = {u_ca_out_353[3:0], u_ca_out_352[7:4]};
assign col_out_354 = {u_ca_out_354[3:0], u_ca_out_353[7:4]};
assign col_out_355 = {u_ca_out_355[3:0], u_ca_out_354[7:4]};
assign col_out_356 = {u_ca_out_356[3:0], u_ca_out_355[7:4]};
assign col_out_357 = {u_ca_out_357[3:0], u_ca_out_356[7:4]};
assign col_out_358 = {u_ca_out_358[3:0], u_ca_out_357[7:4]};
assign col_out_359 = {u_ca_out_359[3:0], u_ca_out_358[7:4]};
assign col_out_360 = {u_ca_out_360[3:0], u_ca_out_359[7:4]};
assign col_out_361 = {u_ca_out_361[3:0], u_ca_out_360[7:4]};
assign col_out_362 = {u_ca_out_362[3:0], u_ca_out_361[7:4]};
assign col_out_363 = {u_ca_out_363[3:0], u_ca_out_362[7:4]};
assign col_out_364 = {u_ca_out_364[3:0], u_ca_out_363[7:4]};
assign col_out_365 = {u_ca_out_365[3:0], u_ca_out_364[7:4]};
assign col_out_366 = {u_ca_out_366[3:0], u_ca_out_365[7:4]};
assign col_out_367 = {u_ca_out_367[3:0], u_ca_out_366[7:4]};
assign col_out_368 = {u_ca_out_368[3:0], u_ca_out_367[7:4]};
assign col_out_369 = {u_ca_out_369[3:0], u_ca_out_368[7:4]};
assign col_out_370 = {u_ca_out_370[3:0], u_ca_out_369[7:4]};
assign col_out_371 = {u_ca_out_371[3:0], u_ca_out_370[7:4]};
assign col_out_372 = {u_ca_out_372[3:0], u_ca_out_371[7:4]};
assign col_out_373 = {u_ca_out_373[3:0], u_ca_out_372[7:4]};
assign col_out_374 = {u_ca_out_374[3:0], u_ca_out_373[7:4]};
assign col_out_375 = {u_ca_out_375[3:0], u_ca_out_374[7:4]};
assign col_out_376 = {u_ca_out_376[3:0], u_ca_out_375[7:4]};
assign col_out_377 = {u_ca_out_377[3:0], u_ca_out_376[7:4]};
assign col_out_378 = {u_ca_out_378[3:0], u_ca_out_377[7:4]};
assign col_out_379 = {u_ca_out_379[3:0], u_ca_out_378[7:4]};
assign col_out_380 = {u_ca_out_380[3:0], u_ca_out_379[7:4]};
assign col_out_381 = {u_ca_out_381[3:0], u_ca_out_380[7:4]};
assign col_out_382 = {u_ca_out_382[3:0], u_ca_out_381[7:4]};
assign col_out_383 = {u_ca_out_383[3:0], u_ca_out_382[7:4]};
assign col_out_384 = {u_ca_out_384[3:0], u_ca_out_383[7:4]};
assign col_out_385 = {u_ca_out_385[3:0], u_ca_out_384[7:4]};
assign col_out_386 = {u_ca_out_386[3:0], u_ca_out_385[7:4]};
assign col_out_387 = {u_ca_out_387[3:0], u_ca_out_386[7:4]};
assign col_out_388 = {u_ca_out_388[3:0], u_ca_out_387[7:4]};
assign col_out_389 = {u_ca_out_389[3:0], u_ca_out_388[7:4]};
assign col_out_390 = {u_ca_out_390[3:0], u_ca_out_389[7:4]};
assign col_out_391 = {u_ca_out_391[3:0], u_ca_out_390[7:4]};
assign col_out_392 = {u_ca_out_392[3:0], u_ca_out_391[7:4]};
assign col_out_393 = {u_ca_out_393[3:0], u_ca_out_392[7:4]};
assign col_out_394 = {u_ca_out_394[3:0], u_ca_out_393[7:4]};
assign col_out_395 = {u_ca_out_395[3:0], u_ca_out_394[7:4]};
assign col_out_396 = {u_ca_out_396[3:0], u_ca_out_395[7:4]};
assign col_out_397 = {u_ca_out_397[3:0], u_ca_out_396[7:4]};
assign col_out_398 = {u_ca_out_398[3:0], u_ca_out_397[7:4]};
assign col_out_399 = {u_ca_out_399[3:0], u_ca_out_398[7:4]};
assign col_out_400 = {u_ca_out_400[3:0], u_ca_out_399[7:4]};
assign col_out_401 = {u_ca_out_401[3:0], u_ca_out_400[7:4]};
assign col_out_402 = {u_ca_out_402[3:0], u_ca_out_401[7:4]};
assign col_out_403 = {u_ca_out_403[3:0], u_ca_out_402[7:4]};
assign col_out_404 = {u_ca_out_404[3:0], u_ca_out_403[7:4]};
assign col_out_405 = {u_ca_out_405[3:0], u_ca_out_404[7:4]};
assign col_out_406 = {u_ca_out_406[3:0], u_ca_out_405[7:4]};
assign col_out_407 = {u_ca_out_407[3:0], u_ca_out_406[7:4]};
assign col_out_408 = {u_ca_out_408[3:0], u_ca_out_407[7:4]};
assign col_out_409 = {u_ca_out_409[3:0], u_ca_out_408[7:4]};
assign col_out_410 = {u_ca_out_410[3:0], u_ca_out_409[7:4]};
assign col_out_411 = {u_ca_out_411[3:0], u_ca_out_410[7:4]};
assign col_out_412 = {u_ca_out_412[3:0], u_ca_out_411[7:4]};
assign col_out_413 = {u_ca_out_413[3:0], u_ca_out_412[7:4]};
assign col_out_414 = {u_ca_out_414[3:0], u_ca_out_413[7:4]};
assign col_out_415 = {u_ca_out_415[3:0], u_ca_out_414[7:4]};
assign col_out_416 = {u_ca_out_416[3:0], u_ca_out_415[7:4]};
assign col_out_417 = {u_ca_out_417[3:0], u_ca_out_416[7:4]};
assign col_out_418 = {u_ca_out_418[3:0], u_ca_out_417[7:4]};
assign col_out_419 = {u_ca_out_419[3:0], u_ca_out_418[7:4]};
assign col_out_420 = {u_ca_out_420[3:0], u_ca_out_419[7:4]};
assign col_out_421 = {u_ca_out_421[3:0], u_ca_out_420[7:4]};
assign col_out_422 = {u_ca_out_422[3:0], u_ca_out_421[7:4]};
assign col_out_423 = {u_ca_out_423[3:0], u_ca_out_422[7:4]};
assign col_out_424 = {u_ca_out_424[3:0], u_ca_out_423[7:4]};
assign col_out_425 = {u_ca_out_425[3:0], u_ca_out_424[7:4]};
assign col_out_426 = {u_ca_out_426[3:0], u_ca_out_425[7:4]};
assign col_out_427 = {u_ca_out_427[3:0], u_ca_out_426[7:4]};
assign col_out_428 = {u_ca_out_428[3:0], u_ca_out_427[7:4]};
assign col_out_429 = {u_ca_out_429[3:0], u_ca_out_428[7:4]};
assign col_out_430 = {u_ca_out_430[3:0], u_ca_out_429[7:4]};
assign col_out_431 = {u_ca_out_431[3:0], u_ca_out_430[7:4]};
assign col_out_432 = {u_ca_out_432[3:0], u_ca_out_431[7:4]};
assign col_out_433 = {u_ca_out_433[3:0], u_ca_out_432[7:4]};
assign col_out_434 = {u_ca_out_434[3:0], u_ca_out_433[7:4]};
assign col_out_435 = {u_ca_out_435[3:0], u_ca_out_434[7:4]};
assign col_out_436 = {u_ca_out_436[3:0], u_ca_out_435[7:4]};
assign col_out_437 = {u_ca_out_437[3:0], u_ca_out_436[7:4]};
assign col_out_438 = {u_ca_out_438[3:0], u_ca_out_437[7:4]};
assign col_out_439 = {u_ca_out_439[3:0], u_ca_out_438[7:4]};
assign col_out_440 = {u_ca_out_440[3:0], u_ca_out_439[7:4]};
assign col_out_441 = {u_ca_out_441[3:0], u_ca_out_440[7:4]};
assign col_out_442 = {u_ca_out_442[3:0], u_ca_out_441[7:4]};
assign col_out_443 = {u_ca_out_443[3:0], u_ca_out_442[7:4]};
assign col_out_444 = {u_ca_out_444[3:0], u_ca_out_443[7:4]};
assign col_out_445 = {u_ca_out_445[3:0], u_ca_out_444[7:4]};
assign col_out_446 = {u_ca_out_446[3:0], u_ca_out_445[7:4]};
assign col_out_447 = {u_ca_out_447[3:0], u_ca_out_446[7:4]};
assign col_out_448 = {u_ca_out_448[3:0], u_ca_out_447[7:4]};
assign col_out_449 = {u_ca_out_449[3:0], u_ca_out_448[7:4]};
assign col_out_450 = {u_ca_out_450[3:0], u_ca_out_449[7:4]};
assign col_out_451 = {u_ca_out_451[3:0], u_ca_out_450[7:4]};
assign col_out_452 = {u_ca_out_452[3:0], u_ca_out_451[7:4]};
assign col_out_453 = {u_ca_out_453[3:0], u_ca_out_452[7:4]};
assign col_out_454 = {u_ca_out_454[3:0], u_ca_out_453[7:4]};
assign col_out_455 = {u_ca_out_455[3:0], u_ca_out_454[7:4]};
assign col_out_456 = {u_ca_out_456[3:0], u_ca_out_455[7:4]};
assign col_out_457 = {u_ca_out_457[3:0], u_ca_out_456[7:4]};
assign col_out_458 = {u_ca_out_458[3:0], u_ca_out_457[7:4]};
assign col_out_459 = {u_ca_out_459[3:0], u_ca_out_458[7:4]};
assign col_out_460 = {u_ca_out_460[3:0], u_ca_out_459[7:4]};
assign col_out_461 = {u_ca_out_461[3:0], u_ca_out_460[7:4]};
assign col_out_462 = {u_ca_out_462[3:0], u_ca_out_461[7:4]};
assign col_out_463 = {u_ca_out_463[3:0], u_ca_out_462[7:4]};
assign col_out_464 = {u_ca_out_464[3:0], u_ca_out_463[7:4]};
assign col_out_465 = {u_ca_out_465[3:0], u_ca_out_464[7:4]};
assign col_out_466 = {u_ca_out_466[3:0], u_ca_out_465[7:4]};
assign col_out_467 = {u_ca_out_467[3:0], u_ca_out_466[7:4]};
assign col_out_468 = {u_ca_out_468[3:0], u_ca_out_467[7:4]};
assign col_out_469 = {u_ca_out_469[3:0], u_ca_out_468[7:4]};
assign col_out_470 = {u_ca_out_470[3:0], u_ca_out_469[7:4]};
assign col_out_471 = {u_ca_out_471[3:0], u_ca_out_470[7:4]};
assign col_out_472 = {u_ca_out_472[3:0], u_ca_out_471[7:4]};
assign col_out_473 = {u_ca_out_473[3:0], u_ca_out_472[7:4]};
assign col_out_474 = {u_ca_out_474[3:0], u_ca_out_473[7:4]};
assign col_out_475 = {u_ca_out_475[3:0], u_ca_out_474[7:4]};
assign col_out_476 = {u_ca_out_476[3:0], u_ca_out_475[7:4]};
assign col_out_477 = {u_ca_out_477[3:0], u_ca_out_476[7:4]};
assign col_out_478 = {u_ca_out_478[3:0], u_ca_out_477[7:4]};
assign col_out_479 = {u_ca_out_479[3:0], u_ca_out_478[7:4]};
assign col_out_480 = {u_ca_out_480[3:0], u_ca_out_479[7:4]};
assign col_out_481 = {u_ca_out_481[3:0], u_ca_out_480[7:4]};
assign col_out_482 = {u_ca_out_482[3:0], u_ca_out_481[7:4]};
assign col_out_483 = {u_ca_out_483[3:0], u_ca_out_482[7:4]};
assign col_out_484 = {u_ca_out_484[3:0], u_ca_out_483[7:4]};
assign col_out_485 = {u_ca_out_485[3:0], u_ca_out_484[7:4]};
assign col_out_486 = {u_ca_out_486[3:0], u_ca_out_485[7:4]};
assign col_out_487 = {u_ca_out_487[3:0], u_ca_out_486[7:4]};
assign col_out_488 = {u_ca_out_488[3:0], u_ca_out_487[7:4]};
assign col_out_489 = {u_ca_out_489[3:0], u_ca_out_488[7:4]};
assign col_out_490 = {u_ca_out_490[3:0], u_ca_out_489[7:4]};
assign col_out_491 = {u_ca_out_491[3:0], u_ca_out_490[7:4]};
assign col_out_492 = {u_ca_out_492[3:0], u_ca_out_491[7:4]};
assign col_out_493 = {u_ca_out_493[3:0], u_ca_out_492[7:4]};
assign col_out_494 = {u_ca_out_494[3:0], u_ca_out_493[7:4]};
assign col_out_495 = {u_ca_out_495[3:0], u_ca_out_494[7:4]};
assign col_out_496 = {u_ca_out_496[3:0], u_ca_out_495[7:4]};
assign col_out_497 = {u_ca_out_497[3:0], u_ca_out_496[7:4]};
assign col_out_498 = {u_ca_out_498[3:0], u_ca_out_497[7:4]};
assign col_out_499 = {u_ca_out_499[3:0], u_ca_out_498[7:4]};
assign col_out_500 = {u_ca_out_500[3:0], u_ca_out_499[7:4]};
assign col_out_501 = {u_ca_out_501[3:0], u_ca_out_500[7:4]};
assign col_out_502 = {u_ca_out_502[3:0], u_ca_out_501[7:4]};
assign col_out_503 = {u_ca_out_503[3:0], u_ca_out_502[7:4]};
assign col_out_504 = {u_ca_out_504[3:0], u_ca_out_503[7:4]};
assign col_out_505 = {u_ca_out_505[3:0], u_ca_out_504[7:4]};
assign col_out_506 = {u_ca_out_506[3:0], u_ca_out_505[7:4]};
assign col_out_507 = {u_ca_out_507[3:0], u_ca_out_506[7:4]};
assign col_out_508 = {u_ca_out_508[3:0], u_ca_out_507[7:4]};
assign col_out_509 = {u_ca_out_509[3:0], u_ca_out_508[7:4]};
assign col_out_510 = {u_ca_out_510[3:0], u_ca_out_509[7:4]};
assign col_out_511 = {u_ca_out_511[3:0], u_ca_out_510[7:4]};
assign col_out_512 = {u_ca_out_512[3:0], u_ca_out_511[7:4]};
assign col_out_513 = {u_ca_out_513[3:0], u_ca_out_512[7:4]};
assign col_out_514 = {u_ca_out_514[3:0], u_ca_out_513[7:4]};
assign col_out_515 = {u_ca_out_515[3:0], u_ca_out_514[7:4]};
assign col_out_516 = {u_ca_out_516[3:0], u_ca_out_515[7:4]};
assign col_out_517 = {u_ca_out_517[3:0], u_ca_out_516[7:4]};
assign col_out_518 = {u_ca_out_518[3:0], u_ca_out_517[7:4]};
assign col_out_519 = {u_ca_out_519[3:0], u_ca_out_518[7:4]};
assign col_out_520 = {u_ca_out_520[3:0], u_ca_out_519[7:4]};
assign col_out_521 = {u_ca_out_521[3:0], u_ca_out_520[7:4]};
assign col_out_522 = {u_ca_out_522[3:0], u_ca_out_521[7:4]};
assign col_out_523 = {u_ca_out_523[3:0], u_ca_out_522[7:4]};
assign col_out_524 = {u_ca_out_524[3:0], u_ca_out_523[7:4]};
assign col_out_525 = {u_ca_out_525[3:0], u_ca_out_524[7:4]};
assign col_out_526 = {u_ca_out_526[3:0], u_ca_out_525[7:4]};
assign col_out_527 = {u_ca_out_527[3:0], u_ca_out_526[7:4]};
assign col_out_528 = {u_ca_out_528[3:0], u_ca_out_527[7:4]};
assign col_out_529 = {u_ca_out_529[3:0], u_ca_out_528[7:4]};
assign col_out_530 = {u_ca_out_530[3:0], u_ca_out_529[7:4]};
assign col_out_531 = {u_ca_out_531[3:0], u_ca_out_530[7:4]};
assign col_out_532 = {u_ca_out_532[3:0], u_ca_out_531[7:4]};
assign col_out_533 = {u_ca_out_533[3:0], u_ca_out_532[7:4]};
assign col_out_534 = {u_ca_out_534[3:0], u_ca_out_533[7:4]};
assign col_out_535 = {u_ca_out_535[3:0], u_ca_out_534[7:4]};
assign col_out_536 = {u_ca_out_536[3:0], u_ca_out_535[7:4]};
assign col_out_537 = {u_ca_out_537[3:0], u_ca_out_536[7:4]};
assign col_out_538 = {u_ca_out_538[3:0], u_ca_out_537[7:4]};
assign col_out_539 = {u_ca_out_539[3:0], u_ca_out_538[7:4]};
assign col_out_540 = {u_ca_out_540[3:0], u_ca_out_539[7:4]};
assign col_out_541 = {u_ca_out_541[3:0], u_ca_out_540[7:4]};
assign col_out_542 = {u_ca_out_542[3:0], u_ca_out_541[7:4]};
assign col_out_543 = {u_ca_out_543[3:0], u_ca_out_542[7:4]};
assign col_out_544 = {u_ca_out_544[3:0], u_ca_out_543[7:4]};
assign col_out_545 = {u_ca_out_545[3:0], u_ca_out_544[7:4]};
assign col_out_546 = {u_ca_out_546[3:0], u_ca_out_545[7:4]};
assign col_out_547 = {u_ca_out_547[3:0], u_ca_out_546[7:4]};
assign col_out_548 = {u_ca_out_548[3:0], u_ca_out_547[7:4]};
assign col_out_549 = {u_ca_out_549[3:0], u_ca_out_548[7:4]};
assign col_out_550 = {u_ca_out_550[3:0], u_ca_out_549[7:4]};
assign col_out_551 = {u_ca_out_551[3:0], u_ca_out_550[7:4]};
assign col_out_552 = {u_ca_out_552[3:0], u_ca_out_551[7:4]};
assign col_out_553 = {u_ca_out_553[3:0], u_ca_out_552[7:4]};
assign col_out_554 = {u_ca_out_554[3:0], u_ca_out_553[7:4]};
assign col_out_555 = {u_ca_out_555[3:0], u_ca_out_554[7:4]};
assign col_out_556 = {u_ca_out_556[3:0], u_ca_out_555[7:4]};
assign col_out_557 = {u_ca_out_557[3:0], u_ca_out_556[7:4]};
assign col_out_558 = {u_ca_out_558[3:0], u_ca_out_557[7:4]};
assign col_out_559 = {u_ca_out_559[3:0], u_ca_out_558[7:4]};
assign col_out_560 = {u_ca_out_560[3:0], u_ca_out_559[7:4]};
assign col_out_561 = {u_ca_out_561[3:0], u_ca_out_560[7:4]};
assign col_out_562 = {u_ca_out_562[3:0], u_ca_out_561[7:4]};
assign col_out_563 = {u_ca_out_563[3:0], u_ca_out_562[7:4]};
assign col_out_564 = {u_ca_out_564[3:0], u_ca_out_563[7:4]};
assign col_out_565 = {u_ca_out_565[3:0], u_ca_out_564[7:4]};
assign col_out_566 = {u_ca_out_566[3:0], u_ca_out_565[7:4]};
assign col_out_567 = {u_ca_out_567[3:0], u_ca_out_566[7:4]};
assign col_out_568 = {u_ca_out_568[3:0], u_ca_out_567[7:4]};
assign col_out_569 = {u_ca_out_569[3:0], u_ca_out_568[7:4]};
assign col_out_570 = {u_ca_out_570[3:0], u_ca_out_569[7:4]};
assign col_out_571 = {u_ca_out_571[3:0], u_ca_out_570[7:4]};
assign col_out_572 = {u_ca_out_572[3:0], u_ca_out_571[7:4]};
assign col_out_573 = {u_ca_out_573[3:0], u_ca_out_572[7:4]};
assign col_out_574 = {u_ca_out_574[3:0], u_ca_out_573[7:4]};
assign col_out_575 = {u_ca_out_575[3:0], u_ca_out_574[7:4]};
assign col_out_576 = {u_ca_out_576[3:0], u_ca_out_575[7:4]};
assign col_out_577 = {u_ca_out_577[3:0], u_ca_out_576[7:4]};
assign col_out_578 = {u_ca_out_578[3:0], u_ca_out_577[7:4]};
assign col_out_579 = {u_ca_out_579[3:0], u_ca_out_578[7:4]};
assign col_out_580 = {u_ca_out_580[3:0], u_ca_out_579[7:4]};
assign col_out_581 = {u_ca_out_581[3:0], u_ca_out_580[7:4]};
assign col_out_582 = {u_ca_out_582[3:0], u_ca_out_581[7:4]};
assign col_out_583 = {u_ca_out_583[3:0], u_ca_out_582[7:4]};
assign col_out_584 = {u_ca_out_584[3:0], u_ca_out_583[7:4]};
assign col_out_585 = {u_ca_out_585[3:0], u_ca_out_584[7:4]};
assign col_out_586 = {u_ca_out_586[3:0], u_ca_out_585[7:4]};
assign col_out_587 = {u_ca_out_587[3:0], u_ca_out_586[7:4]};
assign col_out_588 = {u_ca_out_588[3:0], u_ca_out_587[7:4]};
assign col_out_589 = {u_ca_out_589[3:0], u_ca_out_588[7:4]};
assign col_out_590 = {u_ca_out_590[3:0], u_ca_out_589[7:4]};
assign col_out_591 = {u_ca_out_591[3:0], u_ca_out_590[7:4]};
assign col_out_592 = {u_ca_out_592[3:0], u_ca_out_591[7:4]};
assign col_out_593 = {u_ca_out_593[3:0], u_ca_out_592[7:4]};
assign col_out_594 = {u_ca_out_594[3:0], u_ca_out_593[7:4]};
assign col_out_595 = {u_ca_out_595[3:0], u_ca_out_594[7:4]};
assign col_out_596 = {u_ca_out_596[3:0], u_ca_out_595[7:4]};
assign col_out_597 = {u_ca_out_597[3:0], u_ca_out_596[7:4]};
assign col_out_598 = {u_ca_out_598[3:0], u_ca_out_597[7:4]};
assign col_out_599 = {u_ca_out_599[3:0], u_ca_out_598[7:4]};
assign col_out_600 = {u_ca_out_600[3:0], u_ca_out_599[7:4]};
assign col_out_601 = {u_ca_out_601[3:0], u_ca_out_600[7:4]};
assign col_out_602 = {u_ca_out_602[3:0], u_ca_out_601[7:4]};
assign col_out_603 = {u_ca_out_603[3:0], u_ca_out_602[7:4]};
assign col_out_604 = {u_ca_out_604[3:0], u_ca_out_603[7:4]};
assign col_out_605 = {u_ca_out_605[3:0], u_ca_out_604[7:4]};
assign col_out_606 = {u_ca_out_606[3:0], u_ca_out_605[7:4]};
assign col_out_607 = {u_ca_out_607[3:0], u_ca_out_606[7:4]};
assign col_out_608 = {u_ca_out_608[3:0], u_ca_out_607[7:4]};
assign col_out_609 = {u_ca_out_609[3:0], u_ca_out_608[7:4]};
assign col_out_610 = {u_ca_out_610[3:0], u_ca_out_609[7:4]};
assign col_out_611 = {u_ca_out_611[3:0], u_ca_out_610[7:4]};
assign col_out_612 = {u_ca_out_612[3:0], u_ca_out_611[7:4]};
assign col_out_613 = {u_ca_out_613[3:0], u_ca_out_612[7:4]};
assign col_out_614 = {u_ca_out_614[3:0], u_ca_out_613[7:4]};
assign col_out_615 = {u_ca_out_615[3:0], u_ca_out_614[7:4]};
assign col_out_616 = {u_ca_out_616[3:0], u_ca_out_615[7:4]};
assign col_out_617 = {u_ca_out_617[3:0], u_ca_out_616[7:4]};
assign col_out_618 = {u_ca_out_618[3:0], u_ca_out_617[7:4]};
assign col_out_619 = {u_ca_out_619[3:0], u_ca_out_618[7:4]};
assign col_out_620 = {u_ca_out_620[3:0], u_ca_out_619[7:4]};
assign col_out_621 = {u_ca_out_621[3:0], u_ca_out_620[7:4]};
assign col_out_622 = {u_ca_out_622[3:0], u_ca_out_621[7:4]};
assign col_out_623 = {u_ca_out_623[3:0], u_ca_out_622[7:4]};
assign col_out_624 = {u_ca_out_624[3:0], u_ca_out_623[7:4]};
assign col_out_625 = {u_ca_out_625[3:0], u_ca_out_624[7:4]};
assign col_out_626 = {u_ca_out_626[3:0], u_ca_out_625[7:4]};
assign col_out_627 = {u_ca_out_627[3:0], u_ca_out_626[7:4]};
assign col_out_628 = {u_ca_out_628[3:0], u_ca_out_627[7:4]};
assign col_out_629 = {u_ca_out_629[3:0], u_ca_out_628[7:4]};
assign col_out_630 = {u_ca_out_630[3:0], u_ca_out_629[7:4]};
assign col_out_631 = {u_ca_out_631[3:0], u_ca_out_630[7:4]};
assign col_out_632 = {u_ca_out_632[3:0], u_ca_out_631[7:4]};
assign col_out_633 = {u_ca_out_633[3:0], u_ca_out_632[7:4]};
assign col_out_634 = {u_ca_out_634[3:0], u_ca_out_633[7:4]};
assign col_out_635 = {u_ca_out_635[3:0], u_ca_out_634[7:4]};
assign col_out_636 = {u_ca_out_636[3:0], u_ca_out_635[7:4]};
assign col_out_637 = {u_ca_out_637[3:0], u_ca_out_636[7:4]};
assign col_out_638 = {u_ca_out_638[3:0], u_ca_out_637[7:4]};
assign col_out_639 = {u_ca_out_639[3:0], u_ca_out_638[7:4]};
assign col_out_640 = {u_ca_out_640[3:0], u_ca_out_639[7:4]};
assign col_out_641 = {u_ca_out_641[3:0], u_ca_out_640[7:4]};
assign col_out_642 = {u_ca_out_642[3:0], u_ca_out_641[7:4]};
assign col_out_643 = {u_ca_out_643[3:0], u_ca_out_642[7:4]};
assign col_out_644 = {u_ca_out_644[3:0], u_ca_out_643[7:4]};
assign col_out_645 = {u_ca_out_645[3:0], u_ca_out_644[7:4]};
assign col_out_646 = {u_ca_out_646[3:0], u_ca_out_645[7:4]};
assign col_out_647 = {u_ca_out_647[3:0], u_ca_out_646[7:4]};
assign col_out_648 = {u_ca_out_648[3:0], u_ca_out_647[7:4]};
assign col_out_649 = {u_ca_out_649[3:0], u_ca_out_648[7:4]};
assign col_out_650 = {u_ca_out_650[3:0], u_ca_out_649[7:4]};
assign col_out_651 = {u_ca_out_651[3:0], u_ca_out_650[7:4]};
assign col_out_652 = {u_ca_out_652[3:0], u_ca_out_651[7:4]};
assign col_out_653 = {u_ca_out_653[3:0], u_ca_out_652[7:4]};
assign col_out_654 = {u_ca_out_654[3:0], u_ca_out_653[7:4]};
assign col_out_655 = {u_ca_out_655[3:0], u_ca_out_654[7:4]};
assign col_out_656 = {u_ca_out_656[3:0], u_ca_out_655[7:4]};
assign col_out_657 = {u_ca_out_657[3:0], u_ca_out_656[7:4]};
assign col_out_658 = {u_ca_out_658[3:0], u_ca_out_657[7:4]};
assign col_out_659 = {u_ca_out_659[3:0], u_ca_out_658[7:4]};
assign col_out_660 = {u_ca_out_660[3:0], u_ca_out_659[7:4]};
assign col_out_661 = {u_ca_out_661[3:0], u_ca_out_660[7:4]};
assign col_out_662 = {u_ca_out_662[3:0], u_ca_out_661[7:4]};
assign col_out_663 = {u_ca_out_663[3:0], u_ca_out_662[7:4]};
assign col_out_664 = {u_ca_out_664[3:0], u_ca_out_663[7:4]};
assign col_out_665 = {u_ca_out_665[3:0], u_ca_out_664[7:4]};
assign col_out_666 = {u_ca_out_666[3:0], u_ca_out_665[7:4]};
assign col_out_667 = {u_ca_out_667[3:0], u_ca_out_666[7:4]};
assign col_out_668 = {u_ca_out_668[3:0], u_ca_out_667[7:4]};
assign col_out_669 = {u_ca_out_669[3:0], u_ca_out_668[7:4]};
assign col_out_670 = {u_ca_out_670[3:0], u_ca_out_669[7:4]};
assign col_out_671 = {u_ca_out_671[3:0], u_ca_out_670[7:4]};
assign col_out_672 = {u_ca_out_672[3:0], u_ca_out_671[7:4]};
assign col_out_673 = {u_ca_out_673[3:0], u_ca_out_672[7:4]};
assign col_out_674 = {u_ca_out_674[3:0], u_ca_out_673[7:4]};
assign col_out_675 = {u_ca_out_675[3:0], u_ca_out_674[7:4]};
assign col_out_676 = {u_ca_out_676[3:0], u_ca_out_675[7:4]};
assign col_out_677 = {u_ca_out_677[3:0], u_ca_out_676[7:4]};
assign col_out_678 = {u_ca_out_678[3:0], u_ca_out_677[7:4]};
assign col_out_679 = {u_ca_out_679[3:0], u_ca_out_678[7:4]};
assign col_out_680 = {u_ca_out_680[3:0], u_ca_out_679[7:4]};
assign col_out_681 = {u_ca_out_681[3:0], u_ca_out_680[7:4]};
assign col_out_682 = {u_ca_out_682[3:0], u_ca_out_681[7:4]};
assign col_out_683 = {u_ca_out_683[3:0], u_ca_out_682[7:4]};
assign col_out_684 = {u_ca_out_684[3:0], u_ca_out_683[7:4]};
assign col_out_685 = {u_ca_out_685[3:0], u_ca_out_684[7:4]};
assign col_out_686 = {u_ca_out_686[3:0], u_ca_out_685[7:4]};
assign col_out_687 = {u_ca_out_687[3:0], u_ca_out_686[7:4]};
assign col_out_688 = {u_ca_out_688[3:0], u_ca_out_687[7:4]};
assign col_out_689 = {u_ca_out_689[3:0], u_ca_out_688[7:4]};
assign col_out_690 = {u_ca_out_690[3:0], u_ca_out_689[7:4]};
assign col_out_691 = {u_ca_out_691[3:0], u_ca_out_690[7:4]};
assign col_out_692 = {u_ca_out_692[3:0], u_ca_out_691[7:4]};
assign col_out_693 = {u_ca_out_693[3:0], u_ca_out_692[7:4]};
assign col_out_694 = {u_ca_out_694[3:0], u_ca_out_693[7:4]};
assign col_out_695 = {u_ca_out_695[3:0], u_ca_out_694[7:4]};
assign col_out_696 = {u_ca_out_696[3:0], u_ca_out_695[7:4]};
assign col_out_697 = {u_ca_out_697[3:0], u_ca_out_696[7:4]};
assign col_out_698 = {u_ca_out_698[3:0], u_ca_out_697[7:4]};
assign col_out_699 = {u_ca_out_699[3:0], u_ca_out_698[7:4]};
assign col_out_700 = {u_ca_out_700[3:0], u_ca_out_699[7:4]};
assign col_out_701 = {u_ca_out_701[3:0], u_ca_out_700[7:4]};
assign col_out_702 = {u_ca_out_702[3:0], u_ca_out_701[7:4]};
assign col_out_703 = {u_ca_out_703[3:0], u_ca_out_702[7:4]};
assign col_out_704 = {u_ca_out_704[3:0], u_ca_out_703[7:4]};
assign col_out_705 = {u_ca_out_705[3:0], u_ca_out_704[7:4]};
assign col_out_706 = {u_ca_out_706[3:0], u_ca_out_705[7:4]};
assign col_out_707 = {u_ca_out_707[3:0], u_ca_out_706[7:4]};
assign col_out_708 = {u_ca_out_708[3:0], u_ca_out_707[7:4]};
assign col_out_709 = {u_ca_out_709[3:0], u_ca_out_708[7:4]};
assign col_out_710 = {u_ca_out_710[3:0], u_ca_out_709[7:4]};
assign col_out_711 = {u_ca_out_711[3:0], u_ca_out_710[7:4]};
assign col_out_712 = {u_ca_out_712[3:0], u_ca_out_711[7:4]};
assign col_out_713 = {u_ca_out_713[3:0], u_ca_out_712[7:4]};
assign col_out_714 = {u_ca_out_714[3:0], u_ca_out_713[7:4]};
assign col_out_715 = {u_ca_out_715[3:0], u_ca_out_714[7:4]};
assign col_out_716 = {u_ca_out_716[3:0], u_ca_out_715[7:4]};
assign col_out_717 = {u_ca_out_717[3:0], u_ca_out_716[7:4]};
assign col_out_718 = {u_ca_out_718[3:0], u_ca_out_717[7:4]};
assign col_out_719 = {u_ca_out_719[3:0], u_ca_out_718[7:4]};
assign col_out_720 = {u_ca_out_720[3:0], u_ca_out_719[7:4]};
assign col_out_721 = {u_ca_out_721[3:0], u_ca_out_720[7:4]};
assign col_out_722 = {u_ca_out_722[3:0], u_ca_out_721[7:4]};
assign col_out_723 = {u_ca_out_723[3:0], u_ca_out_722[7:4]};
assign col_out_724 = {u_ca_out_724[3:0], u_ca_out_723[7:4]};
assign col_out_725 = {u_ca_out_725[3:0], u_ca_out_724[7:4]};
assign col_out_726 = {u_ca_out_726[3:0], u_ca_out_725[7:4]};
assign col_out_727 = {u_ca_out_727[3:0], u_ca_out_726[7:4]};
assign col_out_728 = {u_ca_out_728[3:0], u_ca_out_727[7:4]};
assign col_out_729 = {u_ca_out_729[3:0], u_ca_out_728[7:4]};
assign col_out_730 = {u_ca_out_730[3:0], u_ca_out_729[7:4]};
assign col_out_731 = {u_ca_out_731[3:0], u_ca_out_730[7:4]};
assign col_out_732 = {u_ca_out_732[3:0], u_ca_out_731[7:4]};
assign col_out_733 = {u_ca_out_733[3:0], u_ca_out_732[7:4]};
assign col_out_734 = {u_ca_out_734[3:0], u_ca_out_733[7:4]};
assign col_out_735 = {u_ca_out_735[3:0], u_ca_out_734[7:4]};
assign col_out_736 = {u_ca_out_736[3:0], u_ca_out_735[7:4]};
assign col_out_737 = {u_ca_out_737[3:0], u_ca_out_736[7:4]};
assign col_out_738 = {u_ca_out_738[3:0], u_ca_out_737[7:4]};
assign col_out_739 = {u_ca_out_739[3:0], u_ca_out_738[7:4]};
assign col_out_740 = {u_ca_out_740[3:0], u_ca_out_739[7:4]};
assign col_out_741 = {u_ca_out_741[3:0], u_ca_out_740[7:4]};
assign col_out_742 = {u_ca_out_742[3:0], u_ca_out_741[7:4]};
assign col_out_743 = {u_ca_out_743[3:0], u_ca_out_742[7:4]};
assign col_out_744 = {u_ca_out_744[3:0], u_ca_out_743[7:4]};
assign col_out_745 = {u_ca_out_745[3:0], u_ca_out_744[7:4]};
assign col_out_746 = {u_ca_out_746[3:0], u_ca_out_745[7:4]};
assign col_out_747 = {u_ca_out_747[3:0], u_ca_out_746[7:4]};
assign col_out_748 = {u_ca_out_748[3:0], u_ca_out_747[7:4]};
assign col_out_749 = {u_ca_out_749[3:0], u_ca_out_748[7:4]};
assign col_out_750 = {u_ca_out_750[3:0], u_ca_out_749[7:4]};
assign col_out_751 = {u_ca_out_751[3:0], u_ca_out_750[7:4]};
assign col_out_752 = {u_ca_out_752[3:0], u_ca_out_751[7:4]};
assign col_out_753 = {u_ca_out_753[3:0], u_ca_out_752[7:4]};
assign col_out_754 = {u_ca_out_754[3:0], u_ca_out_753[7:4]};
assign col_out_755 = {u_ca_out_755[3:0], u_ca_out_754[7:4]};
assign col_out_756 = {u_ca_out_756[3:0], u_ca_out_755[7:4]};
assign col_out_757 = {u_ca_out_757[3:0], u_ca_out_756[7:4]};
assign col_out_758 = {u_ca_out_758[3:0], u_ca_out_757[7:4]};
assign col_out_759 = {u_ca_out_759[3:0], u_ca_out_758[7:4]};
assign col_out_760 = {u_ca_out_760[3:0], u_ca_out_759[7:4]};
assign col_out_761 = {u_ca_out_761[3:0], u_ca_out_760[7:4]};
assign col_out_762 = {u_ca_out_762[3:0], u_ca_out_761[7:4]};
assign col_out_763 = {u_ca_out_763[3:0], u_ca_out_762[7:4]};
assign col_out_764 = {u_ca_out_764[3:0], u_ca_out_763[7:4]};
assign col_out_765 = {u_ca_out_765[3:0], u_ca_out_764[7:4]};
assign col_out_766 = {u_ca_out_766[3:0], u_ca_out_765[7:4]};
assign col_out_767 = {u_ca_out_767[3:0], u_ca_out_766[7:4]};
assign col_out_768 = {u_ca_out_768[3:0], u_ca_out_767[7:4]};
assign col_out_769 = {u_ca_out_769[3:0], u_ca_out_768[7:4]};
assign col_out_770 = {u_ca_out_770[3:0], u_ca_out_769[7:4]};
assign col_out_771 = {u_ca_out_771[3:0], u_ca_out_770[7:4]};
assign col_out_772 = {u_ca_out_772[3:0], u_ca_out_771[7:4]};
assign col_out_773 = {u_ca_out_773[3:0], u_ca_out_772[7:4]};
assign col_out_774 = {u_ca_out_774[3:0], u_ca_out_773[7:4]};
assign col_out_775 = {u_ca_out_775[3:0], u_ca_out_774[7:4]};
assign col_out_776 = {u_ca_out_776[3:0], u_ca_out_775[7:4]};
assign col_out_777 = {u_ca_out_777[3:0], u_ca_out_776[7:4]};
assign col_out_778 = {u_ca_out_778[3:0], u_ca_out_777[7:4]};
assign col_out_779 = {u_ca_out_779[3:0], u_ca_out_778[7:4]};
assign col_out_780 = {u_ca_out_780[3:0], u_ca_out_779[7:4]};
assign col_out_781 = {u_ca_out_781[3:0], u_ca_out_780[7:4]};
assign col_out_782 = {u_ca_out_782[3:0], u_ca_out_781[7:4]};
assign col_out_783 = {u_ca_out_783[3:0], u_ca_out_782[7:4]};
assign col_out_784 = {u_ca_out_784[3:0], u_ca_out_783[7:4]};
assign col_out_785 = {u_ca_out_785[3:0], u_ca_out_784[7:4]};
assign col_out_786 = {u_ca_out_786[3:0], u_ca_out_785[7:4]};
assign col_out_787 = {u_ca_out_787[3:0], u_ca_out_786[7:4]};
assign col_out_788 = {u_ca_out_788[3:0], u_ca_out_787[7:4]};
assign col_out_789 = {u_ca_out_789[3:0], u_ca_out_788[7:4]};
assign col_out_790 = {u_ca_out_790[3:0], u_ca_out_789[7:4]};
assign col_out_791 = {u_ca_out_791[3:0], u_ca_out_790[7:4]};
assign col_out_792 = {u_ca_out_792[3:0], u_ca_out_791[7:4]};
assign col_out_793 = {u_ca_out_793[3:0], u_ca_out_792[7:4]};
assign col_out_794 = {u_ca_out_794[3:0], u_ca_out_793[7:4]};
assign col_out_795 = {u_ca_out_795[3:0], u_ca_out_794[7:4]};
assign col_out_796 = {u_ca_out_796[3:0], u_ca_out_795[7:4]};
assign col_out_797 = {u_ca_out_797[3:0], u_ca_out_796[7:4]};
assign col_out_798 = {u_ca_out_798[3:0], u_ca_out_797[7:4]};
assign col_out_799 = {u_ca_out_799[3:0], u_ca_out_798[7:4]};
assign col_out_800 = {u_ca_out_800[3:0], u_ca_out_799[7:4]};
assign col_out_801 = {u_ca_out_801[3:0], u_ca_out_800[7:4]};
assign col_out_802 = {u_ca_out_802[3:0], u_ca_out_801[7:4]};
assign col_out_803 = {u_ca_out_803[3:0], u_ca_out_802[7:4]};
assign col_out_804 = {u_ca_out_804[3:0], u_ca_out_803[7:4]};
assign col_out_805 = {u_ca_out_805[3:0], u_ca_out_804[7:4]};
assign col_out_806 = {u_ca_out_806[3:0], u_ca_out_805[7:4]};
assign col_out_807 = {u_ca_out_807[3:0], u_ca_out_806[7:4]};
assign col_out_808 = {u_ca_out_808[3:0], u_ca_out_807[7:4]};
assign col_out_809 = {u_ca_out_809[3:0], u_ca_out_808[7:4]};
assign col_out_810 = {u_ca_out_810[3:0], u_ca_out_809[7:4]};
assign col_out_811 = {u_ca_out_811[3:0], u_ca_out_810[7:4]};
assign col_out_812 = {u_ca_out_812[3:0], u_ca_out_811[7:4]};
assign col_out_813 = {u_ca_out_813[3:0], u_ca_out_812[7:4]};
assign col_out_814 = {u_ca_out_814[3:0], u_ca_out_813[7:4]};
assign col_out_815 = {u_ca_out_815[3:0], u_ca_out_814[7:4]};
assign col_out_816 = {u_ca_out_816[3:0], u_ca_out_815[7:4]};
assign col_out_817 = {u_ca_out_817[3:0], u_ca_out_816[7:4]};
assign col_out_818 = {u_ca_out_818[3:0], u_ca_out_817[7:4]};
assign col_out_819 = {u_ca_out_819[3:0], u_ca_out_818[7:4]};
assign col_out_820 = {u_ca_out_820[3:0], u_ca_out_819[7:4]};
assign col_out_821 = {u_ca_out_821[3:0], u_ca_out_820[7:4]};
assign col_out_822 = {u_ca_out_822[3:0], u_ca_out_821[7:4]};
assign col_out_823 = {u_ca_out_823[3:0], u_ca_out_822[7:4]};
assign col_out_824 = {u_ca_out_824[3:0], u_ca_out_823[7:4]};
assign col_out_825 = {u_ca_out_825[3:0], u_ca_out_824[7:4]};
assign col_out_826 = {u_ca_out_826[3:0], u_ca_out_825[7:4]};
assign col_out_827 = {u_ca_out_827[3:0], u_ca_out_826[7:4]};
assign col_out_828 = {u_ca_out_828[3:0], u_ca_out_827[7:4]};
assign col_out_829 = {u_ca_out_829[3:0], u_ca_out_828[7:4]};
assign col_out_830 = {u_ca_out_830[3:0], u_ca_out_829[7:4]};
assign col_out_831 = {u_ca_out_831[3:0], u_ca_out_830[7:4]};
assign col_out_832 = {u_ca_out_832[3:0], u_ca_out_831[7:4]};
assign col_out_833 = {u_ca_out_833[3:0], u_ca_out_832[7:4]};
assign col_out_834 = {u_ca_out_834[3:0], u_ca_out_833[7:4]};
assign col_out_835 = {u_ca_out_835[3:0], u_ca_out_834[7:4]};
assign col_out_836 = {u_ca_out_836[3:0], u_ca_out_835[7:4]};
assign col_out_837 = {u_ca_out_837[3:0], u_ca_out_836[7:4]};
assign col_out_838 = {u_ca_out_838[3:0], u_ca_out_837[7:4]};
assign col_out_839 = {u_ca_out_839[3:0], u_ca_out_838[7:4]};
assign col_out_840 = {u_ca_out_840[3:0], u_ca_out_839[7:4]};
assign col_out_841 = {u_ca_out_841[3:0], u_ca_out_840[7:4]};
assign col_out_842 = {u_ca_out_842[3:0], u_ca_out_841[7:4]};
assign col_out_843 = {u_ca_out_843[3:0], u_ca_out_842[7:4]};
assign col_out_844 = {u_ca_out_844[3:0], u_ca_out_843[7:4]};
assign col_out_845 = {u_ca_out_845[3:0], u_ca_out_844[7:4]};
assign col_out_846 = {u_ca_out_846[3:0], u_ca_out_845[7:4]};
assign col_out_847 = {u_ca_out_847[3:0], u_ca_out_846[7:4]};
assign col_out_848 = {u_ca_out_848[3:0], u_ca_out_847[7:4]};
assign col_out_849 = {u_ca_out_849[3:0], u_ca_out_848[7:4]};
assign col_out_850 = {u_ca_out_850[3:0], u_ca_out_849[7:4]};
assign col_out_851 = {u_ca_out_851[3:0], u_ca_out_850[7:4]};
assign col_out_852 = {u_ca_out_852[3:0], u_ca_out_851[7:4]};
assign col_out_853 = {u_ca_out_853[3:0], u_ca_out_852[7:4]};
assign col_out_854 = {u_ca_out_854[3:0], u_ca_out_853[7:4]};
assign col_out_855 = {u_ca_out_855[3:0], u_ca_out_854[7:4]};
assign col_out_856 = {u_ca_out_856[3:0], u_ca_out_855[7:4]};
assign col_out_857 = {u_ca_out_857[3:0], u_ca_out_856[7:4]};
assign col_out_858 = {u_ca_out_858[3:0], u_ca_out_857[7:4]};
assign col_out_859 = {u_ca_out_859[3:0], u_ca_out_858[7:4]};
assign col_out_860 = {u_ca_out_860[3:0], u_ca_out_859[7:4]};
assign col_out_861 = {u_ca_out_861[3:0], u_ca_out_860[7:4]};
assign col_out_862 = {u_ca_out_862[3:0], u_ca_out_861[7:4]};
assign col_out_863 = {u_ca_out_863[3:0], u_ca_out_862[7:4]};
assign col_out_864 = {u_ca_out_864[3:0], u_ca_out_863[7:4]};
assign col_out_865 = {u_ca_out_865[3:0], u_ca_out_864[7:4]};
assign col_out_866 = {u_ca_out_866[3:0], u_ca_out_865[7:4]};
assign col_out_867 = {u_ca_out_867[3:0], u_ca_out_866[7:4]};
assign col_out_868 = {u_ca_out_868[3:0], u_ca_out_867[7:4]};
assign col_out_869 = {u_ca_out_869[3:0], u_ca_out_868[7:4]};
assign col_out_870 = {u_ca_out_870[3:0], u_ca_out_869[7:4]};
assign col_out_871 = {u_ca_out_871[3:0], u_ca_out_870[7:4]};
assign col_out_872 = {u_ca_out_872[3:0], u_ca_out_871[7:4]};
assign col_out_873 = {u_ca_out_873[3:0], u_ca_out_872[7:4]};
assign col_out_874 = {u_ca_out_874[3:0], u_ca_out_873[7:4]};
assign col_out_875 = {u_ca_out_875[3:0], u_ca_out_874[7:4]};
assign col_out_876 = {u_ca_out_876[3:0], u_ca_out_875[7:4]};
assign col_out_877 = {u_ca_out_877[3:0], u_ca_out_876[7:4]};
assign col_out_878 = {u_ca_out_878[3:0], u_ca_out_877[7:4]};
assign col_out_879 = {u_ca_out_879[3:0], u_ca_out_878[7:4]};
assign col_out_880 = {u_ca_out_880[3:0], u_ca_out_879[7:4]};
assign col_out_881 = {u_ca_out_881[3:0], u_ca_out_880[7:4]};
assign col_out_882 = {u_ca_out_882[3:0], u_ca_out_881[7:4]};
assign col_out_883 = {u_ca_out_883[3:0], u_ca_out_882[7:4]};
assign col_out_884 = {u_ca_out_884[3:0], u_ca_out_883[7:4]};
assign col_out_885 = {u_ca_out_885[3:0], u_ca_out_884[7:4]};
assign col_out_886 = {u_ca_out_886[3:0], u_ca_out_885[7:4]};
assign col_out_887 = {u_ca_out_887[3:0], u_ca_out_886[7:4]};
assign col_out_888 = {u_ca_out_888[3:0], u_ca_out_887[7:4]};
assign col_out_889 = {u_ca_out_889[3:0], u_ca_out_888[7:4]};
assign col_out_890 = {u_ca_out_890[3:0], u_ca_out_889[7:4]};
assign col_out_891 = {u_ca_out_891[3:0], u_ca_out_890[7:4]};
assign col_out_892 = {u_ca_out_892[3:0], u_ca_out_891[7:4]};
assign col_out_893 = {u_ca_out_893[3:0], u_ca_out_892[7:4]};
assign col_out_894 = {u_ca_out_894[3:0], u_ca_out_893[7:4]};
assign col_out_895 = {u_ca_out_895[3:0], u_ca_out_894[7:4]};
assign col_out_896 = {u_ca_out_896[3:0], u_ca_out_895[7:4]};
assign col_out_897 = {u_ca_out_897[3:0], u_ca_out_896[7:4]};
assign col_out_898 = {u_ca_out_898[3:0], u_ca_out_897[7:4]};
assign col_out_899 = {u_ca_out_899[3:0], u_ca_out_898[7:4]};
assign col_out_900 = {u_ca_out_900[3:0], u_ca_out_899[7:4]};
assign col_out_901 = {u_ca_out_901[3:0], u_ca_out_900[7:4]};
assign col_out_902 = {u_ca_out_902[3:0], u_ca_out_901[7:4]};
assign col_out_903 = {u_ca_out_903[3:0], u_ca_out_902[7:4]};
assign col_out_904 = {u_ca_out_904[3:0], u_ca_out_903[7:4]};
assign col_out_905 = {u_ca_out_905[3:0], u_ca_out_904[7:4]};
assign col_out_906 = {u_ca_out_906[3:0], u_ca_out_905[7:4]};
assign col_out_907 = {u_ca_out_907[3:0], u_ca_out_906[7:4]};
assign col_out_908 = {u_ca_out_908[3:0], u_ca_out_907[7:4]};
assign col_out_909 = {u_ca_out_909[3:0], u_ca_out_908[7:4]};
assign col_out_910 = {u_ca_out_910[3:0], u_ca_out_909[7:4]};
assign col_out_911 = {u_ca_out_911[3:0], u_ca_out_910[7:4]};
assign col_out_912 = {u_ca_out_912[3:0], u_ca_out_911[7:4]};
assign col_out_913 = {u_ca_out_913[3:0], u_ca_out_912[7:4]};
assign col_out_914 = {u_ca_out_914[3:0], u_ca_out_913[7:4]};
assign col_out_915 = {u_ca_out_915[3:0], u_ca_out_914[7:4]};
assign col_out_916 = {u_ca_out_916[3:0], u_ca_out_915[7:4]};
assign col_out_917 = {u_ca_out_917[3:0], u_ca_out_916[7:4]};
assign col_out_918 = {u_ca_out_918[3:0], u_ca_out_917[7:4]};
assign col_out_919 = {u_ca_out_919[3:0], u_ca_out_918[7:4]};
assign col_out_920 = {u_ca_out_920[3:0], u_ca_out_919[7:4]};
assign col_out_921 = {u_ca_out_921[3:0], u_ca_out_920[7:4]};
assign col_out_922 = {u_ca_out_922[3:0], u_ca_out_921[7:4]};
assign col_out_923 = {u_ca_out_923[3:0], u_ca_out_922[7:4]};
assign col_out_924 = {u_ca_out_924[3:0], u_ca_out_923[7:4]};
assign col_out_925 = {u_ca_out_925[3:0], u_ca_out_924[7:4]};
assign col_out_926 = {u_ca_out_926[3:0], u_ca_out_925[7:4]};
assign col_out_927 = {u_ca_out_927[3:0], u_ca_out_926[7:4]};
assign col_out_928 = {u_ca_out_928[3:0], u_ca_out_927[7:4]};
assign col_out_929 = {u_ca_out_929[3:0], u_ca_out_928[7:4]};
assign col_out_930 = {u_ca_out_930[3:0], u_ca_out_929[7:4]};
assign col_out_931 = {u_ca_out_931[3:0], u_ca_out_930[7:4]};
assign col_out_932 = {u_ca_out_932[3:0], u_ca_out_931[7:4]};
assign col_out_933 = {u_ca_out_933[3:0], u_ca_out_932[7:4]};
assign col_out_934 = {u_ca_out_934[3:0], u_ca_out_933[7:4]};
assign col_out_935 = {u_ca_out_935[3:0], u_ca_out_934[7:4]};
assign col_out_936 = {u_ca_out_936[3:0], u_ca_out_935[7:4]};
assign col_out_937 = {u_ca_out_937[3:0], u_ca_out_936[7:4]};
assign col_out_938 = {u_ca_out_938[3:0], u_ca_out_937[7:4]};
assign col_out_939 = {u_ca_out_939[3:0], u_ca_out_938[7:4]};
assign col_out_940 = {u_ca_out_940[3:0], u_ca_out_939[7:4]};
assign col_out_941 = {u_ca_out_941[3:0], u_ca_out_940[7:4]};
assign col_out_942 = {u_ca_out_942[3:0], u_ca_out_941[7:4]};
assign col_out_943 = {u_ca_out_943[3:0], u_ca_out_942[7:4]};
assign col_out_944 = {u_ca_out_944[3:0], u_ca_out_943[7:4]};
assign col_out_945 = {u_ca_out_945[3:0], u_ca_out_944[7:4]};
assign col_out_946 = {u_ca_out_946[3:0], u_ca_out_945[7:4]};
assign col_out_947 = {u_ca_out_947[3:0], u_ca_out_946[7:4]};
assign col_out_948 = {u_ca_out_948[3:0], u_ca_out_947[7:4]};
assign col_out_949 = {u_ca_out_949[3:0], u_ca_out_948[7:4]};
assign col_out_950 = {u_ca_out_950[3:0], u_ca_out_949[7:4]};
assign col_out_951 = {u_ca_out_951[3:0], u_ca_out_950[7:4]};
assign col_out_952 = {u_ca_out_952[3:0], u_ca_out_951[7:4]};
assign col_out_953 = {u_ca_out_953[3:0], u_ca_out_952[7:4]};
assign col_out_954 = {u_ca_out_954[3:0], u_ca_out_953[7:4]};
assign col_out_955 = {u_ca_out_955[3:0], u_ca_out_954[7:4]};
assign col_out_956 = {u_ca_out_956[3:0], u_ca_out_955[7:4]};
assign col_out_957 = {u_ca_out_957[3:0], u_ca_out_956[7:4]};
assign col_out_958 = {u_ca_out_958[3:0], u_ca_out_957[7:4]};
assign col_out_959 = {u_ca_out_959[3:0], u_ca_out_958[7:4]};
assign col_out_960 = {u_ca_out_960[3:0], u_ca_out_959[7:4]};
assign col_out_961 = {u_ca_out_961[3:0], u_ca_out_960[7:4]};
assign col_out_962 = {u_ca_out_962[3:0], u_ca_out_961[7:4]};
assign col_out_963 = {u_ca_out_963[3:0], u_ca_out_962[7:4]};
assign col_out_964 = {u_ca_out_964[3:0], u_ca_out_963[7:4]};
assign col_out_965 = {u_ca_out_965[3:0], u_ca_out_964[7:4]};
assign col_out_966 = {u_ca_out_966[3:0], u_ca_out_965[7:4]};
assign col_out_967 = {u_ca_out_967[3:0], u_ca_out_966[7:4]};
assign col_out_968 = {u_ca_out_968[3:0], u_ca_out_967[7:4]};
assign col_out_969 = {u_ca_out_969[3:0], u_ca_out_968[7:4]};
assign col_out_970 = {u_ca_out_970[3:0], u_ca_out_969[7:4]};
assign col_out_971 = {u_ca_out_971[3:0], u_ca_out_970[7:4]};
assign col_out_972 = {u_ca_out_972[3:0], u_ca_out_971[7:4]};
assign col_out_973 = {u_ca_out_973[3:0], u_ca_out_972[7:4]};
assign col_out_974 = {u_ca_out_974[3:0], u_ca_out_973[7:4]};
assign col_out_975 = {u_ca_out_975[3:0], u_ca_out_974[7:4]};
assign col_out_976 = {u_ca_out_976[3:0], u_ca_out_975[7:4]};
assign col_out_977 = {u_ca_out_977[3:0], u_ca_out_976[7:4]};
assign col_out_978 = {u_ca_out_978[3:0], u_ca_out_977[7:4]};
assign col_out_979 = {u_ca_out_979[3:0], u_ca_out_978[7:4]};
assign col_out_980 = {u_ca_out_980[3:0], u_ca_out_979[7:4]};
assign col_out_981 = {u_ca_out_981[3:0], u_ca_out_980[7:4]};
assign col_out_982 = {u_ca_out_982[3:0], u_ca_out_981[7:4]};
assign col_out_983 = {u_ca_out_983[3:0], u_ca_out_982[7:4]};
assign col_out_984 = {u_ca_out_984[3:0], u_ca_out_983[7:4]};
assign col_out_985 = {u_ca_out_985[3:0], u_ca_out_984[7:4]};
assign col_out_986 = {u_ca_out_986[3:0], u_ca_out_985[7:4]};
assign col_out_987 = {u_ca_out_987[3:0], u_ca_out_986[7:4]};
assign col_out_988 = {u_ca_out_988[3:0], u_ca_out_987[7:4]};
assign col_out_989 = {u_ca_out_989[3:0], u_ca_out_988[7:4]};
assign col_out_990 = {u_ca_out_990[3:0], u_ca_out_989[7:4]};
assign col_out_991 = {u_ca_out_991[3:0], u_ca_out_990[7:4]};
assign col_out_992 = {u_ca_out_992[3:0], u_ca_out_991[7:4]};
assign col_out_993 = {u_ca_out_993[3:0], u_ca_out_992[7:4]};
assign col_out_994 = {u_ca_out_994[3:0], u_ca_out_993[7:4]};
assign col_out_995 = {u_ca_out_995[3:0], u_ca_out_994[7:4]};
assign col_out_996 = {u_ca_out_996[3:0], u_ca_out_995[7:4]};
assign col_out_997 = {u_ca_out_997[3:0], u_ca_out_996[7:4]};
assign col_out_998 = {u_ca_out_998[3:0], u_ca_out_997[7:4]};
assign col_out_999 = {u_ca_out_999[3:0], u_ca_out_998[7:4]};
assign col_out_1000 = {u_ca_out_1000[3:0], u_ca_out_999[7:4]};
assign col_out_1001 = {u_ca_out_1001[3:0], u_ca_out_1000[7:4]};
assign col_out_1002 = {u_ca_out_1002[3:0], u_ca_out_1001[7:4]};
assign col_out_1003 = {u_ca_out_1003[3:0], u_ca_out_1002[7:4]};
assign col_out_1004 = {u_ca_out_1004[3:0], u_ca_out_1003[7:4]};
assign col_out_1005 = {u_ca_out_1005[3:0], u_ca_out_1004[7:4]};
assign col_out_1006 = {u_ca_out_1006[3:0], u_ca_out_1005[7:4]};
assign col_out_1007 = {u_ca_out_1007[3:0], u_ca_out_1006[7:4]};
assign col_out_1008 = {u_ca_out_1008[3:0], u_ca_out_1007[7:4]};
assign col_out_1009 = {u_ca_out_1009[3:0], u_ca_out_1008[7:4]};
assign col_out_1010 = {u_ca_out_1010[3:0], u_ca_out_1009[7:4]};
assign col_out_1011 = {u_ca_out_1011[3:0], u_ca_out_1010[7:4]};
assign col_out_1012 = {u_ca_out_1012[3:0], u_ca_out_1011[7:4]};
assign col_out_1013 = {u_ca_out_1013[3:0], u_ca_out_1012[7:4]};
assign col_out_1014 = {u_ca_out_1014[3:0], u_ca_out_1013[7:4]};
assign col_out_1015 = {u_ca_out_1015[3:0], u_ca_out_1014[7:4]};
assign col_out_1016 = {u_ca_out_1016[3:0], u_ca_out_1015[7:4]};
assign col_out_1017 = {u_ca_out_1017[3:0], u_ca_out_1016[7:4]};
assign col_out_1018 = {u_ca_out_1018[3:0], u_ca_out_1017[7:4]};
assign col_out_1019 = {u_ca_out_1019[3:0], u_ca_out_1018[7:4]};
assign col_out_1020 = {u_ca_out_1020[3:0], u_ca_out_1019[7:4]};
assign col_out_1021 = {u_ca_out_1021[3:0], u_ca_out_1020[7:4]};
assign col_out_1022 = {u_ca_out_1022[3:0], u_ca_out_1021[7:4]};
assign col_out_1023 = {u_ca_out_1023[3:0], u_ca_out_1022[7:4]};
assign col_out_1024 = {u_ca_out_1024[3:0], u_ca_out_1023[7:4]};
assign col_out_1025 = {u_ca_out_1025[3:0], u_ca_out_1024[7:4]};
assign col_out_1026 = {u_ca_out_1026[3:0], u_ca_out_1025[7:4]};
assign col_out_1027 = {u_ca_out_1027[3:0], u_ca_out_1026[7:4]};
assign col_out_1028 = {u_ca_out_1028[3:0], u_ca_out_1027[7:4]};
assign col_out_1029 = {u_ca_out_1029[3:0], u_ca_out_1028[7:4]};
assign col_out_1030 = {u_ca_out_1030[3:0], u_ca_out_1029[7:4]};
assign col_out_1031 = {u_ca_out_1031[3:0], u_ca_out_1030[7:4]};
assign col_out_1032 = {u_ca_out_1032[3:0], u_ca_out_1031[7:4]};
assign col_out_1033 = {{4{1'b0}}, u_ca_out_1032[7:4]};

//---------------------------------------------------------


endmodule
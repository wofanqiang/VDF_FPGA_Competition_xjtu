module xpb_5_1005
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h518f188dc3bcc74e2b05350b884a5649b59b189f07cda47ef7705247e9530f7ad78e543b872a7925d038e47efd60c00c8a63b9b0112fb17789d3d48b0e4d902ef112329e4578cd5e1af4a929bd3c7199f8999c5d7db6c96b6b13f02de8ad5d25ac40a240be5dd29488137ab96686d77be86f7e22c48461b7a18bcd943dbf9d67;
    5'b00010 : xpb = 1024'ha31e311b87798e9c560a6a171094ac936b36313e0f9b48fdeee0a48fd2a61ef5af1ca8770e54f24ba071c8fdfac1801914c77360225f62ef13a7a9161c9b205de224653c8af19abc35e952537a78e333f13338bafb6d92d6d627e05bd15aba4b588144817cbba5291026f572cd0daef7d0defc458908c36f43179b287b7f3ace;
    5'b00011 : xpb = 1024'h4400045389482121b60a274b8884bb8baf5b46ac41f14d0568743d8208f6816883627f39cb58ece2d14c6e3614c42f5b3b11052a10dc441aecdc3e42f0163bdb5ee7632c20d96ad53e43f8da9ed9909cf5c7db7fec9e2f318baf3e8effdd74ded5ba54988a507f30117a894d3bc4604a6a749b85fd41c7f69e33edb8305c71ca;
    5'b00100 : xpb = 1024'h958f1ce14d04e86fe10f5c5710cf11d564f65f4b49bef1845fe48fc9f24990e35af0d37552836608a18552b51224ef67c574beda220bf59276b012cdfe63cc0a4ff995ca665238335938a2045c160236ee6177dd6a54f89cf6c32ebce88ad20481faf6d948ae51c4998e0406a24b37c652e419a8c1c629ae3fbfbb4c6e1c0f31;
    5'b00101 : xpb = 1024'h3670f0194ed37af5410f198b88bf20cda91b74b97c14f58bd97828bc2899f3562f36aa380f87609fd25ff7ed2c279ea9ebbe50a41088d6be4fe4a7fad1dee787ccbc93b9fc3a084c6193488b8076af9ff2f61aa25b8594f7ac4a8cf0170d8c97ff3406f056432bcb9ae197e11101e918ec79b8e935ff2e359adc0ddc22f9462d;
    5'b00110 : xpb = 1024'h880008a7129042436c144e97110977175eb68d5883e29a0ad0e87b0411ed02d106c4fe7396b1d9c5a298dc6c29885eb676220a5421b88835d9b87c85e02c77b6bdcec65841b2d5aa7c87f1b53db32139eb8fb6ffd93c5e63175e7d1dffbae9bdab74a93114a0fe6022f5129a7788c094d4e9370bfa838fed3c67db7060b8e394;
    5'b00111 : xpb = 1024'h28e1dbdf145ed4c8cc140bcb88f9860fa2dba2c6b6389e124a7c13f6483d6543db0ad53653b5d45cd37381a4438b0df89c6b9c1e10356961b2ed11b2b3a793343a91c447d79aa5c384e2983c6213cea2f02459c4ca6cfabdcce5db512e3da45128adb9482235d8672448a674e63f71e76e7ed64c6ebc947497842e0015961a90;
    5'b01000 : xpb = 1024'h7a70f46cd81b9c16f71940d71143dc595876bb65be06429141ec663e319074beb2992971dae04d82a3ac662340ebce0526cf55ce21651ad93cc0e63dc1f523632ba3f6e61d1373219fd741661f50403ce8bdf6224823c42937f9cb7f16eb0176d4ee5b88e093aafbac5c212e4cc6496356ee546f3340f62c390ffb945355b7f7;
    5'b01001 : xpb = 1024'h1b52c7a4d9ea2e9c5718fe0b8933eb519c9bd0d3f05c4698bb7fff3067e0d73186df003497e44819d4870b5b5aee7d474d18e7980fe1fc0515f57b6a95703ee0a866f4d5b2fb433aa831e7ed43b0eda5ed5298e739546083ed8129b2456dbc0a52276b9fee288502adafb508bb7cfab5f083f3afa779fab3942c4e240832eef3;
    5'b01010 : xpb = 1024'h6ce1e0329da6f5ea821e3317117e419b5236e972f829eb17b2f051785133e6ac5e6d54701f0ec13fa4bfefda584f3d53d77ca1482111ad7c9fc94ff5a3bdcf0f99792773f8741098c326911700ed5f3fe5ec3544b70b29ef589519e02e1b192ffe680de0ac86579735c32fc22203d231d8f371d26bfe5c6b35b81bb845f28c5a;
    5'b01011 : xpb = 1024'hdc3b36a9f75886fe21df04b896e5093965bfee12a7fef1f2c83ea6a8784491f32b32b32dc12bbd6d59a95127251ec95fdc633120f8e8ea878fde5227738ea8d163c25638e5be0b1cb81379e254e0ca8ea80d809a83bc64a0e1c78135c9dd3c37ba11df7ba1b319e3716c39c90ba838472891112e03760f290d46e47facfc356;
    5'b01100 : xpb = 1024'h5f52cbf863324fbe0d23255711b8a6dd4bf71780324d939e23f43cb270d7589a0a417f6e633d34fca5d379916fb2aca28829ecc220be402002d1b9ad85867abc074e5801d3d4ae0fe675e0c7e28a7e42e31a746725f28fb579306841454b30e927e1c03878790432bf2a3e55f7415b005af88f35a4bbc2aa32603bdc388f60bd;
    5'b01101 : xpb = 1024'h349f306500e2436d22e28b89a8b5d5901c2cee64a397a59d87d5a4a727bb0cde87563120412f93d6ae1ec989b55be4ae737e8c0f3b214bdc064eda59019639841155f169bc7e28eed0874f06eb2babe7af172c17232c102eb7c67473cdeb7ca51ad04f860dde39c07dd23065f80c52f48e2e7618f4c7318d7c8e6bed6c97b9;
    5'b01110 : xpb = 1024'h51c3b7be28bda9919828179711f30c1f45b7458d6c713c2494f827ec907aca87b615aa6ca76ba8b9a6e7034887161bf138d7383c206ad2c365da2365674f26687523888faf354b8709c53078c4279d45e048b38994d9f57b99cbb6a25c7b48a2515b7290446bb0ce48914ce9cc7ee3cedcfdac98dd7928e92f085c002b2c3520;
    5'b01111 : xpb = 1024'ha352d04bec7a70dfc32d4ca29a3d6268fb525e2c743ee0a38c687a3479cdda028da3fea82e9621df771fe7c78476dbfdc33af1ec319a843aefadf7f0759cb6976635bb2df4ae18e524b9d9a281640edfd8e24fe71290bee704dfa6d04528a5c7fd9c14d102c98362d0a4c7a33305bb4ac56d2abba1fd8aa0d094299468ebd287;
    5'b10000 : xpb = 1024'h4434a383ee490365232d09d7122d71613f77739aa694e4ab05fc1326b01e3c7561e9d56aeb9a1c76a7fa8cff9e798b3fe98483b620176566c8e28d1d4917d214e2f8b91d8a95e8fe2d148029a5c4bc48dd76f2ac03c15b41ba67050373ab605b7ad524e8105e5d69d1f85b7da1bc6c9d5f02c9fc16368f282bb07c241dc90983;
    5'b10001 : xpb = 1024'h95c3bc11b205cab34e323ee29a77c7aaf5128c39ae628929fd6c656e99714bf0397829a672c4959c7833717e9bda4b4c73e83d66314716de52b661a857656243d40aebbbd00eb65c4809295363012de2d6108f09817824ad257af5315c58bd812715c728cebc2ffe5a0bd637084344194772481edabaf0dfcd3c49b85b88a6ea;
    5'b10010 : xpb = 1024'h36a58f49b3d45d38ae31fc171267d6a33937a1a7e0b88d3176fffe60cfc1ae630dbe00692fc89033a90e16b6b5dcfa8e9a31cf301fc3f80a2beaf6d52ae07dc150cde9ab65f686755063cfda8761db4bdaa531ce72a8c107db0253648adb7814a44ed73fdc510a055b5f6a1176f9f56be107e75f4ef3f56728589c481065dde6;
    5'b10011 : xpb = 1024'h8834a7d777912486d93731229ab22ceceed2ba46e88631b06e7050a8b914bddde54c54a4b6f309597946fb35b33dba9b249588e030f3a981b5becb60392e0df041e01c49ab6f53d36b587904449e4ce5d33ece2bf05f8a73461643927388d53a508f79809aaedc99e372e4cadd80cce7c97765821378571ec9e469dc4e257b4d;
    5'b10100 : xpb = 1024'h29167b0f795fb70c3936ee5712a23be532f7cfb51adc35b7e803e99aef652050b9922b6773f703f0aa21a06dcd4069dd4adf1aaa1f708aad8ef3608d0ca9296dbea31a39415723ec73b31f8b68fefa4ed7d370f0e19026cdfb9da1c5a20b8fcdcdc88997a843b6a0e4c678a54c377e3a630d04c287b15ba62500bc6c0302b249;
    5'b10101 : xpb = 1024'h7aa5939d3d1c7e5a643c23629aec922ee892e85422a9da36df743be2d8b82fcb91207fa2fb217d167a5a84eccaa129e9d542d45a30a03c2518c735181af6b99cafb54cd786cff14a8ea7c8b5263b6be8d06d0d4e5f46f03966b191f38ab8ecf37a092bd866a189356cd9f35eb2be55b64b7c82e54c35bd5dc68c8a0040c24fb0;
    5'b10110 : xpb = 1024'h1b8766d53eeb10dfc43be09712dca1272cb7fdc254ffde3e5907d4d50f08923e65665665b82577adab352a24e4a3d92bfb8c66241f1d1d50f1fbca44ee71d51a2c784ac71cb7c16397026f3c4a9c1951d501b01350778c941c38f026b93ba786f7423bef7436633c6e2d873921750708e5122225c06ec1e521a8dc8ff59f86ac;
    5'b10111 : xpb = 1024'h6d167f6302a7d82def4115a29b26f770e25316615ccd82bd5078271cf85ba1b93cf4aaa13f4ff0d37b6e0ea3e204993885f01fd4304ccec87bcf9ecffcbf65491d8a7d6562308ec1b1f7186607d88aebcd9b4c70ce2e55ff874ce054a1e904aca382de30329435d0f64101f287fbde84cd81a04884f3239cc334aa24335f2413;
    5'b11000 : xpb = 1024'hdf8529b04766ab34f40d2d71317066926782bcf8f2386c4ca0bc00f2eac042c113a8163fc53eb6aac48b3dbfc07487aac39b19e1ec9aff4550433fcd03a80c69a4d7b54f8185edaba51beed2c393854d22fef35bf5ef25a3cd43e87d06bbf4020bbee4740290fd7f79495ccf6b28fd767173f88f92c28241e50fcb3e83c5b0f;
    5'b11001 : xpb = 1024'h5f876b28c83332017a4607e29b615cb2dc13446e96f12b43c17c125717ff13a6e8c8d59f837e64907c81985af9680887369d6b4e2ff9616bded80887de8810f58b5fadf33d912c38d5466816e975a9eecac98b933d15bbc5a7e82eb5b9191c65ccfc9087fe86e26c7fa810865d3967534f86bdabbdb089dbbfdcca4825fbf876;
    5'b11010 : xpb = 1024'h693e60ca01c486da45c51713516bab203859dcc9472f4b3b0fab494e4f7619bd0eac6240825f27ad5c3d93136ab7c95ce6fd181e764297b80c9db4b2032c730822abe2d378fc51dda10e9e0dd65757cf5e2e582e4658205d6f8ce8e79bd6f94a35a09f0c1bbc7380fba460cbf018a5e91c5cec31e98e631af91cd7dad92f72;
    5'b11011 : xpb = 1024'h51f856ee8dbe8bd5054afa229b9bc1f4d5d3727bd114d3ca327ffd9137a28594949d009dc7acd84d7d95221210cb77d5e74ab6c82fa5f40f41e0723fc050bca1f934de8118f1c9aff895b7c7cb12c8f1c7f7cab5abfd218bc8837d16d049341ef67642dfca798f08090f1f1a3276f021d18bdb0ef66df01abc84ea6c1898ccd9;
    5'b11100 : xpb = 1024'ha3876f7c517b532330502f2e23e6183e8b6e8b1ad8e2784929f04fd920f5950f6c2b54d94ed751734dce06910e2c37e271ae707840d5a586cbb446cace9e4cd0ea47111f5e6a970e138a60f1884f3a8bc091671329b3eaf733976d44b8f69144a2b6e52088d7619c912299d398fdc79db9fb5931baf251d25e10b80056586a40;
    5'b11101 : xpb = 1024'h446942b45349e5a8904fec629bd62736cf93a0890b387c50a383e8cb5745f78240712b9c0bdb4c0a7ea8abc9282ee72497f802422f5286b2a4e8dbf7a219684e670a0f0ef45267271be50778acafe7f4c52609d81ae48751e91ecb77e7794bd81feff537966c3ba392762dae07b478f05390f8722f2b5659b92d0a900b35a13c;
    5'b11110 : xpb = 1024'h95f85b421706acf6bb55216e24207d80852eb928130620cf9af43b13409906fd17ff7fd79305c5304ee19048258fa731225bbbf24082382a2ebcb082b066f87d581c41ad39cb348536d9b0a269ec598ebdbfa635989b50bd5432bba5d026a8fdcc30977854ca0e381a89a8676e3b506c3c007694f3afb8115ab8d82448f53ea3;
    5'b11111 : xpb = 1024'h36da2e7a18d53f7c1b54dea29c108c78c953ce96455c24d71487d40576e9696fec45569a5009bfc77fbc35803f92567348a54dbc2eff195607f145af83e213fad4df3f9ccfb3049e3f3457298e4d06f7c25448fa89cbed1809ba19d8fea963914969a78f625ee83f1bdd3c41dcf201bed59615d567e8bc98b5d52ab3fdd2759f;
    endcase
end

endmodule

module  modular_square_iterative
(
    input clk,
    input rst,

    input [1023:0] a,
    input start_ms,

    output [1023:0] ms,
    output finish_ms
);


localparam IDLE             = 6'b000001;
localparam TRANS_DATA       = 6'b000010;
localparam COMPRESS_HIGH    = 6'b000100;
localparam COMPRESS_LOW     = 6'b001000;
localparam REDUCTION        = 6'b010000;
localparam FINISH           = 6'b100000;





localparam P1 = 1026'hb0ad4555c1ee34c8cb0577d7105a475171760330d577a0777ddcb955b302ad0803487d78ca267e8e9f5e3f46e35e10ca641a27e622b2d04bb09f3f5e3ad274b1744f34aeaf90fd45129a02a298dbc430f404f9988c862d10b58c91faba2aa2922f079229b0c8f88d86bfe6def7d026294ed9dee2504b5d30466f7b0488e2666b;

localparam P2 = 1026'h1615a8aab83dc6991960aefae20b48ea2e2ec0661aaef40eefbb972ab66055a100690faf1944cfd1d3ebc7e8dc6bc2194c8344fcc4565a097613e7ebc75a4e962e89e695d5f21fa8a2534054531b78861e809f331190c5a216b1923f5745545245e0f24536191f11b0d7fcdbdefa04c529db3bdc4a096ba608cdef60911c4ccd6;

localparam P3 = 1026'h21207d00145ca9e5a61106785310ed5f4546209928066e16679962c011908071809d9786a5e737babde1abdd4aa1a325f2c4e77b2681870e311ddbe1ab0775e145ced9e0c0eb2f7cf37ce07e7ca934c92dc0eecc9a592873220a5b5f02e7fe7b68d16b67d125ae9a8943fb49ce770727bec8d9ca6f0e21790d34e710d9aa73341;

localparam LOOPS = 31'd1073741824;



wire [1026:0] temp_ms0;
wire [1026:0] temp_ms1;
wire [1026:0] temp_ms2;
wire [1026:0] temp_ms3;

reg [1023:0] temp_ms;

reg [1023:0] reg_a;
reg [30:0] counter;
reg reg_start_ms;

reg reg_finish_ms;
reg reg_finish_me;


reg   reg_sel_hp;
reg   [1023:0]  reg_partial_product_high0;
reg   [1023:0]  reg_partial_product_high1;
reg   [1032:0]  reg_partial_product_low0;
reg   [1032:0]  reg_partial_product_low1;
reg   reg_sel_data_in;

reg   [1024:0]  reg_data_out0;
reg   [1024:0]  reg_data_out1;

// data_in_mux Inputs
wire   sel_hp;
wire   [1023:0]  partial_product_high0;
wire   [1023:0]  partial_product_high1;
wire   [1032:0]  partial_product_low0;
wire   [1032:0]  partial_product_low1;
wire   sel_data_in;

assign   sel_hp = reg_sel_hp;
assign   partial_product_high0 = reg_partial_product_high0;
assign   partial_product_high1 = reg_partial_product_high1;
assign   partial_product_low0 = reg_partial_product_low0;
assign   partial_product_low1 = reg_partial_product_low1;
assign   sel_data_in = reg_sel_data_in;


// data_in_mux Outputs
wire  [511:0]  col_out_0;
wire  [511:0]  col_out_1;
wire  [511:0]  col_out_2;
wire  [511:0]  col_out_3;
wire  [511:0]  col_out_4;
wire  [511:0]  col_out_5;
wire  [511:0]  col_out_6;
wire  [511:0]  col_out_7;
wire  [511:0]  col_out_8;
wire  [511:0]  col_out_9;
wire  [511:0]  col_out_10;
wire  [511:0]  col_out_11;
wire  [511:0]  col_out_12;
wire  [511:0]  col_out_13;
wire  [511:0]  col_out_14;
wire  [511:0]  col_out_15;
wire  [511:0]  col_out_16;
wire  [511:0]  col_out_17;
wire  [511:0]  col_out_18;
wire  [511:0]  col_out_19;
wire  [511:0]  col_out_20;
wire  [511:0]  col_out_21;
wire  [511:0]  col_out_22;
wire  [511:0]  col_out_23;
wire  [511:0]  col_out_24;
wire  [511:0]  col_out_25;
wire  [511:0]  col_out_26;
wire  [511:0]  col_out_27;
wire  [511:0]  col_out_28;
wire  [511:0]  col_out_29;
wire  [511:0]  col_out_30;
wire  [511:0]  col_out_31;
wire  [511:0]  col_out_32;
wire  [511:0]  col_out_33;
wire  [511:0]  col_out_34;
wire  [511:0]  col_out_35;
wire  [511:0]  col_out_36;
wire  [511:0]  col_out_37;
wire  [511:0]  col_out_38;
wire  [511:0]  col_out_39;
wire  [511:0]  col_out_40;
wire  [511:0]  col_out_41;
wire  [511:0]  col_out_42;
wire  [511:0]  col_out_43;
wire  [511:0]  col_out_44;
wire  [511:0]  col_out_45;
wire  [511:0]  col_out_46;
wire  [511:0]  col_out_47;
wire  [511:0]  col_out_48;
wire  [511:0]  col_out_49;
wire  [511:0]  col_out_50;
wire  [511:0]  col_out_51;
wire  [511:0]  col_out_52;
wire  [511:0]  col_out_53;
wire  [511:0]  col_out_54;
wire  [511:0]  col_out_55;
wire  [511:0]  col_out_56;
wire  [511:0]  col_out_57;
wire  [511:0]  col_out_58;
wire  [511:0]  col_out_59;
wire  [511:0]  col_out_60;
wire  [511:0]  col_out_61;
wire  [511:0]  col_out_62;
wire  [511:0]  col_out_63;
wire  [511:0]  col_out_64;
wire  [511:0]  col_out_65;
wire  [511:0]  col_out_66;
wire  [511:0]  col_out_67;
wire  [511:0]  col_out_68;
wire  [511:0]  col_out_69;
wire  [511:0]  col_out_70;
wire  [511:0]  col_out_71;
wire  [511:0]  col_out_72;
wire  [511:0]  col_out_73;
wire  [511:0]  col_out_74;
wire  [511:0]  col_out_75;
wire  [511:0]  col_out_76;
wire  [511:0]  col_out_77;
wire  [511:0]  col_out_78;
wire  [511:0]  col_out_79;
wire  [511:0]  col_out_80;
wire  [511:0]  col_out_81;
wire  [511:0]  col_out_82;
wire  [511:0]  col_out_83;
wire  [511:0]  col_out_84;
wire  [511:0]  col_out_85;
wire  [511:0]  col_out_86;
wire  [511:0]  col_out_87;
wire  [511:0]  col_out_88;
wire  [511:0]  col_out_89;
wire  [511:0]  col_out_90;
wire  [511:0]  col_out_91;
wire  [511:0]  col_out_92;
wire  [511:0]  col_out_93;
wire  [511:0]  col_out_94;
wire  [511:0]  col_out_95;
wire  [511:0]  col_out_96;
wire  [511:0]  col_out_97;
wire  [511:0]  col_out_98;
wire  [511:0]  col_out_99;
wire  [511:0]  col_out_100;
wire  [511:0]  col_out_101;
wire  [511:0]  col_out_102;
wire  [511:0]  col_out_103;
wire  [511:0]  col_out_104;
wire  [511:0]  col_out_105;
wire  [511:0]  col_out_106;
wire  [511:0]  col_out_107;
wire  [511:0]  col_out_108;
wire  [511:0]  col_out_109;
wire  [511:0]  col_out_110;
wire  [511:0]  col_out_111;
wire  [511:0]  col_out_112;
wire  [511:0]  col_out_113;
wire  [511:0]  col_out_114;
wire  [511:0]  col_out_115;
wire  [511:0]  col_out_116;
wire  [511:0]  col_out_117;
wire  [511:0]  col_out_118;
wire  [511:0]  col_out_119;
wire  [511:0]  col_out_120;
wire  [511:0]  col_out_121;
wire  [511:0]  col_out_122;
wire  [511:0]  col_out_123;
wire  [511:0]  col_out_124;
wire  [511:0]  col_out_125;
wire  [511:0]  col_out_126;
wire  [511:0]  col_out_127;
wire  [511:0]  col_out_128;
wire  [511:0]  col_out_129;
wire  [511:0]  col_out_130;
wire  [511:0]  col_out_131;
wire  [511:0]  col_out_132;
wire  [511:0]  col_out_133;
wire  [511:0]  col_out_134;
wire  [511:0]  col_out_135;
wire  [511:0]  col_out_136;
wire  [511:0]  col_out_137;
wire  [511:0]  col_out_138;
wire  [511:0]  col_out_139;
wire  [511:0]  col_out_140;
wire  [511:0]  col_out_141;
wire  [511:0]  col_out_142;
wire  [511:0]  col_out_143;
wire  [511:0]  col_out_144;
wire  [511:0]  col_out_145;
wire  [511:0]  col_out_146;
wire  [511:0]  col_out_147;
wire  [511:0]  col_out_148;
wire  [511:0]  col_out_149;
wire  [511:0]  col_out_150;
wire  [511:0]  col_out_151;
wire  [511:0]  col_out_152;
wire  [511:0]  col_out_153;
wire  [511:0]  col_out_154;
wire  [511:0]  col_out_155;
wire  [511:0]  col_out_156;
wire  [511:0]  col_out_157;
wire  [511:0]  col_out_158;
wire  [511:0]  col_out_159;
wire  [511:0]  col_out_160;
wire  [511:0]  col_out_161;
wire  [511:0]  col_out_162;
wire  [511:0]  col_out_163;
wire  [511:0]  col_out_164;
wire  [511:0]  col_out_165;
wire  [511:0]  col_out_166;
wire  [511:0]  col_out_167;
wire  [511:0]  col_out_168;
wire  [511:0]  col_out_169;
wire  [511:0]  col_out_170;
wire  [511:0]  col_out_171;
wire  [511:0]  col_out_172;
wire  [511:0]  col_out_173;
wire  [511:0]  col_out_174;
wire  [511:0]  col_out_175;
wire  [511:0]  col_out_176;
wire  [511:0]  col_out_177;
wire  [511:0]  col_out_178;
wire  [511:0]  col_out_179;
wire  [511:0]  col_out_180;
wire  [511:0]  col_out_181;
wire  [511:0]  col_out_182;
wire  [511:0]  col_out_183;
wire  [511:0]  col_out_184;
wire  [511:0]  col_out_185;
wire  [511:0]  col_out_186;
wire  [511:0]  col_out_187;
wire  [511:0]  col_out_188;
wire  [511:0]  col_out_189;
wire  [511:0]  col_out_190;
wire  [511:0]  col_out_191;
wire  [511:0]  col_out_192;
wire  [511:0]  col_out_193;
wire  [511:0]  col_out_194;
wire  [511:0]  col_out_195;
wire  [511:0]  col_out_196;
wire  [511:0]  col_out_197;
wire  [511:0]  col_out_198;
wire  [511:0]  col_out_199;
wire  [511:0]  col_out_200;
wire  [511:0]  col_out_201;
wire  [511:0]  col_out_202;
wire  [511:0]  col_out_203;
wire  [511:0]  col_out_204;
wire  [511:0]  col_out_205;
wire  [511:0]  col_out_206;
wire  [511:0]  col_out_207;
wire  [511:0]  col_out_208;
wire  [511:0]  col_out_209;
wire  [511:0]  col_out_210;
wire  [511:0]  col_out_211;
wire  [511:0]  col_out_212;
wire  [511:0]  col_out_213;
wire  [511:0]  col_out_214;
wire  [511:0]  col_out_215;
wire  [511:0]  col_out_216;
wire  [511:0]  col_out_217;
wire  [511:0]  col_out_218;
wire  [511:0]  col_out_219;
wire  [511:0]  col_out_220;
wire  [511:0]  col_out_221;
wire  [511:0]  col_out_222;
wire  [511:0]  col_out_223;
wire  [511:0]  col_out_224;
wire  [511:0]  col_out_225;
wire  [511:0]  col_out_226;
wire  [511:0]  col_out_227;
wire  [511:0]  col_out_228;
wire  [511:0]  col_out_229;
wire  [511:0]  col_out_230;
wire  [511:0]  col_out_231;
wire  [511:0]  col_out_232;
wire  [511:0]  col_out_233;
wire  [511:0]  col_out_234;
wire  [511:0]  col_out_235;
wire  [511:0]  col_out_236;
wire  [511:0]  col_out_237;
wire  [511:0]  col_out_238;
wire  [511:0]  col_out_239;
wire  [511:0]  col_out_240;
wire  [511:0]  col_out_241;
wire  [511:0]  col_out_242;
wire  [511:0]  col_out_243;
wire  [511:0]  col_out_244;
wire  [511:0]  col_out_245;
wire  [511:0]  col_out_246;
wire  [511:0]  col_out_247;
wire  [511:0]  col_out_248;
wire  [511:0]  col_out_249;
wire  [511:0]  col_out_250;
wire  [511:0]  col_out_251;
wire  [511:0]  col_out_252;
wire  [511:0]  col_out_253;
wire  [511:0]  col_out_254;
wire  [511:0]  col_out_255;
wire  [511:0]  col_out_256;
wire  [511:0]  col_out_257;
wire  [511:0]  col_out_258;
wire  [511:0]  col_out_259;
wire  [511:0]  col_out_260;
wire  [511:0]  col_out_261;
wire  [511:0]  col_out_262;
wire  [511:0]  col_out_263;
wire  [511:0]  col_out_264;
wire  [511:0]  col_out_265;
wire  [511:0]  col_out_266;
wire  [511:0]  col_out_267;
wire  [511:0]  col_out_268;
wire  [511:0]  col_out_269;
wire  [511:0]  col_out_270;
wire  [511:0]  col_out_271;
wire  [511:0]  col_out_272;
wire  [511:0]  col_out_273;
wire  [511:0]  col_out_274;
wire  [511:0]  col_out_275;
wire  [511:0]  col_out_276;
wire  [511:0]  col_out_277;
wire  [511:0]  col_out_278;
wire  [511:0]  col_out_279;
wire  [511:0]  col_out_280;
wire  [511:0]  col_out_281;
wire  [511:0]  col_out_282;
wire  [511:0]  col_out_283;
wire  [511:0]  col_out_284;
wire  [511:0]  col_out_285;
wire  [511:0]  col_out_286;
wire  [511:0]  col_out_287;
wire  [511:0]  col_out_288;
wire  [511:0]  col_out_289;
wire  [511:0]  col_out_290;
wire  [511:0]  col_out_291;
wire  [511:0]  col_out_292;
wire  [511:0]  col_out_293;
wire  [511:0]  col_out_294;
wire  [511:0]  col_out_295;
wire  [511:0]  col_out_296;
wire  [511:0]  col_out_297;
wire  [511:0]  col_out_298;
wire  [511:0]  col_out_299;
wire  [511:0]  col_out_300;
wire  [511:0]  col_out_301;
wire  [511:0]  col_out_302;
wire  [511:0]  col_out_303;
wire  [511:0]  col_out_304;
wire  [511:0]  col_out_305;
wire  [511:0]  col_out_306;
wire  [511:0]  col_out_307;
wire  [511:0]  col_out_308;
wire  [511:0]  col_out_309;
wire  [511:0]  col_out_310;
wire  [511:0]  col_out_311;
wire  [511:0]  col_out_312;
wire  [511:0]  col_out_313;
wire  [511:0]  col_out_314;
wire  [511:0]  col_out_315;
wire  [511:0]  col_out_316;
wire  [511:0]  col_out_317;
wire  [511:0]  col_out_318;
wire  [511:0]  col_out_319;
wire  [511:0]  col_out_320;
wire  [511:0]  col_out_321;
wire  [511:0]  col_out_322;
wire  [511:0]  col_out_323;
wire  [511:0]  col_out_324;
wire  [511:0]  col_out_325;
wire  [511:0]  col_out_326;
wire  [511:0]  col_out_327;
wire  [511:0]  col_out_328;
wire  [511:0]  col_out_329;
wire  [511:0]  col_out_330;
wire  [511:0]  col_out_331;
wire  [511:0]  col_out_332;
wire  [511:0]  col_out_333;
wire  [511:0]  col_out_334;
wire  [511:0]  col_out_335;
wire  [511:0]  col_out_336;
wire  [511:0]  col_out_337;
wire  [511:0]  col_out_338;
wire  [511:0]  col_out_339;
wire  [511:0]  col_out_340;
wire  [511:0]  col_out_341;
wire  [511:0]  col_out_342;
wire  [511:0]  col_out_343;
wire  [511:0]  col_out_344;
wire  [511:0]  col_out_345;
wire  [511:0]  col_out_346;
wire  [511:0]  col_out_347;
wire  [511:0]  col_out_348;
wire  [511:0]  col_out_349;
wire  [511:0]  col_out_350;
wire  [511:0]  col_out_351;
wire  [511:0]  col_out_352;
wire  [511:0]  col_out_353;
wire  [511:0]  col_out_354;
wire  [511:0]  col_out_355;
wire  [511:0]  col_out_356;
wire  [511:0]  col_out_357;
wire  [511:0]  col_out_358;
wire  [511:0]  col_out_359;
wire  [511:0]  col_out_360;
wire  [511:0]  col_out_361;
wire  [511:0]  col_out_362;
wire  [511:0]  col_out_363;
wire  [511:0]  col_out_364;
wire  [511:0]  col_out_365;
wire  [511:0]  col_out_366;
wire  [511:0]  col_out_367;
wire  [511:0]  col_out_368;
wire  [511:0]  col_out_369;
wire  [511:0]  col_out_370;
wire  [511:0]  col_out_371;
wire  [511:0]  col_out_372;
wire  [511:0]  col_out_373;
wire  [511:0]  col_out_374;
wire  [511:0]  col_out_375;
wire  [511:0]  col_out_376;
wire  [511:0]  col_out_377;
wire  [511:0]  col_out_378;
wire  [511:0]  col_out_379;
wire  [511:0]  col_out_380;
wire  [511:0]  col_out_381;
wire  [511:0]  col_out_382;
wire  [511:0]  col_out_383;
wire  [511:0]  col_out_384;
wire  [511:0]  col_out_385;
wire  [511:0]  col_out_386;
wire  [511:0]  col_out_387;
wire  [511:0]  col_out_388;
wire  [511:0]  col_out_389;
wire  [511:0]  col_out_390;
wire  [511:0]  col_out_391;
wire  [511:0]  col_out_392;
wire  [511:0]  col_out_393;
wire  [511:0]  col_out_394;
wire  [511:0]  col_out_395;
wire  [511:0]  col_out_396;
wire  [511:0]  col_out_397;
wire  [511:0]  col_out_398;
wire  [511:0]  col_out_399;
wire  [511:0]  col_out_400;
wire  [511:0]  col_out_401;
wire  [511:0]  col_out_402;
wire  [511:0]  col_out_403;
wire  [511:0]  col_out_404;
wire  [511:0]  col_out_405;
wire  [511:0]  col_out_406;
wire  [511:0]  col_out_407;
wire  [511:0]  col_out_408;
wire  [511:0]  col_out_409;
wire  [511:0]  col_out_410;
wire  [511:0]  col_out_411;
wire  [511:0]  col_out_412;
wire  [511:0]  col_out_413;
wire  [511:0]  col_out_414;
wire  [511:0]  col_out_415;
wire  [511:0]  col_out_416;
wire  [511:0]  col_out_417;
wire  [511:0]  col_out_418;
wire  [511:0]  col_out_419;
wire  [511:0]  col_out_420;
wire  [511:0]  col_out_421;
wire  [511:0]  col_out_422;
wire  [511:0]  col_out_423;
wire  [511:0]  col_out_424;
wire  [511:0]  col_out_425;
wire  [511:0]  col_out_426;
wire  [511:0]  col_out_427;
wire  [511:0]  col_out_428;
wire  [511:0]  col_out_429;
wire  [511:0]  col_out_430;
wire  [511:0]  col_out_431;
wire  [511:0]  col_out_432;
wire  [511:0]  col_out_433;
wire  [511:0]  col_out_434;
wire  [511:0]  col_out_435;
wire  [511:0]  col_out_436;
wire  [511:0]  col_out_437;
wire  [511:0]  col_out_438;
wire  [511:0]  col_out_439;
wire  [511:0]  col_out_440;
wire  [511:0]  col_out_441;
wire  [511:0]  col_out_442;
wire  [511:0]  col_out_443;
wire  [511:0]  col_out_444;
wire  [511:0]  col_out_445;
wire  [511:0]  col_out_446;
wire  [511:0]  col_out_447;
wire  [511:0]  col_out_448;
wire  [511:0]  col_out_449;
wire  [511:0]  col_out_450;
wire  [511:0]  col_out_451;
wire  [511:0]  col_out_452;
wire  [511:0]  col_out_453;
wire  [511:0]  col_out_454;
wire  [511:0]  col_out_455;
wire  [511:0]  col_out_456;
wire  [511:0]  col_out_457;
wire  [511:0]  col_out_458;
wire  [511:0]  col_out_459;
wire  [511:0]  col_out_460;
wire  [511:0]  col_out_461;
wire  [511:0]  col_out_462;
wire  [511:0]  col_out_463;
wire  [511:0]  col_out_464;
wire  [511:0]  col_out_465;
wire  [511:0]  col_out_466;
wire  [511:0]  col_out_467;
wire  [511:0]  col_out_468;
wire  [511:0]  col_out_469;
wire  [511:0]  col_out_470;
wire  [511:0]  col_out_471;
wire  [511:0]  col_out_472;
wire  [511:0]  col_out_473;
wire  [511:0]  col_out_474;
wire  [511:0]  col_out_475;
wire  [511:0]  col_out_476;
wire  [511:0]  col_out_477;
wire  [511:0]  col_out_478;
wire  [511:0]  col_out_479;
wire  [511:0]  col_out_480;
wire  [511:0]  col_out_481;
wire  [511:0]  col_out_482;
wire  [511:0]  col_out_483;
wire  [511:0]  col_out_484;
wire  [511:0]  col_out_485;
wire  [511:0]  col_out_486;
wire  [511:0]  col_out_487;
wire  [511:0]  col_out_488;
wire  [511:0]  col_out_489;
wire  [511:0]  col_out_490;
wire  [511:0]  col_out_491;
wire  [511:0]  col_out_492;
wire  [511:0]  col_out_493;
wire  [511:0]  col_out_494;
wire  [511:0]  col_out_495;
wire  [511:0]  col_out_496;
wire  [511:0]  col_out_497;
wire  [511:0]  col_out_498;
wire  [511:0]  col_out_499;
wire  [511:0]  col_out_500;
wire  [511:0]  col_out_501;
wire  [511:0]  col_out_502;
wire  [511:0]  col_out_503;
wire  [511:0]  col_out_504;
wire  [511:0]  col_out_505;
wire  [511:0]  col_out_506;
wire  [511:0]  col_out_507;
wire  [511:0]  col_out_508;
wire  [511:0]  col_out_509;
wire  [511:0]  col_out_510;
wire  [511:0]  col_out_511;
wire  [511:0]  col_out_512;
wire  [511:0]  col_out_513;
wire  [511:0]  col_out_514;
wire  [511:0]  col_out_515;
wire  [511:0]  col_out_516;
wire  [511:0]  col_out_517;
wire  [511:0]  col_out_518;
wire  [511:0]  col_out_519;
wire  [511:0]  col_out_520;
wire  [511:0]  col_out_521;
wire  [511:0]  col_out_522;
wire  [511:0]  col_out_523;
wire  [511:0]  col_out_524;
wire  [511:0]  col_out_525;
wire  [511:0]  col_out_526;
wire  [511:0]  col_out_527;
wire  [511:0]  col_out_528;
wire  [511:0]  col_out_529;
wire  [511:0]  col_out_530;
wire  [511:0]  col_out_531;
wire  [511:0]  col_out_532;
wire  [511:0]  col_out_533;
wire  [511:0]  col_out_534;
wire  [511:0]  col_out_535;
wire  [511:0]  col_out_536;
wire  [511:0]  col_out_537;
wire  [511:0]  col_out_538;
wire  [511:0]  col_out_539;
wire  [511:0]  col_out_540;
wire  [511:0]  col_out_541;
wire  [511:0]  col_out_542;
wire  [511:0]  col_out_543;
wire  [511:0]  col_out_544;
wire  [511:0]  col_out_545;
wire  [511:0]  col_out_546;
wire  [511:0]  col_out_547;
wire  [511:0]  col_out_548;
wire  [511:0]  col_out_549;
wire  [511:0]  col_out_550;
wire  [511:0]  col_out_551;
wire  [511:0]  col_out_552;
wire  [511:0]  col_out_553;
wire  [511:0]  col_out_554;
wire  [511:0]  col_out_555;
wire  [511:0]  col_out_556;
wire  [511:0]  col_out_557;
wire  [511:0]  col_out_558;
wire  [511:0]  col_out_559;
wire  [511:0]  col_out_560;
wire  [511:0]  col_out_561;
wire  [511:0]  col_out_562;
wire  [511:0]  col_out_563;
wire  [511:0]  col_out_564;
wire  [511:0]  col_out_565;
wire  [511:0]  col_out_566;
wire  [511:0]  col_out_567;
wire  [511:0]  col_out_568;
wire  [511:0]  col_out_569;
wire  [511:0]  col_out_570;
wire  [511:0]  col_out_571;
wire  [511:0]  col_out_572;
wire  [511:0]  col_out_573;
wire  [511:0]  col_out_574;
wire  [511:0]  col_out_575;
wire  [511:0]  col_out_576;
wire  [511:0]  col_out_577;
wire  [511:0]  col_out_578;
wire  [511:0]  col_out_579;
wire  [511:0]  col_out_580;
wire  [511:0]  col_out_581;
wire  [511:0]  col_out_582;
wire  [511:0]  col_out_583;
wire  [511:0]  col_out_584;
wire  [511:0]  col_out_585;
wire  [511:0]  col_out_586;
wire  [511:0]  col_out_587;
wire  [511:0]  col_out_588;
wire  [511:0]  col_out_589;
wire  [511:0]  col_out_590;
wire  [511:0]  col_out_591;
wire  [511:0]  col_out_592;
wire  [511:0]  col_out_593;
wire  [511:0]  col_out_594;
wire  [511:0]  col_out_595;
wire  [511:0]  col_out_596;
wire  [511:0]  col_out_597;
wire  [511:0]  col_out_598;
wire  [511:0]  col_out_599;
wire  [511:0]  col_out_600;
wire  [511:0]  col_out_601;
wire  [511:0]  col_out_602;
wire  [511:0]  col_out_603;
wire  [511:0]  col_out_604;
wire  [511:0]  col_out_605;
wire  [511:0]  col_out_606;
wire  [511:0]  col_out_607;
wire  [511:0]  col_out_608;
wire  [511:0]  col_out_609;
wire  [511:0]  col_out_610;
wire  [511:0]  col_out_611;
wire  [511:0]  col_out_612;
wire  [511:0]  col_out_613;
wire  [511:0]  col_out_614;
wire  [511:0]  col_out_615;
wire  [511:0]  col_out_616;
wire  [511:0]  col_out_617;
wire  [511:0]  col_out_618;
wire  [511:0]  col_out_619;
wire  [511:0]  col_out_620;
wire  [511:0]  col_out_621;
wire  [511:0]  col_out_622;
wire  [511:0]  col_out_623;
wire  [511:0]  col_out_624;
wire  [511:0]  col_out_625;
wire  [511:0]  col_out_626;
wire  [511:0]  col_out_627;
wire  [511:0]  col_out_628;
wire  [511:0]  col_out_629;
wire  [511:0]  col_out_630;
wire  [511:0]  col_out_631;
wire  [511:0]  col_out_632;
wire  [511:0]  col_out_633;
wire  [511:0]  col_out_634;
wire  [511:0]  col_out_635;
wire  [511:0]  col_out_636;
wire  [511:0]  col_out_637;
wire  [511:0]  col_out_638;
wire  [511:0]  col_out_639;
wire  [511:0]  col_out_640;
wire  [511:0]  col_out_641;
wire  [511:0]  col_out_642;
wire  [511:0]  col_out_643;
wire  [511:0]  col_out_644;
wire  [511:0]  col_out_645;
wire  [511:0]  col_out_646;
wire  [511:0]  col_out_647;
wire  [511:0]  col_out_648;
wire  [511:0]  col_out_649;
wire  [511:0]  col_out_650;
wire  [511:0]  col_out_651;
wire  [511:0]  col_out_652;
wire  [511:0]  col_out_653;
wire  [511:0]  col_out_654;
wire  [511:0]  col_out_655;
wire  [511:0]  col_out_656;
wire  [511:0]  col_out_657;
wire  [511:0]  col_out_658;
wire  [511:0]  col_out_659;
wire  [511:0]  col_out_660;
wire  [511:0]  col_out_661;
wire  [511:0]  col_out_662;
wire  [511:0]  col_out_663;
wire  [511:0]  col_out_664;
wire  [511:0]  col_out_665;
wire  [511:0]  col_out_666;
wire  [511:0]  col_out_667;
wire  [511:0]  col_out_668;
wire  [511:0]  col_out_669;
wire  [511:0]  col_out_670;
wire  [511:0]  col_out_671;
wire  [511:0]  col_out_672;
wire  [511:0]  col_out_673;
wire  [511:0]  col_out_674;
wire  [511:0]  col_out_675;
wire  [511:0]  col_out_676;
wire  [511:0]  col_out_677;
wire  [511:0]  col_out_678;
wire  [511:0]  col_out_679;
wire  [511:0]  col_out_680;
wire  [511:0]  col_out_681;
wire  [511:0]  col_out_682;
wire  [511:0]  col_out_683;
wire  [511:0]  col_out_684;
wire  [511:0]  col_out_685;
wire  [511:0]  col_out_686;
wire  [511:0]  col_out_687;
wire  [511:0]  col_out_688;
wire  [511:0]  col_out_689;
wire  [511:0]  col_out_690;
wire  [511:0]  col_out_691;
wire  [511:0]  col_out_692;
wire  [511:0]  col_out_693;
wire  [511:0]  col_out_694;
wire  [511:0]  col_out_695;
wire  [511:0]  col_out_696;
wire  [511:0]  col_out_697;
wire  [511:0]  col_out_698;
wire  [511:0]  col_out_699;
wire  [511:0]  col_out_700;
wire  [511:0]  col_out_701;
wire  [511:0]  col_out_702;
wire  [511:0]  col_out_703;
wire  [511:0]  col_out_704;
wire  [511:0]  col_out_705;
wire  [511:0]  col_out_706;
wire  [511:0]  col_out_707;
wire  [511:0]  col_out_708;
wire  [511:0]  col_out_709;
wire  [511:0]  col_out_710;
wire  [511:0]  col_out_711;
wire  [511:0]  col_out_712;
wire  [511:0]  col_out_713;
wire  [511:0]  col_out_714;
wire  [511:0]  col_out_715;
wire  [511:0]  col_out_716;
wire  [511:0]  col_out_717;
wire  [511:0]  col_out_718;
wire  [511:0]  col_out_719;
wire  [511:0]  col_out_720;
wire  [511:0]  col_out_721;
wire  [511:0]  col_out_722;
wire  [511:0]  col_out_723;
wire  [511:0]  col_out_724;
wire  [511:0]  col_out_725;
wire  [511:0]  col_out_726;
wire  [511:0]  col_out_727;
wire  [511:0]  col_out_728;
wire  [511:0]  col_out_729;
wire  [511:0]  col_out_730;
wire  [511:0]  col_out_731;
wire  [511:0]  col_out_732;
wire  [511:0]  col_out_733;
wire  [511:0]  col_out_734;
wire  [511:0]  col_out_735;
wire  [511:0]  col_out_736;
wire  [511:0]  col_out_737;
wire  [511:0]  col_out_738;
wire  [511:0]  col_out_739;
wire  [511:0]  col_out_740;
wire  [511:0]  col_out_741;
wire  [511:0]  col_out_742;
wire  [511:0]  col_out_743;
wire  [511:0]  col_out_744;
wire  [511:0]  col_out_745;
wire  [511:0]  col_out_746;
wire  [511:0]  col_out_747;
wire  [511:0]  col_out_748;
wire  [511:0]  col_out_749;
wire  [511:0]  col_out_750;
wire  [511:0]  col_out_751;
wire  [511:0]  col_out_752;
wire  [511:0]  col_out_753;
wire  [511:0]  col_out_754;
wire  [511:0]  col_out_755;
wire  [511:0]  col_out_756;
wire  [511:0]  col_out_757;
wire  [511:0]  col_out_758;
wire  [511:0]  col_out_759;
wire  [511:0]  col_out_760;
wire  [511:0]  col_out_761;
wire  [511:0]  col_out_762;
wire  [511:0]  col_out_763;
wire  [511:0]  col_out_764;
wire  [511:0]  col_out_765;
wire  [511:0]  col_out_766;
wire  [511:0]  col_out_767;
wire  [511:0]  col_out_768;
wire  [511:0]  col_out_769;
wire  [511:0]  col_out_770;
wire  [511:0]  col_out_771;
wire  [511:0]  col_out_772;
wire  [511:0]  col_out_773;
wire  [511:0]  col_out_774;
wire  [511:0]  col_out_775;
wire  [511:0]  col_out_776;
wire  [511:0]  col_out_777;
wire  [511:0]  col_out_778;
wire  [511:0]  col_out_779;
wire  [511:0]  col_out_780;
wire  [511:0]  col_out_781;
wire  [511:0]  col_out_782;
wire  [511:0]  col_out_783;
wire  [511:0]  col_out_784;
wire  [511:0]  col_out_785;
wire  [511:0]  col_out_786;
wire  [511:0]  col_out_787;
wire  [511:0]  col_out_788;
wire  [511:0]  col_out_789;
wire  [511:0]  col_out_790;
wire  [511:0]  col_out_791;
wire  [511:0]  col_out_792;
wire  [511:0]  col_out_793;
wire  [511:0]  col_out_794;
wire  [511:0]  col_out_795;
wire  [511:0]  col_out_796;
wire  [511:0]  col_out_797;
wire  [511:0]  col_out_798;
wire  [511:0]  col_out_799;
wire  [511:0]  col_out_800;
wire  [511:0]  col_out_801;
wire  [511:0]  col_out_802;
wire  [511:0]  col_out_803;
wire  [511:0]  col_out_804;
wire  [511:0]  col_out_805;
wire  [511:0]  col_out_806;
wire  [511:0]  col_out_807;
wire  [511:0]  col_out_808;
wire  [511:0]  col_out_809;
wire  [511:0]  col_out_810;
wire  [511:0]  col_out_811;
wire  [511:0]  col_out_812;
wire  [511:0]  col_out_813;
wire  [511:0]  col_out_814;
wire  [511:0]  col_out_815;
wire  [511:0]  col_out_816;
wire  [511:0]  col_out_817;
wire  [511:0]  col_out_818;
wire  [511:0]  col_out_819;
wire  [511:0]  col_out_820;
wire  [511:0]  col_out_821;
wire  [511:0]  col_out_822;
wire  [511:0]  col_out_823;
wire  [511:0]  col_out_824;
wire  [511:0]  col_out_825;
wire  [511:0]  col_out_826;
wire  [511:0]  col_out_827;
wire  [511:0]  col_out_828;
wire  [511:0]  col_out_829;
wire  [511:0]  col_out_830;
wire  [511:0]  col_out_831;
wire  [511:0]  col_out_832;
wire  [511:0]  col_out_833;
wire  [511:0]  col_out_834;
wire  [511:0]  col_out_835;
wire  [511:0]  col_out_836;
wire  [511:0]  col_out_837;
wire  [511:0]  col_out_838;
wire  [511:0]  col_out_839;
wire  [511:0]  col_out_840;
wire  [511:0]  col_out_841;
wire  [511:0]  col_out_842;
wire  [511:0]  col_out_843;
wire  [511:0]  col_out_844;
wire  [511:0]  col_out_845;
wire  [511:0]  col_out_846;
wire  [511:0]  col_out_847;
wire  [511:0]  col_out_848;
wire  [511:0]  col_out_849;
wire  [511:0]  col_out_850;
wire  [511:0]  col_out_851;
wire  [511:0]  col_out_852;
wire  [511:0]  col_out_853;
wire  [511:0]  col_out_854;
wire  [511:0]  col_out_855;
wire  [511:0]  col_out_856;
wire  [511:0]  col_out_857;
wire  [511:0]  col_out_858;
wire  [511:0]  col_out_859;
wire  [511:0]  col_out_860;
wire  [511:0]  col_out_861;
wire  [511:0]  col_out_862;
wire  [511:0]  col_out_863;
wire  [511:0]  col_out_864;
wire  [511:0]  col_out_865;
wire  [511:0]  col_out_866;
wire  [511:0]  col_out_867;
wire  [511:0]  col_out_868;
wire  [511:0]  col_out_869;
wire  [511:0]  col_out_870;
wire  [511:0]  col_out_871;
wire  [511:0]  col_out_872;
wire  [511:0]  col_out_873;
wire  [511:0]  col_out_874;
wire  [511:0]  col_out_875;
wire  [511:0]  col_out_876;
wire  [511:0]  col_out_877;
wire  [511:0]  col_out_878;
wire  [511:0]  col_out_879;
wire  [511:0]  col_out_880;
wire  [511:0]  col_out_881;
wire  [511:0]  col_out_882;
wire  [511:0]  col_out_883;
wire  [511:0]  col_out_884;
wire  [511:0]  col_out_885;
wire  [511:0]  col_out_886;
wire  [511:0]  col_out_887;
wire  [511:0]  col_out_888;
wire  [511:0]  col_out_889;
wire  [511:0]  col_out_890;
wire  [511:0]  col_out_891;
wire  [511:0]  col_out_892;
wire  [511:0]  col_out_893;
wire  [511:0]  col_out_894;
wire  [511:0]  col_out_895;
wire  [511:0]  col_out_896;
wire  [511:0]  col_out_897;
wire  [511:0]  col_out_898;
wire  [511:0]  col_out_899;
wire  [511:0]  col_out_900;
wire  [511:0]  col_out_901;
wire  [511:0]  col_out_902;
wire  [511:0]  col_out_903;
wire  [511:0]  col_out_904;
wire  [511:0]  col_out_905;
wire  [511:0]  col_out_906;
wire  [511:0]  col_out_907;
wire  [511:0]  col_out_908;
wire  [511:0]  col_out_909;
wire  [511:0]  col_out_910;
wire  [511:0]  col_out_911;
wire  [511:0]  col_out_912;
wire  [511:0]  col_out_913;
wire  [511:0]  col_out_914;
wire  [511:0]  col_out_915;
wire  [511:0]  col_out_916;
wire  [511:0]  col_out_917;
wire  [511:0]  col_out_918;
wire  [511:0]  col_out_919;
wire  [511:0]  col_out_920;
wire  [511:0]  col_out_921;
wire  [511:0]  col_out_922;
wire  [511:0]  col_out_923;
wire  [511:0]  col_out_924;
wire  [511:0]  col_out_925;
wire  [511:0]  col_out_926;
wire  [511:0]  col_out_927;
wire  [511:0]  col_out_928;
wire  [511:0]  col_out_929;
wire  [511:0]  col_out_930;
wire  [511:0]  col_out_931;
wire  [511:0]  col_out_932;
wire  [511:0]  col_out_933;
wire  [511:0]  col_out_934;
wire  [511:0]  col_out_935;
wire  [511:0]  col_out_936;
wire  [511:0]  col_out_937;
wire  [511:0]  col_out_938;
wire  [511:0]  col_out_939;
wire  [511:0]  col_out_940;
wire  [511:0]  col_out_941;
wire  [511:0]  col_out_942;
wire  [511:0]  col_out_943;
wire  [511:0]  col_out_944;
wire  [511:0]  col_out_945;
wire  [511:0]  col_out_946;
wire  [511:0]  col_out_947;
wire  [511:0]  col_out_948;
wire  [511:0]  col_out_949;
wire  [511:0]  col_out_950;
wire  [511:0]  col_out_951;
wire  [511:0]  col_out_952;
wire  [511:0]  col_out_953;
wire  [511:0]  col_out_954;
wire  [511:0]  col_out_955;
wire  [511:0]  col_out_956;
wire  [511:0]  col_out_957;
wire  [511:0]  col_out_958;
wire  [511:0]  col_out_959;
wire  [511:0]  col_out_960;
wire  [511:0]  col_out_961;
wire  [511:0]  col_out_962;
wire  [511:0]  col_out_963;
wire  [511:0]  col_out_964;
wire  [511:0]  col_out_965;
wire  [511:0]  col_out_966;
wire  [511:0]  col_out_967;
wire  [511:0]  col_out_968;
wire  [511:0]  col_out_969;
wire  [511:0]  col_out_970;
wire  [511:0]  col_out_971;
wire  [511:0]  col_out_972;
wire  [511:0]  col_out_973;
wire  [511:0]  col_out_974;
wire  [511:0]  col_out_975;
wire  [511:0]  col_out_976;
wire  [511:0]  col_out_977;
wire  [511:0]  col_out_978;
wire  [511:0]  col_out_979;
wire  [511:0]  col_out_980;
wire  [511:0]  col_out_981;
wire  [511:0]  col_out_982;
wire  [511:0]  col_out_983;
wire  [511:0]  col_out_984;
wire  [511:0]  col_out_985;
wire  [511:0]  col_out_986;
wire  [511:0]  col_out_987;
wire  [511:0]  col_out_988;
wire  [511:0]  col_out_989;
wire  [511:0]  col_out_990;
wire  [511:0]  col_out_991;
wire  [511:0]  col_out_992;
wire  [511:0]  col_out_993;
wire  [511:0]  col_out_994;
wire  [511:0]  col_out_995;
wire  [511:0]  col_out_996;
wire  [511:0]  col_out_997;
wire  [511:0]  col_out_998;
wire  [511:0]  col_out_999;
wire  [511:0]  col_out_1000;
wire  [511:0]  col_out_1001;
wire  [511:0]  col_out_1002;
wire  [511:0]  col_out_1003;
wire  [511:0]  col_out_1004;
wire  [511:0]  col_out_1005;
wire  [511:0]  col_out_1006;
wire  [511:0]  col_out_1007;
wire  [511:0]  col_out_1008;
wire  [511:0]  col_out_1009;
wire  [511:0]  col_out_1010;
wire  [511:0]  col_out_1011;
wire  [511:0]  col_out_1012;
wire  [511:0]  col_out_1013;
wire  [511:0]  col_out_1014;
wire  [511:0]  col_out_1015;
wire  [511:0]  col_out_1016;
wire  [511:0]  col_out_1017;
wire  [511:0]  col_out_1018;
wire  [511:0]  col_out_1019;
wire  [511:0]  col_out_1020;
wire  [511:0]  col_out_1021;
wire  [511:0]  col_out_1022;
wire  [511:0]  col_out_1023;

data_in_mux  u_data_in_mux (
    .a                       ( reg_a                       ),
    .sel_hp                  ( sel_hp                  ),
    .partial_product_high0   ( partial_product_high0   ),
    .partial_product_high1   ( partial_product_high1   ),
    .partial_product_low0    ( partial_product_low0    ),
    .partial_product_low1    ( partial_product_low1    ),
    .sel_data_in             ( sel_data_in             ),

    .col_out_0               ( col_out_0               ),
    .col_out_1               ( col_out_1               ),
    .col_out_2               ( col_out_2               ),
    .col_out_3               ( col_out_3               ),
    .col_out_4               ( col_out_4               ),
    .col_out_5               ( col_out_5               ),
    .col_out_6               ( col_out_6               ),
    .col_out_7               ( col_out_7               ),
    .col_out_8               ( col_out_8               ),
    .col_out_9               ( col_out_9               ),
    .col_out_10              ( col_out_10              ),
    .col_out_11              ( col_out_11              ),
    .col_out_12              ( col_out_12              ),
    .col_out_13              ( col_out_13              ),
    .col_out_14              ( col_out_14              ),
    .col_out_15              ( col_out_15              ),
    .col_out_16              ( col_out_16              ),
    .col_out_17              ( col_out_17              ),
    .col_out_18              ( col_out_18              ),
    .col_out_19              ( col_out_19              ),
    .col_out_20              ( col_out_20              ),
    .col_out_21              ( col_out_21              ),
    .col_out_22              ( col_out_22              ),
    .col_out_23              ( col_out_23              ),
    .col_out_24              ( col_out_24              ),
    .col_out_25              ( col_out_25              ),
    .col_out_26              ( col_out_26              ),
    .col_out_27              ( col_out_27              ),
    .col_out_28              ( col_out_28              ),
    .col_out_29              ( col_out_29              ),
    .col_out_30              ( col_out_30              ),
    .col_out_31              ( col_out_31              ),
    .col_out_32              ( col_out_32              ),
    .col_out_33              ( col_out_33              ),
    .col_out_34              ( col_out_34              ),
    .col_out_35              ( col_out_35              ),
    .col_out_36              ( col_out_36              ),
    .col_out_37              ( col_out_37              ),
    .col_out_38              ( col_out_38              ),
    .col_out_39              ( col_out_39              ),
    .col_out_40              ( col_out_40              ),
    .col_out_41              ( col_out_41              ),
    .col_out_42              ( col_out_42              ),
    .col_out_43              ( col_out_43              ),
    .col_out_44              ( col_out_44              ),
    .col_out_45              ( col_out_45              ),
    .col_out_46              ( col_out_46              ),
    .col_out_47              ( col_out_47              ),
    .col_out_48              ( col_out_48              ),
    .col_out_49              ( col_out_49              ),
    .col_out_50              ( col_out_50              ),
    .col_out_51              ( col_out_51              ),
    .col_out_52              ( col_out_52              ),
    .col_out_53              ( col_out_53              ),
    .col_out_54              ( col_out_54              ),
    .col_out_55              ( col_out_55              ),
    .col_out_56              ( col_out_56              ),
    .col_out_57              ( col_out_57              ),
    .col_out_58              ( col_out_58              ),
    .col_out_59              ( col_out_59              ),
    .col_out_60              ( col_out_60              ),
    .col_out_61              ( col_out_61              ),
    .col_out_62              ( col_out_62              ),
    .col_out_63              ( col_out_63              ),
    .col_out_64              ( col_out_64              ),
    .col_out_65              ( col_out_65              ),
    .col_out_66              ( col_out_66              ),
    .col_out_67              ( col_out_67              ),
    .col_out_68              ( col_out_68              ),
    .col_out_69              ( col_out_69              ),
    .col_out_70              ( col_out_70              ),
    .col_out_71              ( col_out_71              ),
    .col_out_72              ( col_out_72              ),
    .col_out_73              ( col_out_73              ),
    .col_out_74              ( col_out_74              ),
    .col_out_75              ( col_out_75              ),
    .col_out_76              ( col_out_76              ),
    .col_out_77              ( col_out_77              ),
    .col_out_78              ( col_out_78              ),
    .col_out_79              ( col_out_79              ),
    .col_out_80              ( col_out_80              ),
    .col_out_81              ( col_out_81              ),
    .col_out_82              ( col_out_82              ),
    .col_out_83              ( col_out_83              ),
    .col_out_84              ( col_out_84              ),
    .col_out_85              ( col_out_85              ),
    .col_out_86              ( col_out_86              ),
    .col_out_87              ( col_out_87              ),
    .col_out_88              ( col_out_88              ),
    .col_out_89              ( col_out_89              ),
    .col_out_90              ( col_out_90              ),
    .col_out_91              ( col_out_91              ),
    .col_out_92              ( col_out_92              ),
    .col_out_93              ( col_out_93              ),
    .col_out_94              ( col_out_94              ),
    .col_out_95              ( col_out_95              ),
    .col_out_96              ( col_out_96              ),
    .col_out_97              ( col_out_97              ),
    .col_out_98              ( col_out_98              ),
    .col_out_99              ( col_out_99              ),
    .col_out_100             ( col_out_100             ),
    .col_out_101             ( col_out_101             ),
    .col_out_102             ( col_out_102             ),
    .col_out_103             ( col_out_103             ),
    .col_out_104             ( col_out_104             ),
    .col_out_105             ( col_out_105             ),
    .col_out_106             ( col_out_106             ),
    .col_out_107             ( col_out_107             ),
    .col_out_108             ( col_out_108             ),
    .col_out_109             ( col_out_109             ),
    .col_out_110             ( col_out_110             ),
    .col_out_111             ( col_out_111             ),
    .col_out_112             ( col_out_112             ),
    .col_out_113             ( col_out_113             ),
    .col_out_114             ( col_out_114             ),
    .col_out_115             ( col_out_115             ),
    .col_out_116             ( col_out_116             ),
    .col_out_117             ( col_out_117             ),
    .col_out_118             ( col_out_118             ),
    .col_out_119             ( col_out_119             ),
    .col_out_120             ( col_out_120             ),
    .col_out_121             ( col_out_121             ),
    .col_out_122             ( col_out_122             ),
    .col_out_123             ( col_out_123             ),
    .col_out_124             ( col_out_124             ),
    .col_out_125             ( col_out_125             ),
    .col_out_126             ( col_out_126             ),
    .col_out_127             ( col_out_127             ),
    .col_out_128             ( col_out_128             ),
    .col_out_129             ( col_out_129             ),
    .col_out_130             ( col_out_130             ),
    .col_out_131             ( col_out_131             ),
    .col_out_132             ( col_out_132             ),
    .col_out_133             ( col_out_133             ),
    .col_out_134             ( col_out_134             ),
    .col_out_135             ( col_out_135             ),
    .col_out_136             ( col_out_136             ),
    .col_out_137             ( col_out_137             ),
    .col_out_138             ( col_out_138             ),
    .col_out_139             ( col_out_139             ),
    .col_out_140             ( col_out_140             ),
    .col_out_141             ( col_out_141             ),
    .col_out_142             ( col_out_142             ),
    .col_out_143             ( col_out_143             ),
    .col_out_144             ( col_out_144             ),
    .col_out_145             ( col_out_145             ),
    .col_out_146             ( col_out_146             ),
    .col_out_147             ( col_out_147             ),
    .col_out_148             ( col_out_148             ),
    .col_out_149             ( col_out_149             ),
    .col_out_150             ( col_out_150             ),
    .col_out_151             ( col_out_151             ),
    .col_out_152             ( col_out_152             ),
    .col_out_153             ( col_out_153             ),
    .col_out_154             ( col_out_154             ),
    .col_out_155             ( col_out_155             ),
    .col_out_156             ( col_out_156             ),
    .col_out_157             ( col_out_157             ),
    .col_out_158             ( col_out_158             ),
    .col_out_159             ( col_out_159             ),
    .col_out_160             ( col_out_160             ),
    .col_out_161             ( col_out_161             ),
    .col_out_162             ( col_out_162             ),
    .col_out_163             ( col_out_163             ),
    .col_out_164             ( col_out_164             ),
    .col_out_165             ( col_out_165             ),
    .col_out_166             ( col_out_166             ),
    .col_out_167             ( col_out_167             ),
    .col_out_168             ( col_out_168             ),
    .col_out_169             ( col_out_169             ),
    .col_out_170             ( col_out_170             ),
    .col_out_171             ( col_out_171             ),
    .col_out_172             ( col_out_172             ),
    .col_out_173             ( col_out_173             ),
    .col_out_174             ( col_out_174             ),
    .col_out_175             ( col_out_175             ),
    .col_out_176             ( col_out_176             ),
    .col_out_177             ( col_out_177             ),
    .col_out_178             ( col_out_178             ),
    .col_out_179             ( col_out_179             ),
    .col_out_180             ( col_out_180             ),
    .col_out_181             ( col_out_181             ),
    .col_out_182             ( col_out_182             ),
    .col_out_183             ( col_out_183             ),
    .col_out_184             ( col_out_184             ),
    .col_out_185             ( col_out_185             ),
    .col_out_186             ( col_out_186             ),
    .col_out_187             ( col_out_187             ),
    .col_out_188             ( col_out_188             ),
    .col_out_189             ( col_out_189             ),
    .col_out_190             ( col_out_190             ),
    .col_out_191             ( col_out_191             ),
    .col_out_192             ( col_out_192             ),
    .col_out_193             ( col_out_193             ),
    .col_out_194             ( col_out_194             ),
    .col_out_195             ( col_out_195             ),
    .col_out_196             ( col_out_196             ),
    .col_out_197             ( col_out_197             ),
    .col_out_198             ( col_out_198             ),
    .col_out_199             ( col_out_199             ),
    .col_out_200             ( col_out_200             ),
    .col_out_201             ( col_out_201             ),
    .col_out_202             ( col_out_202             ),
    .col_out_203             ( col_out_203             ),
    .col_out_204             ( col_out_204             ),
    .col_out_205             ( col_out_205             ),
    .col_out_206             ( col_out_206             ),
    .col_out_207             ( col_out_207             ),
    .col_out_208             ( col_out_208             ),
    .col_out_209             ( col_out_209             ),
    .col_out_210             ( col_out_210             ),
    .col_out_211             ( col_out_211             ),
    .col_out_212             ( col_out_212             ),
    .col_out_213             ( col_out_213             ),
    .col_out_214             ( col_out_214             ),
    .col_out_215             ( col_out_215             ),
    .col_out_216             ( col_out_216             ),
    .col_out_217             ( col_out_217             ),
    .col_out_218             ( col_out_218             ),
    .col_out_219             ( col_out_219             ),
    .col_out_220             ( col_out_220             ),
    .col_out_221             ( col_out_221             ),
    .col_out_222             ( col_out_222             ),
    .col_out_223             ( col_out_223             ),
    .col_out_224             ( col_out_224             ),
    .col_out_225             ( col_out_225             ),
    .col_out_226             ( col_out_226             ),
    .col_out_227             ( col_out_227             ),
    .col_out_228             ( col_out_228             ),
    .col_out_229             ( col_out_229             ),
    .col_out_230             ( col_out_230             ),
    .col_out_231             ( col_out_231             ),
    .col_out_232             ( col_out_232             ),
    .col_out_233             ( col_out_233             ),
    .col_out_234             ( col_out_234             ),
    .col_out_235             ( col_out_235             ),
    .col_out_236             ( col_out_236             ),
    .col_out_237             ( col_out_237             ),
    .col_out_238             ( col_out_238             ),
    .col_out_239             ( col_out_239             ),
    .col_out_240             ( col_out_240             ),
    .col_out_241             ( col_out_241             ),
    .col_out_242             ( col_out_242             ),
    .col_out_243             ( col_out_243             ),
    .col_out_244             ( col_out_244             ),
    .col_out_245             ( col_out_245             ),
    .col_out_246             ( col_out_246             ),
    .col_out_247             ( col_out_247             ),
    .col_out_248             ( col_out_248             ),
    .col_out_249             ( col_out_249             ),
    .col_out_250             ( col_out_250             ),
    .col_out_251             ( col_out_251             ),
    .col_out_252             ( col_out_252             ),
    .col_out_253             ( col_out_253             ),
    .col_out_254             ( col_out_254             ),
    .col_out_255             ( col_out_255             ),
    .col_out_256             ( col_out_256             ),
    .col_out_257             ( col_out_257             ),
    .col_out_258             ( col_out_258             ),
    .col_out_259             ( col_out_259             ),
    .col_out_260             ( col_out_260             ),
    .col_out_261             ( col_out_261             ),
    .col_out_262             ( col_out_262             ),
    .col_out_263             ( col_out_263             ),
    .col_out_264             ( col_out_264             ),
    .col_out_265             ( col_out_265             ),
    .col_out_266             ( col_out_266             ),
    .col_out_267             ( col_out_267             ),
    .col_out_268             ( col_out_268             ),
    .col_out_269             ( col_out_269             ),
    .col_out_270             ( col_out_270             ),
    .col_out_271             ( col_out_271             ),
    .col_out_272             ( col_out_272             ),
    .col_out_273             ( col_out_273             ),
    .col_out_274             ( col_out_274             ),
    .col_out_275             ( col_out_275             ),
    .col_out_276             ( col_out_276             ),
    .col_out_277             ( col_out_277             ),
    .col_out_278             ( col_out_278             ),
    .col_out_279             ( col_out_279             ),
    .col_out_280             ( col_out_280             ),
    .col_out_281             ( col_out_281             ),
    .col_out_282             ( col_out_282             ),
    .col_out_283             ( col_out_283             ),
    .col_out_284             ( col_out_284             ),
    .col_out_285             ( col_out_285             ),
    .col_out_286             ( col_out_286             ),
    .col_out_287             ( col_out_287             ),
    .col_out_288             ( col_out_288             ),
    .col_out_289             ( col_out_289             ),
    .col_out_290             ( col_out_290             ),
    .col_out_291             ( col_out_291             ),
    .col_out_292             ( col_out_292             ),
    .col_out_293             ( col_out_293             ),
    .col_out_294             ( col_out_294             ),
    .col_out_295             ( col_out_295             ),
    .col_out_296             ( col_out_296             ),
    .col_out_297             ( col_out_297             ),
    .col_out_298             ( col_out_298             ),
    .col_out_299             ( col_out_299             ),
    .col_out_300             ( col_out_300             ),
    .col_out_301             ( col_out_301             ),
    .col_out_302             ( col_out_302             ),
    .col_out_303             ( col_out_303             ),
    .col_out_304             ( col_out_304             ),
    .col_out_305             ( col_out_305             ),
    .col_out_306             ( col_out_306             ),
    .col_out_307             ( col_out_307             ),
    .col_out_308             ( col_out_308             ),
    .col_out_309             ( col_out_309             ),
    .col_out_310             ( col_out_310             ),
    .col_out_311             ( col_out_311             ),
    .col_out_312             ( col_out_312             ),
    .col_out_313             ( col_out_313             ),
    .col_out_314             ( col_out_314             ),
    .col_out_315             ( col_out_315             ),
    .col_out_316             ( col_out_316             ),
    .col_out_317             ( col_out_317             ),
    .col_out_318             ( col_out_318             ),
    .col_out_319             ( col_out_319             ),
    .col_out_320             ( col_out_320             ),
    .col_out_321             ( col_out_321             ),
    .col_out_322             ( col_out_322             ),
    .col_out_323             ( col_out_323             ),
    .col_out_324             ( col_out_324             ),
    .col_out_325             ( col_out_325             ),
    .col_out_326             ( col_out_326             ),
    .col_out_327             ( col_out_327             ),
    .col_out_328             ( col_out_328             ),
    .col_out_329             ( col_out_329             ),
    .col_out_330             ( col_out_330             ),
    .col_out_331             ( col_out_331             ),
    .col_out_332             ( col_out_332             ),
    .col_out_333             ( col_out_333             ),
    .col_out_334             ( col_out_334             ),
    .col_out_335             ( col_out_335             ),
    .col_out_336             ( col_out_336             ),
    .col_out_337             ( col_out_337             ),
    .col_out_338             ( col_out_338             ),
    .col_out_339             ( col_out_339             ),
    .col_out_340             ( col_out_340             ),
    .col_out_341             ( col_out_341             ),
    .col_out_342             ( col_out_342             ),
    .col_out_343             ( col_out_343             ),
    .col_out_344             ( col_out_344             ),
    .col_out_345             ( col_out_345             ),
    .col_out_346             ( col_out_346             ),
    .col_out_347             ( col_out_347             ),
    .col_out_348             ( col_out_348             ),
    .col_out_349             ( col_out_349             ),
    .col_out_350             ( col_out_350             ),
    .col_out_351             ( col_out_351             ),
    .col_out_352             ( col_out_352             ),
    .col_out_353             ( col_out_353             ),
    .col_out_354             ( col_out_354             ),
    .col_out_355             ( col_out_355             ),
    .col_out_356             ( col_out_356             ),
    .col_out_357             ( col_out_357             ),
    .col_out_358             ( col_out_358             ),
    .col_out_359             ( col_out_359             ),
    .col_out_360             ( col_out_360             ),
    .col_out_361             ( col_out_361             ),
    .col_out_362             ( col_out_362             ),
    .col_out_363             ( col_out_363             ),
    .col_out_364             ( col_out_364             ),
    .col_out_365             ( col_out_365             ),
    .col_out_366             ( col_out_366             ),
    .col_out_367             ( col_out_367             ),
    .col_out_368             ( col_out_368             ),
    .col_out_369             ( col_out_369             ),
    .col_out_370             ( col_out_370             ),
    .col_out_371             ( col_out_371             ),
    .col_out_372             ( col_out_372             ),
    .col_out_373             ( col_out_373             ),
    .col_out_374             ( col_out_374             ),
    .col_out_375             ( col_out_375             ),
    .col_out_376             ( col_out_376             ),
    .col_out_377             ( col_out_377             ),
    .col_out_378             ( col_out_378             ),
    .col_out_379             ( col_out_379             ),
    .col_out_380             ( col_out_380             ),
    .col_out_381             ( col_out_381             ),
    .col_out_382             ( col_out_382             ),
    .col_out_383             ( col_out_383             ),
    .col_out_384             ( col_out_384             ),
    .col_out_385             ( col_out_385             ),
    .col_out_386             ( col_out_386             ),
    .col_out_387             ( col_out_387             ),
    .col_out_388             ( col_out_388             ),
    .col_out_389             ( col_out_389             ),
    .col_out_390             ( col_out_390             ),
    .col_out_391             ( col_out_391             ),
    .col_out_392             ( col_out_392             ),
    .col_out_393             ( col_out_393             ),
    .col_out_394             ( col_out_394             ),
    .col_out_395             ( col_out_395             ),
    .col_out_396             ( col_out_396             ),
    .col_out_397             ( col_out_397             ),
    .col_out_398             ( col_out_398             ),
    .col_out_399             ( col_out_399             ),
    .col_out_400             ( col_out_400             ),
    .col_out_401             ( col_out_401             ),
    .col_out_402             ( col_out_402             ),
    .col_out_403             ( col_out_403             ),
    .col_out_404             ( col_out_404             ),
    .col_out_405             ( col_out_405             ),
    .col_out_406             ( col_out_406             ),
    .col_out_407             ( col_out_407             ),
    .col_out_408             ( col_out_408             ),
    .col_out_409             ( col_out_409             ),
    .col_out_410             ( col_out_410             ),
    .col_out_411             ( col_out_411             ),
    .col_out_412             ( col_out_412             ),
    .col_out_413             ( col_out_413             ),
    .col_out_414             ( col_out_414             ),
    .col_out_415             ( col_out_415             ),
    .col_out_416             ( col_out_416             ),
    .col_out_417             ( col_out_417             ),
    .col_out_418             ( col_out_418             ),
    .col_out_419             ( col_out_419             ),
    .col_out_420             ( col_out_420             ),
    .col_out_421             ( col_out_421             ),
    .col_out_422             ( col_out_422             ),
    .col_out_423             ( col_out_423             ),
    .col_out_424             ( col_out_424             ),
    .col_out_425             ( col_out_425             ),
    .col_out_426             ( col_out_426             ),
    .col_out_427             ( col_out_427             ),
    .col_out_428             ( col_out_428             ),
    .col_out_429             ( col_out_429             ),
    .col_out_430             ( col_out_430             ),
    .col_out_431             ( col_out_431             ),
    .col_out_432             ( col_out_432             ),
    .col_out_433             ( col_out_433             ),
    .col_out_434             ( col_out_434             ),
    .col_out_435             ( col_out_435             ),
    .col_out_436             ( col_out_436             ),
    .col_out_437             ( col_out_437             ),
    .col_out_438             ( col_out_438             ),
    .col_out_439             ( col_out_439             ),
    .col_out_440             ( col_out_440             ),
    .col_out_441             ( col_out_441             ),
    .col_out_442             ( col_out_442             ),
    .col_out_443             ( col_out_443             ),
    .col_out_444             ( col_out_444             ),
    .col_out_445             ( col_out_445             ),
    .col_out_446             ( col_out_446             ),
    .col_out_447             ( col_out_447             ),
    .col_out_448             ( col_out_448             ),
    .col_out_449             ( col_out_449             ),
    .col_out_450             ( col_out_450             ),
    .col_out_451             ( col_out_451             ),
    .col_out_452             ( col_out_452             ),
    .col_out_453             ( col_out_453             ),
    .col_out_454             ( col_out_454             ),
    .col_out_455             ( col_out_455             ),
    .col_out_456             ( col_out_456             ),
    .col_out_457             ( col_out_457             ),
    .col_out_458             ( col_out_458             ),
    .col_out_459             ( col_out_459             ),
    .col_out_460             ( col_out_460             ),
    .col_out_461             ( col_out_461             ),
    .col_out_462             ( col_out_462             ),
    .col_out_463             ( col_out_463             ),
    .col_out_464             ( col_out_464             ),
    .col_out_465             ( col_out_465             ),
    .col_out_466             ( col_out_466             ),
    .col_out_467             ( col_out_467             ),
    .col_out_468             ( col_out_468             ),
    .col_out_469             ( col_out_469             ),
    .col_out_470             ( col_out_470             ),
    .col_out_471             ( col_out_471             ),
    .col_out_472             ( col_out_472             ),
    .col_out_473             ( col_out_473             ),
    .col_out_474             ( col_out_474             ),
    .col_out_475             ( col_out_475             ),
    .col_out_476             ( col_out_476             ),
    .col_out_477             ( col_out_477             ),
    .col_out_478             ( col_out_478             ),
    .col_out_479             ( col_out_479             ),
    .col_out_480             ( col_out_480             ),
    .col_out_481             ( col_out_481             ),
    .col_out_482             ( col_out_482             ),
    .col_out_483             ( col_out_483             ),
    .col_out_484             ( col_out_484             ),
    .col_out_485             ( col_out_485             ),
    .col_out_486             ( col_out_486             ),
    .col_out_487             ( col_out_487             ),
    .col_out_488             ( col_out_488             ),
    .col_out_489             ( col_out_489             ),
    .col_out_490             ( col_out_490             ),
    .col_out_491             ( col_out_491             ),
    .col_out_492             ( col_out_492             ),
    .col_out_493             ( col_out_493             ),
    .col_out_494             ( col_out_494             ),
    .col_out_495             ( col_out_495             ),
    .col_out_496             ( col_out_496             ),
    .col_out_497             ( col_out_497             ),
    .col_out_498             ( col_out_498             ),
    .col_out_499             ( col_out_499             ),
    .col_out_500             ( col_out_500             ),
    .col_out_501             ( col_out_501             ),
    .col_out_502             ( col_out_502             ),
    .col_out_503             ( col_out_503             ),
    .col_out_504             ( col_out_504             ),
    .col_out_505             ( col_out_505             ),
    .col_out_506             ( col_out_506             ),
    .col_out_507             ( col_out_507             ),
    .col_out_508             ( col_out_508             ),
    .col_out_509             ( col_out_509             ),
    .col_out_510             ( col_out_510             ),
    .col_out_511             ( col_out_511             ),
    .col_out_512             ( col_out_512             ),
    .col_out_513             ( col_out_513             ),
    .col_out_514             ( col_out_514             ),
    .col_out_515             ( col_out_515             ),
    .col_out_516             ( col_out_516             ),
    .col_out_517             ( col_out_517             ),
    .col_out_518             ( col_out_518             ),
    .col_out_519             ( col_out_519             ),
    .col_out_520             ( col_out_520             ),
    .col_out_521             ( col_out_521             ),
    .col_out_522             ( col_out_522             ),
    .col_out_523             ( col_out_523             ),
    .col_out_524             ( col_out_524             ),
    .col_out_525             ( col_out_525             ),
    .col_out_526             ( col_out_526             ),
    .col_out_527             ( col_out_527             ),
    .col_out_528             ( col_out_528             ),
    .col_out_529             ( col_out_529             ),
    .col_out_530             ( col_out_530             ),
    .col_out_531             ( col_out_531             ),
    .col_out_532             ( col_out_532             ),
    .col_out_533             ( col_out_533             ),
    .col_out_534             ( col_out_534             ),
    .col_out_535             ( col_out_535             ),
    .col_out_536             ( col_out_536             ),
    .col_out_537             ( col_out_537             ),
    .col_out_538             ( col_out_538             ),
    .col_out_539             ( col_out_539             ),
    .col_out_540             ( col_out_540             ),
    .col_out_541             ( col_out_541             ),
    .col_out_542             ( col_out_542             ),
    .col_out_543             ( col_out_543             ),
    .col_out_544             ( col_out_544             ),
    .col_out_545             ( col_out_545             ),
    .col_out_546             ( col_out_546             ),
    .col_out_547             ( col_out_547             ),
    .col_out_548             ( col_out_548             ),
    .col_out_549             ( col_out_549             ),
    .col_out_550             ( col_out_550             ),
    .col_out_551             ( col_out_551             ),
    .col_out_552             ( col_out_552             ),
    .col_out_553             ( col_out_553             ),
    .col_out_554             ( col_out_554             ),
    .col_out_555             ( col_out_555             ),
    .col_out_556             ( col_out_556             ),
    .col_out_557             ( col_out_557             ),
    .col_out_558             ( col_out_558             ),
    .col_out_559             ( col_out_559             ),
    .col_out_560             ( col_out_560             ),
    .col_out_561             ( col_out_561             ),
    .col_out_562             ( col_out_562             ),
    .col_out_563             ( col_out_563             ),
    .col_out_564             ( col_out_564             ),
    .col_out_565             ( col_out_565             ),
    .col_out_566             ( col_out_566             ),
    .col_out_567             ( col_out_567             ),
    .col_out_568             ( col_out_568             ),
    .col_out_569             ( col_out_569             ),
    .col_out_570             ( col_out_570             ),
    .col_out_571             ( col_out_571             ),
    .col_out_572             ( col_out_572             ),
    .col_out_573             ( col_out_573             ),
    .col_out_574             ( col_out_574             ),
    .col_out_575             ( col_out_575             ),
    .col_out_576             ( col_out_576             ),
    .col_out_577             ( col_out_577             ),
    .col_out_578             ( col_out_578             ),
    .col_out_579             ( col_out_579             ),
    .col_out_580             ( col_out_580             ),
    .col_out_581             ( col_out_581             ),
    .col_out_582             ( col_out_582             ),
    .col_out_583             ( col_out_583             ),
    .col_out_584             ( col_out_584             ),
    .col_out_585             ( col_out_585             ),
    .col_out_586             ( col_out_586             ),
    .col_out_587             ( col_out_587             ),
    .col_out_588             ( col_out_588             ),
    .col_out_589             ( col_out_589             ),
    .col_out_590             ( col_out_590             ),
    .col_out_591             ( col_out_591             ),
    .col_out_592             ( col_out_592             ),
    .col_out_593             ( col_out_593             ),
    .col_out_594             ( col_out_594             ),
    .col_out_595             ( col_out_595             ),
    .col_out_596             ( col_out_596             ),
    .col_out_597             ( col_out_597             ),
    .col_out_598             ( col_out_598             ),
    .col_out_599             ( col_out_599             ),
    .col_out_600             ( col_out_600             ),
    .col_out_601             ( col_out_601             ),
    .col_out_602             ( col_out_602             ),
    .col_out_603             ( col_out_603             ),
    .col_out_604             ( col_out_604             ),
    .col_out_605             ( col_out_605             ),
    .col_out_606             ( col_out_606             ),
    .col_out_607             ( col_out_607             ),
    .col_out_608             ( col_out_608             ),
    .col_out_609             ( col_out_609             ),
    .col_out_610             ( col_out_610             ),
    .col_out_611             ( col_out_611             ),
    .col_out_612             ( col_out_612             ),
    .col_out_613             ( col_out_613             ),
    .col_out_614             ( col_out_614             ),
    .col_out_615             ( col_out_615             ),
    .col_out_616             ( col_out_616             ),
    .col_out_617             ( col_out_617             ),
    .col_out_618             ( col_out_618             ),
    .col_out_619             ( col_out_619             ),
    .col_out_620             ( col_out_620             ),
    .col_out_621             ( col_out_621             ),
    .col_out_622             ( col_out_622             ),
    .col_out_623             ( col_out_623             ),
    .col_out_624             ( col_out_624             ),
    .col_out_625             ( col_out_625             ),
    .col_out_626             ( col_out_626             ),
    .col_out_627             ( col_out_627             ),
    .col_out_628             ( col_out_628             ),
    .col_out_629             ( col_out_629             ),
    .col_out_630             ( col_out_630             ),
    .col_out_631             ( col_out_631             ),
    .col_out_632             ( col_out_632             ),
    .col_out_633             ( col_out_633             ),
    .col_out_634             ( col_out_634             ),
    .col_out_635             ( col_out_635             ),
    .col_out_636             ( col_out_636             ),
    .col_out_637             ( col_out_637             ),
    .col_out_638             ( col_out_638             ),
    .col_out_639             ( col_out_639             ),
    .col_out_640             ( col_out_640             ),
    .col_out_641             ( col_out_641             ),
    .col_out_642             ( col_out_642             ),
    .col_out_643             ( col_out_643             ),
    .col_out_644             ( col_out_644             ),
    .col_out_645             ( col_out_645             ),
    .col_out_646             ( col_out_646             ),
    .col_out_647             ( col_out_647             ),
    .col_out_648             ( col_out_648             ),
    .col_out_649             ( col_out_649             ),
    .col_out_650             ( col_out_650             ),
    .col_out_651             ( col_out_651             ),
    .col_out_652             ( col_out_652             ),
    .col_out_653             ( col_out_653             ),
    .col_out_654             ( col_out_654             ),
    .col_out_655             ( col_out_655             ),
    .col_out_656             ( col_out_656             ),
    .col_out_657             ( col_out_657             ),
    .col_out_658             ( col_out_658             ),
    .col_out_659             ( col_out_659             ),
    .col_out_660             ( col_out_660             ),
    .col_out_661             ( col_out_661             ),
    .col_out_662             ( col_out_662             ),
    .col_out_663             ( col_out_663             ),
    .col_out_664             ( col_out_664             ),
    .col_out_665             ( col_out_665             ),
    .col_out_666             ( col_out_666             ),
    .col_out_667             ( col_out_667             ),
    .col_out_668             ( col_out_668             ),
    .col_out_669             ( col_out_669             ),
    .col_out_670             ( col_out_670             ),
    .col_out_671             ( col_out_671             ),
    .col_out_672             ( col_out_672             ),
    .col_out_673             ( col_out_673             ),
    .col_out_674             ( col_out_674             ),
    .col_out_675             ( col_out_675             ),
    .col_out_676             ( col_out_676             ),
    .col_out_677             ( col_out_677             ),
    .col_out_678             ( col_out_678             ),
    .col_out_679             ( col_out_679             ),
    .col_out_680             ( col_out_680             ),
    .col_out_681             ( col_out_681             ),
    .col_out_682             ( col_out_682             ),
    .col_out_683             ( col_out_683             ),
    .col_out_684             ( col_out_684             ),
    .col_out_685             ( col_out_685             ),
    .col_out_686             ( col_out_686             ),
    .col_out_687             ( col_out_687             ),
    .col_out_688             ( col_out_688             ),
    .col_out_689             ( col_out_689             ),
    .col_out_690             ( col_out_690             ),
    .col_out_691             ( col_out_691             ),
    .col_out_692             ( col_out_692             ),
    .col_out_693             ( col_out_693             ),
    .col_out_694             ( col_out_694             ),
    .col_out_695             ( col_out_695             ),
    .col_out_696             ( col_out_696             ),
    .col_out_697             ( col_out_697             ),
    .col_out_698             ( col_out_698             ),
    .col_out_699             ( col_out_699             ),
    .col_out_700             ( col_out_700             ),
    .col_out_701             ( col_out_701             ),
    .col_out_702             ( col_out_702             ),
    .col_out_703             ( col_out_703             ),
    .col_out_704             ( col_out_704             ),
    .col_out_705             ( col_out_705             ),
    .col_out_706             ( col_out_706             ),
    .col_out_707             ( col_out_707             ),
    .col_out_708             ( col_out_708             ),
    .col_out_709             ( col_out_709             ),
    .col_out_710             ( col_out_710             ),
    .col_out_711             ( col_out_711             ),
    .col_out_712             ( col_out_712             ),
    .col_out_713             ( col_out_713             ),
    .col_out_714             ( col_out_714             ),
    .col_out_715             ( col_out_715             ),
    .col_out_716             ( col_out_716             ),
    .col_out_717             ( col_out_717             ),
    .col_out_718             ( col_out_718             ),
    .col_out_719             ( col_out_719             ),
    .col_out_720             ( col_out_720             ),
    .col_out_721             ( col_out_721             ),
    .col_out_722             ( col_out_722             ),
    .col_out_723             ( col_out_723             ),
    .col_out_724             ( col_out_724             ),
    .col_out_725             ( col_out_725             ),
    .col_out_726             ( col_out_726             ),
    .col_out_727             ( col_out_727             ),
    .col_out_728             ( col_out_728             ),
    .col_out_729             ( col_out_729             ),
    .col_out_730             ( col_out_730             ),
    .col_out_731             ( col_out_731             ),
    .col_out_732             ( col_out_732             ),
    .col_out_733             ( col_out_733             ),
    .col_out_734             ( col_out_734             ),
    .col_out_735             ( col_out_735             ),
    .col_out_736             ( col_out_736             ),
    .col_out_737             ( col_out_737             ),
    .col_out_738             ( col_out_738             ),
    .col_out_739             ( col_out_739             ),
    .col_out_740             ( col_out_740             ),
    .col_out_741             ( col_out_741             ),
    .col_out_742             ( col_out_742             ),
    .col_out_743             ( col_out_743             ),
    .col_out_744             ( col_out_744             ),
    .col_out_745             ( col_out_745             ),
    .col_out_746             ( col_out_746             ),
    .col_out_747             ( col_out_747             ),
    .col_out_748             ( col_out_748             ),
    .col_out_749             ( col_out_749             ),
    .col_out_750             ( col_out_750             ),
    .col_out_751             ( col_out_751             ),
    .col_out_752             ( col_out_752             ),
    .col_out_753             ( col_out_753             ),
    .col_out_754             ( col_out_754             ),
    .col_out_755             ( col_out_755             ),
    .col_out_756             ( col_out_756             ),
    .col_out_757             ( col_out_757             ),
    .col_out_758             ( col_out_758             ),
    .col_out_759             ( col_out_759             ),
    .col_out_760             ( col_out_760             ),
    .col_out_761             ( col_out_761             ),
    .col_out_762             ( col_out_762             ),
    .col_out_763             ( col_out_763             ),
    .col_out_764             ( col_out_764             ),
    .col_out_765             ( col_out_765             ),
    .col_out_766             ( col_out_766             ),
    .col_out_767             ( col_out_767             ),
    .col_out_768             ( col_out_768             ),
    .col_out_769             ( col_out_769             ),
    .col_out_770             ( col_out_770             ),
    .col_out_771             ( col_out_771             ),
    .col_out_772             ( col_out_772             ),
    .col_out_773             ( col_out_773             ),
    .col_out_774             ( col_out_774             ),
    .col_out_775             ( col_out_775             ),
    .col_out_776             ( col_out_776             ),
    .col_out_777             ( col_out_777             ),
    .col_out_778             ( col_out_778             ),
    .col_out_779             ( col_out_779             ),
    .col_out_780             ( col_out_780             ),
    .col_out_781             ( col_out_781             ),
    .col_out_782             ( col_out_782             ),
    .col_out_783             ( col_out_783             ),
    .col_out_784             ( col_out_784             ),
    .col_out_785             ( col_out_785             ),
    .col_out_786             ( col_out_786             ),
    .col_out_787             ( col_out_787             ),
    .col_out_788             ( col_out_788             ),
    .col_out_789             ( col_out_789             ),
    .col_out_790             ( col_out_790             ),
    .col_out_791             ( col_out_791             ),
    .col_out_792             ( col_out_792             ),
    .col_out_793             ( col_out_793             ),
    .col_out_794             ( col_out_794             ),
    .col_out_795             ( col_out_795             ),
    .col_out_796             ( col_out_796             ),
    .col_out_797             ( col_out_797             ),
    .col_out_798             ( col_out_798             ),
    .col_out_799             ( col_out_799             ),
    .col_out_800             ( col_out_800             ),
    .col_out_801             ( col_out_801             ),
    .col_out_802             ( col_out_802             ),
    .col_out_803             ( col_out_803             ),
    .col_out_804             ( col_out_804             ),
    .col_out_805             ( col_out_805             ),
    .col_out_806             ( col_out_806             ),
    .col_out_807             ( col_out_807             ),
    .col_out_808             ( col_out_808             ),
    .col_out_809             ( col_out_809             ),
    .col_out_810             ( col_out_810             ),
    .col_out_811             ( col_out_811             ),
    .col_out_812             ( col_out_812             ),
    .col_out_813             ( col_out_813             ),
    .col_out_814             ( col_out_814             ),
    .col_out_815             ( col_out_815             ),
    .col_out_816             ( col_out_816             ),
    .col_out_817             ( col_out_817             ),
    .col_out_818             ( col_out_818             ),
    .col_out_819             ( col_out_819             ),
    .col_out_820             ( col_out_820             ),
    .col_out_821             ( col_out_821             ),
    .col_out_822             ( col_out_822             ),
    .col_out_823             ( col_out_823             ),
    .col_out_824             ( col_out_824             ),
    .col_out_825             ( col_out_825             ),
    .col_out_826             ( col_out_826             ),
    .col_out_827             ( col_out_827             ),
    .col_out_828             ( col_out_828             ),
    .col_out_829             ( col_out_829             ),
    .col_out_830             ( col_out_830             ),
    .col_out_831             ( col_out_831             ),
    .col_out_832             ( col_out_832             ),
    .col_out_833             ( col_out_833             ),
    .col_out_834             ( col_out_834             ),
    .col_out_835             ( col_out_835             ),
    .col_out_836             ( col_out_836             ),
    .col_out_837             ( col_out_837             ),
    .col_out_838             ( col_out_838             ),
    .col_out_839             ( col_out_839             ),
    .col_out_840             ( col_out_840             ),
    .col_out_841             ( col_out_841             ),
    .col_out_842             ( col_out_842             ),
    .col_out_843             ( col_out_843             ),
    .col_out_844             ( col_out_844             ),
    .col_out_845             ( col_out_845             ),
    .col_out_846             ( col_out_846             ),
    .col_out_847             ( col_out_847             ),
    .col_out_848             ( col_out_848             ),
    .col_out_849             ( col_out_849             ),
    .col_out_850             ( col_out_850             ),
    .col_out_851             ( col_out_851             ),
    .col_out_852             ( col_out_852             ),
    .col_out_853             ( col_out_853             ),
    .col_out_854             ( col_out_854             ),
    .col_out_855             ( col_out_855             ),
    .col_out_856             ( col_out_856             ),
    .col_out_857             ( col_out_857             ),
    .col_out_858             ( col_out_858             ),
    .col_out_859             ( col_out_859             ),
    .col_out_860             ( col_out_860             ),
    .col_out_861             ( col_out_861             ),
    .col_out_862             ( col_out_862             ),
    .col_out_863             ( col_out_863             ),
    .col_out_864             ( col_out_864             ),
    .col_out_865             ( col_out_865             ),
    .col_out_866             ( col_out_866             ),
    .col_out_867             ( col_out_867             ),
    .col_out_868             ( col_out_868             ),
    .col_out_869             ( col_out_869             ),
    .col_out_870             ( col_out_870             ),
    .col_out_871             ( col_out_871             ),
    .col_out_872             ( col_out_872             ),
    .col_out_873             ( col_out_873             ),
    .col_out_874             ( col_out_874             ),
    .col_out_875             ( col_out_875             ),
    .col_out_876             ( col_out_876             ),
    .col_out_877             ( col_out_877             ),
    .col_out_878             ( col_out_878             ),
    .col_out_879             ( col_out_879             ),
    .col_out_880             ( col_out_880             ),
    .col_out_881             ( col_out_881             ),
    .col_out_882             ( col_out_882             ),
    .col_out_883             ( col_out_883             ),
    .col_out_884             ( col_out_884             ),
    .col_out_885             ( col_out_885             ),
    .col_out_886             ( col_out_886             ),
    .col_out_887             ( col_out_887             ),
    .col_out_888             ( col_out_888             ),
    .col_out_889             ( col_out_889             ),
    .col_out_890             ( col_out_890             ),
    .col_out_891             ( col_out_891             ),
    .col_out_892             ( col_out_892             ),
    .col_out_893             ( col_out_893             ),
    .col_out_894             ( col_out_894             ),
    .col_out_895             ( col_out_895             ),
    .col_out_896             ( col_out_896             ),
    .col_out_897             ( col_out_897             ),
    .col_out_898             ( col_out_898             ),
    .col_out_899             ( col_out_899             ),
    .col_out_900             ( col_out_900             ),
    .col_out_901             ( col_out_901             ),
    .col_out_902             ( col_out_902             ),
    .col_out_903             ( col_out_903             ),
    .col_out_904             ( col_out_904             ),
    .col_out_905             ( col_out_905             ),
    .col_out_906             ( col_out_906             ),
    .col_out_907             ( col_out_907             ),
    .col_out_908             ( col_out_908             ),
    .col_out_909             ( col_out_909             ),
    .col_out_910             ( col_out_910             ),
    .col_out_911             ( col_out_911             ),
    .col_out_912             ( col_out_912             ),
    .col_out_913             ( col_out_913             ),
    .col_out_914             ( col_out_914             ),
    .col_out_915             ( col_out_915             ),
    .col_out_916             ( col_out_916             ),
    .col_out_917             ( col_out_917             ),
    .col_out_918             ( col_out_918             ),
    .col_out_919             ( col_out_919             ),
    .col_out_920             ( col_out_920             ),
    .col_out_921             ( col_out_921             ),
    .col_out_922             ( col_out_922             ),
    .col_out_923             ( col_out_923             ),
    .col_out_924             ( col_out_924             ),
    .col_out_925             ( col_out_925             ),
    .col_out_926             ( col_out_926             ),
    .col_out_927             ( col_out_927             ),
    .col_out_928             ( col_out_928             ),
    .col_out_929             ( col_out_929             ),
    .col_out_930             ( col_out_930             ),
    .col_out_931             ( col_out_931             ),
    .col_out_932             ( col_out_932             ),
    .col_out_933             ( col_out_933             ),
    .col_out_934             ( col_out_934             ),
    .col_out_935             ( col_out_935             ),
    .col_out_936             ( col_out_936             ),
    .col_out_937             ( col_out_937             ),
    .col_out_938             ( col_out_938             ),
    .col_out_939             ( col_out_939             ),
    .col_out_940             ( col_out_940             ),
    .col_out_941             ( col_out_941             ),
    .col_out_942             ( col_out_942             ),
    .col_out_943             ( col_out_943             ),
    .col_out_944             ( col_out_944             ),
    .col_out_945             ( col_out_945             ),
    .col_out_946             ( col_out_946             ),
    .col_out_947             ( col_out_947             ),
    .col_out_948             ( col_out_948             ),
    .col_out_949             ( col_out_949             ),
    .col_out_950             ( col_out_950             ),
    .col_out_951             ( col_out_951             ),
    .col_out_952             ( col_out_952             ),
    .col_out_953             ( col_out_953             ),
    .col_out_954             ( col_out_954             ),
    .col_out_955             ( col_out_955             ),
    .col_out_956             ( col_out_956             ),
    .col_out_957             ( col_out_957             ),
    .col_out_958             ( col_out_958             ),
    .col_out_959             ( col_out_959             ),
    .col_out_960             ( col_out_960             ),
    .col_out_961             ( col_out_961             ),
    .col_out_962             ( col_out_962             ),
    .col_out_963             ( col_out_963             ),
    .col_out_964             ( col_out_964             ),
    .col_out_965             ( col_out_965             ),
    .col_out_966             ( col_out_966             ),
    .col_out_967             ( col_out_967             ),
    .col_out_968             ( col_out_968             ),
    .col_out_969             ( col_out_969             ),
    .col_out_970             ( col_out_970             ),
    .col_out_971             ( col_out_971             ),
    .col_out_972             ( col_out_972             ),
    .col_out_973             ( col_out_973             ),
    .col_out_974             ( col_out_974             ),
    .col_out_975             ( col_out_975             ),
    .col_out_976             ( col_out_976             ),
    .col_out_977             ( col_out_977             ),
    .col_out_978             ( col_out_978             ),
    .col_out_979             ( col_out_979             ),
    .col_out_980             ( col_out_980             ),
    .col_out_981             ( col_out_981             ),
    .col_out_982             ( col_out_982             ),
    .col_out_983             ( col_out_983             ),
    .col_out_984             ( col_out_984             ),
    .col_out_985             ( col_out_985             ),
    .col_out_986             ( col_out_986             ),
    .col_out_987             ( col_out_987             ),
    .col_out_988             ( col_out_988             ),
    .col_out_989             ( col_out_989             ),
    .col_out_990             ( col_out_990             ),
    .col_out_991             ( col_out_991             ),
    .col_out_992             ( col_out_992             ),
    .col_out_993             ( col_out_993             ),
    .col_out_994             ( col_out_994             ),
    .col_out_995             ( col_out_995             ),
    .col_out_996             ( col_out_996             ),
    .col_out_997             ( col_out_997             ),
    .col_out_998             ( col_out_998             ),
    .col_out_999             ( col_out_999             ),
    .col_out_1000            ( col_out_1000            ),
    .col_out_1001            ( col_out_1001            ),
    .col_out_1002            ( col_out_1002            ),
    .col_out_1003            ( col_out_1003            ),
    .col_out_1004            ( col_out_1004            ),
    .col_out_1005            ( col_out_1005            ),
    .col_out_1006            ( col_out_1006            ),
    .col_out_1007            ( col_out_1007            ),
    .col_out_1008            ( col_out_1008            ),
    .col_out_1009            ( col_out_1009            ),
    .col_out_1010            ( col_out_1010            ),
    .col_out_1011            ( col_out_1011            ),
    .col_out_1012            ( col_out_1012            ),
    .col_out_1013            ( col_out_1013            ),
    .col_out_1014            ( col_out_1014            ),
    .col_out_1015            ( col_out_1015            ),
    .col_out_1016            ( col_out_1016            ),
    .col_out_1017            ( col_out_1017            ),
    .col_out_1018            ( col_out_1018            ),
    .col_out_1019            ( col_out_1019            ),
    .col_out_1020            ( col_out_1020            ),
    .col_out_1021            ( col_out_1021            ),
    .col_out_1022            ( col_out_1022            ),
    .col_out_1023            ( col_out_1023            )
);







// alu Outputs
wire  [1032:0]  compressor_array_512_out0;
wire  [1032:0]  compressor_array_512_out1;
wire  [1024:0]  data_out_0;
wire  [1024:0]  data_out_1;

alu  u_alu (
    .col_in_0                ( col_out_0       ),
    .col_in_1                ( col_out_1       ),
    .col_in_2                ( col_out_2       ),
    .col_in_3                ( col_out_3       ),
    .col_in_4                ( col_out_4       ),
    .col_in_5                ( col_out_5       ),
    .col_in_6                ( col_out_6       ),
    .col_in_7                ( col_out_7       ),
    .col_in_8                ( col_out_8       ),
    .col_in_9                ( col_out_9       ),
    .col_in_10               ( col_out_10      ),
    .col_in_11               ( col_out_11      ),
    .col_in_12               ( col_out_12      ),
    .col_in_13               ( col_out_13      ),
    .col_in_14               ( col_out_14      ),
    .col_in_15               ( col_out_15      ),
    .col_in_16               ( col_out_16      ),
    .col_in_17               ( col_out_17      ),
    .col_in_18               ( col_out_18      ),
    .col_in_19               ( col_out_19      ),
    .col_in_20               ( col_out_20      ),
    .col_in_21               ( col_out_21      ),
    .col_in_22               ( col_out_22      ),
    .col_in_23               ( col_out_23      ),
    .col_in_24               ( col_out_24      ),
    .col_in_25               ( col_out_25      ),
    .col_in_26               ( col_out_26      ),
    .col_in_27               ( col_out_27      ),
    .col_in_28               ( col_out_28      ),
    .col_in_29               ( col_out_29      ),
    .col_in_30               ( col_out_30      ),
    .col_in_31               ( col_out_31      ),
    .col_in_32               ( col_out_32      ),
    .col_in_33               ( col_out_33      ),
    .col_in_34               ( col_out_34      ),
    .col_in_35               ( col_out_35      ),
    .col_in_36               ( col_out_36      ),
    .col_in_37               ( col_out_37      ),
    .col_in_38               ( col_out_38      ),
    .col_in_39               ( col_out_39      ),
    .col_in_40               ( col_out_40      ),
    .col_in_41               ( col_out_41      ),
    .col_in_42               ( col_out_42      ),
    .col_in_43               ( col_out_43      ),
    .col_in_44               ( col_out_44      ),
    .col_in_45               ( col_out_45      ),
    .col_in_46               ( col_out_46      ),
    .col_in_47               ( col_out_47      ),
    .col_in_48               ( col_out_48      ),
    .col_in_49               ( col_out_49      ),
    .col_in_50               ( col_out_50      ),
    .col_in_51               ( col_out_51      ),
    .col_in_52               ( col_out_52      ),
    .col_in_53               ( col_out_53      ),
    .col_in_54               ( col_out_54      ),
    .col_in_55               ( col_out_55      ),
    .col_in_56               ( col_out_56      ),
    .col_in_57               ( col_out_57      ),
    .col_in_58               ( col_out_58      ),
    .col_in_59               ( col_out_59      ),
    .col_in_60               ( col_out_60      ),
    .col_in_61               ( col_out_61      ),
    .col_in_62               ( col_out_62      ),
    .col_in_63               ( col_out_63      ),
    .col_in_64               ( col_out_64      ),
    .col_in_65               ( col_out_65      ),
    .col_in_66               ( col_out_66      ),
    .col_in_67               ( col_out_67      ),
    .col_in_68               ( col_out_68      ),
    .col_in_69               ( col_out_69      ),
    .col_in_70               ( col_out_70      ),
    .col_in_71               ( col_out_71      ),
    .col_in_72               ( col_out_72      ),
    .col_in_73               ( col_out_73      ),
    .col_in_74               ( col_out_74      ),
    .col_in_75               ( col_out_75      ),
    .col_in_76               ( col_out_76      ),
    .col_in_77               ( col_out_77      ),
    .col_in_78               ( col_out_78      ),
    .col_in_79               ( col_out_79      ),
    .col_in_80               ( col_out_80      ),
    .col_in_81               ( col_out_81      ),
    .col_in_82               ( col_out_82      ),
    .col_in_83               ( col_out_83      ),
    .col_in_84               ( col_out_84      ),
    .col_in_85               ( col_out_85      ),
    .col_in_86               ( col_out_86      ),
    .col_in_87               ( col_out_87      ),
    .col_in_88               ( col_out_88      ),
    .col_in_89               ( col_out_89      ),
    .col_in_90               ( col_out_90      ),
    .col_in_91               ( col_out_91      ),
    .col_in_92               ( col_out_92      ),
    .col_in_93               ( col_out_93      ),
    .col_in_94               ( col_out_94      ),
    .col_in_95               ( col_out_95      ),
    .col_in_96               ( col_out_96      ),
    .col_in_97               ( col_out_97      ),
    .col_in_98               ( col_out_98      ),
    .col_in_99               ( col_out_99      ),
    .col_in_100              ( col_out_100     ),
    .col_in_101              ( col_out_101     ),
    .col_in_102              ( col_out_102     ),
    .col_in_103              ( col_out_103     ),
    .col_in_104              ( col_out_104     ),
    .col_in_105              ( col_out_105     ),
    .col_in_106              ( col_out_106     ),
    .col_in_107              ( col_out_107     ),
    .col_in_108              ( col_out_108     ),
    .col_in_109              ( col_out_109     ),
    .col_in_110              ( col_out_110     ),
    .col_in_111              ( col_out_111     ),
    .col_in_112              ( col_out_112     ),
    .col_in_113              ( col_out_113     ),
    .col_in_114              ( col_out_114     ),
    .col_in_115              ( col_out_115     ),
    .col_in_116              ( col_out_116     ),
    .col_in_117              ( col_out_117     ),
    .col_in_118              ( col_out_118     ),
    .col_in_119              ( col_out_119     ),
    .col_in_120              ( col_out_120     ),
    .col_in_121              ( col_out_121     ),
    .col_in_122              ( col_out_122     ),
    .col_in_123              ( col_out_123     ),
    .col_in_124              ( col_out_124     ),
    .col_in_125              ( col_out_125     ),
    .col_in_126              ( col_out_126     ),
    .col_in_127              ( col_out_127     ),
    .col_in_128              ( col_out_128     ),
    .col_in_129              ( col_out_129     ),
    .col_in_130              ( col_out_130     ),
    .col_in_131              ( col_out_131     ),
    .col_in_132              ( col_out_132     ),
    .col_in_133              ( col_out_133     ),
    .col_in_134              ( col_out_134     ),
    .col_in_135              ( col_out_135     ),
    .col_in_136              ( col_out_136     ),
    .col_in_137              ( col_out_137     ),
    .col_in_138              ( col_out_138     ),
    .col_in_139              ( col_out_139     ),
    .col_in_140              ( col_out_140     ),
    .col_in_141              ( col_out_141     ),
    .col_in_142              ( col_out_142     ),
    .col_in_143              ( col_out_143     ),
    .col_in_144              ( col_out_144     ),
    .col_in_145              ( col_out_145     ),
    .col_in_146              ( col_out_146     ),
    .col_in_147              ( col_out_147     ),
    .col_in_148              ( col_out_148     ),
    .col_in_149              ( col_out_149     ),
    .col_in_150              ( col_out_150     ),
    .col_in_151              ( col_out_151     ),
    .col_in_152              ( col_out_152     ),
    .col_in_153              ( col_out_153     ),
    .col_in_154              ( col_out_154     ),
    .col_in_155              ( col_out_155     ),
    .col_in_156              ( col_out_156     ),
    .col_in_157              ( col_out_157     ),
    .col_in_158              ( col_out_158     ),
    .col_in_159              ( col_out_159     ),
    .col_in_160              ( col_out_160     ),
    .col_in_161              ( col_out_161     ),
    .col_in_162              ( col_out_162     ),
    .col_in_163              ( col_out_163     ),
    .col_in_164              ( col_out_164     ),
    .col_in_165              ( col_out_165     ),
    .col_in_166              ( col_out_166     ),
    .col_in_167              ( col_out_167     ),
    .col_in_168              ( col_out_168     ),
    .col_in_169              ( col_out_169     ),
    .col_in_170              ( col_out_170     ),
    .col_in_171              ( col_out_171     ),
    .col_in_172              ( col_out_172     ),
    .col_in_173              ( col_out_173     ),
    .col_in_174              ( col_out_174     ),
    .col_in_175              ( col_out_175     ),
    .col_in_176              ( col_out_176     ),
    .col_in_177              ( col_out_177     ),
    .col_in_178              ( col_out_178     ),
    .col_in_179              ( col_out_179     ),
    .col_in_180              ( col_out_180     ),
    .col_in_181              ( col_out_181     ),
    .col_in_182              ( col_out_182     ),
    .col_in_183              ( col_out_183     ),
    .col_in_184              ( col_out_184     ),
    .col_in_185              ( col_out_185     ),
    .col_in_186              ( col_out_186     ),
    .col_in_187              ( col_out_187     ),
    .col_in_188              ( col_out_188     ),
    .col_in_189              ( col_out_189     ),
    .col_in_190              ( col_out_190     ),
    .col_in_191              ( col_out_191     ),
    .col_in_192              ( col_out_192     ),
    .col_in_193              ( col_out_193     ),
    .col_in_194              ( col_out_194     ),
    .col_in_195              ( col_out_195     ),
    .col_in_196              ( col_out_196     ),
    .col_in_197              ( col_out_197     ),
    .col_in_198              ( col_out_198     ),
    .col_in_199              ( col_out_199     ),
    .col_in_200              ( col_out_200     ),
    .col_in_201              ( col_out_201     ),
    .col_in_202              ( col_out_202     ),
    .col_in_203              ( col_out_203     ),
    .col_in_204              ( col_out_204     ),
    .col_in_205              ( col_out_205     ),
    .col_in_206              ( col_out_206     ),
    .col_in_207              ( col_out_207     ),
    .col_in_208              ( col_out_208     ),
    .col_in_209              ( col_out_209     ),
    .col_in_210              ( col_out_210     ),
    .col_in_211              ( col_out_211     ),
    .col_in_212              ( col_out_212     ),
    .col_in_213              ( col_out_213     ),
    .col_in_214              ( col_out_214     ),
    .col_in_215              ( col_out_215     ),
    .col_in_216              ( col_out_216     ),
    .col_in_217              ( col_out_217     ),
    .col_in_218              ( col_out_218     ),
    .col_in_219              ( col_out_219     ),
    .col_in_220              ( col_out_220     ),
    .col_in_221              ( col_out_221     ),
    .col_in_222              ( col_out_222     ),
    .col_in_223              ( col_out_223     ),
    .col_in_224              ( col_out_224     ),
    .col_in_225              ( col_out_225     ),
    .col_in_226              ( col_out_226     ),
    .col_in_227              ( col_out_227     ),
    .col_in_228              ( col_out_228     ),
    .col_in_229              ( col_out_229     ),
    .col_in_230              ( col_out_230     ),
    .col_in_231              ( col_out_231     ),
    .col_in_232              ( col_out_232     ),
    .col_in_233              ( col_out_233     ),
    .col_in_234              ( col_out_234     ),
    .col_in_235              ( col_out_235     ),
    .col_in_236              ( col_out_236     ),
    .col_in_237              ( col_out_237     ),
    .col_in_238              ( col_out_238     ),
    .col_in_239              ( col_out_239     ),
    .col_in_240              ( col_out_240     ),
    .col_in_241              ( col_out_241     ),
    .col_in_242              ( col_out_242     ),
    .col_in_243              ( col_out_243     ),
    .col_in_244              ( col_out_244     ),
    .col_in_245              ( col_out_245     ),
    .col_in_246              ( col_out_246     ),
    .col_in_247              ( col_out_247     ),
    .col_in_248              ( col_out_248     ),
    .col_in_249              ( col_out_249     ),
    .col_in_250              ( col_out_250     ),
    .col_in_251              ( col_out_251     ),
    .col_in_252              ( col_out_252     ),
    .col_in_253              ( col_out_253     ),
    .col_in_254              ( col_out_254     ),
    .col_in_255              ( col_out_255     ),
    .col_in_256              ( col_out_256     ),
    .col_in_257              ( col_out_257     ),
    .col_in_258              ( col_out_258     ),
    .col_in_259              ( col_out_259     ),
    .col_in_260              ( col_out_260     ),
    .col_in_261              ( col_out_261     ),
    .col_in_262              ( col_out_262     ),
    .col_in_263              ( col_out_263     ),
    .col_in_264              ( col_out_264     ),
    .col_in_265              ( col_out_265     ),
    .col_in_266              ( col_out_266     ),
    .col_in_267              ( col_out_267     ),
    .col_in_268              ( col_out_268     ),
    .col_in_269              ( col_out_269     ),
    .col_in_270              ( col_out_270     ),
    .col_in_271              ( col_out_271     ),
    .col_in_272              ( col_out_272     ),
    .col_in_273              ( col_out_273     ),
    .col_in_274              ( col_out_274     ),
    .col_in_275              ( col_out_275     ),
    .col_in_276              ( col_out_276     ),
    .col_in_277              ( col_out_277     ),
    .col_in_278              ( col_out_278     ),
    .col_in_279              ( col_out_279     ),
    .col_in_280              ( col_out_280     ),
    .col_in_281              ( col_out_281     ),
    .col_in_282              ( col_out_282     ),
    .col_in_283              ( col_out_283     ),
    .col_in_284              ( col_out_284     ),
    .col_in_285              ( col_out_285     ),
    .col_in_286              ( col_out_286     ),
    .col_in_287              ( col_out_287     ),
    .col_in_288              ( col_out_288     ),
    .col_in_289              ( col_out_289     ),
    .col_in_290              ( col_out_290     ),
    .col_in_291              ( col_out_291     ),
    .col_in_292              ( col_out_292     ),
    .col_in_293              ( col_out_293     ),
    .col_in_294              ( col_out_294     ),
    .col_in_295              ( col_out_295     ),
    .col_in_296              ( col_out_296     ),
    .col_in_297              ( col_out_297     ),
    .col_in_298              ( col_out_298     ),
    .col_in_299              ( col_out_299     ),
    .col_in_300              ( col_out_300     ),
    .col_in_301              ( col_out_301     ),
    .col_in_302              ( col_out_302     ),
    .col_in_303              ( col_out_303     ),
    .col_in_304              ( col_out_304     ),
    .col_in_305              ( col_out_305     ),
    .col_in_306              ( col_out_306     ),
    .col_in_307              ( col_out_307     ),
    .col_in_308              ( col_out_308     ),
    .col_in_309              ( col_out_309     ),
    .col_in_310              ( col_out_310     ),
    .col_in_311              ( col_out_311     ),
    .col_in_312              ( col_out_312     ),
    .col_in_313              ( col_out_313     ),
    .col_in_314              ( col_out_314     ),
    .col_in_315              ( col_out_315     ),
    .col_in_316              ( col_out_316     ),
    .col_in_317              ( col_out_317     ),
    .col_in_318              ( col_out_318     ),
    .col_in_319              ( col_out_319     ),
    .col_in_320              ( col_out_320     ),
    .col_in_321              ( col_out_321     ),
    .col_in_322              ( col_out_322     ),
    .col_in_323              ( col_out_323     ),
    .col_in_324              ( col_out_324     ),
    .col_in_325              ( col_out_325     ),
    .col_in_326              ( col_out_326     ),
    .col_in_327              ( col_out_327     ),
    .col_in_328              ( col_out_328     ),
    .col_in_329              ( col_out_329     ),
    .col_in_330              ( col_out_330     ),
    .col_in_331              ( col_out_331     ),
    .col_in_332              ( col_out_332     ),
    .col_in_333              ( col_out_333     ),
    .col_in_334              ( col_out_334     ),
    .col_in_335              ( col_out_335     ),
    .col_in_336              ( col_out_336     ),
    .col_in_337              ( col_out_337     ),
    .col_in_338              ( col_out_338     ),
    .col_in_339              ( col_out_339     ),
    .col_in_340              ( col_out_340     ),
    .col_in_341              ( col_out_341     ),
    .col_in_342              ( col_out_342     ),
    .col_in_343              ( col_out_343     ),
    .col_in_344              ( col_out_344     ),
    .col_in_345              ( col_out_345     ),
    .col_in_346              ( col_out_346     ),
    .col_in_347              ( col_out_347     ),
    .col_in_348              ( col_out_348     ),
    .col_in_349              ( col_out_349     ),
    .col_in_350              ( col_out_350     ),
    .col_in_351              ( col_out_351     ),
    .col_in_352              ( col_out_352     ),
    .col_in_353              ( col_out_353     ),
    .col_in_354              ( col_out_354     ),
    .col_in_355              ( col_out_355     ),
    .col_in_356              ( col_out_356     ),
    .col_in_357              ( col_out_357     ),
    .col_in_358              ( col_out_358     ),
    .col_in_359              ( col_out_359     ),
    .col_in_360              ( col_out_360     ),
    .col_in_361              ( col_out_361     ),
    .col_in_362              ( col_out_362     ),
    .col_in_363              ( col_out_363     ),
    .col_in_364              ( col_out_364     ),
    .col_in_365              ( col_out_365     ),
    .col_in_366              ( col_out_366     ),
    .col_in_367              ( col_out_367     ),
    .col_in_368              ( col_out_368     ),
    .col_in_369              ( col_out_369     ),
    .col_in_370              ( col_out_370     ),
    .col_in_371              ( col_out_371     ),
    .col_in_372              ( col_out_372     ),
    .col_in_373              ( col_out_373     ),
    .col_in_374              ( col_out_374     ),
    .col_in_375              ( col_out_375     ),
    .col_in_376              ( col_out_376     ),
    .col_in_377              ( col_out_377     ),
    .col_in_378              ( col_out_378     ),
    .col_in_379              ( col_out_379     ),
    .col_in_380              ( col_out_380     ),
    .col_in_381              ( col_out_381     ),
    .col_in_382              ( col_out_382     ),
    .col_in_383              ( col_out_383     ),
    .col_in_384              ( col_out_384     ),
    .col_in_385              ( col_out_385     ),
    .col_in_386              ( col_out_386     ),
    .col_in_387              ( col_out_387     ),
    .col_in_388              ( col_out_388     ),
    .col_in_389              ( col_out_389     ),
    .col_in_390              ( col_out_390     ),
    .col_in_391              ( col_out_391     ),
    .col_in_392              ( col_out_392     ),
    .col_in_393              ( col_out_393     ),
    .col_in_394              ( col_out_394     ),
    .col_in_395              ( col_out_395     ),
    .col_in_396              ( col_out_396     ),
    .col_in_397              ( col_out_397     ),
    .col_in_398              ( col_out_398     ),
    .col_in_399              ( col_out_399     ),
    .col_in_400              ( col_out_400     ),
    .col_in_401              ( col_out_401     ),
    .col_in_402              ( col_out_402     ),
    .col_in_403              ( col_out_403     ),
    .col_in_404              ( col_out_404     ),
    .col_in_405              ( col_out_405     ),
    .col_in_406              ( col_out_406     ),
    .col_in_407              ( col_out_407     ),
    .col_in_408              ( col_out_408     ),
    .col_in_409              ( col_out_409     ),
    .col_in_410              ( col_out_410     ),
    .col_in_411              ( col_out_411     ),
    .col_in_412              ( col_out_412     ),
    .col_in_413              ( col_out_413     ),
    .col_in_414              ( col_out_414     ),
    .col_in_415              ( col_out_415     ),
    .col_in_416              ( col_out_416     ),
    .col_in_417              ( col_out_417     ),
    .col_in_418              ( col_out_418     ),
    .col_in_419              ( col_out_419     ),
    .col_in_420              ( col_out_420     ),
    .col_in_421              ( col_out_421     ),
    .col_in_422              ( col_out_422     ),
    .col_in_423              ( col_out_423     ),
    .col_in_424              ( col_out_424     ),
    .col_in_425              ( col_out_425     ),
    .col_in_426              ( col_out_426     ),
    .col_in_427              ( col_out_427     ),
    .col_in_428              ( col_out_428     ),
    .col_in_429              ( col_out_429     ),
    .col_in_430              ( col_out_430     ),
    .col_in_431              ( col_out_431     ),
    .col_in_432              ( col_out_432     ),
    .col_in_433              ( col_out_433     ),
    .col_in_434              ( col_out_434     ),
    .col_in_435              ( col_out_435     ),
    .col_in_436              ( col_out_436     ),
    .col_in_437              ( col_out_437     ),
    .col_in_438              ( col_out_438     ),
    .col_in_439              ( col_out_439     ),
    .col_in_440              ( col_out_440     ),
    .col_in_441              ( col_out_441     ),
    .col_in_442              ( col_out_442     ),
    .col_in_443              ( col_out_443     ),
    .col_in_444              ( col_out_444     ),
    .col_in_445              ( col_out_445     ),
    .col_in_446              ( col_out_446     ),
    .col_in_447              ( col_out_447     ),
    .col_in_448              ( col_out_448     ),
    .col_in_449              ( col_out_449     ),
    .col_in_450              ( col_out_450     ),
    .col_in_451              ( col_out_451     ),
    .col_in_452              ( col_out_452     ),
    .col_in_453              ( col_out_453     ),
    .col_in_454              ( col_out_454     ),
    .col_in_455              ( col_out_455     ),
    .col_in_456              ( col_out_456     ),
    .col_in_457              ( col_out_457     ),
    .col_in_458              ( col_out_458     ),
    .col_in_459              ( col_out_459     ),
    .col_in_460              ( col_out_460     ),
    .col_in_461              ( col_out_461     ),
    .col_in_462              ( col_out_462     ),
    .col_in_463              ( col_out_463     ),
    .col_in_464              ( col_out_464     ),
    .col_in_465              ( col_out_465     ),
    .col_in_466              ( col_out_466     ),
    .col_in_467              ( col_out_467     ),
    .col_in_468              ( col_out_468     ),
    .col_in_469              ( col_out_469     ),
    .col_in_470              ( col_out_470     ),
    .col_in_471              ( col_out_471     ),
    .col_in_472              ( col_out_472     ),
    .col_in_473              ( col_out_473     ),
    .col_in_474              ( col_out_474     ),
    .col_in_475              ( col_out_475     ),
    .col_in_476              ( col_out_476     ),
    .col_in_477              ( col_out_477     ),
    .col_in_478              ( col_out_478     ),
    .col_in_479              ( col_out_479     ),
    .col_in_480              ( col_out_480     ),
    .col_in_481              ( col_out_481     ),
    .col_in_482              ( col_out_482     ),
    .col_in_483              ( col_out_483     ),
    .col_in_484              ( col_out_484     ),
    .col_in_485              ( col_out_485     ),
    .col_in_486              ( col_out_486     ),
    .col_in_487              ( col_out_487     ),
    .col_in_488              ( col_out_488     ),
    .col_in_489              ( col_out_489     ),
    .col_in_490              ( col_out_490     ),
    .col_in_491              ( col_out_491     ),
    .col_in_492              ( col_out_492     ),
    .col_in_493              ( col_out_493     ),
    .col_in_494              ( col_out_494     ),
    .col_in_495              ( col_out_495     ),
    .col_in_496              ( col_out_496     ),
    .col_in_497              ( col_out_497     ),
    .col_in_498              ( col_out_498     ),
    .col_in_499              ( col_out_499     ),
    .col_in_500              ( col_out_500     ),
    .col_in_501              ( col_out_501     ),
    .col_in_502              ( col_out_502     ),
    .col_in_503              ( col_out_503     ),
    .col_in_504              ( col_out_504     ),
    .col_in_505              ( col_out_505     ),
    .col_in_506              ( col_out_506     ),
    .col_in_507              ( col_out_507     ),
    .col_in_508              ( col_out_508     ),
    .col_in_509              ( col_out_509     ),
    .col_in_510              ( col_out_510     ),
    .col_in_511              ( col_out_511     ),
    .col_in_512              ( col_out_512     ),
    .col_in_513              ( col_out_513     ),
    .col_in_514              ( col_out_514     ),
    .col_in_515              ( col_out_515     ),
    .col_in_516              ( col_out_516     ),
    .col_in_517              ( col_out_517     ),
    .col_in_518              ( col_out_518     ),
    .col_in_519              ( col_out_519     ),
    .col_in_520              ( col_out_520     ),
    .col_in_521              ( col_out_521     ),
    .col_in_522              ( col_out_522     ),
    .col_in_523              ( col_out_523     ),
    .col_in_524              ( col_out_524     ),
    .col_in_525              ( col_out_525     ),
    .col_in_526              ( col_out_526     ),
    .col_in_527              ( col_out_527     ),
    .col_in_528              ( col_out_528     ),
    .col_in_529              ( col_out_529     ),
    .col_in_530              ( col_out_530     ),
    .col_in_531              ( col_out_531     ),
    .col_in_532              ( col_out_532     ),
    .col_in_533              ( col_out_533     ),
    .col_in_534              ( col_out_534     ),
    .col_in_535              ( col_out_535     ),
    .col_in_536              ( col_out_536     ),
    .col_in_537              ( col_out_537     ),
    .col_in_538              ( col_out_538     ),
    .col_in_539              ( col_out_539     ),
    .col_in_540              ( col_out_540     ),
    .col_in_541              ( col_out_541     ),
    .col_in_542              ( col_out_542     ),
    .col_in_543              ( col_out_543     ),
    .col_in_544              ( col_out_544     ),
    .col_in_545              ( col_out_545     ),
    .col_in_546              ( col_out_546     ),
    .col_in_547              ( col_out_547     ),
    .col_in_548              ( col_out_548     ),
    .col_in_549              ( col_out_549     ),
    .col_in_550              ( col_out_550     ),
    .col_in_551              ( col_out_551     ),
    .col_in_552              ( col_out_552     ),
    .col_in_553              ( col_out_553     ),
    .col_in_554              ( col_out_554     ),
    .col_in_555              ( col_out_555     ),
    .col_in_556              ( col_out_556     ),
    .col_in_557              ( col_out_557     ),
    .col_in_558              ( col_out_558     ),
    .col_in_559              ( col_out_559     ),
    .col_in_560              ( col_out_560     ),
    .col_in_561              ( col_out_561     ),
    .col_in_562              ( col_out_562     ),
    .col_in_563              ( col_out_563     ),
    .col_in_564              ( col_out_564     ),
    .col_in_565              ( col_out_565     ),
    .col_in_566              ( col_out_566     ),
    .col_in_567              ( col_out_567     ),
    .col_in_568              ( col_out_568     ),
    .col_in_569              ( col_out_569     ),
    .col_in_570              ( col_out_570     ),
    .col_in_571              ( col_out_571     ),
    .col_in_572              ( col_out_572     ),
    .col_in_573              ( col_out_573     ),
    .col_in_574              ( col_out_574     ),
    .col_in_575              ( col_out_575     ),
    .col_in_576              ( col_out_576     ),
    .col_in_577              ( col_out_577     ),
    .col_in_578              ( col_out_578     ),
    .col_in_579              ( col_out_579     ),
    .col_in_580              ( col_out_580     ),
    .col_in_581              ( col_out_581     ),
    .col_in_582              ( col_out_582     ),
    .col_in_583              ( col_out_583     ),
    .col_in_584              ( col_out_584     ),
    .col_in_585              ( col_out_585     ),
    .col_in_586              ( col_out_586     ),
    .col_in_587              ( col_out_587     ),
    .col_in_588              ( col_out_588     ),
    .col_in_589              ( col_out_589     ),
    .col_in_590              ( col_out_590     ),
    .col_in_591              ( col_out_591     ),
    .col_in_592              ( col_out_592     ),
    .col_in_593              ( col_out_593     ),
    .col_in_594              ( col_out_594     ),
    .col_in_595              ( col_out_595     ),
    .col_in_596              ( col_out_596     ),
    .col_in_597              ( col_out_597     ),
    .col_in_598              ( col_out_598     ),
    .col_in_599              ( col_out_599     ),
    .col_in_600              ( col_out_600     ),
    .col_in_601              ( col_out_601     ),
    .col_in_602              ( col_out_602     ),
    .col_in_603              ( col_out_603     ),
    .col_in_604              ( col_out_604     ),
    .col_in_605              ( col_out_605     ),
    .col_in_606              ( col_out_606     ),
    .col_in_607              ( col_out_607     ),
    .col_in_608              ( col_out_608     ),
    .col_in_609              ( col_out_609     ),
    .col_in_610              ( col_out_610     ),
    .col_in_611              ( col_out_611     ),
    .col_in_612              ( col_out_612     ),
    .col_in_613              ( col_out_613     ),
    .col_in_614              ( col_out_614     ),
    .col_in_615              ( col_out_615     ),
    .col_in_616              ( col_out_616     ),
    .col_in_617              ( col_out_617     ),
    .col_in_618              ( col_out_618     ),
    .col_in_619              ( col_out_619     ),
    .col_in_620              ( col_out_620     ),
    .col_in_621              ( col_out_621     ),
    .col_in_622              ( col_out_622     ),
    .col_in_623              ( col_out_623     ),
    .col_in_624              ( col_out_624     ),
    .col_in_625              ( col_out_625     ),
    .col_in_626              ( col_out_626     ),
    .col_in_627              ( col_out_627     ),
    .col_in_628              ( col_out_628     ),
    .col_in_629              ( col_out_629     ),
    .col_in_630              ( col_out_630     ),
    .col_in_631              ( col_out_631     ),
    .col_in_632              ( col_out_632     ),
    .col_in_633              ( col_out_633     ),
    .col_in_634              ( col_out_634     ),
    .col_in_635              ( col_out_635     ),
    .col_in_636              ( col_out_636     ),
    .col_in_637              ( col_out_637     ),
    .col_in_638              ( col_out_638     ),
    .col_in_639              ( col_out_639     ),
    .col_in_640              ( col_out_640     ),
    .col_in_641              ( col_out_641     ),
    .col_in_642              ( col_out_642     ),
    .col_in_643              ( col_out_643     ),
    .col_in_644              ( col_out_644     ),
    .col_in_645              ( col_out_645     ),
    .col_in_646              ( col_out_646     ),
    .col_in_647              ( col_out_647     ),
    .col_in_648              ( col_out_648     ),
    .col_in_649              ( col_out_649     ),
    .col_in_650              ( col_out_650     ),
    .col_in_651              ( col_out_651     ),
    .col_in_652              ( col_out_652     ),
    .col_in_653              ( col_out_653     ),
    .col_in_654              ( col_out_654     ),
    .col_in_655              ( col_out_655     ),
    .col_in_656              ( col_out_656     ),
    .col_in_657              ( col_out_657     ),
    .col_in_658              ( col_out_658     ),
    .col_in_659              ( col_out_659     ),
    .col_in_660              ( col_out_660     ),
    .col_in_661              ( col_out_661     ),
    .col_in_662              ( col_out_662     ),
    .col_in_663              ( col_out_663     ),
    .col_in_664              ( col_out_664     ),
    .col_in_665              ( col_out_665     ),
    .col_in_666              ( col_out_666     ),
    .col_in_667              ( col_out_667     ),
    .col_in_668              ( col_out_668     ),
    .col_in_669              ( col_out_669     ),
    .col_in_670              ( col_out_670     ),
    .col_in_671              ( col_out_671     ),
    .col_in_672              ( col_out_672     ),
    .col_in_673              ( col_out_673     ),
    .col_in_674              ( col_out_674     ),
    .col_in_675              ( col_out_675     ),
    .col_in_676              ( col_out_676     ),
    .col_in_677              ( col_out_677     ),
    .col_in_678              ( col_out_678     ),
    .col_in_679              ( col_out_679     ),
    .col_in_680              ( col_out_680     ),
    .col_in_681              ( col_out_681     ),
    .col_in_682              ( col_out_682     ),
    .col_in_683              ( col_out_683     ),
    .col_in_684              ( col_out_684     ),
    .col_in_685              ( col_out_685     ),
    .col_in_686              ( col_out_686     ),
    .col_in_687              ( col_out_687     ),
    .col_in_688              ( col_out_688     ),
    .col_in_689              ( col_out_689     ),
    .col_in_690              ( col_out_690     ),
    .col_in_691              ( col_out_691     ),
    .col_in_692              ( col_out_692     ),
    .col_in_693              ( col_out_693     ),
    .col_in_694              ( col_out_694     ),
    .col_in_695              ( col_out_695     ),
    .col_in_696              ( col_out_696     ),
    .col_in_697              ( col_out_697     ),
    .col_in_698              ( col_out_698     ),
    .col_in_699              ( col_out_699     ),
    .col_in_700              ( col_out_700     ),
    .col_in_701              ( col_out_701     ),
    .col_in_702              ( col_out_702     ),
    .col_in_703              ( col_out_703     ),
    .col_in_704              ( col_out_704     ),
    .col_in_705              ( col_out_705     ),
    .col_in_706              ( col_out_706     ),
    .col_in_707              ( col_out_707     ),
    .col_in_708              ( col_out_708     ),
    .col_in_709              ( col_out_709     ),
    .col_in_710              ( col_out_710     ),
    .col_in_711              ( col_out_711     ),
    .col_in_712              ( col_out_712     ),
    .col_in_713              ( col_out_713     ),
    .col_in_714              ( col_out_714     ),
    .col_in_715              ( col_out_715     ),
    .col_in_716              ( col_out_716     ),
    .col_in_717              ( col_out_717     ),
    .col_in_718              ( col_out_718     ),
    .col_in_719              ( col_out_719     ),
    .col_in_720              ( col_out_720     ),
    .col_in_721              ( col_out_721     ),
    .col_in_722              ( col_out_722     ),
    .col_in_723              ( col_out_723     ),
    .col_in_724              ( col_out_724     ),
    .col_in_725              ( col_out_725     ),
    .col_in_726              ( col_out_726     ),
    .col_in_727              ( col_out_727     ),
    .col_in_728              ( col_out_728     ),
    .col_in_729              ( col_out_729     ),
    .col_in_730              ( col_out_730     ),
    .col_in_731              ( col_out_731     ),
    .col_in_732              ( col_out_732     ),
    .col_in_733              ( col_out_733     ),
    .col_in_734              ( col_out_734     ),
    .col_in_735              ( col_out_735     ),
    .col_in_736              ( col_out_736     ),
    .col_in_737              ( col_out_737     ),
    .col_in_738              ( col_out_738     ),
    .col_in_739              ( col_out_739     ),
    .col_in_740              ( col_out_740     ),
    .col_in_741              ( col_out_741     ),
    .col_in_742              ( col_out_742     ),
    .col_in_743              ( col_out_743     ),
    .col_in_744              ( col_out_744     ),
    .col_in_745              ( col_out_745     ),
    .col_in_746              ( col_out_746     ),
    .col_in_747              ( col_out_747     ),
    .col_in_748              ( col_out_748     ),
    .col_in_749              ( col_out_749     ),
    .col_in_750              ( col_out_750     ),
    .col_in_751              ( col_out_751     ),
    .col_in_752              ( col_out_752     ),
    .col_in_753              ( col_out_753     ),
    .col_in_754              ( col_out_754     ),
    .col_in_755              ( col_out_755     ),
    .col_in_756              ( col_out_756     ),
    .col_in_757              ( col_out_757     ),
    .col_in_758              ( col_out_758     ),
    .col_in_759              ( col_out_759     ),
    .col_in_760              ( col_out_760     ),
    .col_in_761              ( col_out_761     ),
    .col_in_762              ( col_out_762     ),
    .col_in_763              ( col_out_763     ),
    .col_in_764              ( col_out_764     ),
    .col_in_765              ( col_out_765     ),
    .col_in_766              ( col_out_766     ),
    .col_in_767              ( col_out_767     ),
    .col_in_768              ( col_out_768     ),
    .col_in_769              ( col_out_769     ),
    .col_in_770              ( col_out_770     ),
    .col_in_771              ( col_out_771     ),
    .col_in_772              ( col_out_772     ),
    .col_in_773              ( col_out_773     ),
    .col_in_774              ( col_out_774     ),
    .col_in_775              ( col_out_775     ),
    .col_in_776              ( col_out_776     ),
    .col_in_777              ( col_out_777     ),
    .col_in_778              ( col_out_778     ),
    .col_in_779              ( col_out_779     ),
    .col_in_780              ( col_out_780     ),
    .col_in_781              ( col_out_781     ),
    .col_in_782              ( col_out_782     ),
    .col_in_783              ( col_out_783     ),
    .col_in_784              ( col_out_784     ),
    .col_in_785              ( col_out_785     ),
    .col_in_786              ( col_out_786     ),
    .col_in_787              ( col_out_787     ),
    .col_in_788              ( col_out_788     ),
    .col_in_789              ( col_out_789     ),
    .col_in_790              ( col_out_790     ),
    .col_in_791              ( col_out_791     ),
    .col_in_792              ( col_out_792     ),
    .col_in_793              ( col_out_793     ),
    .col_in_794              ( col_out_794     ),
    .col_in_795              ( col_out_795     ),
    .col_in_796              ( col_out_796     ),
    .col_in_797              ( col_out_797     ),
    .col_in_798              ( col_out_798     ),
    .col_in_799              ( col_out_799     ),
    .col_in_800              ( col_out_800     ),
    .col_in_801              ( col_out_801     ),
    .col_in_802              ( col_out_802     ),
    .col_in_803              ( col_out_803     ),
    .col_in_804              ( col_out_804     ),
    .col_in_805              ( col_out_805     ),
    .col_in_806              ( col_out_806     ),
    .col_in_807              ( col_out_807     ),
    .col_in_808              ( col_out_808     ),
    .col_in_809              ( col_out_809     ),
    .col_in_810              ( col_out_810     ),
    .col_in_811              ( col_out_811     ),
    .col_in_812              ( col_out_812     ),
    .col_in_813              ( col_out_813     ),
    .col_in_814              ( col_out_814     ),
    .col_in_815              ( col_out_815     ),
    .col_in_816              ( col_out_816     ),
    .col_in_817              ( col_out_817     ),
    .col_in_818              ( col_out_818     ),
    .col_in_819              ( col_out_819     ),
    .col_in_820              ( col_out_820     ),
    .col_in_821              ( col_out_821     ),
    .col_in_822              ( col_out_822     ),
    .col_in_823              ( col_out_823     ),
    .col_in_824              ( col_out_824     ),
    .col_in_825              ( col_out_825     ),
    .col_in_826              ( col_out_826     ),
    .col_in_827              ( col_out_827     ),
    .col_in_828              ( col_out_828     ),
    .col_in_829              ( col_out_829     ),
    .col_in_830              ( col_out_830     ),
    .col_in_831              ( col_out_831     ),
    .col_in_832              ( col_out_832     ),
    .col_in_833              ( col_out_833     ),
    .col_in_834              ( col_out_834     ),
    .col_in_835              ( col_out_835     ),
    .col_in_836              ( col_out_836     ),
    .col_in_837              ( col_out_837     ),
    .col_in_838              ( col_out_838     ),
    .col_in_839              ( col_out_839     ),
    .col_in_840              ( col_out_840     ),
    .col_in_841              ( col_out_841     ),
    .col_in_842              ( col_out_842     ),
    .col_in_843              ( col_out_843     ),
    .col_in_844              ( col_out_844     ),
    .col_in_845              ( col_out_845     ),
    .col_in_846              ( col_out_846     ),
    .col_in_847              ( col_out_847     ),
    .col_in_848              ( col_out_848     ),
    .col_in_849              ( col_out_849     ),
    .col_in_850              ( col_out_850     ),
    .col_in_851              ( col_out_851     ),
    .col_in_852              ( col_out_852     ),
    .col_in_853              ( col_out_853     ),
    .col_in_854              ( col_out_854     ),
    .col_in_855              ( col_out_855     ),
    .col_in_856              ( col_out_856     ),
    .col_in_857              ( col_out_857     ),
    .col_in_858              ( col_out_858     ),
    .col_in_859              ( col_out_859     ),
    .col_in_860              ( col_out_860     ),
    .col_in_861              ( col_out_861     ),
    .col_in_862              ( col_out_862     ),
    .col_in_863              ( col_out_863     ),
    .col_in_864              ( col_out_864     ),
    .col_in_865              ( col_out_865     ),
    .col_in_866              ( col_out_866     ),
    .col_in_867              ( col_out_867     ),
    .col_in_868              ( col_out_868     ),
    .col_in_869              ( col_out_869     ),
    .col_in_870              ( col_out_870     ),
    .col_in_871              ( col_out_871     ),
    .col_in_872              ( col_out_872     ),
    .col_in_873              ( col_out_873     ),
    .col_in_874              ( col_out_874     ),
    .col_in_875              ( col_out_875     ),
    .col_in_876              ( col_out_876     ),
    .col_in_877              ( col_out_877     ),
    .col_in_878              ( col_out_878     ),
    .col_in_879              ( col_out_879     ),
    .col_in_880              ( col_out_880     ),
    .col_in_881              ( col_out_881     ),
    .col_in_882              ( col_out_882     ),
    .col_in_883              ( col_out_883     ),
    .col_in_884              ( col_out_884     ),
    .col_in_885              ( col_out_885     ),
    .col_in_886              ( col_out_886     ),
    .col_in_887              ( col_out_887     ),
    .col_in_888              ( col_out_888     ),
    .col_in_889              ( col_out_889     ),
    .col_in_890              ( col_out_890     ),
    .col_in_891              ( col_out_891     ),
    .col_in_892              ( col_out_892     ),
    .col_in_893              ( col_out_893     ),
    .col_in_894              ( col_out_894     ),
    .col_in_895              ( col_out_895     ),
    .col_in_896              ( col_out_896     ),
    .col_in_897              ( col_out_897     ),
    .col_in_898              ( col_out_898     ),
    .col_in_899              ( col_out_899     ),
    .col_in_900              ( col_out_900     ),
    .col_in_901              ( col_out_901     ),
    .col_in_902              ( col_out_902     ),
    .col_in_903              ( col_out_903     ),
    .col_in_904              ( col_out_904     ),
    .col_in_905              ( col_out_905     ),
    .col_in_906              ( col_out_906     ),
    .col_in_907              ( col_out_907     ),
    .col_in_908              ( col_out_908     ),
    .col_in_909              ( col_out_909     ),
    .col_in_910              ( col_out_910     ),
    .col_in_911              ( col_out_911     ),
    .col_in_912              ( col_out_912     ),
    .col_in_913              ( col_out_913     ),
    .col_in_914              ( col_out_914     ),
    .col_in_915              ( col_out_915     ),
    .col_in_916              ( col_out_916     ),
    .col_in_917              ( col_out_917     ),
    .col_in_918              ( col_out_918     ),
    .col_in_919              ( col_out_919     ),
    .col_in_920              ( col_out_920     ),
    .col_in_921              ( col_out_921     ),
    .col_in_922              ( col_out_922     ),
    .col_in_923              ( col_out_923     ),
    .col_in_924              ( col_out_924     ),
    .col_in_925              ( col_out_925     ),
    .col_in_926              ( col_out_926     ),
    .col_in_927              ( col_out_927     ),
    .col_in_928              ( col_out_928     ),
    .col_in_929              ( col_out_929     ),
    .col_in_930              ( col_out_930     ),
    .col_in_931              ( col_out_931     ),
    .col_in_932              ( col_out_932     ),
    .col_in_933              ( col_out_933     ),
    .col_in_934              ( col_out_934     ),
    .col_in_935              ( col_out_935     ),
    .col_in_936              ( col_out_936     ),
    .col_in_937              ( col_out_937     ),
    .col_in_938              ( col_out_938     ),
    .col_in_939              ( col_out_939     ),
    .col_in_940              ( col_out_940     ),
    .col_in_941              ( col_out_941     ),
    .col_in_942              ( col_out_942     ),
    .col_in_943              ( col_out_943     ),
    .col_in_944              ( col_out_944     ),
    .col_in_945              ( col_out_945     ),
    .col_in_946              ( col_out_946     ),
    .col_in_947              ( col_out_947     ),
    .col_in_948              ( col_out_948     ),
    .col_in_949              ( col_out_949     ),
    .col_in_950              ( col_out_950     ),
    .col_in_951              ( col_out_951     ),
    .col_in_952              ( col_out_952     ),
    .col_in_953              ( col_out_953     ),
    .col_in_954              ( col_out_954     ),
    .col_in_955              ( col_out_955     ),
    .col_in_956              ( col_out_956     ),
    .col_in_957              ( col_out_957     ),
    .col_in_958              ( col_out_958     ),
    .col_in_959              ( col_out_959     ),
    .col_in_960              ( col_out_960     ),
    .col_in_961              ( col_out_961     ),
    .col_in_962              ( col_out_962     ),
    .col_in_963              ( col_out_963     ),
    .col_in_964              ( col_out_964     ),
    .col_in_965              ( col_out_965     ),
    .col_in_966              ( col_out_966     ),
    .col_in_967              ( col_out_967     ),
    .col_in_968              ( col_out_968     ),
    .col_in_969              ( col_out_969     ),
    .col_in_970              ( col_out_970     ),
    .col_in_971              ( col_out_971     ),
    .col_in_972              ( col_out_972     ),
    .col_in_973              ( col_out_973     ),
    .col_in_974              ( col_out_974     ),
    .col_in_975              ( col_out_975     ),
    .col_in_976              ( col_out_976     ),
    .col_in_977              ( col_out_977     ),
    .col_in_978              ( col_out_978     ),
    .col_in_979              ( col_out_979     ),
    .col_in_980              ( col_out_980     ),
    .col_in_981              ( col_out_981     ),
    .col_in_982              ( col_out_982     ),
    .col_in_983              ( col_out_983     ),
    .col_in_984              ( col_out_984     ),
    .col_in_985              ( col_out_985     ),
    .col_in_986              ( col_out_986     ),
    .col_in_987              ( col_out_987     ),
    .col_in_988              ( col_out_988     ),
    .col_in_989              ( col_out_989     ),
    .col_in_990              ( col_out_990     ),
    .col_in_991              ( col_out_991     ),
    .col_in_992              ( col_out_992     ),
    .col_in_993              ( col_out_993     ),
    .col_in_994              ( col_out_994     ),
    .col_in_995              ( col_out_995     ),
    .col_in_996              ( col_out_996     ),
    .col_in_997              ( col_out_997     ),
    .col_in_998              ( col_out_998     ),
    .col_in_999              ( col_out_999     ),
    .col_in_1000             ( col_out_1000    ),
    .col_in_1001             ( col_out_1001    ),
    .col_in_1002             ( col_out_1002    ),
    .col_in_1003             ( col_out_1003    ),
    .col_in_1004             ( col_out_1004    ),
    .col_in_1005             ( col_out_1005    ),
    .col_in_1006             ( col_out_1006    ),
    .col_in_1007             ( col_out_1007    ),
    .col_in_1008             ( col_out_1008    ),
    .col_in_1009             ( col_out_1009    ),
    .col_in_1010             ( col_out_1010    ),
    .col_in_1011             ( col_out_1011    ),
    .col_in_1012             ( col_out_1012    ),
    .col_in_1013             ( col_out_1013    ),
    .col_in_1014             ( col_out_1014    ),
    .col_in_1015             ( col_out_1015    ),
    .col_in_1016             ( col_out_1016    ),
    .col_in_1017             ( col_out_1017    ),
    .col_in_1018             ( col_out_1018    ),
    .col_in_1019             ( col_out_1019    ),
    .col_in_1020             ( col_out_1020    ),
    .col_in_1021             ( col_out_1021    ),
    .col_in_1022             ( col_out_1022    ),
    .col_in_1023             ( col_out_1023    ),

    .compressor_array_512_out0 ( compressor_array_512_out0   ),
    .compressor_array_512_out1 ( compressor_array_512_out1   ),
    .data_out_0              ( data_out_0     ),
    .data_out_1              ( data_out_1     )
);


reg [5:0] state_current;
reg [5:0] state_next;


always@(posedge clk) begin
    if(rst) begin 
        state_current <= IDLE;
    end
    else begin
        state_current <= state_next;
    end
end

always@(posedge clk) begin
    if(rst) begin 
        counter <= 31'b0;
    end
    else begin
        if(finish_ms) counter <= counter + 1'b1;
        else counter <= counter;

    end
end


always@(*)begin
    case(state_current)
    IDLE: 
        begin
            if(reg_start_ms)
                state_next <= TRANS_DATA;
            else
                state_next <= IDLE;
        end

    TRANS_DATA: 
        begin
            state_next <= COMPRESS_HIGH;
        end

    COMPRESS_HIGH:
        begin 
            state_next <= COMPRESS_LOW;
        end

    COMPRESS_LOW: 
        begin
            state_next <= REDUCTION;
        end

    REDUCTION: 
        begin
            state_next <= FINISH;
        end

    FINISH: 
        begin
            if(counter < LOOPS)
                state_next <= COMPRESS_HIGH;
            else
                state_next <= IDLE;
        end

    default: 
        begin
            state_next <= IDLE;
        end
    endcase
end




always@(posedge clk)begin
    case(state_next)
    IDLE: 
        begin
            reg_start_ms                <= start_ms;
            reg_a                       <= 1024'b0;
            reg_partial_product_high0   <= 1024'b0;
            reg_partial_product_high1   <= 1024'b0;
            reg_partial_product_low0    <= 1033'b0;
            reg_partial_product_low1    <= 1033'b0;
            reg_sel_hp                  <= 1'b0;
            reg_sel_data_in             <= 1'b0;
            reg_data_out0               <= 1025'b0;
            reg_data_out1               <= 1025'b0;
            reg_finish_ms               <= 1'b0;
        end

    TRANS_DATA: 
        begin
            reg_start_ms                <= start_ms;
            reg_a                       <= a;
            reg_partial_product_high0   <= reg_partial_product_high0;
            reg_partial_product_high1   <= reg_partial_product_high1;
            reg_partial_product_low0    <= reg_partial_product_low0;
            reg_partial_product_low1    <= reg_partial_product_low1;
            reg_sel_hp                  <= 1'b1;
            reg_sel_data_in             <= 1'b1;
            reg_data_out0               <= data_out_0;
            reg_data_out1               <= data_out_1;
            reg_finish_ms               <= 1'b0;
        end

    COMPRESS_HIGH: 
        begin
            reg_start_ms                <= start_ms;
            reg_a                       <= reg_a;
            reg_partial_product_high0   <= compressor_array_512_out0[1023:0];
            reg_partial_product_high1   <= compressor_array_512_out1[1023:0];
            reg_partial_product_low0    <= reg_partial_product_low0;
            reg_partial_product_low1    <= reg_partial_product_low1;
            reg_sel_hp                  <= 1'b0;
            reg_sel_data_in             <= 1'b1;
            reg_data_out0               <= reg_data_out0;
            reg_data_out1               <= reg_data_out1;
            reg_finish_ms               <= 1'b0;
        end


    COMPRESS_LOW: 
        begin
            reg_start_ms                <= start_ms;
            reg_a                       <= reg_a;
            reg_partial_product_high0   <= reg_partial_product_high0;
            reg_partial_product_high1   <= reg_partial_product_high1;
            reg_partial_product_low0    <= compressor_array_512_out0;
            reg_partial_product_low1    <= compressor_array_512_out1;
            reg_sel_hp                  <= 1'b1;
            reg_sel_data_in             <= 1'b0;
            reg_data_out0               <= reg_data_out0;
            reg_data_out1               <= reg_data_out1;
            reg_finish_ms               <= 1'b0;
        end

    REDUCTION: 
        begin
            reg_start_ms                <= start_ms;
            reg_a                       <= reg_a;
            reg_partial_product_high0   <= reg_partial_product_high0;
            reg_partial_product_high1   <= reg_partial_product_high1;
            reg_partial_product_low0    <= reg_partial_product_low0;
            reg_partial_product_low1    <= reg_partial_product_low1;
            reg_sel_hp                  <= 1'b1;
            reg_sel_data_in             <= 1'b0;
            reg_data_out0               <= data_out_0;
            reg_data_out1               <= data_out_1;
            reg_finish_ms               <= 1'b0;
        end
    
    FINISH: 
        begin
            reg_start_ms                <= start_ms;
            reg_a                       <= ms;
            reg_partial_product_high0   <= reg_partial_product_high0;
            reg_partial_product_high1   <= reg_partial_product_high1;
            reg_partial_product_low0    <= reg_partial_product_low0;
            reg_partial_product_low1    <= reg_partial_product_low1;
            reg_sel_hp                  <= 1'b1;
            reg_sel_data_in             <= 1'b1;
            reg_data_out0               <= reg_data_out0;
            reg_data_out1               <= reg_data_out1;
            reg_finish_ms               <= 1'b1;
        end

    default: 
        begin
            reg_start_ms                <= start_ms;
            reg_a                       <= 1024'b0;
            reg_partial_product_high0   <= 1024'b0;
            reg_partial_product_high1   <= 1024'b0;
            reg_partial_product_low0    <= 1033'b0;
            reg_partial_product_low1    <= 1033'b0;
            reg_sel_hp                  <= 1'b1;
            reg_sel_data_in             <= 1'b1;
            reg_data_out0               <= 1025'b0;
            reg_data_out1               <= 1025'b0;
            reg_finish_ms               <= 1'b0;
        end
    endcase
end




assign finish_ms = reg_finish_ms;

assign temp_ms0 = reg_data_out0 + reg_data_out1;
assign temp_ms1 = reg_data_out0 + reg_data_out1 - P1;
assign temp_ms2 = reg_data_out0 + reg_data_out1 - P2;
assign temp_ms3 = reg_data_out0 + reg_data_out1 - P3;


always@(*)begin
    if(!temp_ms3[1026]) temp_ms = temp_ms3[1023:0];
    else if(!temp_ms2[1026]) temp_ms = temp_ms2[1023:0];
    else if(!temp_ms1[1026]) temp_ms = temp_ms1[1023:0];
    else temp_ms = temp_ms0[1023:0];
end

assign ms = temp_ms;



endmodule
module xpb_5_695
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h7b0ec66fec2a1f679d76b3b5bcaadd0ac423ba7912b9be0463ce511a797938a87f8233232388586e7d4665cef26d395ce9a60a446a3b9abc0c9466bead3bdbe805dae0ab1319ec063d2393e5ac140f0138966640e5ebbd62b0c585f5e0c7581a41d040de8f4b181e50dae94f1bdb23204c77c31b4316d7cc1c53a72ce664f99e;
    5'b00010 : xpb = 1024'h4570478a16660a066fe7ef9468fb72c416d171c14ffbdb9149bfe8df3fefc448fbbbe8cd7cea324e5b2e8c57017c61ef6f31eca2b1c4652c68898e1f1fa5431e97668ca776a2dac767ad2528bf4c59d17d27d2e93f514db4abfe79f107640da25498ef936dcd37af1af5ebbf3fe620174a15a75435e25267f237d35543e78cd1;
    5'b00011 : xpb = 1024'hfd1c8a440a1f4a542592b73154c087d697f29098d3df91e2fb180a406664fe977f59e77d64c0c2e3916b2df108b8a81f4bdcf00f94d2f9cc47eb57f920eaa5528f238a3da2bc9889236b66bd284a4a1c1b93f9198b6de06a7376dec2e00c32a67619e484c4f573fe510ee2f63f11d0e47b38b8d28adcd03c81bff7da16a2004;
    5'b00100 : xpb = 1024'h8ae08f142ccc140cdfcfdf28d1f6e5882da2e3829ff7b722937fd1be7fdf8891f777d19af9d4649cb65d18ae02f8c3dede63d9456388ca58d1131c3e3f4a863d2ecd194eed45b58ecf5a4a517e98b3a2fa4fa5d27ea29b6957fcf3e20ec81b44a931df26db9a6f5e35ebd77e7fcc402e942b4ea86bc4a4cfe46fa6aa87cf19a2;
    5'b00101 : xpb = 1024'h5542102e5707feabb2411b077e477b4180509acadd39d4af797169834656143273b1874553363e7c94453f361207ec7163efbba3ab1194c92d08439eb1b3ed73c058c54b50cea44ff9e3db9491d0fe733ee1127ad8082bbb5335e7dd3564d0ccbbfa8ddbba1c8eef0006d9eea3d73d2591c932e15e901f6bba53d2d2e551acd5;
    5'b00110 : xpb = 1024'h1fa391488143e94a84b256e62a9810fad2fe52131a7bf23c5f6301480ccc9fd2efeb3cefac98185c722d65be21171503e97b9e01f29a5f3988fd6aff241d54aa51e47147b4579311246d6cd7a509494383727f23316dbc0d4e6edbd85c018654cec33c90989eae7fca21dc5ec7e23a1c8f67171a515b9a079037fefb42d44008;
    5'b00111 : xpb = 1024'h9ab257b86d6e08b222290a9be742ee0597220c8c2d35b040c33152628645d87b6f6d7012d02070caef73cb8d13844e60d321a8465cd5f9f59591d1bdd159309257bf51f2c7717f17619100bd511d5844bc08e5641759796fff3461ce3cc8de6f10937d6f27e9c69e1afcc5ade3bd5d3cdbdeda35947271d3ac8ba628293939a6;
    5'b01000 : xpb = 1024'h6513d8d297a9f350f49a467a939383bee9cfc3d46a77cdcda922ea274cbc641beba725bd29824aaacd5bf215229376f358ad8aa4a45ec465f186f91e43c297c8e94afdef2afa6dd88c1a92006455a315009a520c70bf09c1fa6d55c9636593f7235c2c24066be62ee517c81e07c85a33d97cbe6e873dec6f826fd25086bbccd9;
    5'b01001 : xpb = 1024'h2f7559ecc1e5ddefc70b82593fe419783c7d7b1ca7b9eb5a8f1481ec1332efbc67e0db6782e4248aab44189d31a29f85de396d02ebe78ed64d7c207eb62bfeff7ad6a9eb8e835c99b6a42343778dede5452bbeb4ca249a13f5a649c48a02497f3624dad8e4ee05bfaf32ca8e2bd3572ad71aa2a77a09670b5853fe78e43e600c;
    5'b01010 : xpb = 1024'haa84205cae0ffd576482360efc8ef68300a13595ba73a95ef2e2d3068cac2864e7630e8aa66c7cf9288a7e6c240fd8e2c7df7747562329925a10873d6367dae780b18a96a19d489ff3c7b72923a1fce67dc224f5b0105776a66bcfba6ac9a19977f51bb774391dde000db3dd47ae7a4b239265c2bd203ed774a7a5a5caa359aa;
    5'b01011 : xpb = 1024'h74e5a176d84be7f636f371eda8df8c3c534eecddf7b5c6ebd8d46acb5322b405639cc434ffce56d90672a4f4331f01754d6b59a59dabf402b605ae9dd5d1421e123d3693052637611e51486c36da47b6c253919e0975e7c8a1a4c3b5916657218abdca6c52bb3d6eca28b64d6bb97742213049fbafebb9734a8bd1ce2825ecdd;
    5'b01100 : xpb = 1024'h3f4722910287d2950964adcc553021f5a5fca42634f7e478bec6029019993fa5dfd679df593030b8e45acb7c422e2a07d2f73c03e534be7311fad5fe483aa954a3c8e28f68af262248dad9af4a12928706e4fe4662db781a9cddb7b0b8030ca99d867921313d5cff9443b8bd8fc474391ece2e34a2b7340f206ffdf685a88010;
    5'b01101 : xpb = 1024'h9a8a3ab2cc3bd33dbd5e9ab0180b7aef8aa5b6e723a0205a4b79a54e00fcb465c102f89b2920a98c242f204513d529a58831e622cbd88e36deffd5ebaa4108b35548e8bcc3814e373646af25d4add574b766aeebc41086c9816ababde9fc231b04f27d60fbf7c905e5ebb2db3cf71301c6c126d9582aeaaf6542a1ee32b1343;
    5'b01110 : xpb = 1024'h84b76a1b18eddc9b794c9d60be2b94b9bcce15e784f3c00a0885eb6f598903eedb9262acd61a63073f8957d343aa8bf7422928a696f9239f7a84641d67dfec733b2f6f36df5200e9b087fed8095eec58840cd12fa22cc5cf48dc31a1bf671a4bf21f68b49f0a94aeaf39a47ccfaa945068e3d588d899867712a7d14bc9900ce1;
    5'b01111 : xpb = 1024'h4f18eb354329c73a4bbdd93f6a7c2a730f7bcd2fc235dd96ee7783341fff8f8f57cc18572f7c3ce71d717e5b52b9b489c7b50b04de81ee0fd6798b7dda4953a9ccbb1b3342daefaadb11901b1c973728c89e3dd7fb9256214415259ce603cfd404e817697d8cb43f7954a6ecf3b591476681b9c1cb650112e88bfd742712a014;
    5'b10000 : xpb = 1024'h197a6c4f6d65b1d91e2f151e16ccc02c62298477ff77fb23d4691af8e6761b2fd405ce0188de16c6fb59a4e361c8dd1c4d40ed63260ab880326eb2de4cb2bae05e46c72fa663de6c059b215e2fcf81f90d2faa8054f7e6733f4e19980ca0855c17b0c61e5c0ed3d0436fa95d17c08e3e641f9dfabe307baebe70299c84953347;
    5'b10001 : xpb = 1024'h948932bf598fd140bba5c8d3d3779d37264d3ef11231b92838376c135fef53d853880124ac666f3578a00ab25436167936e6f7a79046533c3f03199cf9ee96c86421a7dab97dca7242beb543dbe390fa45c610c13ae3a3d5f0139f8ded67dd76598106fceb59ebee944a92ac339bb15eb09761160147537adac3d0c96afa2ce5;
    5'b10010 : xpb = 1024'h5eeab3d983cbbbdf8e1704b27fc832f078faf6394f73d6b51e2903d82665df78cfc1b6cf05c849155688313a63453f0bbc72da05d7cf1dac9af840fd6c57fdfef5ad53d71d06b9336d484686ef1bdbca8a577d6994493427eb4c9389140492fe6c49b5b1c9dc0b7f5e65951c57a6ae55ae35454ef412ce16b0a7fcf1c87cc018;
    5'b10011 : xpb = 1024'h294c34f3ae07a67e608840912c18c8a9cba8ad818cb5f442041a9b9cecdc6b194bfb6c795f2a22f5347057c27254679e41febc641f57e81cf6ed685ddec165358738ffd3808fa7f497d1d7ca0254269acee8ea11edaec479e68587843aa148867f126466a85e2b102880978c7bb1ab4cabd32987e6de48b2868c291a25ff534b;
    5'b10100 : xpb = 1024'ha45afb639a31c5e5fdfef446e8c3a5b48fcc67fa9f6fb24667e8ecb76655a3c1cb7d9f9c82b27b63b1b6bd9164c1a0fb2ba4c6a8899382d90381cf1c8bfd411d8d13e07e93a993fad4f56bafae68359c077f5052d39a81dc974b0d7a1b68a0a0c0e2a54537a9432e795b80db978cce6cf84aeca329f5207ea2dfd0470c644ce9;
    5'b10101 : xpb = 1024'h6ebc7c7dc46db084d070302595143b6de27a1f42dcb1cfd34dda847c2ccc2f6247b75546dc1455438f9ee41973d0c98db130a906d11c4d495f76f67cfe66a8541e9f8c7af73282bbff7efcf2c1a0806c4c10bcfb2d00122e9284017542055628d3ab53fa162b62bf4376834bbb97cb63f5e8d0dc1cc09b1a78c3fc6f69e6e01c;
    5'b10110 : xpb = 1024'h391dfd97eea99b23a2e16c044164d1273527d68b19f3ed6033cc1c40f342bb02c3f10af135762f236d870aa182dff22036bc8b6518a517b9bb6c1ddd70d00f8ab02b38775abb717d2a088e35d4d8cb3c90a229a38665a2808dbcf57068a20bb0e67402aef4ad82500d9185bbdfa2c85af386b5150f8c15b64ea82897c769734f;
    5'b10111 : xpb = 1024'h37f7eb218e585c27552a7e2edb566e087d58dd357360aed19bdb405b9b946a3402ac09b8ed809034b6f312991ef1ab2bc486dc3602de22a1761453de33976c141b6e473be44603e54921f78e811160cd533964bdfcb32d288f5e96b8f3ec138f93cb163d32fa1e0d7ac882c03adc551f124994e02579052248c54c024ec0682;
    5'b11000 : xpb = 1024'h7e8e4522050fa52a12c95b98aa6043eb4bf9484c69efc8f17d8c052033327f4bbfacf3beb2606171c8b596f8845c540fa5ee7807ca697ce623f5abfc907552a94791c51ed15e4c4491b5b35e9425250e0dc9fc8cc5b6f03539bb6f61700619533b0cf242627ab9ff2887717b1f88e8723d9c5c69456e681e40dffbed0b510020;
    5'b11001 : xpb = 1024'h48efc63c2f4b8fc8e53a977756b0d9a49ea6ff94a731e67e637d9ce4f9a90aec3be6a9690bc23b51a69dbd80936b7ca22b7a5a6611f247567fead35d02deb9dfd91d711b34e73b05bc3f44a1a75d6fde525b69351f1c808734f4635c96a2cedb4dd5a0f740fcd98ff2a273eb4393e5693b3a40a23839e2ba16c4281568d39353;
    5'b11010 : xpb = 1024'h1351475659877a67b7abd35603016f5df154b6dce474040b496f34a9c01f968cb8205f13652415318485e408a27aa534b1063cc4597b11c6dbdffabd754821166aa91d17987029c6e6c8d5e4ba95baae96ecd5dd788210d9302d5757bd3f8463609e4fac1f7ef920bcbd765b679ee26038d824db2b055d55eca8543dc6562686;
    5'b11011 : xpb = 1024'h8e600dc645b199cf5522870bbfac4c68b5787155f72dc20fad3d85c43998cf3537a2923688ac6da001cc49d794e7de919aac4708c3b6ac82e874617c2283fcfe7083fdc2ab8a15cd23ec69ca66a9c9afcf833c1e5e6dce3be0f2dd4d9e06dc7da26e908aaeca113f0d985faa837a0580854fe7f66e1c352208fbfb6aacbb2024;
    5'b11100 : xpb = 1024'h58c18ee06fed846e2793c2ea6bfce2220826289e346fdf9c932f1d89000f5ad5b3dc47e0e20e477fdfb4705fa3f70724203829670b3f76f3446988dc94ed6435020fa9bf0f13048e4e75fb0d79e214801414a8c6b7d35e8ddc2bd148c4a39205b5373f3f8d4c30cfd7b3621aa785027782edcc2f60e7afbddee027930a3db357;
    5'b11101 : xpb = 1024'h23230ffa9a296f0cfa04fec9184d77db5ad3dfe671b1fd297920b54dc685e6763015fd8b3b70215fbd9c96e7b3062fb6a5c40bc552c84163a05eb03d0756cb6b939b55bb729bf34f78ff8c508d1a5f5058a6156f1138eedfd764c543eb40478dc7ffedf46bce5060a1ce648acb8fff6e808bb06853b32a59b4c453bb67c0468a;
    5'b11110 : xpb = 1024'h9e31d66a86538e74977bb27ed4f854e61ef79a5f846bbb2ddcef06683fff1f1eaf9830ae5ef879ce3ae2fcb6a57369138f6a1609bd03dc1facf316fbb492a7539976366685b5df55b6232036392e6e51913c7baff724ac42882a4b39cc079fa809d02ed2fb19687ef2a94dd9e76b228ecd03738396ca0225d117fae84e254028;
    5'b11111 : xpb = 1024'h68935784b08f791369ecee5d8148ea9f71a551a7c1add8bac2e09e2d0675aabf2bd1e658b85a53ae18cb233eb48291a614f5f868048ca69008e83e5c26fc0e8a2b01e262e93ece16e0acb1794c66b921d5cde858508a3c9483633f34f2a455301c98dd87d99b880fbcc4504a0b761f85caa157bc89957cc1a6fc2710aba7d35b;
    endcase
end

endmodule

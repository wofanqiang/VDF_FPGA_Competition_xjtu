module xpb_5_430
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h4b02701ce7c564b930e1e987d6ed5c48e342c12ef16ca65172a7b4cc3bba46124570b5d23d0a54af07fcb00e3b782cc688018164b6712725dfce9d0bfeb766482d68259deac58c374f2b03daebf03bd1ea98104736fcb9f0454631a0a29535704a5ee8823cb9252f93b1921ff22618c63820cdbe2fed3d686df692e3172b06a;
    5'b00010 : xpb = 1024'h9604e039cf8ac97261c3d30faddab891c685825de2d94ca2e54f699877748c248ae16ba47a14a95e0ff9601c76f0598d100302c96ce24e4bbf9d3a17fd6ecc905ad04b3bd58b186e9e5607b5d7e077a3d530208e6df973e08a8c6341452a6ae094bdd10479724a5f2763243fe44c318c70419b7c5fda7ad0dbed25c62e560d4;
    5'b00011 : xpb = 1024'he1075056b7502e2b92a5bc9784c814daa9c8438cd445f2f457f71e64b32ed236d0522176b71efe0d17f6102ab26886539804842e235375719f6bd723fc2632d8883870d9c050a4a5ed810b90c3d0b375bfc830d5a4f62dd0cfd294e1e7bfa050df1cb986b62b6f8ebb14b65fd6724a52a862693a8fc7b83949e3b8a9458113e;
    5'b00100 : xpb = 1024'h12c09c0739f1592e4c387a61f5bb571238d0b04bbc5b29945ca9ed330eee9184915c2d748f42952bc1ff2c038ede0b31a20060592d9c49c977f3a742ffadd9920b5a09677ab1630dd3cac0f6bafc0ef47aa60411cdbf2e7c11518c6828a54d5c1297ba208f2e494be4ec6487fc8986318e08336f8bfb4f5a1b7da4b8c5cac1a8;
    5'b00101 : xpb = 1024'h1770c309086daf79df4698fa732a2cd6c704dc5eab71f3f973d4687fd2aa35e5b5b338d1b3133a76b27ef70472958dfe0a80786f79035c3bd5f09113bf994ff68e308bc1595dbbd148bd713469bb12b1994f8516412efa1b15a5ef8232cea0b3173da8a8b2f9db9ede277da9fbabe7bdf18a404b6efa2330a25d0de6f73d7212;
    5'b00110 : xpb = 1024'h1c20ea0ad6ea05c57254b792f099029b553908719a88be5e8afee3cc9665da46da0a442ed6e3dfc1a2fec205564d10ca73009085c46a6eae33ed7ae47f84c65b11070e1b380a1494bdb02172187a166eb7f9061ab49ec5ba19fa529c3cf7f40a1be39730d6c56df1d76296cbface494a550c4d2751f8f707293c771528b0227c;
    5'b00111 : xpb = 1024'h20d1110ca5665c110562d62b6e07d85fe36d3484899f88c3a2295f195a217ea7fe614f8bfab4850c937e8d063a049396db80a89c0fd1812091ea64b53f703cbf93dd907516b66d5832a2d1afc7391a2bd6a2871f280e91591e4eb5b647214761208985b8fa910044d09dafedf9f0aad6b88e5a0334f7caddb01be0435a22d2e6;
    5'b01000 : xpb = 1024'h2581380e73e2b25c9870f4c3eb76ae2471a1609778b65328b953da661ddd230922b85ae91e852a5783fe58071dbc16634400c0b25b389392efe74e85ff5bb32416b412cef562c61ba79581ed75f81de8f54c08239b7e5cf822a318d0514a9ab8252f74411e5c9297c9d8c90ff9130c631c1066df17f69eb436fb49718b958350;
    5'b01001 : xpb = 1024'h2a315f10425f08a82b7f135c68e583e8ffd58caa67cd1d8dd07e55b2e198c76a470f66464255cfa2747e23080173992fac80d8c8a69fa6054de43856bf472988998a9528d40f1edf1c88322b24b721a613f589280eee289726f77bea5b73ee0f29d562c9422824eac313e231f8356def7f9273bafaf5728abddab29fbd0833ba;
    5'b01010 : xpb = 1024'h2ee1861210db5ef3be8d31f4e65459ad8e09b8bd56e3e7f2e7a8d0ffa5546bcb6b6671a3662674ed64fdee08e52b1bfc1500f0def206b877abe122277f329fed1c611782b2bb77a2917ae268d3762563329f0a2c825df4362b4bdf04659d41662e7b515165f3b73dbc4efb53f757cf7be3148096ddf4466144ba1bcdee7ae424;
    5'b01011 : xpb = 1024'h3391ad13df57b53f519b508d63c32f721c3de4d045fab257fed34c4c6910102c8fbd7d0089f71a38557db909c8e29ec87d8108f53d6dcaea09de0bf83f1e16519f3799dc9167d066066d92a68235292051488b30f5cdbfd52fa0421e6fc694bd33213fd989bf4990b58a1475f67a310846968d72c0f31a37cb9984fc1fed948e;
    5'b01100 : xpb = 1024'h3841d415add40b8ae4a96f25e1320536aa7210e335117cbd15fdc7992ccbb48db414885dadc7bf8345fd840aac9a2194e601210b88d4dd5c67daf5c8ff098cb6220e1c36701429297b6042e430f42cdd6ff20c35693d8b7433f4a53879efe81437c72e61ad8adbe3aec52d97f59c9294aa189a4ea3f1ee0e5278ee2a516044f8;
    5'b01101 : xpb = 1024'h3cf1fb177c5061d677b78dbe5ea0dafb38a63cf6242847222d2842e5f08758eed86b93bad19864ce367d4f0b9051a4614e813921d43befcec5d7df99bef5031aa4e49e904ec081ecf052f321dfb3309a8e9b8d39dcad57133849085284193b6b3c6d1ce9d1566e36a80046b9f4bef4210d9aa72a86f0c1e4d958575882d2f562;
    5'b01110 : xpb = 1024'h41a222194accb8220ac5ac56dc0fb0bfc6da6909133f11874452be32b442fd4ffcc29f17f5690a1926fd1a0c7409272db70151381fa3024123d4c96a7ee0797f27bb20ea2d6cdab06545a35f8e723457ad450e3e501d22b23c9d6b6c8e428ec241130b71f5220089a13b5fdbf3e155ad711cb40669ef95bb6037c086b445a5cc;
    5'b01111 : xpb = 1024'h4652491b19490e6d9dd3caef597e8684550e951c0255dbec5b7d397f77fea1b12119aa751939af64177ce50d57c0a9fa1f81694e6b0a14b381d1b33b3ecbefe3aa91a3440c193373da38539d3d313814cbee8f42c38cee5140f1ce86986be21945b8f9fa18ed92dc9a7678fdf303b739d49ec0e24cee6991e71729b4e5b85636;
    5'b10000 : xpb = 1024'h4b02701ce7c564b930e1e987d6ed5c48e342c12ef16ca65172a7b4cc3bba46124570b5d23d0a54af07fcb00e3b782cc688018164b6712725dfce9d0bfeb766482d68259deac58c374f2b03daebf03bd1ea98104736fcb9f0454631a0a29535704a5ee8823cb9252f93b1921ff22618c63820cdbe2fed3d686df692e3172b06a0;
    5'b10001 : xpb = 1024'h4fb2971eb641bb04c3f00820545c320d7176ed41e08370b689d23018ff75ea7369c7c12f60daf9f9f87c7b0f1f2faf92f081997b01d839983dcb86dcbea2dcacb03ea7f7c971e4fac41db4189aaf3f8f0941914baa6c858f499a94baacbe88c74f04d70a6084b7828cecab41f1487a529ba2da9a12ec113ef4d5fc11489db70a;
    5'b10010 : xpb = 1024'h5462be2084be115056fe26b8d1cb07d1ffab1954cf9a3b1ba0fcab65c3318ed48e1ecc8c84ab9f44e8fc461002e7325f5901b1914d3f4c0a9bc870ad7e8e531133152a51a81e3dbe39106456496e434c27eb12501ddc512e4deef7d4b6e7dc1e53aac592845049d58627c463f06adbdeff24e775f5eae5157bb5653f7a106774;
    5'b10011 : xpb = 1024'h5912e522533a679bea0c45514f39dd968ddf4567beb10580b82726b286ed3335b275d7e9a87c448fd97c1110e69eb52bc181c9a798a65e7cf9c55a7e3e79c975b5ebacab86ca9681ae031493f82d470946949354914c1ccd52435aeec1112f755850b41aa81bdc287f62dd85ef8d3d6b62a6f451d8e9b8ec0294ce6dab8317de;
    5'b10100 : xpb = 1024'h5dc30c2421b6bde77d1a63e9cca8b35b1c13717aadc7cfe5cf51a1ff4aa8d796d6cce346cc4ce9dac9fbdc11ca5637f82a01e1bde40d70ef57c2444efe653fda38c22f056576ef4522f5c4d1a6ec4ac6653e145904bbe86c5697be08cb3a82cc5cf6a2a2cbe76e7b789df6a7eeaf9ef7c629012dbbe88cc28974379bdcf5c848;
    5'b10101 : xpb = 1024'h62733325f0331433102882824a17891faa479d8d9cde9a4ae67c1d4c0e647bf7fb23eea3f01d8f25ba7ba712ae0dbac49281f9d42f748361b5bf2e1fbe50b63ebb98b15f4423480897e8750f55ab4e8383e7955d782bb40b5aec2122d563d623619c912aefb300ce71d90fc9edd2008429ab0e099ee760991053a0ca0e6878b2;
    5'b10110 : xpb = 1024'h67235a27beaf6a7ea336a11ac7865ee4387bc9a08bf564affda69898d22020591f7afa0113ee3470aafb721391c53d90fb0211ea7adb95d413bc17f07e3c2ca33e6f33b922cfa0cc0cdb254d046a5240a2911661eb9b7faa5f40843cdf8d297a66427fb3137e93216b1428ebecf462108d2d1ae581e6346f973309f83fdb291c;
    5'b10111 : xpb = 1024'h6bd381298d2bc0ca3644bfb344f534a8c6aff5b37b0c2f1514d113e595dbc4ba43d2055e37bed9bb9b7b3d14757cc05d63822a00c642a84671b901c13e27a307c145b613017bf98f81cdd58ab32955fdc13a97665f0b4b496394e756e9b67cd16ae86e3b374a2574644f420dec16c39cf0af27c164e508461e127326714dd986;
    5'b11000 : xpb = 1024'h7083a82b5ba81715c952de4bc2640a6d54e421c66a22f97a2bfb8f325997691b682910bb5b8f7f068bfb081559344329cc02421711a9bab8cfb5eb91fe13196c441c386ce0285252f6c085c861e859badfe4186ad27b16e867e94a70f3dfd0286f8e5cc35b15b7c75d8a5b2feb3925295431349d47e3dc1ca4f1dc54a2c089f0;
    5'b11001 : xpb = 1024'h7533cf2d2a246d615c60fce43fd2e031e3184dd95939c3df43260a7f1d530d7c8c801c187f6024517c7ad3163cebc5f634825a2d5d10cd2b2db2d562bdfe8fd0c6f2bac6bed4ab166bb3360610a75d77fe8d996f45eae2876c3dad8afe09237f74344b4b7ee14a1a56c57451ea5b86b5b7b341792ae2aff32bd14582d4333a5a;
    5'b11010 : xpb = 1024'h79e3f62ef8a0c3acef6f1b7cbd41b5f6714c79ec48508e445a5085cbe10eb1ddb0d72775a330c99c6cfa9e1720a348c29d027243a877df9d8bafbf337dea063549c93d209d8103d9e0a5e643bf6661351d371a73b95aae26709210a5083276d678da39d3a2acdc6d50008d73e97de8421b354e550de183c9b2b0aeb105a5eac4;
    5'b11011 : xpb = 1024'h7e941d30c71d19f8827d3a153ab08bbaff80a5ff376758a9717b0118a4ca563ed52e32d2c7016ee75d7a6918045acb8f05828a59f3def20fe9aca9043dd57c99cc9fbf7a7c2d5c9d559896816e2564f23be09b782cca79c574e673bf125bca2d7d80285bc6786ec0493ba695e8a049ce7eb75b30f0e057a0399017df37189b2e;
    5'b11100 : xpb = 1024'h8344443295997044158b58adb81f617f8db4d212267e230e88a57c656885fa9ff9853e2fead214324dfa3418e8124e5b6e02a2703f46048247a992d4fdc0f2fe4f7641d45ad9b560ca8b46bf1ce468af5a8a1c7ca03a4564793ad6d91c851d84822616e3ea4401134276bfb7e7c2ab5ae239680cd3df2b76c06f810d688b4b98;
    5'b11101 : xpb = 1024'h87f46b346415c68fa8997746358e37441be8fe251594ed739fcff7b22c419f011ddc498d0ea2b97d3e79ff19cbc9d127d682ba868aad16f4a5a67ca5bdac6962d24cc42e39860e243f7df6fccba36c6c79339d8113aa11037d8f39f326ae70db86cc056c0e0f93663bb1d8d9e6e50ce745bb74e8b6ddff4d474eea3b99fdfc02;
    5'b11110 : xpb = 1024'h8ca4923632921cdb3ba795deb2fd0d08aa1d2a3804abb7d8b6fa72feeffd4362423354ea32735ec82ef9ca1aaf8153f43f02d29cd614296703a366767d97dfc755234688183266e7b470a73a7a62702997dd1e858719dca281e39d0d30d7c4328b71f3f431db25b934ecf1fbe6076e73a93d81c499dcd323ce2e5369cb70ac6c;
    5'b11111 : xpb = 1024'h9154b938010e7326ceb5b477306be2cd3851564af3c2823dce24ee4bb3b8e7c3668a6047564404131f79951b9338d6c0a782eab3217b3bd961a050473d83562bd7f9c8e1f6debfab29635778292173e6b6869f89fa89a841863800273b0117899017e27c55a6b80c2e280b1de529d0000cbf8ea07cdba6fa550dbc97fce35cd6;
    endcase
end

endmodule

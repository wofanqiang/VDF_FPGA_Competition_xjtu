module xpb_4_1020
(
    input [4:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    4'b0000 : xpb = 1024'h0;
    4'b0001 : xpb = 1024'h6e6828cdd3044576e56ee6e4f4f2f4a7996efc81e7fc27717975470a87a1b4552cf8249cfe1929200790b83228122ebb3b6690d1a75c6cb408fb5d7f391c8b7ad95c5942e5da5e413cbd2b6a6fb2d7dab03b235c64cafc42f85d9fe2db712cb987ca33db66bc49d1eea978fd270f277ec1fa124debe7ae6427db80efdda409ce;
    4'b0010 : xpb = 1024'h2c230c45e41a5624ffd855f2d98ba1fdc167f5d2fa80ae6b750dd4bf5c40bba256a7cbc1320bd3b16fc3311d6cc64cac12b2f9bd2c06091c61577ba03766a2443e697dd71c23bf3d66e054324689eb846c714d203d0fcb753b2eadcafcb7b6e0e08cd58d1caf9b1656930b1b564e28d4351a45b98783ff98094786db3265ad31;
    4'b0011 : xpb = 1024'h9a8b3513b71e9b9be5473cd7ce7e96a55ad6f254e27cd5dcee831bc9e3e26ff7839ff05e3024fcd17753e94f94d87b674e198a8ed36275d06a52d91f70832dbf17c5d71a01fe1d7ea39d7f9cb63cc35f1cac707ca1dac7b8338c4dadd828e39a68570968836be4e8453c84187d5d5052f7145807736badfc312307cb1009b6ff;
    4'b0100 : xpb = 1024'h5846188bc834ac49ffb0abe5b31743fb82cfeba5f5015cd6ea1ba97eb8817744ad4f97826417a762df86623ad98c99582565f37a580c1238c2aef7406ecd44887cd2fbae38477e7acdc0a8648d13d708d8e29a407a1f96ea765d5b95f96f6dc1c119ab1a395f362cad261636ac9c51a86a348b730f07ff30128f0db664cb5a62;
    4'b0101 : xpb = 1024'h1600fc03d94abcf81a1a1af397aff151aac8e4f70785e3d0e5b437338d207e91d6ff3ea6980a51f447b8db261e40b748fcb25c65dcb5aea11b0b15616d175b51e1e020426e90df76f7e3d12c63eaeab29518c4045264661cb92e697e1ab5f7e919dc4ccbef528771150fa854dbdb52fddd54bedeaaa45063f3fb13a1b98cfdc5;
    4'b0110 : xpb = 1024'h846924d1ac4f026eff8901d88ca2e5f94437e178ef820b425f297e3e14c232e703f7634396237b144f4993584652e6043818ed3784121b55240672e0a633e6ccbb3c7985546b3db834a0fc96d39dc28d4553e760b72f625fb18c0960f62724a2a1a680a7560ed14303b9215202ea7a7c9f4ed12c968bfec81bd6949197310793;
    4'b0111 : xpb = 1024'h42240849bd65131d19f270e6713b934f6c30daca0206923c5ac20bf2e9613a342da70a67ca1625a5b77c0c438b0703f50f65562308bbb7bd7c629101a47dfd9620499e198ab49eb45ec4255eaa74d637018a11248f743191f45d1749176daec9fa6922590c0222876ba2b37032297bd2126f049832284ffbfd429a7cebf2aaf6;
    4'b1000 : xpb = 1024'hb08c311790695893ff6157cb662e87f7059fd74bea02b9add43752fd7102ee895a9f2f04c82f4ec5bf0cc475b31932b04acbe6f4b0182471855dee80dd9a8910f9a5f75c708efcf59b8150c91a27ae11b1c53480f43f2dd4ecbab72bf2dedb838233563472be6c595a4c2c6d5938a350d46916e61e0ffe60251e1b6cc996b4c4;
    4'b1001 : xpb = 1024'h6e47148fa17f694219cac6d94ac7354d2d98d09cfc8740a7cfcfe0b245a1f5d6844ed628fc21f957273f3d60f7cd50a122184fe034c1c0d9ddba0ca1dbe49fda5eb31bf0a6d85df1c5a47990f0fec1bb6dfb5e44cc83fd072f8bc514142565aadaf5f7e628b1bd9dc235be8b8877a4a647894a51b9ac4f94068a21581e585827;
    4'b1010 : xpb = 1024'h2c01f807b29579f0343435e72f5fe2a35591c9ee0f0bc7a1cb686e671a40fd23adfe7d4d3014a3e88f71b64c3c816e91f964b8cbb96b5d4236162ac2da2eb6a3c3c04084dd21beedefc7a258c7d5d5652a318808a4c8cc39725cd2fc356befd233b89997dea50ee22a1f50a9b7b6a5fbbaa97dbd5548a0c7e7f627437319fb8a;
    4'b1011 : xpb = 1024'h9a6a20d58599bf6719a31ccc2452d74aef00c66ff707ef1344ddb571a1e2b178daf6a1ea2e2dcd0897026e7e64939d4d34cb499d60c7c9f63f118842134b421e9d1c99c7c2fc1d2f2c84cdc33788ad3fda6cab650993c87c6aba72df10dd1c8bbb82cd73456158b418c8c9a6dec5cd7a7ca3900b41304f2c0fd1a83350be0558;
    4'b1100 : xpb = 1024'h5825044d96afd015340c8bda08eb84a116f9bfc1098c760d407643267681b8c604a6490e62207799ff34e769a947bb3e0c17b288e571665e976da663119558e80229be5bf9457e2b56a7f68b0e5fc0e996a2d528e1d897aead8b80c73223a6b314456f24fb54a9f880b25bc50e04cecfefc3c376dccca05ff13dae1ea57fa8bb;
    4'b1101 : xpb = 1024'h15dfe7c5a7c5e0c34e75fae7ed8431f73ef2b9121c10fd073c0ed0db4b20c0132e55f0329613222b67676054edfbd92ee3641b746a1b02c6efc9c4840fdf6fb16736e2f02f8edf2780cb1f52e536d49352d8feecba1d66e0f05c8eaf536a30da6d0810d6b147fb3ce89bede33d43d02562e3f6e27868f193d2a9b409fa414c1e;
    4'b1110 : xpb = 1024'h844810937aca263a33e4e1cce277269ed861b594040d2478b58417e5d2c274685b4e14cf942c4b4b6ef81887160e07ea1ecaac4611776f7af8c5220348fbfb2c40933c3315693d68bd884abd54e9ac6e031422491ee86323e8ba2e922edb5d93f4d244b21804450ed74566e06452f7a424de093064509ff7fa8534f9d7e555ec;
    4'b1111 : xpb = 1024'h4202f40b8be036e84e4e50dac70fd3f5005aaee51691ab72b11ca59aa7617bb584fdbbf3c81ef5dcd72a91725ac225daf617153196210be351214024474611f5a5a060c74bb29e64e7ab73852bc0c017bf4a4c0cf72d32562b8b3c7a5021e7bb4d94e663cdf796533f2ef8fe9391f8f997fe3c9bffecf12bdbf13ae52ca6f94f;
    endcase
end

endmodule

module xpb_5_400
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h2cc260305d9dd832cb85ba8243f2bd2ee8f445a16a42656d11598f3a8a2f25bf5abcefc06d4d075222fd29c62dc3965d3bf03bbf42892461b8e189d67892284b8b024ef5d3c6f7f4574b5a5ea998da95f7fa4197293619dead2a04c54810aad06f1ace4015fdb915c21f2a491ca8a4187f78a309e2874a8db7f580742e2da392;
    5'b00010 : xpb = 1024'h5984c060bb3bb065970b750487e57a5dd1e88b42d484cada22b31e75145e4b7eb579df80da9a0ea445fa538c5b872cba77e0777e851248c371c313acf124509716049deba78defe8ae96b4bd5331b52beff4832e526c33bd5a54098a902155a0de359c802bfb722b843e549239514830fef14613c50e951b6feb00e85c5b4724;
    5'b00011 : xpb = 1024'h8647209118d9889862912f86cbd8378cbadcd0e43ec73047340cadaf9e8d713e1036cf4147e715f668f77d52894ac317b3d0b33dc79b6d252aa49d8369b678e2a106ece17b54e7dd05e20f1bfcca8fc1e7eec4c57ba24d9c077e0e4fd83200714d506ac041f92b41465d7edb55f9ec497e69e91da795dfa927e0815c8a88eab6;
    5'b00100 : xpb = 1024'h25c3b6bb4892c0263117231ff70ad6a325b1354d391f53cc789839475b9e9f567ab4188eb0d9eb9ec9667d1d3b048aa8ba6c716e771c13b32e6e7fba7762c7cb7ba07289f8ae28c4a9366d80d87a626ebe40cc418523a69ff1b811a661808af8d63a6d6a72debc981bcc2457ad26a38af08ad4539d1cd06996686cc2fd427dd;
    5'b00101 : xpb = 1024'h2f1e9b9c122704352e972cb443636a991b4f58f63dd45aa9d8e312ceffe90fb4c2683149585aa60c0f9391980173df07c79702d629fae59cebc871d2200854c842bc561e7351da80a1dec136b72080bce3de4e5b41885448ac4585dfae28b37ffc7e7516bd2ba4df43dbec8e977b0e512e81504f1c591794515c07405e01cb6f;
    5'b00110 : xpb = 1024'h5be0fbcc6fc4dc67fa1ce736875627c804439e97a816c016ea3ca2098a1835741d252109c5a7ad5e3290bb5e2f37756503873e956c8409fea4a9fba8989a7d13cdbea5144718d274f92a1b9560b95b52dbd88ff26abe6e27596f8aa4f6395e506b994356d3295df505fb16d7b423b269adf9f358fee06222095187b48c2f6f01;
    5'b00111 : xpb = 1024'h88a35bfccd62b49ac5a2a1b8cb48e4f6ed37e43912592583fb96314414475b3377e210ca32f4b4b0558de5245cfb0bc23f777a54af0d2e605d8b857f112ca55f58c0f40a1adfca69507575f40a5235e8d3d2d18993f4880606998f6a3e4a0920dab41196e927170ac81a4120d0cc56822d729662e167acafc1470828ba5d1293;
    5'b01000 : xpb = 1024'h4b876d769125804c622e463fee15ad464b626a9a723ea798f130728eb73d3eacf568311d61b3d73d92ccfa3a7609155174d8e2dcee3827665cdcff74eec58f96f740e513f15c5189526cdb01b0f4c4dd7c8198830a474d3fe370234cc30115f1ac74dad4e5bd7930379848af5a4d4715e115a8a73a39a0d32cd0d985fa84fba;
    5'b01001 : xpb = 1024'h317ad707c6b0303791a89ee642d418034daa6c4b11664fe6a06c966375a2f9aa2a1372d2436844c5fc29f969d52427b2533dc9ed116ca6d81eaf59cdc77e8144fa765d4712dcbd0cec72280ec4a826e3cfc25b1f59da8eb2ab6106fa1440bc2f89e21bed645990a8c598aed4124d7889dd89fd94562ae49aeac28e0c8dd5f34c;
    5'b01010 : xpb = 1024'h5e3d3738244e086a5d2e596886c6d532369eb1ec7ba8b553b1c6259dffd21f6984d06292b0b54c181f27233002e7be0f8f2e05ac53f5cb39d790e3a44010a9908578ac3ce6a3b50143bd826d6e410179c7bc9cb68310a891588b0bbf5c5166fff8fcea2d7a5749be87b7d91d2ef61ca25d02a09e38b22f28a2b80e80bc0396de;
    5'b01011 : xpb = 1024'h8aff976881ebe09d28b413eacab992611f92f78de5eb1ac0c31fb4d88a014528df8d52531e02536a42244cf630ab546ccb1e416b967eef9b90726d7ab8a2d1dc107afb32ba6aacf59b08dccc17d9dc0fbfb6de4dac46c27005b51084a46211d06817b86d905502d449d703664b9ec0badc7b43a81b3979b65aad8ef4ea313a70;
    5'b01100 : xpb = 1024'h714b2431d9b840729345695fe52083e971139fe7ab5dfb6569c8abd612dbde03701c49ac128dc2dc5c337757b10d9ffa2f45544b65543b198b4b7f2f6628576272e1579dea0a7a4dfba34882896f274c3ac264c48f6af3dfd52834f32481a0ea82af483f589c35c853646d070773eaa0d1a07cfad756713cc3394648f7c7797;
    5'b01101 : xpb = 1024'h33d712737b395c39f4ba11184244c56d80057f9fe4f8452367f619f7eb5ce39f91beb45b2e75e37fe8c0613ba8d4705cdee49103f8de6813519641c96ef4adc1b230646fb2679f9937058ee6d22fcd0abba667e3722cc91caa7c88147a58c4df1745c2c40b877c72475571198d1fe2c28c92aad98ffcb1a1842914d8bdaa1b29;
    5'b01110 : xpb = 1024'h609972a3d8d7346cc03fcb9a8637829c68f9c5414f3aaa90794fa932758c095eec7ba41b9bc2ead20bbd8b01d69806ba1ad4ccc33b678c750a77cb9fe786d60d3d32b365862e978d8e50e9457bc8a7a0b3a0a97a9b62e2fb57a68cd9c2696faf866091042185358809749b62a9c886db0c0b4de37283fc2f3c1e954cebd7bebb;
    5'b01111 : xpb = 1024'h8d5bd2d436750c9f8bc5861cca2a3fcb51ee0ae2b97d0ffd8aa9386cffbb2f1e473893dc090ff2242ebab4c8045b9d1756c508827df0b0d6c35955766018fe58c835025b59f58f81e59c43a425618236ab9aeb11c498fcda04d0919f0a7a1a7ff57b5f443782ee9dcb93c5abc6712af38b83f0ed550b46bcf41415c11a05624d;
    5'b10000 : xpb = 1024'h970edaed224b0098c45c8c7fdc2b5a8c96c4d534e47d4f31e260e51d6e7a7d59ead0623ac367ae7b2599f474ec122aa2e9b1c5b9dc704eccb9b9fee9dd8b1f2dee81ca27e2b8a312a4d9b60361e989baf9033106148e9a7fc6e0469986022be358e9b5a9cb7af2606f30915eb49a8e2bc22b514e747341a659a1b30bf509f74;
    5'b10001 : xpb = 1024'h36334ddf2fc2883c57cb834a41b572d7b26092f4b88a3a602f7f9d8c6116cd94f969f5e419838239d556c90d7c84b9076a8b581ae050294e847d29c5166ada3e69ea6b9851f282258198f5bedfb77331a78a74a78a7f0386a998092ee070cd8ea4a9699ab2b5683bc912335f07f24cfb3b9b581ec9ce7ea81d8f9ba4ed7e4306;
    5'b10010 : xpb = 1024'h62f5ae0f8d60606f23513dcc85a830069b54d89622cc9fcd40d92cc6eb45f3545426e5a486d0898bf853f2d3aa484f64a67b93da22d94db03d5eb39b8efd0289f4ecba8e25b97a19d8e4501d89504dc79f84b63eb3b51d6556c20df42881785f13c437dac8b321518b315da8249af113bb13fb28ac55c935d5851c191babe698;
    5'b10011 : xpb = 1024'h8fb80e3feafe38a1eed6f84ec99aed3584491e378d0f053a5232bc0175751913aee3d564f41d90de1b511c99d80be5c1e26bcf9965627211f6403d72078f2ad57fef0983f980720e302faa7c32e9285d977ef7d5dceb374403ec12b97092232f82df061adeb0da674d5087f14143952c3a8c9e328edd13c38d7a9c8d49d98a2a;
    5'b10100 : xpb = 1024'hbcd291a86addc0bef573af9fd336312fbc760a821d9ca2fe5af91e64ca191cb065847ac974419a19ef0071922716b54ba41e3728538c627fe8287ea454ede6f96a223cb1db66cbd74e1023843a63ec29b743fd4799b2411fb898583fe782b6dc2f2423143e59aef88afcb5b661c131b6b2b625a21190120ff00a1fcef24c751;
    5'b10101 : xpb = 1024'h388f894ae44bb43ebadcf57c41262041e4bba6498c1c2f9cf7092120d6d0b78a6115376d049120f3c1ed30df503501b1f6321f31c7c1ea89b76411c0bde106bb21a472c0f17d64b1cc2c5c96ed3f1958936e816ba2d13df0a8b38a494688d63e320d107159e354054acef5a482c4b733eaa4056403a04baeb6f622711d526ae3;
    5'b10110 : xpb = 1024'h6551e97b41e98c718662affe8518dd70cdafebeaf65e950a0862b05b60ffdd49bbd2272d71de2845e4ea5aa57df8980f32225af10a4b0eeb70459b9736732f06aca6c1b6c5445ca62377b6f596d7f3ee8b68c302cc0757cf55dd8f0e8e99810ea127deb16fe10d1b0cee1fed9f6d5b4c6a1ca86de627963c6eeba2e54b800e75;
    5'b10111 : xpb = 1024'h921449ab9f8764a451e86a80c90b9a9fb6a4318c60a0fa7719bc3f95eb2f0309168f16eddf2b2f9807e7846babbc2e6c6e1296b04cd4334d2927256daf05575237a910ac990b549a7ac311544070ce8483630499f53d71ae030793d3d6aa2bdf1042acf185dec630cf0d4a36bc15ff64e9954b77c8aee0ca26e1235979adb207;
    5'b11000 : xpb = 1024'he2964863b37080e5268ad2bfca4107d2e2273fcf56bbf6cad39157ac25b7bc06e0389358251b85b8b866eeaf621b3ff45e8aa896caa876331696fe5ecc50aec4e5c2af3bd414f49bf746910512de4e987584c9891ed5e7bfaa5069e6490341d5055e907eb1386b90a6c8da0e0ee7d541a340f9f5aeace27986728c91ef8ef2e;
    5'b11001 : xpb = 1024'h3aebc4b698d4e0411dee67ae4096cdac1716b99e5fae24d9be92a4b54c8aa17fc8c078f5ef9ebfadae8398b123e54a5c81d8e648af33abc4ea4af9bc65573337d95e79e99108473e16bfc36efac6bf7f7f528e2fbb23785aa7cf0b63aca0deedbf70b74801113fcecc8bb7e9fd97216c99acb2a93d7218b5505ca93d4d2692c0;
    5'b11010 : xpb = 1024'h67ae24e6f672b873e974223084898adb000aff3fc9f08a46cfec33efd6b9c73f237d68b65cebc6ffd180c27751a8e0b9bdc92207f1bcd026a32c8392dde95b836460c8df64cf3f326e0b1dcda45f9a15774ccfc6e459923954f91028f4b189be2e8b8588170ef8e48eaae2331a3fc585192555b31ff96343085229b17b543652;
    5'b11011 : xpb = 1024'h94708517541090a6b4f9dcb2c87c4809e8ff44e13432efb3e145c32a60e8ecfe7e3a5876ca38ce51f47dec3d7f6c7716f9b95dc73445f4885c0e0d69567b83ceef6317d538963726c556782c4df874ab6f47115e0d8fac18022314ee3cc2348e9da653c82d0cb1fa50ca0c7c36e8699d989df8bd0280add0c047aa25a981d9e4;
    5'b11100 : xpb = 1024'h10859ff1efc03410b57a1f5dfc14bde7607d8751c8fdb4a974c2990f381565b5d5aecabe6d5f5715781cd6bcc9d1fca9d18f71a0541c489e645057e1943b37690616321c5ccc31d60a07cfe85eb58b10733c595caa3f98e5f9c087b8caa83cccddb98fde924172828c294fe65bc0e78cc93cbce494bc9b2e31cdaf954ecd170b;
    5'b11101 : xpb = 1024'h3d4800224d5e0c4380ffd9e040077b164971ccf333401a16861c2849c2448b75306bba7edaac5e679b1a0082f79593070d7fad5f96a56d001d31e1b80ccd5fb491188112309329ca61532a47084e65a66b369af3d375b2c4a6ea8c7e12b8e79d4cd45e1ea83f2b984e487a2f78698ba548b55fee7743e5bbe9c330097cfaba9d;
    5'b11110 : xpb = 1024'h6a0a6052aafbe4764c85946283fa3845326612949d827f839775b7844c73b1348b28aa3f47f965b9be172a4925592964496fe91ed92e9161d6136b8e855f88001c1ad008045a21beb89e84a5b1e7403c6330dc8afcabcca3541491435ac9926dbbef2c5ebe3ce4ae1067a47895122fbdc82e02f859cb3049a1b8b07dab285e2f;
    5'b11111 : xpb = 1024'h96ccc0830899bca9180b4ee4c7ecf5741b5a583607c4e4f0a8cf46bed6a2d6f3e5e599ffb5466d0be114540f531cbfc1856024de1bb7b5c38ef4f564fdf1b04ba71d1efdd82119b30fe9df045b801ad25b2b1e2225e1e682013e9608a2da3d3e2b09fa9ed43a9dc3d286cec1b1bad3d647a6a6023c527ad759ae30f1d95601c1;
    endcase
end

endmodule

module xpb_5_645
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h72d7f7163bb1a02e5884115adc5234034af942a4cd466096e3e0f3b2099f67461233fa8c8632d154b5d2032fe429a83b71ecd774542034adb003e3504264b87cfe2256b69769803d4f431a88f211c37b7b0e23502a99000ec99ea900518a9de60fc2e46dd47616ee01424cae6698432b0fce35edaa44bc74a5d0e0cea6f99a1a;
    5'b00010 : xpb = 1024'h3502a8d6b5750b93e602aadea84a20b5247c8218c51520b649e52e0e603c2184211f77a0423f241acc45c718e4f53fac7fbf8702858d990faf68874249f6fc4887f578be7f4203358bec326f4b47c2c602174d07c8abd30cddb0c005e8ea9939f07e36b1f823354e7bc4b27dd560602cd0c28cf9043e1bb905324698c510cdc9;
    5'b00011 : xpb = 1024'ha7da9fecf126abc23e86bc39849c54b86f75c4bd925b814d2dc621c069db88ca3353722cc871f56f8217ca48c91ee7e7f1ac5e76d9adcdbd5f6c6a928c5bb4c58617cf7516ab8372db2f4cf83d5986417d257057f344d31ba74f69063a75372000411b1fcc994c3c7d06ff2c3bf8a357e090c2e6ae82d82dab0327676c0a67e3;
    5'b00100 : xpb = 1024'h6a0551ad6aea1727cc0555bd5094416a48f904318a2a416c93ca5c1cc0784308423eef40847e4835988b8e31c9ea7f58ff7f0e050b1b321f5ed10e8493edf8910feaf17cfe84066b17d864de968f858c042e9a0f9157a619bb61800bd1d53273e0fc6d63f0466a9cf78964fbaac0c059a18519f2087c37720a648d318a219b92;
    5'b00101 : xpb = 1024'h2c30036de4ad828d5983ef411c8c2e1c227c43a581f9018bf9ce96791714fd46512a6c54408a9afbaeff521acab616ca0d51bd933c8896815e35b2769b803c5c99be1384e65c896354817cc4efc584d68b37c3c72f6a7917cf73971169352dc7c1b7bfa813f388fd720bcacb1988dd5b627970fd627596b669c5f2fba838cf41;
    5'b00110 : xpb = 1024'h9f07fa84205f22bbb208009bf8de621f6d75864a4f3f6222ddaf8a2b20b4648c635e66e0c6bd6c5064d1554aaedfbf057f3e950790a8cb2f0e3995c6dde4f4d997e06a3b7dc609a0a3c4974de1d748520645e7175a03792699124011babfcbadd17aa415e8699feb734e1779802120867247a6eb0cba532b0f96d3ca4f32695b;
    5'b00111 : xpb = 1024'h6132ac449a228e213f869a1fc4d64ed146f8c5be470e224243b3c48777511eca7249e3f482c9bf167b451933afab56768d114495c2162f910d9e39b8e57738a521b38c43659e8c98e06daf343b0d479c8d4f10cef8164c24ad245717521fc701b235f65a0c16be4bedd07d48eee93d88333bfdf666b3b26f6ef839946d499d0a;
    5'b01000 : xpb = 1024'h235d5e0513e5f986cd0533a390ce3b83207c05323edce261a9b7fee3cdedd908813561083ed611dc91b8dd1cb076ede79ae3f423f38393f30d02ddaaed097c70ab86ae4b4d770f911d16c71a944346e714583a8696291f22c1366e1ce97fc25592f1489e2fc3dcac6852e3185db15a89f4305501c0ad11b3ce599f5e8b60d0b9;
    5'b01001 : xpb = 1024'h9635551b4f9799b5258944fe6d206f866b7547d70c2342f88d98f295d78d404e93695b94c508e331478ae04c94a096230cd0cb9847a3c8a0bd06c0fb2f6e34eda9a90501e4e08fce6c59e1a386550a628f665dd6c0c21f318ad5171d3b0a603ba2b42d0c0439f39a69952fc6c4499db503fe8aef6af1ce28742a802d325a6ad3;
    5'b01010 : xpb = 1024'h586006dbc95b051ab307de8239185c3844f8874b03f20317f39d2cf22e29fa8ca254d8a8811535f75dfea435956c2d941aa37b2679112d02bc6b64ed370078b9337c2709ccb912c6a902f989df8b09ad166f878e5ed4f22f9ee72e22d26a5b8f836f7f5027e711fae41795963311bab6c4f2e1fac4eb2d6cd38be5f750719e82;
    5'b01011 : xpb = 1024'h1a8ab89c431e708040867806051048ea1e7bc6befbc0c33759a1674e84c6b4cab14055bc3d2188bd7472681e9637c50528762ab4aa7e9164bbd008df3e92bc84bd4f4911b49195bee5ac117038c108f79d78b145fce7c52db2f9452869ca56e3642ad1944b94305b5e99fb65a1d9d7b885e739061ee48cb132ed4bc16e88d231;
    5'b01100 : xpb = 1024'h8d62afb27ed010ae990a8960e1627ced69750963c90723ce3d825b008e661c10c3745048c3545a122a446b4e7a616d409a630228fe9ec6126bd3ec2f80f77501bb719fc84bfb15fc34ef2bf92ad2cc731886d4962780c53c7c97ee28bb54f4c973edb602200a47495fdc481408721ae395b56ef3c9294925d8be2c9015826c4b;
    5'b01101 : xpb = 1024'h4f8d6172f8937c14268922e4ad5a699f42f848d7c0d5e3eda386955ce502d64ed25fcd5c7f60acd840b82f377b2d04b1a835b1b7300c2a746b3890218889b8cd4544c1d033d398f4719843df8408cbbd9f8ffe4dc593983a90aa052e52b4f01d54a9084643b765a9da5eade3773a37e556a9c5ff2322a86a381f925a33999ffa;
    5'b01110 : xpb = 1024'h11b813337256e779b407bc68795256511c7b884bb8a4a40d098acfb93b9f908ce14b4a703b6cff9e572bf3207bf89c22b608614561798ed66a9d3413901bfc98cf17e3d81bac1becae415bc5dd3ecb082699280563a66b38a4bc1c33ea14eb7135645a8a6764840a54e113b2e60254e7179e1d0a7d1c07ae9780f82451b0d3a9;
    5'b01111 : xpb = 1024'h84900a49ae0887a80c8bcdc355a48a546774caf085eb04a3ed6bc36b453ef7d2f37f44fcc19fd0f30cfdf6506022445e27f538b9b599c3841aa11763d280b515cd3a3a8eb3159c29fd84764ecf508e83a1a74b558e3f6b476e5ac5343b9f895745273ef83bda9af8562360614c9a9812276c52f82760c4233d51d8f2f8aa6dc3;
    5'b10000 : xpb = 1024'h46babc0a27cbf30d9a0a6747219c770640f80a647db9c4c3536ffdc79bdbb211026ac2107dac23b92371ba3960eddbcf35c7e847e70727e61a05bb55da12f8e1570d5c969aee1f223a2d8e3528868dce28b0750d2c523e45826cdc39d2ff84ab25e2913c5f87b958d0a5c630bb62b513e860aa03815a23679cb33ebd16c1a172;
    5'b10001 : xpb = 1024'h8e56dcaa18f5e73278900caed9463b81a7b49d8758884e2b9743823f2786c4f11563f2439b8767f39e57e2261b97340439a97d618748c48196a5f47e1a53cace0e07e9e82c6a21a76d6a61b81bc8d18afb99ec4ca651143967ef33f6a5f7fff069de3808334d7b94b282c002a2ad215a955010edb5382abfc14a48734d8d521;
    5'b10010 : xpb = 1024'h7bbd64e0dd40fea1800d1225c9e697bb65748c7d42cee5799d552bd5fc17d395238a39b0bfeb47d3efb7815245e31b7bb5876f4a6c94c0f5c96e42982409f529df02d5551a302257c619c0a473ce50942ac7c214f4fe1152601d9c3fbbea1de51660c7ee57aaeea74c6a78ae90c31540b92336fc85983f20a1e58555dbd26f3b;
    5'b10011 : xpb = 1024'h3de816a157046a070d8baba995de846d3ef7cbf13a9da5990359663252b48dd33275b6c47bf79a9a062b453b46aeb2ecc35a1ed89e022557c8d2e68a2b9c38f568d5f75d0208a55002c2d88acd044fdeb1d0ebcc9310e450742fb345534a1938f71c1a327b580d07c6ecde7dff8b32427a178e07df919e650146eb1ff9e9a2ea;
    5'b10100 : xpb = 1024'h12c861d0c7d56c9b0a452d61d6711f187b0b65326c65b8695da08ea9514811416133d83803ed601c9f0924477a4a5dd12cce66cf6f89b9c8378a7c332e7cc0f2a91964e9e128483f6bf071263a4f2938da15843123b74e8841ca4aeaaa148cd7d76c769f052b68416f444d6e534f443b0be513398afda960a850ea1800d699;
    5'b10101 : xpb = 1024'h72eabf780c79759af38e56883e28a52263744e09ffb2c64f4d3e9440b2f0af5753952e64be36beb4d2710c542ba3f2994319a5db238fbe67783b6dcc7593353df0cb701b814aa8858eaf0afa184c12a4b3e838d45bbcb75d51e0734b3c34b272e79a50e4737b425642b190fbd4eb926f4ada1b00e3cfba1e067931b8befa70b3;
    5'b10110 : xpb = 1024'h35157138863ce100810cf00c0a2091d43cf78d7df781866eb342ce9d098d69956280ab787a43117ae8e4d03d2c6f8a0a50ec556954fd22c977a011be7d2579097a9e922369232b7dcb5822e0718211ef3af1628bf9cf8a5b65f28a50d394adc6c855a328972860b6bd33f6cb43b3af710bce720c3dc9196265da9782dd11a462;
    5'b10111 : xpb = 1024'ha7ed684ec1ee812ed9910166e672c5d787f0d022c4c7e7059723c24f132cd0db74b4a6050075e2cf9eb6d36d10993245c2d92cdda91d577727a3f50ebf8a318678c0e8da008cabbb1a9b3d696393d56ab5ff85dc24688a6a2f913351251f4bacd81887966b9e77a4be764379aa4bf29c1b9ca7f9e80dd5d70bab7851840b3e7c;
    5'b11000 : xpb = 1024'h6a181a0f3bb1ec94670f9aeab26ab28961740f96bc96a724fd27fcab69c98b1983a02318bc823595b52a97561164c9b6d0abdc6bda8abbd927089900c71c755202940ae1e8652eb35744554fbcc9d4b53d08af93c27b5d6843a34a56bc7f4700b8d3d9da8f4b960538f8a94919140f9ddc90ff054207351b6b0cde1ba222722b;
    5'b11001 : xpb = 1024'h2c42cbcfb57557f9f48e346e7e629f3b3af74f0ab4656744632c3707c0664557928ba02c788e885bcb9e5b3f12306127de7e8bfa0bf8203b266d3cf2ceaeb91d8c672ce9d03db1ab93ed6d3615ffd3ffc411d94b608e306657b5615c53df4254998f2c1eb2f8b465b37b0f1887dc2c9f9d8556109c00945fca6e43e5c039a5da;
    5'b11010 : xpb = 1024'h9f1ac2e5f126f8284d1245c95ab4d33e85f091af81abc7db470d2ab9ca05ac9da4bf9ab8fec159b081705e6ef65a0963506b636e601854e8d67120431113719a8a8983a067a731e8e33087bf0811977b3f1ffc9b8b27307521540a5ca569e03aa952108c876ecb53b4bd5bc6ee746fcaad538bfe464550d4703f24b467333ff4;
    5'b11011 : xpb = 1024'h614574a66aea638dda90df4d26acbff05f73d123797a87faad11651620a266dbb3ab17ccbacdac7697e42257f725a0d45e3e12fc9185b94ad5d5c43518a5b566145ca5a84f7fb4e11fd99fa5614796c5c6292653293a0373356621623cc9db8e8a0d62d0ab1be9b42f3fc1965d3c8ccc6e47e309a03eb018cfa08a7e854a73a3;
    5'b11100 : xpb = 1024'h23702666e4adcef3680f78d0f2a4aca238f710977149481a13159f72773f2119c29694e076d9ff3cae57e640f7f138456c10c28ac2f31dacd53a68272037f9319e2fc7b0375837d95c82b78bba7d96104d32500ac74cd67149783867d429d6e26ac8b514cec90814a9c22765cc04a9ce2f3c3a14fa380f5d2f01f048a361a752;
    5'b11101 : xpb = 1024'h96481d7d205f6f21c0938a2bcef6e0a583f0533c3e8fa8b0f6f6932480de885fd4ca8f6cfd0cd0916429e970dc1ae080ddfd99ff1713525a853e4b77629cb1ae9c521e66cec1b816abc5d214ac8f598bc840735af1e5d6801316e16825b474c87a8b9982a33f1f02ab047414329cecf93f0a7002a47ccbd1d4d2d1174a5b416c;
    5'b11110 : xpb = 1024'h5872cf3d9a22da874e1223af9aeecd575d7392b0365e68d05cfacd80d77b429de3b60c80b91923577a9dad59dce677f1ebd0498d4880b6bc84a2ef696a2ef57a2625406eb69a3b0ee86ee9fb05c558d64f499d128ff8a97e2728f86dbd14701c5b46ebc6c6ec3d632586d9e3a16509fafffec70dfe762b16343436e16872751b;
    5'b11111 : xpb = 1024'h1a9d80fe13e645ecdb90bd3366e6ba0936f6d2242e2d28efc2ff07dd2e17fcdbf2a189947525761d91117142ddb20f62f9a2f91b79ee1b1e8407935b71c13945aff862769e72be07251801e15efb5820d652c6ca2e0b7c7c3b3b0f7354746b703c023e0aea995bc3a0093fb3102d26fcc0f31e19586f8a5a93959cab8689a8ca;
    endcase
end

endmodule

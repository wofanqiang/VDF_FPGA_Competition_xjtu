module xpb_5_975
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h80fb1db1364c0318a055539b87f9424cb447214c88b2cffc1d8e362971547263d6d61267d99c3e05fa5d5122d58dff836784187f34bf6e65362963a18d75d78fbc0e2c3ebf28ccb9d45a40ef39ac6c3652d342d8066b61933c4195c4b3aa9cfea3eb5fd5d27b4e9bdf5aea08eca1bbdd2aceb43b454c1d36cfb838a095c5e97b;
    5'b00010 : xpb = 1024'h5148f60caaa9d16875a52f5fff983d47f7183f683bedff80bd3fb2fd2fa637bfaa63a756e911fd7d555c62fec7bdee3c6aee091846cc0c7ebbb387e4e0193a6e03cd23cecec09c2e961a7f3bda7d143bb1a18c1780509615c2f6998ead2a976b18cf2d81f42da4aa37f5ed32e173519106c389943a4cdd3d5900f63ca2a96c8b;
    5'b00011 : xpb = 1024'h2196ce681f079fb84af50b247737384339e95d83ef292f055cf12fd0edf7fd1b7df13c45f887bcf4b05b74dab9eddcf56e57f9b158d8aa98413dac2832bc9d4c4b8c1b5ede586ba357dabd887b4dbc41106fd556fa35ca9849ab9d58a6aa91d78db2fb2e15dffab89090f05cd644e744e2b85eed2f4d9d43e249b3d8af8cef9b;
    5'b00100 : xpb = 1024'ha291ec195553a2d0eb4a5ebfff307a8fee307ed077dbff017a7f65fa5f4c6f7f54c74eadd223fafaaab8c5fd8f7bdc78d5dc12308d9818fd77670fc9c03274dc079a479d9d81385d2c34fe77b4fa28776343182f00a12c2b85ed331d5a552ed6319e5b03e85b49546febda65c2e6a3220d8713287499ba7ab201ec794552d916;
    5'b00101 : xpb = 1024'h72dfc474c9b17120c09a3a8476cf758b31019cec2b172e861a30e2ce1d9e34db2854e39ce199ba7205b7d7d981abcb31d94602c99fa4b716fcf1340d12d5d7ba4f593f2dad1907d1edf53cc455cad07cc211616e7a8660ae0ca236e753d52942a68228b00a0d9f62c886dd8fb7b838d5e97be881699a7a813b4aaa1552365c26;
    5'b00110 : xpb = 1024'h432d9cd03e0f3f7095ea1648ee6e708673d2bb07de525e0ab9e25fa1dbeffa36fbe2788bf10f79e960b6e9b573dbb9eadcaff362b1b15530827b585065793a98971836bdbcb0d746afb57b10f69b788220dfaaadf46b953093573ab14d5523af1b65f65c2bbff5712121e0b9ac89ce89c570bdda5e9b3a87c49367b15f19df36;
    5'b00111 : xpb = 1024'h137b752bb26d0dc06b39f20d660d6b81b6a3d923918d8d8f5993dc759a41bf92cf700d7b00853960bbb5fb91660ba8a3e019e3fbc3bdf34a08057c93b81c9d76ded72e4dcc48a6bb7175b95d976c20877fadf3ed6e50c9b31a0c3e7b46d51e1b9049c4084d724b7f79bce3e3a15b643da1659333539bfa8e4ddc254d6bfd6246;
    5'b01000 : xpb = 1024'h947692dce8b910d90b8f45a8ee06adce6aeafa701a405d8b7722129f0b9631f6a6461fe2da217766b6134cb43b99a827479dfc7af87d61af3e2ee035459275069ae55a8c8b71737545cffa4cd1188cbdd28136c574bc2b46564dd43ffa7fbb1a343523de1fed9a1b5917cdec8dfd201acc34476e98e817c51d945dee01c34bc1;
    5'b01001 : xpb = 1024'h64c46b385d16df28e0df216d65a5a8c9adbc188bcd7b8d1016d38f72c9e7f75279d3b4d1e99736de11125e902dc996e04b07ed140a89ffc8c3b904789835d7e4e2a4521c9b0942ea0790389971e934c3314f8004eea15fc8dd02d809f3ffb586a918f18a419ff029b1b2d11682ceb5cea8291cc78de8d7cba6dd1b8a0ea6ced1;
    5'b01010 : xpb = 1024'h35124393d174ad78b62efd31dd44a3c4f08d36a780b6bc94b6850c468839bcae4d6149c0f90cf6556c11706c1ff985994e71ddad1c969de2494328bbead93ac32a6349acaaa1125ec95076e612b9dcc8901dc9446886944b63b7dbd3ed7faff31dfcbf36635246380a4dd44077a04b82841df22082e997d23025d9261b8a51e1;
    5'b01011 : xpb = 1024'h5601bef45d27bc88b7ed8f654e39ec0335e54c333f1ec195636891a468b820a20eedeb00882b5ccc71082481229745251dbce462ea33bfbcecd4cff3d7c9da17222413cba38e1d38b10b532b38a84cdeeec1283e26bc8cdea6cdf9de6ffaa5f92e08ce285049c4662e8d76a6c71e1366012c77977ea57d8b96e96c2286dd4f1;
    5'b01100 : xpb = 1024'h865b39a07c1e7ee12bd42c91dcdce10ce7a5760fbca4bc1573c4bf43b7dff46df7c4f117e21ef3d2c16dd36ae7b773d5b95fe6c56362aa6104f6b0a0caf275312e306d7b7961ae8d5f6af621ed36f10441bf555be8d72a6126ae75629aaa475e36cbecb8577feae24243c17359139d138ae17bb4bd36750f8926cf62be33be6c;
    5'b01101 : xpb = 1024'h56a911fbf07c4d3101240856547bdc082a76942b6fdfeb9a13763c177631b9c9cb528606f194b34a1c6ce546d9e7628ebcc9d75e756f487a8a80d4e41d95d80f75ef650b88f97e02212b346e8e079909a08d9e9b62bc5ee3ad63792c942a41caabafba64793240f09adec49d4de532c766d6510db2373516126f8cfecb17417c;
    5'b01110 : xpb = 1024'h26f6ea5764da1b80d673e41acc1ad7036d47b247231b1b1eb327b8eb34837f259ee01af6010a72c1776bf722cc175147c033c7f7877be694100af92770393aedbdae5c9b98914d76e2eb72bb2ed8410eff5be7dadca1936634187cf68daa3c37209388109ae496fef379c7c742b6c87b42cb2666a737f51c9bb84a9ad7fac48c;
    5'b01111 : xpb = 1024'ha7f208089b261e9976c937b654141950218ed393abcdeb1ad0b5ef14a5d7f18975b62d5ddaa6b0c771c94845a1a550cb27b7e076bc3b54f946345cc8fdaf127d79bc88da57ba1a30b745b3aa6884ad45522f2ab2e30cf4f9705a12bb4154d935c47ee7e66d5fe59ad2d4b1d02f5884586d99daa1ec8412536b70833b6dc0ae07;
    5'b10000 : xpb = 1024'h783fe0640f83ece94c19137acbb3144b645ff1af5f091a9f70676be86429b6e54943c24cea1c703eccc85a2193d53f842b21d10fce47f312cbbe810c5052755bc17b806a6751e9a57905f1f70955554ab0fd73f25cf2297bf70f16853ad4d3a23962b5928f123ba92b6fb4fa242a1a0c498eaffae184d259f4b940d77aa43117;
    5'b10001 : xpb = 1024'h488db8bf83e1bb392168ef3f43520f46a7310fcb12444a241018e8bc227b7c411cd1573bf9922fb627c76bfd86052e3d2e8bc1a8e054912c5148a54fa2f5d83a093a77fa76e9b91a3ac63043aa25fd500fcbbd31d6d75dfe7dc41a4f3454ce0eae46833eb0c491b7840ab82418fbafc025838553d68592607e01fe738787b427;
    5'b10010 : xpb = 1024'h18db911af83f8988f6b8cb03baf10a41ea022de6c57f79a8afca658fe0cd419cf05eec2b0907ef2d82c67dd978351cf631f5b241f2612f45d6d2c992f5993b1850f96f8a8681888efc866e904af6a5556e9a067150bc928104791e192dd4c87b232a50ead276e7c5dca5bb4e0dcd457401785aaccb865267074abc0f946b3737;
    5'b10011 : xpb = 1024'h99d6aecc2e8b8ca1970e1e9f42ea4c8e9e494f334e3249a4cd589bb95221b400c734fe92e2a42d337d23cefc4dc31c799979cac127209dab0cfc2d34830f12a80d079bc945aa5548d0e0af7f84a3118bc16d49495727f41440bab3dde17f6579c715b0c0a4f23661bc00a556fa6f01512c470ee810d26f9dd702f4b02a3120b2;
    5'b10100 : xpb = 1024'h6a248727a2e95af16c5dfa63ba894789e11a6d4f016d79296d0a188d1073795c9ac29381f219ecaad822e0d83ff30b329ce3bb5a392d3bc492865177d5b2758654c69359554224bd92a0edcc2573b991203b9288d10d2896c76fb7a7daff5fe63bf97e6cc6a48c70149ba880ef409705083be44105d32fa4604bb24c3714a3c2;
    5'b10101 : xpb = 1024'h3a725f831747294141add6283228428523eb8b6ab4a8a8ae0cbb9560cec53eb86e502871018fac223321f2b43222f9eba04dabf34b39d9de181075bb2855d8649c858ae964d9f43254612c18c64461967f09dbc84af25d194e24bb71d47f5a52b0dd4c18e856e27e6d36abaae4122cb8e430b999fad3efaae9946fe843f826d2;
    5'b10110 : xpb = 1024'hac037de8ba4f79116fdb1eca9c73d8066bca98667e3d832ac6d12348d17041441ddbd6011056b998e2104902452e8a4a3b79c8c5d4677f79d9a99fe7af93b42e44482797471c3a716216a656715099bddd82507c4d7919bd4d9bf3bcdff54bf25c119c50a09388cc5d1aed4d8e3c26cc0258ef2efd4afb172dd2d8450dba9e2;
    5'b10111 : xpb = 1024'h8bbb558fc1f0faa9b753058831c07fcd1b03cad2f096a82ec9fb485dfe6b767818b3cfc7eaa1a99f887e55b2f9e0e8280b3bb50b9205e65cd3c3fda0086f12d2a052aeb8339a9060ea7bab54a0c175d230ab67dfcb42f32f111b550081a9f1bdc9ac799adc848728a52c98ddc5857e49eaf4432e3520cce842956624e6a1935d;
    5'b11000 : xpb = 1024'h5c092deb364ec8f98ca2e14ca95f7ac85dd4e8eea3d1d7b369acc531bcbd3bd3ec4164b6fa176916e37d678eec10d6e10ea5a5a4a4128476594e21e35b1275b0e811a64843325fd5ac3be9a141921dd78f79b11f452827b197d058ca7b29ec2a3e904746fe36dd36fdc79c07ba5713fdc6e918872a218ceecbde23c0f385166d;
    5'b11001 : xpb = 1024'h2c570646aaac974961f2bd1120fe75c3a0a6070a570d0738095e42057b0f012fbfcef9a6098d288e3e7c796ade40c59a120f963db61f228fded84626adb5d88f2fd09dd852ca2f4a6dfc27ede262c5dcee47fa5ebf0d5c341e855c9474a9e696b37414f31fe9334556629f31af28a9b1a2ddede01f224cf55526e15d0068997d;
    5'b11010 : xpb = 1024'had5223f7e0f89a62024810aca8f7b81054ed2856dfbfd73426ec782eec63739396a50c0de329669438d9ca8db3cec51d7993aebceade90f51501a9c83b2bb01eebdeca1711f2fc04425668dd1c0f3213411b3d36c578bdc75ac6f25928548395575f74c8f26481e135bd893a9bca658ecdaca21b646e6a2c24df19fd962e82f8;
    5'b11011 : xpb = 1024'h7d9ffc53555668b1d797ec712096b30b97be467292fb06b8c69df502aab538ef6a32a0fcf29f260b93d8dc69a5feb3d67cfd9f55fceb2f0e9a8bce0b8dcf12fd339dc1a7218acb790416a729bcdfda189fe986763f5df249e17bf62321d47e01cc4342751416d7ef8e588c64909bfb42a9a17774596f2a32ae27d799a3120608;
    5'b11100 : xpb = 1024'h4dedd4aec9b43701ace7c8359835ae06da8f648e4636363d664f71d66906fe4b3dc035ec0214e582eed7ee45982ea28f80678fef0ef7cd282015f24ee07275db7b5cb93731229aedc5d6e5765db0821dfeb7cfb5b94326cc6830f9ed1b54786e4127102135c92dfde6f38f8e856d90f685964ccd4e6fea3937709535aff58918;
    5'b11101 : xpb = 1024'h1e3bad0a3e1205518237a3fa0fd4a9021d6082a9f97165c20600eeaa2758c3a7114dcadb118aa4fa49d700218a5e914883d1808821046b41a5a016923315d8b9c31bb0c740ba6a62879723c2fe812a235d8618f533285b4eeee5fdb714d472dab60addcd577b840c3f8e92b87a3f26aa618b22264370aa3fc0b952d1bcd90c28;
    5'b11110 : xpb = 1024'h9f36cabb745e086a228cf79597cdeb4ed1a7a3f6822435be238f24d398ad360ae823dd42eb26e300443451445fec90cbeb55990755c3d9a6dbc97a33c08bb0497f29dd05ffe3371c5bf164b2382d9659b0595bcd3993bce22b27937bc87f0fd959f63da329f6d2a81ee97cc166e0e2878c59d66188bcc77690718b72529ef5a3;
    5'b11111 : xpb = 1024'h6f84a316e8bbd6b9f7dcd35a0f6ce64a1478c212355f6542c340a1a756fefb66bbb17231fa9ca2779f336320521c7f84eebf89a067d077c061539e77132f1327c6e8d4960f7b06911db1a2fed8fe3e5f0f27a50cb378f164b1dc9745c1ff0a45ceda0b4f4ba928b677847feb5bb2783b684eabba7dbd877d19ba490e5f8278b3;
    endcase
end

endmodule

module xpb_5_1010
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h88694707dc9206ca465a13ae245ae2c27eeee7354d29c9560bf8264d603c78eac3d3aad5d73438ed4ff519ff3cf3167fd309076c402ecacd91c51a3a922fa429c5f1723b152bd1fc5a2900534b897891baede5580782b68374ce0a06e756c0b6f5aa49d020bcbad3a3f0b6fb4378d93abe0593f82c6d1e505760f8483b921306;
    5'b00010 : xpb = 1024'h602548b9f735d8cbc1aeaf85385b7e338c67cb39c4dbf2349a1393450d7644cd845ed832e441f34c008bf4b796881c3541f7e6f25daac54f72eaf516e98cd3a21793afc77ac6a6b3a1b7fe03fe372cf281d6d117827f3ff6340f82131482dedbbc4d017690b07d19c12187178f218c4c2d31490e088edf706852758bee41bfa1;
    5'b00011 : xpb = 1024'h37e14a6c11d9aacd3d034b5c4c5c19a499e0af3e3c8e1b13282f003cbab010b044ea058ff14fadaab122cf6ff01d21eab0e6c6787b26bfd15410cff340ea031a6935ed53e0617b6ae946fbb4b0e4e15348bfbcd6fd7bc968f350fa1f41aefd0082efb91d00a43f5fde525733daca3f5d9c5cfe23e4b0a0907943f2cfa0f16c3c;
    5'b00100 : xpb = 1024'hf9d4c1e2c7d7cceb857e733605cb515a7599342b44043f1b64a6d3467e9dc93057532ecfe5d680961b9aa2849b227a01fd5a5fe98a2ba533536aacf98473292bad82ae045fc502230d5f965639295b40fa8a896787852dbb292722b6edb1b25499270c3709801a5fb8327502672f26f0b88b339c0d261b08a35701353a118d7;
    5'b00101 : xpb = 1024'h98069326090f8398feb1fae184b797d826487a78016a0d47c2429381c826557dc948ddc2d591a0f6b1aec42786a53e1ff2dead6ad8d18520c6fbc50a2a76d6bc80c99d1b5b28221e8afef9b8af1c0e45ca968dee7ffb095f27607c325631dbdc3f3cba939154bc799f73de4b69ebcba9c98e4731ed3f8000e196685b8f332bdd;
    5'b00110 : xpb = 1024'h6fc294d823b3559a7a0696b898b8334933c15e7c791c3626505e00797560216089d40b1fe29f5b5562459edfe03a43d561cd8cf0f64d7fa2a8219fe681d40634d26bdaa7c0c2f6d5d28df76961c9c2a6917f79adfaf792d1e6a1f43e835dfa0105df723a01487ebfbca4ae67b5947ebb38b9fc47c9614120f287e59f41e2d878;
    5'b00111 : xpb = 1024'h477e968a3e57279bf55b328facb8ceba413a4280f0ce5f04de796d712299ed434a5f387cefad15b412dc799839cf498ad0bc6c7713c97a2489477ac2d93135ad240e1834265dcb8d1a1cf51a147777075868656d75f41c44a5e36c4ab08a1825cc8229e0713c4105d9d57e84013d31cca7e5b15da5830241037962e2f4928513;
    5'b01000 : xpb = 1024'h1f3a983c58faf99d70afce66c0b96a2b4eb32685688087e36c94da68cfd3b9260aea65d9fcbad012c373545093644f403fab4bfd314574a66a6d559f308e652575b055c08bf8a04461abf2cac7252b681f51512cf0f0a5b76524e456ddb6364a9324e186e130034bf7064ea04ce5e4de1711667381a4c361146ae026a74231ae;
    5'b01001 : xpb = 1024'ha7a3df44358d0067b709e214e5144cedcda20dbab5aa5139788d00b630103210cebe10afd3ef090013686e4fd05765c012b4536971743f73fc326fd9c2be094f3ba1c7fba1247240bbd4f31e12aea3f9da3f3684f8735c3ad9f2ee5dc50cf70188cf2b5701ecbe1f9af7059b905ebe18d516fa6bae11e1b16bcbd86ee2d444b4;
    5'b01010 : xpb = 1024'h7f5fe0f65030d269325e7debf914e85edb1af1bf2d5c7a1806a86daddd49fdf38f493e0ce0fcc35ec3ff490829ec6b7581a332ef8ef039f5dd584ab61a1b38c78d44058806bf46f80363f0cec55c585aa1282244736fe5ad99346669f23915264f71e2fd71e08065b827d5b7dc07712a4442af818a33a2d17cbd55b29583f14f;
    5'b01011 : xpb = 1024'h571be2a86ad4a46aadb319c30d1583cfe893d5c3a50ea2f694c3daa58a83c9d64fd46b69ee0a7dbd749623c08381712af0921275ac6c3477be7e25927178683fdee643146c5a1baf4af2ee7f780a0cbb68110e03ee6c6f205875de761f65334b16149aa3e1d442abd558a5d427b0243bb36e6497665563f18daed2f648339dea;
    5'b01100 : xpb = 1024'h2ed7e45a8578766c2907b59a21161f40f60cb9c81cc0cbd522df479d37bd95b9105f98c6fb18381c252cfe78dd1676e05f80f1fbc9e82ef99fa4006ec8d597b8308880a0d1f4f0669281ec302ab7c11c2ef9f9c36968f89317b756824c91516fdcb7524a51c804f1f28975f07358d74d229a19ad427725119ea05039fae34a85;
    5'b01101 : xpb = 1024'h693e60ca01c486da45c51713516bab203859dcc9472f4b3b0fab494e4f7619bd0eac6240825f27ad5c3d93136ab7c95ce6fd181e764297b80c9db4b2032c730822abe2d378fc51dda10e9e0dd65757cf5e2e582e4658205d6f8ce8e79bd6f94a35a09f0c1bbc7380fba460cbf018a5e91c5cec31e98e631af91cd7dad92f720;
    5'b01110 : xpb = 1024'h8efd2d147cae4f37eab6651f59719d7482748501e19cbe09bcf2dae24533da8694be70f9df5a2b6825b8f330739e9315a178d8ee2792f449128ef585b2626b5a481c30684cbb971a3439ea3428eeee0eb0d0cadaebe838894bc6d8956114304b990453c0e278820bb3aafd08027a63994fcb62bb4b06048206f2c5c5e9250a26;
    5'b01111 : xpb = 1024'h66b92ec697522139660b00f66d7238e58fed6906594ee6e84b0e47d9f26da66955499e56ec67e5c6d64fcde8cd3398cb1067b874450eeecaf3b4d06209bf9ad299be6df4b2566bd17bc8e7e4db9ca26f77b9b69a66e4c1fc0b0850a18e404e705fa70b67526c4451d0dbcd244e2316aabef717d12727c5a217e443099bd4b6c1;
    5'b10000 : xpb = 1024'h3e753078b1f5f33ae15f9ccd8172d4569d664d0ad1010fc6d929b4d19fa7724c15d4cbb3f975a02586e6a8a126c89e807f5697fa628ae94cd4daab3e611cca4aeb60ab8117f14088c357e5958e4a56d03ea2a259e1e14b6eca49c8adbb6c6c952649c30dc2600697ee0c9d4099cbc9bc2e22cce7034986c228d5c04d4e84635c;
    5'b10001 : xpb = 1024'h1631322acc99c53c5cb438a495736fc7aadf310f48b338a5674521c94ce13e2ed65ff91106835a84377d8359805da435ee4577808006e3ceb600861ab879f9c33d02e90d7d8c15400ae6e34640f80b31058b8e195cddd4e1898b40b9e8988ab9ecec7ab43253c8de0b3d6d5ce5747ccd9d4e81fcdf6b47e239c73d9101340ff7;
    5'b10010 : xpb = 1024'h9e9a7932a92bcc06a30e4c52b9ce528a29ce184495dd01fb733d4816ad1db7199a33a3e6ddb7937187729d58bd50bab5c14e7eecc035ae9c47c5a0554aa99ded02f45b4892b7e73c650fe3998c8183c2c079737164608b64fe594ac0cfef4b70e296c484531083b1af2e245828ed56085b5415f50bd86632912835d93cc622fd;
    5'b10011 : xpb = 1024'h76567ae4c3cf9e081e62e829cdceedfb3746fc490d8f2ada0158b50e5a5782fc5abed143eac54dd03809781116e5c06b303d5e72ddb1a91e28eb7b31a206cd65549698d4f852bbf3ac9ee14a3f2f382387625f30df5d14d7bd9ac2ccfd1b6995a9397c2ac30445f7cc5ef47474960919ca7fcb0ae7fa2752a219b31cef75cf98;
    5'b10100 : xpb = 1024'h4e127c96de73700999b78400e1cf896c44bfe04d854153b88f74220607914edf1b49fea0f7d3082ee8a052c9707ac6209f2c3df8fb2da3a00a11560df963fcdda638d6615ded90aaf42ddefaf1dcec844e4b4af05a599e4a7cdc3ad92a4787ba6fdc33d132f8083de98fc490c03ebc2b39ab8020c41be872b30b3060a2257c33;
    5'b10101 : xpb = 1024'h25ce7e48f917420b150c1fd7f5d024dd5238c451fcf37c971d8f8efdb4cb1ac1dbd52bfe04e0c28d99372d81ca0fcbd60e1b1d7f18a99e21eb3730ea50c12c55f7db13edc38865623bbcdcaba48aa0e5153436afd55627bd3c1db2e55773a5df367eeb77a2ebca8406c094ad0be76f3ca8d73536a03da992c3fcada454d528ce;
    5'b10110 : xpb = 1024'hae37c550d5a948d55b6633861a2b079fd127ab874a1d45ed2987b54b150793ac9fa8d6d3dc14fb7ae92c47810702e255e12424eb58d868ef7cfc4b24e2f0d07fbdcc8628d8b4375e95e5dcfef0141976d0221c07dcd8de40b0ebbcec3eca66962c293547c3a88557aab14ba84f60487766dcc92eccaac7e31b5da5ec90673bd4;
    5'b10111 : xpb = 1024'h85f3c702f04d1ad6d6bacf5d2e2ba310dea08f8bc1cf6ecbb7a32242c2415f8f60340430e922b5d999c322396097e80b50130471765463715e2226013a4dfff80f6ec3b53e4f0c15dd74daafa2c1cdd7970b07c757d567b3702d34f86bf684baf2cbecee339c479dc7e21bc49b08fb88d6087e44a8cc89032c4f23304316e86f;
    5'b11000 : xpb = 1024'h5dafc8b50af0ecd8520f6b34422c3e81ec197390398197aa45be8f3a6f7b2b7220bf318df63070384a59fcf1ba2cedc0bf01e3f793d05df33f4800dd91ab2f7061110141a3e9e0cd2503d860556f82385df3f386d2d1f1262f6ead049922a2dfb96ea494a39009e3e512ebe0e6b1ae9a4534335a84ee4a233d40a073f5c6950a;
    5'b11001 : xpb = 1024'h356bca672594bed9cd64070b562cd9f2f9925794b133c088d3d9fc321cb4f754e14a5eeb033e2a96faf0d7aa13c1f3762df0c37db14c5875206ddbb9e9085ee8b2b33ece0984b5846c92d611081d369924dcdf464dce7a98eeb02510c64ec10480115c3b1383cc2a0243bbfd325a61abb45fe87061100b434e321db7a87641a5;
    5'b11010 : xpb = 1024'hd27cc19403890db48b8a2e26a2d7564070b3b9928e5e96761f56929c9eec337a1d58c48104be4f5ab87b2626d56f92b9cdfa303cec852f70193b69640658e6104557c5a6f1f8a3bb421d3c1bacaeaf9ebc5cb05c8cb040badf19d1cf37adf2946b413e183778e701f748c197e0314bd238b9d863d31cc635f239afb5b25ee40;
    5'b11011 : xpb = 1024'h959113211cca97a58f12b6908e88582685fa22ce760fb2bd6ded8f772a2b3c2265a9371de7801de2fb7ccc61aa4a0fab6fe8aa700ef71dc49358d0d0d295328aca46ee95844b5c380e4ad4150654638ba6b3b05dd04dba8f22bfa723dad19fe03c5e5db1a4344943c3654314c17bedf7e191317e699eeab3b684934396b80146;
    5'b11100 : xpb = 1024'h6d4d14d3376e69a70a675267a288f397937306d2edc1db9bfc08fc6ed76508052634647af48dd841ac13a71a03df1560ded789f62c731846747eabad29f262031be92c21e9e630ef55d9d1c5b90217ec6d9c9c1d4b4a4401e2011f3007fdbe050301155814280b89e09613310d24a10950bce69445c0abd3c77610874967ade1;
    5'b11101 : xpb = 1024'h4509168552123ba885bbee3eb6898f08a0ebead76574047a8a246966849ed3e7e6bf91d8019b92a05caa81d25d741b164dc6697c49ef12c855a48689814f917b6d8b69ae4f8105a69d68cf766bafcc4d348587dcc646cd74a142973c3529dc29c9a3ccfe841bcdcffdc6e34d58cd541abfe89baa21e26cf3d8678dcafc175a7c;
    5'b11110 : xpb = 1024'h1cc518376cb60daa01108a15ca8a2a79ae64cedbdd262d59183fd65e31d89fcaa74abf350ea94cff0d415c8ab70920cbbcb54902676b0d4a36ca6165d8acc0f3bf2da73ab51bda5de4f7cd271e5d80adfb6e739c414356e760840f486255fa4e904684a4f40f90161af7b369a476072c2f1450bffe042e13e9590b0eaec70717;
    5'b11111 : xpb = 1024'ha52e5f3f49481474476a9dc3eee50d3c2d53b6112a4ff6af2437fcab921518b56b1e6a0ae5dd85ec5d367689f3fc374b8fbe506ea799d817c88f7ba06adc651d851f1975ca47ac5a3f20cd7a69e6f93fb65c58f448c60d6ad552194f49acbb0585f0ce7514cc4ae9bee86a64e7eee066ed19e4b82a714c6440ba0356ea591a1d;
    endcase
end

endmodule

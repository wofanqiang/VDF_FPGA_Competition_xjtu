module xpb_5_820
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h4cc2ce3dd76451bbdcbf10e86a91a569db2dd1b2bb25200d3f1e2985c7722aed48d26cbca911f90c98fa27d984d87a6d14c73c806afc82d9155488e039b25cadb9ad45ed90477ce7a088be67bb882d14d5dfddd970d859d5bd1a534e4e15a35a8fb012e6327993b6d1e8aee3bba9936197e41b327e7646b01771897da2d35eb6;
    5'b00010 : xpb = 1024'h99859c7baec8a377b97e21d0d5234ad3b65ba365764a401a7e3c530b8ee455da91a4d9795223f21931f44fb309b0f4da298e7900d5f905b22aa911c07364b95b735a8bdb208ef9cf41117ccf77105a29abbfbbb2e1b0b3ab7a34a69c9c2b46b51f6025cc64f3276da3d15dc7775326c32fc83664fcec8d602ee312fb45a6bd6c;
    5'b00011 : xpb = 1024'h359b2563c43ec06acb37bae22f5aa8ec201371e75bf7bfb03f7dc33ba353d3bfd72ec8bd310f6c972b903845ab2b5e7cda3b8d9b1e42b83f8f5e5b427244a157b8b89d1a01457971cf00389499bcc30d8d9a9ff3c602e07081c267f03016477d8008a688e6a3c296eefa25cc3b2c93fb78d272b52b1776dfffe521745f97b5b7;
    5'b00100 : xpb = 1024'h825df3a19ba31226a7f6cbca99ec4e55fb41439a171cdfbd7e9becc16ac5fead20013579da2165a3c48a601f3003d8e9ef02ca1b893f3b18a4b2e422abf6fe057265e307918cf6596f88f6fc5544f022637a7dcd36db3a463edcbb3e7e2bead80fb8b96f191d564dc0e2d4aff6d6275d10b68de7a98dbd901756aaf2026b146d;
    5'b00101 : xpb = 1024'h1e737c89b1192f19b9b064dbf423ac6e64f9121bfcca5f533fdd5cf17f357c92658b24bdb90ce021be2648b1d17e428c9fafdeb5d188eda609682da4aad6e601b7c3f446724375fbfd77b2c177f159064555620e1b2d670b466a7c921216eba070613a2b9acdf1770c0b9cb4baaf949559c0ca37d7b8a70fe858b96b1c5c0cb8;
    5'b00110 : xpb = 1024'h6b364ac7887d80d5966f75c45eb551d84026e3ceb7ef7f607efb867746a7a77fae5d917a621ed92e5720708b5656bcf9b4771b363c85707f1ebcb684e48942af71713a34028af2e39e0071293379861b1b353fe78c05c0e10384cfe0602c8efb00114d11cd47852dddf44b98765927f6f1a4e56a562eedbfffca42e8bf2f6b6e;
    5'b00111 : xpb = 1024'h74bd3af9df39dc8a8290ed5b8ecaff0a9deb2509d9cfef6403cf6a75b172564f3e780be410a53ac50bc591df7d1269c65242fd084cf230c83720006e3692aabb6cf4b72e34172862bef2cee5625eefefd1024287057eda60b129133f4178fc360b9cdce4ef82057291d139d3a32952f3aaf21ba8459d73fd0cc5161d92063b9;
    5'b01000 : xpb = 1024'h540ea1ed7557ef8484e81fbe237e555a850c840358c21f037f5b202d228950523cb9ed7aea1c4cb8e9b680f77ca9a10979eb6c50efcba5e598c688e71d1b8759707c91607388ef6dcc77eb5611ae1c13d2f00201e130477bc82ce482422d331df069e0b48171b40dfb05c280f5dc2890d2933ced02d01defe83ddadf7bf3c26f;
    5'b01001 : xpb = 1024'ha0d1702b4cbc414061a730a68e0ffac4603a55b613e73f10be7949b2e9fb7b3f858c5a37932e45c582b0a8d101821b768eb2a8d15ac828beae1b11c756cde4072a29d74e03d06c556d00a9bdcd364928a8cfdfdb5208a151854737d09042d6788019f39ab3eb47c4ccee7164b185bbf26a77581f8146649fffaf645d1ec72125;
    5'b01010 : xpb = 1024'h3ce6f91362325e337360c9b7e84758dcc9f22437f994bea67fbab9e2fe6af924cb16497b7219c0437c4c9163a2fc85193f5fbd6ba311db4c12d05b4955adcc036f87e88ce486ebf7faef6582efe2b20c8aaac41c365ace168cd4f924242dd740e0c27457359be2ee18173969755f292ab381946faf714e1fd0b172d638b81970;
    5'b01011 : xpb = 1024'h89a9c7513996afef501fdaa052d8fe46a51ff5eab4b9deb3bed8e368c5dd241213e8b6381b2bb9501546b93d27d4ff865426f9ec0e0e5e252824e4298f6028b129352e7a74ce68df9b7823eaab6adf21608aa1f5a73327ec49ef4c7272437a9b7072873d681576a4e9ffe84d3108bc8c4b65afa22de794cfe822fc53db8b7826;
    5'b01100 : xpb = 1024'h25bf50394f0ccce261d973b1ad105c5f0ed7c46c9a675e49801a5398da4ca1f75972a57bfa1733ce0ee2a1cfc94f692904d40e86565810b28cda2dab8e4010ad6e933fb95584e8822966dfafce174805426586368b8554b1517d0dc6062e7b63d11b07f9e9c611ce3528b051f4e229c4946febf25c127e4fb9250accf57c7071;
    5'b01101 : xpb = 1024'h72821e7726711e9e3e98849a17a201c8ea05961f558c7e56bf387d1ea1becce4a2451238a3292cdaa7dcc9a94e27e396199b4b06c154938ba22eb68bc7f26d5b284085a6e5cc6569c9ef9e17899f751a1845640ffc5dae870e97611454441ebe60cb1ae01c3fa58507115f35b08bbd262c540724da88c4ffd096944a984fcf27;
    5'b01110 : xpb = 1024'he97a75f3be73b9150521dab71d95fe153bd64a13b39fdec8079ed4eb62e4ac9e7cf017c8214a758a178b23befa24d38ca485fa1099e461906e4000dc6d255576d9e96e5c682e50c57de59dcac4bddfdfa204850e0afdb4c16252267e82f1f86c1739b9c9df040ae523a273a74652a5e755e437508b3ae7fa198a2c3b240c772;
    5'b01111 : xpb = 1024'h5b5a759d134b8d4d2d112e93dc6b054b2eeb3653f65f1df9bf9816d47da075b730a16e392b26a0653a72da15747ac7a5df0f9c21749ac8f21c3888ee0084b205274bdcd356ca61f3f867184467d40b12d000262a51883521d33f75b63644c2e15123ae82d069d4652422d61e300ebdc00d425ea78729f52fb90a2c4155142628;
    5'b10000 : xpb = 1024'ha81d43daeaafdf0909d03f7c46fcaab50a190806b1843e06feb6405a4512a0a47973daf5d4389971d36d01eef9534212f3d6d8a1df974bcb318d11ce3a370eb2e0f922c0e711dedb98efd6ac235c3827a5e00403c2608ef79059c904845a663be0d3c16902e3681bf60b8501ebb85121a52679da05a03bdfd07bb5bef7e784de;
    5'b10001 : xpb = 1024'h4432ccc30025fbfc1b89d88da13408cd73d0d6889731bd9cbff7b08a59821e89befdca39b32413efcd08ea819acdabb5a483ed3c27e0fe5896425b503916f6af265733ffc7c85e7e26de92714608a10b87bae844a6b2bbbc97e78a5818456704417c42258494034541344d06af91be59ee30b62a33cb255fa17dc43811d87d29;
    5'b10010 : xpb = 1024'h90f59b00d78a4db7f848e9760bc5ae374efea83b5256dda9ff15da1020f4497707d036f65c360cfc6603125b1fa62622b94b29bc92dd8131ab96e43072c9535ce00479ed580fdb65c76750d90190ce205d9ac61e178b15925501dda6665b0a5ed12c550bb70d96fc131cfbea6b3b51bb8614d15cb2416c0fb8ef4db5b4abdbdf;
    5'b10011 : xpb = 1024'h2d0b23e8ed006aab0a02828765fd0c4fb8b676bd38045d3fc0574a403563c75c4d5a263a3b21877a5f9efaedc1208fc569f83e56db2733bf104c2db271a93b5925628b2c38c65b0855560c9e243d37043f75aa5efbdd42575c8f9ef9fa460b2731d4d5c838be32255e45c3ef2f14bef3cf1f0dace06c558f89f15c2ece9cd42a;
    5'b10100 : xpb = 1024'h79cdf226c464bc66e6c1936fd08eb1b993e4486ff3297d4cff7573c5fcd5f249962c92f6e4338086f89922c745f90a327ebf7ad74623b69825a0b692ab5b9806df0fd119c90dd7eff5decb05dfc56419155588386cb59c2d19a9f248485bae81c184e8ae6b37c5dc302e72d2eabe5255670328df5ee29c3fa162e5ac717032e0;
    5'b10101 : xpb = 1024'h15e37b0ed9dad959f87b2c812ac60fd1fd9c16f1d8d6fce2c0b6e3f61145702edbb6823ac31efb04f2350b59e77373d52f6c8f718e6d69258a560014aa3b8003246de258a9c4579283cd86cb0271ccfcf7306c795107c8f22137b39bdc46af4a222d696aece861057b573ad7ae97bf8db00d652f8d0d85bf7264f4258b612b2b;
    5'b10110 : xpb = 1024'h62a6494cb13f2b15d53a3d699557b53bd8c9e8a493fc1cefffd50d7bd8b79b1c2488eef76c30f4118b2f33336c4bee424433cbf1f969ebfe9faa88f4e3eddcb0de1b28463a0bd47a24564532bdf9fa11cd104a52c1e022c7de5206ea2a5c52a4b1dd7c511f61f4bc4d3fe9bb6a4152ef47f180620b83cc6f89d67da32e3489e1;
    5'b10111 : xpb = 1024'haf69178a88a37cd1b1f94e51ffe95aa5b3f7ba574f213cfd3ef33701a029c6096d5b5bb41542ed1e24295b0cf12468af58fb087264666ed7b4ff11d51da0395e97c86e33ca535161c4df039a79822726a2f0282c32b87c9d9b6c5a387871f5ff418d8f3751db88731f28989f25eae650dfd59b9489fa131fa1480720d107e897;
    5'b11000 : xpb = 1024'h4b7ea0729e1999c4c3b2e7635a20b8be1daf88d934cebc930034a731b49943eeb2e54af7f42e679c1dc5439f929ed25209a81d0cacb0216519b45b571c80215add267f72ab09d10452cdbf5f9c2e900a84cb0c6d170aa962a2fa1b8c0c5cf6c7a2360ff3d38c239c6a5160a3e9c4538928dfd7e4b824fc9f724a1599eaf8e0e2;
    5'b11001 : xpb = 1024'h98416eb0757deb80a071f84bc4b25e27f8dd5a8beff3dca03f52d0b77c0b6edbfbb7b7b49d4060a8b6bf6b7917774cbf1e6f598d17aca43e2f08e43756327e0896d3c5603b514debf3567dc757b6bd1f5aaaea4687e3033860146eda5a729a2231e622da0605b7533c3a0f87a56de6eac0c3f317369b434f89bb9f178dcc3f98;
    5'b11010 : xpb = 1024'h3456f7988af40873b22b915d1ee9bc406295290dd5a15c36009440e7907aecc14141a6f87c2bdb26b05b540bb8f1b661cf1c6e275ff656cb93be2db955126604dc31d69f1c07cd8e8145398c7a6326033c85ce876c352ffd67a2302dee5d9aea928ea39687b6527c8762d78c6947542309ce2f6764c62ccf5abdad90a7bd37e3;
    5'b11011 : xpb = 1024'h8119c5d662585a2f8eeaa245897b61aa3dc2fac090c67c433fb26a6d57ed17ae8a1413b5253dd43349557be53dca30cee3e3aaa7caf2d9a4a912b6998ec4c2b295df1c8cac4f4a7621cdf7f435eb53181265ac60dd0d89d324bc837c3c733e45223eb67cba2fe633594b867024f0e784a1b24a99e33c737f722f370e4a909699;
    5'b11100 : xpb = 1024'h1d2f4ebe77ce7722a0a43b56e3b2bfc2a77ac9427673fbd900f3da9d6c5c9593cf9e02f904294eb142f16477df449a719490bf42133c8c320dc8001b8da4aaaedb3d2dcb8d05ca18afbcb3b95897bbfbf44090a1c15fb6982c4a44cfd05e3f0d82e737393be0815ca4744e74e8ca54bceabc86ea11675cff4331458764818ee4;
    5'b11101 : xpb = 1024'h69f21cfc4f32c8de7d634c3f4e44652c82a89af531991be64012042333cec08118706fb5ad3b47bddbeb8c51641d14dea957fbc27e390f0b231c88fbc757075c94ea73b91d4d470050457221141fe910ca206e7b3238106de964981e1e73e26812974a1f6e5a1513765cfd58a473e81e82a0a21c8fdda3af5aa2cf050754ed9a;
    5'b11110 : xpb = 1024'h607a5e464a8e5d18f1ce550a87bc344ec60697717469b7c01537453483e3e665dfa5ef98c26c23bd58774e405977e815a05105cc682c19887d1d27dc636ef58da4884f7fe03c6a2de342de636cc51f4abfb52bc168a3d32f0f25971b25ee330733fcadbf00ab03cc185c55d684d5556cbaade6cbe088d2f2ba4dd7e2145e5e5;
    5'b11111 : xpb = 1024'h52ca74223c0d378d6bdbf639130d68aec78e3b29d26bbb8940719dd90fb06953a6cccbb63538bb486e819cbd8a6ff8ee6ecc4cdd317f44719d265b5dffe94c0693f5cae58e4b438a7ebcec4df2547f0981db309587629708ae0cacc00074868b02efddc2228443f3936e744123f6e8b8638ef99f3c7ed3df431666fbc419449b;
    endcase
end

endmodule

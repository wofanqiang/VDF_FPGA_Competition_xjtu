module xpb_5_890
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h76ce70b7605ce3e2f3a80a002a70481fec8c2c41c8412d07c3c01364c0835fc988cb772ca8611e5002e1855539eadfbeed02ba80c73f02a4a304503409df0e63d055a23cd8643ed6d29c5cb6965178bc15eb11fac84c55a3d20c7115765ae08fa2a3bb54ba83c8d1ee03a6bf09f2e1e69e290a3a078eda12cd05000a169165e5;
    5'b00010 : xpb = 1024'h3cef9c18fecb92fd1c4a9c29448648ee67a25552bb0ab99809a36d73ce04128b0e4e70e0869bbe116664cb639077aeb375eb4d1b6bcb34fd95696109d8eba8162c5c0fcb01378068929eb6ca93c72d4737d12a5d04127e36ee8c5030328b1e8d163fe47fc43e99165547669f1c159da3ed783591bed256f5539a850fa440655f;
    5'b00011 : xpb = 1024'h310c77a9d3a421744ed2e525e9c49bce2b87e63add446284f86c782db84c54c93d16a9464d65dd2c9e81171e7047da7fed3dfb61057675687ce71dfa7f841c888627d592a0ac1fa52a110de913ce1d259b742bf3fd8a6ca0b0c2f4aeebb5c8a89dc0daacdf9695abc8b267f2e3859613cc760e97615d3d7da300a1531ef64d9;
    5'b00100 : xpb = 1024'h79df3831fd9725fa38953852890c91dccf44aaa5761573301346dae79c0825161c9ce1c10d377c22ccc996c720ef5d66ebd69a36d79669fb2ad2c213b1d7502c58b81f96026f00d1253d6d95278e5a8e6fa254ba0824fc6ddd18a06065163d1a2c7fc8ff887d322caa8ecd3e382b3b47daf06b237da4adeaa7350a1f4880cabe;
    5'b00101 : xpb = 1024'h400063939c05d5146137ca7ba32292ab4a5ad3b668deffc0592a34f6a988d7d7a21fdb74eb721be4304cdcd5777c2c5b74bf2cd17c229c541d37d2e980e3e9deb4be8d242b424262e53fc7a925040f1991886d1c43eb2500f9987f7b21467b17a01bf22a9238027111d28d1e4a4df7052a3f967b34e82acd2dca8f24d62fca38;
    5'b00110 : xpb = 1024'h6218ef53a74842e89da5ca4bd389379c570fcc75ba88c509f0d8f05b7098a9927a2d528c9acbba593d022e3ce08fb4ffda7bf6c20aecead0f9ce3bf4ff0839110c4fab2541583f4a54221bd2279c3a4b36e857e7fb14d9416185e95dd76b91513b81b559bf2d2b579164cfe5c70b2c2798ec1d2ec2ba7afb460142a63dec9b2;
    5'b00111 : xpb = 1024'h7cefffac9ad168117d8266a4e7a8db99b1fd290923e9b95862cda26a778cea62b06e4c55720dd9f596b1a83907f3db0eeaaa79ece7edd151b2a133f359cf91f4e11a9cef2c79c2cb77de7e73b8cb3c60c959977947fda337e824cfab53d199a4b65bd6aa56769b876719f3bd666394a917b7cc0cf3ba81c2816514347a702f97;
    5'b01000 : xpb = 1024'h43112b0e3940172ba624f8ce01bedc682d13521a16b345e8a8b0fc79850d9d2435f14609504879b6fa34ee475e80aa0373930c878c7a03aaa50644c928dc2ba73d210a7d554d045d37e0d887b640f0ebeb3fafdb83c3cbcb04a4aec61001d7a229f7ffd560316bcbce5db39d788650666706f764aafdfea507fa993a081f2f11;
    5'b01001 : xpb = 1024'h932566fd7aec645cec78af71bd4dd36a8297b2b097cd278ee945688928e4fe5bb743fbd2e8319785db83455b50d78f7fc7b9f2231063603976b559ef7e8c5599927780b7e2045eef7e3329bb3b6a5770d25c83dbf89f45e21248de0cc32159f9d94290069ec3c1035a1737d8aa90c23b65622bc62417b878e901e3f95ce2e8b;
    5'b01010 : xpb = 1024'h8000c727380baa28c26f94f74645255694b5a76cd1bdff80b25469ed5311afaf443fb6e9d6e437c86099b9aaeef858b6e97e59a2f84538a83a6fa5d301c7d3bd697d1a48568484c5ca7f8f524a081e332310da3887d64a01f330fef6428cf62f4037e455247004e223a51a3c949bee0a547f2cf669d0559a5b951e49ac5f9470;
    5'b01011 : xpb = 1024'h4621f288d67a5942eb122720605b26250fcbd07dc4878c10f837c3fc60926270c9c2b09db51ed789c41cffb9458527ab7266ec3d9cd16b012cd4b6a8d0d46d6fc58387d67f57c6578a81e966477dd2be44f6f29ac39c72950fb0de10febd342cb3d40d802e2ad5268ae8da1ca6bea9c7a3ce584e2113d27ce22aa34f3a0e93ea;
    5'b01100 : xpb = 1024'hc431dea74e9085d13b4b9497a7126f38ae1f98eb75118a13e1b1e0b6e1315324f45aa519359774b27a045c79c11f69ffb4f7ed8415d9d5a1f39c77e9fe107222189f564a82b07e94a84437a44f3874966dd0afcff629b282c30bd2bbaed722a277036ab37e5a56af22c99fcb8e16584f31d83a5d8574f5f68c02854c7bd9364;
    5'b01101 : xpb = 1024'h83118ea1d545ec40075cc349a4e16f13776e25d07f9245a901db31702e9674fbd811217e3bba959b2a81cb1cd5fcd65ee8523959089c9ffec23e17b2a9c01585f1df97a1808f46c01d20a030db4500057cc81cf7c7aef0cbfe3d2e41314852b9ca13f1fff2696e3ce03040bbc2d4476b91468ddfdfe6297235c5285ede4ef949;
    5'b01110 : xpb = 1024'h4932ba0373b49b5a2fff5572bef76fe1f2844ee1725bd23947be8b7f3c1727bd5d941b3219f5355c8e05112b2c89a553713acbf3ad28d257b4a3288878ccaf384de6052fa9628851dd22fa44d8bab4909eae355a0375195f1abd0d5bed7890b73db01b2afc243e814774009bd4f70328e095b9379729a654bc5aad646bfdf8c3;
    5'b01111 : xpb = 1024'hf53e56512234a7458a1e79bd90d70b06d9a77f265255ec98da1e58e4997da7ee31714e5f82fd51df188573983167447fa235e8e51b504b0a708395e47d948eaa9ec72bdd235c9e39d255458d630691bc0944dbc3f3b41f2373cec76a9a8ceb4b14c445605df0ec5aeb7c07be719bee62fe4e48f4e6d233742f03269f9acf83d;
    5'b10000 : xpb = 1024'h8622561c72802e574c49f19c037db8d05a26a4342d668bd15161f8f30a1b3a486be28c12a090f36df469dc8ebd015406e726190f18f407554a0c899251b8574e7a4214faaa9a08ba6fc1b10f6c81e1d7d67f5fb70787979609495d8c2003af4453efffaac062d7979cbb673af10ca0ccce0deec955fbfd4a0ff53274103e5e22;
    5'b10001 : xpb = 1024'h4c43817e10eedd7174ec83c51d93b99ed53ccd452030186197455302179bed09f16585c67ecb932f57ed229d138e22fb700eaba9bd8039ae3c719a6820c4f100d6488288d36d4a4c2fc40b2369f79662f8657819434dc02925c93ca6dc33ed41c78c28d5ca1da7dc03ff271b032f5c8a1d5d1a210d3f7a2c968ab7799ded5d9c;
    5'b10010 : xpb = 1024'h1264acdfaf5d8c8b9d8f15ee37a9ba6d5052f65612f9a4f1dd28ad11251c9fcb76e87f7a5d0632f0bb7068ab6a1af1eff8f73e44620c6c072ed6ab3defd18ab3324ef016fc408bddefc66537676d4aee1a4b907b7f13e8bc42491bc198642b3f3b285200d3d878206b42e6fb155218476cac4578c482f70f1d203c7f2b9c5d16;
    5'b10011 : xpb = 1024'h89331d970fba706e91371fee621a028d3cdf2297db3ad1f9a0e8c075e59fff94ffb3f6a705675140be51ee00a405d1aee5f9f8c5294b6eabd1dafb71f9b0991702a49253d4a4cab4c262c1edfdbec3aa3036a27647603e6014558cd70ebf0bceddcc0d558e5c40f259468dba1f44fa2e0ad54fb2cc11d121ea253c89422dc2fb;
    5'b10100 : xpb = 1024'h4f5448f8ae291f88b9d9b2177c30035bb7f54ba8ce045e89e6cc1a84f320b2568536f05ae3a1f10221d5340efa92a0a36ee28b5fcdd7a104c4400c47c8bd32c95eaaffe1fd780c4682651c01fb347835521cbad8832666f330d56bf1caef49cc5168368098171136c08a4d9a3167b5eb5a247b0a83554e0470bac18ecfdcc275;
    5'b10101 : xpb = 1024'h1575745a4c97cea2e27c44409646042a330b74b9c0cdeb1a2caf749400a165180ab9ea0ec1dc90c385587a1d511f6f97f7cb1dfa7263d35db6a51d1d97c9cc7bbab16d70264b4dd842677615f8aa2cc07402d33abeec8f864d554b0c871f87c9c5045faba1d1e17b27ce0d7a438a71a8a973a6623a98cae6f75046945d8bc1ef;
    5'b10110 : xpb = 1024'h8c43e511acf4b285d6244e40c0b64c4a1f97a0fb890f1821f06f87f8c124c4e19385613b6a3daf138839ff728b0a4f56e4cdd87b39a2d60259a96d51a1a8dadf8b070facfeaf8caf1503d2cc8efba57c89ede5358738e52a1f61bc21fd7a685967a81b005c55aa4d15d1b4394d7d538f479cb09c4227a4f9c455469e741d27d4;
    5'b10111 : xpb = 1024'h526510734b63619ffec6e069dacc4d189aadca0c7bd8a4b23652e207cea577a319085aef48784ed4ebbd4580e1971e4b6db66b15de2f085b4c0e7e2770b57491e70d7d3b2782ce40d5062ce08c715a07abd3fd97c2ff0dbd3be19b3cb9aaa656db44442b66107a917d1574195fa00f4c96ebdbf3f96b21dc4aeacba401cc274e;
    5'b11000 : xpb = 1024'h18863bd4e9d210ba27697292f4e24de715c3f31d6ea231427c363c16dc262a649e8b54a326b2ee964f408b8f3823ed3ff69efdb082bb3ab43e738efd3fc20e444313eac950560fd2950886f489e70e92cdba15f9fec5365058617a5775dae4544ee06d566fcb4ad5e45933f971c2cb09e63b074bb0ae9ebed18050a98f7b26c8;
    5'b11001 : xpb = 1024'h8f54ac8c4a2ef49d1b117c931f52960702501f5f36e35e4a3ff64f7b9ca98a2e2756cbcfcf140ce6522210e4720eccfee3a1b83149fa3d58e177df3149a11ca813698d0628ba4ea967a4e3ab2038874ee3a527f4c7118bf42a6deb6cec35c4e3f18428ab2a4f13a7d25cdab87bb5acf084641185b83d78d19e8550b3a60c8cad;
    5'b11010 : xpb = 1024'h5575d7ede89da3b743b40ebc396896d57d66487029aceada85d9a98aaa2a3cefacd9c583ad4eaca7b5a556f2c89b9bf36c8a4acbee866fb1d3dcf00718adb65a6f6ffa94518d903b27a73dbf1dae3bda058b405702d7b48746edca87a86602e1652051d63409e3ec39a09a988dd868add3b33cdd6f80f5b4251ad5b933bb8c27;
    5'b11011 : xpb = 1024'h1b97034f870c52d16c56a0e5537e97a3f87c71811c76776acbbd0399b7aaefb1325cbf378b894c6919289d011f286ae7f572dd669312a20ac64200dce7ba500ccb7668227a60d1cce7a997d31b23f065277158b93e9ddd1a636da9a2649640ded8bc7b013dc4b430a0e45a789ffb246b2302683526c47296abb05abec16a8ba1;
    5'b11100 : xpb = 1024'h92657406e76936b45ffeaae57deedfc3e5089dc2e4b7a4728f7d16fe782e4f7abb28366433ea6ab91c0a225659134aa6e27597e75a51a4af69465110f1995e709bcc0a5f52c510a3ba45f489b17569213d5c6ab406ea32be357a1ab7daf1216e7b603655f8487d028ee80137a9ee0651c12b726f2e534ca978b55ac8d7fbf186;
    5'b11101 : xpb = 1024'h58869f6885d7e5ce88a13d0e9804e092601ec6d3d7813102d560710d85af023c40ab301812250a7a7f8d6864afa0199b6b5e2a81feddd7085bab61e6c0a5f822f7d277ed7b9852357a484e9daeeb1dac5f42831642b05b5151f9f9d297215f6beefc5f8102034d46f62bc117bc10c20f107a9dc6e596c98bff4adfce65aaf100;
    5'b11110 : xpb = 1024'h1ea7caca244694e8b143cf37b21ae160db34efe4ca4abd931b43cb1c932fb4fdc62e29cbf05faa3be310ae73062ce88ff446bd1ca36a09614e1072bc8fb291d553d8e57ba46b93c73a4aa8b1ac60d23781289b787e7683e46e79d8ed53519d69629888ac0bbe1d8b5d6f80f7ce337dcc5fc9c91e9cda466e85e064d3f359f07a;
    5'b11111 : xpb = 1024'h95763b8184a378cba4ebd937dc8b2980c7c11c26928bea9adf03de8153b314c74ef9a0f898c0c88be5f233c84017c84ee149779d6aa90c05f114c2f09991a039242e87b87ccfd29e0ce7056842b24af39713ad7346c2d98840864a02c9ac7df9053c4400c641e65d4b7327b6d8265fb2fdf2d358a469208152e564de09eb565f;
    endcase
end

endmodule

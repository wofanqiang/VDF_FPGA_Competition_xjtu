module xpb_5_545
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h421865244a32a4e143a4a0dfa3b7d34732f1989a76551b69f192d88ceb89bbf559b64d24159ddb5d8cd6a8fbf30b1994dba825ab64eaa6e0360aa2f982e60bac4ddc698529ee63e2dd08f8976f9c773300956d5047f0cad22b1b817b2059ec4d79755ad6f127c5b489e8999dc1594fc5f34464e802cf3650840d05ab3e7749b6;
    5'b00010 : xpb = 1024'h8430ca48946549c2874941bf476fa68e65e33134ecaa36d3e325b119d71377eab36c9a482b3bb6bb19ad51f7e6163329b7504b56c9d54dc06c1545f305cc17589bb8d30a53dcc7c5ba11f12edf38ee66012adaa08fe195a4563702f640b3d89af2eab5ade24f8b6913d1333b82b29f8be688c9d0059e6ca1081a0b567cee936c;
    5'b00011 : xpb = 1024'h159bea171ca9b9daffe86ac7dacd3284275ec69e8d87b1c656dbd0510f9a86d809da69f376b3138a0725bbacf5c33bf42ede491c0c0d2454f180a98e4ddfae53754607e0ce3a2e638480e723b5f9a1680dbb4e584b4c3365cbc5f276a6e322563d587e5b22ae589016f9e5fa4c3bc9288af34fd5b82245c145b795fd328376b7;
    5'b00100 : xpb = 1024'h57b44f3b66dc5ebc438d0ba77e8505cb5a505f3903dccd30486ea8ddfb2442cd6390b7178c50eee793fc64a8e8ce55890a866ec770f7cb35278b4c87d0c5b9ffc3227165f82892466189dfbb2596189b0e50bba8933cfe37f6e173f1c73d0ea3b6cdd93213d61e44a0e27f980d9518ee7e37b4bdbaf17c11c9c49ba870fac06d;
    5'b00101 : xpb = 1024'h99ccb45fb10f039d8731ac87223cd9128d41f7d37a31e89a3a01816ae6adfec2bd47043ba1eeca4520d30da4dbd96f1de62e9472d5e272155d95ef8153abc5ac10fedaeb2216f6293e92d85295328fce0ee628f8db2dc90a21fcf56ce796faf13043340904fde3f92acb1935ceee68b4717c19a5bdc0b2624dd1a153af720a23;
    5'b00110 : xpb = 1024'h2b37d42e395373b5ffd0d58fb59a65084ebd8d3d1b0f638cadb7a0a21f350db013b4d3e6ed6627140e4b7759eb8677e85dbc9238181a48a9e301531c9bbf5ca6ea8c0fc19c745cc70901ce476bf342d01b769cb0969866cb978be4ed4dc644ac7ab0fcb6455cb1202df3cbf49877925115e69fab70448b828b6f2bfa6506ed6e;
    5'b00111 : xpb = 1024'h6d503952838618974375766f5952384f81af25d791647ef69f4a792f0abec9a56d6b210b030402719b222055de91917d3964b7e37d04ef8a190bf6161ea5685338687946c662c0a9e60ac6dedb8fba031c0c0a00de89319dc2a766686e2030f9f426578d368476d4b7dc659259d0e217092b04937313c1d30f7c31a5a37e3724;
    5'b01000 : xpb = 1024'haf689e76cdb8bd78871a174efd0a0b96b4a0be7207b99a6090dd51bbf648859ac7216e2f18a1ddcf27f8c951d19cab12150cdd8ee1ef966a4f16990fa18b73ff8644e2cbf051248cc313bf764b2c31361ca177512679fc6fedc2e7e38e7a1d476d9bb26427ac3c8941c4ff301b2a31dcfc6f697b75e2f82393893750e1f580da;
    5'b01001 : xpb = 1024'h40d3be4555fd2d90ffb940579067978c761c53dba8971553049370f32ecf94881d8f3dda64193a9e15713306e149b3dc8c9adb5424276cfed481fcaae99f0afa5fd217a26aae8b2a8d82b56b21ece4382931eb08e1e49a316351d763f4a96702b8097b11680b09b044edb1eee4b35b79a0d9ef812866d143d126c1f7978a6425;
    5'b01010 : xpb = 1024'h82ec2369a02fd272435de137341f6ad3a90dec761eec30bcf62649801a59507d77458afe79b715fba247dc02d454cd71684300ff891213df0a8c9fa46c8516a6adae8127949cef0d6a8bae0291895b6b29c7585929d565038e6d58df15035350317ed5e85932cf64ced64b8ca60cab3f941e54692b3607945533c7a2d601addb;
    5'b01011 : xpb = 1024'h145743382874428abbfd0a3fc77cf6c96a8981dfbfc9abaf69dc68b752e05f6acdb35aa9c52e72ca8fc045b7e401d63bdfd0fec4cb49ea738ff8033fb498ada1873bb5fe0efa55ab34faa3f7684a0e6d3657cc10e54002c503fc485f7b329d0b7bec9e9599919c8bd1fefe4b6f95d4dc3888da6eddb9e0b492d152498b969126;
    5'b01100 : xpb = 1024'h566fa85c72a6e76bffa1ab1f6b34ca109d7b1a7a361ec7195b6f41443e6a1b602769a7cddacc4e281c96eeb3d70cefd0bb79247030349153c602a639377eb94dd5181f8338e8b98e12039c8ed7e685a036ed39612d30cd972f17c9da9b8c8958f561f96c8ab962405be797e930ef24a22bcd3f56e089170516de57f4ca0ddadc;
    5'b01101 : xpb = 1024'h98880d80bcd98c4d43464bff0eec9d57d06cb314ac73e2834d0219d129f3d755811ff4f1f06a2985a96d97afca18096597214a1b951f3833fc0d4932ba64c4fa22f4890862d71d70ef0c95264782fcd33782a6b1752198695a334b55bbe675a66ed754437be127f4e5d03186f24874681f11a43ee3584d559aeb5da008852492;
    5'b01110 : xpb = 1024'h29f32d4f451dfc65bbe57507a24a294d91e8487e4d515d75c0b83908627ae642d78dc49d3be1865496e60164d9c512300eaf47e0d7570ec88178acce02785bf4fc81bddedd34840eb97b8b1b1e43afd544131a69308c362acfc23ad62215bf61b9451cf0bc3ff51be8f8e445bbd19e04c37c2a4495dc2675d888e846be1a07dd;
    5'b01111 : xpb = 1024'h6c0b92738f50a146ff8a15e74601fc94c4d9e118c3a678dfb24b11954e04a238314411c1517f61b223bcaa60ccd02bc4ea576d8c3c41b5a8b7834fc7855e67a14a5e27640722e7f1968483b28de0270844a887b9787d00fcfaddbc51426fabaf32ba77c7ad67bad072e17de37d2aedcab6c08f2c98ab5cc65c95edf1fc915193;
    5'b10000 : xpb = 1024'hae23f797d9834628432eb6c6e9b9cfdbf7cb79b339fb9449a3ddea22398e5e2d8afa5ee5671d3d0fb093535cbfdb4559c5ff9337a12c5c88ed8df2c10844734d983a90e931114bd4738d7c49fd7c9e3b453df509c06dcbcf25f93dcc62c997fcac2fd29e9e8f8084fcca17813e843d90aa04f4149b7a9316e0a2f39d3b089b49;
    5'b10001 : xpb = 1024'h3f8f176661c7b640bbcddfcf7d175bd1b9470f1cdad90f3c1794095972156d1ae1682e90b29499de9e0bbd11cf884e243d8d90fce364331d72f9565c50580a4871c7c5bfab6eb2723dfc723ed43d513d51ce68c17bd869909b882d4cc8f8e1b7f69d9b4bdeee4dabfff2ca40080d672d4e6f7a1a4dfe6c371e407e43f09d7e94;
    5'b10010 : xpb = 1024'h81a77c8aabfa5b21ff7280af20cf2f18ec38a7b7512e2aa60926e1e65d9f29103b1e7bb4c832753c2ae2660dc29367b91935b6a8484ed9fda903f955d33e15f4bfa42f44d55d16551b056ad643d9c8705263d611c3c93462c6a3aec7e952ce057012f622d016136089db63ddc966b6f341b3df0250cda287a24d83ef2f14c84a;
    5'b10011 : xpb = 1024'h13129c59343ecb3a7811a9b7b42cbb0eadb43d20f20ba5987cdd011d962637fd918c4b6013a9d20b185acfc2d240708390c3b46d8a86b0922e6f5cf11b51acef9931641b4fba7cf2e57460cb1a9a7b725ef449c97f33d2243c329e484f8217c0ba80bed01074e0878d04169c92efe08fe61e650803517ba7dfeb0e95e4a9ab95;
    5'b10100 : xpb = 1024'h552b017d7e71701bbbb64a9757e48e55e0a5d5bb6860c1026e6fd9aa81aff3f2eb4298842947ad68a53178bec54b8a186c6bda18ef7157726479ffea9e37b89be70dcda079a8e0d5c27d59628a36f2a55f89b719c7249cf6674e1fc36fdc040e33f619a7019ca63c16ecb03a54493055d962c9f00620b1f863f814412320f54b;
    5'b10101 : xpb = 1024'h974366a1c8a414fcff5aeb76fb9c619d13976e55deb5dc6c6002b2376d39afe844f8e5a83ee588c6320821bab856a3ad4813ffc4545bfe529a84a2e4211dc44834ea3725a39744b89f8651f9f9d369d8601f246a0f1567c89269a13e9035f05bad6b747df2c46bf0a0d549d815a2801bcca72ed808efe848e80519ec61983f01;
    5'b10110 : xpb = 1024'h28ae867050e8851577fa147f8ef9ed92d51303bf7f93575ed3b8d16ea5c0bed59b66b5538a5ce5951f808b6fc803ac77bfa1fd899693d4e71ff0067f69315b430e776bfc1df4ab5669f547eed0941cda6caf9821ca80058a07f890bef6653a16f7d93d2b33233917a3fdfc96df2ba9b87111b4ddbb73c16925a2a493172d224c;
    5'b10111 : xpb = 1024'h6ac6eb949b1b29f6bb9eb55f32b1c0da08049c59f5e872c8c54ba9fb914a7acaf51d02779ffac0f2ac57346bbb0ec60c9b4a2334fb7e7bc755faa978ec1766ef5c53d58147e30f3946fe40864030940d6d4505721270d05c3314123a16bf2664714e9802244afecc2de69634a084f97e645619c5be42f7b9a9afaa3e55a46c02;
    5'b11000 : xpb = 1024'hacdf50b8e54dced7ff43563ed66994213af634f46c3d8e32b6de82887cd436c04ed34f9bb5989c50392ddd67ae19dfa176f248e0606922a78c054c726efd729baa303f0671d1731c2407391dafcd0b406dda72c25a619b2e5e2f93b5371912b1eac3f2d91572c480b7cf2fd261de4944579a7eadc1122e0a2dbcafe9941bb5b8;
    5'b11001 : xpb = 1024'h3e4a70876d923ef077e27f4769c72016fc71ca5e0d1b09252a94a1bfb55b45ada5411f47010ff91f26a6471cbdc6e86bee8046a5a2a0f93c1170b00db711099683bd73dcec2ed9b9ee762f12868dbe427a6ae67a15cc38efd3be83359d485c6d3531bb8655d191a7baf7e2912b6772e0fc0504b37396072a6b5a3a9049b09903;
    5'b11010 : xpb = 1024'h8062d5abb7c4e3d1bb8720270d7ef35e2f6362f88370248f1c277a4ca0e501a2fef76c6b16add47cb37cf018b0d20200ca286c51078ba01c477b530739f71542d199dd62161d3d9ccb7f27a9f62a35757b0053ca5dbd03c1feda04b0bda248baaea7165d46f9575c44e07c2eecc0c2a6ef49699b76653d7aef67403b8827e2b9;
    5'b11011 : xpb = 1024'h11cdf57a400953ea3426492fa0dc7f53f0def862244d9f818fdd9983d96c109055653c166225314ba0f559cdc07f0acb41b66a1649c376b0cce6b6a2820aac3dab271238907aa43a95ee1d9ecceae8778790c7821927a1837468f43123d19275f914df0a8758248348092eedb649ec4393b3efa128e9169b2d04cae23dbcc604;
    5'b11100 : xpb = 1024'h53e65a9e8a3bf8cb77caea0f4494529b23d090fc9aa2baeb81707210c4f5cc85af1b893a77c30ca92dcc02c9b38a24601d5e8fc1aeae1d9102f1599c04f0b7e9f9037bbdba69081d72f716363c875faa882634d261186c559f8475ac442b7ec3728a39e1787fea37d1f1c88b77a33c0986f854892bb84cebb111d08d7c340fba;
    5'b11101 : xpb = 1024'h95febfc2d46e9dacbb6f8aeee84c25e256c2299710f7d65573034a9db07f887b08d1d65e8d60e806baa2abc5a6953df4f906b56d1398c47138fbfc9587d6c39646dfe542e4576c0050000ecdac23d6dd88bba222a9093727ca9ff72764856b10ebff94b869a7afec5bda622938fc8bcf7a3cb9712e87833c351ed638baab5970;
    5'b11110 : xpb = 1024'h2769df915cb30dc5340eb3f77ba9b1d8183dbf00b1d55147e6b969d4e90697685f3fa609d8d844d5a81b157ab64246bf7094b33255d09b05be676030cfea5a91206d1a195eb4d29e1a6f04c282e489df954c15da6473d4e9402ee6a7cab4b4cc366d5d65aa067d135f0314e80285b56c1ea73f76e10b5c5c72bc60df70403cbb;
    5'b11111 : xpb = 1024'h698244b5a6e5b2a677b354d71f61851f4b2f579b282a6cb1d84c4261d490535db8f5f32dee76203334f1be76a94d60544c3cd8ddbabb41e5f472032a52d0663d6e49839e88a33680f777fd59f281011295e1832aac649fbb6b4a6822eb0ea119afe2b83c9b2e42c7e8ebae85c3df053211eba45ee3da92acf6c9668aaeb78671;
    endcase
end

endmodule

module alu
(
    input clk,
    input rst,   //needing a clear signal "clear_reg", usage: .rst(rst_sys & clear_reg)
    input [127:0] col_in_0,
    input [127:0] col_in_1,
    input [127:0] col_in_2,
    input [127:0] col_in_3,
    input [127:0] col_in_4,
    input [127:0] col_in_5,
    input [127:0] col_in_6,
    input [127:0] col_in_7,
    input [127:0] col_in_8,
    input [127:0] col_in_9,
    input [127:0] col_in_10,
    input [127:0] col_in_11,
    input [127:0] col_in_12,
    input [127:0] col_in_13,
    input [127:0] col_in_14,
    input [127:0] col_in_15,
    input [127:0] col_in_16,
    input [127:0] col_in_17,
    input [127:0] col_in_18,
    input [127:0] col_in_19,
    input [127:0] col_in_20,
    input [127:0] col_in_21,
    input [127:0] col_in_22,
    input [127:0] col_in_23,
    input [127:0] col_in_24,
    input [127:0] col_in_25,
    input [127:0] col_in_26,
    input [127:0] col_in_27,
    input [127:0] col_in_28,
    input [127:0] col_in_29,
    input [127:0] col_in_30,
    input [127:0] col_in_31,
    input [127:0] col_in_32,
    input [127:0] col_in_33,
    input [127:0] col_in_34,
    input [127:0] col_in_35,
    input [127:0] col_in_36,
    input [127:0] col_in_37,
    input [127:0] col_in_38,
    input [127:0] col_in_39,
    input [127:0] col_in_40,
    input [127:0] col_in_41,
    input [127:0] col_in_42,
    input [127:0] col_in_43,
    input [127:0] col_in_44,
    input [127:0] col_in_45,
    input [127:0] col_in_46,
    input [127:0] col_in_47,
    input [127:0] col_in_48,
    input [127:0] col_in_49,
    input [127:0] col_in_50,
    input [127:0] col_in_51,
    input [127:0] col_in_52,
    input [127:0] col_in_53,
    input [127:0] col_in_54,
    input [127:0] col_in_55,
    input [127:0] col_in_56,
    input [127:0] col_in_57,
    input [127:0] col_in_58,
    input [127:0] col_in_59,
    input [127:0] col_in_60,
    input [127:0] col_in_61,
    input [127:0] col_in_62,
    input [127:0] col_in_63,
    input [127:0] col_in_64,
    input [127:0] col_in_65,
    input [127:0] col_in_66,
    input [127:0] col_in_67,
    input [127:0] col_in_68,
    input [127:0] col_in_69,
    input [127:0] col_in_70,
    input [127:0] col_in_71,
    input [127:0] col_in_72,
    input [127:0] col_in_73,
    input [127:0] col_in_74,
    input [127:0] col_in_75,
    input [127:0] col_in_76,
    input [127:0] col_in_77,
    input [127:0] col_in_78,
    input [127:0] col_in_79,
    input [127:0] col_in_80,
    input [127:0] col_in_81,
    input [127:0] col_in_82,
    input [127:0] col_in_83,
    input [127:0] col_in_84,
    input [127:0] col_in_85,
    input [127:0] col_in_86,
    input [127:0] col_in_87,
    input [127:0] col_in_88,
    input [127:0] col_in_89,
    input [127:0] col_in_90,
    input [127:0] col_in_91,
    input [127:0] col_in_92,
    input [127:0] col_in_93,
    input [127:0] col_in_94,
    input [127:0] col_in_95,
    input [127:0] col_in_96,
    input [127:0] col_in_97,
    input [127:0] col_in_98,
    input [127:0] col_in_99,
    input [127:0] col_in_100,
    input [127:0] col_in_101,
    input [127:0] col_in_102,
    input [127:0] col_in_103,
    input [127:0] col_in_104,
    input [127:0] col_in_105,
    input [127:0] col_in_106,
    input [127:0] col_in_107,
    input [127:0] col_in_108,
    input [127:0] col_in_109,
    input [127:0] col_in_110,
    input [127:0] col_in_111,
    input [127:0] col_in_112,
    input [127:0] col_in_113,
    input [127:0] col_in_114,
    input [127:0] col_in_115,
    input [127:0] col_in_116,
    input [127:0] col_in_117,
    input [127:0] col_in_118,
    input [127:0] col_in_119,
    input [127:0] col_in_120,
    input [127:0] col_in_121,
    input [127:0] col_in_122,
    input [127:0] col_in_123,
    input [127:0] col_in_124,
    input [127:0] col_in_125,
    input [127:0] col_in_126,
    input [127:0] col_in_127,
    input [127:0] col_in_128,
    input [127:0] col_in_129,
    input [127:0] col_in_130,
    input [127:0] col_in_131,
    input [127:0] col_in_132,
    input [127:0] col_in_133,
    input [127:0] col_in_134,
    input [127:0] col_in_135,
    input [127:0] col_in_136,
    input [127:0] col_in_137,
    input [127:0] col_in_138,
    input [127:0] col_in_139,
    input [127:0] col_in_140,
    input [127:0] col_in_141,
    input [127:0] col_in_142,
    input [127:0] col_in_143,
    input [127:0] col_in_144,
    input [127:0] col_in_145,
    input [127:0] col_in_146,
    input [127:0] col_in_147,
    input [127:0] col_in_148,
    input [127:0] col_in_149,
    input [127:0] col_in_150,
    input [127:0] col_in_151,
    input [127:0] col_in_152,
    input [127:0] col_in_153,
    input [127:0] col_in_154,
    input [127:0] col_in_155,
    input [127:0] col_in_156,
    input [127:0] col_in_157,
    input [127:0] col_in_158,
    input [127:0] col_in_159,
    input [127:0] col_in_160,
    input [127:0] col_in_161,
    input [127:0] col_in_162,
    input [127:0] col_in_163,
    input [127:0] col_in_164,
    input [127:0] col_in_165,
    input [127:0] col_in_166,
    input [127:0] col_in_167,
    input [127:0] col_in_168,
    input [127:0] col_in_169,
    input [127:0] col_in_170,
    input [127:0] col_in_171,
    input [127:0] col_in_172,
    input [127:0] col_in_173,
    input [127:0] col_in_174,
    input [127:0] col_in_175,
    input [127:0] col_in_176,
    input [127:0] col_in_177,
    input [127:0] col_in_178,
    input [127:0] col_in_179,
    input [127:0] col_in_180,
    input [127:0] col_in_181,
    input [127:0] col_in_182,
    input [127:0] col_in_183,
    input [127:0] col_in_184,
    input [127:0] col_in_185,
    input [127:0] col_in_186,
    input [127:0] col_in_187,
    input [127:0] col_in_188,
    input [127:0] col_in_189,
    input [127:0] col_in_190,
    input [127:0] col_in_191,
    input [127:0] col_in_192,
    input [127:0] col_in_193,
    input [127:0] col_in_194,
    input [127:0] col_in_195,
    input [127:0] col_in_196,
    input [127:0] col_in_197,
    input [127:0] col_in_198,
    input [127:0] col_in_199,
    input [127:0] col_in_200,
    input [127:0] col_in_201,
    input [127:0] col_in_202,
    input [127:0] col_in_203,
    input [127:0] col_in_204,
    input [127:0] col_in_205,
    input [127:0] col_in_206,
    input [127:0] col_in_207,
    input [127:0] col_in_208,
    input [127:0] col_in_209,
    input [127:0] col_in_210,
    input [127:0] col_in_211,
    input [127:0] col_in_212,
    input [127:0] col_in_213,
    input [127:0] col_in_214,
    input [127:0] col_in_215,
    input [127:0] col_in_216,
    input [127:0] col_in_217,
    input [127:0] col_in_218,
    input [127:0] col_in_219,
    input [127:0] col_in_220,
    input [127:0] col_in_221,
    input [127:0] col_in_222,
    input [127:0] col_in_223,
    input [127:0] col_in_224,
    input [127:0] col_in_225,
    input [127:0] col_in_226,
    input [127:0] col_in_227,
    input [127:0] col_in_228,
    input [127:0] col_in_229,
    input [127:0] col_in_230,
    input [127:0] col_in_231,
    input [127:0] col_in_232,
    input [127:0] col_in_233,
    input [127:0] col_in_234,
    input [127:0] col_in_235,
    input [127:0] col_in_236,
    input [127:0] col_in_237,
    input [127:0] col_in_238,
    input [127:0] col_in_239,
    input [127:0] col_in_240,
    input [127:0] col_in_241,
    input [127:0] col_in_242,
    input [127:0] col_in_243,
    input [127:0] col_in_244,
    input [127:0] col_in_245,
    input [127:0] col_in_246,
    input [127:0] col_in_247,
    input [127:0] col_in_248,
    input [127:0] col_in_249,
    input [127:0] col_in_250,
    input [127:0] col_in_251,
    input [127:0] col_in_252,
    input [127:0] col_in_253,
    input [127:0] col_in_254,
    input [127:0] col_in_255,
    input [127:0] col_in_256,
    input [127:0] col_in_257,
    input [127:0] col_in_258,
    input [127:0] col_in_259,
    input [127:0] col_in_260,
    input [127:0] col_in_261,
    input [127:0] col_in_262,
    input [127:0] col_in_263,
    input [127:0] col_in_264,
    input [127:0] col_in_265,
    input [127:0] col_in_266,
    input [127:0] col_in_267,
    input [127:0] col_in_268,
    input [127:0] col_in_269,
    input [127:0] col_in_270,
    input [127:0] col_in_271,
    input [127:0] col_in_272,
    input [127:0] col_in_273,
    input [127:0] col_in_274,
    input [127:0] col_in_275,
    input [127:0] col_in_276,
    input [127:0] col_in_277,
    input [127:0] col_in_278,
    input [127:0] col_in_279,
    input [127:0] col_in_280,
    input [127:0] col_in_281,
    input [127:0] col_in_282,
    input [127:0] col_in_283,
    input [127:0] col_in_284,
    input [127:0] col_in_285,
    input [127:0] col_in_286,
    input [127:0] col_in_287,
    input [127:0] col_in_288,
    input [127:0] col_in_289,
    input [127:0] col_in_290,
    input [127:0] col_in_291,
    input [127:0] col_in_292,
    input [127:0] col_in_293,
    input [127:0] col_in_294,
    input [127:0] col_in_295,
    input [127:0] col_in_296,
    input [127:0] col_in_297,
    input [127:0] col_in_298,
    input [127:0] col_in_299,
    input [127:0] col_in_300,
    input [127:0] col_in_301,
    input [127:0] col_in_302,
    input [127:0] col_in_303,
    input [127:0] col_in_304,
    input [127:0] col_in_305,
    input [127:0] col_in_306,
    input [127:0] col_in_307,
    input [127:0] col_in_308,
    input [127:0] col_in_309,
    input [127:0] col_in_310,
    input [127:0] col_in_311,
    input [127:0] col_in_312,
    input [127:0] col_in_313,
    input [127:0] col_in_314,
    input [127:0] col_in_315,
    input [127:0] col_in_316,
    input [127:0] col_in_317,
    input [127:0] col_in_318,
    input [127:0] col_in_319,
    input [127:0] col_in_320,
    input [127:0] col_in_321,
    input [127:0] col_in_322,
    input [127:0] col_in_323,
    input [127:0] col_in_324,
    input [127:0] col_in_325,
    input [127:0] col_in_326,
    input [127:0] col_in_327,
    input [127:0] col_in_328,
    input [127:0] col_in_329,
    input [127:0] col_in_330,
    input [127:0] col_in_331,
    input [127:0] col_in_332,
    input [127:0] col_in_333,
    input [127:0] col_in_334,
    input [127:0] col_in_335,
    input [127:0] col_in_336,
    input [127:0] col_in_337,
    input [127:0] col_in_338,
    input [127:0] col_in_339,
    input [127:0] col_in_340,
    input [127:0] col_in_341,
    input [127:0] col_in_342,
    input [127:0] col_in_343,
    input [127:0] col_in_344,
    input [127:0] col_in_345,
    input [127:0] col_in_346,
    input [127:0] col_in_347,
    input [127:0] col_in_348,
    input [127:0] col_in_349,
    input [127:0] col_in_350,
    input [127:0] col_in_351,
    input [127:0] col_in_352,
    input [127:0] col_in_353,
    input [127:0] col_in_354,
    input [127:0] col_in_355,
    input [127:0] col_in_356,
    input [127:0] col_in_357,
    input [127:0] col_in_358,
    input [127:0] col_in_359,
    input [127:0] col_in_360,
    input [127:0] col_in_361,
    input [127:0] col_in_362,
    input [127:0] col_in_363,
    input [127:0] col_in_364,
    input [127:0] col_in_365,
    input [127:0] col_in_366,
    input [127:0] col_in_367,
    input [127:0] col_in_368,
    input [127:0] col_in_369,
    input [127:0] col_in_370,
    input [127:0] col_in_371,
    input [127:0] col_in_372,
    input [127:0] col_in_373,
    input [127:0] col_in_374,
    input [127:0] col_in_375,
    input [127:0] col_in_376,
    input [127:0] col_in_377,
    input [127:0] col_in_378,
    input [127:0] col_in_379,
    input [127:0] col_in_380,
    input [127:0] col_in_381,
    input [127:0] col_in_382,
    input [127:0] col_in_383,
    input [127:0] col_in_384,
    input [127:0] col_in_385,
    input [127:0] col_in_386,
    input [127:0] col_in_387,
    input [127:0] col_in_388,
    input [127:0] col_in_389,
    input [127:0] col_in_390,
    input [127:0] col_in_391,
    input [127:0] col_in_392,
    input [127:0] col_in_393,
    input [127:0] col_in_394,
    input [127:0] col_in_395,
    input [127:0] col_in_396,
    input [127:0] col_in_397,
    input [127:0] col_in_398,
    input [127:0] col_in_399,
    input [127:0] col_in_400,
    input [127:0] col_in_401,
    input [127:0] col_in_402,
    input [127:0] col_in_403,
    input [127:0] col_in_404,
    input [127:0] col_in_405,
    input [127:0] col_in_406,
    input [127:0] col_in_407,
    input [127:0] col_in_408,
    input [127:0] col_in_409,
    input [127:0] col_in_410,
    input [127:0] col_in_411,
    input [127:0] col_in_412,
    input [127:0] col_in_413,
    input [127:0] col_in_414,
    input [127:0] col_in_415,
    input [127:0] col_in_416,
    input [127:0] col_in_417,
    input [127:0] col_in_418,
    input [127:0] col_in_419,
    input [127:0] col_in_420,
    input [127:0] col_in_421,
    input [127:0] col_in_422,
    input [127:0] col_in_423,
    input [127:0] col_in_424,
    input [127:0] col_in_425,
    input [127:0] col_in_426,
    input [127:0] col_in_427,
    input [127:0] col_in_428,
    input [127:0] col_in_429,
    input [127:0] col_in_430,
    input [127:0] col_in_431,
    input [127:0] col_in_432,
    input [127:0] col_in_433,
    input [127:0] col_in_434,
    input [127:0] col_in_435,
    input [127:0] col_in_436,
    input [127:0] col_in_437,
    input [127:0] col_in_438,
    input [127:0] col_in_439,
    input [127:0] col_in_440,
    input [127:0] col_in_441,
    input [127:0] col_in_442,
    input [127:0] col_in_443,
    input [127:0] col_in_444,
    input [127:0] col_in_445,
    input [127:0] col_in_446,
    input [127:0] col_in_447,
    input [127:0] col_in_448,
    input [127:0] col_in_449,
    input [127:0] col_in_450,
    input [127:0] col_in_451,
    input [127:0] col_in_452,
    input [127:0] col_in_453,
    input [127:0] col_in_454,
    input [127:0] col_in_455,
    input [127:0] col_in_456,
    input [127:0] col_in_457,
    input [127:0] col_in_458,
    input [127:0] col_in_459,
    input [127:0] col_in_460,
    input [127:0] col_in_461,
    input [127:0] col_in_462,
    input [127:0] col_in_463,
    input [127:0] col_in_464,
    input [127:0] col_in_465,
    input [127:0] col_in_466,
    input [127:0] col_in_467,
    input [127:0] col_in_468,
    input [127:0] col_in_469,
    input [127:0] col_in_470,
    input [127:0] col_in_471,
    input [127:0] col_in_472,
    input [127:0] col_in_473,
    input [127:0] col_in_474,
    input [127:0] col_in_475,
    input [127:0] col_in_476,
    input [127:0] col_in_477,
    input [127:0] col_in_478,
    input [127:0] col_in_479,
    input [127:0] col_in_480,
    input [127:0] col_in_481,
    input [127:0] col_in_482,
    input [127:0] col_in_483,
    input [127:0] col_in_484,
    input [127:0] col_in_485,
    input [127:0] col_in_486,
    input [127:0] col_in_487,
    input [127:0] col_in_488,
    input [127:0] col_in_489,
    input [127:0] col_in_490,
    input [127:0] col_in_491,
    input [127:0] col_in_492,
    input [127:0] col_in_493,
    input [127:0] col_in_494,
    input [127:0] col_in_495,
    input [127:0] col_in_496,
    input [127:0] col_in_497,
    input [127:0] col_in_498,
    input [127:0] col_in_499,
    input [127:0] col_in_500,
    input [127:0] col_in_501,
    input [127:0] col_in_502,
    input [127:0] col_in_503,
    input [127:0] col_in_504,
    input [127:0] col_in_505,
    input [127:0] col_in_506,
    input [127:0] col_in_507,
    input [127:0] col_in_508,
    input [127:0] col_in_509,
    input [127:0] col_in_510,
    input [127:0] col_in_511,
    input [127:0] col_in_512,
    input [127:0] col_in_513,
    input [127:0] col_in_514,
    input [127:0] col_in_515,
    input [127:0] col_in_516,
    input [127:0] col_in_517,
    input [127:0] col_in_518,
    input [127:0] col_in_519,
    input [127:0] col_in_520,
    input [127:0] col_in_521,
    input [127:0] col_in_522,
    input [127:0] col_in_523,
    input [127:0] col_in_524,
    input [127:0] col_in_525,
    input [127:0] col_in_526,
    input [127:0] col_in_527,
    input [127:0] col_in_528,
    input [127:0] col_in_529,
    input [127:0] col_in_530,
    input [127:0] col_in_531,
    input [127:0] col_in_532,
    input [127:0] col_in_533,
    input [127:0] col_in_534,
    input [127:0] col_in_535,
    input [127:0] col_in_536,
    input [127:0] col_in_537,
    input [127:0] col_in_538,
    input [127:0] col_in_539,
    input [127:0] col_in_540,
    input [127:0] col_in_541,
    input [127:0] col_in_542,
    input [127:0] col_in_543,
    input [127:0] col_in_544,
    input [127:0] col_in_545,
    input [127:0] col_in_546,
    input [127:0] col_in_547,
    input [127:0] col_in_548,
    input [127:0] col_in_549,
    input [127:0] col_in_550,
    input [127:0] col_in_551,
    input [127:0] col_in_552,
    input [127:0] col_in_553,
    input [127:0] col_in_554,
    input [127:0] col_in_555,
    input [127:0] col_in_556,
    input [127:0] col_in_557,
    input [127:0] col_in_558,
    input [127:0] col_in_559,
    input [127:0] col_in_560,
    input [127:0] col_in_561,
    input [127:0] col_in_562,
    input [127:0] col_in_563,
    input [127:0] col_in_564,
    input [127:0] col_in_565,
    input [127:0] col_in_566,
    input [127:0] col_in_567,
    input [127:0] col_in_568,
    input [127:0] col_in_569,
    input [127:0] col_in_570,
    input [127:0] col_in_571,
    input [127:0] col_in_572,
    input [127:0] col_in_573,
    input [127:0] col_in_574,
    input [127:0] col_in_575,
    input [127:0] col_in_576,
    input [127:0] col_in_577,
    input [127:0] col_in_578,
    input [127:0] col_in_579,
    input [127:0] col_in_580,
    input [127:0] col_in_581,
    input [127:0] col_in_582,
    input [127:0] col_in_583,
    input [127:0] col_in_584,
    input [127:0] col_in_585,
    input [127:0] col_in_586,
    input [127:0] col_in_587,
    input [127:0] col_in_588,
    input [127:0] col_in_589,
    input [127:0] col_in_590,
    input [127:0] col_in_591,
    input [127:0] col_in_592,
    input [127:0] col_in_593,
    input [127:0] col_in_594,
    input [127:0] col_in_595,
    input [127:0] col_in_596,
    input [127:0] col_in_597,
    input [127:0] col_in_598,
    input [127:0] col_in_599,
    input [127:0] col_in_600,
    input [127:0] col_in_601,
    input [127:0] col_in_602,
    input [127:0] col_in_603,
    input [127:0] col_in_604,
    input [127:0] col_in_605,
    input [127:0] col_in_606,
    input [127:0] col_in_607,
    input [127:0] col_in_608,
    input [127:0] col_in_609,
    input [127:0] col_in_610,
    input [127:0] col_in_611,
    input [127:0] col_in_612,
    input [127:0] col_in_613,
    input [127:0] col_in_614,
    input [127:0] col_in_615,
    input [127:0] col_in_616,
    input [127:0] col_in_617,
    input [127:0] col_in_618,
    input [127:0] col_in_619,
    input [127:0] col_in_620,
    input [127:0] col_in_621,
    input [127:0] col_in_622,
    input [127:0] col_in_623,
    input [127:0] col_in_624,
    input [127:0] col_in_625,
    input [127:0] col_in_626,
    input [127:0] col_in_627,
    input [127:0] col_in_628,
    input [127:0] col_in_629,
    input [127:0] col_in_630,
    input [127:0] col_in_631,
    input [127:0] col_in_632,
    input [127:0] col_in_633,
    input [127:0] col_in_634,
    input [127:0] col_in_635,
    input [127:0] col_in_636,
    input [127:0] col_in_637,
    input [127:0] col_in_638,
    input [127:0] col_in_639,
    input [127:0] col_in_640,
    input [127:0] col_in_641,
    input [127:0] col_in_642,
    input [127:0] col_in_643,
    input [127:0] col_in_644,
    input [127:0] col_in_645,
    input [127:0] col_in_646,
    input [127:0] col_in_647,
    input [127:0] col_in_648,
    input [127:0] col_in_649,
    input [127:0] col_in_650,
    input [127:0] col_in_651,
    input [127:0] col_in_652,
    input [127:0] col_in_653,
    input [127:0] col_in_654,
    input [127:0] col_in_655,
    input [127:0] col_in_656,
    input [127:0] col_in_657,
    input [127:0] col_in_658,
    input [127:0] col_in_659,
    input [127:0] col_in_660,
    input [127:0] col_in_661,
    input [127:0] col_in_662,
    input [127:0] col_in_663,
    input [127:0] col_in_664,
    input [127:0] col_in_665,
    input [127:0] col_in_666,
    input [127:0] col_in_667,
    input [127:0] col_in_668,
    input [127:0] col_in_669,
    input [127:0] col_in_670,
    input [127:0] col_in_671,
    input [127:0] col_in_672,
    input [127:0] col_in_673,
    input [127:0] col_in_674,
    input [127:0] col_in_675,
    input [127:0] col_in_676,
    input [127:0] col_in_677,
    input [127:0] col_in_678,
    input [127:0] col_in_679,
    input [127:0] col_in_680,
    input [127:0] col_in_681,
    input [127:0] col_in_682,
    input [127:0] col_in_683,
    input [127:0] col_in_684,
    input [127:0] col_in_685,
    input [127:0] col_in_686,
    input [127:0] col_in_687,
    input [127:0] col_in_688,
    input [127:0] col_in_689,
    input [127:0] col_in_690,
    input [127:0] col_in_691,
    input [127:0] col_in_692,
    input [127:0] col_in_693,
    input [127:0] col_in_694,
    input [127:0] col_in_695,
    input [127:0] col_in_696,
    input [127:0] col_in_697,
    input [127:0] col_in_698,
    input [127:0] col_in_699,
    input [127:0] col_in_700,
    input [127:0] col_in_701,
    input [127:0] col_in_702,
    input [127:0] col_in_703,
    input [127:0] col_in_704,
    input [127:0] col_in_705,
    input [127:0] col_in_706,
    input [127:0] col_in_707,
    input [127:0] col_in_708,
    input [127:0] col_in_709,
    input [127:0] col_in_710,
    input [127:0] col_in_711,
    input [127:0] col_in_712,
    input [127:0] col_in_713,
    input [127:0] col_in_714,
    input [127:0] col_in_715,
    input [127:0] col_in_716,
    input [127:0] col_in_717,
    input [127:0] col_in_718,
    input [127:0] col_in_719,
    input [127:0] col_in_720,
    input [127:0] col_in_721,
    input [127:0] col_in_722,
    input [127:0] col_in_723,
    input [127:0] col_in_724,
    input [127:0] col_in_725,
    input [127:0] col_in_726,
    input [127:0] col_in_727,
    input [127:0] col_in_728,
    input [127:0] col_in_729,
    input [127:0] col_in_730,
    input [127:0] col_in_731,
    input [127:0] col_in_732,
    input [127:0] col_in_733,
    input [127:0] col_in_734,
    input [127:0] col_in_735,
    input [127:0] col_in_736,
    input [127:0] col_in_737,
    input [127:0] col_in_738,
    input [127:0] col_in_739,
    input [127:0] col_in_740,
    input [127:0] col_in_741,
    input [127:0] col_in_742,
    input [127:0] col_in_743,
    input [127:0] col_in_744,
    input [127:0] col_in_745,
    input [127:0] col_in_746,
    input [127:0] col_in_747,
    input [127:0] col_in_748,
    input [127:0] col_in_749,
    input [127:0] col_in_750,
    input [127:0] col_in_751,
    input [127:0] col_in_752,
    input [127:0] col_in_753,
    input [127:0] col_in_754,
    input [127:0] col_in_755,
    input [127:0] col_in_756,
    input [127:0] col_in_757,
    input [127:0] col_in_758,
    input [127:0] col_in_759,
    input [127:0] col_in_760,
    input [127:0] col_in_761,
    input [127:0] col_in_762,
    input [127:0] col_in_763,
    input [127:0] col_in_764,
    input [127:0] col_in_765,
    input [127:0] col_in_766,
    input [127:0] col_in_767,
    input [127:0] col_in_768,
    input [127:0] col_in_769,
    input [127:0] col_in_770,
    input [127:0] col_in_771,
    input [127:0] col_in_772,
    input [127:0] col_in_773,
    input [127:0] col_in_774,
    input [127:0] col_in_775,
    input [127:0] col_in_776,
    input [127:0] col_in_777,
    input [127:0] col_in_778,
    input [127:0] col_in_779,
    input [127:0] col_in_780,
    input [127:0] col_in_781,
    input [127:0] col_in_782,
    input [127:0] col_in_783,
    input [127:0] col_in_784,
    input [127:0] col_in_785,
    input [127:0] col_in_786,
    input [127:0] col_in_787,
    input [127:0] col_in_788,
    input [127:0] col_in_789,
    input [127:0] col_in_790,
    input [127:0] col_in_791,
    input [127:0] col_in_792,
    input [127:0] col_in_793,
    input [127:0] col_in_794,
    input [127:0] col_in_795,
    input [127:0] col_in_796,
    input [127:0] col_in_797,
    input [127:0] col_in_798,
    input [127:0] col_in_799,
    input [127:0] col_in_800,
    input [127:0] col_in_801,
    input [127:0] col_in_802,
    input [127:0] col_in_803,
    input [127:0] col_in_804,
    input [127:0] col_in_805,
    input [127:0] col_in_806,
    input [127:0] col_in_807,
    input [127:0] col_in_808,
    input [127:0] col_in_809,
    input [127:0] col_in_810,
    input [127:0] col_in_811,
    input [127:0] col_in_812,
    input [127:0] col_in_813,
    input [127:0] col_in_814,
    input [127:0] col_in_815,
    input [127:0] col_in_816,
    input [127:0] col_in_817,
    input [127:0] col_in_818,
    input [127:0] col_in_819,
    input [127:0] col_in_820,
    input [127:0] col_in_821,
    input [127:0] col_in_822,
    input [127:0] col_in_823,
    input [127:0] col_in_824,
    input [127:0] col_in_825,
    input [127:0] col_in_826,
    input [127:0] col_in_827,
    input [127:0] col_in_828,
    input [127:0] col_in_829,
    input [127:0] col_in_830,
    input [127:0] col_in_831,
    input [127:0] col_in_832,
    input [127:0] col_in_833,
    input [127:0] col_in_834,
    input [127:0] col_in_835,
    input [127:0] col_in_836,
    input [127:0] col_in_837,
    input [127:0] col_in_838,
    input [127:0] col_in_839,
    input [127:0] col_in_840,
    input [127:0] col_in_841,
    input [127:0] col_in_842,
    input [127:0] col_in_843,
    input [127:0] col_in_844,
    input [127:0] col_in_845,
    input [127:0] col_in_846,
    input [127:0] col_in_847,
    input [127:0] col_in_848,
    input [127:0] col_in_849,
    input [127:0] col_in_850,
    input [127:0] col_in_851,
    input [127:0] col_in_852,
    input [127:0] col_in_853,
    input [127:0] col_in_854,
    input [127:0] col_in_855,
    input [127:0] col_in_856,
    input [127:0] col_in_857,
    input [127:0] col_in_858,
    input [127:0] col_in_859,
    input [127:0] col_in_860,
    input [127:0] col_in_861,
    input [127:0] col_in_862,
    input [127:0] col_in_863,
    input [127:0] col_in_864,
    input [127:0] col_in_865,
    input [127:0] col_in_866,
    input [127:0] col_in_867,
    input [127:0] col_in_868,
    input [127:0] col_in_869,
    input [127:0] col_in_870,
    input [127:0] col_in_871,
    input [127:0] col_in_872,
    input [127:0] col_in_873,
    input [127:0] col_in_874,
    input [127:0] col_in_875,
    input [127:0] col_in_876,
    input [127:0] col_in_877,
    input [127:0] col_in_878,
    input [127:0] col_in_879,
    input [127:0] col_in_880,
    input [127:0] col_in_881,
    input [127:0] col_in_882,
    input [127:0] col_in_883,
    input [127:0] col_in_884,
    input [127:0] col_in_885,
    input [127:0] col_in_886,
    input [127:0] col_in_887,
    input [127:0] col_in_888,
    input [127:0] col_in_889,
    input [127:0] col_in_890,
    input [127:0] col_in_891,
    input [127:0] col_in_892,
    input [127:0] col_in_893,
    input [127:0] col_in_894,
    input [127:0] col_in_895,
    input [127:0] col_in_896,
    input [127:0] col_in_897,
    input [127:0] col_in_898,
    input [127:0] col_in_899,
    input [127:0] col_in_900,
    input [127:0] col_in_901,
    input [127:0] col_in_902,
    input [127:0] col_in_903,
    input [127:0] col_in_904,
    input [127:0] col_in_905,
    input [127:0] col_in_906,
    input [127:0] col_in_907,
    input [127:0] col_in_908,
    input [127:0] col_in_909,
    input [127:0] col_in_910,
    input [127:0] col_in_911,
    input [127:0] col_in_912,
    input [127:0] col_in_913,
    input [127:0] col_in_914,
    input [127:0] col_in_915,
    input [127:0] col_in_916,
    input [127:0] col_in_917,
    input [127:0] col_in_918,
    input [127:0] col_in_919,
    input [127:0] col_in_920,
    input [127:0] col_in_921,
    input [127:0] col_in_922,
    input [127:0] col_in_923,
    input [127:0] col_in_924,
    input [127:0] col_in_925,
    input [127:0] col_in_926,
    input [127:0] col_in_927,
    input [127:0] col_in_928,
    input [127:0] col_in_929,
    input [127:0] col_in_930,
    input [127:0] col_in_931,
    input [127:0] col_in_932,
    input [127:0] col_in_933,
    input [127:0] col_in_934,
    input [127:0] col_in_935,
    input [127:0] col_in_936,
    input [127:0] col_in_937,
    input [127:0] col_in_938,
    input [127:0] col_in_939,
    input [127:0] col_in_940,
    input [127:0] col_in_941,
    input [127:0] col_in_942,
    input [127:0] col_in_943,
    input [127:0] col_in_944,
    input [127:0] col_in_945,
    input [127:0] col_in_946,
    input [127:0] col_in_947,
    input [127:0] col_in_948,
    input [127:0] col_in_949,
    input [127:0] col_in_950,
    input [127:0] col_in_951,
    input [127:0] col_in_952,
    input [127:0] col_in_953,
    input [127:0] col_in_954,
    input [127:0] col_in_955,
    input [127:0] col_in_956,
    input [127:0] col_in_957,
    input [127:0] col_in_958,
    input [127:0] col_in_959,
    input [127:0] col_in_960,
    input [127:0] col_in_961,
    input [127:0] col_in_962,
    input [127:0] col_in_963,
    input [127:0] col_in_964,
    input [127:0] col_in_965,
    input [127:0] col_in_966,
    input [127:0] col_in_967,
    input [127:0] col_in_968,
    input [127:0] col_in_969,
    input [127:0] col_in_970,
    input [127:0] col_in_971,
    input [127:0] col_in_972,
    input [127:0] col_in_973,
    input [127:0] col_in_974,
    input [127:0] col_in_975,
    input [127:0] col_in_976,
    input [127:0] col_in_977,
    input [127:0] col_in_978,
    input [127:0] col_in_979,
    input [127:0] col_in_980,
    input [127:0] col_in_981,
    input [127:0] col_in_982,
    input [127:0] col_in_983,
    input [127:0] col_in_984,
    input [127:0] col_in_985,
    input [127:0] col_in_986,
    input [127:0] col_in_987,
    input [127:0] col_in_988,
    input [127:0] col_in_989,
    input [127:0] col_in_990,
    input [127:0] col_in_991,
    input [127:0] col_in_992,
    input [127:0] col_in_993,
    input [127:0] col_in_994,
    input [127:0] col_in_995,
    input [127:0] col_in_996,
    input [127:0] col_in_997,
    input [127:0] col_in_998,
    input [127:0] col_in_999,
    input [127:0] col_in_1000,
    input [127:0] col_in_1001,
    input [127:0] col_in_1002,
    input [127:0] col_in_1003,
    input [127:0] col_in_1004,
    input [127:0] col_in_1005,
    input [127:0] col_in_1006,
    input [127:0] col_in_1007,
    input [127:0] col_in_1008,
    input [127:0] col_in_1009,
    input [127:0] col_in_1010,
    input [127:0] col_in_1011,
    input [127:0] col_in_1012,
    input [127:0] col_in_1013,
    input [127:0] col_in_1014,
    input [127:0] col_in_1015,
    input [127:0] col_in_1016,
    input [127:0] col_in_1017,
    input [127:0] col_in_1018,
    input [127:0] col_in_1019,
    input [127:0] col_in_1020,
    input [127:0] col_in_1021,
    input [127:0] col_in_1022,
    input [127:0] col_in_1023,
    input [127:0] col_in_1024,
    input [127:0] col_in_1025,
    input [127:0] col_in_1026,
    input [127:0] col_in_1027,
    input [127:0] col_in_1028,
    input [127:0] col_in_1029,
    input [127:0] col_in_1030,
    input [127:0] col_in_1031,
    input [127:0] col_in_1032,
    input [127:0] col_in_1033,
    input [127:0] col_in_1034,
    input [127:0] col_in_1035,
    input [127:0] col_in_1036,
    input [127:0] col_in_1037,
    input [127:0] col_in_1038,
    input [127:0] col_in_1039,
    input [127:0] col_in_1040,
    input [127:0] col_in_1041,
    input [127:0] col_in_1042,
    input [127:0] col_in_1043,
    input [127:0] col_in_1044,
    input [127:0] col_in_1045,
    input [127:0] col_in_1046,
    input [127:0] col_in_1047,
    input [127:0] col_in_1048,
    input [127:0] col_in_1049,
    input [127:0] col_in_1050,
    input [127:0] col_in_1051,
    input [127:0] col_in_1052,
    input [127:0] col_in_1053,
    input [127:0] col_in_1054,
    input [127:0] col_in_1055,
    input [127:0] col_in_1056,
    input [127:0] col_in_1057,
    input [127:0] col_in_1058,
    input [127:0] col_in_1059,
    input [127:0] col_in_1060,
    input [127:0] col_in_1061,
    input [127:0] col_in_1062,
    input [127:0] col_in_1063,
    input [127:0] col_in_1064,
    input [127:0] col_in_1065,
    input [127:0] col_in_1066,
    input [127:0] col_in_1067,
    input [127:0] col_in_1068,
    input [127:0] col_in_1069,
    input [127:0] col_in_1070,
    input [127:0] col_in_1071,
    input [127:0] col_in_1072,
    input [127:0] col_in_1073,
    input [127:0] col_in_1074,
    input [127:0] col_in_1075,
    input [127:0] col_in_1076,
    input [127:0] col_in_1077,
    input [127:0] col_in_1078,
    input [127:0] col_in_1079,
    input [127:0] col_in_1080,
    input [127:0] col_in_1081,
    input [127:0] col_in_1082,
    input [127:0] col_in_1083,
    input [127:0] col_in_1084,
    input [127:0] col_in_1085,
    input [127:0] col_in_1086,
    input [127:0] col_in_1087,
    input [127:0] col_in_1088,
    input [127:0] col_in_1089,
    input [127:0] col_in_1090,
    input [127:0] col_in_1091,
    input [127:0] col_in_1092,
    input [127:0] col_in_1093,
    input [127:0] col_in_1094,
    input [127:0] col_in_1095,
    input [127:0] col_in_1096,
    input [127:0] col_in_1097,
    input [127:0] col_in_1098,
    input [127:0] col_in_1099,
    input [127:0] col_in_1100,
    input [127:0] col_in_1101,
    input [127:0] col_in_1102,
    input [127:0] col_in_1103,
    input [127:0] col_in_1104,
    input [127:0] col_in_1105,
    input [127:0] col_in_1106,
    input [127:0] col_in_1107,
    input [127:0] col_in_1108,
    input [127:0] col_in_1109,
    input [127:0] col_in_1110,
    input [127:0] col_in_1111,
    input [127:0] col_in_1112,
    input [127:0] col_in_1113,
    input [127:0] col_in_1114,
    input [127:0] col_in_1115,
    input [127:0] col_in_1116,
    input [127:0] col_in_1117,
    input [127:0] col_in_1118,
    input [127:0] col_in_1119,
    input [127:0] col_in_1120,
    input [127:0] col_in_1121,
    input [127:0] col_in_1122,
    input [127:0] col_in_1123,
    input [127:0] col_in_1124,
    input [127:0] col_in_1125,
    input [127:0] col_in_1126,
    input [127:0] col_in_1127,
    input [127:0] col_in_1128,
    input [127:0] col_in_1129,
    input [127:0] col_in_1130,
    input [127:0] col_in_1131,
    input [127:0] col_in_1132,
    input [127:0] col_in_1133,
    input [127:0] col_in_1134,
    input [127:0] col_in_1135,
    input [127:0] col_in_1136,
    input [127:0] col_in_1137,
    input [127:0] col_in_1138,
    input [127:0] col_in_1139,
    input [127:0] col_in_1140,
    input [127:0] col_in_1141,
    input [127:0] col_in_1142,
    input [127:0] col_in_1143,
    input [127:0] col_in_1144,
    input [127:0] col_in_1145,
    input [127:0] col_in_1146,
    input [127:0] col_in_1147,
    input [127:0] col_in_1148,
    input [127:0] col_in_1149,
    input [127:0] col_in_1150,
    input [127:0] col_in_1151,
    input [127:0] col_in_1152,
    input [127:0] col_in_1153,
    input [127:0] col_in_1154,
    input [127:0] col_in_1155,
    input [127:0] col_in_1156,
    input [127:0] col_in_1157,
    input [127:0] col_in_1158,
    input [127:0] col_in_1159,
    input [127:0] col_in_1160,
    input [127:0] col_in_1161,
    input [127:0] col_in_1162,
    input [127:0] col_in_1163,
    input [127:0] col_in_1164,
    input [127:0] col_in_1165,
    input [127:0] col_in_1166,
    input [127:0] col_in_1167,
    input [127:0] col_in_1168,
    input [127:0] col_in_1169,
    input [127:0] col_in_1170,
    input [127:0] col_in_1171,
    input [127:0] col_in_1172,
    input [127:0] col_in_1173,
    input [127:0] col_in_1174,
    input [127:0] col_in_1175,
    input [127:0] col_in_1176,
    input [127:0] col_in_1177,
    input [127:0] col_in_1178,
    input [127:0] col_in_1179,
    input [127:0] col_in_1180,
    input [127:0] col_in_1181,
    input [127:0] col_in_1182,
    input [127:0] col_in_1183,
    input [127:0] col_in_1184,
    input [127:0] col_in_1185,
    input [127:0] col_in_1186,
    input [127:0] col_in_1187,
    input [127:0] col_in_1188,
    input [127:0] col_in_1189,
    input [127:0] col_in_1190,
    input [127:0] col_in_1191,
    input [127:0] col_in_1192,
    input [127:0] col_in_1193,
    input [127:0] col_in_1194,
    input [127:0] col_in_1195,
    input [127:0] col_in_1196,
    input [127:0] col_in_1197,
    input [127:0] col_in_1198,
    input [127:0] col_in_1199,
    input [127:0] col_in_1200,
    input [127:0] col_in_1201,
    input [127:0] col_in_1202,
    input [127:0] col_in_1203,
    input [127:0] col_in_1204,
    input [127:0] col_in_1205,
    input [127:0] col_in_1206,
    input [127:0] col_in_1207,
    input [127:0] col_in_1208,
    input [127:0] col_in_1209,
    input [127:0] col_in_1210,
    input [127:0] col_in_1211,
    input [127:0] col_in_1212,
    input [127:0] col_in_1213,
    input [127:0] col_in_1214,
    input [127:0] col_in_1215,
    input [127:0] col_in_1216,
    input [127:0] col_in_1217,
    input [127:0] col_in_1218,
    input [127:0] col_in_1219,
    input [127:0] col_in_1220,
    input [127:0] col_in_1221,
    input [127:0] col_in_1222,
    input [127:0] col_in_1223,
    input [127:0] col_in_1224,
    input [127:0] col_in_1225,
    input [127:0] col_in_1226,
    input [127:0] col_in_1227,
    input [127:0] col_in_1228,
    input [127:0] col_in_1229,
    input [127:0] col_in_1230,
    input [127:0] col_in_1231,
    input [127:0] col_in_1232,
    input [127:0] col_in_1233,
    input [127:0] col_in_1234,
    input [127:0] col_in_1235,
    input [127:0] col_in_1236,
    input [127:0] col_in_1237,
    input [127:0] col_in_1238,
    input [127:0] col_in_1239,
    input [127:0] col_in_1240,
    input [127:0] col_in_1241,
    input [127:0] col_in_1242,
    input [127:0] col_in_1243,
    input [127:0] col_in_1244,
    input [127:0] col_in_1245,
    input [127:0] col_in_1246,
    input [127:0] col_in_1247,
    input [127:0] col_in_1248,
    input [127:0] col_in_1249,
    input [127:0] col_in_1250,
    input [127:0] col_in_1251,
    input [127:0] col_in_1252,
    input [127:0] col_in_1253,
    input [127:0] col_in_1254,
    input [127:0] col_in_1255,
    input [127:0] col_in_1256,
    input [127:0] col_in_1257,
    input [127:0] col_in_1258,
    input [127:0] col_in_1259,
    input [127:0] col_in_1260,
    input [127:0] col_in_1261,
    input [127:0] col_in_1262,
    input [127:0] col_in_1263,
    input [127:0] col_in_1264,
    input [127:0] col_in_1265,
    input [127:0] col_in_1266,
    input [127:0] col_in_1267,
    input [127:0] col_in_1268,
    input [127:0] col_in_1269,
    input [127:0] col_in_1270,
    input [127:0] col_in_1271,
    input [127:0] col_in_1272,
    input [127:0] col_in_1273,
    input [127:0] col_in_1274,
    input [127:0] col_in_1275,
    input [127:0] col_in_1276,
    input [127:0] col_in_1277,
    input [127:0] col_in_1278,
    input [127:0] col_in_1279,


    output [1023:0] ms
);


localparam P1 = 1026'hb0ad4555c1ee34c8cb0577d7105a475171760330d577a0777ddcb955b302ad0803487d78ca267e8e9f5e3f46e35e10ca641a27e622b2d04bb09f3f5e3ad274b1744f34aeaf90fd45129a02a298dbc430f404f9988c862d10b58c91faba2aa2922f079229b0c8f88d86bfe6def7d026294ed9dee2504b5d30466f7b0488e2666b;

localparam P2 = 1026'h1615a8aab83dc6991960aefae20b48ea2e2ec0661aaef40eefbb972ab66055a100690faf1944cfd1d3ebc7e8dc6bc2194c8344fcc4565a097613e7ebc75a4e962e89e695d5f21fa8a2534054531b78861e809f331190c5a216b1923f5745545245e0f24536191f11b0d7fcdbdefa04c529db3bdc4a096ba608cdef60911c4ccd6;

localparam P3 = 1026'h21207d00145ca9e5a61106785310ed5f4546209928066e16679962c011908071809d9786a5e737babde1abdd4aa1a325f2c4e77b2681870e311ddbe1ab0775e145ced9e0c0eb2f7cf37ce07e7ca934c92dc0eecc9a592873220a5b5f02e7fe7b68d16b67d125ae9a8943fb49ce770727bec8d9ca6f0e21790d34e710d9aa73341;

//-----------------------Stage 1------------------------------------

(* max_fanout = 50 *)reg [1287:0] reg_intermediate0;
(* max_fanout = 50 *)reg [1287:0] reg_intermediate1;


wire [1026:0] temp_ms0;
wire [1026:0] temp_ms1;
wire [1026:0] temp_ms2;
wire [1026:0] temp_ms3;

(* max_fanout = 50 *)reg [1023:0] temp_ms;


wire [105:0] u0_col_out_0;
wire [105:0] u0_col_out_1;
wire [105:0] u0_col_out_2;
wire [105:0] u0_col_out_3;
wire [105:0] u0_col_out_4;
wire [105:0] u0_col_out_5;
wire [105:0] u0_col_out_6;
wire [105:0] u0_col_out_7;
wire [105:0] u0_col_out_8;
wire [105:0] u0_col_out_9;
wire [105:0] u0_col_out_10;
wire [105:0] u0_col_out_11;
wire [105:0] u0_col_out_12;
wire [105:0] u0_col_out_13;
wire [105:0] u0_col_out_14;
wire [105:0] u0_col_out_15;
wire [105:0] u0_col_out_16;
wire [105:0] u0_col_out_17;
wire [105:0] u0_col_out_18;
wire [105:0] u0_col_out_19;
wire [105:0] u0_col_out_20;
wire [105:0] u0_col_out_21;
wire [105:0] u0_col_out_22;
wire [105:0] u0_col_out_23;
wire [105:0] u0_col_out_24;
wire [105:0] u0_col_out_25;
wire [105:0] u0_col_out_26;
wire [105:0] u0_col_out_27;
wire [105:0] u0_col_out_28;
wire [105:0] u0_col_out_29;
wire [105:0] u0_col_out_30;
wire [105:0] u0_col_out_31;
wire [105:0] u0_col_out_32;
wire [105:0] u0_col_out_33;
wire [105:0] u0_col_out_34;
wire [105:0] u0_col_out_35;
wire [105:0] u0_col_out_36;
wire [105:0] u0_col_out_37;
wire [105:0] u0_col_out_38;
wire [105:0] u0_col_out_39;
wire [105:0] u0_col_out_40;
wire [105:0] u0_col_out_41;
wire [105:0] u0_col_out_42;
wire [105:0] u0_col_out_43;
wire [105:0] u0_col_out_44;
wire [105:0] u0_col_out_45;
wire [105:0] u0_col_out_46;
wire [105:0] u0_col_out_47;
wire [105:0] u0_col_out_48;
wire [105:0] u0_col_out_49;
wire [105:0] u0_col_out_50;
wire [105:0] u0_col_out_51;
wire [105:0] u0_col_out_52;
wire [105:0] u0_col_out_53;
wire [105:0] u0_col_out_54;
wire [105:0] u0_col_out_55;
wire [105:0] u0_col_out_56;
wire [105:0] u0_col_out_57;
wire [105:0] u0_col_out_58;
wire [105:0] u0_col_out_59;
wire [105:0] u0_col_out_60;
wire [105:0] u0_col_out_61;
wire [105:0] u0_col_out_62;
wire [105:0] u0_col_out_63;
wire [105:0] u0_col_out_64;
wire [105:0] u0_col_out_65;
wire [105:0] u0_col_out_66;
wire [105:0] u0_col_out_67;
wire [105:0] u0_col_out_68;
wire [105:0] u0_col_out_69;
wire [105:0] u0_col_out_70;
wire [105:0] u0_col_out_71;
wire [105:0] u0_col_out_72;
wire [105:0] u0_col_out_73;
wire [105:0] u0_col_out_74;
wire [105:0] u0_col_out_75;
wire [105:0] u0_col_out_76;
wire [105:0] u0_col_out_77;
wire [105:0] u0_col_out_78;
wire [105:0] u0_col_out_79;
wire [105:0] u0_col_out_80;
wire [105:0] u0_col_out_81;
wire [105:0] u0_col_out_82;
wire [105:0] u0_col_out_83;
wire [105:0] u0_col_out_84;
wire [105:0] u0_col_out_85;
wire [105:0] u0_col_out_86;
wire [105:0] u0_col_out_87;
wire [105:0] u0_col_out_88;
wire [105:0] u0_col_out_89;
wire [105:0] u0_col_out_90;
wire [105:0] u0_col_out_91;
wire [105:0] u0_col_out_92;
wire [105:0] u0_col_out_93;
wire [105:0] u0_col_out_94;
wire [105:0] u0_col_out_95;
wire [105:0] u0_col_out_96;
wire [105:0] u0_col_out_97;
wire [105:0] u0_col_out_98;
wire [105:0] u0_col_out_99;
wire [105:0] u0_col_out_100;
wire [105:0] u0_col_out_101;
wire [105:0] u0_col_out_102;
wire [105:0] u0_col_out_103;
wire [105:0] u0_col_out_104;
wire [105:0] u0_col_out_105;
wire [105:0] u0_col_out_106;
wire [105:0] u0_col_out_107;
wire [105:0] u0_col_out_108;
wire [105:0] u0_col_out_109;
wire [105:0] u0_col_out_110;
wire [105:0] u0_col_out_111;
wire [105:0] u0_col_out_112;
wire [105:0] u0_col_out_113;
wire [105:0] u0_col_out_114;
wire [105:0] u0_col_out_115;
wire [105:0] u0_col_out_116;
wire [105:0] u0_col_out_117;
wire [105:0] u0_col_out_118;
wire [105:0] u0_col_out_119;
wire [105:0] u0_col_out_120;
wire [105:0] u0_col_out_121;
wire [105:0] u0_col_out_122;
wire [105:0] u0_col_out_123;
wire [105:0] u0_col_out_124;
wire [105:0] u0_col_out_125;
wire [105:0] u0_col_out_126;
wire [105:0] u0_col_out_127;
wire [105:0] u0_col_out_128;
wire [105:0] u0_col_out_129;
wire [105:0] u0_col_out_130;
wire [105:0] u0_col_out_131;
wire [105:0] u0_col_out_132;
wire [105:0] u0_col_out_133;
wire [105:0] u0_col_out_134;
wire [105:0] u0_col_out_135;
wire [105:0] u0_col_out_136;
wire [105:0] u0_col_out_137;
wire [105:0] u0_col_out_138;
wire [105:0] u0_col_out_139;
wire [105:0] u0_col_out_140;
wire [105:0] u0_col_out_141;
wire [105:0] u0_col_out_142;
wire [105:0] u0_col_out_143;
wire [105:0] u0_col_out_144;
wire [105:0] u0_col_out_145;
wire [105:0] u0_col_out_146;
wire [105:0] u0_col_out_147;
wire [105:0] u0_col_out_148;
wire [105:0] u0_col_out_149;
wire [105:0] u0_col_out_150;
wire [105:0] u0_col_out_151;
wire [105:0] u0_col_out_152;
wire [105:0] u0_col_out_153;
wire [105:0] u0_col_out_154;
wire [105:0] u0_col_out_155;
wire [105:0] u0_col_out_156;
wire [105:0] u0_col_out_157;
wire [105:0] u0_col_out_158;
wire [105:0] u0_col_out_159;
wire [105:0] u0_col_out_160;
wire [105:0] u0_col_out_161;
wire [105:0] u0_col_out_162;
wire [105:0] u0_col_out_163;
wire [105:0] u0_col_out_164;
wire [105:0] u0_col_out_165;
wire [105:0] u0_col_out_166;
wire [105:0] u0_col_out_167;
wire [105:0] u0_col_out_168;
wire [105:0] u0_col_out_169;
wire [105:0] u0_col_out_170;
wire [105:0] u0_col_out_171;
wire [105:0] u0_col_out_172;
wire [105:0] u0_col_out_173;
wire [105:0] u0_col_out_174;
wire [105:0] u0_col_out_175;
wire [105:0] u0_col_out_176;
wire [105:0] u0_col_out_177;
wire [105:0] u0_col_out_178;
wire [105:0] u0_col_out_179;
wire [105:0] u0_col_out_180;
wire [105:0] u0_col_out_181;
wire [105:0] u0_col_out_182;
wire [105:0] u0_col_out_183;
wire [105:0] u0_col_out_184;
wire [105:0] u0_col_out_185;
wire [105:0] u0_col_out_186;
wire [105:0] u0_col_out_187;
wire [105:0] u0_col_out_188;
wire [105:0] u0_col_out_189;
wire [105:0] u0_col_out_190;
wire [105:0] u0_col_out_191;
wire [105:0] u0_col_out_192;
wire [105:0] u0_col_out_193;
wire [105:0] u0_col_out_194;
wire [105:0] u0_col_out_195;
wire [105:0] u0_col_out_196;
wire [105:0] u0_col_out_197;
wire [105:0] u0_col_out_198;
wire [105:0] u0_col_out_199;
wire [105:0] u0_col_out_200;
wire [105:0] u0_col_out_201;
wire [105:0] u0_col_out_202;
wire [105:0] u0_col_out_203;
wire [105:0] u0_col_out_204;
wire [105:0] u0_col_out_205;
wire [105:0] u0_col_out_206;
wire [105:0] u0_col_out_207;
wire [105:0] u0_col_out_208;
wire [105:0] u0_col_out_209;
wire [105:0] u0_col_out_210;
wire [105:0] u0_col_out_211;
wire [105:0] u0_col_out_212;
wire [105:0] u0_col_out_213;
wire [105:0] u0_col_out_214;
wire [105:0] u0_col_out_215;
wire [105:0] u0_col_out_216;
wire [105:0] u0_col_out_217;
wire [105:0] u0_col_out_218;
wire [105:0] u0_col_out_219;
wire [105:0] u0_col_out_220;
wire [105:0] u0_col_out_221;
wire [105:0] u0_col_out_222;
wire [105:0] u0_col_out_223;
wire [105:0] u0_col_out_224;
wire [105:0] u0_col_out_225;
wire [105:0] u0_col_out_226;
wire [105:0] u0_col_out_227;
wire [105:0] u0_col_out_228;
wire [105:0] u0_col_out_229;
wire [105:0] u0_col_out_230;
wire [105:0] u0_col_out_231;
wire [105:0] u0_col_out_232;
wire [105:0] u0_col_out_233;
wire [105:0] u0_col_out_234;
wire [105:0] u0_col_out_235;
wire [105:0] u0_col_out_236;
wire [105:0] u0_col_out_237;
wire [105:0] u0_col_out_238;
wire [105:0] u0_col_out_239;
wire [105:0] u0_col_out_240;
wire [105:0] u0_col_out_241;
wire [105:0] u0_col_out_242;
wire [105:0] u0_col_out_243;
wire [105:0] u0_col_out_244;
wire [105:0] u0_col_out_245;
wire [105:0] u0_col_out_246;
wire [105:0] u0_col_out_247;
wire [105:0] u0_col_out_248;
wire [105:0] u0_col_out_249;
wire [105:0] u0_col_out_250;
wire [105:0] u0_col_out_251;
wire [105:0] u0_col_out_252;
wire [105:0] u0_col_out_253;
wire [105:0] u0_col_out_254;
wire [105:0] u0_col_out_255;
wire [105:0] u0_col_out_256;
wire [105:0] u0_col_out_257;
wire [105:0] u0_col_out_258;
wire [105:0] u0_col_out_259;
wire [105:0] u0_col_out_260;
wire [105:0] u0_col_out_261;
wire [105:0] u0_col_out_262;
wire [105:0] u0_col_out_263;
wire [105:0] u0_col_out_264;
wire [105:0] u0_col_out_265;
wire [105:0] u0_col_out_266;
wire [105:0] u0_col_out_267;
wire [105:0] u0_col_out_268;
wire [105:0] u0_col_out_269;
wire [105:0] u0_col_out_270;
wire [105:0] u0_col_out_271;
wire [105:0] u0_col_out_272;
wire [105:0] u0_col_out_273;
wire [105:0] u0_col_out_274;
wire [105:0] u0_col_out_275;
wire [105:0] u0_col_out_276;
wire [105:0] u0_col_out_277;
wire [105:0] u0_col_out_278;
wire [105:0] u0_col_out_279;
wire [105:0] u0_col_out_280;
wire [105:0] u0_col_out_281;
wire [105:0] u0_col_out_282;
wire [105:0] u0_col_out_283;
wire [105:0] u0_col_out_284;
wire [105:0] u0_col_out_285;
wire [105:0] u0_col_out_286;
wire [105:0] u0_col_out_287;
wire [105:0] u0_col_out_288;
wire [105:0] u0_col_out_289;
wire [105:0] u0_col_out_290;
wire [105:0] u0_col_out_291;
wire [105:0] u0_col_out_292;
wire [105:0] u0_col_out_293;
wire [105:0] u0_col_out_294;
wire [105:0] u0_col_out_295;
wire [105:0] u0_col_out_296;
wire [105:0] u0_col_out_297;
wire [105:0] u0_col_out_298;
wire [105:0] u0_col_out_299;
wire [105:0] u0_col_out_300;
wire [105:0] u0_col_out_301;
wire [105:0] u0_col_out_302;
wire [105:0] u0_col_out_303;
wire [105:0] u0_col_out_304;
wire [105:0] u0_col_out_305;
wire [105:0] u0_col_out_306;
wire [105:0] u0_col_out_307;
wire [105:0] u0_col_out_308;
wire [105:0] u0_col_out_309;
wire [105:0] u0_col_out_310;
wire [105:0] u0_col_out_311;
wire [105:0] u0_col_out_312;
wire [105:0] u0_col_out_313;
wire [105:0] u0_col_out_314;
wire [105:0] u0_col_out_315;
wire [105:0] u0_col_out_316;
wire [105:0] u0_col_out_317;
wire [105:0] u0_col_out_318;
wire [105:0] u0_col_out_319;
wire [105:0] u0_col_out_320;
wire [105:0] u0_col_out_321;
wire [105:0] u0_col_out_322;
wire [105:0] u0_col_out_323;
wire [105:0] u0_col_out_324;
wire [105:0] u0_col_out_325;
wire [105:0] u0_col_out_326;
wire [105:0] u0_col_out_327;
wire [105:0] u0_col_out_328;
wire [105:0] u0_col_out_329;
wire [105:0] u0_col_out_330;
wire [105:0] u0_col_out_331;
wire [105:0] u0_col_out_332;
wire [105:0] u0_col_out_333;
wire [105:0] u0_col_out_334;
wire [105:0] u0_col_out_335;
wire [105:0] u0_col_out_336;
wire [105:0] u0_col_out_337;
wire [105:0] u0_col_out_338;
wire [105:0] u0_col_out_339;
wire [105:0] u0_col_out_340;
wire [105:0] u0_col_out_341;
wire [105:0] u0_col_out_342;
wire [105:0] u0_col_out_343;
wire [105:0] u0_col_out_344;
wire [105:0] u0_col_out_345;
wire [105:0] u0_col_out_346;
wire [105:0] u0_col_out_347;
wire [105:0] u0_col_out_348;
wire [105:0] u0_col_out_349;
wire [105:0] u0_col_out_350;
wire [105:0] u0_col_out_351;
wire [105:0] u0_col_out_352;
wire [105:0] u0_col_out_353;
wire [105:0] u0_col_out_354;
wire [105:0] u0_col_out_355;
wire [105:0] u0_col_out_356;
wire [105:0] u0_col_out_357;
wire [105:0] u0_col_out_358;
wire [105:0] u0_col_out_359;
wire [105:0] u0_col_out_360;
wire [105:0] u0_col_out_361;
wire [105:0] u0_col_out_362;
wire [105:0] u0_col_out_363;
wire [105:0] u0_col_out_364;
wire [105:0] u0_col_out_365;
wire [105:0] u0_col_out_366;
wire [105:0] u0_col_out_367;
wire [105:0] u0_col_out_368;
wire [105:0] u0_col_out_369;
wire [105:0] u0_col_out_370;
wire [105:0] u0_col_out_371;
wire [105:0] u0_col_out_372;
wire [105:0] u0_col_out_373;
wire [105:0] u0_col_out_374;
wire [105:0] u0_col_out_375;
wire [105:0] u0_col_out_376;
wire [105:0] u0_col_out_377;
wire [105:0] u0_col_out_378;
wire [105:0] u0_col_out_379;
wire [105:0] u0_col_out_380;
wire [105:0] u0_col_out_381;
wire [105:0] u0_col_out_382;
wire [105:0] u0_col_out_383;
wire [105:0] u0_col_out_384;
wire [105:0] u0_col_out_385;
wire [105:0] u0_col_out_386;
wire [105:0] u0_col_out_387;
wire [105:0] u0_col_out_388;
wire [105:0] u0_col_out_389;
wire [105:0] u0_col_out_390;
wire [105:0] u0_col_out_391;
wire [105:0] u0_col_out_392;
wire [105:0] u0_col_out_393;
wire [105:0] u0_col_out_394;
wire [105:0] u0_col_out_395;
wire [105:0] u0_col_out_396;
wire [105:0] u0_col_out_397;
wire [105:0] u0_col_out_398;
wire [105:0] u0_col_out_399;
wire [105:0] u0_col_out_400;
wire [105:0] u0_col_out_401;
wire [105:0] u0_col_out_402;
wire [105:0] u0_col_out_403;
wire [105:0] u0_col_out_404;
wire [105:0] u0_col_out_405;
wire [105:0] u0_col_out_406;
wire [105:0] u0_col_out_407;
wire [105:0] u0_col_out_408;
wire [105:0] u0_col_out_409;
wire [105:0] u0_col_out_410;
wire [105:0] u0_col_out_411;
wire [105:0] u0_col_out_412;
wire [105:0] u0_col_out_413;
wire [105:0] u0_col_out_414;
wire [105:0] u0_col_out_415;
wire [105:0] u0_col_out_416;
wire [105:0] u0_col_out_417;
wire [105:0] u0_col_out_418;
wire [105:0] u0_col_out_419;
wire [105:0] u0_col_out_420;
wire [105:0] u0_col_out_421;
wire [105:0] u0_col_out_422;
wire [105:0] u0_col_out_423;
wire [105:0] u0_col_out_424;
wire [105:0] u0_col_out_425;
wire [105:0] u0_col_out_426;
wire [105:0] u0_col_out_427;
wire [105:0] u0_col_out_428;
wire [105:0] u0_col_out_429;
wire [105:0] u0_col_out_430;
wire [105:0] u0_col_out_431;
wire [105:0] u0_col_out_432;
wire [105:0] u0_col_out_433;
wire [105:0] u0_col_out_434;
wire [105:0] u0_col_out_435;
wire [105:0] u0_col_out_436;
wire [105:0] u0_col_out_437;
wire [105:0] u0_col_out_438;
wire [105:0] u0_col_out_439;
wire [105:0] u0_col_out_440;
wire [105:0] u0_col_out_441;
wire [105:0] u0_col_out_442;
wire [105:0] u0_col_out_443;
wire [105:0] u0_col_out_444;
wire [105:0] u0_col_out_445;
wire [105:0] u0_col_out_446;
wire [105:0] u0_col_out_447;
wire [105:0] u0_col_out_448;
wire [105:0] u0_col_out_449;
wire [105:0] u0_col_out_450;
wire [105:0] u0_col_out_451;
wire [105:0] u0_col_out_452;
wire [105:0] u0_col_out_453;
wire [105:0] u0_col_out_454;
wire [105:0] u0_col_out_455;
wire [105:0] u0_col_out_456;
wire [105:0] u0_col_out_457;
wire [105:0] u0_col_out_458;
wire [105:0] u0_col_out_459;
wire [105:0] u0_col_out_460;
wire [105:0] u0_col_out_461;
wire [105:0] u0_col_out_462;
wire [105:0] u0_col_out_463;
wire [105:0] u0_col_out_464;
wire [105:0] u0_col_out_465;
wire [105:0] u0_col_out_466;
wire [105:0] u0_col_out_467;
wire [105:0] u0_col_out_468;
wire [105:0] u0_col_out_469;
wire [105:0] u0_col_out_470;
wire [105:0] u0_col_out_471;
wire [105:0] u0_col_out_472;
wire [105:0] u0_col_out_473;
wire [105:0] u0_col_out_474;
wire [105:0] u0_col_out_475;
wire [105:0] u0_col_out_476;
wire [105:0] u0_col_out_477;
wire [105:0] u0_col_out_478;
wire [105:0] u0_col_out_479;
wire [105:0] u0_col_out_480;
wire [105:0] u0_col_out_481;
wire [105:0] u0_col_out_482;
wire [105:0] u0_col_out_483;
wire [105:0] u0_col_out_484;
wire [105:0] u0_col_out_485;
wire [105:0] u0_col_out_486;
wire [105:0] u0_col_out_487;
wire [105:0] u0_col_out_488;
wire [105:0] u0_col_out_489;
wire [105:0] u0_col_out_490;
wire [105:0] u0_col_out_491;
wire [105:0] u0_col_out_492;
wire [105:0] u0_col_out_493;
wire [105:0] u0_col_out_494;
wire [105:0] u0_col_out_495;
wire [105:0] u0_col_out_496;
wire [105:0] u0_col_out_497;
wire [105:0] u0_col_out_498;
wire [105:0] u0_col_out_499;
wire [105:0] u0_col_out_500;
wire [105:0] u0_col_out_501;
wire [105:0] u0_col_out_502;
wire [105:0] u0_col_out_503;
wire [105:0] u0_col_out_504;
wire [105:0] u0_col_out_505;
wire [105:0] u0_col_out_506;
wire [105:0] u0_col_out_507;
wire [105:0] u0_col_out_508;
wire [105:0] u0_col_out_509;
wire [105:0] u0_col_out_510;
wire [105:0] u0_col_out_511;
wire [105:0] u0_col_out_512;
wire [105:0] u0_col_out_513;
wire [105:0] u0_col_out_514;
wire [105:0] u0_col_out_515;
wire [105:0] u0_col_out_516;
wire [105:0] u0_col_out_517;
wire [105:0] u0_col_out_518;
wire [105:0] u0_col_out_519;
wire [105:0] u0_col_out_520;
wire [105:0] u0_col_out_521;
wire [105:0] u0_col_out_522;
wire [105:0] u0_col_out_523;
wire [105:0] u0_col_out_524;
wire [105:0] u0_col_out_525;
wire [105:0] u0_col_out_526;
wire [105:0] u0_col_out_527;
wire [105:0] u0_col_out_528;
wire [105:0] u0_col_out_529;
wire [105:0] u0_col_out_530;
wire [105:0] u0_col_out_531;
wire [105:0] u0_col_out_532;
wire [105:0] u0_col_out_533;
wire [105:0] u0_col_out_534;
wire [105:0] u0_col_out_535;
wire [105:0] u0_col_out_536;
wire [105:0] u0_col_out_537;
wire [105:0] u0_col_out_538;
wire [105:0] u0_col_out_539;
wire [105:0] u0_col_out_540;
wire [105:0] u0_col_out_541;
wire [105:0] u0_col_out_542;
wire [105:0] u0_col_out_543;
wire [105:0] u0_col_out_544;
wire [105:0] u0_col_out_545;
wire [105:0] u0_col_out_546;
wire [105:0] u0_col_out_547;
wire [105:0] u0_col_out_548;
wire [105:0] u0_col_out_549;
wire [105:0] u0_col_out_550;
wire [105:0] u0_col_out_551;
wire [105:0] u0_col_out_552;
wire [105:0] u0_col_out_553;
wire [105:0] u0_col_out_554;
wire [105:0] u0_col_out_555;
wire [105:0] u0_col_out_556;
wire [105:0] u0_col_out_557;
wire [105:0] u0_col_out_558;
wire [105:0] u0_col_out_559;
wire [105:0] u0_col_out_560;
wire [105:0] u0_col_out_561;
wire [105:0] u0_col_out_562;
wire [105:0] u0_col_out_563;
wire [105:0] u0_col_out_564;
wire [105:0] u0_col_out_565;
wire [105:0] u0_col_out_566;
wire [105:0] u0_col_out_567;
wire [105:0] u0_col_out_568;
wire [105:0] u0_col_out_569;
wire [105:0] u0_col_out_570;
wire [105:0] u0_col_out_571;
wire [105:0] u0_col_out_572;
wire [105:0] u0_col_out_573;
wire [105:0] u0_col_out_574;
wire [105:0] u0_col_out_575;
wire [105:0] u0_col_out_576;
wire [105:0] u0_col_out_577;
wire [105:0] u0_col_out_578;
wire [105:0] u0_col_out_579;
wire [105:0] u0_col_out_580;
wire [105:0] u0_col_out_581;
wire [105:0] u0_col_out_582;
wire [105:0] u0_col_out_583;
wire [105:0] u0_col_out_584;
wire [105:0] u0_col_out_585;
wire [105:0] u0_col_out_586;
wire [105:0] u0_col_out_587;
wire [105:0] u0_col_out_588;
wire [105:0] u0_col_out_589;
wire [105:0] u0_col_out_590;
wire [105:0] u0_col_out_591;
wire [105:0] u0_col_out_592;
wire [105:0] u0_col_out_593;
wire [105:0] u0_col_out_594;
wire [105:0] u0_col_out_595;
wire [105:0] u0_col_out_596;
wire [105:0] u0_col_out_597;
wire [105:0] u0_col_out_598;
wire [105:0] u0_col_out_599;
wire [105:0] u0_col_out_600;
wire [105:0] u0_col_out_601;
wire [105:0] u0_col_out_602;
wire [105:0] u0_col_out_603;
wire [105:0] u0_col_out_604;
wire [105:0] u0_col_out_605;
wire [105:0] u0_col_out_606;
wire [105:0] u0_col_out_607;
wire [105:0] u0_col_out_608;
wire [105:0] u0_col_out_609;
wire [105:0] u0_col_out_610;
wire [105:0] u0_col_out_611;
wire [105:0] u0_col_out_612;
wire [105:0] u0_col_out_613;
wire [105:0] u0_col_out_614;
wire [105:0] u0_col_out_615;
wire [105:0] u0_col_out_616;
wire [105:0] u0_col_out_617;
wire [105:0] u0_col_out_618;
wire [105:0] u0_col_out_619;
wire [105:0] u0_col_out_620;
wire [105:0] u0_col_out_621;
wire [105:0] u0_col_out_622;
wire [105:0] u0_col_out_623;
wire [105:0] u0_col_out_624;
wire [105:0] u0_col_out_625;
wire [105:0] u0_col_out_626;
wire [105:0] u0_col_out_627;
wire [105:0] u0_col_out_628;
wire [105:0] u0_col_out_629;
wire [105:0] u0_col_out_630;
wire [105:0] u0_col_out_631;
wire [105:0] u0_col_out_632;
wire [105:0] u0_col_out_633;
wire [105:0] u0_col_out_634;
wire [105:0] u0_col_out_635;
wire [105:0] u0_col_out_636;
wire [105:0] u0_col_out_637;
wire [105:0] u0_col_out_638;
wire [105:0] u0_col_out_639;
wire [105:0] u0_col_out_640;
wire [105:0] u0_col_out_641;
wire [105:0] u0_col_out_642;
wire [105:0] u0_col_out_643;
wire [105:0] u0_col_out_644;
wire [105:0] u0_col_out_645;
wire [105:0] u0_col_out_646;
wire [105:0] u0_col_out_647;
wire [105:0] u0_col_out_648;
wire [105:0] u0_col_out_649;
wire [105:0] u0_col_out_650;
wire [105:0] u0_col_out_651;
wire [105:0] u0_col_out_652;
wire [105:0] u0_col_out_653;
wire [105:0] u0_col_out_654;
wire [105:0] u0_col_out_655;
wire [105:0] u0_col_out_656;
wire [105:0] u0_col_out_657;
wire [105:0] u0_col_out_658;
wire [105:0] u0_col_out_659;
wire [105:0] u0_col_out_660;
wire [105:0] u0_col_out_661;
wire [105:0] u0_col_out_662;
wire [105:0] u0_col_out_663;
wire [105:0] u0_col_out_664;
wire [105:0] u0_col_out_665;
wire [105:0] u0_col_out_666;
wire [105:0] u0_col_out_667;
wire [105:0] u0_col_out_668;
wire [105:0] u0_col_out_669;
wire [105:0] u0_col_out_670;
wire [105:0] u0_col_out_671;
wire [105:0] u0_col_out_672;
wire [105:0] u0_col_out_673;
wire [105:0] u0_col_out_674;
wire [105:0] u0_col_out_675;
wire [105:0] u0_col_out_676;
wire [105:0] u0_col_out_677;
wire [105:0] u0_col_out_678;
wire [105:0] u0_col_out_679;
wire [105:0] u0_col_out_680;
wire [105:0] u0_col_out_681;
wire [105:0] u0_col_out_682;
wire [105:0] u0_col_out_683;
wire [105:0] u0_col_out_684;
wire [105:0] u0_col_out_685;
wire [105:0] u0_col_out_686;
wire [105:0] u0_col_out_687;
wire [105:0] u0_col_out_688;
wire [105:0] u0_col_out_689;
wire [105:0] u0_col_out_690;
wire [105:0] u0_col_out_691;
wire [105:0] u0_col_out_692;
wire [105:0] u0_col_out_693;
wire [105:0] u0_col_out_694;
wire [105:0] u0_col_out_695;
wire [105:0] u0_col_out_696;
wire [105:0] u0_col_out_697;
wire [105:0] u0_col_out_698;
wire [105:0] u0_col_out_699;
wire [105:0] u0_col_out_700;
wire [105:0] u0_col_out_701;
wire [105:0] u0_col_out_702;
wire [105:0] u0_col_out_703;
wire [105:0] u0_col_out_704;
wire [105:0] u0_col_out_705;
wire [105:0] u0_col_out_706;
wire [105:0] u0_col_out_707;
wire [105:0] u0_col_out_708;
wire [105:0] u0_col_out_709;
wire [105:0] u0_col_out_710;
wire [105:0] u0_col_out_711;
wire [105:0] u0_col_out_712;
wire [105:0] u0_col_out_713;
wire [105:0] u0_col_out_714;
wire [105:0] u0_col_out_715;
wire [105:0] u0_col_out_716;
wire [105:0] u0_col_out_717;
wire [105:0] u0_col_out_718;
wire [105:0] u0_col_out_719;
wire [105:0] u0_col_out_720;
wire [105:0] u0_col_out_721;
wire [105:0] u0_col_out_722;
wire [105:0] u0_col_out_723;
wire [105:0] u0_col_out_724;
wire [105:0] u0_col_out_725;
wire [105:0] u0_col_out_726;
wire [105:0] u0_col_out_727;
wire [105:0] u0_col_out_728;
wire [105:0] u0_col_out_729;
wire [105:0] u0_col_out_730;
wire [105:0] u0_col_out_731;
wire [105:0] u0_col_out_732;
wire [105:0] u0_col_out_733;
wire [105:0] u0_col_out_734;
wire [105:0] u0_col_out_735;
wire [105:0] u0_col_out_736;
wire [105:0] u0_col_out_737;
wire [105:0] u0_col_out_738;
wire [105:0] u0_col_out_739;
wire [105:0] u0_col_out_740;
wire [105:0] u0_col_out_741;
wire [105:0] u0_col_out_742;
wire [105:0] u0_col_out_743;
wire [105:0] u0_col_out_744;
wire [105:0] u0_col_out_745;
wire [105:0] u0_col_out_746;
wire [105:0] u0_col_out_747;
wire [105:0] u0_col_out_748;
wire [105:0] u0_col_out_749;
wire [105:0] u0_col_out_750;
wire [105:0] u0_col_out_751;
wire [105:0] u0_col_out_752;
wire [105:0] u0_col_out_753;
wire [105:0] u0_col_out_754;
wire [105:0] u0_col_out_755;
wire [105:0] u0_col_out_756;
wire [105:0] u0_col_out_757;
wire [105:0] u0_col_out_758;
wire [105:0] u0_col_out_759;
wire [105:0] u0_col_out_760;
wire [105:0] u0_col_out_761;
wire [105:0] u0_col_out_762;
wire [105:0] u0_col_out_763;
wire [105:0] u0_col_out_764;
wire [105:0] u0_col_out_765;
wire [105:0] u0_col_out_766;
wire [105:0] u0_col_out_767;
wire [105:0] u0_col_out_768;
wire [105:0] u0_col_out_769;
wire [105:0] u0_col_out_770;
wire [105:0] u0_col_out_771;
wire [105:0] u0_col_out_772;
wire [105:0] u0_col_out_773;
wire [105:0] u0_col_out_774;
wire [105:0] u0_col_out_775;
wire [105:0] u0_col_out_776;
wire [105:0] u0_col_out_777;
wire [105:0] u0_col_out_778;
wire [105:0] u0_col_out_779;
wire [105:0] u0_col_out_780;
wire [105:0] u0_col_out_781;
wire [105:0] u0_col_out_782;
wire [105:0] u0_col_out_783;
wire [105:0] u0_col_out_784;
wire [105:0] u0_col_out_785;
wire [105:0] u0_col_out_786;
wire [105:0] u0_col_out_787;
wire [105:0] u0_col_out_788;
wire [105:0] u0_col_out_789;
wire [105:0] u0_col_out_790;
wire [105:0] u0_col_out_791;
wire [105:0] u0_col_out_792;
wire [105:0] u0_col_out_793;
wire [105:0] u0_col_out_794;
wire [105:0] u0_col_out_795;
wire [105:0] u0_col_out_796;
wire [105:0] u0_col_out_797;
wire [105:0] u0_col_out_798;
wire [105:0] u0_col_out_799;
wire [105:0] u0_col_out_800;
wire [105:0] u0_col_out_801;
wire [105:0] u0_col_out_802;
wire [105:0] u0_col_out_803;
wire [105:0] u0_col_out_804;
wire [105:0] u0_col_out_805;
wire [105:0] u0_col_out_806;
wire [105:0] u0_col_out_807;
wire [105:0] u0_col_out_808;
wire [105:0] u0_col_out_809;
wire [105:0] u0_col_out_810;
wire [105:0] u0_col_out_811;
wire [105:0] u0_col_out_812;
wire [105:0] u0_col_out_813;
wire [105:0] u0_col_out_814;
wire [105:0] u0_col_out_815;
wire [105:0] u0_col_out_816;
wire [105:0] u0_col_out_817;
wire [105:0] u0_col_out_818;
wire [105:0] u0_col_out_819;
wire [105:0] u0_col_out_820;
wire [105:0] u0_col_out_821;
wire [105:0] u0_col_out_822;
wire [105:0] u0_col_out_823;
wire [105:0] u0_col_out_824;
wire [105:0] u0_col_out_825;
wire [105:0] u0_col_out_826;
wire [105:0] u0_col_out_827;
wire [105:0] u0_col_out_828;
wire [105:0] u0_col_out_829;
wire [105:0] u0_col_out_830;
wire [105:0] u0_col_out_831;
wire [105:0] u0_col_out_832;
wire [105:0] u0_col_out_833;
wire [105:0] u0_col_out_834;
wire [105:0] u0_col_out_835;
wire [105:0] u0_col_out_836;
wire [105:0] u0_col_out_837;
wire [105:0] u0_col_out_838;
wire [105:0] u0_col_out_839;
wire [105:0] u0_col_out_840;
wire [105:0] u0_col_out_841;
wire [105:0] u0_col_out_842;
wire [105:0] u0_col_out_843;
wire [105:0] u0_col_out_844;
wire [105:0] u0_col_out_845;
wire [105:0] u0_col_out_846;
wire [105:0] u0_col_out_847;
wire [105:0] u0_col_out_848;
wire [105:0] u0_col_out_849;
wire [105:0] u0_col_out_850;
wire [105:0] u0_col_out_851;
wire [105:0] u0_col_out_852;
wire [105:0] u0_col_out_853;
wire [105:0] u0_col_out_854;
wire [105:0] u0_col_out_855;
wire [105:0] u0_col_out_856;
wire [105:0] u0_col_out_857;
wire [105:0] u0_col_out_858;
wire [105:0] u0_col_out_859;
wire [105:0] u0_col_out_860;
wire [105:0] u0_col_out_861;
wire [105:0] u0_col_out_862;
wire [105:0] u0_col_out_863;
wire [105:0] u0_col_out_864;
wire [105:0] u0_col_out_865;
wire [105:0] u0_col_out_866;
wire [105:0] u0_col_out_867;
wire [105:0] u0_col_out_868;
wire [105:0] u0_col_out_869;
wire [105:0] u0_col_out_870;
wire [105:0] u0_col_out_871;
wire [105:0] u0_col_out_872;
wire [105:0] u0_col_out_873;
wire [105:0] u0_col_out_874;
wire [105:0] u0_col_out_875;
wire [105:0] u0_col_out_876;
wire [105:0] u0_col_out_877;
wire [105:0] u0_col_out_878;
wire [105:0] u0_col_out_879;
wire [105:0] u0_col_out_880;
wire [105:0] u0_col_out_881;
wire [105:0] u0_col_out_882;
wire [105:0] u0_col_out_883;
wire [105:0] u0_col_out_884;
wire [105:0] u0_col_out_885;
wire [105:0] u0_col_out_886;
wire [105:0] u0_col_out_887;
wire [105:0] u0_col_out_888;
wire [105:0] u0_col_out_889;
wire [105:0] u0_col_out_890;
wire [105:0] u0_col_out_891;
wire [105:0] u0_col_out_892;
wire [105:0] u0_col_out_893;
wire [105:0] u0_col_out_894;
wire [105:0] u0_col_out_895;
wire [105:0] u0_col_out_896;
wire [105:0] u0_col_out_897;
wire [105:0] u0_col_out_898;
wire [105:0] u0_col_out_899;
wire [105:0] u0_col_out_900;
wire [105:0] u0_col_out_901;
wire [105:0] u0_col_out_902;
wire [105:0] u0_col_out_903;
wire [105:0] u0_col_out_904;
wire [105:0] u0_col_out_905;
wire [105:0] u0_col_out_906;
wire [105:0] u0_col_out_907;
wire [105:0] u0_col_out_908;
wire [105:0] u0_col_out_909;
wire [105:0] u0_col_out_910;
wire [105:0] u0_col_out_911;
wire [105:0] u0_col_out_912;
wire [105:0] u0_col_out_913;
wire [105:0] u0_col_out_914;
wire [105:0] u0_col_out_915;
wire [105:0] u0_col_out_916;
wire [105:0] u0_col_out_917;
wire [105:0] u0_col_out_918;
wire [105:0] u0_col_out_919;
wire [105:0] u0_col_out_920;
wire [105:0] u0_col_out_921;
wire [105:0] u0_col_out_922;
wire [105:0] u0_col_out_923;
wire [105:0] u0_col_out_924;
wire [105:0] u0_col_out_925;
wire [105:0] u0_col_out_926;
wire [105:0] u0_col_out_927;
wire [105:0] u0_col_out_928;
wire [105:0] u0_col_out_929;
wire [105:0] u0_col_out_930;
wire [105:0] u0_col_out_931;
wire [105:0] u0_col_out_932;
wire [105:0] u0_col_out_933;
wire [105:0] u0_col_out_934;
wire [105:0] u0_col_out_935;
wire [105:0] u0_col_out_936;
wire [105:0] u0_col_out_937;
wire [105:0] u0_col_out_938;
wire [105:0] u0_col_out_939;
wire [105:0] u0_col_out_940;
wire [105:0] u0_col_out_941;
wire [105:0] u0_col_out_942;
wire [105:0] u0_col_out_943;
wire [105:0] u0_col_out_944;
wire [105:0] u0_col_out_945;
wire [105:0] u0_col_out_946;
wire [105:0] u0_col_out_947;
wire [105:0] u0_col_out_948;
wire [105:0] u0_col_out_949;
wire [105:0] u0_col_out_950;
wire [105:0] u0_col_out_951;
wire [105:0] u0_col_out_952;
wire [105:0] u0_col_out_953;
wire [105:0] u0_col_out_954;
wire [105:0] u0_col_out_955;
wire [105:0] u0_col_out_956;
wire [105:0] u0_col_out_957;
wire [105:0] u0_col_out_958;
wire [105:0] u0_col_out_959;
wire [105:0] u0_col_out_960;
wire [105:0] u0_col_out_961;
wire [105:0] u0_col_out_962;
wire [105:0] u0_col_out_963;
wire [105:0] u0_col_out_964;
wire [105:0] u0_col_out_965;
wire [105:0] u0_col_out_966;
wire [105:0] u0_col_out_967;
wire [105:0] u0_col_out_968;
wire [105:0] u0_col_out_969;
wire [105:0] u0_col_out_970;
wire [105:0] u0_col_out_971;
wire [105:0] u0_col_out_972;
wire [105:0] u0_col_out_973;
wire [105:0] u0_col_out_974;
wire [105:0] u0_col_out_975;
wire [105:0] u0_col_out_976;
wire [105:0] u0_col_out_977;
wire [105:0] u0_col_out_978;
wire [105:0] u0_col_out_979;
wire [105:0] u0_col_out_980;
wire [105:0] u0_col_out_981;
wire [105:0] u0_col_out_982;
wire [105:0] u0_col_out_983;
wire [105:0] u0_col_out_984;
wire [105:0] u0_col_out_985;
wire [105:0] u0_col_out_986;
wire [105:0] u0_col_out_987;
wire [105:0] u0_col_out_988;
wire [105:0] u0_col_out_989;
wire [105:0] u0_col_out_990;
wire [105:0] u0_col_out_991;
wire [105:0] u0_col_out_992;
wire [105:0] u0_col_out_993;
wire [105:0] u0_col_out_994;
wire [105:0] u0_col_out_995;
wire [105:0] u0_col_out_996;
wire [105:0] u0_col_out_997;
wire [105:0] u0_col_out_998;
wire [105:0] u0_col_out_999;
wire [105:0] u0_col_out_1000;
wire [105:0] u0_col_out_1001;
wire [105:0] u0_col_out_1002;
wire [105:0] u0_col_out_1003;
wire [105:0] u0_col_out_1004;
wire [105:0] u0_col_out_1005;
wire [105:0] u0_col_out_1006;
wire [105:0] u0_col_out_1007;
wire [105:0] u0_col_out_1008;
wire [105:0] u0_col_out_1009;
wire [105:0] u0_col_out_1010;
wire [105:0] u0_col_out_1011;
wire [105:0] u0_col_out_1012;
wire [105:0] u0_col_out_1013;
wire [105:0] u0_col_out_1014;
wire [105:0] u0_col_out_1015;
wire [105:0] u0_col_out_1016;
wire [105:0] u0_col_out_1017;
wire [105:0] u0_col_out_1018;
wire [105:0] u0_col_out_1019;
wire [105:0] u0_col_out_1020;
wire [105:0] u0_col_out_1021;
wire [105:0] u0_col_out_1022;
wire [105:0] u0_col_out_1023;
wire [105:0] u0_col_out_1024;
wire [105:0] u0_col_out_1025;
wire [105:0] u0_col_out_1026;
wire [105:0] u0_col_out_1027;
wire [105:0] u0_col_out_1028;
wire [105:0] u0_col_out_1029;
wire [105:0] u0_col_out_1030;
wire [105:0] u0_col_out_1031;
wire [105:0] u0_col_out_1032;
wire [105:0] u0_col_out_1033;
wire [105:0] u0_col_out_1034;
wire [105:0] u0_col_out_1035;
wire [105:0] u0_col_out_1036;
wire [105:0] u0_col_out_1037;
wire [105:0] u0_col_out_1038;
wire [105:0] u0_col_out_1039;
wire [105:0] u0_col_out_1040;
wire [105:0] u0_col_out_1041;
wire [105:0] u0_col_out_1042;
wire [105:0] u0_col_out_1043;
wire [105:0] u0_col_out_1044;
wire [105:0] u0_col_out_1045;
wire [105:0] u0_col_out_1046;
wire [105:0] u0_col_out_1047;
wire [105:0] u0_col_out_1048;
wire [105:0] u0_col_out_1049;
wire [105:0] u0_col_out_1050;
wire [105:0] u0_col_out_1051;
wire [105:0] u0_col_out_1052;
wire [105:0] u0_col_out_1053;
wire [105:0] u0_col_out_1054;
wire [105:0] u0_col_out_1055;
wire [105:0] u0_col_out_1056;
wire [105:0] u0_col_out_1057;
wire [105:0] u0_col_out_1058;
wire [105:0] u0_col_out_1059;
wire [105:0] u0_col_out_1060;
wire [105:0] u0_col_out_1061;
wire [105:0] u0_col_out_1062;
wire [105:0] u0_col_out_1063;
wire [105:0] u0_col_out_1064;
wire [105:0] u0_col_out_1065;
wire [105:0] u0_col_out_1066;
wire [105:0] u0_col_out_1067;
wire [105:0] u0_col_out_1068;
wire [105:0] u0_col_out_1069;
wire [105:0] u0_col_out_1070;
wire [105:0] u0_col_out_1071;
wire [105:0] u0_col_out_1072;
wire [105:0] u0_col_out_1073;
wire [105:0] u0_col_out_1074;
wire [105:0] u0_col_out_1075;
wire [105:0] u0_col_out_1076;
wire [105:0] u0_col_out_1077;
wire [105:0] u0_col_out_1078;
wire [105:0] u0_col_out_1079;
wire [105:0] u0_col_out_1080;
wire [105:0] u0_col_out_1081;
wire [105:0] u0_col_out_1082;
wire [105:0] u0_col_out_1083;
wire [105:0] u0_col_out_1084;
wire [105:0] u0_col_out_1085;
wire [105:0] u0_col_out_1086;
wire [105:0] u0_col_out_1087;
wire [105:0] u0_col_out_1088;
wire [105:0] u0_col_out_1089;
wire [105:0] u0_col_out_1090;
wire [105:0] u0_col_out_1091;
wire [105:0] u0_col_out_1092;
wire [105:0] u0_col_out_1093;
wire [105:0] u0_col_out_1094;
wire [105:0] u0_col_out_1095;
wire [105:0] u0_col_out_1096;
wire [105:0] u0_col_out_1097;
wire [105:0] u0_col_out_1098;
wire [105:0] u0_col_out_1099;
wire [105:0] u0_col_out_1100;
wire [105:0] u0_col_out_1101;
wire [105:0] u0_col_out_1102;
wire [105:0] u0_col_out_1103;
wire [105:0] u0_col_out_1104;
wire [105:0] u0_col_out_1105;
wire [105:0] u0_col_out_1106;
wire [105:0] u0_col_out_1107;
wire [105:0] u0_col_out_1108;
wire [105:0] u0_col_out_1109;
wire [105:0] u0_col_out_1110;
wire [105:0] u0_col_out_1111;
wire [105:0] u0_col_out_1112;
wire [105:0] u0_col_out_1113;
wire [105:0] u0_col_out_1114;
wire [105:0] u0_col_out_1115;
wire [105:0] u0_col_out_1116;
wire [105:0] u0_col_out_1117;
wire [105:0] u0_col_out_1118;
wire [105:0] u0_col_out_1119;
wire [105:0] u0_col_out_1120;
wire [105:0] u0_col_out_1121;
wire [105:0] u0_col_out_1122;
wire [105:0] u0_col_out_1123;
wire [105:0] u0_col_out_1124;
wire [105:0] u0_col_out_1125;
wire [105:0] u0_col_out_1126;
wire [105:0] u0_col_out_1127;
wire [105:0] u0_col_out_1128;
wire [105:0] u0_col_out_1129;
wire [105:0] u0_col_out_1130;
wire [105:0] u0_col_out_1131;
wire [105:0] u0_col_out_1132;
wire [105:0] u0_col_out_1133;
wire [105:0] u0_col_out_1134;
wire [105:0] u0_col_out_1135;
wire [105:0] u0_col_out_1136;
wire [105:0] u0_col_out_1137;
wire [105:0] u0_col_out_1138;
wire [105:0] u0_col_out_1139;
wire [105:0] u0_col_out_1140;
wire [105:0] u0_col_out_1141;
wire [105:0] u0_col_out_1142;
wire [105:0] u0_col_out_1143;
wire [105:0] u0_col_out_1144;
wire [105:0] u0_col_out_1145;
wire [105:0] u0_col_out_1146;
wire [105:0] u0_col_out_1147;
wire [105:0] u0_col_out_1148;
wire [105:0] u0_col_out_1149;
wire [105:0] u0_col_out_1150;
wire [105:0] u0_col_out_1151;
wire [105:0] u0_col_out_1152;
wire [105:0] u0_col_out_1153;
wire [105:0] u0_col_out_1154;
wire [105:0] u0_col_out_1155;
wire [105:0] u0_col_out_1156;
wire [105:0] u0_col_out_1157;
wire [105:0] u0_col_out_1158;
wire [105:0] u0_col_out_1159;
wire [105:0] u0_col_out_1160;
wire [105:0] u0_col_out_1161;
wire [105:0] u0_col_out_1162;
wire [105:0] u0_col_out_1163;
wire [105:0] u0_col_out_1164;
wire [105:0] u0_col_out_1165;
wire [105:0] u0_col_out_1166;
wire [105:0] u0_col_out_1167;
wire [105:0] u0_col_out_1168;
wire [105:0] u0_col_out_1169;
wire [105:0] u0_col_out_1170;
wire [105:0] u0_col_out_1171;
wire [105:0] u0_col_out_1172;
wire [105:0] u0_col_out_1173;
wire [105:0] u0_col_out_1174;
wire [105:0] u0_col_out_1175;
wire [105:0] u0_col_out_1176;
wire [105:0] u0_col_out_1177;
wire [105:0] u0_col_out_1178;
wire [105:0] u0_col_out_1179;
wire [105:0] u0_col_out_1180;
wire [105:0] u0_col_out_1181;
wire [105:0] u0_col_out_1182;
wire [105:0] u0_col_out_1183;
wire [105:0] u0_col_out_1184;
wire [105:0] u0_col_out_1185;
wire [105:0] u0_col_out_1186;
wire [105:0] u0_col_out_1187;
wire [105:0] u0_col_out_1188;
wire [105:0] u0_col_out_1189;
wire [105:0] u0_col_out_1190;
wire [105:0] u0_col_out_1191;
wire [105:0] u0_col_out_1192;
wire [105:0] u0_col_out_1193;
wire [105:0] u0_col_out_1194;
wire [105:0] u0_col_out_1195;
wire [105:0] u0_col_out_1196;
wire [105:0] u0_col_out_1197;
wire [105:0] u0_col_out_1198;
wire [105:0] u0_col_out_1199;
wire [105:0] u0_col_out_1200;
wire [105:0] u0_col_out_1201;
wire [105:0] u0_col_out_1202;
wire [105:0] u0_col_out_1203;
wire [105:0] u0_col_out_1204;
wire [105:0] u0_col_out_1205;
wire [105:0] u0_col_out_1206;
wire [105:0] u0_col_out_1207;
wire [105:0] u0_col_out_1208;
wire [105:0] u0_col_out_1209;
wire [105:0] u0_col_out_1210;
wire [105:0] u0_col_out_1211;
wire [105:0] u0_col_out_1212;
wire [105:0] u0_col_out_1213;
wire [105:0] u0_col_out_1214;
wire [105:0] u0_col_out_1215;
wire [105:0] u0_col_out_1216;
wire [105:0] u0_col_out_1217;
wire [105:0] u0_col_out_1218;
wire [105:0] u0_col_out_1219;
wire [105:0] u0_col_out_1220;
wire [105:0] u0_col_out_1221;
wire [105:0] u0_col_out_1222;
wire [105:0] u0_col_out_1223;
wire [105:0] u0_col_out_1224;
wire [105:0] u0_col_out_1225;
wire [105:0] u0_col_out_1226;
wire [105:0] u0_col_out_1227;
wire [105:0] u0_col_out_1228;
wire [105:0] u0_col_out_1229;
wire [105:0] u0_col_out_1230;
wire [105:0] u0_col_out_1231;
wire [105:0] u0_col_out_1232;
wire [105:0] u0_col_out_1233;
wire [105:0] u0_col_out_1234;
wire [105:0] u0_col_out_1235;
wire [105:0] u0_col_out_1236;
wire [105:0] u0_col_out_1237;
wire [105:0] u0_col_out_1238;
wire [105:0] u0_col_out_1239;
wire [105:0] u0_col_out_1240;
wire [105:0] u0_col_out_1241;
wire [105:0] u0_col_out_1242;
wire [105:0] u0_col_out_1243;
wire [105:0] u0_col_out_1244;
wire [105:0] u0_col_out_1245;
wire [105:0] u0_col_out_1246;
wire [105:0] u0_col_out_1247;
wire [105:0] u0_col_out_1248;
wire [105:0] u0_col_out_1249;
wire [105:0] u0_col_out_1250;
wire [105:0] u0_col_out_1251;
wire [105:0] u0_col_out_1252;
wire [105:0] u0_col_out_1253;
wire [105:0] u0_col_out_1254;
wire [105:0] u0_col_out_1255;
wire [105:0] u0_col_out_1256;
wire [105:0] u0_col_out_1257;
wire [105:0] u0_col_out_1258;
wire [105:0] u0_col_out_1259;
wire [105:0] u0_col_out_1260;
wire [105:0] u0_col_out_1261;
wire [105:0] u0_col_out_1262;
wire [105:0] u0_col_out_1263;
wire [105:0] u0_col_out_1264;
wire [105:0] u0_col_out_1265;
wire [105:0] u0_col_out_1266;
wire [105:0] u0_col_out_1267;
wire [105:0] u0_col_out_1268;
wire [105:0] u0_col_out_1269;
wire [105:0] u0_col_out_1270;
wire [105:0] u0_col_out_1271;
wire [105:0] u0_col_out_1272;
wire [105:0] u0_col_out_1273;
wire [105:0] u0_col_out_1274;
wire [105:0] u0_col_out_1275;
wire [105:0] u0_col_out_1276;
wire [105:0] u0_col_out_1277;
wire [105:0] u0_col_out_1278;
wire [105:0] u0_col_out_1279;
wire [105:0] u0_col_out_1280;
wire [105:0] u0_col_out_1281;
wire [105:0] u0_col_out_1282;
wire [105:0] u0_col_out_1283;
wire [105:0] u0_col_out_1284;
wire [105:0] u0_col_out_1285;
wire [105:0] u0_col_out_1286;
wire [105:0] u0_col_out_1287;


xpb_first u0_xpb_first
(
    .data_in0(reg_intermediate0[1287:1024]),
    .data_in1(reg_intermediate1[1287:1024]),


    .col_out_0(u0_col_out_0),
    .col_out_1(u0_col_out_1),
    .col_out_2(u0_col_out_2),
    .col_out_3(u0_col_out_3),
    .col_out_4(u0_col_out_4),
    .col_out_5(u0_col_out_5),
    .col_out_6(u0_col_out_6),
    .col_out_7(u0_col_out_7),
    .col_out_8(u0_col_out_8),
    .col_out_9(u0_col_out_9),
    .col_out_10(u0_col_out_10),
    .col_out_11(u0_col_out_11),
    .col_out_12(u0_col_out_12),
    .col_out_13(u0_col_out_13),
    .col_out_14(u0_col_out_14),
    .col_out_15(u0_col_out_15),
    .col_out_16(u0_col_out_16),
    .col_out_17(u0_col_out_17),
    .col_out_18(u0_col_out_18),
    .col_out_19(u0_col_out_19),
    .col_out_20(u0_col_out_20),
    .col_out_21(u0_col_out_21),
    .col_out_22(u0_col_out_22),
    .col_out_23(u0_col_out_23),
    .col_out_24(u0_col_out_24),
    .col_out_25(u0_col_out_25),
    .col_out_26(u0_col_out_26),
    .col_out_27(u0_col_out_27),
    .col_out_28(u0_col_out_28),
    .col_out_29(u0_col_out_29),
    .col_out_30(u0_col_out_30),
    .col_out_31(u0_col_out_31),
    .col_out_32(u0_col_out_32),
    .col_out_33(u0_col_out_33),
    .col_out_34(u0_col_out_34),
    .col_out_35(u0_col_out_35),
    .col_out_36(u0_col_out_36),
    .col_out_37(u0_col_out_37),
    .col_out_38(u0_col_out_38),
    .col_out_39(u0_col_out_39),
    .col_out_40(u0_col_out_40),
    .col_out_41(u0_col_out_41),
    .col_out_42(u0_col_out_42),
    .col_out_43(u0_col_out_43),
    .col_out_44(u0_col_out_44),
    .col_out_45(u0_col_out_45),
    .col_out_46(u0_col_out_46),
    .col_out_47(u0_col_out_47),
    .col_out_48(u0_col_out_48),
    .col_out_49(u0_col_out_49),
    .col_out_50(u0_col_out_50),
    .col_out_51(u0_col_out_51),
    .col_out_52(u0_col_out_52),
    .col_out_53(u0_col_out_53),
    .col_out_54(u0_col_out_54),
    .col_out_55(u0_col_out_55),
    .col_out_56(u0_col_out_56),
    .col_out_57(u0_col_out_57),
    .col_out_58(u0_col_out_58),
    .col_out_59(u0_col_out_59),
    .col_out_60(u0_col_out_60),
    .col_out_61(u0_col_out_61),
    .col_out_62(u0_col_out_62),
    .col_out_63(u0_col_out_63),
    .col_out_64(u0_col_out_64),
    .col_out_65(u0_col_out_65),
    .col_out_66(u0_col_out_66),
    .col_out_67(u0_col_out_67),
    .col_out_68(u0_col_out_68),
    .col_out_69(u0_col_out_69),
    .col_out_70(u0_col_out_70),
    .col_out_71(u0_col_out_71),
    .col_out_72(u0_col_out_72),
    .col_out_73(u0_col_out_73),
    .col_out_74(u0_col_out_74),
    .col_out_75(u0_col_out_75),
    .col_out_76(u0_col_out_76),
    .col_out_77(u0_col_out_77),
    .col_out_78(u0_col_out_78),
    .col_out_79(u0_col_out_79),
    .col_out_80(u0_col_out_80),
    .col_out_81(u0_col_out_81),
    .col_out_82(u0_col_out_82),
    .col_out_83(u0_col_out_83),
    .col_out_84(u0_col_out_84),
    .col_out_85(u0_col_out_85),
    .col_out_86(u0_col_out_86),
    .col_out_87(u0_col_out_87),
    .col_out_88(u0_col_out_88),
    .col_out_89(u0_col_out_89),
    .col_out_90(u0_col_out_90),
    .col_out_91(u0_col_out_91),
    .col_out_92(u0_col_out_92),
    .col_out_93(u0_col_out_93),
    .col_out_94(u0_col_out_94),
    .col_out_95(u0_col_out_95),
    .col_out_96(u0_col_out_96),
    .col_out_97(u0_col_out_97),
    .col_out_98(u0_col_out_98),
    .col_out_99(u0_col_out_99),
    .col_out_100(u0_col_out_100),
    .col_out_101(u0_col_out_101),
    .col_out_102(u0_col_out_102),
    .col_out_103(u0_col_out_103),
    .col_out_104(u0_col_out_104),
    .col_out_105(u0_col_out_105),
    .col_out_106(u0_col_out_106),
    .col_out_107(u0_col_out_107),
    .col_out_108(u0_col_out_108),
    .col_out_109(u0_col_out_109),
    .col_out_110(u0_col_out_110),
    .col_out_111(u0_col_out_111),
    .col_out_112(u0_col_out_112),
    .col_out_113(u0_col_out_113),
    .col_out_114(u0_col_out_114),
    .col_out_115(u0_col_out_115),
    .col_out_116(u0_col_out_116),
    .col_out_117(u0_col_out_117),
    .col_out_118(u0_col_out_118),
    .col_out_119(u0_col_out_119),
    .col_out_120(u0_col_out_120),
    .col_out_121(u0_col_out_121),
    .col_out_122(u0_col_out_122),
    .col_out_123(u0_col_out_123),
    .col_out_124(u0_col_out_124),
    .col_out_125(u0_col_out_125),
    .col_out_126(u0_col_out_126),
    .col_out_127(u0_col_out_127),
    .col_out_128(u0_col_out_128),
    .col_out_129(u0_col_out_129),
    .col_out_130(u0_col_out_130),
    .col_out_131(u0_col_out_131),
    .col_out_132(u0_col_out_132),
    .col_out_133(u0_col_out_133),
    .col_out_134(u0_col_out_134),
    .col_out_135(u0_col_out_135),
    .col_out_136(u0_col_out_136),
    .col_out_137(u0_col_out_137),
    .col_out_138(u0_col_out_138),
    .col_out_139(u0_col_out_139),
    .col_out_140(u0_col_out_140),
    .col_out_141(u0_col_out_141),
    .col_out_142(u0_col_out_142),
    .col_out_143(u0_col_out_143),
    .col_out_144(u0_col_out_144),
    .col_out_145(u0_col_out_145),
    .col_out_146(u0_col_out_146),
    .col_out_147(u0_col_out_147),
    .col_out_148(u0_col_out_148),
    .col_out_149(u0_col_out_149),
    .col_out_150(u0_col_out_150),
    .col_out_151(u0_col_out_151),
    .col_out_152(u0_col_out_152),
    .col_out_153(u0_col_out_153),
    .col_out_154(u0_col_out_154),
    .col_out_155(u0_col_out_155),
    .col_out_156(u0_col_out_156),
    .col_out_157(u0_col_out_157),
    .col_out_158(u0_col_out_158),
    .col_out_159(u0_col_out_159),
    .col_out_160(u0_col_out_160),
    .col_out_161(u0_col_out_161),
    .col_out_162(u0_col_out_162),
    .col_out_163(u0_col_out_163),
    .col_out_164(u0_col_out_164),
    .col_out_165(u0_col_out_165),
    .col_out_166(u0_col_out_166),
    .col_out_167(u0_col_out_167),
    .col_out_168(u0_col_out_168),
    .col_out_169(u0_col_out_169),
    .col_out_170(u0_col_out_170),
    .col_out_171(u0_col_out_171),
    .col_out_172(u0_col_out_172),
    .col_out_173(u0_col_out_173),
    .col_out_174(u0_col_out_174),
    .col_out_175(u0_col_out_175),
    .col_out_176(u0_col_out_176),
    .col_out_177(u0_col_out_177),
    .col_out_178(u0_col_out_178),
    .col_out_179(u0_col_out_179),
    .col_out_180(u0_col_out_180),
    .col_out_181(u0_col_out_181),
    .col_out_182(u0_col_out_182),
    .col_out_183(u0_col_out_183),
    .col_out_184(u0_col_out_184),
    .col_out_185(u0_col_out_185),
    .col_out_186(u0_col_out_186),
    .col_out_187(u0_col_out_187),
    .col_out_188(u0_col_out_188),
    .col_out_189(u0_col_out_189),
    .col_out_190(u0_col_out_190),
    .col_out_191(u0_col_out_191),
    .col_out_192(u0_col_out_192),
    .col_out_193(u0_col_out_193),
    .col_out_194(u0_col_out_194),
    .col_out_195(u0_col_out_195),
    .col_out_196(u0_col_out_196),
    .col_out_197(u0_col_out_197),
    .col_out_198(u0_col_out_198),
    .col_out_199(u0_col_out_199),
    .col_out_200(u0_col_out_200),
    .col_out_201(u0_col_out_201),
    .col_out_202(u0_col_out_202),
    .col_out_203(u0_col_out_203),
    .col_out_204(u0_col_out_204),
    .col_out_205(u0_col_out_205),
    .col_out_206(u0_col_out_206),
    .col_out_207(u0_col_out_207),
    .col_out_208(u0_col_out_208),
    .col_out_209(u0_col_out_209),
    .col_out_210(u0_col_out_210),
    .col_out_211(u0_col_out_211),
    .col_out_212(u0_col_out_212),
    .col_out_213(u0_col_out_213),
    .col_out_214(u0_col_out_214),
    .col_out_215(u0_col_out_215),
    .col_out_216(u0_col_out_216),
    .col_out_217(u0_col_out_217),
    .col_out_218(u0_col_out_218),
    .col_out_219(u0_col_out_219),
    .col_out_220(u0_col_out_220),
    .col_out_221(u0_col_out_221),
    .col_out_222(u0_col_out_222),
    .col_out_223(u0_col_out_223),
    .col_out_224(u0_col_out_224),
    .col_out_225(u0_col_out_225),
    .col_out_226(u0_col_out_226),
    .col_out_227(u0_col_out_227),
    .col_out_228(u0_col_out_228),
    .col_out_229(u0_col_out_229),
    .col_out_230(u0_col_out_230),
    .col_out_231(u0_col_out_231),
    .col_out_232(u0_col_out_232),
    .col_out_233(u0_col_out_233),
    .col_out_234(u0_col_out_234),
    .col_out_235(u0_col_out_235),
    .col_out_236(u0_col_out_236),
    .col_out_237(u0_col_out_237),
    .col_out_238(u0_col_out_238),
    .col_out_239(u0_col_out_239),
    .col_out_240(u0_col_out_240),
    .col_out_241(u0_col_out_241),
    .col_out_242(u0_col_out_242),
    .col_out_243(u0_col_out_243),
    .col_out_244(u0_col_out_244),
    .col_out_245(u0_col_out_245),
    .col_out_246(u0_col_out_246),
    .col_out_247(u0_col_out_247),
    .col_out_248(u0_col_out_248),
    .col_out_249(u0_col_out_249),
    .col_out_250(u0_col_out_250),
    .col_out_251(u0_col_out_251),
    .col_out_252(u0_col_out_252),
    .col_out_253(u0_col_out_253),
    .col_out_254(u0_col_out_254),
    .col_out_255(u0_col_out_255),
    .col_out_256(u0_col_out_256),
    .col_out_257(u0_col_out_257),
    .col_out_258(u0_col_out_258),
    .col_out_259(u0_col_out_259),
    .col_out_260(u0_col_out_260),
    .col_out_261(u0_col_out_261),
    .col_out_262(u0_col_out_262),
    .col_out_263(u0_col_out_263),
    .col_out_264(u0_col_out_264),
    .col_out_265(u0_col_out_265),
    .col_out_266(u0_col_out_266),
    .col_out_267(u0_col_out_267),
    .col_out_268(u0_col_out_268),
    .col_out_269(u0_col_out_269),
    .col_out_270(u0_col_out_270),
    .col_out_271(u0_col_out_271),
    .col_out_272(u0_col_out_272),
    .col_out_273(u0_col_out_273),
    .col_out_274(u0_col_out_274),
    .col_out_275(u0_col_out_275),
    .col_out_276(u0_col_out_276),
    .col_out_277(u0_col_out_277),
    .col_out_278(u0_col_out_278),
    .col_out_279(u0_col_out_279),
    .col_out_280(u0_col_out_280),
    .col_out_281(u0_col_out_281),
    .col_out_282(u0_col_out_282),
    .col_out_283(u0_col_out_283),
    .col_out_284(u0_col_out_284),
    .col_out_285(u0_col_out_285),
    .col_out_286(u0_col_out_286),
    .col_out_287(u0_col_out_287),
    .col_out_288(u0_col_out_288),
    .col_out_289(u0_col_out_289),
    .col_out_290(u0_col_out_290),
    .col_out_291(u0_col_out_291),
    .col_out_292(u0_col_out_292),
    .col_out_293(u0_col_out_293),
    .col_out_294(u0_col_out_294),
    .col_out_295(u0_col_out_295),
    .col_out_296(u0_col_out_296),
    .col_out_297(u0_col_out_297),
    .col_out_298(u0_col_out_298),
    .col_out_299(u0_col_out_299),
    .col_out_300(u0_col_out_300),
    .col_out_301(u0_col_out_301),
    .col_out_302(u0_col_out_302),
    .col_out_303(u0_col_out_303),
    .col_out_304(u0_col_out_304),
    .col_out_305(u0_col_out_305),
    .col_out_306(u0_col_out_306),
    .col_out_307(u0_col_out_307),
    .col_out_308(u0_col_out_308),
    .col_out_309(u0_col_out_309),
    .col_out_310(u0_col_out_310),
    .col_out_311(u0_col_out_311),
    .col_out_312(u0_col_out_312),
    .col_out_313(u0_col_out_313),
    .col_out_314(u0_col_out_314),
    .col_out_315(u0_col_out_315),
    .col_out_316(u0_col_out_316),
    .col_out_317(u0_col_out_317),
    .col_out_318(u0_col_out_318),
    .col_out_319(u0_col_out_319),
    .col_out_320(u0_col_out_320),
    .col_out_321(u0_col_out_321),
    .col_out_322(u0_col_out_322),
    .col_out_323(u0_col_out_323),
    .col_out_324(u0_col_out_324),
    .col_out_325(u0_col_out_325),
    .col_out_326(u0_col_out_326),
    .col_out_327(u0_col_out_327),
    .col_out_328(u0_col_out_328),
    .col_out_329(u0_col_out_329),
    .col_out_330(u0_col_out_330),
    .col_out_331(u0_col_out_331),
    .col_out_332(u0_col_out_332),
    .col_out_333(u0_col_out_333),
    .col_out_334(u0_col_out_334),
    .col_out_335(u0_col_out_335),
    .col_out_336(u0_col_out_336),
    .col_out_337(u0_col_out_337),
    .col_out_338(u0_col_out_338),
    .col_out_339(u0_col_out_339),
    .col_out_340(u0_col_out_340),
    .col_out_341(u0_col_out_341),
    .col_out_342(u0_col_out_342),
    .col_out_343(u0_col_out_343),
    .col_out_344(u0_col_out_344),
    .col_out_345(u0_col_out_345),
    .col_out_346(u0_col_out_346),
    .col_out_347(u0_col_out_347),
    .col_out_348(u0_col_out_348),
    .col_out_349(u0_col_out_349),
    .col_out_350(u0_col_out_350),
    .col_out_351(u0_col_out_351),
    .col_out_352(u0_col_out_352),
    .col_out_353(u0_col_out_353),
    .col_out_354(u0_col_out_354),
    .col_out_355(u0_col_out_355),
    .col_out_356(u0_col_out_356),
    .col_out_357(u0_col_out_357),
    .col_out_358(u0_col_out_358),
    .col_out_359(u0_col_out_359),
    .col_out_360(u0_col_out_360),
    .col_out_361(u0_col_out_361),
    .col_out_362(u0_col_out_362),
    .col_out_363(u0_col_out_363),
    .col_out_364(u0_col_out_364),
    .col_out_365(u0_col_out_365),
    .col_out_366(u0_col_out_366),
    .col_out_367(u0_col_out_367),
    .col_out_368(u0_col_out_368),
    .col_out_369(u0_col_out_369),
    .col_out_370(u0_col_out_370),
    .col_out_371(u0_col_out_371),
    .col_out_372(u0_col_out_372),
    .col_out_373(u0_col_out_373),
    .col_out_374(u0_col_out_374),
    .col_out_375(u0_col_out_375),
    .col_out_376(u0_col_out_376),
    .col_out_377(u0_col_out_377),
    .col_out_378(u0_col_out_378),
    .col_out_379(u0_col_out_379),
    .col_out_380(u0_col_out_380),
    .col_out_381(u0_col_out_381),
    .col_out_382(u0_col_out_382),
    .col_out_383(u0_col_out_383),
    .col_out_384(u0_col_out_384),
    .col_out_385(u0_col_out_385),
    .col_out_386(u0_col_out_386),
    .col_out_387(u0_col_out_387),
    .col_out_388(u0_col_out_388),
    .col_out_389(u0_col_out_389),
    .col_out_390(u0_col_out_390),
    .col_out_391(u0_col_out_391),
    .col_out_392(u0_col_out_392),
    .col_out_393(u0_col_out_393),
    .col_out_394(u0_col_out_394),
    .col_out_395(u0_col_out_395),
    .col_out_396(u0_col_out_396),
    .col_out_397(u0_col_out_397),
    .col_out_398(u0_col_out_398),
    .col_out_399(u0_col_out_399),
    .col_out_400(u0_col_out_400),
    .col_out_401(u0_col_out_401),
    .col_out_402(u0_col_out_402),
    .col_out_403(u0_col_out_403),
    .col_out_404(u0_col_out_404),
    .col_out_405(u0_col_out_405),
    .col_out_406(u0_col_out_406),
    .col_out_407(u0_col_out_407),
    .col_out_408(u0_col_out_408),
    .col_out_409(u0_col_out_409),
    .col_out_410(u0_col_out_410),
    .col_out_411(u0_col_out_411),
    .col_out_412(u0_col_out_412),
    .col_out_413(u0_col_out_413),
    .col_out_414(u0_col_out_414),
    .col_out_415(u0_col_out_415),
    .col_out_416(u0_col_out_416),
    .col_out_417(u0_col_out_417),
    .col_out_418(u0_col_out_418),
    .col_out_419(u0_col_out_419),
    .col_out_420(u0_col_out_420),
    .col_out_421(u0_col_out_421),
    .col_out_422(u0_col_out_422),
    .col_out_423(u0_col_out_423),
    .col_out_424(u0_col_out_424),
    .col_out_425(u0_col_out_425),
    .col_out_426(u0_col_out_426),
    .col_out_427(u0_col_out_427),
    .col_out_428(u0_col_out_428),
    .col_out_429(u0_col_out_429),
    .col_out_430(u0_col_out_430),
    .col_out_431(u0_col_out_431),
    .col_out_432(u0_col_out_432),
    .col_out_433(u0_col_out_433),
    .col_out_434(u0_col_out_434),
    .col_out_435(u0_col_out_435),
    .col_out_436(u0_col_out_436),
    .col_out_437(u0_col_out_437),
    .col_out_438(u0_col_out_438),
    .col_out_439(u0_col_out_439),
    .col_out_440(u0_col_out_440),
    .col_out_441(u0_col_out_441),
    .col_out_442(u0_col_out_442),
    .col_out_443(u0_col_out_443),
    .col_out_444(u0_col_out_444),
    .col_out_445(u0_col_out_445),
    .col_out_446(u0_col_out_446),
    .col_out_447(u0_col_out_447),
    .col_out_448(u0_col_out_448),
    .col_out_449(u0_col_out_449),
    .col_out_450(u0_col_out_450),
    .col_out_451(u0_col_out_451),
    .col_out_452(u0_col_out_452),
    .col_out_453(u0_col_out_453),
    .col_out_454(u0_col_out_454),
    .col_out_455(u0_col_out_455),
    .col_out_456(u0_col_out_456),
    .col_out_457(u0_col_out_457),
    .col_out_458(u0_col_out_458),
    .col_out_459(u0_col_out_459),
    .col_out_460(u0_col_out_460),
    .col_out_461(u0_col_out_461),
    .col_out_462(u0_col_out_462),
    .col_out_463(u0_col_out_463),
    .col_out_464(u0_col_out_464),
    .col_out_465(u0_col_out_465),
    .col_out_466(u0_col_out_466),
    .col_out_467(u0_col_out_467),
    .col_out_468(u0_col_out_468),
    .col_out_469(u0_col_out_469),
    .col_out_470(u0_col_out_470),
    .col_out_471(u0_col_out_471),
    .col_out_472(u0_col_out_472),
    .col_out_473(u0_col_out_473),
    .col_out_474(u0_col_out_474),
    .col_out_475(u0_col_out_475),
    .col_out_476(u0_col_out_476),
    .col_out_477(u0_col_out_477),
    .col_out_478(u0_col_out_478),
    .col_out_479(u0_col_out_479),
    .col_out_480(u0_col_out_480),
    .col_out_481(u0_col_out_481),
    .col_out_482(u0_col_out_482),
    .col_out_483(u0_col_out_483),
    .col_out_484(u0_col_out_484),
    .col_out_485(u0_col_out_485),
    .col_out_486(u0_col_out_486),
    .col_out_487(u0_col_out_487),
    .col_out_488(u0_col_out_488),
    .col_out_489(u0_col_out_489),
    .col_out_490(u0_col_out_490),
    .col_out_491(u0_col_out_491),
    .col_out_492(u0_col_out_492),
    .col_out_493(u0_col_out_493),
    .col_out_494(u0_col_out_494),
    .col_out_495(u0_col_out_495),
    .col_out_496(u0_col_out_496),
    .col_out_497(u0_col_out_497),
    .col_out_498(u0_col_out_498),
    .col_out_499(u0_col_out_499),
    .col_out_500(u0_col_out_500),
    .col_out_501(u0_col_out_501),
    .col_out_502(u0_col_out_502),
    .col_out_503(u0_col_out_503),
    .col_out_504(u0_col_out_504),
    .col_out_505(u0_col_out_505),
    .col_out_506(u0_col_out_506),
    .col_out_507(u0_col_out_507),
    .col_out_508(u0_col_out_508),
    .col_out_509(u0_col_out_509),
    .col_out_510(u0_col_out_510),
    .col_out_511(u0_col_out_511),
    .col_out_512(u0_col_out_512),
    .col_out_513(u0_col_out_513),
    .col_out_514(u0_col_out_514),
    .col_out_515(u0_col_out_515),
    .col_out_516(u0_col_out_516),
    .col_out_517(u0_col_out_517),
    .col_out_518(u0_col_out_518),
    .col_out_519(u0_col_out_519),
    .col_out_520(u0_col_out_520),
    .col_out_521(u0_col_out_521),
    .col_out_522(u0_col_out_522),
    .col_out_523(u0_col_out_523),
    .col_out_524(u0_col_out_524),
    .col_out_525(u0_col_out_525),
    .col_out_526(u0_col_out_526),
    .col_out_527(u0_col_out_527),
    .col_out_528(u0_col_out_528),
    .col_out_529(u0_col_out_529),
    .col_out_530(u0_col_out_530),
    .col_out_531(u0_col_out_531),
    .col_out_532(u0_col_out_532),
    .col_out_533(u0_col_out_533),
    .col_out_534(u0_col_out_534),
    .col_out_535(u0_col_out_535),
    .col_out_536(u0_col_out_536),
    .col_out_537(u0_col_out_537),
    .col_out_538(u0_col_out_538),
    .col_out_539(u0_col_out_539),
    .col_out_540(u0_col_out_540),
    .col_out_541(u0_col_out_541),
    .col_out_542(u0_col_out_542),
    .col_out_543(u0_col_out_543),
    .col_out_544(u0_col_out_544),
    .col_out_545(u0_col_out_545),
    .col_out_546(u0_col_out_546),
    .col_out_547(u0_col_out_547),
    .col_out_548(u0_col_out_548),
    .col_out_549(u0_col_out_549),
    .col_out_550(u0_col_out_550),
    .col_out_551(u0_col_out_551),
    .col_out_552(u0_col_out_552),
    .col_out_553(u0_col_out_553),
    .col_out_554(u0_col_out_554),
    .col_out_555(u0_col_out_555),
    .col_out_556(u0_col_out_556),
    .col_out_557(u0_col_out_557),
    .col_out_558(u0_col_out_558),
    .col_out_559(u0_col_out_559),
    .col_out_560(u0_col_out_560),
    .col_out_561(u0_col_out_561),
    .col_out_562(u0_col_out_562),
    .col_out_563(u0_col_out_563),
    .col_out_564(u0_col_out_564),
    .col_out_565(u0_col_out_565),
    .col_out_566(u0_col_out_566),
    .col_out_567(u0_col_out_567),
    .col_out_568(u0_col_out_568),
    .col_out_569(u0_col_out_569),
    .col_out_570(u0_col_out_570),
    .col_out_571(u0_col_out_571),
    .col_out_572(u0_col_out_572),
    .col_out_573(u0_col_out_573),
    .col_out_574(u0_col_out_574),
    .col_out_575(u0_col_out_575),
    .col_out_576(u0_col_out_576),
    .col_out_577(u0_col_out_577),
    .col_out_578(u0_col_out_578),
    .col_out_579(u0_col_out_579),
    .col_out_580(u0_col_out_580),
    .col_out_581(u0_col_out_581),
    .col_out_582(u0_col_out_582),
    .col_out_583(u0_col_out_583),
    .col_out_584(u0_col_out_584),
    .col_out_585(u0_col_out_585),
    .col_out_586(u0_col_out_586),
    .col_out_587(u0_col_out_587),
    .col_out_588(u0_col_out_588),
    .col_out_589(u0_col_out_589),
    .col_out_590(u0_col_out_590),
    .col_out_591(u0_col_out_591),
    .col_out_592(u0_col_out_592),
    .col_out_593(u0_col_out_593),
    .col_out_594(u0_col_out_594),
    .col_out_595(u0_col_out_595),
    .col_out_596(u0_col_out_596),
    .col_out_597(u0_col_out_597),
    .col_out_598(u0_col_out_598),
    .col_out_599(u0_col_out_599),
    .col_out_600(u0_col_out_600),
    .col_out_601(u0_col_out_601),
    .col_out_602(u0_col_out_602),
    .col_out_603(u0_col_out_603),
    .col_out_604(u0_col_out_604),
    .col_out_605(u0_col_out_605),
    .col_out_606(u0_col_out_606),
    .col_out_607(u0_col_out_607),
    .col_out_608(u0_col_out_608),
    .col_out_609(u0_col_out_609),
    .col_out_610(u0_col_out_610),
    .col_out_611(u0_col_out_611),
    .col_out_612(u0_col_out_612),
    .col_out_613(u0_col_out_613),
    .col_out_614(u0_col_out_614),
    .col_out_615(u0_col_out_615),
    .col_out_616(u0_col_out_616),
    .col_out_617(u0_col_out_617),
    .col_out_618(u0_col_out_618),
    .col_out_619(u0_col_out_619),
    .col_out_620(u0_col_out_620),
    .col_out_621(u0_col_out_621),
    .col_out_622(u0_col_out_622),
    .col_out_623(u0_col_out_623),
    .col_out_624(u0_col_out_624),
    .col_out_625(u0_col_out_625),
    .col_out_626(u0_col_out_626),
    .col_out_627(u0_col_out_627),
    .col_out_628(u0_col_out_628),
    .col_out_629(u0_col_out_629),
    .col_out_630(u0_col_out_630),
    .col_out_631(u0_col_out_631),
    .col_out_632(u0_col_out_632),
    .col_out_633(u0_col_out_633),
    .col_out_634(u0_col_out_634),
    .col_out_635(u0_col_out_635),
    .col_out_636(u0_col_out_636),
    .col_out_637(u0_col_out_637),
    .col_out_638(u0_col_out_638),
    .col_out_639(u0_col_out_639),
    .col_out_640(u0_col_out_640),
    .col_out_641(u0_col_out_641),
    .col_out_642(u0_col_out_642),
    .col_out_643(u0_col_out_643),
    .col_out_644(u0_col_out_644),
    .col_out_645(u0_col_out_645),
    .col_out_646(u0_col_out_646),
    .col_out_647(u0_col_out_647),
    .col_out_648(u0_col_out_648),
    .col_out_649(u0_col_out_649),
    .col_out_650(u0_col_out_650),
    .col_out_651(u0_col_out_651),
    .col_out_652(u0_col_out_652),
    .col_out_653(u0_col_out_653),
    .col_out_654(u0_col_out_654),
    .col_out_655(u0_col_out_655),
    .col_out_656(u0_col_out_656),
    .col_out_657(u0_col_out_657),
    .col_out_658(u0_col_out_658),
    .col_out_659(u0_col_out_659),
    .col_out_660(u0_col_out_660),
    .col_out_661(u0_col_out_661),
    .col_out_662(u0_col_out_662),
    .col_out_663(u0_col_out_663),
    .col_out_664(u0_col_out_664),
    .col_out_665(u0_col_out_665),
    .col_out_666(u0_col_out_666),
    .col_out_667(u0_col_out_667),
    .col_out_668(u0_col_out_668),
    .col_out_669(u0_col_out_669),
    .col_out_670(u0_col_out_670),
    .col_out_671(u0_col_out_671),
    .col_out_672(u0_col_out_672),
    .col_out_673(u0_col_out_673),
    .col_out_674(u0_col_out_674),
    .col_out_675(u0_col_out_675),
    .col_out_676(u0_col_out_676),
    .col_out_677(u0_col_out_677),
    .col_out_678(u0_col_out_678),
    .col_out_679(u0_col_out_679),
    .col_out_680(u0_col_out_680),
    .col_out_681(u0_col_out_681),
    .col_out_682(u0_col_out_682),
    .col_out_683(u0_col_out_683),
    .col_out_684(u0_col_out_684),
    .col_out_685(u0_col_out_685),
    .col_out_686(u0_col_out_686),
    .col_out_687(u0_col_out_687),
    .col_out_688(u0_col_out_688),
    .col_out_689(u0_col_out_689),
    .col_out_690(u0_col_out_690),
    .col_out_691(u0_col_out_691),
    .col_out_692(u0_col_out_692),
    .col_out_693(u0_col_out_693),
    .col_out_694(u0_col_out_694),
    .col_out_695(u0_col_out_695),
    .col_out_696(u0_col_out_696),
    .col_out_697(u0_col_out_697),
    .col_out_698(u0_col_out_698),
    .col_out_699(u0_col_out_699),
    .col_out_700(u0_col_out_700),
    .col_out_701(u0_col_out_701),
    .col_out_702(u0_col_out_702),
    .col_out_703(u0_col_out_703),
    .col_out_704(u0_col_out_704),
    .col_out_705(u0_col_out_705),
    .col_out_706(u0_col_out_706),
    .col_out_707(u0_col_out_707),
    .col_out_708(u0_col_out_708),
    .col_out_709(u0_col_out_709),
    .col_out_710(u0_col_out_710),
    .col_out_711(u0_col_out_711),
    .col_out_712(u0_col_out_712),
    .col_out_713(u0_col_out_713),
    .col_out_714(u0_col_out_714),
    .col_out_715(u0_col_out_715),
    .col_out_716(u0_col_out_716),
    .col_out_717(u0_col_out_717),
    .col_out_718(u0_col_out_718),
    .col_out_719(u0_col_out_719),
    .col_out_720(u0_col_out_720),
    .col_out_721(u0_col_out_721),
    .col_out_722(u0_col_out_722),
    .col_out_723(u0_col_out_723),
    .col_out_724(u0_col_out_724),
    .col_out_725(u0_col_out_725),
    .col_out_726(u0_col_out_726),
    .col_out_727(u0_col_out_727),
    .col_out_728(u0_col_out_728),
    .col_out_729(u0_col_out_729),
    .col_out_730(u0_col_out_730),
    .col_out_731(u0_col_out_731),
    .col_out_732(u0_col_out_732),
    .col_out_733(u0_col_out_733),
    .col_out_734(u0_col_out_734),
    .col_out_735(u0_col_out_735),
    .col_out_736(u0_col_out_736),
    .col_out_737(u0_col_out_737),
    .col_out_738(u0_col_out_738),
    .col_out_739(u0_col_out_739),
    .col_out_740(u0_col_out_740),
    .col_out_741(u0_col_out_741),
    .col_out_742(u0_col_out_742),
    .col_out_743(u0_col_out_743),
    .col_out_744(u0_col_out_744),
    .col_out_745(u0_col_out_745),
    .col_out_746(u0_col_out_746),
    .col_out_747(u0_col_out_747),
    .col_out_748(u0_col_out_748),
    .col_out_749(u0_col_out_749),
    .col_out_750(u0_col_out_750),
    .col_out_751(u0_col_out_751),
    .col_out_752(u0_col_out_752),
    .col_out_753(u0_col_out_753),
    .col_out_754(u0_col_out_754),
    .col_out_755(u0_col_out_755),
    .col_out_756(u0_col_out_756),
    .col_out_757(u0_col_out_757),
    .col_out_758(u0_col_out_758),
    .col_out_759(u0_col_out_759),
    .col_out_760(u0_col_out_760),
    .col_out_761(u0_col_out_761),
    .col_out_762(u0_col_out_762),
    .col_out_763(u0_col_out_763),
    .col_out_764(u0_col_out_764),
    .col_out_765(u0_col_out_765),
    .col_out_766(u0_col_out_766),
    .col_out_767(u0_col_out_767),
    .col_out_768(u0_col_out_768),
    .col_out_769(u0_col_out_769),
    .col_out_770(u0_col_out_770),
    .col_out_771(u0_col_out_771),
    .col_out_772(u0_col_out_772),
    .col_out_773(u0_col_out_773),
    .col_out_774(u0_col_out_774),
    .col_out_775(u0_col_out_775),
    .col_out_776(u0_col_out_776),
    .col_out_777(u0_col_out_777),
    .col_out_778(u0_col_out_778),
    .col_out_779(u0_col_out_779),
    .col_out_780(u0_col_out_780),
    .col_out_781(u0_col_out_781),
    .col_out_782(u0_col_out_782),
    .col_out_783(u0_col_out_783),
    .col_out_784(u0_col_out_784),
    .col_out_785(u0_col_out_785),
    .col_out_786(u0_col_out_786),
    .col_out_787(u0_col_out_787),
    .col_out_788(u0_col_out_788),
    .col_out_789(u0_col_out_789),
    .col_out_790(u0_col_out_790),
    .col_out_791(u0_col_out_791),
    .col_out_792(u0_col_out_792),
    .col_out_793(u0_col_out_793),
    .col_out_794(u0_col_out_794),
    .col_out_795(u0_col_out_795),
    .col_out_796(u0_col_out_796),
    .col_out_797(u0_col_out_797),
    .col_out_798(u0_col_out_798),
    .col_out_799(u0_col_out_799),
    .col_out_800(u0_col_out_800),
    .col_out_801(u0_col_out_801),
    .col_out_802(u0_col_out_802),
    .col_out_803(u0_col_out_803),
    .col_out_804(u0_col_out_804),
    .col_out_805(u0_col_out_805),
    .col_out_806(u0_col_out_806),
    .col_out_807(u0_col_out_807),
    .col_out_808(u0_col_out_808),
    .col_out_809(u0_col_out_809),
    .col_out_810(u0_col_out_810),
    .col_out_811(u0_col_out_811),
    .col_out_812(u0_col_out_812),
    .col_out_813(u0_col_out_813),
    .col_out_814(u0_col_out_814),
    .col_out_815(u0_col_out_815),
    .col_out_816(u0_col_out_816),
    .col_out_817(u0_col_out_817),
    .col_out_818(u0_col_out_818),
    .col_out_819(u0_col_out_819),
    .col_out_820(u0_col_out_820),
    .col_out_821(u0_col_out_821),
    .col_out_822(u0_col_out_822),
    .col_out_823(u0_col_out_823),
    .col_out_824(u0_col_out_824),
    .col_out_825(u0_col_out_825),
    .col_out_826(u0_col_out_826),
    .col_out_827(u0_col_out_827),
    .col_out_828(u0_col_out_828),
    .col_out_829(u0_col_out_829),
    .col_out_830(u0_col_out_830),
    .col_out_831(u0_col_out_831),
    .col_out_832(u0_col_out_832),
    .col_out_833(u0_col_out_833),
    .col_out_834(u0_col_out_834),
    .col_out_835(u0_col_out_835),
    .col_out_836(u0_col_out_836),
    .col_out_837(u0_col_out_837),
    .col_out_838(u0_col_out_838),
    .col_out_839(u0_col_out_839),
    .col_out_840(u0_col_out_840),
    .col_out_841(u0_col_out_841),
    .col_out_842(u0_col_out_842),
    .col_out_843(u0_col_out_843),
    .col_out_844(u0_col_out_844),
    .col_out_845(u0_col_out_845),
    .col_out_846(u0_col_out_846),
    .col_out_847(u0_col_out_847),
    .col_out_848(u0_col_out_848),
    .col_out_849(u0_col_out_849),
    .col_out_850(u0_col_out_850),
    .col_out_851(u0_col_out_851),
    .col_out_852(u0_col_out_852),
    .col_out_853(u0_col_out_853),
    .col_out_854(u0_col_out_854),
    .col_out_855(u0_col_out_855),
    .col_out_856(u0_col_out_856),
    .col_out_857(u0_col_out_857),
    .col_out_858(u0_col_out_858),
    .col_out_859(u0_col_out_859),
    .col_out_860(u0_col_out_860),
    .col_out_861(u0_col_out_861),
    .col_out_862(u0_col_out_862),
    .col_out_863(u0_col_out_863),
    .col_out_864(u0_col_out_864),
    .col_out_865(u0_col_out_865),
    .col_out_866(u0_col_out_866),
    .col_out_867(u0_col_out_867),
    .col_out_868(u0_col_out_868),
    .col_out_869(u0_col_out_869),
    .col_out_870(u0_col_out_870),
    .col_out_871(u0_col_out_871),
    .col_out_872(u0_col_out_872),
    .col_out_873(u0_col_out_873),
    .col_out_874(u0_col_out_874),
    .col_out_875(u0_col_out_875),
    .col_out_876(u0_col_out_876),
    .col_out_877(u0_col_out_877),
    .col_out_878(u0_col_out_878),
    .col_out_879(u0_col_out_879),
    .col_out_880(u0_col_out_880),
    .col_out_881(u0_col_out_881),
    .col_out_882(u0_col_out_882),
    .col_out_883(u0_col_out_883),
    .col_out_884(u0_col_out_884),
    .col_out_885(u0_col_out_885),
    .col_out_886(u0_col_out_886),
    .col_out_887(u0_col_out_887),
    .col_out_888(u0_col_out_888),
    .col_out_889(u0_col_out_889),
    .col_out_890(u0_col_out_890),
    .col_out_891(u0_col_out_891),
    .col_out_892(u0_col_out_892),
    .col_out_893(u0_col_out_893),
    .col_out_894(u0_col_out_894),
    .col_out_895(u0_col_out_895),
    .col_out_896(u0_col_out_896),
    .col_out_897(u0_col_out_897),
    .col_out_898(u0_col_out_898),
    .col_out_899(u0_col_out_899),
    .col_out_900(u0_col_out_900),
    .col_out_901(u0_col_out_901),
    .col_out_902(u0_col_out_902),
    .col_out_903(u0_col_out_903),
    .col_out_904(u0_col_out_904),
    .col_out_905(u0_col_out_905),
    .col_out_906(u0_col_out_906),
    .col_out_907(u0_col_out_907),
    .col_out_908(u0_col_out_908),
    .col_out_909(u0_col_out_909),
    .col_out_910(u0_col_out_910),
    .col_out_911(u0_col_out_911),
    .col_out_912(u0_col_out_912),
    .col_out_913(u0_col_out_913),
    .col_out_914(u0_col_out_914),
    .col_out_915(u0_col_out_915),
    .col_out_916(u0_col_out_916),
    .col_out_917(u0_col_out_917),
    .col_out_918(u0_col_out_918),
    .col_out_919(u0_col_out_919),
    .col_out_920(u0_col_out_920),
    .col_out_921(u0_col_out_921),
    .col_out_922(u0_col_out_922),
    .col_out_923(u0_col_out_923),
    .col_out_924(u0_col_out_924),
    .col_out_925(u0_col_out_925),
    .col_out_926(u0_col_out_926),
    .col_out_927(u0_col_out_927),
    .col_out_928(u0_col_out_928),
    .col_out_929(u0_col_out_929),
    .col_out_930(u0_col_out_930),
    .col_out_931(u0_col_out_931),
    .col_out_932(u0_col_out_932),
    .col_out_933(u0_col_out_933),
    .col_out_934(u0_col_out_934),
    .col_out_935(u0_col_out_935),
    .col_out_936(u0_col_out_936),
    .col_out_937(u0_col_out_937),
    .col_out_938(u0_col_out_938),
    .col_out_939(u0_col_out_939),
    .col_out_940(u0_col_out_940),
    .col_out_941(u0_col_out_941),
    .col_out_942(u0_col_out_942),
    .col_out_943(u0_col_out_943),
    .col_out_944(u0_col_out_944),
    .col_out_945(u0_col_out_945),
    .col_out_946(u0_col_out_946),
    .col_out_947(u0_col_out_947),
    .col_out_948(u0_col_out_948),
    .col_out_949(u0_col_out_949),
    .col_out_950(u0_col_out_950),
    .col_out_951(u0_col_out_951),
    .col_out_952(u0_col_out_952),
    .col_out_953(u0_col_out_953),
    .col_out_954(u0_col_out_954),
    .col_out_955(u0_col_out_955),
    .col_out_956(u0_col_out_956),
    .col_out_957(u0_col_out_957),
    .col_out_958(u0_col_out_958),
    .col_out_959(u0_col_out_959),
    .col_out_960(u0_col_out_960),
    .col_out_961(u0_col_out_961),
    .col_out_962(u0_col_out_962),
    .col_out_963(u0_col_out_963),
    .col_out_964(u0_col_out_964),
    .col_out_965(u0_col_out_965),
    .col_out_966(u0_col_out_966),
    .col_out_967(u0_col_out_967),
    .col_out_968(u0_col_out_968),
    .col_out_969(u0_col_out_969),
    .col_out_970(u0_col_out_970),
    .col_out_971(u0_col_out_971),
    .col_out_972(u0_col_out_972),
    .col_out_973(u0_col_out_973),
    .col_out_974(u0_col_out_974),
    .col_out_975(u0_col_out_975),
    .col_out_976(u0_col_out_976),
    .col_out_977(u0_col_out_977),
    .col_out_978(u0_col_out_978),
    .col_out_979(u0_col_out_979),
    .col_out_980(u0_col_out_980),
    .col_out_981(u0_col_out_981),
    .col_out_982(u0_col_out_982),
    .col_out_983(u0_col_out_983),
    .col_out_984(u0_col_out_984),
    .col_out_985(u0_col_out_985),
    .col_out_986(u0_col_out_986),
    .col_out_987(u0_col_out_987),
    .col_out_988(u0_col_out_988),
    .col_out_989(u0_col_out_989),
    .col_out_990(u0_col_out_990),
    .col_out_991(u0_col_out_991),
    .col_out_992(u0_col_out_992),
    .col_out_993(u0_col_out_993),
    .col_out_994(u0_col_out_994),
    .col_out_995(u0_col_out_995),
    .col_out_996(u0_col_out_996),
    .col_out_997(u0_col_out_997),
    .col_out_998(u0_col_out_998),
    .col_out_999(u0_col_out_999),
    .col_out_1000(u0_col_out_1000),
    .col_out_1001(u0_col_out_1001),
    .col_out_1002(u0_col_out_1002),
    .col_out_1003(u0_col_out_1003),
    .col_out_1004(u0_col_out_1004),
    .col_out_1005(u0_col_out_1005),
    .col_out_1006(u0_col_out_1006),
    .col_out_1007(u0_col_out_1007),
    .col_out_1008(u0_col_out_1008),
    .col_out_1009(u0_col_out_1009),
    .col_out_1010(u0_col_out_1010),
    .col_out_1011(u0_col_out_1011),
    .col_out_1012(u0_col_out_1012),
    .col_out_1013(u0_col_out_1013),
    .col_out_1014(u0_col_out_1014),
    .col_out_1015(u0_col_out_1015),
    .col_out_1016(u0_col_out_1016),
    .col_out_1017(u0_col_out_1017),
    .col_out_1018(u0_col_out_1018),
    .col_out_1019(u0_col_out_1019),
    .col_out_1020(u0_col_out_1020),
    .col_out_1021(u0_col_out_1021),
    .col_out_1022(u0_col_out_1022),
    .col_out_1023(u0_col_out_1023)
);


wire [235:0] u1_col_in_0;
wire [235:0] u1_col_in_1;
wire [235:0] u1_col_in_2;
wire [235:0] u1_col_in_3;
wire [235:0] u1_col_in_4;
wire [235:0] u1_col_in_5;
wire [235:0] u1_col_in_6;
wire [235:0] u1_col_in_7;
wire [235:0] u1_col_in_8;
wire [235:0] u1_col_in_9;
wire [235:0] u1_col_in_10;
wire [235:0] u1_col_in_11;
wire [235:0] u1_col_in_12;
wire [235:0] u1_col_in_13;
wire [235:0] u1_col_in_14;
wire [235:0] u1_col_in_15;
wire [235:0] u1_col_in_16;
wire [235:0] u1_col_in_17;
wire [235:0] u1_col_in_18;
wire [235:0] u1_col_in_19;
wire [235:0] u1_col_in_20;
wire [235:0] u1_col_in_21;
wire [235:0] u1_col_in_22;
wire [235:0] u1_col_in_23;
wire [235:0] u1_col_in_24;
wire [235:0] u1_col_in_25;
wire [235:0] u1_col_in_26;
wire [235:0] u1_col_in_27;
wire [235:0] u1_col_in_28;
wire [235:0] u1_col_in_29;
wire [235:0] u1_col_in_30;
wire [235:0] u1_col_in_31;
wire [235:0] u1_col_in_32;
wire [235:0] u1_col_in_33;
wire [235:0] u1_col_in_34;
wire [235:0] u1_col_in_35;
wire [235:0] u1_col_in_36;
wire [235:0] u1_col_in_37;
wire [235:0] u1_col_in_38;
wire [235:0] u1_col_in_39;
wire [235:0] u1_col_in_40;
wire [235:0] u1_col_in_41;
wire [235:0] u1_col_in_42;
wire [235:0] u1_col_in_43;
wire [235:0] u1_col_in_44;
wire [235:0] u1_col_in_45;
wire [235:0] u1_col_in_46;
wire [235:0] u1_col_in_47;
wire [235:0] u1_col_in_48;
wire [235:0] u1_col_in_49;
wire [235:0] u1_col_in_50;
wire [235:0] u1_col_in_51;
wire [235:0] u1_col_in_52;
wire [235:0] u1_col_in_53;
wire [235:0] u1_col_in_54;
wire [235:0] u1_col_in_55;
wire [235:0] u1_col_in_56;
wire [235:0] u1_col_in_57;
wire [235:0] u1_col_in_58;
wire [235:0] u1_col_in_59;
wire [235:0] u1_col_in_60;
wire [235:0] u1_col_in_61;
wire [235:0] u1_col_in_62;
wire [235:0] u1_col_in_63;
wire [235:0] u1_col_in_64;
wire [235:0] u1_col_in_65;
wire [235:0] u1_col_in_66;
wire [235:0] u1_col_in_67;
wire [235:0] u1_col_in_68;
wire [235:0] u1_col_in_69;
wire [235:0] u1_col_in_70;
wire [235:0] u1_col_in_71;
wire [235:0] u1_col_in_72;
wire [235:0] u1_col_in_73;
wire [235:0] u1_col_in_74;
wire [235:0] u1_col_in_75;
wire [235:0] u1_col_in_76;
wire [235:0] u1_col_in_77;
wire [235:0] u1_col_in_78;
wire [235:0] u1_col_in_79;
wire [235:0] u1_col_in_80;
wire [235:0] u1_col_in_81;
wire [235:0] u1_col_in_82;
wire [235:0] u1_col_in_83;
wire [235:0] u1_col_in_84;
wire [235:0] u1_col_in_85;
wire [235:0] u1_col_in_86;
wire [235:0] u1_col_in_87;
wire [235:0] u1_col_in_88;
wire [235:0] u1_col_in_89;
wire [235:0] u1_col_in_90;
wire [235:0] u1_col_in_91;
wire [235:0] u1_col_in_92;
wire [235:0] u1_col_in_93;
wire [235:0] u1_col_in_94;
wire [235:0] u1_col_in_95;
wire [235:0] u1_col_in_96;
wire [235:0] u1_col_in_97;
wire [235:0] u1_col_in_98;
wire [235:0] u1_col_in_99;
wire [235:0] u1_col_in_100;
wire [235:0] u1_col_in_101;
wire [235:0] u1_col_in_102;
wire [235:0] u1_col_in_103;
wire [235:0] u1_col_in_104;
wire [235:0] u1_col_in_105;
wire [235:0] u1_col_in_106;
wire [235:0] u1_col_in_107;
wire [235:0] u1_col_in_108;
wire [235:0] u1_col_in_109;
wire [235:0] u1_col_in_110;
wire [235:0] u1_col_in_111;
wire [235:0] u1_col_in_112;
wire [235:0] u1_col_in_113;
wire [235:0] u1_col_in_114;
wire [235:0] u1_col_in_115;
wire [235:0] u1_col_in_116;
wire [235:0] u1_col_in_117;
wire [235:0] u1_col_in_118;
wire [235:0] u1_col_in_119;
wire [235:0] u1_col_in_120;
wire [235:0] u1_col_in_121;
wire [235:0] u1_col_in_122;
wire [235:0] u1_col_in_123;
wire [235:0] u1_col_in_124;
wire [235:0] u1_col_in_125;
wire [235:0] u1_col_in_126;
wire [235:0] u1_col_in_127;
wire [235:0] u1_col_in_128;
wire [235:0] u1_col_in_129;
wire [235:0] u1_col_in_130;
wire [235:0] u1_col_in_131;
wire [235:0] u1_col_in_132;
wire [235:0] u1_col_in_133;
wire [235:0] u1_col_in_134;
wire [235:0] u1_col_in_135;
wire [235:0] u1_col_in_136;
wire [235:0] u1_col_in_137;
wire [235:0] u1_col_in_138;
wire [235:0] u1_col_in_139;
wire [235:0] u1_col_in_140;
wire [235:0] u1_col_in_141;
wire [235:0] u1_col_in_142;
wire [235:0] u1_col_in_143;
wire [235:0] u1_col_in_144;
wire [235:0] u1_col_in_145;
wire [235:0] u1_col_in_146;
wire [235:0] u1_col_in_147;
wire [235:0] u1_col_in_148;
wire [235:0] u1_col_in_149;
wire [235:0] u1_col_in_150;
wire [235:0] u1_col_in_151;
wire [235:0] u1_col_in_152;
wire [235:0] u1_col_in_153;
wire [235:0] u1_col_in_154;
wire [235:0] u1_col_in_155;
wire [235:0] u1_col_in_156;
wire [235:0] u1_col_in_157;
wire [235:0] u1_col_in_158;
wire [235:0] u1_col_in_159;
wire [235:0] u1_col_in_160;
wire [235:0] u1_col_in_161;
wire [235:0] u1_col_in_162;
wire [235:0] u1_col_in_163;
wire [235:0] u1_col_in_164;
wire [235:0] u1_col_in_165;
wire [235:0] u1_col_in_166;
wire [235:0] u1_col_in_167;
wire [235:0] u1_col_in_168;
wire [235:0] u1_col_in_169;
wire [235:0] u1_col_in_170;
wire [235:0] u1_col_in_171;
wire [235:0] u1_col_in_172;
wire [235:0] u1_col_in_173;
wire [235:0] u1_col_in_174;
wire [235:0] u1_col_in_175;
wire [235:0] u1_col_in_176;
wire [235:0] u1_col_in_177;
wire [235:0] u1_col_in_178;
wire [235:0] u1_col_in_179;
wire [235:0] u1_col_in_180;
wire [235:0] u1_col_in_181;
wire [235:0] u1_col_in_182;
wire [235:0] u1_col_in_183;
wire [235:0] u1_col_in_184;
wire [235:0] u1_col_in_185;
wire [235:0] u1_col_in_186;
wire [235:0] u1_col_in_187;
wire [235:0] u1_col_in_188;
wire [235:0] u1_col_in_189;
wire [235:0] u1_col_in_190;
wire [235:0] u1_col_in_191;
wire [235:0] u1_col_in_192;
wire [235:0] u1_col_in_193;
wire [235:0] u1_col_in_194;
wire [235:0] u1_col_in_195;
wire [235:0] u1_col_in_196;
wire [235:0] u1_col_in_197;
wire [235:0] u1_col_in_198;
wire [235:0] u1_col_in_199;
wire [235:0] u1_col_in_200;
wire [235:0] u1_col_in_201;
wire [235:0] u1_col_in_202;
wire [235:0] u1_col_in_203;
wire [235:0] u1_col_in_204;
wire [235:0] u1_col_in_205;
wire [235:0] u1_col_in_206;
wire [235:0] u1_col_in_207;
wire [235:0] u1_col_in_208;
wire [235:0] u1_col_in_209;
wire [235:0] u1_col_in_210;
wire [235:0] u1_col_in_211;
wire [235:0] u1_col_in_212;
wire [235:0] u1_col_in_213;
wire [235:0] u1_col_in_214;
wire [235:0] u1_col_in_215;
wire [235:0] u1_col_in_216;
wire [235:0] u1_col_in_217;
wire [235:0] u1_col_in_218;
wire [235:0] u1_col_in_219;
wire [235:0] u1_col_in_220;
wire [235:0] u1_col_in_221;
wire [235:0] u1_col_in_222;
wire [235:0] u1_col_in_223;
wire [235:0] u1_col_in_224;
wire [235:0] u1_col_in_225;
wire [235:0] u1_col_in_226;
wire [235:0] u1_col_in_227;
wire [235:0] u1_col_in_228;
wire [235:0] u1_col_in_229;
wire [235:0] u1_col_in_230;
wire [235:0] u1_col_in_231;
wire [235:0] u1_col_in_232;
wire [235:0] u1_col_in_233;
wire [235:0] u1_col_in_234;
wire [235:0] u1_col_in_235;
wire [235:0] u1_col_in_236;
wire [235:0] u1_col_in_237;
wire [235:0] u1_col_in_238;
wire [235:0] u1_col_in_239;
wire [235:0] u1_col_in_240;
wire [235:0] u1_col_in_241;
wire [235:0] u1_col_in_242;
wire [235:0] u1_col_in_243;
wire [235:0] u1_col_in_244;
wire [235:0] u1_col_in_245;
wire [235:0] u1_col_in_246;
wire [235:0] u1_col_in_247;
wire [235:0] u1_col_in_248;
wire [235:0] u1_col_in_249;
wire [235:0] u1_col_in_250;
wire [235:0] u1_col_in_251;
wire [235:0] u1_col_in_252;
wire [235:0] u1_col_in_253;
wire [235:0] u1_col_in_254;
wire [235:0] u1_col_in_255;
wire [235:0] u1_col_in_256;
wire [235:0] u1_col_in_257;
wire [235:0] u1_col_in_258;
wire [235:0] u1_col_in_259;
wire [235:0] u1_col_in_260;
wire [235:0] u1_col_in_261;
wire [235:0] u1_col_in_262;
wire [235:0] u1_col_in_263;
wire [235:0] u1_col_in_264;
wire [235:0] u1_col_in_265;
wire [235:0] u1_col_in_266;
wire [235:0] u1_col_in_267;
wire [235:0] u1_col_in_268;
wire [235:0] u1_col_in_269;
wire [235:0] u1_col_in_270;
wire [235:0] u1_col_in_271;
wire [235:0] u1_col_in_272;
wire [235:0] u1_col_in_273;
wire [235:0] u1_col_in_274;
wire [235:0] u1_col_in_275;
wire [235:0] u1_col_in_276;
wire [235:0] u1_col_in_277;
wire [235:0] u1_col_in_278;
wire [235:0] u1_col_in_279;
wire [235:0] u1_col_in_280;
wire [235:0] u1_col_in_281;
wire [235:0] u1_col_in_282;
wire [235:0] u1_col_in_283;
wire [235:0] u1_col_in_284;
wire [235:0] u1_col_in_285;
wire [235:0] u1_col_in_286;
wire [235:0] u1_col_in_287;
wire [235:0] u1_col_in_288;
wire [235:0] u1_col_in_289;
wire [235:0] u1_col_in_290;
wire [235:0] u1_col_in_291;
wire [235:0] u1_col_in_292;
wire [235:0] u1_col_in_293;
wire [235:0] u1_col_in_294;
wire [235:0] u1_col_in_295;
wire [235:0] u1_col_in_296;
wire [235:0] u1_col_in_297;
wire [235:0] u1_col_in_298;
wire [235:0] u1_col_in_299;
wire [235:0] u1_col_in_300;
wire [235:0] u1_col_in_301;
wire [235:0] u1_col_in_302;
wire [235:0] u1_col_in_303;
wire [235:0] u1_col_in_304;
wire [235:0] u1_col_in_305;
wire [235:0] u1_col_in_306;
wire [235:0] u1_col_in_307;
wire [235:0] u1_col_in_308;
wire [235:0] u1_col_in_309;
wire [235:0] u1_col_in_310;
wire [235:0] u1_col_in_311;
wire [235:0] u1_col_in_312;
wire [235:0] u1_col_in_313;
wire [235:0] u1_col_in_314;
wire [235:0] u1_col_in_315;
wire [235:0] u1_col_in_316;
wire [235:0] u1_col_in_317;
wire [235:0] u1_col_in_318;
wire [235:0] u1_col_in_319;
wire [235:0] u1_col_in_320;
wire [235:0] u1_col_in_321;
wire [235:0] u1_col_in_322;
wire [235:0] u1_col_in_323;
wire [235:0] u1_col_in_324;
wire [235:0] u1_col_in_325;
wire [235:0] u1_col_in_326;
wire [235:0] u1_col_in_327;
wire [235:0] u1_col_in_328;
wire [235:0] u1_col_in_329;
wire [235:0] u1_col_in_330;
wire [235:0] u1_col_in_331;
wire [235:0] u1_col_in_332;
wire [235:0] u1_col_in_333;
wire [235:0] u1_col_in_334;
wire [235:0] u1_col_in_335;
wire [235:0] u1_col_in_336;
wire [235:0] u1_col_in_337;
wire [235:0] u1_col_in_338;
wire [235:0] u1_col_in_339;
wire [235:0] u1_col_in_340;
wire [235:0] u1_col_in_341;
wire [235:0] u1_col_in_342;
wire [235:0] u1_col_in_343;
wire [235:0] u1_col_in_344;
wire [235:0] u1_col_in_345;
wire [235:0] u1_col_in_346;
wire [235:0] u1_col_in_347;
wire [235:0] u1_col_in_348;
wire [235:0] u1_col_in_349;
wire [235:0] u1_col_in_350;
wire [235:0] u1_col_in_351;
wire [235:0] u1_col_in_352;
wire [235:0] u1_col_in_353;
wire [235:0] u1_col_in_354;
wire [235:0] u1_col_in_355;
wire [235:0] u1_col_in_356;
wire [235:0] u1_col_in_357;
wire [235:0] u1_col_in_358;
wire [235:0] u1_col_in_359;
wire [235:0] u1_col_in_360;
wire [235:0] u1_col_in_361;
wire [235:0] u1_col_in_362;
wire [235:0] u1_col_in_363;
wire [235:0] u1_col_in_364;
wire [235:0] u1_col_in_365;
wire [235:0] u1_col_in_366;
wire [235:0] u1_col_in_367;
wire [235:0] u1_col_in_368;
wire [235:0] u1_col_in_369;
wire [235:0] u1_col_in_370;
wire [235:0] u1_col_in_371;
wire [235:0] u1_col_in_372;
wire [235:0] u1_col_in_373;
wire [235:0] u1_col_in_374;
wire [235:0] u1_col_in_375;
wire [235:0] u1_col_in_376;
wire [235:0] u1_col_in_377;
wire [235:0] u1_col_in_378;
wire [235:0] u1_col_in_379;
wire [235:0] u1_col_in_380;
wire [235:0] u1_col_in_381;
wire [235:0] u1_col_in_382;
wire [235:0] u1_col_in_383;
wire [235:0] u1_col_in_384;
wire [235:0] u1_col_in_385;
wire [235:0] u1_col_in_386;
wire [235:0] u1_col_in_387;
wire [235:0] u1_col_in_388;
wire [235:0] u1_col_in_389;
wire [235:0] u1_col_in_390;
wire [235:0] u1_col_in_391;
wire [235:0] u1_col_in_392;
wire [235:0] u1_col_in_393;
wire [235:0] u1_col_in_394;
wire [235:0] u1_col_in_395;
wire [235:0] u1_col_in_396;
wire [235:0] u1_col_in_397;
wire [235:0] u1_col_in_398;
wire [235:0] u1_col_in_399;
wire [235:0] u1_col_in_400;
wire [235:0] u1_col_in_401;
wire [235:0] u1_col_in_402;
wire [235:0] u1_col_in_403;
wire [235:0] u1_col_in_404;
wire [235:0] u1_col_in_405;
wire [235:0] u1_col_in_406;
wire [235:0] u1_col_in_407;
wire [235:0] u1_col_in_408;
wire [235:0] u1_col_in_409;
wire [235:0] u1_col_in_410;
wire [235:0] u1_col_in_411;
wire [235:0] u1_col_in_412;
wire [235:0] u1_col_in_413;
wire [235:0] u1_col_in_414;
wire [235:0] u1_col_in_415;
wire [235:0] u1_col_in_416;
wire [235:0] u1_col_in_417;
wire [235:0] u1_col_in_418;
wire [235:0] u1_col_in_419;
wire [235:0] u1_col_in_420;
wire [235:0] u1_col_in_421;
wire [235:0] u1_col_in_422;
wire [235:0] u1_col_in_423;
wire [235:0] u1_col_in_424;
wire [235:0] u1_col_in_425;
wire [235:0] u1_col_in_426;
wire [235:0] u1_col_in_427;
wire [235:0] u1_col_in_428;
wire [235:0] u1_col_in_429;
wire [235:0] u1_col_in_430;
wire [235:0] u1_col_in_431;
wire [235:0] u1_col_in_432;
wire [235:0] u1_col_in_433;
wire [235:0] u1_col_in_434;
wire [235:0] u1_col_in_435;
wire [235:0] u1_col_in_436;
wire [235:0] u1_col_in_437;
wire [235:0] u1_col_in_438;
wire [235:0] u1_col_in_439;
wire [235:0] u1_col_in_440;
wire [235:0] u1_col_in_441;
wire [235:0] u1_col_in_442;
wire [235:0] u1_col_in_443;
wire [235:0] u1_col_in_444;
wire [235:0] u1_col_in_445;
wire [235:0] u1_col_in_446;
wire [235:0] u1_col_in_447;
wire [235:0] u1_col_in_448;
wire [235:0] u1_col_in_449;
wire [235:0] u1_col_in_450;
wire [235:0] u1_col_in_451;
wire [235:0] u1_col_in_452;
wire [235:0] u1_col_in_453;
wire [235:0] u1_col_in_454;
wire [235:0] u1_col_in_455;
wire [235:0] u1_col_in_456;
wire [235:0] u1_col_in_457;
wire [235:0] u1_col_in_458;
wire [235:0] u1_col_in_459;
wire [235:0] u1_col_in_460;
wire [235:0] u1_col_in_461;
wire [235:0] u1_col_in_462;
wire [235:0] u1_col_in_463;
wire [235:0] u1_col_in_464;
wire [235:0] u1_col_in_465;
wire [235:0] u1_col_in_466;
wire [235:0] u1_col_in_467;
wire [235:0] u1_col_in_468;
wire [235:0] u1_col_in_469;
wire [235:0] u1_col_in_470;
wire [235:0] u1_col_in_471;
wire [235:0] u1_col_in_472;
wire [235:0] u1_col_in_473;
wire [235:0] u1_col_in_474;
wire [235:0] u1_col_in_475;
wire [235:0] u1_col_in_476;
wire [235:0] u1_col_in_477;
wire [235:0] u1_col_in_478;
wire [235:0] u1_col_in_479;
wire [235:0] u1_col_in_480;
wire [235:0] u1_col_in_481;
wire [235:0] u1_col_in_482;
wire [235:0] u1_col_in_483;
wire [235:0] u1_col_in_484;
wire [235:0] u1_col_in_485;
wire [235:0] u1_col_in_486;
wire [235:0] u1_col_in_487;
wire [235:0] u1_col_in_488;
wire [235:0] u1_col_in_489;
wire [235:0] u1_col_in_490;
wire [235:0] u1_col_in_491;
wire [235:0] u1_col_in_492;
wire [235:0] u1_col_in_493;
wire [235:0] u1_col_in_494;
wire [235:0] u1_col_in_495;
wire [235:0] u1_col_in_496;
wire [235:0] u1_col_in_497;
wire [235:0] u1_col_in_498;
wire [235:0] u1_col_in_499;
wire [235:0] u1_col_in_500;
wire [235:0] u1_col_in_501;
wire [235:0] u1_col_in_502;
wire [235:0] u1_col_in_503;
wire [235:0] u1_col_in_504;
wire [235:0] u1_col_in_505;
wire [235:0] u1_col_in_506;
wire [235:0] u1_col_in_507;
wire [235:0] u1_col_in_508;
wire [235:0] u1_col_in_509;
wire [235:0] u1_col_in_510;
wire [235:0] u1_col_in_511;
wire [235:0] u1_col_in_512;
wire [235:0] u1_col_in_513;
wire [235:0] u1_col_in_514;
wire [235:0] u1_col_in_515;
wire [235:0] u1_col_in_516;
wire [235:0] u1_col_in_517;
wire [235:0] u1_col_in_518;
wire [235:0] u1_col_in_519;
wire [235:0] u1_col_in_520;
wire [235:0] u1_col_in_521;
wire [235:0] u1_col_in_522;
wire [235:0] u1_col_in_523;
wire [235:0] u1_col_in_524;
wire [235:0] u1_col_in_525;
wire [235:0] u1_col_in_526;
wire [235:0] u1_col_in_527;
wire [235:0] u1_col_in_528;
wire [235:0] u1_col_in_529;
wire [235:0] u1_col_in_530;
wire [235:0] u1_col_in_531;
wire [235:0] u1_col_in_532;
wire [235:0] u1_col_in_533;
wire [235:0] u1_col_in_534;
wire [235:0] u1_col_in_535;
wire [235:0] u1_col_in_536;
wire [235:0] u1_col_in_537;
wire [235:0] u1_col_in_538;
wire [235:0] u1_col_in_539;
wire [235:0] u1_col_in_540;
wire [235:0] u1_col_in_541;
wire [235:0] u1_col_in_542;
wire [235:0] u1_col_in_543;
wire [235:0] u1_col_in_544;
wire [235:0] u1_col_in_545;
wire [235:0] u1_col_in_546;
wire [235:0] u1_col_in_547;
wire [235:0] u1_col_in_548;
wire [235:0] u1_col_in_549;
wire [235:0] u1_col_in_550;
wire [235:0] u1_col_in_551;
wire [235:0] u1_col_in_552;
wire [235:0] u1_col_in_553;
wire [235:0] u1_col_in_554;
wire [235:0] u1_col_in_555;
wire [235:0] u1_col_in_556;
wire [235:0] u1_col_in_557;
wire [235:0] u1_col_in_558;
wire [235:0] u1_col_in_559;
wire [235:0] u1_col_in_560;
wire [235:0] u1_col_in_561;
wire [235:0] u1_col_in_562;
wire [235:0] u1_col_in_563;
wire [235:0] u1_col_in_564;
wire [235:0] u1_col_in_565;
wire [235:0] u1_col_in_566;
wire [235:0] u1_col_in_567;
wire [235:0] u1_col_in_568;
wire [235:0] u1_col_in_569;
wire [235:0] u1_col_in_570;
wire [235:0] u1_col_in_571;
wire [235:0] u1_col_in_572;
wire [235:0] u1_col_in_573;
wire [235:0] u1_col_in_574;
wire [235:0] u1_col_in_575;
wire [235:0] u1_col_in_576;
wire [235:0] u1_col_in_577;
wire [235:0] u1_col_in_578;
wire [235:0] u1_col_in_579;
wire [235:0] u1_col_in_580;
wire [235:0] u1_col_in_581;
wire [235:0] u1_col_in_582;
wire [235:0] u1_col_in_583;
wire [235:0] u1_col_in_584;
wire [235:0] u1_col_in_585;
wire [235:0] u1_col_in_586;
wire [235:0] u1_col_in_587;
wire [235:0] u1_col_in_588;
wire [235:0] u1_col_in_589;
wire [235:0] u1_col_in_590;
wire [235:0] u1_col_in_591;
wire [235:0] u1_col_in_592;
wire [235:0] u1_col_in_593;
wire [235:0] u1_col_in_594;
wire [235:0] u1_col_in_595;
wire [235:0] u1_col_in_596;
wire [235:0] u1_col_in_597;
wire [235:0] u1_col_in_598;
wire [235:0] u1_col_in_599;
wire [235:0] u1_col_in_600;
wire [235:0] u1_col_in_601;
wire [235:0] u1_col_in_602;
wire [235:0] u1_col_in_603;
wire [235:0] u1_col_in_604;
wire [235:0] u1_col_in_605;
wire [235:0] u1_col_in_606;
wire [235:0] u1_col_in_607;
wire [235:0] u1_col_in_608;
wire [235:0] u1_col_in_609;
wire [235:0] u1_col_in_610;
wire [235:0] u1_col_in_611;
wire [235:0] u1_col_in_612;
wire [235:0] u1_col_in_613;
wire [235:0] u1_col_in_614;
wire [235:0] u1_col_in_615;
wire [235:0] u1_col_in_616;
wire [235:0] u1_col_in_617;
wire [235:0] u1_col_in_618;
wire [235:0] u1_col_in_619;
wire [235:0] u1_col_in_620;
wire [235:0] u1_col_in_621;
wire [235:0] u1_col_in_622;
wire [235:0] u1_col_in_623;
wire [235:0] u1_col_in_624;
wire [235:0] u1_col_in_625;
wire [235:0] u1_col_in_626;
wire [235:0] u1_col_in_627;
wire [235:0] u1_col_in_628;
wire [235:0] u1_col_in_629;
wire [235:0] u1_col_in_630;
wire [235:0] u1_col_in_631;
wire [235:0] u1_col_in_632;
wire [235:0] u1_col_in_633;
wire [235:0] u1_col_in_634;
wire [235:0] u1_col_in_635;
wire [235:0] u1_col_in_636;
wire [235:0] u1_col_in_637;
wire [235:0] u1_col_in_638;
wire [235:0] u1_col_in_639;
wire [235:0] u1_col_in_640;
wire [235:0] u1_col_in_641;
wire [235:0] u1_col_in_642;
wire [235:0] u1_col_in_643;
wire [235:0] u1_col_in_644;
wire [235:0] u1_col_in_645;
wire [235:0] u1_col_in_646;
wire [235:0] u1_col_in_647;
wire [235:0] u1_col_in_648;
wire [235:0] u1_col_in_649;
wire [235:0] u1_col_in_650;
wire [235:0] u1_col_in_651;
wire [235:0] u1_col_in_652;
wire [235:0] u1_col_in_653;
wire [235:0] u1_col_in_654;
wire [235:0] u1_col_in_655;
wire [235:0] u1_col_in_656;
wire [235:0] u1_col_in_657;
wire [235:0] u1_col_in_658;
wire [235:0] u1_col_in_659;
wire [235:0] u1_col_in_660;
wire [235:0] u1_col_in_661;
wire [235:0] u1_col_in_662;
wire [235:0] u1_col_in_663;
wire [235:0] u1_col_in_664;
wire [235:0] u1_col_in_665;
wire [235:0] u1_col_in_666;
wire [235:0] u1_col_in_667;
wire [235:0] u1_col_in_668;
wire [235:0] u1_col_in_669;
wire [235:0] u1_col_in_670;
wire [235:0] u1_col_in_671;
wire [235:0] u1_col_in_672;
wire [235:0] u1_col_in_673;
wire [235:0] u1_col_in_674;
wire [235:0] u1_col_in_675;
wire [235:0] u1_col_in_676;
wire [235:0] u1_col_in_677;
wire [235:0] u1_col_in_678;
wire [235:0] u1_col_in_679;
wire [235:0] u1_col_in_680;
wire [235:0] u1_col_in_681;
wire [235:0] u1_col_in_682;
wire [235:0] u1_col_in_683;
wire [235:0] u1_col_in_684;
wire [235:0] u1_col_in_685;
wire [235:0] u1_col_in_686;
wire [235:0] u1_col_in_687;
wire [235:0] u1_col_in_688;
wire [235:0] u1_col_in_689;
wire [235:0] u1_col_in_690;
wire [235:0] u1_col_in_691;
wire [235:0] u1_col_in_692;
wire [235:0] u1_col_in_693;
wire [235:0] u1_col_in_694;
wire [235:0] u1_col_in_695;
wire [235:0] u1_col_in_696;
wire [235:0] u1_col_in_697;
wire [235:0] u1_col_in_698;
wire [235:0] u1_col_in_699;
wire [235:0] u1_col_in_700;
wire [235:0] u1_col_in_701;
wire [235:0] u1_col_in_702;
wire [235:0] u1_col_in_703;
wire [235:0] u1_col_in_704;
wire [235:0] u1_col_in_705;
wire [235:0] u1_col_in_706;
wire [235:0] u1_col_in_707;
wire [235:0] u1_col_in_708;
wire [235:0] u1_col_in_709;
wire [235:0] u1_col_in_710;
wire [235:0] u1_col_in_711;
wire [235:0] u1_col_in_712;
wire [235:0] u1_col_in_713;
wire [235:0] u1_col_in_714;
wire [235:0] u1_col_in_715;
wire [235:0] u1_col_in_716;
wire [235:0] u1_col_in_717;
wire [235:0] u1_col_in_718;
wire [235:0] u1_col_in_719;
wire [235:0] u1_col_in_720;
wire [235:0] u1_col_in_721;
wire [235:0] u1_col_in_722;
wire [235:0] u1_col_in_723;
wire [235:0] u1_col_in_724;
wire [235:0] u1_col_in_725;
wire [235:0] u1_col_in_726;
wire [235:0] u1_col_in_727;
wire [235:0] u1_col_in_728;
wire [235:0] u1_col_in_729;
wire [235:0] u1_col_in_730;
wire [235:0] u1_col_in_731;
wire [235:0] u1_col_in_732;
wire [235:0] u1_col_in_733;
wire [235:0] u1_col_in_734;
wire [235:0] u1_col_in_735;
wire [235:0] u1_col_in_736;
wire [235:0] u1_col_in_737;
wire [235:0] u1_col_in_738;
wire [235:0] u1_col_in_739;
wire [235:0] u1_col_in_740;
wire [235:0] u1_col_in_741;
wire [235:0] u1_col_in_742;
wire [235:0] u1_col_in_743;
wire [235:0] u1_col_in_744;
wire [235:0] u1_col_in_745;
wire [235:0] u1_col_in_746;
wire [235:0] u1_col_in_747;
wire [235:0] u1_col_in_748;
wire [235:0] u1_col_in_749;
wire [235:0] u1_col_in_750;
wire [235:0] u1_col_in_751;
wire [235:0] u1_col_in_752;
wire [235:0] u1_col_in_753;
wire [235:0] u1_col_in_754;
wire [235:0] u1_col_in_755;
wire [235:0] u1_col_in_756;
wire [235:0] u1_col_in_757;
wire [235:0] u1_col_in_758;
wire [235:0] u1_col_in_759;
wire [235:0] u1_col_in_760;
wire [235:0] u1_col_in_761;
wire [235:0] u1_col_in_762;
wire [235:0] u1_col_in_763;
wire [235:0] u1_col_in_764;
wire [235:0] u1_col_in_765;
wire [235:0] u1_col_in_766;
wire [235:0] u1_col_in_767;
wire [235:0] u1_col_in_768;
wire [235:0] u1_col_in_769;
wire [235:0] u1_col_in_770;
wire [235:0] u1_col_in_771;
wire [235:0] u1_col_in_772;
wire [235:0] u1_col_in_773;
wire [235:0] u1_col_in_774;
wire [235:0] u1_col_in_775;
wire [235:0] u1_col_in_776;
wire [235:0] u1_col_in_777;
wire [235:0] u1_col_in_778;
wire [235:0] u1_col_in_779;
wire [235:0] u1_col_in_780;
wire [235:0] u1_col_in_781;
wire [235:0] u1_col_in_782;
wire [235:0] u1_col_in_783;
wire [235:0] u1_col_in_784;
wire [235:0] u1_col_in_785;
wire [235:0] u1_col_in_786;
wire [235:0] u1_col_in_787;
wire [235:0] u1_col_in_788;
wire [235:0] u1_col_in_789;
wire [235:0] u1_col_in_790;
wire [235:0] u1_col_in_791;
wire [235:0] u1_col_in_792;
wire [235:0] u1_col_in_793;
wire [235:0] u1_col_in_794;
wire [235:0] u1_col_in_795;
wire [235:0] u1_col_in_796;
wire [235:0] u1_col_in_797;
wire [235:0] u1_col_in_798;
wire [235:0] u1_col_in_799;
wire [235:0] u1_col_in_800;
wire [235:0] u1_col_in_801;
wire [235:0] u1_col_in_802;
wire [235:0] u1_col_in_803;
wire [235:0] u1_col_in_804;
wire [235:0] u1_col_in_805;
wire [235:0] u1_col_in_806;
wire [235:0] u1_col_in_807;
wire [235:0] u1_col_in_808;
wire [235:0] u1_col_in_809;
wire [235:0] u1_col_in_810;
wire [235:0] u1_col_in_811;
wire [235:0] u1_col_in_812;
wire [235:0] u1_col_in_813;
wire [235:0] u1_col_in_814;
wire [235:0] u1_col_in_815;
wire [235:0] u1_col_in_816;
wire [235:0] u1_col_in_817;
wire [235:0] u1_col_in_818;
wire [235:0] u1_col_in_819;
wire [235:0] u1_col_in_820;
wire [235:0] u1_col_in_821;
wire [235:0] u1_col_in_822;
wire [235:0] u1_col_in_823;
wire [235:0] u1_col_in_824;
wire [235:0] u1_col_in_825;
wire [235:0] u1_col_in_826;
wire [235:0] u1_col_in_827;
wire [235:0] u1_col_in_828;
wire [235:0] u1_col_in_829;
wire [235:0] u1_col_in_830;
wire [235:0] u1_col_in_831;
wire [235:0] u1_col_in_832;
wire [235:0] u1_col_in_833;
wire [235:0] u1_col_in_834;
wire [235:0] u1_col_in_835;
wire [235:0] u1_col_in_836;
wire [235:0] u1_col_in_837;
wire [235:0] u1_col_in_838;
wire [235:0] u1_col_in_839;
wire [235:0] u1_col_in_840;
wire [235:0] u1_col_in_841;
wire [235:0] u1_col_in_842;
wire [235:0] u1_col_in_843;
wire [235:0] u1_col_in_844;
wire [235:0] u1_col_in_845;
wire [235:0] u1_col_in_846;
wire [235:0] u1_col_in_847;
wire [235:0] u1_col_in_848;
wire [235:0] u1_col_in_849;
wire [235:0] u1_col_in_850;
wire [235:0] u1_col_in_851;
wire [235:0] u1_col_in_852;
wire [235:0] u1_col_in_853;
wire [235:0] u1_col_in_854;
wire [235:0] u1_col_in_855;
wire [235:0] u1_col_in_856;
wire [235:0] u1_col_in_857;
wire [235:0] u1_col_in_858;
wire [235:0] u1_col_in_859;
wire [235:0] u1_col_in_860;
wire [235:0] u1_col_in_861;
wire [235:0] u1_col_in_862;
wire [235:0] u1_col_in_863;
wire [235:0] u1_col_in_864;
wire [235:0] u1_col_in_865;
wire [235:0] u1_col_in_866;
wire [235:0] u1_col_in_867;
wire [235:0] u1_col_in_868;
wire [235:0] u1_col_in_869;
wire [235:0] u1_col_in_870;
wire [235:0] u1_col_in_871;
wire [235:0] u1_col_in_872;
wire [235:0] u1_col_in_873;
wire [235:0] u1_col_in_874;
wire [235:0] u1_col_in_875;
wire [235:0] u1_col_in_876;
wire [235:0] u1_col_in_877;
wire [235:0] u1_col_in_878;
wire [235:0] u1_col_in_879;
wire [235:0] u1_col_in_880;
wire [235:0] u1_col_in_881;
wire [235:0] u1_col_in_882;
wire [235:0] u1_col_in_883;
wire [235:0] u1_col_in_884;
wire [235:0] u1_col_in_885;
wire [235:0] u1_col_in_886;
wire [235:0] u1_col_in_887;
wire [235:0] u1_col_in_888;
wire [235:0] u1_col_in_889;
wire [235:0] u1_col_in_890;
wire [235:0] u1_col_in_891;
wire [235:0] u1_col_in_892;
wire [235:0] u1_col_in_893;
wire [235:0] u1_col_in_894;
wire [235:0] u1_col_in_895;
wire [235:0] u1_col_in_896;
wire [235:0] u1_col_in_897;
wire [235:0] u1_col_in_898;
wire [235:0] u1_col_in_899;
wire [235:0] u1_col_in_900;
wire [235:0] u1_col_in_901;
wire [235:0] u1_col_in_902;
wire [235:0] u1_col_in_903;
wire [235:0] u1_col_in_904;
wire [235:0] u1_col_in_905;
wire [235:0] u1_col_in_906;
wire [235:0] u1_col_in_907;
wire [235:0] u1_col_in_908;
wire [235:0] u1_col_in_909;
wire [235:0] u1_col_in_910;
wire [235:0] u1_col_in_911;
wire [235:0] u1_col_in_912;
wire [235:0] u1_col_in_913;
wire [235:0] u1_col_in_914;
wire [235:0] u1_col_in_915;
wire [235:0] u1_col_in_916;
wire [235:0] u1_col_in_917;
wire [235:0] u1_col_in_918;
wire [235:0] u1_col_in_919;
wire [235:0] u1_col_in_920;
wire [235:0] u1_col_in_921;
wire [235:0] u1_col_in_922;
wire [235:0] u1_col_in_923;
wire [235:0] u1_col_in_924;
wire [235:0] u1_col_in_925;
wire [235:0] u1_col_in_926;
wire [235:0] u1_col_in_927;
wire [235:0] u1_col_in_928;
wire [235:0] u1_col_in_929;
wire [235:0] u1_col_in_930;
wire [235:0] u1_col_in_931;
wire [235:0] u1_col_in_932;
wire [235:0] u1_col_in_933;
wire [235:0] u1_col_in_934;
wire [235:0] u1_col_in_935;
wire [235:0] u1_col_in_936;
wire [235:0] u1_col_in_937;
wire [235:0] u1_col_in_938;
wire [235:0] u1_col_in_939;
wire [235:0] u1_col_in_940;
wire [235:0] u1_col_in_941;
wire [235:0] u1_col_in_942;
wire [235:0] u1_col_in_943;
wire [235:0] u1_col_in_944;
wire [235:0] u1_col_in_945;
wire [235:0] u1_col_in_946;
wire [235:0] u1_col_in_947;
wire [235:0] u1_col_in_948;
wire [235:0] u1_col_in_949;
wire [235:0] u1_col_in_950;
wire [235:0] u1_col_in_951;
wire [235:0] u1_col_in_952;
wire [235:0] u1_col_in_953;
wire [235:0] u1_col_in_954;
wire [235:0] u1_col_in_955;
wire [235:0] u1_col_in_956;
wire [235:0] u1_col_in_957;
wire [235:0] u1_col_in_958;
wire [235:0] u1_col_in_959;
wire [235:0] u1_col_in_960;
wire [235:0] u1_col_in_961;
wire [235:0] u1_col_in_962;
wire [235:0] u1_col_in_963;
wire [235:0] u1_col_in_964;
wire [235:0] u1_col_in_965;
wire [235:0] u1_col_in_966;
wire [235:0] u1_col_in_967;
wire [235:0] u1_col_in_968;
wire [235:0] u1_col_in_969;
wire [235:0] u1_col_in_970;
wire [235:0] u1_col_in_971;
wire [235:0] u1_col_in_972;
wire [235:0] u1_col_in_973;
wire [235:0] u1_col_in_974;
wire [235:0] u1_col_in_975;
wire [235:0] u1_col_in_976;
wire [235:0] u1_col_in_977;
wire [235:0] u1_col_in_978;
wire [235:0] u1_col_in_979;
wire [235:0] u1_col_in_980;
wire [235:0] u1_col_in_981;
wire [235:0] u1_col_in_982;
wire [235:0] u1_col_in_983;
wire [235:0] u1_col_in_984;
wire [235:0] u1_col_in_985;
wire [235:0] u1_col_in_986;
wire [235:0] u1_col_in_987;
wire [235:0] u1_col_in_988;
wire [235:0] u1_col_in_989;
wire [235:0] u1_col_in_990;
wire [235:0] u1_col_in_991;
wire [235:0] u1_col_in_992;
wire [235:0] u1_col_in_993;
wire [235:0] u1_col_in_994;
wire [235:0] u1_col_in_995;
wire [235:0] u1_col_in_996;
wire [235:0] u1_col_in_997;
wire [235:0] u1_col_in_998;
wire [235:0] u1_col_in_999;
wire [235:0] u1_col_in_1000;
wire [235:0] u1_col_in_1001;
wire [235:0] u1_col_in_1002;
wire [235:0] u1_col_in_1003;
wire [235:0] u1_col_in_1004;
wire [235:0] u1_col_in_1005;
wire [235:0] u1_col_in_1006;
wire [235:0] u1_col_in_1007;
wire [235:0] u1_col_in_1008;
wire [235:0] u1_col_in_1009;
wire [235:0] u1_col_in_1010;
wire [235:0] u1_col_in_1011;
wire [235:0] u1_col_in_1012;
wire [235:0] u1_col_in_1013;
wire [235:0] u1_col_in_1014;
wire [235:0] u1_col_in_1015;
wire [235:0] u1_col_in_1016;
wire [235:0] u1_col_in_1017;
wire [235:0] u1_col_in_1018;
wire [235:0] u1_col_in_1019;
wire [235:0] u1_col_in_1020;
wire [235:0] u1_col_in_1021;
wire [235:0] u1_col_in_1022;
wire [235:0] u1_col_in_1023;
wire [235:0] u1_col_in_1024;
wire [235:0] u1_col_in_1025;
wire [235:0] u1_col_in_1026;
wire [235:0] u1_col_in_1027;
wire [235:0] u1_col_in_1028;
wire [235:0] u1_col_in_1029;
wire [235:0] u1_col_in_1030;
wire [235:0] u1_col_in_1031;
wire [235:0] u1_col_in_1032;
wire [235:0] u1_col_in_1033;
wire [235:0] u1_col_in_1034;
wire [235:0] u1_col_in_1035;
wire [235:0] u1_col_in_1036;
wire [235:0] u1_col_in_1037;
wire [235:0] u1_col_in_1038;
wire [235:0] u1_col_in_1039;
wire [235:0] u1_col_in_1040;
wire [235:0] u1_col_in_1041;
wire [235:0] u1_col_in_1042;
wire [235:0] u1_col_in_1043;
wire [235:0] u1_col_in_1044;
wire [235:0] u1_col_in_1045;
wire [235:0] u1_col_in_1046;
wire [235:0] u1_col_in_1047;
wire [235:0] u1_col_in_1048;
wire [235:0] u1_col_in_1049;
wire [235:0] u1_col_in_1050;
wire [235:0] u1_col_in_1051;
wire [235:0] u1_col_in_1052;
wire [235:0] u1_col_in_1053;
wire [235:0] u1_col_in_1054;
wire [235:0] u1_col_in_1055;
wire [235:0] u1_col_in_1056;
wire [235:0] u1_col_in_1057;
wire [235:0] u1_col_in_1058;
wire [235:0] u1_col_in_1059;
wire [235:0] u1_col_in_1060;
wire [235:0] u1_col_in_1061;
wire [235:0] u1_col_in_1062;
wire [235:0] u1_col_in_1063;
wire [235:0] u1_col_in_1064;
wire [235:0] u1_col_in_1065;
wire [235:0] u1_col_in_1066;
wire [235:0] u1_col_in_1067;
wire [235:0] u1_col_in_1068;
wire [235:0] u1_col_in_1069;
wire [235:0] u1_col_in_1070;
wire [235:0] u1_col_in_1071;
wire [235:0] u1_col_in_1072;
wire [235:0] u1_col_in_1073;
wire [235:0] u1_col_in_1074;
wire [235:0] u1_col_in_1075;
wire [235:0] u1_col_in_1076;
wire [235:0] u1_col_in_1077;
wire [235:0] u1_col_in_1078;
wire [235:0] u1_col_in_1079;
wire [235:0] u1_col_in_1080;
wire [235:0] u1_col_in_1081;
wire [235:0] u1_col_in_1082;
wire [235:0] u1_col_in_1083;
wire [235:0] u1_col_in_1084;
wire [235:0] u1_col_in_1085;
wire [235:0] u1_col_in_1086;
wire [235:0] u1_col_in_1087;
wire [235:0] u1_col_in_1088;
wire [235:0] u1_col_in_1089;
wire [235:0] u1_col_in_1090;
wire [235:0] u1_col_in_1091;
wire [235:0] u1_col_in_1092;
wire [235:0] u1_col_in_1093;
wire [235:0] u1_col_in_1094;
wire [235:0] u1_col_in_1095;
wire [235:0] u1_col_in_1096;
wire [235:0] u1_col_in_1097;
wire [235:0] u1_col_in_1098;
wire [235:0] u1_col_in_1099;
wire [235:0] u1_col_in_1100;
wire [235:0] u1_col_in_1101;
wire [235:0] u1_col_in_1102;
wire [235:0] u1_col_in_1103;
wire [235:0] u1_col_in_1104;
wire [235:0] u1_col_in_1105;
wire [235:0] u1_col_in_1106;
wire [235:0] u1_col_in_1107;
wire [235:0] u1_col_in_1108;
wire [235:0] u1_col_in_1109;
wire [235:0] u1_col_in_1110;
wire [235:0] u1_col_in_1111;
wire [235:0] u1_col_in_1112;
wire [235:0] u1_col_in_1113;
wire [235:0] u1_col_in_1114;
wire [235:0] u1_col_in_1115;
wire [235:0] u1_col_in_1116;
wire [235:0] u1_col_in_1117;
wire [235:0] u1_col_in_1118;
wire [235:0] u1_col_in_1119;
wire [235:0] u1_col_in_1120;
wire [235:0] u1_col_in_1121;
wire [235:0] u1_col_in_1122;
wire [235:0] u1_col_in_1123;
wire [235:0] u1_col_in_1124;
wire [235:0] u1_col_in_1125;
wire [235:0] u1_col_in_1126;
wire [235:0] u1_col_in_1127;
wire [235:0] u1_col_in_1128;
wire [235:0] u1_col_in_1129;
wire [235:0] u1_col_in_1130;
wire [235:0] u1_col_in_1131;
wire [235:0] u1_col_in_1132;
wire [235:0] u1_col_in_1133;
wire [235:0] u1_col_in_1134;
wire [235:0] u1_col_in_1135;
wire [235:0] u1_col_in_1136;
wire [235:0] u1_col_in_1137;
wire [235:0] u1_col_in_1138;
wire [235:0] u1_col_in_1139;
wire [235:0] u1_col_in_1140;
wire [235:0] u1_col_in_1141;
wire [235:0] u1_col_in_1142;
wire [235:0] u1_col_in_1143;
wire [235:0] u1_col_in_1144;
wire [235:0] u1_col_in_1145;
wire [235:0] u1_col_in_1146;
wire [235:0] u1_col_in_1147;
wire [235:0] u1_col_in_1148;
wire [235:0] u1_col_in_1149;
wire [235:0] u1_col_in_1150;
wire [235:0] u1_col_in_1151;
wire [235:0] u1_col_in_1152;
wire [235:0] u1_col_in_1153;
wire [235:0] u1_col_in_1154;
wire [235:0] u1_col_in_1155;
wire [235:0] u1_col_in_1156;
wire [235:0] u1_col_in_1157;
wire [235:0] u1_col_in_1158;
wire [235:0] u1_col_in_1159;
wire [235:0] u1_col_in_1160;
wire [235:0] u1_col_in_1161;
wire [235:0] u1_col_in_1162;
wire [235:0] u1_col_in_1163;
wire [235:0] u1_col_in_1164;
wire [235:0] u1_col_in_1165;
wire [235:0] u1_col_in_1166;
wire [235:0] u1_col_in_1167;
wire [235:0] u1_col_in_1168;
wire [235:0] u1_col_in_1169;
wire [235:0] u1_col_in_1170;
wire [235:0] u1_col_in_1171;
wire [235:0] u1_col_in_1172;
wire [235:0] u1_col_in_1173;
wire [235:0] u1_col_in_1174;
wire [235:0] u1_col_in_1175;
wire [235:0] u1_col_in_1176;
wire [235:0] u1_col_in_1177;
wire [235:0] u1_col_in_1178;
wire [235:0] u1_col_in_1179;
wire [235:0] u1_col_in_1180;
wire [235:0] u1_col_in_1181;
wire [235:0] u1_col_in_1182;
wire [235:0] u1_col_in_1183;
wire [235:0] u1_col_in_1184;
wire [235:0] u1_col_in_1185;
wire [235:0] u1_col_in_1186;
wire [235:0] u1_col_in_1187;
wire [235:0] u1_col_in_1188;
wire [235:0] u1_col_in_1189;
wire [235:0] u1_col_in_1190;
wire [235:0] u1_col_in_1191;
wire [235:0] u1_col_in_1192;
wire [235:0] u1_col_in_1193;
wire [235:0] u1_col_in_1194;
wire [235:0] u1_col_in_1195;
wire [235:0] u1_col_in_1196;
wire [235:0] u1_col_in_1197;
wire [235:0] u1_col_in_1198;
wire [235:0] u1_col_in_1199;
wire [235:0] u1_col_in_1200;
wire [235:0] u1_col_in_1201;
wire [235:0] u1_col_in_1202;
wire [235:0] u1_col_in_1203;
wire [235:0] u1_col_in_1204;
wire [235:0] u1_col_in_1205;
wire [235:0] u1_col_in_1206;
wire [235:0] u1_col_in_1207;
wire [235:0] u1_col_in_1208;
wire [235:0] u1_col_in_1209;
wire [235:0] u1_col_in_1210;
wire [235:0] u1_col_in_1211;
wire [235:0] u1_col_in_1212;
wire [235:0] u1_col_in_1213;
wire [235:0] u1_col_in_1214;
wire [235:0] u1_col_in_1215;
wire [235:0] u1_col_in_1216;
wire [235:0] u1_col_in_1217;
wire [235:0] u1_col_in_1218;
wire [235:0] u1_col_in_1219;
wire [235:0] u1_col_in_1220;
wire [235:0] u1_col_in_1221;
wire [235:0] u1_col_in_1222;
wire [235:0] u1_col_in_1223;
wire [235:0] u1_col_in_1224;
wire [235:0] u1_col_in_1225;
wire [235:0] u1_col_in_1226;
wire [235:0] u1_col_in_1227;
wire [235:0] u1_col_in_1228;
wire [235:0] u1_col_in_1229;
wire [235:0] u1_col_in_1230;
wire [235:0] u1_col_in_1231;
wire [235:0] u1_col_in_1232;
wire [235:0] u1_col_in_1233;
wire [235:0] u1_col_in_1234;
wire [235:0] u1_col_in_1235;
wire [235:0] u1_col_in_1236;
wire [235:0] u1_col_in_1237;
wire [235:0] u1_col_in_1238;
wire [235:0] u1_col_in_1239;
wire [235:0] u1_col_in_1240;
wire [235:0] u1_col_in_1241;
wire [235:0] u1_col_in_1242;
wire [235:0] u1_col_in_1243;
wire [235:0] u1_col_in_1244;
wire [235:0] u1_col_in_1245;
wire [235:0] u1_col_in_1246;
wire [235:0] u1_col_in_1247;
wire [235:0] u1_col_in_1248;
wire [235:0] u1_col_in_1249;
wire [235:0] u1_col_in_1250;
wire [235:0] u1_col_in_1251;
wire [235:0] u1_col_in_1252;
wire [235:0] u1_col_in_1253;
wire [235:0] u1_col_in_1254;
wire [235:0] u1_col_in_1255;
wire [235:0] u1_col_in_1256;
wire [235:0] u1_col_in_1257;
wire [235:0] u1_col_in_1258;
wire [235:0] u1_col_in_1259;
wire [235:0] u1_col_in_1260;
wire [235:0] u1_col_in_1261;
wire [235:0] u1_col_in_1262;
wire [235:0] u1_col_in_1263;
wire [235:0] u1_col_in_1264;
wire [235:0] u1_col_in_1265;
wire [235:0] u1_col_in_1266;
wire [235:0] u1_col_in_1267;
wire [235:0] u1_col_in_1268;
wire [235:0] u1_col_in_1269;
wire [235:0] u1_col_in_1270;
wire [235:0] u1_col_in_1271;
wire [235:0] u1_col_in_1272;
wire [235:0] u1_col_in_1273;
wire [235:0] u1_col_in_1274;
wire [235:0] u1_col_in_1275;
wire [235:0] u1_col_in_1276;
wire [235:0] u1_col_in_1277;
wire [235:0] u1_col_in_1278;
wire [235:0] u1_col_in_1279;


wire [1287:0] u1_row_out_0;
wire [1287:0] u1_row_out_1;


assign u1_col_in_0 = {col_in_0, 108'h0};
assign u1_col_in_1 = {col_in_1, 108'h0};
assign u1_col_in_2 = {col_in_2, 108'h0};
assign u1_col_in_3 = {col_in_3, 108'h0};
assign u1_col_in_4 = {col_in_4, 108'h0};
assign u1_col_in_5 = {col_in_5, 108'h0};
assign u1_col_in_6 = {col_in_6, 108'h0};
assign u1_col_in_7 = {col_in_7, 108'h0};
assign u1_col_in_8 = {col_in_8, 108'h0};
assign u1_col_in_9 = {col_in_9, 108'h0};
assign u1_col_in_10 = {col_in_10, 108'h0};
assign u1_col_in_11 = {col_in_11, 108'h0};
assign u1_col_in_12 = {col_in_12, 108'h0};
assign u1_col_in_13 = {col_in_13, 108'h0};
assign u1_col_in_14 = {col_in_14, 108'h0};
assign u1_col_in_15 = {col_in_15, 108'h0};
assign u1_col_in_16 = {col_in_16, 108'h0};
assign u1_col_in_17 = {col_in_17, 108'h0};
assign u1_col_in_18 = {col_in_18, 108'h0};
assign u1_col_in_19 = {col_in_19, 108'h0};
assign u1_col_in_20 = {col_in_20, 108'h0};
assign u1_col_in_21 = {col_in_21, 108'h0};
assign u1_col_in_22 = {col_in_22, 108'h0};
assign u1_col_in_23 = {col_in_23, 108'h0};
assign u1_col_in_24 = {col_in_24, 108'h0};
assign u1_col_in_25 = {col_in_25, 108'h0};
assign u1_col_in_26 = {col_in_26, 108'h0};
assign u1_col_in_27 = {col_in_27, 108'h0};
assign u1_col_in_28 = {col_in_28, 108'h0};
assign u1_col_in_29 = {col_in_29, 108'h0};
assign u1_col_in_30 = {col_in_30, 108'h0};
assign u1_col_in_31 = {col_in_31, 108'h0};
assign u1_col_in_32 = {col_in_32, 108'h0};
assign u1_col_in_33 = {col_in_33, 108'h0};
assign u1_col_in_34 = {col_in_34, 108'h0};
assign u1_col_in_35 = {col_in_35, 108'h0};
assign u1_col_in_36 = {col_in_36, 108'h0};
assign u1_col_in_37 = {col_in_37, 108'h0};
assign u1_col_in_38 = {col_in_38, 108'h0};
assign u1_col_in_39 = {col_in_39, 108'h0};
assign u1_col_in_40 = {col_in_40, 108'h0};
assign u1_col_in_41 = {col_in_41, 108'h0};
assign u1_col_in_42 = {col_in_42, 108'h0};
assign u1_col_in_43 = {col_in_43, 108'h0};
assign u1_col_in_44 = {col_in_44, 108'h0};
assign u1_col_in_45 = {col_in_45, 108'h0};
assign u1_col_in_46 = {col_in_46, 108'h0};
assign u1_col_in_47 = {col_in_47, 108'h0};
assign u1_col_in_48 = {col_in_48, 108'h0};
assign u1_col_in_49 = {col_in_49, 108'h0};
assign u1_col_in_50 = {col_in_50, 108'h0};
assign u1_col_in_51 = {col_in_51, 108'h0};
assign u1_col_in_52 = {col_in_52, 108'h0};
assign u1_col_in_53 = {col_in_53, 108'h0};
assign u1_col_in_54 = {col_in_54, 108'h0};
assign u1_col_in_55 = {col_in_55, 108'h0};
assign u1_col_in_56 = {col_in_56, 108'h0};
assign u1_col_in_57 = {col_in_57, 108'h0};
assign u1_col_in_58 = {col_in_58, 108'h0};
assign u1_col_in_59 = {col_in_59, 108'h0};
assign u1_col_in_60 = {col_in_60, 108'h0};
assign u1_col_in_61 = {col_in_61, 108'h0};
assign u1_col_in_62 = {col_in_62, 108'h0};
assign u1_col_in_63 = {col_in_63, 108'h0};
assign u1_col_in_64 = {col_in_64, 108'h0};
assign u1_col_in_65 = {col_in_65, 108'h0};
assign u1_col_in_66 = {col_in_66, 108'h0};
assign u1_col_in_67 = {col_in_67, 108'h0};
assign u1_col_in_68 = {col_in_68, 108'h0};
assign u1_col_in_69 = {col_in_69, 108'h0};
assign u1_col_in_70 = {col_in_70, 108'h0};
assign u1_col_in_71 = {col_in_71, 108'h0};
assign u1_col_in_72 = {col_in_72, 108'h0};
assign u1_col_in_73 = {col_in_73, 108'h0};
assign u1_col_in_74 = {col_in_74, 108'h0};
assign u1_col_in_75 = {col_in_75, 108'h0};
assign u1_col_in_76 = {col_in_76, 108'h0};
assign u1_col_in_77 = {col_in_77, 108'h0};
assign u1_col_in_78 = {col_in_78, 108'h0};
assign u1_col_in_79 = {col_in_79, 108'h0};
assign u1_col_in_80 = {col_in_80, 108'h0};
assign u1_col_in_81 = {col_in_81, 108'h0};
assign u1_col_in_82 = {col_in_82, 108'h0};
assign u1_col_in_83 = {col_in_83, 108'h0};
assign u1_col_in_84 = {col_in_84, 108'h0};
assign u1_col_in_85 = {col_in_85, 108'h0};
assign u1_col_in_86 = {col_in_86, 108'h0};
assign u1_col_in_87 = {col_in_87, 108'h0};
assign u1_col_in_88 = {col_in_88, 108'h0};
assign u1_col_in_89 = {col_in_89, 108'h0};
assign u1_col_in_90 = {col_in_90, 108'h0};
assign u1_col_in_91 = {col_in_91, 108'h0};
assign u1_col_in_92 = {col_in_92, 108'h0};
assign u1_col_in_93 = {col_in_93, 108'h0};
assign u1_col_in_94 = {col_in_94, 108'h0};
assign u1_col_in_95 = {col_in_95, 108'h0};
assign u1_col_in_96 = {col_in_96, 108'h0};
assign u1_col_in_97 = {col_in_97, 108'h0};
assign u1_col_in_98 = {col_in_98, 108'h0};
assign u1_col_in_99 = {col_in_99, 108'h0};
assign u1_col_in_100 = {col_in_100, 108'h0};
assign u1_col_in_101 = {col_in_101, 108'h0};
assign u1_col_in_102 = {col_in_102, 108'h0};
assign u1_col_in_103 = {col_in_103, 108'h0};
assign u1_col_in_104 = {col_in_104, 108'h0};
assign u1_col_in_105 = {col_in_105, 108'h0};
assign u1_col_in_106 = {col_in_106, 108'h0};
assign u1_col_in_107 = {col_in_107, 108'h0};
assign u1_col_in_108 = {col_in_108, 108'h0};
assign u1_col_in_109 = {col_in_109, 108'h0};
assign u1_col_in_110 = {col_in_110, 108'h0};
assign u1_col_in_111 = {col_in_111, 108'h0};
assign u1_col_in_112 = {col_in_112, 108'h0};
assign u1_col_in_113 = {col_in_113, 108'h0};
assign u1_col_in_114 = {col_in_114, 108'h0};
assign u1_col_in_115 = {col_in_115, 108'h0};
assign u1_col_in_116 = {col_in_116, 108'h0};
assign u1_col_in_117 = {col_in_117, 108'h0};
assign u1_col_in_118 = {col_in_118, 108'h0};
assign u1_col_in_119 = {col_in_119, 108'h0};
assign u1_col_in_120 = {col_in_120, 108'h0};
assign u1_col_in_121 = {col_in_121, 108'h0};
assign u1_col_in_122 = {col_in_122, 108'h0};
assign u1_col_in_123 = {col_in_123, 108'h0};
assign u1_col_in_124 = {col_in_124, 108'h0};
assign u1_col_in_125 = {col_in_125, 108'h0};
assign u1_col_in_126 = {col_in_126, 108'h0};
assign u1_col_in_127 = {col_in_127, 108'h0};
assign u1_col_in_128 = {col_in_128, 108'h0};
assign u1_col_in_129 = {col_in_129, 108'h0};
assign u1_col_in_130 = {col_in_130, 108'h0};
assign u1_col_in_131 = {col_in_131, 108'h0};
assign u1_col_in_132 = {col_in_132, 108'h0};
assign u1_col_in_133 = {col_in_133, 108'h0};
assign u1_col_in_134 = {col_in_134, 108'h0};
assign u1_col_in_135 = {col_in_135, 108'h0};
assign u1_col_in_136 = {col_in_136, 108'h0};
assign u1_col_in_137 = {col_in_137, 108'h0};
assign u1_col_in_138 = {col_in_138, 108'h0};
assign u1_col_in_139 = {col_in_139, 108'h0};
assign u1_col_in_140 = {col_in_140, 108'h0};
assign u1_col_in_141 = {col_in_141, 108'h0};
assign u1_col_in_142 = {col_in_142, 108'h0};
assign u1_col_in_143 = {col_in_143, 108'h0};
assign u1_col_in_144 = {col_in_144, 108'h0};
assign u1_col_in_145 = {col_in_145, 108'h0};
assign u1_col_in_146 = {col_in_146, 108'h0};
assign u1_col_in_147 = {col_in_147, 108'h0};
assign u1_col_in_148 = {col_in_148, 108'h0};
assign u1_col_in_149 = {col_in_149, 108'h0};
assign u1_col_in_150 = {col_in_150, 108'h0};
assign u1_col_in_151 = {col_in_151, 108'h0};
assign u1_col_in_152 = {col_in_152, 108'h0};
assign u1_col_in_153 = {col_in_153, 108'h0};
assign u1_col_in_154 = {col_in_154, 108'h0};
assign u1_col_in_155 = {col_in_155, 108'h0};
assign u1_col_in_156 = {col_in_156, 108'h0};
assign u1_col_in_157 = {col_in_157, 108'h0};
assign u1_col_in_158 = {col_in_158, 108'h0};
assign u1_col_in_159 = {col_in_159, 108'h0};
assign u1_col_in_160 = {col_in_160, 108'h0};
assign u1_col_in_161 = {col_in_161, 108'h0};
assign u1_col_in_162 = {col_in_162, 108'h0};
assign u1_col_in_163 = {col_in_163, 108'h0};
assign u1_col_in_164 = {col_in_164, 108'h0};
assign u1_col_in_165 = {col_in_165, 108'h0};
assign u1_col_in_166 = {col_in_166, 108'h0};
assign u1_col_in_167 = {col_in_167, 108'h0};
assign u1_col_in_168 = {col_in_168, 108'h0};
assign u1_col_in_169 = {col_in_169, 108'h0};
assign u1_col_in_170 = {col_in_170, 108'h0};
assign u1_col_in_171 = {col_in_171, 108'h0};
assign u1_col_in_172 = {col_in_172, 108'h0};
assign u1_col_in_173 = {col_in_173, 108'h0};
assign u1_col_in_174 = {col_in_174, 108'h0};
assign u1_col_in_175 = {col_in_175, 108'h0};
assign u1_col_in_176 = {col_in_176, 108'h0};
assign u1_col_in_177 = {col_in_177, 108'h0};
assign u1_col_in_178 = {col_in_178, 108'h0};
assign u1_col_in_179 = {col_in_179, 108'h0};
assign u1_col_in_180 = {col_in_180, 108'h0};
assign u1_col_in_181 = {col_in_181, 108'h0};
assign u1_col_in_182 = {col_in_182, 108'h0};
assign u1_col_in_183 = {col_in_183, 108'h0};
assign u1_col_in_184 = {col_in_184, 108'h0};
assign u1_col_in_185 = {col_in_185, 108'h0};
assign u1_col_in_186 = {col_in_186, 108'h0};
assign u1_col_in_187 = {col_in_187, 108'h0};
assign u1_col_in_188 = {col_in_188, 108'h0};
assign u1_col_in_189 = {col_in_189, 108'h0};
assign u1_col_in_190 = {col_in_190, 108'h0};
assign u1_col_in_191 = {col_in_191, 108'h0};
assign u1_col_in_192 = {col_in_192, 108'h0};
assign u1_col_in_193 = {col_in_193, 108'h0};
assign u1_col_in_194 = {col_in_194, 108'h0};
assign u1_col_in_195 = {col_in_195, 108'h0};
assign u1_col_in_196 = {col_in_196, 108'h0};
assign u1_col_in_197 = {col_in_197, 108'h0};
assign u1_col_in_198 = {col_in_198, 108'h0};
assign u1_col_in_199 = {col_in_199, 108'h0};
assign u1_col_in_200 = {col_in_200, 108'h0};
assign u1_col_in_201 = {col_in_201, 108'h0};
assign u1_col_in_202 = {col_in_202, 108'h0};
assign u1_col_in_203 = {col_in_203, 108'h0};
assign u1_col_in_204 = {col_in_204, 108'h0};
assign u1_col_in_205 = {col_in_205, 108'h0};
assign u1_col_in_206 = {col_in_206, 108'h0};
assign u1_col_in_207 = {col_in_207, 108'h0};
assign u1_col_in_208 = {col_in_208, 108'h0};
assign u1_col_in_209 = {col_in_209, 108'h0};
assign u1_col_in_210 = {col_in_210, 108'h0};
assign u1_col_in_211 = {col_in_211, 108'h0};
assign u1_col_in_212 = {col_in_212, 108'h0};
assign u1_col_in_213 = {col_in_213, 108'h0};
assign u1_col_in_214 = {col_in_214, 108'h0};
assign u1_col_in_215 = {col_in_215, 108'h0};
assign u1_col_in_216 = {col_in_216, 108'h0};
assign u1_col_in_217 = {col_in_217, 108'h0};
assign u1_col_in_218 = {col_in_218, 108'h0};
assign u1_col_in_219 = {col_in_219, 108'h0};
assign u1_col_in_220 = {col_in_220, 108'h0};
assign u1_col_in_221 = {col_in_221, 108'h0};
assign u1_col_in_222 = {col_in_222, 108'h0};
assign u1_col_in_223 = {col_in_223, 108'h0};
assign u1_col_in_224 = {col_in_224, 108'h0};
assign u1_col_in_225 = {col_in_225, 108'h0};
assign u1_col_in_226 = {col_in_226, 108'h0};
assign u1_col_in_227 = {col_in_227, 108'h0};
assign u1_col_in_228 = {col_in_228, 108'h0};
assign u1_col_in_229 = {col_in_229, 108'h0};
assign u1_col_in_230 = {col_in_230, 108'h0};
assign u1_col_in_231 = {col_in_231, 108'h0};
assign u1_col_in_232 = {col_in_232, 108'h0};
assign u1_col_in_233 = {col_in_233, 108'h0};
assign u1_col_in_234 = {col_in_234, 108'h0};
assign u1_col_in_235 = {col_in_235, 108'h0};
assign u1_col_in_236 = {col_in_236, 108'h0};
assign u1_col_in_237 = {col_in_237, 108'h0};
assign u1_col_in_238 = {col_in_238, 108'h0};
assign u1_col_in_239 = {col_in_239, 108'h0};
assign u1_col_in_240 = {col_in_240, 108'h0};
assign u1_col_in_241 = {col_in_241, 108'h0};
assign u1_col_in_242 = {col_in_242, 108'h0};
assign u1_col_in_243 = {col_in_243, 108'h0};
assign u1_col_in_244 = {col_in_244, 108'h0};
assign u1_col_in_245 = {col_in_245, 108'h0};
assign u1_col_in_246 = {col_in_246, 108'h0};
assign u1_col_in_247 = {col_in_247, 108'h0};
assign u1_col_in_248 = {col_in_248, 108'h0};
assign u1_col_in_249 = {col_in_249, 108'h0};
assign u1_col_in_250 = {col_in_250, 108'h0};
assign u1_col_in_251 = {col_in_251, 108'h0};
assign u1_col_in_252 = {col_in_252, 108'h0};
assign u1_col_in_253 = {col_in_253, 108'h0};
assign u1_col_in_254 = {col_in_254, 108'h0};
assign u1_col_in_255 = {col_in_255, 108'h0};
assign u1_col_in_256 = {col_in_256, u0_col_out_0, reg_intermediate0[0], reg_intermediate1[0]};
assign u1_col_in_257 = {col_in_257, u0_col_out_1, reg_intermediate0[1], reg_intermediate1[1]};
assign u1_col_in_258 = {col_in_258, u0_col_out_2, reg_intermediate0[2], reg_intermediate1[2]};
assign u1_col_in_259 = {col_in_259, u0_col_out_3, reg_intermediate0[3], reg_intermediate1[3]};
assign u1_col_in_260 = {col_in_260, u0_col_out_4, reg_intermediate0[4], reg_intermediate1[4]};
assign u1_col_in_261 = {col_in_261, u0_col_out_5, reg_intermediate0[5], reg_intermediate1[5]};
assign u1_col_in_262 = {col_in_262, u0_col_out_6, reg_intermediate0[6], reg_intermediate1[6]};
assign u1_col_in_263 = {col_in_263, u0_col_out_7, reg_intermediate0[7], reg_intermediate1[7]};
assign u1_col_in_264 = {col_in_264, u0_col_out_8, reg_intermediate0[8], reg_intermediate1[8]};
assign u1_col_in_265 = {col_in_265, u0_col_out_9, reg_intermediate0[9], reg_intermediate1[9]};
assign u1_col_in_266 = {col_in_266, u0_col_out_10, reg_intermediate0[10], reg_intermediate1[10]};
assign u1_col_in_267 = {col_in_267, u0_col_out_11, reg_intermediate0[11], reg_intermediate1[11]};
assign u1_col_in_268 = {col_in_268, u0_col_out_12, reg_intermediate0[12], reg_intermediate1[12]};
assign u1_col_in_269 = {col_in_269, u0_col_out_13, reg_intermediate0[13], reg_intermediate1[13]};
assign u1_col_in_270 = {col_in_270, u0_col_out_14, reg_intermediate0[14], reg_intermediate1[14]};
assign u1_col_in_271 = {col_in_271, u0_col_out_15, reg_intermediate0[15], reg_intermediate1[15]};
assign u1_col_in_272 = {col_in_272, u0_col_out_16, reg_intermediate0[16], reg_intermediate1[16]};
assign u1_col_in_273 = {col_in_273, u0_col_out_17, reg_intermediate0[17], reg_intermediate1[17]};
assign u1_col_in_274 = {col_in_274, u0_col_out_18, reg_intermediate0[18], reg_intermediate1[18]};
assign u1_col_in_275 = {col_in_275, u0_col_out_19, reg_intermediate0[19], reg_intermediate1[19]};
assign u1_col_in_276 = {col_in_276, u0_col_out_20, reg_intermediate0[20], reg_intermediate1[20]};
assign u1_col_in_277 = {col_in_277, u0_col_out_21, reg_intermediate0[21], reg_intermediate1[21]};
assign u1_col_in_278 = {col_in_278, u0_col_out_22, reg_intermediate0[22], reg_intermediate1[22]};
assign u1_col_in_279 = {col_in_279, u0_col_out_23, reg_intermediate0[23], reg_intermediate1[23]};
assign u1_col_in_280 = {col_in_280, u0_col_out_24, reg_intermediate0[24], reg_intermediate1[24]};
assign u1_col_in_281 = {col_in_281, u0_col_out_25, reg_intermediate0[25], reg_intermediate1[25]};
assign u1_col_in_282 = {col_in_282, u0_col_out_26, reg_intermediate0[26], reg_intermediate1[26]};
assign u1_col_in_283 = {col_in_283, u0_col_out_27, reg_intermediate0[27], reg_intermediate1[27]};
assign u1_col_in_284 = {col_in_284, u0_col_out_28, reg_intermediate0[28], reg_intermediate1[28]};
assign u1_col_in_285 = {col_in_285, u0_col_out_29, reg_intermediate0[29], reg_intermediate1[29]};
assign u1_col_in_286 = {col_in_286, u0_col_out_30, reg_intermediate0[30], reg_intermediate1[30]};
assign u1_col_in_287 = {col_in_287, u0_col_out_31, reg_intermediate0[31], reg_intermediate1[31]};
assign u1_col_in_288 = {col_in_288, u0_col_out_32, reg_intermediate0[32], reg_intermediate1[32]};
assign u1_col_in_289 = {col_in_289, u0_col_out_33, reg_intermediate0[33], reg_intermediate1[33]};
assign u1_col_in_290 = {col_in_290, u0_col_out_34, reg_intermediate0[34], reg_intermediate1[34]};
assign u1_col_in_291 = {col_in_291, u0_col_out_35, reg_intermediate0[35], reg_intermediate1[35]};
assign u1_col_in_292 = {col_in_292, u0_col_out_36, reg_intermediate0[36], reg_intermediate1[36]};
assign u1_col_in_293 = {col_in_293, u0_col_out_37, reg_intermediate0[37], reg_intermediate1[37]};
assign u1_col_in_294 = {col_in_294, u0_col_out_38, reg_intermediate0[38], reg_intermediate1[38]};
assign u1_col_in_295 = {col_in_295, u0_col_out_39, reg_intermediate0[39], reg_intermediate1[39]};
assign u1_col_in_296 = {col_in_296, u0_col_out_40, reg_intermediate0[40], reg_intermediate1[40]};
assign u1_col_in_297 = {col_in_297, u0_col_out_41, reg_intermediate0[41], reg_intermediate1[41]};
assign u1_col_in_298 = {col_in_298, u0_col_out_42, reg_intermediate0[42], reg_intermediate1[42]};
assign u1_col_in_299 = {col_in_299, u0_col_out_43, reg_intermediate0[43], reg_intermediate1[43]};
assign u1_col_in_300 = {col_in_300, u0_col_out_44, reg_intermediate0[44], reg_intermediate1[44]};
assign u1_col_in_301 = {col_in_301, u0_col_out_45, reg_intermediate0[45], reg_intermediate1[45]};
assign u1_col_in_302 = {col_in_302, u0_col_out_46, reg_intermediate0[46], reg_intermediate1[46]};
assign u1_col_in_303 = {col_in_303, u0_col_out_47, reg_intermediate0[47], reg_intermediate1[47]};
assign u1_col_in_304 = {col_in_304, u0_col_out_48, reg_intermediate0[48], reg_intermediate1[48]};
assign u1_col_in_305 = {col_in_305, u0_col_out_49, reg_intermediate0[49], reg_intermediate1[49]};
assign u1_col_in_306 = {col_in_306, u0_col_out_50, reg_intermediate0[50], reg_intermediate1[50]};
assign u1_col_in_307 = {col_in_307, u0_col_out_51, reg_intermediate0[51], reg_intermediate1[51]};
assign u1_col_in_308 = {col_in_308, u0_col_out_52, reg_intermediate0[52], reg_intermediate1[52]};
assign u1_col_in_309 = {col_in_309, u0_col_out_53, reg_intermediate0[53], reg_intermediate1[53]};
assign u1_col_in_310 = {col_in_310, u0_col_out_54, reg_intermediate0[54], reg_intermediate1[54]};
assign u1_col_in_311 = {col_in_311, u0_col_out_55, reg_intermediate0[55], reg_intermediate1[55]};
assign u1_col_in_312 = {col_in_312, u0_col_out_56, reg_intermediate0[56], reg_intermediate1[56]};
assign u1_col_in_313 = {col_in_313, u0_col_out_57, reg_intermediate0[57], reg_intermediate1[57]};
assign u1_col_in_314 = {col_in_314, u0_col_out_58, reg_intermediate0[58], reg_intermediate1[58]};
assign u1_col_in_315 = {col_in_315, u0_col_out_59, reg_intermediate0[59], reg_intermediate1[59]};
assign u1_col_in_316 = {col_in_316, u0_col_out_60, reg_intermediate0[60], reg_intermediate1[60]};
assign u1_col_in_317 = {col_in_317, u0_col_out_61, reg_intermediate0[61], reg_intermediate1[61]};
assign u1_col_in_318 = {col_in_318, u0_col_out_62, reg_intermediate0[62], reg_intermediate1[62]};
assign u1_col_in_319 = {col_in_319, u0_col_out_63, reg_intermediate0[63], reg_intermediate1[63]};
assign u1_col_in_320 = {col_in_320, u0_col_out_64, reg_intermediate0[64], reg_intermediate1[64]};
assign u1_col_in_321 = {col_in_321, u0_col_out_65, reg_intermediate0[65], reg_intermediate1[65]};
assign u1_col_in_322 = {col_in_322, u0_col_out_66, reg_intermediate0[66], reg_intermediate1[66]};
assign u1_col_in_323 = {col_in_323, u0_col_out_67, reg_intermediate0[67], reg_intermediate1[67]};
assign u1_col_in_324 = {col_in_324, u0_col_out_68, reg_intermediate0[68], reg_intermediate1[68]};
assign u1_col_in_325 = {col_in_325, u0_col_out_69, reg_intermediate0[69], reg_intermediate1[69]};
assign u1_col_in_326 = {col_in_326, u0_col_out_70, reg_intermediate0[70], reg_intermediate1[70]};
assign u1_col_in_327 = {col_in_327, u0_col_out_71, reg_intermediate0[71], reg_intermediate1[71]};
assign u1_col_in_328 = {col_in_328, u0_col_out_72, reg_intermediate0[72], reg_intermediate1[72]};
assign u1_col_in_329 = {col_in_329, u0_col_out_73, reg_intermediate0[73], reg_intermediate1[73]};
assign u1_col_in_330 = {col_in_330, u0_col_out_74, reg_intermediate0[74], reg_intermediate1[74]};
assign u1_col_in_331 = {col_in_331, u0_col_out_75, reg_intermediate0[75], reg_intermediate1[75]};
assign u1_col_in_332 = {col_in_332, u0_col_out_76, reg_intermediate0[76], reg_intermediate1[76]};
assign u1_col_in_333 = {col_in_333, u0_col_out_77, reg_intermediate0[77], reg_intermediate1[77]};
assign u1_col_in_334 = {col_in_334, u0_col_out_78, reg_intermediate0[78], reg_intermediate1[78]};
assign u1_col_in_335 = {col_in_335, u0_col_out_79, reg_intermediate0[79], reg_intermediate1[79]};
assign u1_col_in_336 = {col_in_336, u0_col_out_80, reg_intermediate0[80], reg_intermediate1[80]};
assign u1_col_in_337 = {col_in_337, u0_col_out_81, reg_intermediate0[81], reg_intermediate1[81]};
assign u1_col_in_338 = {col_in_338, u0_col_out_82, reg_intermediate0[82], reg_intermediate1[82]};
assign u1_col_in_339 = {col_in_339, u0_col_out_83, reg_intermediate0[83], reg_intermediate1[83]};
assign u1_col_in_340 = {col_in_340, u0_col_out_84, reg_intermediate0[84], reg_intermediate1[84]};
assign u1_col_in_341 = {col_in_341, u0_col_out_85, reg_intermediate0[85], reg_intermediate1[85]};
assign u1_col_in_342 = {col_in_342, u0_col_out_86, reg_intermediate0[86], reg_intermediate1[86]};
assign u1_col_in_343 = {col_in_343, u0_col_out_87, reg_intermediate0[87], reg_intermediate1[87]};
assign u1_col_in_344 = {col_in_344, u0_col_out_88, reg_intermediate0[88], reg_intermediate1[88]};
assign u1_col_in_345 = {col_in_345, u0_col_out_89, reg_intermediate0[89], reg_intermediate1[89]};
assign u1_col_in_346 = {col_in_346, u0_col_out_90, reg_intermediate0[90], reg_intermediate1[90]};
assign u1_col_in_347 = {col_in_347, u0_col_out_91, reg_intermediate0[91], reg_intermediate1[91]};
assign u1_col_in_348 = {col_in_348, u0_col_out_92, reg_intermediate0[92], reg_intermediate1[92]};
assign u1_col_in_349 = {col_in_349, u0_col_out_93, reg_intermediate0[93], reg_intermediate1[93]};
assign u1_col_in_350 = {col_in_350, u0_col_out_94, reg_intermediate0[94], reg_intermediate1[94]};
assign u1_col_in_351 = {col_in_351, u0_col_out_95, reg_intermediate0[95], reg_intermediate1[95]};
assign u1_col_in_352 = {col_in_352, u0_col_out_96, reg_intermediate0[96], reg_intermediate1[96]};
assign u1_col_in_353 = {col_in_353, u0_col_out_97, reg_intermediate0[97], reg_intermediate1[97]};
assign u1_col_in_354 = {col_in_354, u0_col_out_98, reg_intermediate0[98], reg_intermediate1[98]};
assign u1_col_in_355 = {col_in_355, u0_col_out_99, reg_intermediate0[99], reg_intermediate1[99]};
assign u1_col_in_356 = {col_in_356, u0_col_out_100, reg_intermediate0[100], reg_intermediate1[100]};
assign u1_col_in_357 = {col_in_357, u0_col_out_101, reg_intermediate0[101], reg_intermediate1[101]};
assign u1_col_in_358 = {col_in_358, u0_col_out_102, reg_intermediate0[102], reg_intermediate1[102]};
assign u1_col_in_359 = {col_in_359, u0_col_out_103, reg_intermediate0[103], reg_intermediate1[103]};
assign u1_col_in_360 = {col_in_360, u0_col_out_104, reg_intermediate0[104], reg_intermediate1[104]};
assign u1_col_in_361 = {col_in_361, u0_col_out_105, reg_intermediate0[105], reg_intermediate1[105]};
assign u1_col_in_362 = {col_in_362, u0_col_out_106, reg_intermediate0[106], reg_intermediate1[106]};
assign u1_col_in_363 = {col_in_363, u0_col_out_107, reg_intermediate0[107], reg_intermediate1[107]};
assign u1_col_in_364 = {col_in_364, u0_col_out_108, reg_intermediate0[108], reg_intermediate1[108]};
assign u1_col_in_365 = {col_in_365, u0_col_out_109, reg_intermediate0[109], reg_intermediate1[109]};
assign u1_col_in_366 = {col_in_366, u0_col_out_110, reg_intermediate0[110], reg_intermediate1[110]};
assign u1_col_in_367 = {col_in_367, u0_col_out_111, reg_intermediate0[111], reg_intermediate1[111]};
assign u1_col_in_368 = {col_in_368, u0_col_out_112, reg_intermediate0[112], reg_intermediate1[112]};
assign u1_col_in_369 = {col_in_369, u0_col_out_113, reg_intermediate0[113], reg_intermediate1[113]};
assign u1_col_in_370 = {col_in_370, u0_col_out_114, reg_intermediate0[114], reg_intermediate1[114]};
assign u1_col_in_371 = {col_in_371, u0_col_out_115, reg_intermediate0[115], reg_intermediate1[115]};
assign u1_col_in_372 = {col_in_372, u0_col_out_116, reg_intermediate0[116], reg_intermediate1[116]};
assign u1_col_in_373 = {col_in_373, u0_col_out_117, reg_intermediate0[117], reg_intermediate1[117]};
assign u1_col_in_374 = {col_in_374, u0_col_out_118, reg_intermediate0[118], reg_intermediate1[118]};
assign u1_col_in_375 = {col_in_375, u0_col_out_119, reg_intermediate0[119], reg_intermediate1[119]};
assign u1_col_in_376 = {col_in_376, u0_col_out_120, reg_intermediate0[120], reg_intermediate1[120]};
assign u1_col_in_377 = {col_in_377, u0_col_out_121, reg_intermediate0[121], reg_intermediate1[121]};
assign u1_col_in_378 = {col_in_378, u0_col_out_122, reg_intermediate0[122], reg_intermediate1[122]};
assign u1_col_in_379 = {col_in_379, u0_col_out_123, reg_intermediate0[123], reg_intermediate1[123]};
assign u1_col_in_380 = {col_in_380, u0_col_out_124, reg_intermediate0[124], reg_intermediate1[124]};
assign u1_col_in_381 = {col_in_381, u0_col_out_125, reg_intermediate0[125], reg_intermediate1[125]};
assign u1_col_in_382 = {col_in_382, u0_col_out_126, reg_intermediate0[126], reg_intermediate1[126]};
assign u1_col_in_383 = {col_in_383, u0_col_out_127, reg_intermediate0[127], reg_intermediate1[127]};
assign u1_col_in_384 = {col_in_384, u0_col_out_128, reg_intermediate0[128], reg_intermediate1[128]};
assign u1_col_in_385 = {col_in_385, u0_col_out_129, reg_intermediate0[129], reg_intermediate1[129]};
assign u1_col_in_386 = {col_in_386, u0_col_out_130, reg_intermediate0[130], reg_intermediate1[130]};
assign u1_col_in_387 = {col_in_387, u0_col_out_131, reg_intermediate0[131], reg_intermediate1[131]};
assign u1_col_in_388 = {col_in_388, u0_col_out_132, reg_intermediate0[132], reg_intermediate1[132]};
assign u1_col_in_389 = {col_in_389, u0_col_out_133, reg_intermediate0[133], reg_intermediate1[133]};
assign u1_col_in_390 = {col_in_390, u0_col_out_134, reg_intermediate0[134], reg_intermediate1[134]};
assign u1_col_in_391 = {col_in_391, u0_col_out_135, reg_intermediate0[135], reg_intermediate1[135]};
assign u1_col_in_392 = {col_in_392, u0_col_out_136, reg_intermediate0[136], reg_intermediate1[136]};
assign u1_col_in_393 = {col_in_393, u0_col_out_137, reg_intermediate0[137], reg_intermediate1[137]};
assign u1_col_in_394 = {col_in_394, u0_col_out_138, reg_intermediate0[138], reg_intermediate1[138]};
assign u1_col_in_395 = {col_in_395, u0_col_out_139, reg_intermediate0[139], reg_intermediate1[139]};
assign u1_col_in_396 = {col_in_396, u0_col_out_140, reg_intermediate0[140], reg_intermediate1[140]};
assign u1_col_in_397 = {col_in_397, u0_col_out_141, reg_intermediate0[141], reg_intermediate1[141]};
assign u1_col_in_398 = {col_in_398, u0_col_out_142, reg_intermediate0[142], reg_intermediate1[142]};
assign u1_col_in_399 = {col_in_399, u0_col_out_143, reg_intermediate0[143], reg_intermediate1[143]};
assign u1_col_in_400 = {col_in_400, u0_col_out_144, reg_intermediate0[144], reg_intermediate1[144]};
assign u1_col_in_401 = {col_in_401, u0_col_out_145, reg_intermediate0[145], reg_intermediate1[145]};
assign u1_col_in_402 = {col_in_402, u0_col_out_146, reg_intermediate0[146], reg_intermediate1[146]};
assign u1_col_in_403 = {col_in_403, u0_col_out_147, reg_intermediate0[147], reg_intermediate1[147]};
assign u1_col_in_404 = {col_in_404, u0_col_out_148, reg_intermediate0[148], reg_intermediate1[148]};
assign u1_col_in_405 = {col_in_405, u0_col_out_149, reg_intermediate0[149], reg_intermediate1[149]};
assign u1_col_in_406 = {col_in_406, u0_col_out_150, reg_intermediate0[150], reg_intermediate1[150]};
assign u1_col_in_407 = {col_in_407, u0_col_out_151, reg_intermediate0[151], reg_intermediate1[151]};
assign u1_col_in_408 = {col_in_408, u0_col_out_152, reg_intermediate0[152], reg_intermediate1[152]};
assign u1_col_in_409 = {col_in_409, u0_col_out_153, reg_intermediate0[153], reg_intermediate1[153]};
assign u1_col_in_410 = {col_in_410, u0_col_out_154, reg_intermediate0[154], reg_intermediate1[154]};
assign u1_col_in_411 = {col_in_411, u0_col_out_155, reg_intermediate0[155], reg_intermediate1[155]};
assign u1_col_in_412 = {col_in_412, u0_col_out_156, reg_intermediate0[156], reg_intermediate1[156]};
assign u1_col_in_413 = {col_in_413, u0_col_out_157, reg_intermediate0[157], reg_intermediate1[157]};
assign u1_col_in_414 = {col_in_414, u0_col_out_158, reg_intermediate0[158], reg_intermediate1[158]};
assign u1_col_in_415 = {col_in_415, u0_col_out_159, reg_intermediate0[159], reg_intermediate1[159]};
assign u1_col_in_416 = {col_in_416, u0_col_out_160, reg_intermediate0[160], reg_intermediate1[160]};
assign u1_col_in_417 = {col_in_417, u0_col_out_161, reg_intermediate0[161], reg_intermediate1[161]};
assign u1_col_in_418 = {col_in_418, u0_col_out_162, reg_intermediate0[162], reg_intermediate1[162]};
assign u1_col_in_419 = {col_in_419, u0_col_out_163, reg_intermediate0[163], reg_intermediate1[163]};
assign u1_col_in_420 = {col_in_420, u0_col_out_164, reg_intermediate0[164], reg_intermediate1[164]};
assign u1_col_in_421 = {col_in_421, u0_col_out_165, reg_intermediate0[165], reg_intermediate1[165]};
assign u1_col_in_422 = {col_in_422, u0_col_out_166, reg_intermediate0[166], reg_intermediate1[166]};
assign u1_col_in_423 = {col_in_423, u0_col_out_167, reg_intermediate0[167], reg_intermediate1[167]};
assign u1_col_in_424 = {col_in_424, u0_col_out_168, reg_intermediate0[168], reg_intermediate1[168]};
assign u1_col_in_425 = {col_in_425, u0_col_out_169, reg_intermediate0[169], reg_intermediate1[169]};
assign u1_col_in_426 = {col_in_426, u0_col_out_170, reg_intermediate0[170], reg_intermediate1[170]};
assign u1_col_in_427 = {col_in_427, u0_col_out_171, reg_intermediate0[171], reg_intermediate1[171]};
assign u1_col_in_428 = {col_in_428, u0_col_out_172, reg_intermediate0[172], reg_intermediate1[172]};
assign u1_col_in_429 = {col_in_429, u0_col_out_173, reg_intermediate0[173], reg_intermediate1[173]};
assign u1_col_in_430 = {col_in_430, u0_col_out_174, reg_intermediate0[174], reg_intermediate1[174]};
assign u1_col_in_431 = {col_in_431, u0_col_out_175, reg_intermediate0[175], reg_intermediate1[175]};
assign u1_col_in_432 = {col_in_432, u0_col_out_176, reg_intermediate0[176], reg_intermediate1[176]};
assign u1_col_in_433 = {col_in_433, u0_col_out_177, reg_intermediate0[177], reg_intermediate1[177]};
assign u1_col_in_434 = {col_in_434, u0_col_out_178, reg_intermediate0[178], reg_intermediate1[178]};
assign u1_col_in_435 = {col_in_435, u0_col_out_179, reg_intermediate0[179], reg_intermediate1[179]};
assign u1_col_in_436 = {col_in_436, u0_col_out_180, reg_intermediate0[180], reg_intermediate1[180]};
assign u1_col_in_437 = {col_in_437, u0_col_out_181, reg_intermediate0[181], reg_intermediate1[181]};
assign u1_col_in_438 = {col_in_438, u0_col_out_182, reg_intermediate0[182], reg_intermediate1[182]};
assign u1_col_in_439 = {col_in_439, u0_col_out_183, reg_intermediate0[183], reg_intermediate1[183]};
assign u1_col_in_440 = {col_in_440, u0_col_out_184, reg_intermediate0[184], reg_intermediate1[184]};
assign u1_col_in_441 = {col_in_441, u0_col_out_185, reg_intermediate0[185], reg_intermediate1[185]};
assign u1_col_in_442 = {col_in_442, u0_col_out_186, reg_intermediate0[186], reg_intermediate1[186]};
assign u1_col_in_443 = {col_in_443, u0_col_out_187, reg_intermediate0[187], reg_intermediate1[187]};
assign u1_col_in_444 = {col_in_444, u0_col_out_188, reg_intermediate0[188], reg_intermediate1[188]};
assign u1_col_in_445 = {col_in_445, u0_col_out_189, reg_intermediate0[189], reg_intermediate1[189]};
assign u1_col_in_446 = {col_in_446, u0_col_out_190, reg_intermediate0[190], reg_intermediate1[190]};
assign u1_col_in_447 = {col_in_447, u0_col_out_191, reg_intermediate0[191], reg_intermediate1[191]};
assign u1_col_in_448 = {col_in_448, u0_col_out_192, reg_intermediate0[192], reg_intermediate1[192]};
assign u1_col_in_449 = {col_in_449, u0_col_out_193, reg_intermediate0[193], reg_intermediate1[193]};
assign u1_col_in_450 = {col_in_450, u0_col_out_194, reg_intermediate0[194], reg_intermediate1[194]};
assign u1_col_in_451 = {col_in_451, u0_col_out_195, reg_intermediate0[195], reg_intermediate1[195]};
assign u1_col_in_452 = {col_in_452, u0_col_out_196, reg_intermediate0[196], reg_intermediate1[196]};
assign u1_col_in_453 = {col_in_453, u0_col_out_197, reg_intermediate0[197], reg_intermediate1[197]};
assign u1_col_in_454 = {col_in_454, u0_col_out_198, reg_intermediate0[198], reg_intermediate1[198]};
assign u1_col_in_455 = {col_in_455, u0_col_out_199, reg_intermediate0[199], reg_intermediate1[199]};
assign u1_col_in_456 = {col_in_456, u0_col_out_200, reg_intermediate0[200], reg_intermediate1[200]};
assign u1_col_in_457 = {col_in_457, u0_col_out_201, reg_intermediate0[201], reg_intermediate1[201]};
assign u1_col_in_458 = {col_in_458, u0_col_out_202, reg_intermediate0[202], reg_intermediate1[202]};
assign u1_col_in_459 = {col_in_459, u0_col_out_203, reg_intermediate0[203], reg_intermediate1[203]};
assign u1_col_in_460 = {col_in_460, u0_col_out_204, reg_intermediate0[204], reg_intermediate1[204]};
assign u1_col_in_461 = {col_in_461, u0_col_out_205, reg_intermediate0[205], reg_intermediate1[205]};
assign u1_col_in_462 = {col_in_462, u0_col_out_206, reg_intermediate0[206], reg_intermediate1[206]};
assign u1_col_in_463 = {col_in_463, u0_col_out_207, reg_intermediate0[207], reg_intermediate1[207]};
assign u1_col_in_464 = {col_in_464, u0_col_out_208, reg_intermediate0[208], reg_intermediate1[208]};
assign u1_col_in_465 = {col_in_465, u0_col_out_209, reg_intermediate0[209], reg_intermediate1[209]};
assign u1_col_in_466 = {col_in_466, u0_col_out_210, reg_intermediate0[210], reg_intermediate1[210]};
assign u1_col_in_467 = {col_in_467, u0_col_out_211, reg_intermediate0[211], reg_intermediate1[211]};
assign u1_col_in_468 = {col_in_468, u0_col_out_212, reg_intermediate0[212], reg_intermediate1[212]};
assign u1_col_in_469 = {col_in_469, u0_col_out_213, reg_intermediate0[213], reg_intermediate1[213]};
assign u1_col_in_470 = {col_in_470, u0_col_out_214, reg_intermediate0[214], reg_intermediate1[214]};
assign u1_col_in_471 = {col_in_471, u0_col_out_215, reg_intermediate0[215], reg_intermediate1[215]};
assign u1_col_in_472 = {col_in_472, u0_col_out_216, reg_intermediate0[216], reg_intermediate1[216]};
assign u1_col_in_473 = {col_in_473, u0_col_out_217, reg_intermediate0[217], reg_intermediate1[217]};
assign u1_col_in_474 = {col_in_474, u0_col_out_218, reg_intermediate0[218], reg_intermediate1[218]};
assign u1_col_in_475 = {col_in_475, u0_col_out_219, reg_intermediate0[219], reg_intermediate1[219]};
assign u1_col_in_476 = {col_in_476, u0_col_out_220, reg_intermediate0[220], reg_intermediate1[220]};
assign u1_col_in_477 = {col_in_477, u0_col_out_221, reg_intermediate0[221], reg_intermediate1[221]};
assign u1_col_in_478 = {col_in_478, u0_col_out_222, reg_intermediate0[222], reg_intermediate1[222]};
assign u1_col_in_479 = {col_in_479, u0_col_out_223, reg_intermediate0[223], reg_intermediate1[223]};
assign u1_col_in_480 = {col_in_480, u0_col_out_224, reg_intermediate0[224], reg_intermediate1[224]};
assign u1_col_in_481 = {col_in_481, u0_col_out_225, reg_intermediate0[225], reg_intermediate1[225]};
assign u1_col_in_482 = {col_in_482, u0_col_out_226, reg_intermediate0[226], reg_intermediate1[226]};
assign u1_col_in_483 = {col_in_483, u0_col_out_227, reg_intermediate0[227], reg_intermediate1[227]};
assign u1_col_in_484 = {col_in_484, u0_col_out_228, reg_intermediate0[228], reg_intermediate1[228]};
assign u1_col_in_485 = {col_in_485, u0_col_out_229, reg_intermediate0[229], reg_intermediate1[229]};
assign u1_col_in_486 = {col_in_486, u0_col_out_230, reg_intermediate0[230], reg_intermediate1[230]};
assign u1_col_in_487 = {col_in_487, u0_col_out_231, reg_intermediate0[231], reg_intermediate1[231]};
assign u1_col_in_488 = {col_in_488, u0_col_out_232, reg_intermediate0[232], reg_intermediate1[232]};
assign u1_col_in_489 = {col_in_489, u0_col_out_233, reg_intermediate0[233], reg_intermediate1[233]};
assign u1_col_in_490 = {col_in_490, u0_col_out_234, reg_intermediate0[234], reg_intermediate1[234]};
assign u1_col_in_491 = {col_in_491, u0_col_out_235, reg_intermediate0[235], reg_intermediate1[235]};
assign u1_col_in_492 = {col_in_492, u0_col_out_236, reg_intermediate0[236], reg_intermediate1[236]};
assign u1_col_in_493 = {col_in_493, u0_col_out_237, reg_intermediate0[237], reg_intermediate1[237]};
assign u1_col_in_494 = {col_in_494, u0_col_out_238, reg_intermediate0[238], reg_intermediate1[238]};
assign u1_col_in_495 = {col_in_495, u0_col_out_239, reg_intermediate0[239], reg_intermediate1[239]};
assign u1_col_in_496 = {col_in_496, u0_col_out_240, reg_intermediate0[240], reg_intermediate1[240]};
assign u1_col_in_497 = {col_in_497, u0_col_out_241, reg_intermediate0[241], reg_intermediate1[241]};
assign u1_col_in_498 = {col_in_498, u0_col_out_242, reg_intermediate0[242], reg_intermediate1[242]};
assign u1_col_in_499 = {col_in_499, u0_col_out_243, reg_intermediate0[243], reg_intermediate1[243]};
assign u1_col_in_500 = {col_in_500, u0_col_out_244, reg_intermediate0[244], reg_intermediate1[244]};
assign u1_col_in_501 = {col_in_501, u0_col_out_245, reg_intermediate0[245], reg_intermediate1[245]};
assign u1_col_in_502 = {col_in_502, u0_col_out_246, reg_intermediate0[246], reg_intermediate1[246]};
assign u1_col_in_503 = {col_in_503, u0_col_out_247, reg_intermediate0[247], reg_intermediate1[247]};
assign u1_col_in_504 = {col_in_504, u0_col_out_248, reg_intermediate0[248], reg_intermediate1[248]};
assign u1_col_in_505 = {col_in_505, u0_col_out_249, reg_intermediate0[249], reg_intermediate1[249]};
assign u1_col_in_506 = {col_in_506, u0_col_out_250, reg_intermediate0[250], reg_intermediate1[250]};
assign u1_col_in_507 = {col_in_507, u0_col_out_251, reg_intermediate0[251], reg_intermediate1[251]};
assign u1_col_in_508 = {col_in_508, u0_col_out_252, reg_intermediate0[252], reg_intermediate1[252]};
assign u1_col_in_509 = {col_in_509, u0_col_out_253, reg_intermediate0[253], reg_intermediate1[253]};
assign u1_col_in_510 = {col_in_510, u0_col_out_254, reg_intermediate0[254], reg_intermediate1[254]};
assign u1_col_in_511 = {col_in_511, u0_col_out_255, reg_intermediate0[255], reg_intermediate1[255]};
assign u1_col_in_512 = {col_in_512, u0_col_out_256, reg_intermediate0[256], reg_intermediate1[256]};
assign u1_col_in_513 = {col_in_513, u0_col_out_257, reg_intermediate0[257], reg_intermediate1[257]};
assign u1_col_in_514 = {col_in_514, u0_col_out_258, reg_intermediate0[258], reg_intermediate1[258]};
assign u1_col_in_515 = {col_in_515, u0_col_out_259, reg_intermediate0[259], reg_intermediate1[259]};
assign u1_col_in_516 = {col_in_516, u0_col_out_260, reg_intermediate0[260], reg_intermediate1[260]};
assign u1_col_in_517 = {col_in_517, u0_col_out_261, reg_intermediate0[261], reg_intermediate1[261]};
assign u1_col_in_518 = {col_in_518, u0_col_out_262, reg_intermediate0[262], reg_intermediate1[262]};
assign u1_col_in_519 = {col_in_519, u0_col_out_263, reg_intermediate0[263], reg_intermediate1[263]};
assign u1_col_in_520 = {col_in_520, u0_col_out_264, reg_intermediate0[264], reg_intermediate1[264]};
assign u1_col_in_521 = {col_in_521, u0_col_out_265, reg_intermediate0[265], reg_intermediate1[265]};
assign u1_col_in_522 = {col_in_522, u0_col_out_266, reg_intermediate0[266], reg_intermediate1[266]};
assign u1_col_in_523 = {col_in_523, u0_col_out_267, reg_intermediate0[267], reg_intermediate1[267]};
assign u1_col_in_524 = {col_in_524, u0_col_out_268, reg_intermediate0[268], reg_intermediate1[268]};
assign u1_col_in_525 = {col_in_525, u0_col_out_269, reg_intermediate0[269], reg_intermediate1[269]};
assign u1_col_in_526 = {col_in_526, u0_col_out_270, reg_intermediate0[270], reg_intermediate1[270]};
assign u1_col_in_527 = {col_in_527, u0_col_out_271, reg_intermediate0[271], reg_intermediate1[271]};
assign u1_col_in_528 = {col_in_528, u0_col_out_272, reg_intermediate0[272], reg_intermediate1[272]};
assign u1_col_in_529 = {col_in_529, u0_col_out_273, reg_intermediate0[273], reg_intermediate1[273]};
assign u1_col_in_530 = {col_in_530, u0_col_out_274, reg_intermediate0[274], reg_intermediate1[274]};
assign u1_col_in_531 = {col_in_531, u0_col_out_275, reg_intermediate0[275], reg_intermediate1[275]};
assign u1_col_in_532 = {col_in_532, u0_col_out_276, reg_intermediate0[276], reg_intermediate1[276]};
assign u1_col_in_533 = {col_in_533, u0_col_out_277, reg_intermediate0[277], reg_intermediate1[277]};
assign u1_col_in_534 = {col_in_534, u0_col_out_278, reg_intermediate0[278], reg_intermediate1[278]};
assign u1_col_in_535 = {col_in_535, u0_col_out_279, reg_intermediate0[279], reg_intermediate1[279]};
assign u1_col_in_536 = {col_in_536, u0_col_out_280, reg_intermediate0[280], reg_intermediate1[280]};
assign u1_col_in_537 = {col_in_537, u0_col_out_281, reg_intermediate0[281], reg_intermediate1[281]};
assign u1_col_in_538 = {col_in_538, u0_col_out_282, reg_intermediate0[282], reg_intermediate1[282]};
assign u1_col_in_539 = {col_in_539, u0_col_out_283, reg_intermediate0[283], reg_intermediate1[283]};
assign u1_col_in_540 = {col_in_540, u0_col_out_284, reg_intermediate0[284], reg_intermediate1[284]};
assign u1_col_in_541 = {col_in_541, u0_col_out_285, reg_intermediate0[285], reg_intermediate1[285]};
assign u1_col_in_542 = {col_in_542, u0_col_out_286, reg_intermediate0[286], reg_intermediate1[286]};
assign u1_col_in_543 = {col_in_543, u0_col_out_287, reg_intermediate0[287], reg_intermediate1[287]};
assign u1_col_in_544 = {col_in_544, u0_col_out_288, reg_intermediate0[288], reg_intermediate1[288]};
assign u1_col_in_545 = {col_in_545, u0_col_out_289, reg_intermediate0[289], reg_intermediate1[289]};
assign u1_col_in_546 = {col_in_546, u0_col_out_290, reg_intermediate0[290], reg_intermediate1[290]};
assign u1_col_in_547 = {col_in_547, u0_col_out_291, reg_intermediate0[291], reg_intermediate1[291]};
assign u1_col_in_548 = {col_in_548, u0_col_out_292, reg_intermediate0[292], reg_intermediate1[292]};
assign u1_col_in_549 = {col_in_549, u0_col_out_293, reg_intermediate0[293], reg_intermediate1[293]};
assign u1_col_in_550 = {col_in_550, u0_col_out_294, reg_intermediate0[294], reg_intermediate1[294]};
assign u1_col_in_551 = {col_in_551, u0_col_out_295, reg_intermediate0[295], reg_intermediate1[295]};
assign u1_col_in_552 = {col_in_552, u0_col_out_296, reg_intermediate0[296], reg_intermediate1[296]};
assign u1_col_in_553 = {col_in_553, u0_col_out_297, reg_intermediate0[297], reg_intermediate1[297]};
assign u1_col_in_554 = {col_in_554, u0_col_out_298, reg_intermediate0[298], reg_intermediate1[298]};
assign u1_col_in_555 = {col_in_555, u0_col_out_299, reg_intermediate0[299], reg_intermediate1[299]};
assign u1_col_in_556 = {col_in_556, u0_col_out_300, reg_intermediate0[300], reg_intermediate1[300]};
assign u1_col_in_557 = {col_in_557, u0_col_out_301, reg_intermediate0[301], reg_intermediate1[301]};
assign u1_col_in_558 = {col_in_558, u0_col_out_302, reg_intermediate0[302], reg_intermediate1[302]};
assign u1_col_in_559 = {col_in_559, u0_col_out_303, reg_intermediate0[303], reg_intermediate1[303]};
assign u1_col_in_560 = {col_in_560, u0_col_out_304, reg_intermediate0[304], reg_intermediate1[304]};
assign u1_col_in_561 = {col_in_561, u0_col_out_305, reg_intermediate0[305], reg_intermediate1[305]};
assign u1_col_in_562 = {col_in_562, u0_col_out_306, reg_intermediate0[306], reg_intermediate1[306]};
assign u1_col_in_563 = {col_in_563, u0_col_out_307, reg_intermediate0[307], reg_intermediate1[307]};
assign u1_col_in_564 = {col_in_564, u0_col_out_308, reg_intermediate0[308], reg_intermediate1[308]};
assign u1_col_in_565 = {col_in_565, u0_col_out_309, reg_intermediate0[309], reg_intermediate1[309]};
assign u1_col_in_566 = {col_in_566, u0_col_out_310, reg_intermediate0[310], reg_intermediate1[310]};
assign u1_col_in_567 = {col_in_567, u0_col_out_311, reg_intermediate0[311], reg_intermediate1[311]};
assign u1_col_in_568 = {col_in_568, u0_col_out_312, reg_intermediate0[312], reg_intermediate1[312]};
assign u1_col_in_569 = {col_in_569, u0_col_out_313, reg_intermediate0[313], reg_intermediate1[313]};
assign u1_col_in_570 = {col_in_570, u0_col_out_314, reg_intermediate0[314], reg_intermediate1[314]};
assign u1_col_in_571 = {col_in_571, u0_col_out_315, reg_intermediate0[315], reg_intermediate1[315]};
assign u1_col_in_572 = {col_in_572, u0_col_out_316, reg_intermediate0[316], reg_intermediate1[316]};
assign u1_col_in_573 = {col_in_573, u0_col_out_317, reg_intermediate0[317], reg_intermediate1[317]};
assign u1_col_in_574 = {col_in_574, u0_col_out_318, reg_intermediate0[318], reg_intermediate1[318]};
assign u1_col_in_575 = {col_in_575, u0_col_out_319, reg_intermediate0[319], reg_intermediate1[319]};
assign u1_col_in_576 = {col_in_576, u0_col_out_320, reg_intermediate0[320], reg_intermediate1[320]};
assign u1_col_in_577 = {col_in_577, u0_col_out_321, reg_intermediate0[321], reg_intermediate1[321]};
assign u1_col_in_578 = {col_in_578, u0_col_out_322, reg_intermediate0[322], reg_intermediate1[322]};
assign u1_col_in_579 = {col_in_579, u0_col_out_323, reg_intermediate0[323], reg_intermediate1[323]};
assign u1_col_in_580 = {col_in_580, u0_col_out_324, reg_intermediate0[324], reg_intermediate1[324]};
assign u1_col_in_581 = {col_in_581, u0_col_out_325, reg_intermediate0[325], reg_intermediate1[325]};
assign u1_col_in_582 = {col_in_582, u0_col_out_326, reg_intermediate0[326], reg_intermediate1[326]};
assign u1_col_in_583 = {col_in_583, u0_col_out_327, reg_intermediate0[327], reg_intermediate1[327]};
assign u1_col_in_584 = {col_in_584, u0_col_out_328, reg_intermediate0[328], reg_intermediate1[328]};
assign u1_col_in_585 = {col_in_585, u0_col_out_329, reg_intermediate0[329], reg_intermediate1[329]};
assign u1_col_in_586 = {col_in_586, u0_col_out_330, reg_intermediate0[330], reg_intermediate1[330]};
assign u1_col_in_587 = {col_in_587, u0_col_out_331, reg_intermediate0[331], reg_intermediate1[331]};
assign u1_col_in_588 = {col_in_588, u0_col_out_332, reg_intermediate0[332], reg_intermediate1[332]};
assign u1_col_in_589 = {col_in_589, u0_col_out_333, reg_intermediate0[333], reg_intermediate1[333]};
assign u1_col_in_590 = {col_in_590, u0_col_out_334, reg_intermediate0[334], reg_intermediate1[334]};
assign u1_col_in_591 = {col_in_591, u0_col_out_335, reg_intermediate0[335], reg_intermediate1[335]};
assign u1_col_in_592 = {col_in_592, u0_col_out_336, reg_intermediate0[336], reg_intermediate1[336]};
assign u1_col_in_593 = {col_in_593, u0_col_out_337, reg_intermediate0[337], reg_intermediate1[337]};
assign u1_col_in_594 = {col_in_594, u0_col_out_338, reg_intermediate0[338], reg_intermediate1[338]};
assign u1_col_in_595 = {col_in_595, u0_col_out_339, reg_intermediate0[339], reg_intermediate1[339]};
assign u1_col_in_596 = {col_in_596, u0_col_out_340, reg_intermediate0[340], reg_intermediate1[340]};
assign u1_col_in_597 = {col_in_597, u0_col_out_341, reg_intermediate0[341], reg_intermediate1[341]};
assign u1_col_in_598 = {col_in_598, u0_col_out_342, reg_intermediate0[342], reg_intermediate1[342]};
assign u1_col_in_599 = {col_in_599, u0_col_out_343, reg_intermediate0[343], reg_intermediate1[343]};
assign u1_col_in_600 = {col_in_600, u0_col_out_344, reg_intermediate0[344], reg_intermediate1[344]};
assign u1_col_in_601 = {col_in_601, u0_col_out_345, reg_intermediate0[345], reg_intermediate1[345]};
assign u1_col_in_602 = {col_in_602, u0_col_out_346, reg_intermediate0[346], reg_intermediate1[346]};
assign u1_col_in_603 = {col_in_603, u0_col_out_347, reg_intermediate0[347], reg_intermediate1[347]};
assign u1_col_in_604 = {col_in_604, u0_col_out_348, reg_intermediate0[348], reg_intermediate1[348]};
assign u1_col_in_605 = {col_in_605, u0_col_out_349, reg_intermediate0[349], reg_intermediate1[349]};
assign u1_col_in_606 = {col_in_606, u0_col_out_350, reg_intermediate0[350], reg_intermediate1[350]};
assign u1_col_in_607 = {col_in_607, u0_col_out_351, reg_intermediate0[351], reg_intermediate1[351]};
assign u1_col_in_608 = {col_in_608, u0_col_out_352, reg_intermediate0[352], reg_intermediate1[352]};
assign u1_col_in_609 = {col_in_609, u0_col_out_353, reg_intermediate0[353], reg_intermediate1[353]};
assign u1_col_in_610 = {col_in_610, u0_col_out_354, reg_intermediate0[354], reg_intermediate1[354]};
assign u1_col_in_611 = {col_in_611, u0_col_out_355, reg_intermediate0[355], reg_intermediate1[355]};
assign u1_col_in_612 = {col_in_612, u0_col_out_356, reg_intermediate0[356], reg_intermediate1[356]};
assign u1_col_in_613 = {col_in_613, u0_col_out_357, reg_intermediate0[357], reg_intermediate1[357]};
assign u1_col_in_614 = {col_in_614, u0_col_out_358, reg_intermediate0[358], reg_intermediate1[358]};
assign u1_col_in_615 = {col_in_615, u0_col_out_359, reg_intermediate0[359], reg_intermediate1[359]};
assign u1_col_in_616 = {col_in_616, u0_col_out_360, reg_intermediate0[360], reg_intermediate1[360]};
assign u1_col_in_617 = {col_in_617, u0_col_out_361, reg_intermediate0[361], reg_intermediate1[361]};
assign u1_col_in_618 = {col_in_618, u0_col_out_362, reg_intermediate0[362], reg_intermediate1[362]};
assign u1_col_in_619 = {col_in_619, u0_col_out_363, reg_intermediate0[363], reg_intermediate1[363]};
assign u1_col_in_620 = {col_in_620, u0_col_out_364, reg_intermediate0[364], reg_intermediate1[364]};
assign u1_col_in_621 = {col_in_621, u0_col_out_365, reg_intermediate0[365], reg_intermediate1[365]};
assign u1_col_in_622 = {col_in_622, u0_col_out_366, reg_intermediate0[366], reg_intermediate1[366]};
assign u1_col_in_623 = {col_in_623, u0_col_out_367, reg_intermediate0[367], reg_intermediate1[367]};
assign u1_col_in_624 = {col_in_624, u0_col_out_368, reg_intermediate0[368], reg_intermediate1[368]};
assign u1_col_in_625 = {col_in_625, u0_col_out_369, reg_intermediate0[369], reg_intermediate1[369]};
assign u1_col_in_626 = {col_in_626, u0_col_out_370, reg_intermediate0[370], reg_intermediate1[370]};
assign u1_col_in_627 = {col_in_627, u0_col_out_371, reg_intermediate0[371], reg_intermediate1[371]};
assign u1_col_in_628 = {col_in_628, u0_col_out_372, reg_intermediate0[372], reg_intermediate1[372]};
assign u1_col_in_629 = {col_in_629, u0_col_out_373, reg_intermediate0[373], reg_intermediate1[373]};
assign u1_col_in_630 = {col_in_630, u0_col_out_374, reg_intermediate0[374], reg_intermediate1[374]};
assign u1_col_in_631 = {col_in_631, u0_col_out_375, reg_intermediate0[375], reg_intermediate1[375]};
assign u1_col_in_632 = {col_in_632, u0_col_out_376, reg_intermediate0[376], reg_intermediate1[376]};
assign u1_col_in_633 = {col_in_633, u0_col_out_377, reg_intermediate0[377], reg_intermediate1[377]};
assign u1_col_in_634 = {col_in_634, u0_col_out_378, reg_intermediate0[378], reg_intermediate1[378]};
assign u1_col_in_635 = {col_in_635, u0_col_out_379, reg_intermediate0[379], reg_intermediate1[379]};
assign u1_col_in_636 = {col_in_636, u0_col_out_380, reg_intermediate0[380], reg_intermediate1[380]};
assign u1_col_in_637 = {col_in_637, u0_col_out_381, reg_intermediate0[381], reg_intermediate1[381]};
assign u1_col_in_638 = {col_in_638, u0_col_out_382, reg_intermediate0[382], reg_intermediate1[382]};
assign u1_col_in_639 = {col_in_639, u0_col_out_383, reg_intermediate0[383], reg_intermediate1[383]};
assign u1_col_in_640 = {col_in_640, u0_col_out_384, reg_intermediate0[384], reg_intermediate1[384]};
assign u1_col_in_641 = {col_in_641, u0_col_out_385, reg_intermediate0[385], reg_intermediate1[385]};
assign u1_col_in_642 = {col_in_642, u0_col_out_386, reg_intermediate0[386], reg_intermediate1[386]};
assign u1_col_in_643 = {col_in_643, u0_col_out_387, reg_intermediate0[387], reg_intermediate1[387]};
assign u1_col_in_644 = {col_in_644, u0_col_out_388, reg_intermediate0[388], reg_intermediate1[388]};
assign u1_col_in_645 = {col_in_645, u0_col_out_389, reg_intermediate0[389], reg_intermediate1[389]};
assign u1_col_in_646 = {col_in_646, u0_col_out_390, reg_intermediate0[390], reg_intermediate1[390]};
assign u1_col_in_647 = {col_in_647, u0_col_out_391, reg_intermediate0[391], reg_intermediate1[391]};
assign u1_col_in_648 = {col_in_648, u0_col_out_392, reg_intermediate0[392], reg_intermediate1[392]};
assign u1_col_in_649 = {col_in_649, u0_col_out_393, reg_intermediate0[393], reg_intermediate1[393]};
assign u1_col_in_650 = {col_in_650, u0_col_out_394, reg_intermediate0[394], reg_intermediate1[394]};
assign u1_col_in_651 = {col_in_651, u0_col_out_395, reg_intermediate0[395], reg_intermediate1[395]};
assign u1_col_in_652 = {col_in_652, u0_col_out_396, reg_intermediate0[396], reg_intermediate1[396]};
assign u1_col_in_653 = {col_in_653, u0_col_out_397, reg_intermediate0[397], reg_intermediate1[397]};
assign u1_col_in_654 = {col_in_654, u0_col_out_398, reg_intermediate0[398], reg_intermediate1[398]};
assign u1_col_in_655 = {col_in_655, u0_col_out_399, reg_intermediate0[399], reg_intermediate1[399]};
assign u1_col_in_656 = {col_in_656, u0_col_out_400, reg_intermediate0[400], reg_intermediate1[400]};
assign u1_col_in_657 = {col_in_657, u0_col_out_401, reg_intermediate0[401], reg_intermediate1[401]};
assign u1_col_in_658 = {col_in_658, u0_col_out_402, reg_intermediate0[402], reg_intermediate1[402]};
assign u1_col_in_659 = {col_in_659, u0_col_out_403, reg_intermediate0[403], reg_intermediate1[403]};
assign u1_col_in_660 = {col_in_660, u0_col_out_404, reg_intermediate0[404], reg_intermediate1[404]};
assign u1_col_in_661 = {col_in_661, u0_col_out_405, reg_intermediate0[405], reg_intermediate1[405]};
assign u1_col_in_662 = {col_in_662, u0_col_out_406, reg_intermediate0[406], reg_intermediate1[406]};
assign u1_col_in_663 = {col_in_663, u0_col_out_407, reg_intermediate0[407], reg_intermediate1[407]};
assign u1_col_in_664 = {col_in_664, u0_col_out_408, reg_intermediate0[408], reg_intermediate1[408]};
assign u1_col_in_665 = {col_in_665, u0_col_out_409, reg_intermediate0[409], reg_intermediate1[409]};
assign u1_col_in_666 = {col_in_666, u0_col_out_410, reg_intermediate0[410], reg_intermediate1[410]};
assign u1_col_in_667 = {col_in_667, u0_col_out_411, reg_intermediate0[411], reg_intermediate1[411]};
assign u1_col_in_668 = {col_in_668, u0_col_out_412, reg_intermediate0[412], reg_intermediate1[412]};
assign u1_col_in_669 = {col_in_669, u0_col_out_413, reg_intermediate0[413], reg_intermediate1[413]};
assign u1_col_in_670 = {col_in_670, u0_col_out_414, reg_intermediate0[414], reg_intermediate1[414]};
assign u1_col_in_671 = {col_in_671, u0_col_out_415, reg_intermediate0[415], reg_intermediate1[415]};
assign u1_col_in_672 = {col_in_672, u0_col_out_416, reg_intermediate0[416], reg_intermediate1[416]};
assign u1_col_in_673 = {col_in_673, u0_col_out_417, reg_intermediate0[417], reg_intermediate1[417]};
assign u1_col_in_674 = {col_in_674, u0_col_out_418, reg_intermediate0[418], reg_intermediate1[418]};
assign u1_col_in_675 = {col_in_675, u0_col_out_419, reg_intermediate0[419], reg_intermediate1[419]};
assign u1_col_in_676 = {col_in_676, u0_col_out_420, reg_intermediate0[420], reg_intermediate1[420]};
assign u1_col_in_677 = {col_in_677, u0_col_out_421, reg_intermediate0[421], reg_intermediate1[421]};
assign u1_col_in_678 = {col_in_678, u0_col_out_422, reg_intermediate0[422], reg_intermediate1[422]};
assign u1_col_in_679 = {col_in_679, u0_col_out_423, reg_intermediate0[423], reg_intermediate1[423]};
assign u1_col_in_680 = {col_in_680, u0_col_out_424, reg_intermediate0[424], reg_intermediate1[424]};
assign u1_col_in_681 = {col_in_681, u0_col_out_425, reg_intermediate0[425], reg_intermediate1[425]};
assign u1_col_in_682 = {col_in_682, u0_col_out_426, reg_intermediate0[426], reg_intermediate1[426]};
assign u1_col_in_683 = {col_in_683, u0_col_out_427, reg_intermediate0[427], reg_intermediate1[427]};
assign u1_col_in_684 = {col_in_684, u0_col_out_428, reg_intermediate0[428], reg_intermediate1[428]};
assign u1_col_in_685 = {col_in_685, u0_col_out_429, reg_intermediate0[429], reg_intermediate1[429]};
assign u1_col_in_686 = {col_in_686, u0_col_out_430, reg_intermediate0[430], reg_intermediate1[430]};
assign u1_col_in_687 = {col_in_687, u0_col_out_431, reg_intermediate0[431], reg_intermediate1[431]};
assign u1_col_in_688 = {col_in_688, u0_col_out_432, reg_intermediate0[432], reg_intermediate1[432]};
assign u1_col_in_689 = {col_in_689, u0_col_out_433, reg_intermediate0[433], reg_intermediate1[433]};
assign u1_col_in_690 = {col_in_690, u0_col_out_434, reg_intermediate0[434], reg_intermediate1[434]};
assign u1_col_in_691 = {col_in_691, u0_col_out_435, reg_intermediate0[435], reg_intermediate1[435]};
assign u1_col_in_692 = {col_in_692, u0_col_out_436, reg_intermediate0[436], reg_intermediate1[436]};
assign u1_col_in_693 = {col_in_693, u0_col_out_437, reg_intermediate0[437], reg_intermediate1[437]};
assign u1_col_in_694 = {col_in_694, u0_col_out_438, reg_intermediate0[438], reg_intermediate1[438]};
assign u1_col_in_695 = {col_in_695, u0_col_out_439, reg_intermediate0[439], reg_intermediate1[439]};
assign u1_col_in_696 = {col_in_696, u0_col_out_440, reg_intermediate0[440], reg_intermediate1[440]};
assign u1_col_in_697 = {col_in_697, u0_col_out_441, reg_intermediate0[441], reg_intermediate1[441]};
assign u1_col_in_698 = {col_in_698, u0_col_out_442, reg_intermediate0[442], reg_intermediate1[442]};
assign u1_col_in_699 = {col_in_699, u0_col_out_443, reg_intermediate0[443], reg_intermediate1[443]};
assign u1_col_in_700 = {col_in_700, u0_col_out_444, reg_intermediate0[444], reg_intermediate1[444]};
assign u1_col_in_701 = {col_in_701, u0_col_out_445, reg_intermediate0[445], reg_intermediate1[445]};
assign u1_col_in_702 = {col_in_702, u0_col_out_446, reg_intermediate0[446], reg_intermediate1[446]};
assign u1_col_in_703 = {col_in_703, u0_col_out_447, reg_intermediate0[447], reg_intermediate1[447]};
assign u1_col_in_704 = {col_in_704, u0_col_out_448, reg_intermediate0[448], reg_intermediate1[448]};
assign u1_col_in_705 = {col_in_705, u0_col_out_449, reg_intermediate0[449], reg_intermediate1[449]};
assign u1_col_in_706 = {col_in_706, u0_col_out_450, reg_intermediate0[450], reg_intermediate1[450]};
assign u1_col_in_707 = {col_in_707, u0_col_out_451, reg_intermediate0[451], reg_intermediate1[451]};
assign u1_col_in_708 = {col_in_708, u0_col_out_452, reg_intermediate0[452], reg_intermediate1[452]};
assign u1_col_in_709 = {col_in_709, u0_col_out_453, reg_intermediate0[453], reg_intermediate1[453]};
assign u1_col_in_710 = {col_in_710, u0_col_out_454, reg_intermediate0[454], reg_intermediate1[454]};
assign u1_col_in_711 = {col_in_711, u0_col_out_455, reg_intermediate0[455], reg_intermediate1[455]};
assign u1_col_in_712 = {col_in_712, u0_col_out_456, reg_intermediate0[456], reg_intermediate1[456]};
assign u1_col_in_713 = {col_in_713, u0_col_out_457, reg_intermediate0[457], reg_intermediate1[457]};
assign u1_col_in_714 = {col_in_714, u0_col_out_458, reg_intermediate0[458], reg_intermediate1[458]};
assign u1_col_in_715 = {col_in_715, u0_col_out_459, reg_intermediate0[459], reg_intermediate1[459]};
assign u1_col_in_716 = {col_in_716, u0_col_out_460, reg_intermediate0[460], reg_intermediate1[460]};
assign u1_col_in_717 = {col_in_717, u0_col_out_461, reg_intermediate0[461], reg_intermediate1[461]};
assign u1_col_in_718 = {col_in_718, u0_col_out_462, reg_intermediate0[462], reg_intermediate1[462]};
assign u1_col_in_719 = {col_in_719, u0_col_out_463, reg_intermediate0[463], reg_intermediate1[463]};
assign u1_col_in_720 = {col_in_720, u0_col_out_464, reg_intermediate0[464], reg_intermediate1[464]};
assign u1_col_in_721 = {col_in_721, u0_col_out_465, reg_intermediate0[465], reg_intermediate1[465]};
assign u1_col_in_722 = {col_in_722, u0_col_out_466, reg_intermediate0[466], reg_intermediate1[466]};
assign u1_col_in_723 = {col_in_723, u0_col_out_467, reg_intermediate0[467], reg_intermediate1[467]};
assign u1_col_in_724 = {col_in_724, u0_col_out_468, reg_intermediate0[468], reg_intermediate1[468]};
assign u1_col_in_725 = {col_in_725, u0_col_out_469, reg_intermediate0[469], reg_intermediate1[469]};
assign u1_col_in_726 = {col_in_726, u0_col_out_470, reg_intermediate0[470], reg_intermediate1[470]};
assign u1_col_in_727 = {col_in_727, u0_col_out_471, reg_intermediate0[471], reg_intermediate1[471]};
assign u1_col_in_728 = {col_in_728, u0_col_out_472, reg_intermediate0[472], reg_intermediate1[472]};
assign u1_col_in_729 = {col_in_729, u0_col_out_473, reg_intermediate0[473], reg_intermediate1[473]};
assign u1_col_in_730 = {col_in_730, u0_col_out_474, reg_intermediate0[474], reg_intermediate1[474]};
assign u1_col_in_731 = {col_in_731, u0_col_out_475, reg_intermediate0[475], reg_intermediate1[475]};
assign u1_col_in_732 = {col_in_732, u0_col_out_476, reg_intermediate0[476], reg_intermediate1[476]};
assign u1_col_in_733 = {col_in_733, u0_col_out_477, reg_intermediate0[477], reg_intermediate1[477]};
assign u1_col_in_734 = {col_in_734, u0_col_out_478, reg_intermediate0[478], reg_intermediate1[478]};
assign u1_col_in_735 = {col_in_735, u0_col_out_479, reg_intermediate0[479], reg_intermediate1[479]};
assign u1_col_in_736 = {col_in_736, u0_col_out_480, reg_intermediate0[480], reg_intermediate1[480]};
assign u1_col_in_737 = {col_in_737, u0_col_out_481, reg_intermediate0[481], reg_intermediate1[481]};
assign u1_col_in_738 = {col_in_738, u0_col_out_482, reg_intermediate0[482], reg_intermediate1[482]};
assign u1_col_in_739 = {col_in_739, u0_col_out_483, reg_intermediate0[483], reg_intermediate1[483]};
assign u1_col_in_740 = {col_in_740, u0_col_out_484, reg_intermediate0[484], reg_intermediate1[484]};
assign u1_col_in_741 = {col_in_741, u0_col_out_485, reg_intermediate0[485], reg_intermediate1[485]};
assign u1_col_in_742 = {col_in_742, u0_col_out_486, reg_intermediate0[486], reg_intermediate1[486]};
assign u1_col_in_743 = {col_in_743, u0_col_out_487, reg_intermediate0[487], reg_intermediate1[487]};
assign u1_col_in_744 = {col_in_744, u0_col_out_488, reg_intermediate0[488], reg_intermediate1[488]};
assign u1_col_in_745 = {col_in_745, u0_col_out_489, reg_intermediate0[489], reg_intermediate1[489]};
assign u1_col_in_746 = {col_in_746, u0_col_out_490, reg_intermediate0[490], reg_intermediate1[490]};
assign u1_col_in_747 = {col_in_747, u0_col_out_491, reg_intermediate0[491], reg_intermediate1[491]};
assign u1_col_in_748 = {col_in_748, u0_col_out_492, reg_intermediate0[492], reg_intermediate1[492]};
assign u1_col_in_749 = {col_in_749, u0_col_out_493, reg_intermediate0[493], reg_intermediate1[493]};
assign u1_col_in_750 = {col_in_750, u0_col_out_494, reg_intermediate0[494], reg_intermediate1[494]};
assign u1_col_in_751 = {col_in_751, u0_col_out_495, reg_intermediate0[495], reg_intermediate1[495]};
assign u1_col_in_752 = {col_in_752, u0_col_out_496, reg_intermediate0[496], reg_intermediate1[496]};
assign u1_col_in_753 = {col_in_753, u0_col_out_497, reg_intermediate0[497], reg_intermediate1[497]};
assign u1_col_in_754 = {col_in_754, u0_col_out_498, reg_intermediate0[498], reg_intermediate1[498]};
assign u1_col_in_755 = {col_in_755, u0_col_out_499, reg_intermediate0[499], reg_intermediate1[499]};
assign u1_col_in_756 = {col_in_756, u0_col_out_500, reg_intermediate0[500], reg_intermediate1[500]};
assign u1_col_in_757 = {col_in_757, u0_col_out_501, reg_intermediate0[501], reg_intermediate1[501]};
assign u1_col_in_758 = {col_in_758, u0_col_out_502, reg_intermediate0[502], reg_intermediate1[502]};
assign u1_col_in_759 = {col_in_759, u0_col_out_503, reg_intermediate0[503], reg_intermediate1[503]};
assign u1_col_in_760 = {col_in_760, u0_col_out_504, reg_intermediate0[504], reg_intermediate1[504]};
assign u1_col_in_761 = {col_in_761, u0_col_out_505, reg_intermediate0[505], reg_intermediate1[505]};
assign u1_col_in_762 = {col_in_762, u0_col_out_506, reg_intermediate0[506], reg_intermediate1[506]};
assign u1_col_in_763 = {col_in_763, u0_col_out_507, reg_intermediate0[507], reg_intermediate1[507]};
assign u1_col_in_764 = {col_in_764, u0_col_out_508, reg_intermediate0[508], reg_intermediate1[508]};
assign u1_col_in_765 = {col_in_765, u0_col_out_509, reg_intermediate0[509], reg_intermediate1[509]};
assign u1_col_in_766 = {col_in_766, u0_col_out_510, reg_intermediate0[510], reg_intermediate1[510]};
assign u1_col_in_767 = {col_in_767, u0_col_out_511, reg_intermediate0[511], reg_intermediate1[511]};
assign u1_col_in_768 = {col_in_768, u0_col_out_512, reg_intermediate0[512], reg_intermediate1[512]};
assign u1_col_in_769 = {col_in_769, u0_col_out_513, reg_intermediate0[513], reg_intermediate1[513]};
assign u1_col_in_770 = {col_in_770, u0_col_out_514, reg_intermediate0[514], reg_intermediate1[514]};
assign u1_col_in_771 = {col_in_771, u0_col_out_515, reg_intermediate0[515], reg_intermediate1[515]};
assign u1_col_in_772 = {col_in_772, u0_col_out_516, reg_intermediate0[516], reg_intermediate1[516]};
assign u1_col_in_773 = {col_in_773, u0_col_out_517, reg_intermediate0[517], reg_intermediate1[517]};
assign u1_col_in_774 = {col_in_774, u0_col_out_518, reg_intermediate0[518], reg_intermediate1[518]};
assign u1_col_in_775 = {col_in_775, u0_col_out_519, reg_intermediate0[519], reg_intermediate1[519]};
assign u1_col_in_776 = {col_in_776, u0_col_out_520, reg_intermediate0[520], reg_intermediate1[520]};
assign u1_col_in_777 = {col_in_777, u0_col_out_521, reg_intermediate0[521], reg_intermediate1[521]};
assign u1_col_in_778 = {col_in_778, u0_col_out_522, reg_intermediate0[522], reg_intermediate1[522]};
assign u1_col_in_779 = {col_in_779, u0_col_out_523, reg_intermediate0[523], reg_intermediate1[523]};
assign u1_col_in_780 = {col_in_780, u0_col_out_524, reg_intermediate0[524], reg_intermediate1[524]};
assign u1_col_in_781 = {col_in_781, u0_col_out_525, reg_intermediate0[525], reg_intermediate1[525]};
assign u1_col_in_782 = {col_in_782, u0_col_out_526, reg_intermediate0[526], reg_intermediate1[526]};
assign u1_col_in_783 = {col_in_783, u0_col_out_527, reg_intermediate0[527], reg_intermediate1[527]};
assign u1_col_in_784 = {col_in_784, u0_col_out_528, reg_intermediate0[528], reg_intermediate1[528]};
assign u1_col_in_785 = {col_in_785, u0_col_out_529, reg_intermediate0[529], reg_intermediate1[529]};
assign u1_col_in_786 = {col_in_786, u0_col_out_530, reg_intermediate0[530], reg_intermediate1[530]};
assign u1_col_in_787 = {col_in_787, u0_col_out_531, reg_intermediate0[531], reg_intermediate1[531]};
assign u1_col_in_788 = {col_in_788, u0_col_out_532, reg_intermediate0[532], reg_intermediate1[532]};
assign u1_col_in_789 = {col_in_789, u0_col_out_533, reg_intermediate0[533], reg_intermediate1[533]};
assign u1_col_in_790 = {col_in_790, u0_col_out_534, reg_intermediate0[534], reg_intermediate1[534]};
assign u1_col_in_791 = {col_in_791, u0_col_out_535, reg_intermediate0[535], reg_intermediate1[535]};
assign u1_col_in_792 = {col_in_792, u0_col_out_536, reg_intermediate0[536], reg_intermediate1[536]};
assign u1_col_in_793 = {col_in_793, u0_col_out_537, reg_intermediate0[537], reg_intermediate1[537]};
assign u1_col_in_794 = {col_in_794, u0_col_out_538, reg_intermediate0[538], reg_intermediate1[538]};
assign u1_col_in_795 = {col_in_795, u0_col_out_539, reg_intermediate0[539], reg_intermediate1[539]};
assign u1_col_in_796 = {col_in_796, u0_col_out_540, reg_intermediate0[540], reg_intermediate1[540]};
assign u1_col_in_797 = {col_in_797, u0_col_out_541, reg_intermediate0[541], reg_intermediate1[541]};
assign u1_col_in_798 = {col_in_798, u0_col_out_542, reg_intermediate0[542], reg_intermediate1[542]};
assign u1_col_in_799 = {col_in_799, u0_col_out_543, reg_intermediate0[543], reg_intermediate1[543]};
assign u1_col_in_800 = {col_in_800, u0_col_out_544, reg_intermediate0[544], reg_intermediate1[544]};
assign u1_col_in_801 = {col_in_801, u0_col_out_545, reg_intermediate0[545], reg_intermediate1[545]};
assign u1_col_in_802 = {col_in_802, u0_col_out_546, reg_intermediate0[546], reg_intermediate1[546]};
assign u1_col_in_803 = {col_in_803, u0_col_out_547, reg_intermediate0[547], reg_intermediate1[547]};
assign u1_col_in_804 = {col_in_804, u0_col_out_548, reg_intermediate0[548], reg_intermediate1[548]};
assign u1_col_in_805 = {col_in_805, u0_col_out_549, reg_intermediate0[549], reg_intermediate1[549]};
assign u1_col_in_806 = {col_in_806, u0_col_out_550, reg_intermediate0[550], reg_intermediate1[550]};
assign u1_col_in_807 = {col_in_807, u0_col_out_551, reg_intermediate0[551], reg_intermediate1[551]};
assign u1_col_in_808 = {col_in_808, u0_col_out_552, reg_intermediate0[552], reg_intermediate1[552]};
assign u1_col_in_809 = {col_in_809, u0_col_out_553, reg_intermediate0[553], reg_intermediate1[553]};
assign u1_col_in_810 = {col_in_810, u0_col_out_554, reg_intermediate0[554], reg_intermediate1[554]};
assign u1_col_in_811 = {col_in_811, u0_col_out_555, reg_intermediate0[555], reg_intermediate1[555]};
assign u1_col_in_812 = {col_in_812, u0_col_out_556, reg_intermediate0[556], reg_intermediate1[556]};
assign u1_col_in_813 = {col_in_813, u0_col_out_557, reg_intermediate0[557], reg_intermediate1[557]};
assign u1_col_in_814 = {col_in_814, u0_col_out_558, reg_intermediate0[558], reg_intermediate1[558]};
assign u1_col_in_815 = {col_in_815, u0_col_out_559, reg_intermediate0[559], reg_intermediate1[559]};
assign u1_col_in_816 = {col_in_816, u0_col_out_560, reg_intermediate0[560], reg_intermediate1[560]};
assign u1_col_in_817 = {col_in_817, u0_col_out_561, reg_intermediate0[561], reg_intermediate1[561]};
assign u1_col_in_818 = {col_in_818, u0_col_out_562, reg_intermediate0[562], reg_intermediate1[562]};
assign u1_col_in_819 = {col_in_819, u0_col_out_563, reg_intermediate0[563], reg_intermediate1[563]};
assign u1_col_in_820 = {col_in_820, u0_col_out_564, reg_intermediate0[564], reg_intermediate1[564]};
assign u1_col_in_821 = {col_in_821, u0_col_out_565, reg_intermediate0[565], reg_intermediate1[565]};
assign u1_col_in_822 = {col_in_822, u0_col_out_566, reg_intermediate0[566], reg_intermediate1[566]};
assign u1_col_in_823 = {col_in_823, u0_col_out_567, reg_intermediate0[567], reg_intermediate1[567]};
assign u1_col_in_824 = {col_in_824, u0_col_out_568, reg_intermediate0[568], reg_intermediate1[568]};
assign u1_col_in_825 = {col_in_825, u0_col_out_569, reg_intermediate0[569], reg_intermediate1[569]};
assign u1_col_in_826 = {col_in_826, u0_col_out_570, reg_intermediate0[570], reg_intermediate1[570]};
assign u1_col_in_827 = {col_in_827, u0_col_out_571, reg_intermediate0[571], reg_intermediate1[571]};
assign u1_col_in_828 = {col_in_828, u0_col_out_572, reg_intermediate0[572], reg_intermediate1[572]};
assign u1_col_in_829 = {col_in_829, u0_col_out_573, reg_intermediate0[573], reg_intermediate1[573]};
assign u1_col_in_830 = {col_in_830, u0_col_out_574, reg_intermediate0[574], reg_intermediate1[574]};
assign u1_col_in_831 = {col_in_831, u0_col_out_575, reg_intermediate0[575], reg_intermediate1[575]};
assign u1_col_in_832 = {col_in_832, u0_col_out_576, reg_intermediate0[576], reg_intermediate1[576]};
assign u1_col_in_833 = {col_in_833, u0_col_out_577, reg_intermediate0[577], reg_intermediate1[577]};
assign u1_col_in_834 = {col_in_834, u0_col_out_578, reg_intermediate0[578], reg_intermediate1[578]};
assign u1_col_in_835 = {col_in_835, u0_col_out_579, reg_intermediate0[579], reg_intermediate1[579]};
assign u1_col_in_836 = {col_in_836, u0_col_out_580, reg_intermediate0[580], reg_intermediate1[580]};
assign u1_col_in_837 = {col_in_837, u0_col_out_581, reg_intermediate0[581], reg_intermediate1[581]};
assign u1_col_in_838 = {col_in_838, u0_col_out_582, reg_intermediate0[582], reg_intermediate1[582]};
assign u1_col_in_839 = {col_in_839, u0_col_out_583, reg_intermediate0[583], reg_intermediate1[583]};
assign u1_col_in_840 = {col_in_840, u0_col_out_584, reg_intermediate0[584], reg_intermediate1[584]};
assign u1_col_in_841 = {col_in_841, u0_col_out_585, reg_intermediate0[585], reg_intermediate1[585]};
assign u1_col_in_842 = {col_in_842, u0_col_out_586, reg_intermediate0[586], reg_intermediate1[586]};
assign u1_col_in_843 = {col_in_843, u0_col_out_587, reg_intermediate0[587], reg_intermediate1[587]};
assign u1_col_in_844 = {col_in_844, u0_col_out_588, reg_intermediate0[588], reg_intermediate1[588]};
assign u1_col_in_845 = {col_in_845, u0_col_out_589, reg_intermediate0[589], reg_intermediate1[589]};
assign u1_col_in_846 = {col_in_846, u0_col_out_590, reg_intermediate0[590], reg_intermediate1[590]};
assign u1_col_in_847 = {col_in_847, u0_col_out_591, reg_intermediate0[591], reg_intermediate1[591]};
assign u1_col_in_848 = {col_in_848, u0_col_out_592, reg_intermediate0[592], reg_intermediate1[592]};
assign u1_col_in_849 = {col_in_849, u0_col_out_593, reg_intermediate0[593], reg_intermediate1[593]};
assign u1_col_in_850 = {col_in_850, u0_col_out_594, reg_intermediate0[594], reg_intermediate1[594]};
assign u1_col_in_851 = {col_in_851, u0_col_out_595, reg_intermediate0[595], reg_intermediate1[595]};
assign u1_col_in_852 = {col_in_852, u0_col_out_596, reg_intermediate0[596], reg_intermediate1[596]};
assign u1_col_in_853 = {col_in_853, u0_col_out_597, reg_intermediate0[597], reg_intermediate1[597]};
assign u1_col_in_854 = {col_in_854, u0_col_out_598, reg_intermediate0[598], reg_intermediate1[598]};
assign u1_col_in_855 = {col_in_855, u0_col_out_599, reg_intermediate0[599], reg_intermediate1[599]};
assign u1_col_in_856 = {col_in_856, u0_col_out_600, reg_intermediate0[600], reg_intermediate1[600]};
assign u1_col_in_857 = {col_in_857, u0_col_out_601, reg_intermediate0[601], reg_intermediate1[601]};
assign u1_col_in_858 = {col_in_858, u0_col_out_602, reg_intermediate0[602], reg_intermediate1[602]};
assign u1_col_in_859 = {col_in_859, u0_col_out_603, reg_intermediate0[603], reg_intermediate1[603]};
assign u1_col_in_860 = {col_in_860, u0_col_out_604, reg_intermediate0[604], reg_intermediate1[604]};
assign u1_col_in_861 = {col_in_861, u0_col_out_605, reg_intermediate0[605], reg_intermediate1[605]};
assign u1_col_in_862 = {col_in_862, u0_col_out_606, reg_intermediate0[606], reg_intermediate1[606]};
assign u1_col_in_863 = {col_in_863, u0_col_out_607, reg_intermediate0[607], reg_intermediate1[607]};
assign u1_col_in_864 = {col_in_864, u0_col_out_608, reg_intermediate0[608], reg_intermediate1[608]};
assign u1_col_in_865 = {col_in_865, u0_col_out_609, reg_intermediate0[609], reg_intermediate1[609]};
assign u1_col_in_866 = {col_in_866, u0_col_out_610, reg_intermediate0[610], reg_intermediate1[610]};
assign u1_col_in_867 = {col_in_867, u0_col_out_611, reg_intermediate0[611], reg_intermediate1[611]};
assign u1_col_in_868 = {col_in_868, u0_col_out_612, reg_intermediate0[612], reg_intermediate1[612]};
assign u1_col_in_869 = {col_in_869, u0_col_out_613, reg_intermediate0[613], reg_intermediate1[613]};
assign u1_col_in_870 = {col_in_870, u0_col_out_614, reg_intermediate0[614], reg_intermediate1[614]};
assign u1_col_in_871 = {col_in_871, u0_col_out_615, reg_intermediate0[615], reg_intermediate1[615]};
assign u1_col_in_872 = {col_in_872, u0_col_out_616, reg_intermediate0[616], reg_intermediate1[616]};
assign u1_col_in_873 = {col_in_873, u0_col_out_617, reg_intermediate0[617], reg_intermediate1[617]};
assign u1_col_in_874 = {col_in_874, u0_col_out_618, reg_intermediate0[618], reg_intermediate1[618]};
assign u1_col_in_875 = {col_in_875, u0_col_out_619, reg_intermediate0[619], reg_intermediate1[619]};
assign u1_col_in_876 = {col_in_876, u0_col_out_620, reg_intermediate0[620], reg_intermediate1[620]};
assign u1_col_in_877 = {col_in_877, u0_col_out_621, reg_intermediate0[621], reg_intermediate1[621]};
assign u1_col_in_878 = {col_in_878, u0_col_out_622, reg_intermediate0[622], reg_intermediate1[622]};
assign u1_col_in_879 = {col_in_879, u0_col_out_623, reg_intermediate0[623], reg_intermediate1[623]};
assign u1_col_in_880 = {col_in_880, u0_col_out_624, reg_intermediate0[624], reg_intermediate1[624]};
assign u1_col_in_881 = {col_in_881, u0_col_out_625, reg_intermediate0[625], reg_intermediate1[625]};
assign u1_col_in_882 = {col_in_882, u0_col_out_626, reg_intermediate0[626], reg_intermediate1[626]};
assign u1_col_in_883 = {col_in_883, u0_col_out_627, reg_intermediate0[627], reg_intermediate1[627]};
assign u1_col_in_884 = {col_in_884, u0_col_out_628, reg_intermediate0[628], reg_intermediate1[628]};
assign u1_col_in_885 = {col_in_885, u0_col_out_629, reg_intermediate0[629], reg_intermediate1[629]};
assign u1_col_in_886 = {col_in_886, u0_col_out_630, reg_intermediate0[630], reg_intermediate1[630]};
assign u1_col_in_887 = {col_in_887, u0_col_out_631, reg_intermediate0[631], reg_intermediate1[631]};
assign u1_col_in_888 = {col_in_888, u0_col_out_632, reg_intermediate0[632], reg_intermediate1[632]};
assign u1_col_in_889 = {col_in_889, u0_col_out_633, reg_intermediate0[633], reg_intermediate1[633]};
assign u1_col_in_890 = {col_in_890, u0_col_out_634, reg_intermediate0[634], reg_intermediate1[634]};
assign u1_col_in_891 = {col_in_891, u0_col_out_635, reg_intermediate0[635], reg_intermediate1[635]};
assign u1_col_in_892 = {col_in_892, u0_col_out_636, reg_intermediate0[636], reg_intermediate1[636]};
assign u1_col_in_893 = {col_in_893, u0_col_out_637, reg_intermediate0[637], reg_intermediate1[637]};
assign u1_col_in_894 = {col_in_894, u0_col_out_638, reg_intermediate0[638], reg_intermediate1[638]};
assign u1_col_in_895 = {col_in_895, u0_col_out_639, reg_intermediate0[639], reg_intermediate1[639]};
assign u1_col_in_896 = {col_in_896, u0_col_out_640, reg_intermediate0[640], reg_intermediate1[640]};
assign u1_col_in_897 = {col_in_897, u0_col_out_641, reg_intermediate0[641], reg_intermediate1[641]};
assign u1_col_in_898 = {col_in_898, u0_col_out_642, reg_intermediate0[642], reg_intermediate1[642]};
assign u1_col_in_899 = {col_in_899, u0_col_out_643, reg_intermediate0[643], reg_intermediate1[643]};
assign u1_col_in_900 = {col_in_900, u0_col_out_644, reg_intermediate0[644], reg_intermediate1[644]};
assign u1_col_in_901 = {col_in_901, u0_col_out_645, reg_intermediate0[645], reg_intermediate1[645]};
assign u1_col_in_902 = {col_in_902, u0_col_out_646, reg_intermediate0[646], reg_intermediate1[646]};
assign u1_col_in_903 = {col_in_903, u0_col_out_647, reg_intermediate0[647], reg_intermediate1[647]};
assign u1_col_in_904 = {col_in_904, u0_col_out_648, reg_intermediate0[648], reg_intermediate1[648]};
assign u1_col_in_905 = {col_in_905, u0_col_out_649, reg_intermediate0[649], reg_intermediate1[649]};
assign u1_col_in_906 = {col_in_906, u0_col_out_650, reg_intermediate0[650], reg_intermediate1[650]};
assign u1_col_in_907 = {col_in_907, u0_col_out_651, reg_intermediate0[651], reg_intermediate1[651]};
assign u1_col_in_908 = {col_in_908, u0_col_out_652, reg_intermediate0[652], reg_intermediate1[652]};
assign u1_col_in_909 = {col_in_909, u0_col_out_653, reg_intermediate0[653], reg_intermediate1[653]};
assign u1_col_in_910 = {col_in_910, u0_col_out_654, reg_intermediate0[654], reg_intermediate1[654]};
assign u1_col_in_911 = {col_in_911, u0_col_out_655, reg_intermediate0[655], reg_intermediate1[655]};
assign u1_col_in_912 = {col_in_912, u0_col_out_656, reg_intermediate0[656], reg_intermediate1[656]};
assign u1_col_in_913 = {col_in_913, u0_col_out_657, reg_intermediate0[657], reg_intermediate1[657]};
assign u1_col_in_914 = {col_in_914, u0_col_out_658, reg_intermediate0[658], reg_intermediate1[658]};
assign u1_col_in_915 = {col_in_915, u0_col_out_659, reg_intermediate0[659], reg_intermediate1[659]};
assign u1_col_in_916 = {col_in_916, u0_col_out_660, reg_intermediate0[660], reg_intermediate1[660]};
assign u1_col_in_917 = {col_in_917, u0_col_out_661, reg_intermediate0[661], reg_intermediate1[661]};
assign u1_col_in_918 = {col_in_918, u0_col_out_662, reg_intermediate0[662], reg_intermediate1[662]};
assign u1_col_in_919 = {col_in_919, u0_col_out_663, reg_intermediate0[663], reg_intermediate1[663]};
assign u1_col_in_920 = {col_in_920, u0_col_out_664, reg_intermediate0[664], reg_intermediate1[664]};
assign u1_col_in_921 = {col_in_921, u0_col_out_665, reg_intermediate0[665], reg_intermediate1[665]};
assign u1_col_in_922 = {col_in_922, u0_col_out_666, reg_intermediate0[666], reg_intermediate1[666]};
assign u1_col_in_923 = {col_in_923, u0_col_out_667, reg_intermediate0[667], reg_intermediate1[667]};
assign u1_col_in_924 = {col_in_924, u0_col_out_668, reg_intermediate0[668], reg_intermediate1[668]};
assign u1_col_in_925 = {col_in_925, u0_col_out_669, reg_intermediate0[669], reg_intermediate1[669]};
assign u1_col_in_926 = {col_in_926, u0_col_out_670, reg_intermediate0[670], reg_intermediate1[670]};
assign u1_col_in_927 = {col_in_927, u0_col_out_671, reg_intermediate0[671], reg_intermediate1[671]};
assign u1_col_in_928 = {col_in_928, u0_col_out_672, reg_intermediate0[672], reg_intermediate1[672]};
assign u1_col_in_929 = {col_in_929, u0_col_out_673, reg_intermediate0[673], reg_intermediate1[673]};
assign u1_col_in_930 = {col_in_930, u0_col_out_674, reg_intermediate0[674], reg_intermediate1[674]};
assign u1_col_in_931 = {col_in_931, u0_col_out_675, reg_intermediate0[675], reg_intermediate1[675]};
assign u1_col_in_932 = {col_in_932, u0_col_out_676, reg_intermediate0[676], reg_intermediate1[676]};
assign u1_col_in_933 = {col_in_933, u0_col_out_677, reg_intermediate0[677], reg_intermediate1[677]};
assign u1_col_in_934 = {col_in_934, u0_col_out_678, reg_intermediate0[678], reg_intermediate1[678]};
assign u1_col_in_935 = {col_in_935, u0_col_out_679, reg_intermediate0[679], reg_intermediate1[679]};
assign u1_col_in_936 = {col_in_936, u0_col_out_680, reg_intermediate0[680], reg_intermediate1[680]};
assign u1_col_in_937 = {col_in_937, u0_col_out_681, reg_intermediate0[681], reg_intermediate1[681]};
assign u1_col_in_938 = {col_in_938, u0_col_out_682, reg_intermediate0[682], reg_intermediate1[682]};
assign u1_col_in_939 = {col_in_939, u0_col_out_683, reg_intermediate0[683], reg_intermediate1[683]};
assign u1_col_in_940 = {col_in_940, u0_col_out_684, reg_intermediate0[684], reg_intermediate1[684]};
assign u1_col_in_941 = {col_in_941, u0_col_out_685, reg_intermediate0[685], reg_intermediate1[685]};
assign u1_col_in_942 = {col_in_942, u0_col_out_686, reg_intermediate0[686], reg_intermediate1[686]};
assign u1_col_in_943 = {col_in_943, u0_col_out_687, reg_intermediate0[687], reg_intermediate1[687]};
assign u1_col_in_944 = {col_in_944, u0_col_out_688, reg_intermediate0[688], reg_intermediate1[688]};
assign u1_col_in_945 = {col_in_945, u0_col_out_689, reg_intermediate0[689], reg_intermediate1[689]};
assign u1_col_in_946 = {col_in_946, u0_col_out_690, reg_intermediate0[690], reg_intermediate1[690]};
assign u1_col_in_947 = {col_in_947, u0_col_out_691, reg_intermediate0[691], reg_intermediate1[691]};
assign u1_col_in_948 = {col_in_948, u0_col_out_692, reg_intermediate0[692], reg_intermediate1[692]};
assign u1_col_in_949 = {col_in_949, u0_col_out_693, reg_intermediate0[693], reg_intermediate1[693]};
assign u1_col_in_950 = {col_in_950, u0_col_out_694, reg_intermediate0[694], reg_intermediate1[694]};
assign u1_col_in_951 = {col_in_951, u0_col_out_695, reg_intermediate0[695], reg_intermediate1[695]};
assign u1_col_in_952 = {col_in_952, u0_col_out_696, reg_intermediate0[696], reg_intermediate1[696]};
assign u1_col_in_953 = {col_in_953, u0_col_out_697, reg_intermediate0[697], reg_intermediate1[697]};
assign u1_col_in_954 = {col_in_954, u0_col_out_698, reg_intermediate0[698], reg_intermediate1[698]};
assign u1_col_in_955 = {col_in_955, u0_col_out_699, reg_intermediate0[699], reg_intermediate1[699]};
assign u1_col_in_956 = {col_in_956, u0_col_out_700, reg_intermediate0[700], reg_intermediate1[700]};
assign u1_col_in_957 = {col_in_957, u0_col_out_701, reg_intermediate0[701], reg_intermediate1[701]};
assign u1_col_in_958 = {col_in_958, u0_col_out_702, reg_intermediate0[702], reg_intermediate1[702]};
assign u1_col_in_959 = {col_in_959, u0_col_out_703, reg_intermediate0[703], reg_intermediate1[703]};
assign u1_col_in_960 = {col_in_960, u0_col_out_704, reg_intermediate0[704], reg_intermediate1[704]};
assign u1_col_in_961 = {col_in_961, u0_col_out_705, reg_intermediate0[705], reg_intermediate1[705]};
assign u1_col_in_962 = {col_in_962, u0_col_out_706, reg_intermediate0[706], reg_intermediate1[706]};
assign u1_col_in_963 = {col_in_963, u0_col_out_707, reg_intermediate0[707], reg_intermediate1[707]};
assign u1_col_in_964 = {col_in_964, u0_col_out_708, reg_intermediate0[708], reg_intermediate1[708]};
assign u1_col_in_965 = {col_in_965, u0_col_out_709, reg_intermediate0[709], reg_intermediate1[709]};
assign u1_col_in_966 = {col_in_966, u0_col_out_710, reg_intermediate0[710], reg_intermediate1[710]};
assign u1_col_in_967 = {col_in_967, u0_col_out_711, reg_intermediate0[711], reg_intermediate1[711]};
assign u1_col_in_968 = {col_in_968, u0_col_out_712, reg_intermediate0[712], reg_intermediate1[712]};
assign u1_col_in_969 = {col_in_969, u0_col_out_713, reg_intermediate0[713], reg_intermediate1[713]};
assign u1_col_in_970 = {col_in_970, u0_col_out_714, reg_intermediate0[714], reg_intermediate1[714]};
assign u1_col_in_971 = {col_in_971, u0_col_out_715, reg_intermediate0[715], reg_intermediate1[715]};
assign u1_col_in_972 = {col_in_972, u0_col_out_716, reg_intermediate0[716], reg_intermediate1[716]};
assign u1_col_in_973 = {col_in_973, u0_col_out_717, reg_intermediate0[717], reg_intermediate1[717]};
assign u1_col_in_974 = {col_in_974, u0_col_out_718, reg_intermediate0[718], reg_intermediate1[718]};
assign u1_col_in_975 = {col_in_975, u0_col_out_719, reg_intermediate0[719], reg_intermediate1[719]};
assign u1_col_in_976 = {col_in_976, u0_col_out_720, reg_intermediate0[720], reg_intermediate1[720]};
assign u1_col_in_977 = {col_in_977, u0_col_out_721, reg_intermediate0[721], reg_intermediate1[721]};
assign u1_col_in_978 = {col_in_978, u0_col_out_722, reg_intermediate0[722], reg_intermediate1[722]};
assign u1_col_in_979 = {col_in_979, u0_col_out_723, reg_intermediate0[723], reg_intermediate1[723]};
assign u1_col_in_980 = {col_in_980, u0_col_out_724, reg_intermediate0[724], reg_intermediate1[724]};
assign u1_col_in_981 = {col_in_981, u0_col_out_725, reg_intermediate0[725], reg_intermediate1[725]};
assign u1_col_in_982 = {col_in_982, u0_col_out_726, reg_intermediate0[726], reg_intermediate1[726]};
assign u1_col_in_983 = {col_in_983, u0_col_out_727, reg_intermediate0[727], reg_intermediate1[727]};
assign u1_col_in_984 = {col_in_984, u0_col_out_728, reg_intermediate0[728], reg_intermediate1[728]};
assign u1_col_in_985 = {col_in_985, u0_col_out_729, reg_intermediate0[729], reg_intermediate1[729]};
assign u1_col_in_986 = {col_in_986, u0_col_out_730, reg_intermediate0[730], reg_intermediate1[730]};
assign u1_col_in_987 = {col_in_987, u0_col_out_731, reg_intermediate0[731], reg_intermediate1[731]};
assign u1_col_in_988 = {col_in_988, u0_col_out_732, reg_intermediate0[732], reg_intermediate1[732]};
assign u1_col_in_989 = {col_in_989, u0_col_out_733, reg_intermediate0[733], reg_intermediate1[733]};
assign u1_col_in_990 = {col_in_990, u0_col_out_734, reg_intermediate0[734], reg_intermediate1[734]};
assign u1_col_in_991 = {col_in_991, u0_col_out_735, reg_intermediate0[735], reg_intermediate1[735]};
assign u1_col_in_992 = {col_in_992, u0_col_out_736, reg_intermediate0[736], reg_intermediate1[736]};
assign u1_col_in_993 = {col_in_993, u0_col_out_737, reg_intermediate0[737], reg_intermediate1[737]};
assign u1_col_in_994 = {col_in_994, u0_col_out_738, reg_intermediate0[738], reg_intermediate1[738]};
assign u1_col_in_995 = {col_in_995, u0_col_out_739, reg_intermediate0[739], reg_intermediate1[739]};
assign u1_col_in_996 = {col_in_996, u0_col_out_740, reg_intermediate0[740], reg_intermediate1[740]};
assign u1_col_in_997 = {col_in_997, u0_col_out_741, reg_intermediate0[741], reg_intermediate1[741]};
assign u1_col_in_998 = {col_in_998, u0_col_out_742, reg_intermediate0[742], reg_intermediate1[742]};
assign u1_col_in_999 = {col_in_999, u0_col_out_743, reg_intermediate0[743], reg_intermediate1[743]};
assign u1_col_in_1000 = {col_in_1000, u0_col_out_744, reg_intermediate0[744], reg_intermediate1[744]};
assign u1_col_in_1001 = {col_in_1001, u0_col_out_745, reg_intermediate0[745], reg_intermediate1[745]};
assign u1_col_in_1002 = {col_in_1002, u0_col_out_746, reg_intermediate0[746], reg_intermediate1[746]};
assign u1_col_in_1003 = {col_in_1003, u0_col_out_747, reg_intermediate0[747], reg_intermediate1[747]};
assign u1_col_in_1004 = {col_in_1004, u0_col_out_748, reg_intermediate0[748], reg_intermediate1[748]};
assign u1_col_in_1005 = {col_in_1005, u0_col_out_749, reg_intermediate0[749], reg_intermediate1[749]};
assign u1_col_in_1006 = {col_in_1006, u0_col_out_750, reg_intermediate0[750], reg_intermediate1[750]};
assign u1_col_in_1007 = {col_in_1007, u0_col_out_751, reg_intermediate0[751], reg_intermediate1[751]};
assign u1_col_in_1008 = {col_in_1008, u0_col_out_752, reg_intermediate0[752], reg_intermediate1[752]};
assign u1_col_in_1009 = {col_in_1009, u0_col_out_753, reg_intermediate0[753], reg_intermediate1[753]};
assign u1_col_in_1010 = {col_in_1010, u0_col_out_754, reg_intermediate0[754], reg_intermediate1[754]};
assign u1_col_in_1011 = {col_in_1011, u0_col_out_755, reg_intermediate0[755], reg_intermediate1[755]};
assign u1_col_in_1012 = {col_in_1012, u0_col_out_756, reg_intermediate0[756], reg_intermediate1[756]};
assign u1_col_in_1013 = {col_in_1013, u0_col_out_757, reg_intermediate0[757], reg_intermediate1[757]};
assign u1_col_in_1014 = {col_in_1014, u0_col_out_758, reg_intermediate0[758], reg_intermediate1[758]};
assign u1_col_in_1015 = {col_in_1015, u0_col_out_759, reg_intermediate0[759], reg_intermediate1[759]};
assign u1_col_in_1016 = {col_in_1016, u0_col_out_760, reg_intermediate0[760], reg_intermediate1[760]};
assign u1_col_in_1017 = {col_in_1017, u0_col_out_761, reg_intermediate0[761], reg_intermediate1[761]};
assign u1_col_in_1018 = {col_in_1018, u0_col_out_762, reg_intermediate0[762], reg_intermediate1[762]};
assign u1_col_in_1019 = {col_in_1019, u0_col_out_763, reg_intermediate0[763], reg_intermediate1[763]};
assign u1_col_in_1020 = {col_in_1020, u0_col_out_764, reg_intermediate0[764], reg_intermediate1[764]};
assign u1_col_in_1021 = {col_in_1021, u0_col_out_765, reg_intermediate0[765], reg_intermediate1[765]};
assign u1_col_in_1022 = {col_in_1022, u0_col_out_766, reg_intermediate0[766], reg_intermediate1[766]};
assign u1_col_in_1023 = {col_in_1023, u0_col_out_767, reg_intermediate0[767], reg_intermediate1[767]};
assign u1_col_in_1024 = {col_in_1024, u0_col_out_768, reg_intermediate0[768], reg_intermediate1[768]};
assign u1_col_in_1025 = {col_in_1025, u0_col_out_769, reg_intermediate0[769], reg_intermediate1[769]};
assign u1_col_in_1026 = {col_in_1026, u0_col_out_770, reg_intermediate0[770], reg_intermediate1[770]};
assign u1_col_in_1027 = {col_in_1027, u0_col_out_771, reg_intermediate0[771], reg_intermediate1[771]};
assign u1_col_in_1028 = {col_in_1028, u0_col_out_772, reg_intermediate0[772], reg_intermediate1[772]};
assign u1_col_in_1029 = {col_in_1029, u0_col_out_773, reg_intermediate0[773], reg_intermediate1[773]};
assign u1_col_in_1030 = {col_in_1030, u0_col_out_774, reg_intermediate0[774], reg_intermediate1[774]};
assign u1_col_in_1031 = {col_in_1031, u0_col_out_775, reg_intermediate0[775], reg_intermediate1[775]};
assign u1_col_in_1032 = {col_in_1032, u0_col_out_776, reg_intermediate0[776], reg_intermediate1[776]};
assign u1_col_in_1033 = {col_in_1033, u0_col_out_777, reg_intermediate0[777], reg_intermediate1[777]};
assign u1_col_in_1034 = {col_in_1034, u0_col_out_778, reg_intermediate0[778], reg_intermediate1[778]};
assign u1_col_in_1035 = {col_in_1035, u0_col_out_779, reg_intermediate0[779], reg_intermediate1[779]};
assign u1_col_in_1036 = {col_in_1036, u0_col_out_780, reg_intermediate0[780], reg_intermediate1[780]};
assign u1_col_in_1037 = {col_in_1037, u0_col_out_781, reg_intermediate0[781], reg_intermediate1[781]};
assign u1_col_in_1038 = {col_in_1038, u0_col_out_782, reg_intermediate0[782], reg_intermediate1[782]};
assign u1_col_in_1039 = {col_in_1039, u0_col_out_783, reg_intermediate0[783], reg_intermediate1[783]};
assign u1_col_in_1040 = {col_in_1040, u0_col_out_784, reg_intermediate0[784], reg_intermediate1[784]};
assign u1_col_in_1041 = {col_in_1041, u0_col_out_785, reg_intermediate0[785], reg_intermediate1[785]};
assign u1_col_in_1042 = {col_in_1042, u0_col_out_786, reg_intermediate0[786], reg_intermediate1[786]};
assign u1_col_in_1043 = {col_in_1043, u0_col_out_787, reg_intermediate0[787], reg_intermediate1[787]};
assign u1_col_in_1044 = {col_in_1044, u0_col_out_788, reg_intermediate0[788], reg_intermediate1[788]};
assign u1_col_in_1045 = {col_in_1045, u0_col_out_789, reg_intermediate0[789], reg_intermediate1[789]};
assign u1_col_in_1046 = {col_in_1046, u0_col_out_790, reg_intermediate0[790], reg_intermediate1[790]};
assign u1_col_in_1047 = {col_in_1047, u0_col_out_791, reg_intermediate0[791], reg_intermediate1[791]};
assign u1_col_in_1048 = {col_in_1048, u0_col_out_792, reg_intermediate0[792], reg_intermediate1[792]};
assign u1_col_in_1049 = {col_in_1049, u0_col_out_793, reg_intermediate0[793], reg_intermediate1[793]};
assign u1_col_in_1050 = {col_in_1050, u0_col_out_794, reg_intermediate0[794], reg_intermediate1[794]};
assign u1_col_in_1051 = {col_in_1051, u0_col_out_795, reg_intermediate0[795], reg_intermediate1[795]};
assign u1_col_in_1052 = {col_in_1052, u0_col_out_796, reg_intermediate0[796], reg_intermediate1[796]};
assign u1_col_in_1053 = {col_in_1053, u0_col_out_797, reg_intermediate0[797], reg_intermediate1[797]};
assign u1_col_in_1054 = {col_in_1054, u0_col_out_798, reg_intermediate0[798], reg_intermediate1[798]};
assign u1_col_in_1055 = {col_in_1055, u0_col_out_799, reg_intermediate0[799], reg_intermediate1[799]};
assign u1_col_in_1056 = {col_in_1056, u0_col_out_800, reg_intermediate0[800], reg_intermediate1[800]};
assign u1_col_in_1057 = {col_in_1057, u0_col_out_801, reg_intermediate0[801], reg_intermediate1[801]};
assign u1_col_in_1058 = {col_in_1058, u0_col_out_802, reg_intermediate0[802], reg_intermediate1[802]};
assign u1_col_in_1059 = {col_in_1059, u0_col_out_803, reg_intermediate0[803], reg_intermediate1[803]};
assign u1_col_in_1060 = {col_in_1060, u0_col_out_804, reg_intermediate0[804], reg_intermediate1[804]};
assign u1_col_in_1061 = {col_in_1061, u0_col_out_805, reg_intermediate0[805], reg_intermediate1[805]};
assign u1_col_in_1062 = {col_in_1062, u0_col_out_806, reg_intermediate0[806], reg_intermediate1[806]};
assign u1_col_in_1063 = {col_in_1063, u0_col_out_807, reg_intermediate0[807], reg_intermediate1[807]};
assign u1_col_in_1064 = {col_in_1064, u0_col_out_808, reg_intermediate0[808], reg_intermediate1[808]};
assign u1_col_in_1065 = {col_in_1065, u0_col_out_809, reg_intermediate0[809], reg_intermediate1[809]};
assign u1_col_in_1066 = {col_in_1066, u0_col_out_810, reg_intermediate0[810], reg_intermediate1[810]};
assign u1_col_in_1067 = {col_in_1067, u0_col_out_811, reg_intermediate0[811], reg_intermediate1[811]};
assign u1_col_in_1068 = {col_in_1068, u0_col_out_812, reg_intermediate0[812], reg_intermediate1[812]};
assign u1_col_in_1069 = {col_in_1069, u0_col_out_813, reg_intermediate0[813], reg_intermediate1[813]};
assign u1_col_in_1070 = {col_in_1070, u0_col_out_814, reg_intermediate0[814], reg_intermediate1[814]};
assign u1_col_in_1071 = {col_in_1071, u0_col_out_815, reg_intermediate0[815], reg_intermediate1[815]};
assign u1_col_in_1072 = {col_in_1072, u0_col_out_816, reg_intermediate0[816], reg_intermediate1[816]};
assign u1_col_in_1073 = {col_in_1073, u0_col_out_817, reg_intermediate0[817], reg_intermediate1[817]};
assign u1_col_in_1074 = {col_in_1074, u0_col_out_818, reg_intermediate0[818], reg_intermediate1[818]};
assign u1_col_in_1075 = {col_in_1075, u0_col_out_819, reg_intermediate0[819], reg_intermediate1[819]};
assign u1_col_in_1076 = {col_in_1076, u0_col_out_820, reg_intermediate0[820], reg_intermediate1[820]};
assign u1_col_in_1077 = {col_in_1077, u0_col_out_821, reg_intermediate0[821], reg_intermediate1[821]};
assign u1_col_in_1078 = {col_in_1078, u0_col_out_822, reg_intermediate0[822], reg_intermediate1[822]};
assign u1_col_in_1079 = {col_in_1079, u0_col_out_823, reg_intermediate0[823], reg_intermediate1[823]};
assign u1_col_in_1080 = {col_in_1080, u0_col_out_824, reg_intermediate0[824], reg_intermediate1[824]};
assign u1_col_in_1081 = {col_in_1081, u0_col_out_825, reg_intermediate0[825], reg_intermediate1[825]};
assign u1_col_in_1082 = {col_in_1082, u0_col_out_826, reg_intermediate0[826], reg_intermediate1[826]};
assign u1_col_in_1083 = {col_in_1083, u0_col_out_827, reg_intermediate0[827], reg_intermediate1[827]};
assign u1_col_in_1084 = {col_in_1084, u0_col_out_828, reg_intermediate0[828], reg_intermediate1[828]};
assign u1_col_in_1085 = {col_in_1085, u0_col_out_829, reg_intermediate0[829], reg_intermediate1[829]};
assign u1_col_in_1086 = {col_in_1086, u0_col_out_830, reg_intermediate0[830], reg_intermediate1[830]};
assign u1_col_in_1087 = {col_in_1087, u0_col_out_831, reg_intermediate0[831], reg_intermediate1[831]};
assign u1_col_in_1088 = {col_in_1088, u0_col_out_832, reg_intermediate0[832], reg_intermediate1[832]};
assign u1_col_in_1089 = {col_in_1089, u0_col_out_833, reg_intermediate0[833], reg_intermediate1[833]};
assign u1_col_in_1090 = {col_in_1090, u0_col_out_834, reg_intermediate0[834], reg_intermediate1[834]};
assign u1_col_in_1091 = {col_in_1091, u0_col_out_835, reg_intermediate0[835], reg_intermediate1[835]};
assign u1_col_in_1092 = {col_in_1092, u0_col_out_836, reg_intermediate0[836], reg_intermediate1[836]};
assign u1_col_in_1093 = {col_in_1093, u0_col_out_837, reg_intermediate0[837], reg_intermediate1[837]};
assign u1_col_in_1094 = {col_in_1094, u0_col_out_838, reg_intermediate0[838], reg_intermediate1[838]};
assign u1_col_in_1095 = {col_in_1095, u0_col_out_839, reg_intermediate0[839], reg_intermediate1[839]};
assign u1_col_in_1096 = {col_in_1096, u0_col_out_840, reg_intermediate0[840], reg_intermediate1[840]};
assign u1_col_in_1097 = {col_in_1097, u0_col_out_841, reg_intermediate0[841], reg_intermediate1[841]};
assign u1_col_in_1098 = {col_in_1098, u0_col_out_842, reg_intermediate0[842], reg_intermediate1[842]};
assign u1_col_in_1099 = {col_in_1099, u0_col_out_843, reg_intermediate0[843], reg_intermediate1[843]};
assign u1_col_in_1100 = {col_in_1100, u0_col_out_844, reg_intermediate0[844], reg_intermediate1[844]};
assign u1_col_in_1101 = {col_in_1101, u0_col_out_845, reg_intermediate0[845], reg_intermediate1[845]};
assign u1_col_in_1102 = {col_in_1102, u0_col_out_846, reg_intermediate0[846], reg_intermediate1[846]};
assign u1_col_in_1103 = {col_in_1103, u0_col_out_847, reg_intermediate0[847], reg_intermediate1[847]};
assign u1_col_in_1104 = {col_in_1104, u0_col_out_848, reg_intermediate0[848], reg_intermediate1[848]};
assign u1_col_in_1105 = {col_in_1105, u0_col_out_849, reg_intermediate0[849], reg_intermediate1[849]};
assign u1_col_in_1106 = {col_in_1106, u0_col_out_850, reg_intermediate0[850], reg_intermediate1[850]};
assign u1_col_in_1107 = {col_in_1107, u0_col_out_851, reg_intermediate0[851], reg_intermediate1[851]};
assign u1_col_in_1108 = {col_in_1108, u0_col_out_852, reg_intermediate0[852], reg_intermediate1[852]};
assign u1_col_in_1109 = {col_in_1109, u0_col_out_853, reg_intermediate0[853], reg_intermediate1[853]};
assign u1_col_in_1110 = {col_in_1110, u0_col_out_854, reg_intermediate0[854], reg_intermediate1[854]};
assign u1_col_in_1111 = {col_in_1111, u0_col_out_855, reg_intermediate0[855], reg_intermediate1[855]};
assign u1_col_in_1112 = {col_in_1112, u0_col_out_856, reg_intermediate0[856], reg_intermediate1[856]};
assign u1_col_in_1113 = {col_in_1113, u0_col_out_857, reg_intermediate0[857], reg_intermediate1[857]};
assign u1_col_in_1114 = {col_in_1114, u0_col_out_858, reg_intermediate0[858], reg_intermediate1[858]};
assign u1_col_in_1115 = {col_in_1115, u0_col_out_859, reg_intermediate0[859], reg_intermediate1[859]};
assign u1_col_in_1116 = {col_in_1116, u0_col_out_860, reg_intermediate0[860], reg_intermediate1[860]};
assign u1_col_in_1117 = {col_in_1117, u0_col_out_861, reg_intermediate0[861], reg_intermediate1[861]};
assign u1_col_in_1118 = {col_in_1118, u0_col_out_862, reg_intermediate0[862], reg_intermediate1[862]};
assign u1_col_in_1119 = {col_in_1119, u0_col_out_863, reg_intermediate0[863], reg_intermediate1[863]};
assign u1_col_in_1120 = {col_in_1120, u0_col_out_864, reg_intermediate0[864], reg_intermediate1[864]};
assign u1_col_in_1121 = {col_in_1121, u0_col_out_865, reg_intermediate0[865], reg_intermediate1[865]};
assign u1_col_in_1122 = {col_in_1122, u0_col_out_866, reg_intermediate0[866], reg_intermediate1[866]};
assign u1_col_in_1123 = {col_in_1123, u0_col_out_867, reg_intermediate0[867], reg_intermediate1[867]};
assign u1_col_in_1124 = {col_in_1124, u0_col_out_868, reg_intermediate0[868], reg_intermediate1[868]};
assign u1_col_in_1125 = {col_in_1125, u0_col_out_869, reg_intermediate0[869], reg_intermediate1[869]};
assign u1_col_in_1126 = {col_in_1126, u0_col_out_870, reg_intermediate0[870], reg_intermediate1[870]};
assign u1_col_in_1127 = {col_in_1127, u0_col_out_871, reg_intermediate0[871], reg_intermediate1[871]};
assign u1_col_in_1128 = {col_in_1128, u0_col_out_872, reg_intermediate0[872], reg_intermediate1[872]};
assign u1_col_in_1129 = {col_in_1129, u0_col_out_873, reg_intermediate0[873], reg_intermediate1[873]};
assign u1_col_in_1130 = {col_in_1130, u0_col_out_874, reg_intermediate0[874], reg_intermediate1[874]};
assign u1_col_in_1131 = {col_in_1131, u0_col_out_875, reg_intermediate0[875], reg_intermediate1[875]};
assign u1_col_in_1132 = {col_in_1132, u0_col_out_876, reg_intermediate0[876], reg_intermediate1[876]};
assign u1_col_in_1133 = {col_in_1133, u0_col_out_877, reg_intermediate0[877], reg_intermediate1[877]};
assign u1_col_in_1134 = {col_in_1134, u0_col_out_878, reg_intermediate0[878], reg_intermediate1[878]};
assign u1_col_in_1135 = {col_in_1135, u0_col_out_879, reg_intermediate0[879], reg_intermediate1[879]};
assign u1_col_in_1136 = {col_in_1136, u0_col_out_880, reg_intermediate0[880], reg_intermediate1[880]};
assign u1_col_in_1137 = {col_in_1137, u0_col_out_881, reg_intermediate0[881], reg_intermediate1[881]};
assign u1_col_in_1138 = {col_in_1138, u0_col_out_882, reg_intermediate0[882], reg_intermediate1[882]};
assign u1_col_in_1139 = {col_in_1139, u0_col_out_883, reg_intermediate0[883], reg_intermediate1[883]};
assign u1_col_in_1140 = {col_in_1140, u0_col_out_884, reg_intermediate0[884], reg_intermediate1[884]};
assign u1_col_in_1141 = {col_in_1141, u0_col_out_885, reg_intermediate0[885], reg_intermediate1[885]};
assign u1_col_in_1142 = {col_in_1142, u0_col_out_886, reg_intermediate0[886], reg_intermediate1[886]};
assign u1_col_in_1143 = {col_in_1143, u0_col_out_887, reg_intermediate0[887], reg_intermediate1[887]};
assign u1_col_in_1144 = {col_in_1144, u0_col_out_888, reg_intermediate0[888], reg_intermediate1[888]};
assign u1_col_in_1145 = {col_in_1145, u0_col_out_889, reg_intermediate0[889], reg_intermediate1[889]};
assign u1_col_in_1146 = {col_in_1146, u0_col_out_890, reg_intermediate0[890], reg_intermediate1[890]};
assign u1_col_in_1147 = {col_in_1147, u0_col_out_891, reg_intermediate0[891], reg_intermediate1[891]};
assign u1_col_in_1148 = {col_in_1148, u0_col_out_892, reg_intermediate0[892], reg_intermediate1[892]};
assign u1_col_in_1149 = {col_in_1149, u0_col_out_893, reg_intermediate0[893], reg_intermediate1[893]};
assign u1_col_in_1150 = {col_in_1150, u0_col_out_894, reg_intermediate0[894], reg_intermediate1[894]};
assign u1_col_in_1151 = {col_in_1151, u0_col_out_895, reg_intermediate0[895], reg_intermediate1[895]};
assign u1_col_in_1152 = {col_in_1152, u0_col_out_896, reg_intermediate0[896], reg_intermediate1[896]};
assign u1_col_in_1153 = {col_in_1153, u0_col_out_897, reg_intermediate0[897], reg_intermediate1[897]};
assign u1_col_in_1154 = {col_in_1154, u0_col_out_898, reg_intermediate0[898], reg_intermediate1[898]};
assign u1_col_in_1155 = {col_in_1155, u0_col_out_899, reg_intermediate0[899], reg_intermediate1[899]};
assign u1_col_in_1156 = {col_in_1156, u0_col_out_900, reg_intermediate0[900], reg_intermediate1[900]};
assign u1_col_in_1157 = {col_in_1157, u0_col_out_901, reg_intermediate0[901], reg_intermediate1[901]};
assign u1_col_in_1158 = {col_in_1158, u0_col_out_902, reg_intermediate0[902], reg_intermediate1[902]};
assign u1_col_in_1159 = {col_in_1159, u0_col_out_903, reg_intermediate0[903], reg_intermediate1[903]};
assign u1_col_in_1160 = {col_in_1160, u0_col_out_904, reg_intermediate0[904], reg_intermediate1[904]};
assign u1_col_in_1161 = {col_in_1161, u0_col_out_905, reg_intermediate0[905], reg_intermediate1[905]};
assign u1_col_in_1162 = {col_in_1162, u0_col_out_906, reg_intermediate0[906], reg_intermediate1[906]};
assign u1_col_in_1163 = {col_in_1163, u0_col_out_907, reg_intermediate0[907], reg_intermediate1[907]};
assign u1_col_in_1164 = {col_in_1164, u0_col_out_908, reg_intermediate0[908], reg_intermediate1[908]};
assign u1_col_in_1165 = {col_in_1165, u0_col_out_909, reg_intermediate0[909], reg_intermediate1[909]};
assign u1_col_in_1166 = {col_in_1166, u0_col_out_910, reg_intermediate0[910], reg_intermediate1[910]};
assign u1_col_in_1167 = {col_in_1167, u0_col_out_911, reg_intermediate0[911], reg_intermediate1[911]};
assign u1_col_in_1168 = {col_in_1168, u0_col_out_912, reg_intermediate0[912], reg_intermediate1[912]};
assign u1_col_in_1169 = {col_in_1169, u0_col_out_913, reg_intermediate0[913], reg_intermediate1[913]};
assign u1_col_in_1170 = {col_in_1170, u0_col_out_914, reg_intermediate0[914], reg_intermediate1[914]};
assign u1_col_in_1171 = {col_in_1171, u0_col_out_915, reg_intermediate0[915], reg_intermediate1[915]};
assign u1_col_in_1172 = {col_in_1172, u0_col_out_916, reg_intermediate0[916], reg_intermediate1[916]};
assign u1_col_in_1173 = {col_in_1173, u0_col_out_917, reg_intermediate0[917], reg_intermediate1[917]};
assign u1_col_in_1174 = {col_in_1174, u0_col_out_918, reg_intermediate0[918], reg_intermediate1[918]};
assign u1_col_in_1175 = {col_in_1175, u0_col_out_919, reg_intermediate0[919], reg_intermediate1[919]};
assign u1_col_in_1176 = {col_in_1176, u0_col_out_920, reg_intermediate0[920], reg_intermediate1[920]};
assign u1_col_in_1177 = {col_in_1177, u0_col_out_921, reg_intermediate0[921], reg_intermediate1[921]};
assign u1_col_in_1178 = {col_in_1178, u0_col_out_922, reg_intermediate0[922], reg_intermediate1[922]};
assign u1_col_in_1179 = {col_in_1179, u0_col_out_923, reg_intermediate0[923], reg_intermediate1[923]};
assign u1_col_in_1180 = {col_in_1180, u0_col_out_924, reg_intermediate0[924], reg_intermediate1[924]};
assign u1_col_in_1181 = {col_in_1181, u0_col_out_925, reg_intermediate0[925], reg_intermediate1[925]};
assign u1_col_in_1182 = {col_in_1182, u0_col_out_926, reg_intermediate0[926], reg_intermediate1[926]};
assign u1_col_in_1183 = {col_in_1183, u0_col_out_927, reg_intermediate0[927], reg_intermediate1[927]};
assign u1_col_in_1184 = {col_in_1184, u0_col_out_928, reg_intermediate0[928], reg_intermediate1[928]};
assign u1_col_in_1185 = {col_in_1185, u0_col_out_929, reg_intermediate0[929], reg_intermediate1[929]};
assign u1_col_in_1186 = {col_in_1186, u0_col_out_930, reg_intermediate0[930], reg_intermediate1[930]};
assign u1_col_in_1187 = {col_in_1187, u0_col_out_931, reg_intermediate0[931], reg_intermediate1[931]};
assign u1_col_in_1188 = {col_in_1188, u0_col_out_932, reg_intermediate0[932], reg_intermediate1[932]};
assign u1_col_in_1189 = {col_in_1189, u0_col_out_933, reg_intermediate0[933], reg_intermediate1[933]};
assign u1_col_in_1190 = {col_in_1190, u0_col_out_934, reg_intermediate0[934], reg_intermediate1[934]};
assign u1_col_in_1191 = {col_in_1191, u0_col_out_935, reg_intermediate0[935], reg_intermediate1[935]};
assign u1_col_in_1192 = {col_in_1192, u0_col_out_936, reg_intermediate0[936], reg_intermediate1[936]};
assign u1_col_in_1193 = {col_in_1193, u0_col_out_937, reg_intermediate0[937], reg_intermediate1[937]};
assign u1_col_in_1194 = {col_in_1194, u0_col_out_938, reg_intermediate0[938], reg_intermediate1[938]};
assign u1_col_in_1195 = {col_in_1195, u0_col_out_939, reg_intermediate0[939], reg_intermediate1[939]};
assign u1_col_in_1196 = {col_in_1196, u0_col_out_940, reg_intermediate0[940], reg_intermediate1[940]};
assign u1_col_in_1197 = {col_in_1197, u0_col_out_941, reg_intermediate0[941], reg_intermediate1[941]};
assign u1_col_in_1198 = {col_in_1198, u0_col_out_942, reg_intermediate0[942], reg_intermediate1[942]};
assign u1_col_in_1199 = {col_in_1199, u0_col_out_943, reg_intermediate0[943], reg_intermediate1[943]};
assign u1_col_in_1200 = {col_in_1200, u0_col_out_944, reg_intermediate0[944], reg_intermediate1[944]};
assign u1_col_in_1201 = {col_in_1201, u0_col_out_945, reg_intermediate0[945], reg_intermediate1[945]};
assign u1_col_in_1202 = {col_in_1202, u0_col_out_946, reg_intermediate0[946], reg_intermediate1[946]};
assign u1_col_in_1203 = {col_in_1203, u0_col_out_947, reg_intermediate0[947], reg_intermediate1[947]};
assign u1_col_in_1204 = {col_in_1204, u0_col_out_948, reg_intermediate0[948], reg_intermediate1[948]};
assign u1_col_in_1205 = {col_in_1205, u0_col_out_949, reg_intermediate0[949], reg_intermediate1[949]};
assign u1_col_in_1206 = {col_in_1206, u0_col_out_950, reg_intermediate0[950], reg_intermediate1[950]};
assign u1_col_in_1207 = {col_in_1207, u0_col_out_951, reg_intermediate0[951], reg_intermediate1[951]};
assign u1_col_in_1208 = {col_in_1208, u0_col_out_952, reg_intermediate0[952], reg_intermediate1[952]};
assign u1_col_in_1209 = {col_in_1209, u0_col_out_953, reg_intermediate0[953], reg_intermediate1[953]};
assign u1_col_in_1210 = {col_in_1210, u0_col_out_954, reg_intermediate0[954], reg_intermediate1[954]};
assign u1_col_in_1211 = {col_in_1211, u0_col_out_955, reg_intermediate0[955], reg_intermediate1[955]};
assign u1_col_in_1212 = {col_in_1212, u0_col_out_956, reg_intermediate0[956], reg_intermediate1[956]};
assign u1_col_in_1213 = {col_in_1213, u0_col_out_957, reg_intermediate0[957], reg_intermediate1[957]};
assign u1_col_in_1214 = {col_in_1214, u0_col_out_958, reg_intermediate0[958], reg_intermediate1[958]};
assign u1_col_in_1215 = {col_in_1215, u0_col_out_959, reg_intermediate0[959], reg_intermediate1[959]};
assign u1_col_in_1216 = {col_in_1216, u0_col_out_960, reg_intermediate0[960], reg_intermediate1[960]};
assign u1_col_in_1217 = {col_in_1217, u0_col_out_961, reg_intermediate0[961], reg_intermediate1[961]};
assign u1_col_in_1218 = {col_in_1218, u0_col_out_962, reg_intermediate0[962], reg_intermediate1[962]};
assign u1_col_in_1219 = {col_in_1219, u0_col_out_963, reg_intermediate0[963], reg_intermediate1[963]};
assign u1_col_in_1220 = {col_in_1220, u0_col_out_964, reg_intermediate0[964], reg_intermediate1[964]};
assign u1_col_in_1221 = {col_in_1221, u0_col_out_965, reg_intermediate0[965], reg_intermediate1[965]};
assign u1_col_in_1222 = {col_in_1222, u0_col_out_966, reg_intermediate0[966], reg_intermediate1[966]};
assign u1_col_in_1223 = {col_in_1223, u0_col_out_967, reg_intermediate0[967], reg_intermediate1[967]};
assign u1_col_in_1224 = {col_in_1224, u0_col_out_968, reg_intermediate0[968], reg_intermediate1[968]};
assign u1_col_in_1225 = {col_in_1225, u0_col_out_969, reg_intermediate0[969], reg_intermediate1[969]};
assign u1_col_in_1226 = {col_in_1226, u0_col_out_970, reg_intermediate0[970], reg_intermediate1[970]};
assign u1_col_in_1227 = {col_in_1227, u0_col_out_971, reg_intermediate0[971], reg_intermediate1[971]};
assign u1_col_in_1228 = {col_in_1228, u0_col_out_972, reg_intermediate0[972], reg_intermediate1[972]};
assign u1_col_in_1229 = {col_in_1229, u0_col_out_973, reg_intermediate0[973], reg_intermediate1[973]};
assign u1_col_in_1230 = {col_in_1230, u0_col_out_974, reg_intermediate0[974], reg_intermediate1[974]};
assign u1_col_in_1231 = {col_in_1231, u0_col_out_975, reg_intermediate0[975], reg_intermediate1[975]};
assign u1_col_in_1232 = {col_in_1232, u0_col_out_976, reg_intermediate0[976], reg_intermediate1[976]};
assign u1_col_in_1233 = {col_in_1233, u0_col_out_977, reg_intermediate0[977], reg_intermediate1[977]};
assign u1_col_in_1234 = {col_in_1234, u0_col_out_978, reg_intermediate0[978], reg_intermediate1[978]};
assign u1_col_in_1235 = {col_in_1235, u0_col_out_979, reg_intermediate0[979], reg_intermediate1[979]};
assign u1_col_in_1236 = {col_in_1236, u0_col_out_980, reg_intermediate0[980], reg_intermediate1[980]};
assign u1_col_in_1237 = {col_in_1237, u0_col_out_981, reg_intermediate0[981], reg_intermediate1[981]};
assign u1_col_in_1238 = {col_in_1238, u0_col_out_982, reg_intermediate0[982], reg_intermediate1[982]};
assign u1_col_in_1239 = {col_in_1239, u0_col_out_983, reg_intermediate0[983], reg_intermediate1[983]};
assign u1_col_in_1240 = {col_in_1240, u0_col_out_984, reg_intermediate0[984], reg_intermediate1[984]};
assign u1_col_in_1241 = {col_in_1241, u0_col_out_985, reg_intermediate0[985], reg_intermediate1[985]};
assign u1_col_in_1242 = {col_in_1242, u0_col_out_986, reg_intermediate0[986], reg_intermediate1[986]};
assign u1_col_in_1243 = {col_in_1243, u0_col_out_987, reg_intermediate0[987], reg_intermediate1[987]};
assign u1_col_in_1244 = {col_in_1244, u0_col_out_988, reg_intermediate0[988], reg_intermediate1[988]};
assign u1_col_in_1245 = {col_in_1245, u0_col_out_989, reg_intermediate0[989], reg_intermediate1[989]};
assign u1_col_in_1246 = {col_in_1246, u0_col_out_990, reg_intermediate0[990], reg_intermediate1[990]};
assign u1_col_in_1247 = {col_in_1247, u0_col_out_991, reg_intermediate0[991], reg_intermediate1[991]};
assign u1_col_in_1248 = {col_in_1248, u0_col_out_992, reg_intermediate0[992], reg_intermediate1[992]};
assign u1_col_in_1249 = {col_in_1249, u0_col_out_993, reg_intermediate0[993], reg_intermediate1[993]};
assign u1_col_in_1250 = {col_in_1250, u0_col_out_994, reg_intermediate0[994], reg_intermediate1[994]};
assign u1_col_in_1251 = {col_in_1251, u0_col_out_995, reg_intermediate0[995], reg_intermediate1[995]};
assign u1_col_in_1252 = {col_in_1252, u0_col_out_996, reg_intermediate0[996], reg_intermediate1[996]};
assign u1_col_in_1253 = {col_in_1253, u0_col_out_997, reg_intermediate0[997], reg_intermediate1[997]};
assign u1_col_in_1254 = {col_in_1254, u0_col_out_998, reg_intermediate0[998], reg_intermediate1[998]};
assign u1_col_in_1255 = {col_in_1255, u0_col_out_999, reg_intermediate0[999], reg_intermediate1[999]};
assign u1_col_in_1256 = {col_in_1256, u0_col_out_1000, reg_intermediate0[1000], reg_intermediate1[1000]};
assign u1_col_in_1257 = {col_in_1257, u0_col_out_1001, reg_intermediate0[1001], reg_intermediate1[1001]};
assign u1_col_in_1258 = {col_in_1258, u0_col_out_1002, reg_intermediate0[1002], reg_intermediate1[1002]};
assign u1_col_in_1259 = {col_in_1259, u0_col_out_1003, reg_intermediate0[1003], reg_intermediate1[1003]};
assign u1_col_in_1260 = {col_in_1260, u0_col_out_1004, reg_intermediate0[1004], reg_intermediate1[1004]};
assign u1_col_in_1261 = {col_in_1261, u0_col_out_1005, reg_intermediate0[1005], reg_intermediate1[1005]};
assign u1_col_in_1262 = {col_in_1262, u0_col_out_1006, reg_intermediate0[1006], reg_intermediate1[1006]};
assign u1_col_in_1263 = {col_in_1263, u0_col_out_1007, reg_intermediate0[1007], reg_intermediate1[1007]};
assign u1_col_in_1264 = {col_in_1264, u0_col_out_1008, reg_intermediate0[1008], reg_intermediate1[1008]};
assign u1_col_in_1265 = {col_in_1265, u0_col_out_1009, reg_intermediate0[1009], reg_intermediate1[1009]};
assign u1_col_in_1266 = {col_in_1266, u0_col_out_1010, reg_intermediate0[1010], reg_intermediate1[1010]};
assign u1_col_in_1267 = {col_in_1267, u0_col_out_1011, reg_intermediate0[1011], reg_intermediate1[1011]};
assign u1_col_in_1268 = {col_in_1268, u0_col_out_1012, reg_intermediate0[1012], reg_intermediate1[1012]};
assign u1_col_in_1269 = {col_in_1269, u0_col_out_1013, reg_intermediate0[1013], reg_intermediate1[1013]};
assign u1_col_in_1270 = {col_in_1270, u0_col_out_1014, reg_intermediate0[1014], reg_intermediate1[1014]};
assign u1_col_in_1271 = {col_in_1271, u0_col_out_1015, reg_intermediate0[1015], reg_intermediate1[1015]};
assign u1_col_in_1272 = {col_in_1272, u0_col_out_1016, reg_intermediate0[1016], reg_intermediate1[1016]};
assign u1_col_in_1273 = {col_in_1273, u0_col_out_1017, reg_intermediate0[1017], reg_intermediate1[1017]};
assign u1_col_in_1274 = {col_in_1274, u0_col_out_1018, reg_intermediate0[1018], reg_intermediate1[1018]};
assign u1_col_in_1275 = {col_in_1275, u0_col_out_1019, reg_intermediate0[1019], reg_intermediate1[1019]};
assign u1_col_in_1276 = {col_in_1276, u0_col_out_1020, reg_intermediate0[1020], reg_intermediate1[1020]};
assign u1_col_in_1277 = {col_in_1277, u0_col_out_1021, reg_intermediate0[1021], reg_intermediate1[1021]};
assign u1_col_in_1278 = {col_in_1278, u0_col_out_1022, reg_intermediate0[1022], reg_intermediate1[1022]};
assign u1_col_in_1279 = {col_in_1279, u0_col_out_1023, reg_intermediate0[1023], reg_intermediate1[1023]};


compressor_array_236_2_1280_row u1_compressor_array_236_2_1280_row
(
    .col_in_0(u1_col_in_0),
    .col_in_1(u1_col_in_1),
    .col_in_2(u1_col_in_2),
    .col_in_3(u1_col_in_3),
    .col_in_4(u1_col_in_4),
    .col_in_5(u1_col_in_5),
    .col_in_6(u1_col_in_6),
    .col_in_7(u1_col_in_7),
    .col_in_8(u1_col_in_8),
    .col_in_9(u1_col_in_9),
    .col_in_10(u1_col_in_10),
    .col_in_11(u1_col_in_11),
    .col_in_12(u1_col_in_12),
    .col_in_13(u1_col_in_13),
    .col_in_14(u1_col_in_14),
    .col_in_15(u1_col_in_15),
    .col_in_16(u1_col_in_16),
    .col_in_17(u1_col_in_17),
    .col_in_18(u1_col_in_18),
    .col_in_19(u1_col_in_19),
    .col_in_20(u1_col_in_20),
    .col_in_21(u1_col_in_21),
    .col_in_22(u1_col_in_22),
    .col_in_23(u1_col_in_23),
    .col_in_24(u1_col_in_24),
    .col_in_25(u1_col_in_25),
    .col_in_26(u1_col_in_26),
    .col_in_27(u1_col_in_27),
    .col_in_28(u1_col_in_28),
    .col_in_29(u1_col_in_29),
    .col_in_30(u1_col_in_30),
    .col_in_31(u1_col_in_31),
    .col_in_32(u1_col_in_32),
    .col_in_33(u1_col_in_33),
    .col_in_34(u1_col_in_34),
    .col_in_35(u1_col_in_35),
    .col_in_36(u1_col_in_36),
    .col_in_37(u1_col_in_37),
    .col_in_38(u1_col_in_38),
    .col_in_39(u1_col_in_39),
    .col_in_40(u1_col_in_40),
    .col_in_41(u1_col_in_41),
    .col_in_42(u1_col_in_42),
    .col_in_43(u1_col_in_43),
    .col_in_44(u1_col_in_44),
    .col_in_45(u1_col_in_45),
    .col_in_46(u1_col_in_46),
    .col_in_47(u1_col_in_47),
    .col_in_48(u1_col_in_48),
    .col_in_49(u1_col_in_49),
    .col_in_50(u1_col_in_50),
    .col_in_51(u1_col_in_51),
    .col_in_52(u1_col_in_52),
    .col_in_53(u1_col_in_53),
    .col_in_54(u1_col_in_54),
    .col_in_55(u1_col_in_55),
    .col_in_56(u1_col_in_56),
    .col_in_57(u1_col_in_57),
    .col_in_58(u1_col_in_58),
    .col_in_59(u1_col_in_59),
    .col_in_60(u1_col_in_60),
    .col_in_61(u1_col_in_61),
    .col_in_62(u1_col_in_62),
    .col_in_63(u1_col_in_63),
    .col_in_64(u1_col_in_64),
    .col_in_65(u1_col_in_65),
    .col_in_66(u1_col_in_66),
    .col_in_67(u1_col_in_67),
    .col_in_68(u1_col_in_68),
    .col_in_69(u1_col_in_69),
    .col_in_70(u1_col_in_70),
    .col_in_71(u1_col_in_71),
    .col_in_72(u1_col_in_72),
    .col_in_73(u1_col_in_73),
    .col_in_74(u1_col_in_74),
    .col_in_75(u1_col_in_75),
    .col_in_76(u1_col_in_76),
    .col_in_77(u1_col_in_77),
    .col_in_78(u1_col_in_78),
    .col_in_79(u1_col_in_79),
    .col_in_80(u1_col_in_80),
    .col_in_81(u1_col_in_81),
    .col_in_82(u1_col_in_82),
    .col_in_83(u1_col_in_83),
    .col_in_84(u1_col_in_84),
    .col_in_85(u1_col_in_85),
    .col_in_86(u1_col_in_86),
    .col_in_87(u1_col_in_87),
    .col_in_88(u1_col_in_88),
    .col_in_89(u1_col_in_89),
    .col_in_90(u1_col_in_90),
    .col_in_91(u1_col_in_91),
    .col_in_92(u1_col_in_92),
    .col_in_93(u1_col_in_93),
    .col_in_94(u1_col_in_94),
    .col_in_95(u1_col_in_95),
    .col_in_96(u1_col_in_96),
    .col_in_97(u1_col_in_97),
    .col_in_98(u1_col_in_98),
    .col_in_99(u1_col_in_99),
    .col_in_100(u1_col_in_100),
    .col_in_101(u1_col_in_101),
    .col_in_102(u1_col_in_102),
    .col_in_103(u1_col_in_103),
    .col_in_104(u1_col_in_104),
    .col_in_105(u1_col_in_105),
    .col_in_106(u1_col_in_106),
    .col_in_107(u1_col_in_107),
    .col_in_108(u1_col_in_108),
    .col_in_109(u1_col_in_109),
    .col_in_110(u1_col_in_110),
    .col_in_111(u1_col_in_111),
    .col_in_112(u1_col_in_112),
    .col_in_113(u1_col_in_113),
    .col_in_114(u1_col_in_114),
    .col_in_115(u1_col_in_115),
    .col_in_116(u1_col_in_116),
    .col_in_117(u1_col_in_117),
    .col_in_118(u1_col_in_118),
    .col_in_119(u1_col_in_119),
    .col_in_120(u1_col_in_120),
    .col_in_121(u1_col_in_121),
    .col_in_122(u1_col_in_122),
    .col_in_123(u1_col_in_123),
    .col_in_124(u1_col_in_124),
    .col_in_125(u1_col_in_125),
    .col_in_126(u1_col_in_126),
    .col_in_127(u1_col_in_127),
    .col_in_128(u1_col_in_128),
    .col_in_129(u1_col_in_129),
    .col_in_130(u1_col_in_130),
    .col_in_131(u1_col_in_131),
    .col_in_132(u1_col_in_132),
    .col_in_133(u1_col_in_133),
    .col_in_134(u1_col_in_134),
    .col_in_135(u1_col_in_135),
    .col_in_136(u1_col_in_136),
    .col_in_137(u1_col_in_137),
    .col_in_138(u1_col_in_138),
    .col_in_139(u1_col_in_139),
    .col_in_140(u1_col_in_140),
    .col_in_141(u1_col_in_141),
    .col_in_142(u1_col_in_142),
    .col_in_143(u1_col_in_143),
    .col_in_144(u1_col_in_144),
    .col_in_145(u1_col_in_145),
    .col_in_146(u1_col_in_146),
    .col_in_147(u1_col_in_147),
    .col_in_148(u1_col_in_148),
    .col_in_149(u1_col_in_149),
    .col_in_150(u1_col_in_150),
    .col_in_151(u1_col_in_151),
    .col_in_152(u1_col_in_152),
    .col_in_153(u1_col_in_153),
    .col_in_154(u1_col_in_154),
    .col_in_155(u1_col_in_155),
    .col_in_156(u1_col_in_156),
    .col_in_157(u1_col_in_157),
    .col_in_158(u1_col_in_158),
    .col_in_159(u1_col_in_159),
    .col_in_160(u1_col_in_160),
    .col_in_161(u1_col_in_161),
    .col_in_162(u1_col_in_162),
    .col_in_163(u1_col_in_163),
    .col_in_164(u1_col_in_164),
    .col_in_165(u1_col_in_165),
    .col_in_166(u1_col_in_166),
    .col_in_167(u1_col_in_167),
    .col_in_168(u1_col_in_168),
    .col_in_169(u1_col_in_169),
    .col_in_170(u1_col_in_170),
    .col_in_171(u1_col_in_171),
    .col_in_172(u1_col_in_172),
    .col_in_173(u1_col_in_173),
    .col_in_174(u1_col_in_174),
    .col_in_175(u1_col_in_175),
    .col_in_176(u1_col_in_176),
    .col_in_177(u1_col_in_177),
    .col_in_178(u1_col_in_178),
    .col_in_179(u1_col_in_179),
    .col_in_180(u1_col_in_180),
    .col_in_181(u1_col_in_181),
    .col_in_182(u1_col_in_182),
    .col_in_183(u1_col_in_183),
    .col_in_184(u1_col_in_184),
    .col_in_185(u1_col_in_185),
    .col_in_186(u1_col_in_186),
    .col_in_187(u1_col_in_187),
    .col_in_188(u1_col_in_188),
    .col_in_189(u1_col_in_189),
    .col_in_190(u1_col_in_190),
    .col_in_191(u1_col_in_191),
    .col_in_192(u1_col_in_192),
    .col_in_193(u1_col_in_193),
    .col_in_194(u1_col_in_194),
    .col_in_195(u1_col_in_195),
    .col_in_196(u1_col_in_196),
    .col_in_197(u1_col_in_197),
    .col_in_198(u1_col_in_198),
    .col_in_199(u1_col_in_199),
    .col_in_200(u1_col_in_200),
    .col_in_201(u1_col_in_201),
    .col_in_202(u1_col_in_202),
    .col_in_203(u1_col_in_203),
    .col_in_204(u1_col_in_204),
    .col_in_205(u1_col_in_205),
    .col_in_206(u1_col_in_206),
    .col_in_207(u1_col_in_207),
    .col_in_208(u1_col_in_208),
    .col_in_209(u1_col_in_209),
    .col_in_210(u1_col_in_210),
    .col_in_211(u1_col_in_211),
    .col_in_212(u1_col_in_212),
    .col_in_213(u1_col_in_213),
    .col_in_214(u1_col_in_214),
    .col_in_215(u1_col_in_215),
    .col_in_216(u1_col_in_216),
    .col_in_217(u1_col_in_217),
    .col_in_218(u1_col_in_218),
    .col_in_219(u1_col_in_219),
    .col_in_220(u1_col_in_220),
    .col_in_221(u1_col_in_221),
    .col_in_222(u1_col_in_222),
    .col_in_223(u1_col_in_223),
    .col_in_224(u1_col_in_224),
    .col_in_225(u1_col_in_225),
    .col_in_226(u1_col_in_226),
    .col_in_227(u1_col_in_227),
    .col_in_228(u1_col_in_228),
    .col_in_229(u1_col_in_229),
    .col_in_230(u1_col_in_230),
    .col_in_231(u1_col_in_231),
    .col_in_232(u1_col_in_232),
    .col_in_233(u1_col_in_233),
    .col_in_234(u1_col_in_234),
    .col_in_235(u1_col_in_235),
    .col_in_236(u1_col_in_236),
    .col_in_237(u1_col_in_237),
    .col_in_238(u1_col_in_238),
    .col_in_239(u1_col_in_239),
    .col_in_240(u1_col_in_240),
    .col_in_241(u1_col_in_241),
    .col_in_242(u1_col_in_242),
    .col_in_243(u1_col_in_243),
    .col_in_244(u1_col_in_244),
    .col_in_245(u1_col_in_245),
    .col_in_246(u1_col_in_246),
    .col_in_247(u1_col_in_247),
    .col_in_248(u1_col_in_248),
    .col_in_249(u1_col_in_249),
    .col_in_250(u1_col_in_250),
    .col_in_251(u1_col_in_251),
    .col_in_252(u1_col_in_252),
    .col_in_253(u1_col_in_253),
    .col_in_254(u1_col_in_254),
    .col_in_255(u1_col_in_255),
    .col_in_256(u1_col_in_256),
    .col_in_257(u1_col_in_257),
    .col_in_258(u1_col_in_258),
    .col_in_259(u1_col_in_259),
    .col_in_260(u1_col_in_260),
    .col_in_261(u1_col_in_261),
    .col_in_262(u1_col_in_262),
    .col_in_263(u1_col_in_263),
    .col_in_264(u1_col_in_264),
    .col_in_265(u1_col_in_265),
    .col_in_266(u1_col_in_266),
    .col_in_267(u1_col_in_267),
    .col_in_268(u1_col_in_268),
    .col_in_269(u1_col_in_269),
    .col_in_270(u1_col_in_270),
    .col_in_271(u1_col_in_271),
    .col_in_272(u1_col_in_272),
    .col_in_273(u1_col_in_273),
    .col_in_274(u1_col_in_274),
    .col_in_275(u1_col_in_275),
    .col_in_276(u1_col_in_276),
    .col_in_277(u1_col_in_277),
    .col_in_278(u1_col_in_278),
    .col_in_279(u1_col_in_279),
    .col_in_280(u1_col_in_280),
    .col_in_281(u1_col_in_281),
    .col_in_282(u1_col_in_282),
    .col_in_283(u1_col_in_283),
    .col_in_284(u1_col_in_284),
    .col_in_285(u1_col_in_285),
    .col_in_286(u1_col_in_286),
    .col_in_287(u1_col_in_287),
    .col_in_288(u1_col_in_288),
    .col_in_289(u1_col_in_289),
    .col_in_290(u1_col_in_290),
    .col_in_291(u1_col_in_291),
    .col_in_292(u1_col_in_292),
    .col_in_293(u1_col_in_293),
    .col_in_294(u1_col_in_294),
    .col_in_295(u1_col_in_295),
    .col_in_296(u1_col_in_296),
    .col_in_297(u1_col_in_297),
    .col_in_298(u1_col_in_298),
    .col_in_299(u1_col_in_299),
    .col_in_300(u1_col_in_300),
    .col_in_301(u1_col_in_301),
    .col_in_302(u1_col_in_302),
    .col_in_303(u1_col_in_303),
    .col_in_304(u1_col_in_304),
    .col_in_305(u1_col_in_305),
    .col_in_306(u1_col_in_306),
    .col_in_307(u1_col_in_307),
    .col_in_308(u1_col_in_308),
    .col_in_309(u1_col_in_309),
    .col_in_310(u1_col_in_310),
    .col_in_311(u1_col_in_311),
    .col_in_312(u1_col_in_312),
    .col_in_313(u1_col_in_313),
    .col_in_314(u1_col_in_314),
    .col_in_315(u1_col_in_315),
    .col_in_316(u1_col_in_316),
    .col_in_317(u1_col_in_317),
    .col_in_318(u1_col_in_318),
    .col_in_319(u1_col_in_319),
    .col_in_320(u1_col_in_320),
    .col_in_321(u1_col_in_321),
    .col_in_322(u1_col_in_322),
    .col_in_323(u1_col_in_323),
    .col_in_324(u1_col_in_324),
    .col_in_325(u1_col_in_325),
    .col_in_326(u1_col_in_326),
    .col_in_327(u1_col_in_327),
    .col_in_328(u1_col_in_328),
    .col_in_329(u1_col_in_329),
    .col_in_330(u1_col_in_330),
    .col_in_331(u1_col_in_331),
    .col_in_332(u1_col_in_332),
    .col_in_333(u1_col_in_333),
    .col_in_334(u1_col_in_334),
    .col_in_335(u1_col_in_335),
    .col_in_336(u1_col_in_336),
    .col_in_337(u1_col_in_337),
    .col_in_338(u1_col_in_338),
    .col_in_339(u1_col_in_339),
    .col_in_340(u1_col_in_340),
    .col_in_341(u1_col_in_341),
    .col_in_342(u1_col_in_342),
    .col_in_343(u1_col_in_343),
    .col_in_344(u1_col_in_344),
    .col_in_345(u1_col_in_345),
    .col_in_346(u1_col_in_346),
    .col_in_347(u1_col_in_347),
    .col_in_348(u1_col_in_348),
    .col_in_349(u1_col_in_349),
    .col_in_350(u1_col_in_350),
    .col_in_351(u1_col_in_351),
    .col_in_352(u1_col_in_352),
    .col_in_353(u1_col_in_353),
    .col_in_354(u1_col_in_354),
    .col_in_355(u1_col_in_355),
    .col_in_356(u1_col_in_356),
    .col_in_357(u1_col_in_357),
    .col_in_358(u1_col_in_358),
    .col_in_359(u1_col_in_359),
    .col_in_360(u1_col_in_360),
    .col_in_361(u1_col_in_361),
    .col_in_362(u1_col_in_362),
    .col_in_363(u1_col_in_363),
    .col_in_364(u1_col_in_364),
    .col_in_365(u1_col_in_365),
    .col_in_366(u1_col_in_366),
    .col_in_367(u1_col_in_367),
    .col_in_368(u1_col_in_368),
    .col_in_369(u1_col_in_369),
    .col_in_370(u1_col_in_370),
    .col_in_371(u1_col_in_371),
    .col_in_372(u1_col_in_372),
    .col_in_373(u1_col_in_373),
    .col_in_374(u1_col_in_374),
    .col_in_375(u1_col_in_375),
    .col_in_376(u1_col_in_376),
    .col_in_377(u1_col_in_377),
    .col_in_378(u1_col_in_378),
    .col_in_379(u1_col_in_379),
    .col_in_380(u1_col_in_380),
    .col_in_381(u1_col_in_381),
    .col_in_382(u1_col_in_382),
    .col_in_383(u1_col_in_383),
    .col_in_384(u1_col_in_384),
    .col_in_385(u1_col_in_385),
    .col_in_386(u1_col_in_386),
    .col_in_387(u1_col_in_387),
    .col_in_388(u1_col_in_388),
    .col_in_389(u1_col_in_389),
    .col_in_390(u1_col_in_390),
    .col_in_391(u1_col_in_391),
    .col_in_392(u1_col_in_392),
    .col_in_393(u1_col_in_393),
    .col_in_394(u1_col_in_394),
    .col_in_395(u1_col_in_395),
    .col_in_396(u1_col_in_396),
    .col_in_397(u1_col_in_397),
    .col_in_398(u1_col_in_398),
    .col_in_399(u1_col_in_399),
    .col_in_400(u1_col_in_400),
    .col_in_401(u1_col_in_401),
    .col_in_402(u1_col_in_402),
    .col_in_403(u1_col_in_403),
    .col_in_404(u1_col_in_404),
    .col_in_405(u1_col_in_405),
    .col_in_406(u1_col_in_406),
    .col_in_407(u1_col_in_407),
    .col_in_408(u1_col_in_408),
    .col_in_409(u1_col_in_409),
    .col_in_410(u1_col_in_410),
    .col_in_411(u1_col_in_411),
    .col_in_412(u1_col_in_412),
    .col_in_413(u1_col_in_413),
    .col_in_414(u1_col_in_414),
    .col_in_415(u1_col_in_415),
    .col_in_416(u1_col_in_416),
    .col_in_417(u1_col_in_417),
    .col_in_418(u1_col_in_418),
    .col_in_419(u1_col_in_419),
    .col_in_420(u1_col_in_420),
    .col_in_421(u1_col_in_421),
    .col_in_422(u1_col_in_422),
    .col_in_423(u1_col_in_423),
    .col_in_424(u1_col_in_424),
    .col_in_425(u1_col_in_425),
    .col_in_426(u1_col_in_426),
    .col_in_427(u1_col_in_427),
    .col_in_428(u1_col_in_428),
    .col_in_429(u1_col_in_429),
    .col_in_430(u1_col_in_430),
    .col_in_431(u1_col_in_431),
    .col_in_432(u1_col_in_432),
    .col_in_433(u1_col_in_433),
    .col_in_434(u1_col_in_434),
    .col_in_435(u1_col_in_435),
    .col_in_436(u1_col_in_436),
    .col_in_437(u1_col_in_437),
    .col_in_438(u1_col_in_438),
    .col_in_439(u1_col_in_439),
    .col_in_440(u1_col_in_440),
    .col_in_441(u1_col_in_441),
    .col_in_442(u1_col_in_442),
    .col_in_443(u1_col_in_443),
    .col_in_444(u1_col_in_444),
    .col_in_445(u1_col_in_445),
    .col_in_446(u1_col_in_446),
    .col_in_447(u1_col_in_447),
    .col_in_448(u1_col_in_448),
    .col_in_449(u1_col_in_449),
    .col_in_450(u1_col_in_450),
    .col_in_451(u1_col_in_451),
    .col_in_452(u1_col_in_452),
    .col_in_453(u1_col_in_453),
    .col_in_454(u1_col_in_454),
    .col_in_455(u1_col_in_455),
    .col_in_456(u1_col_in_456),
    .col_in_457(u1_col_in_457),
    .col_in_458(u1_col_in_458),
    .col_in_459(u1_col_in_459),
    .col_in_460(u1_col_in_460),
    .col_in_461(u1_col_in_461),
    .col_in_462(u1_col_in_462),
    .col_in_463(u1_col_in_463),
    .col_in_464(u1_col_in_464),
    .col_in_465(u1_col_in_465),
    .col_in_466(u1_col_in_466),
    .col_in_467(u1_col_in_467),
    .col_in_468(u1_col_in_468),
    .col_in_469(u1_col_in_469),
    .col_in_470(u1_col_in_470),
    .col_in_471(u1_col_in_471),
    .col_in_472(u1_col_in_472),
    .col_in_473(u1_col_in_473),
    .col_in_474(u1_col_in_474),
    .col_in_475(u1_col_in_475),
    .col_in_476(u1_col_in_476),
    .col_in_477(u1_col_in_477),
    .col_in_478(u1_col_in_478),
    .col_in_479(u1_col_in_479),
    .col_in_480(u1_col_in_480),
    .col_in_481(u1_col_in_481),
    .col_in_482(u1_col_in_482),
    .col_in_483(u1_col_in_483),
    .col_in_484(u1_col_in_484),
    .col_in_485(u1_col_in_485),
    .col_in_486(u1_col_in_486),
    .col_in_487(u1_col_in_487),
    .col_in_488(u1_col_in_488),
    .col_in_489(u1_col_in_489),
    .col_in_490(u1_col_in_490),
    .col_in_491(u1_col_in_491),
    .col_in_492(u1_col_in_492),
    .col_in_493(u1_col_in_493),
    .col_in_494(u1_col_in_494),
    .col_in_495(u1_col_in_495),
    .col_in_496(u1_col_in_496),
    .col_in_497(u1_col_in_497),
    .col_in_498(u1_col_in_498),
    .col_in_499(u1_col_in_499),
    .col_in_500(u1_col_in_500),
    .col_in_501(u1_col_in_501),
    .col_in_502(u1_col_in_502),
    .col_in_503(u1_col_in_503),
    .col_in_504(u1_col_in_504),
    .col_in_505(u1_col_in_505),
    .col_in_506(u1_col_in_506),
    .col_in_507(u1_col_in_507),
    .col_in_508(u1_col_in_508),
    .col_in_509(u1_col_in_509),
    .col_in_510(u1_col_in_510),
    .col_in_511(u1_col_in_511),
    .col_in_512(u1_col_in_512),
    .col_in_513(u1_col_in_513),
    .col_in_514(u1_col_in_514),
    .col_in_515(u1_col_in_515),
    .col_in_516(u1_col_in_516),
    .col_in_517(u1_col_in_517),
    .col_in_518(u1_col_in_518),
    .col_in_519(u1_col_in_519),
    .col_in_520(u1_col_in_520),
    .col_in_521(u1_col_in_521),
    .col_in_522(u1_col_in_522),
    .col_in_523(u1_col_in_523),
    .col_in_524(u1_col_in_524),
    .col_in_525(u1_col_in_525),
    .col_in_526(u1_col_in_526),
    .col_in_527(u1_col_in_527),
    .col_in_528(u1_col_in_528),
    .col_in_529(u1_col_in_529),
    .col_in_530(u1_col_in_530),
    .col_in_531(u1_col_in_531),
    .col_in_532(u1_col_in_532),
    .col_in_533(u1_col_in_533),
    .col_in_534(u1_col_in_534),
    .col_in_535(u1_col_in_535),
    .col_in_536(u1_col_in_536),
    .col_in_537(u1_col_in_537),
    .col_in_538(u1_col_in_538),
    .col_in_539(u1_col_in_539),
    .col_in_540(u1_col_in_540),
    .col_in_541(u1_col_in_541),
    .col_in_542(u1_col_in_542),
    .col_in_543(u1_col_in_543),
    .col_in_544(u1_col_in_544),
    .col_in_545(u1_col_in_545),
    .col_in_546(u1_col_in_546),
    .col_in_547(u1_col_in_547),
    .col_in_548(u1_col_in_548),
    .col_in_549(u1_col_in_549),
    .col_in_550(u1_col_in_550),
    .col_in_551(u1_col_in_551),
    .col_in_552(u1_col_in_552),
    .col_in_553(u1_col_in_553),
    .col_in_554(u1_col_in_554),
    .col_in_555(u1_col_in_555),
    .col_in_556(u1_col_in_556),
    .col_in_557(u1_col_in_557),
    .col_in_558(u1_col_in_558),
    .col_in_559(u1_col_in_559),
    .col_in_560(u1_col_in_560),
    .col_in_561(u1_col_in_561),
    .col_in_562(u1_col_in_562),
    .col_in_563(u1_col_in_563),
    .col_in_564(u1_col_in_564),
    .col_in_565(u1_col_in_565),
    .col_in_566(u1_col_in_566),
    .col_in_567(u1_col_in_567),
    .col_in_568(u1_col_in_568),
    .col_in_569(u1_col_in_569),
    .col_in_570(u1_col_in_570),
    .col_in_571(u1_col_in_571),
    .col_in_572(u1_col_in_572),
    .col_in_573(u1_col_in_573),
    .col_in_574(u1_col_in_574),
    .col_in_575(u1_col_in_575),
    .col_in_576(u1_col_in_576),
    .col_in_577(u1_col_in_577),
    .col_in_578(u1_col_in_578),
    .col_in_579(u1_col_in_579),
    .col_in_580(u1_col_in_580),
    .col_in_581(u1_col_in_581),
    .col_in_582(u1_col_in_582),
    .col_in_583(u1_col_in_583),
    .col_in_584(u1_col_in_584),
    .col_in_585(u1_col_in_585),
    .col_in_586(u1_col_in_586),
    .col_in_587(u1_col_in_587),
    .col_in_588(u1_col_in_588),
    .col_in_589(u1_col_in_589),
    .col_in_590(u1_col_in_590),
    .col_in_591(u1_col_in_591),
    .col_in_592(u1_col_in_592),
    .col_in_593(u1_col_in_593),
    .col_in_594(u1_col_in_594),
    .col_in_595(u1_col_in_595),
    .col_in_596(u1_col_in_596),
    .col_in_597(u1_col_in_597),
    .col_in_598(u1_col_in_598),
    .col_in_599(u1_col_in_599),
    .col_in_600(u1_col_in_600),
    .col_in_601(u1_col_in_601),
    .col_in_602(u1_col_in_602),
    .col_in_603(u1_col_in_603),
    .col_in_604(u1_col_in_604),
    .col_in_605(u1_col_in_605),
    .col_in_606(u1_col_in_606),
    .col_in_607(u1_col_in_607),
    .col_in_608(u1_col_in_608),
    .col_in_609(u1_col_in_609),
    .col_in_610(u1_col_in_610),
    .col_in_611(u1_col_in_611),
    .col_in_612(u1_col_in_612),
    .col_in_613(u1_col_in_613),
    .col_in_614(u1_col_in_614),
    .col_in_615(u1_col_in_615),
    .col_in_616(u1_col_in_616),
    .col_in_617(u1_col_in_617),
    .col_in_618(u1_col_in_618),
    .col_in_619(u1_col_in_619),
    .col_in_620(u1_col_in_620),
    .col_in_621(u1_col_in_621),
    .col_in_622(u1_col_in_622),
    .col_in_623(u1_col_in_623),
    .col_in_624(u1_col_in_624),
    .col_in_625(u1_col_in_625),
    .col_in_626(u1_col_in_626),
    .col_in_627(u1_col_in_627),
    .col_in_628(u1_col_in_628),
    .col_in_629(u1_col_in_629),
    .col_in_630(u1_col_in_630),
    .col_in_631(u1_col_in_631),
    .col_in_632(u1_col_in_632),
    .col_in_633(u1_col_in_633),
    .col_in_634(u1_col_in_634),
    .col_in_635(u1_col_in_635),
    .col_in_636(u1_col_in_636),
    .col_in_637(u1_col_in_637),
    .col_in_638(u1_col_in_638),
    .col_in_639(u1_col_in_639),
    .col_in_640(u1_col_in_640),
    .col_in_641(u1_col_in_641),
    .col_in_642(u1_col_in_642),
    .col_in_643(u1_col_in_643),
    .col_in_644(u1_col_in_644),
    .col_in_645(u1_col_in_645),
    .col_in_646(u1_col_in_646),
    .col_in_647(u1_col_in_647),
    .col_in_648(u1_col_in_648),
    .col_in_649(u1_col_in_649),
    .col_in_650(u1_col_in_650),
    .col_in_651(u1_col_in_651),
    .col_in_652(u1_col_in_652),
    .col_in_653(u1_col_in_653),
    .col_in_654(u1_col_in_654),
    .col_in_655(u1_col_in_655),
    .col_in_656(u1_col_in_656),
    .col_in_657(u1_col_in_657),
    .col_in_658(u1_col_in_658),
    .col_in_659(u1_col_in_659),
    .col_in_660(u1_col_in_660),
    .col_in_661(u1_col_in_661),
    .col_in_662(u1_col_in_662),
    .col_in_663(u1_col_in_663),
    .col_in_664(u1_col_in_664),
    .col_in_665(u1_col_in_665),
    .col_in_666(u1_col_in_666),
    .col_in_667(u1_col_in_667),
    .col_in_668(u1_col_in_668),
    .col_in_669(u1_col_in_669),
    .col_in_670(u1_col_in_670),
    .col_in_671(u1_col_in_671),
    .col_in_672(u1_col_in_672),
    .col_in_673(u1_col_in_673),
    .col_in_674(u1_col_in_674),
    .col_in_675(u1_col_in_675),
    .col_in_676(u1_col_in_676),
    .col_in_677(u1_col_in_677),
    .col_in_678(u1_col_in_678),
    .col_in_679(u1_col_in_679),
    .col_in_680(u1_col_in_680),
    .col_in_681(u1_col_in_681),
    .col_in_682(u1_col_in_682),
    .col_in_683(u1_col_in_683),
    .col_in_684(u1_col_in_684),
    .col_in_685(u1_col_in_685),
    .col_in_686(u1_col_in_686),
    .col_in_687(u1_col_in_687),
    .col_in_688(u1_col_in_688),
    .col_in_689(u1_col_in_689),
    .col_in_690(u1_col_in_690),
    .col_in_691(u1_col_in_691),
    .col_in_692(u1_col_in_692),
    .col_in_693(u1_col_in_693),
    .col_in_694(u1_col_in_694),
    .col_in_695(u1_col_in_695),
    .col_in_696(u1_col_in_696),
    .col_in_697(u1_col_in_697),
    .col_in_698(u1_col_in_698),
    .col_in_699(u1_col_in_699),
    .col_in_700(u1_col_in_700),
    .col_in_701(u1_col_in_701),
    .col_in_702(u1_col_in_702),
    .col_in_703(u1_col_in_703),
    .col_in_704(u1_col_in_704),
    .col_in_705(u1_col_in_705),
    .col_in_706(u1_col_in_706),
    .col_in_707(u1_col_in_707),
    .col_in_708(u1_col_in_708),
    .col_in_709(u1_col_in_709),
    .col_in_710(u1_col_in_710),
    .col_in_711(u1_col_in_711),
    .col_in_712(u1_col_in_712),
    .col_in_713(u1_col_in_713),
    .col_in_714(u1_col_in_714),
    .col_in_715(u1_col_in_715),
    .col_in_716(u1_col_in_716),
    .col_in_717(u1_col_in_717),
    .col_in_718(u1_col_in_718),
    .col_in_719(u1_col_in_719),
    .col_in_720(u1_col_in_720),
    .col_in_721(u1_col_in_721),
    .col_in_722(u1_col_in_722),
    .col_in_723(u1_col_in_723),
    .col_in_724(u1_col_in_724),
    .col_in_725(u1_col_in_725),
    .col_in_726(u1_col_in_726),
    .col_in_727(u1_col_in_727),
    .col_in_728(u1_col_in_728),
    .col_in_729(u1_col_in_729),
    .col_in_730(u1_col_in_730),
    .col_in_731(u1_col_in_731),
    .col_in_732(u1_col_in_732),
    .col_in_733(u1_col_in_733),
    .col_in_734(u1_col_in_734),
    .col_in_735(u1_col_in_735),
    .col_in_736(u1_col_in_736),
    .col_in_737(u1_col_in_737),
    .col_in_738(u1_col_in_738),
    .col_in_739(u1_col_in_739),
    .col_in_740(u1_col_in_740),
    .col_in_741(u1_col_in_741),
    .col_in_742(u1_col_in_742),
    .col_in_743(u1_col_in_743),
    .col_in_744(u1_col_in_744),
    .col_in_745(u1_col_in_745),
    .col_in_746(u1_col_in_746),
    .col_in_747(u1_col_in_747),
    .col_in_748(u1_col_in_748),
    .col_in_749(u1_col_in_749),
    .col_in_750(u1_col_in_750),
    .col_in_751(u1_col_in_751),
    .col_in_752(u1_col_in_752),
    .col_in_753(u1_col_in_753),
    .col_in_754(u1_col_in_754),
    .col_in_755(u1_col_in_755),
    .col_in_756(u1_col_in_756),
    .col_in_757(u1_col_in_757),
    .col_in_758(u1_col_in_758),
    .col_in_759(u1_col_in_759),
    .col_in_760(u1_col_in_760),
    .col_in_761(u1_col_in_761),
    .col_in_762(u1_col_in_762),
    .col_in_763(u1_col_in_763),
    .col_in_764(u1_col_in_764),
    .col_in_765(u1_col_in_765),
    .col_in_766(u1_col_in_766),
    .col_in_767(u1_col_in_767),
    .col_in_768(u1_col_in_768),
    .col_in_769(u1_col_in_769),
    .col_in_770(u1_col_in_770),
    .col_in_771(u1_col_in_771),
    .col_in_772(u1_col_in_772),
    .col_in_773(u1_col_in_773),
    .col_in_774(u1_col_in_774),
    .col_in_775(u1_col_in_775),
    .col_in_776(u1_col_in_776),
    .col_in_777(u1_col_in_777),
    .col_in_778(u1_col_in_778),
    .col_in_779(u1_col_in_779),
    .col_in_780(u1_col_in_780),
    .col_in_781(u1_col_in_781),
    .col_in_782(u1_col_in_782),
    .col_in_783(u1_col_in_783),
    .col_in_784(u1_col_in_784),
    .col_in_785(u1_col_in_785),
    .col_in_786(u1_col_in_786),
    .col_in_787(u1_col_in_787),
    .col_in_788(u1_col_in_788),
    .col_in_789(u1_col_in_789),
    .col_in_790(u1_col_in_790),
    .col_in_791(u1_col_in_791),
    .col_in_792(u1_col_in_792),
    .col_in_793(u1_col_in_793),
    .col_in_794(u1_col_in_794),
    .col_in_795(u1_col_in_795),
    .col_in_796(u1_col_in_796),
    .col_in_797(u1_col_in_797),
    .col_in_798(u1_col_in_798),
    .col_in_799(u1_col_in_799),
    .col_in_800(u1_col_in_800),
    .col_in_801(u1_col_in_801),
    .col_in_802(u1_col_in_802),
    .col_in_803(u1_col_in_803),
    .col_in_804(u1_col_in_804),
    .col_in_805(u1_col_in_805),
    .col_in_806(u1_col_in_806),
    .col_in_807(u1_col_in_807),
    .col_in_808(u1_col_in_808),
    .col_in_809(u1_col_in_809),
    .col_in_810(u1_col_in_810),
    .col_in_811(u1_col_in_811),
    .col_in_812(u1_col_in_812),
    .col_in_813(u1_col_in_813),
    .col_in_814(u1_col_in_814),
    .col_in_815(u1_col_in_815),
    .col_in_816(u1_col_in_816),
    .col_in_817(u1_col_in_817),
    .col_in_818(u1_col_in_818),
    .col_in_819(u1_col_in_819),
    .col_in_820(u1_col_in_820),
    .col_in_821(u1_col_in_821),
    .col_in_822(u1_col_in_822),
    .col_in_823(u1_col_in_823),
    .col_in_824(u1_col_in_824),
    .col_in_825(u1_col_in_825),
    .col_in_826(u1_col_in_826),
    .col_in_827(u1_col_in_827),
    .col_in_828(u1_col_in_828),
    .col_in_829(u1_col_in_829),
    .col_in_830(u1_col_in_830),
    .col_in_831(u1_col_in_831),
    .col_in_832(u1_col_in_832),
    .col_in_833(u1_col_in_833),
    .col_in_834(u1_col_in_834),
    .col_in_835(u1_col_in_835),
    .col_in_836(u1_col_in_836),
    .col_in_837(u1_col_in_837),
    .col_in_838(u1_col_in_838),
    .col_in_839(u1_col_in_839),
    .col_in_840(u1_col_in_840),
    .col_in_841(u1_col_in_841),
    .col_in_842(u1_col_in_842),
    .col_in_843(u1_col_in_843),
    .col_in_844(u1_col_in_844),
    .col_in_845(u1_col_in_845),
    .col_in_846(u1_col_in_846),
    .col_in_847(u1_col_in_847),
    .col_in_848(u1_col_in_848),
    .col_in_849(u1_col_in_849),
    .col_in_850(u1_col_in_850),
    .col_in_851(u1_col_in_851),
    .col_in_852(u1_col_in_852),
    .col_in_853(u1_col_in_853),
    .col_in_854(u1_col_in_854),
    .col_in_855(u1_col_in_855),
    .col_in_856(u1_col_in_856),
    .col_in_857(u1_col_in_857),
    .col_in_858(u1_col_in_858),
    .col_in_859(u1_col_in_859),
    .col_in_860(u1_col_in_860),
    .col_in_861(u1_col_in_861),
    .col_in_862(u1_col_in_862),
    .col_in_863(u1_col_in_863),
    .col_in_864(u1_col_in_864),
    .col_in_865(u1_col_in_865),
    .col_in_866(u1_col_in_866),
    .col_in_867(u1_col_in_867),
    .col_in_868(u1_col_in_868),
    .col_in_869(u1_col_in_869),
    .col_in_870(u1_col_in_870),
    .col_in_871(u1_col_in_871),
    .col_in_872(u1_col_in_872),
    .col_in_873(u1_col_in_873),
    .col_in_874(u1_col_in_874),
    .col_in_875(u1_col_in_875),
    .col_in_876(u1_col_in_876),
    .col_in_877(u1_col_in_877),
    .col_in_878(u1_col_in_878),
    .col_in_879(u1_col_in_879),
    .col_in_880(u1_col_in_880),
    .col_in_881(u1_col_in_881),
    .col_in_882(u1_col_in_882),
    .col_in_883(u1_col_in_883),
    .col_in_884(u1_col_in_884),
    .col_in_885(u1_col_in_885),
    .col_in_886(u1_col_in_886),
    .col_in_887(u1_col_in_887),
    .col_in_888(u1_col_in_888),
    .col_in_889(u1_col_in_889),
    .col_in_890(u1_col_in_890),
    .col_in_891(u1_col_in_891),
    .col_in_892(u1_col_in_892),
    .col_in_893(u1_col_in_893),
    .col_in_894(u1_col_in_894),
    .col_in_895(u1_col_in_895),
    .col_in_896(u1_col_in_896),
    .col_in_897(u1_col_in_897),
    .col_in_898(u1_col_in_898),
    .col_in_899(u1_col_in_899),
    .col_in_900(u1_col_in_900),
    .col_in_901(u1_col_in_901),
    .col_in_902(u1_col_in_902),
    .col_in_903(u1_col_in_903),
    .col_in_904(u1_col_in_904),
    .col_in_905(u1_col_in_905),
    .col_in_906(u1_col_in_906),
    .col_in_907(u1_col_in_907),
    .col_in_908(u1_col_in_908),
    .col_in_909(u1_col_in_909),
    .col_in_910(u1_col_in_910),
    .col_in_911(u1_col_in_911),
    .col_in_912(u1_col_in_912),
    .col_in_913(u1_col_in_913),
    .col_in_914(u1_col_in_914),
    .col_in_915(u1_col_in_915),
    .col_in_916(u1_col_in_916),
    .col_in_917(u1_col_in_917),
    .col_in_918(u1_col_in_918),
    .col_in_919(u1_col_in_919),
    .col_in_920(u1_col_in_920),
    .col_in_921(u1_col_in_921),
    .col_in_922(u1_col_in_922),
    .col_in_923(u1_col_in_923),
    .col_in_924(u1_col_in_924),
    .col_in_925(u1_col_in_925),
    .col_in_926(u1_col_in_926),
    .col_in_927(u1_col_in_927),
    .col_in_928(u1_col_in_928),
    .col_in_929(u1_col_in_929),
    .col_in_930(u1_col_in_930),
    .col_in_931(u1_col_in_931),
    .col_in_932(u1_col_in_932),
    .col_in_933(u1_col_in_933),
    .col_in_934(u1_col_in_934),
    .col_in_935(u1_col_in_935),
    .col_in_936(u1_col_in_936),
    .col_in_937(u1_col_in_937),
    .col_in_938(u1_col_in_938),
    .col_in_939(u1_col_in_939),
    .col_in_940(u1_col_in_940),
    .col_in_941(u1_col_in_941),
    .col_in_942(u1_col_in_942),
    .col_in_943(u1_col_in_943),
    .col_in_944(u1_col_in_944),
    .col_in_945(u1_col_in_945),
    .col_in_946(u1_col_in_946),
    .col_in_947(u1_col_in_947),
    .col_in_948(u1_col_in_948),
    .col_in_949(u1_col_in_949),
    .col_in_950(u1_col_in_950),
    .col_in_951(u1_col_in_951),
    .col_in_952(u1_col_in_952),
    .col_in_953(u1_col_in_953),
    .col_in_954(u1_col_in_954),
    .col_in_955(u1_col_in_955),
    .col_in_956(u1_col_in_956),
    .col_in_957(u1_col_in_957),
    .col_in_958(u1_col_in_958),
    .col_in_959(u1_col_in_959),
    .col_in_960(u1_col_in_960),
    .col_in_961(u1_col_in_961),
    .col_in_962(u1_col_in_962),
    .col_in_963(u1_col_in_963),
    .col_in_964(u1_col_in_964),
    .col_in_965(u1_col_in_965),
    .col_in_966(u1_col_in_966),
    .col_in_967(u1_col_in_967),
    .col_in_968(u1_col_in_968),
    .col_in_969(u1_col_in_969),
    .col_in_970(u1_col_in_970),
    .col_in_971(u1_col_in_971),
    .col_in_972(u1_col_in_972),
    .col_in_973(u1_col_in_973),
    .col_in_974(u1_col_in_974),
    .col_in_975(u1_col_in_975),
    .col_in_976(u1_col_in_976),
    .col_in_977(u1_col_in_977),
    .col_in_978(u1_col_in_978),
    .col_in_979(u1_col_in_979),
    .col_in_980(u1_col_in_980),
    .col_in_981(u1_col_in_981),
    .col_in_982(u1_col_in_982),
    .col_in_983(u1_col_in_983),
    .col_in_984(u1_col_in_984),
    .col_in_985(u1_col_in_985),
    .col_in_986(u1_col_in_986),
    .col_in_987(u1_col_in_987),
    .col_in_988(u1_col_in_988),
    .col_in_989(u1_col_in_989),
    .col_in_990(u1_col_in_990),
    .col_in_991(u1_col_in_991),
    .col_in_992(u1_col_in_992),
    .col_in_993(u1_col_in_993),
    .col_in_994(u1_col_in_994),
    .col_in_995(u1_col_in_995),
    .col_in_996(u1_col_in_996),
    .col_in_997(u1_col_in_997),
    .col_in_998(u1_col_in_998),
    .col_in_999(u1_col_in_999),
    .col_in_1000(u1_col_in_1000),
    .col_in_1001(u1_col_in_1001),
    .col_in_1002(u1_col_in_1002),
    .col_in_1003(u1_col_in_1003),
    .col_in_1004(u1_col_in_1004),
    .col_in_1005(u1_col_in_1005),
    .col_in_1006(u1_col_in_1006),
    .col_in_1007(u1_col_in_1007),
    .col_in_1008(u1_col_in_1008),
    .col_in_1009(u1_col_in_1009),
    .col_in_1010(u1_col_in_1010),
    .col_in_1011(u1_col_in_1011),
    .col_in_1012(u1_col_in_1012),
    .col_in_1013(u1_col_in_1013),
    .col_in_1014(u1_col_in_1014),
    .col_in_1015(u1_col_in_1015),
    .col_in_1016(u1_col_in_1016),
    .col_in_1017(u1_col_in_1017),
    .col_in_1018(u1_col_in_1018),
    .col_in_1019(u1_col_in_1019),
    .col_in_1020(u1_col_in_1020),
    .col_in_1021(u1_col_in_1021),
    .col_in_1022(u1_col_in_1022),
    .col_in_1023(u1_col_in_1023),
    .col_in_1024(u1_col_in_1024),
    .col_in_1025(u1_col_in_1025),
    .col_in_1026(u1_col_in_1026),
    .col_in_1027(u1_col_in_1027),
    .col_in_1028(u1_col_in_1028),
    .col_in_1029(u1_col_in_1029),
    .col_in_1030(u1_col_in_1030),
    .col_in_1031(u1_col_in_1031),
    .col_in_1032(u1_col_in_1032),
    .col_in_1033(u1_col_in_1033),
    .col_in_1034(u1_col_in_1034),
    .col_in_1035(u1_col_in_1035),
    .col_in_1036(u1_col_in_1036),
    .col_in_1037(u1_col_in_1037),
    .col_in_1038(u1_col_in_1038),
    .col_in_1039(u1_col_in_1039),
    .col_in_1040(u1_col_in_1040),
    .col_in_1041(u1_col_in_1041),
    .col_in_1042(u1_col_in_1042),
    .col_in_1043(u1_col_in_1043),
    .col_in_1044(u1_col_in_1044),
    .col_in_1045(u1_col_in_1045),
    .col_in_1046(u1_col_in_1046),
    .col_in_1047(u1_col_in_1047),
    .col_in_1048(u1_col_in_1048),
    .col_in_1049(u1_col_in_1049),
    .col_in_1050(u1_col_in_1050),
    .col_in_1051(u1_col_in_1051),
    .col_in_1052(u1_col_in_1052),
    .col_in_1053(u1_col_in_1053),
    .col_in_1054(u1_col_in_1054),
    .col_in_1055(u1_col_in_1055),
    .col_in_1056(u1_col_in_1056),
    .col_in_1057(u1_col_in_1057),
    .col_in_1058(u1_col_in_1058),
    .col_in_1059(u1_col_in_1059),
    .col_in_1060(u1_col_in_1060),
    .col_in_1061(u1_col_in_1061),
    .col_in_1062(u1_col_in_1062),
    .col_in_1063(u1_col_in_1063),
    .col_in_1064(u1_col_in_1064),
    .col_in_1065(u1_col_in_1065),
    .col_in_1066(u1_col_in_1066),
    .col_in_1067(u1_col_in_1067),
    .col_in_1068(u1_col_in_1068),
    .col_in_1069(u1_col_in_1069),
    .col_in_1070(u1_col_in_1070),
    .col_in_1071(u1_col_in_1071),
    .col_in_1072(u1_col_in_1072),
    .col_in_1073(u1_col_in_1073),
    .col_in_1074(u1_col_in_1074),
    .col_in_1075(u1_col_in_1075),
    .col_in_1076(u1_col_in_1076),
    .col_in_1077(u1_col_in_1077),
    .col_in_1078(u1_col_in_1078),
    .col_in_1079(u1_col_in_1079),
    .col_in_1080(u1_col_in_1080),
    .col_in_1081(u1_col_in_1081),
    .col_in_1082(u1_col_in_1082),
    .col_in_1083(u1_col_in_1083),
    .col_in_1084(u1_col_in_1084),
    .col_in_1085(u1_col_in_1085),
    .col_in_1086(u1_col_in_1086),
    .col_in_1087(u1_col_in_1087),
    .col_in_1088(u1_col_in_1088),
    .col_in_1089(u1_col_in_1089),
    .col_in_1090(u1_col_in_1090),
    .col_in_1091(u1_col_in_1091),
    .col_in_1092(u1_col_in_1092),
    .col_in_1093(u1_col_in_1093),
    .col_in_1094(u1_col_in_1094),
    .col_in_1095(u1_col_in_1095),
    .col_in_1096(u1_col_in_1096),
    .col_in_1097(u1_col_in_1097),
    .col_in_1098(u1_col_in_1098),
    .col_in_1099(u1_col_in_1099),
    .col_in_1100(u1_col_in_1100),
    .col_in_1101(u1_col_in_1101),
    .col_in_1102(u1_col_in_1102),
    .col_in_1103(u1_col_in_1103),
    .col_in_1104(u1_col_in_1104),
    .col_in_1105(u1_col_in_1105),
    .col_in_1106(u1_col_in_1106),
    .col_in_1107(u1_col_in_1107),
    .col_in_1108(u1_col_in_1108),
    .col_in_1109(u1_col_in_1109),
    .col_in_1110(u1_col_in_1110),
    .col_in_1111(u1_col_in_1111),
    .col_in_1112(u1_col_in_1112),
    .col_in_1113(u1_col_in_1113),
    .col_in_1114(u1_col_in_1114),
    .col_in_1115(u1_col_in_1115),
    .col_in_1116(u1_col_in_1116),
    .col_in_1117(u1_col_in_1117),
    .col_in_1118(u1_col_in_1118),
    .col_in_1119(u1_col_in_1119),
    .col_in_1120(u1_col_in_1120),
    .col_in_1121(u1_col_in_1121),
    .col_in_1122(u1_col_in_1122),
    .col_in_1123(u1_col_in_1123),
    .col_in_1124(u1_col_in_1124),
    .col_in_1125(u1_col_in_1125),
    .col_in_1126(u1_col_in_1126),
    .col_in_1127(u1_col_in_1127),
    .col_in_1128(u1_col_in_1128),
    .col_in_1129(u1_col_in_1129),
    .col_in_1130(u1_col_in_1130),
    .col_in_1131(u1_col_in_1131),
    .col_in_1132(u1_col_in_1132),
    .col_in_1133(u1_col_in_1133),
    .col_in_1134(u1_col_in_1134),
    .col_in_1135(u1_col_in_1135),
    .col_in_1136(u1_col_in_1136),
    .col_in_1137(u1_col_in_1137),
    .col_in_1138(u1_col_in_1138),
    .col_in_1139(u1_col_in_1139),
    .col_in_1140(u1_col_in_1140),
    .col_in_1141(u1_col_in_1141),
    .col_in_1142(u1_col_in_1142),
    .col_in_1143(u1_col_in_1143),
    .col_in_1144(u1_col_in_1144),
    .col_in_1145(u1_col_in_1145),
    .col_in_1146(u1_col_in_1146),
    .col_in_1147(u1_col_in_1147),
    .col_in_1148(u1_col_in_1148),
    .col_in_1149(u1_col_in_1149),
    .col_in_1150(u1_col_in_1150),
    .col_in_1151(u1_col_in_1151),
    .col_in_1152(u1_col_in_1152),
    .col_in_1153(u1_col_in_1153),
    .col_in_1154(u1_col_in_1154),
    .col_in_1155(u1_col_in_1155),
    .col_in_1156(u1_col_in_1156),
    .col_in_1157(u1_col_in_1157),
    .col_in_1158(u1_col_in_1158),
    .col_in_1159(u1_col_in_1159),
    .col_in_1160(u1_col_in_1160),
    .col_in_1161(u1_col_in_1161),
    .col_in_1162(u1_col_in_1162),
    .col_in_1163(u1_col_in_1163),
    .col_in_1164(u1_col_in_1164),
    .col_in_1165(u1_col_in_1165),
    .col_in_1166(u1_col_in_1166),
    .col_in_1167(u1_col_in_1167),
    .col_in_1168(u1_col_in_1168),
    .col_in_1169(u1_col_in_1169),
    .col_in_1170(u1_col_in_1170),
    .col_in_1171(u1_col_in_1171),
    .col_in_1172(u1_col_in_1172),
    .col_in_1173(u1_col_in_1173),
    .col_in_1174(u1_col_in_1174),
    .col_in_1175(u1_col_in_1175),
    .col_in_1176(u1_col_in_1176),
    .col_in_1177(u1_col_in_1177),
    .col_in_1178(u1_col_in_1178),
    .col_in_1179(u1_col_in_1179),
    .col_in_1180(u1_col_in_1180),
    .col_in_1181(u1_col_in_1181),
    .col_in_1182(u1_col_in_1182),
    .col_in_1183(u1_col_in_1183),
    .col_in_1184(u1_col_in_1184),
    .col_in_1185(u1_col_in_1185),
    .col_in_1186(u1_col_in_1186),
    .col_in_1187(u1_col_in_1187),
    .col_in_1188(u1_col_in_1188),
    .col_in_1189(u1_col_in_1189),
    .col_in_1190(u1_col_in_1190),
    .col_in_1191(u1_col_in_1191),
    .col_in_1192(u1_col_in_1192),
    .col_in_1193(u1_col_in_1193),
    .col_in_1194(u1_col_in_1194),
    .col_in_1195(u1_col_in_1195),
    .col_in_1196(u1_col_in_1196),
    .col_in_1197(u1_col_in_1197),
    .col_in_1198(u1_col_in_1198),
    .col_in_1199(u1_col_in_1199),
    .col_in_1200(u1_col_in_1200),
    .col_in_1201(u1_col_in_1201),
    .col_in_1202(u1_col_in_1202),
    .col_in_1203(u1_col_in_1203),
    .col_in_1204(u1_col_in_1204),
    .col_in_1205(u1_col_in_1205),
    .col_in_1206(u1_col_in_1206),
    .col_in_1207(u1_col_in_1207),
    .col_in_1208(u1_col_in_1208),
    .col_in_1209(u1_col_in_1209),
    .col_in_1210(u1_col_in_1210),
    .col_in_1211(u1_col_in_1211),
    .col_in_1212(u1_col_in_1212),
    .col_in_1213(u1_col_in_1213),
    .col_in_1214(u1_col_in_1214),
    .col_in_1215(u1_col_in_1215),
    .col_in_1216(u1_col_in_1216),
    .col_in_1217(u1_col_in_1217),
    .col_in_1218(u1_col_in_1218),
    .col_in_1219(u1_col_in_1219),
    .col_in_1220(u1_col_in_1220),
    .col_in_1221(u1_col_in_1221),
    .col_in_1222(u1_col_in_1222),
    .col_in_1223(u1_col_in_1223),
    .col_in_1224(u1_col_in_1224),
    .col_in_1225(u1_col_in_1225),
    .col_in_1226(u1_col_in_1226),
    .col_in_1227(u1_col_in_1227),
    .col_in_1228(u1_col_in_1228),
    .col_in_1229(u1_col_in_1229),
    .col_in_1230(u1_col_in_1230),
    .col_in_1231(u1_col_in_1231),
    .col_in_1232(u1_col_in_1232),
    .col_in_1233(u1_col_in_1233),
    .col_in_1234(u1_col_in_1234),
    .col_in_1235(u1_col_in_1235),
    .col_in_1236(u1_col_in_1236),
    .col_in_1237(u1_col_in_1237),
    .col_in_1238(u1_col_in_1238),
    .col_in_1239(u1_col_in_1239),
    .col_in_1240(u1_col_in_1240),
    .col_in_1241(u1_col_in_1241),
    .col_in_1242(u1_col_in_1242),
    .col_in_1243(u1_col_in_1243),
    .col_in_1244(u1_col_in_1244),
    .col_in_1245(u1_col_in_1245),
    .col_in_1246(u1_col_in_1246),
    .col_in_1247(u1_col_in_1247),
    .col_in_1248(u1_col_in_1248),
    .col_in_1249(u1_col_in_1249),
    .col_in_1250(u1_col_in_1250),
    .col_in_1251(u1_col_in_1251),
    .col_in_1252(u1_col_in_1252),
    .col_in_1253(u1_col_in_1253),
    .col_in_1254(u1_col_in_1254),
    .col_in_1255(u1_col_in_1255),
    .col_in_1256(u1_col_in_1256),
    .col_in_1257(u1_col_in_1257),
    .col_in_1258(u1_col_in_1258),
    .col_in_1259(u1_col_in_1259),
    .col_in_1260(u1_col_in_1260),
    .col_in_1261(u1_col_in_1261),
    .col_in_1262(u1_col_in_1262),
    .col_in_1263(u1_col_in_1263),
    .col_in_1264(u1_col_in_1264),
    .col_in_1265(u1_col_in_1265),
    .col_in_1266(u1_col_in_1266),
    .col_in_1267(u1_col_in_1267),
    .col_in_1268(u1_col_in_1268),
    .col_in_1269(u1_col_in_1269),
    .col_in_1270(u1_col_in_1270),
    .col_in_1271(u1_col_in_1271),
    .col_in_1272(u1_col_in_1272),
    .col_in_1273(u1_col_in_1273),
    .col_in_1274(u1_col_in_1274),
    .col_in_1275(u1_col_in_1275),
    .col_in_1276(u1_col_in_1276),
    .col_in_1277(u1_col_in_1277),
    .col_in_1278(u1_col_in_1278),
    .col_in_1279(u1_col_in_1279),


    .row_out_0(u1_row_out_0),
    .row_out_1(u1_row_out_1)
);


always@(posedge clk)begin
    if(rst)begin
        reg_intermediate0 <= 1288'h0;
        reg_intermediate1 <= 1288'h0;
    end
    else begin
        reg_intermediate0 <= u1_row_out_0;
        reg_intermediate1 <= u1_row_out_1;
    end
end









wire [6:0] u2_data_in;
wire [1023:0] u2_data_out;

assign u2_data_in = u1_row_out_0[1286:1280]  + u1_row_out_1[1286:1280];

xpb_7_0 u2_xpb_7_0
(
    .data_in(u2_data_in),
    .data_out(u2_data_out)
);

wire [1023:0] u3_d_out_c;
wire [1023:0] u3_d_out_s;

compressor_array_3_2_DW #(.DW(1024)) u3_compressor_array_3_2_1024
(
    .d_in0(u1_row_out_0[1279:256]),
    .d_in1(u1_row_out_1[1279:256]),
    .d_in2(u2_data_out),
    .d_out_c(u3_d_out_c),
    .d_out_s(u3_d_out_s)
);

(* max_fanout = 50 *)reg [1024:0] reg_c;
(* max_fanout = 50 *)reg [1023:0] reg_s;
always@(posedge clk)begin
    reg_c <= {u3_d_out_c, 1'b0};
    reg_s <= u3_d_out_s;
end



//-----------------------Stage 2------------------------------------

assign temp_ms0 = reg_c + reg_s;
assign temp_ms1 = reg_c + reg_s - P1;
assign temp_ms2 = reg_c + reg_s - P2;
assign temp_ms3 = reg_c + reg_s - P3;
always@(*)begin
    if(!temp_ms3[1026]) temp_ms = temp_ms3[1023:0];
    else if(!temp_ms2[1026]) temp_ms = temp_ms2[1023:0];
    else if(!temp_ms1[1026]) temp_ms = temp_ms1[1023:0];
    else temp_ms = temp_ms0[1023:0];
end


assign ms = temp_ms;



endmodule



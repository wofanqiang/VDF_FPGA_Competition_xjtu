module xpb_5_250
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h4d9f652598c5bb15f880b5de67467905bff3772cd5fee691d73553f1f2ce2392084561333ca35e044719c8993600fc1fb9b47cbc226c0522fdee91b7602801edb4a366e736efd50fc23d0aadf8fda46aab609a2924657e6fd6f4003ae6da2828f9f9896d96e33add4fe17e33d7285ff9616c03598d63fad1863e4122094e963c;
    5'b00010 : xpb = 1024'h9b3eca4b318b762bf1016bbcce8cf20b7fe6ee59abfdcd23ae6aa7e3e59c4724108ac2667946bc088e3391326c01f83f7368f97844d80a45fbdd236ec05003db6946cdce6ddfaa1f847a155bf1fb48d556c1345248cafcdfade80075cdb45051f3f312db2dc675ba9fc2fc67ae50bff2c2d806b31ac7f5a30c7c8244129d2c78;
    5'b00011 : xpb = 1024'h3830ea1b0862fc791e7ca9c4257923bfce646255ac85133e07c342802567bdae1587a620ebc39b7e35ef1a84bea4e394c9034e4e44913f1d492c75c7e5a59117a99b0006f53e81ea341d1d67521d290f0e1cd4e2e0aa4e3ecf4f6eb5fa63d5e8bee50a1f13e0b80a68e493bc8da8f9c2d56a2b2a57e093444c4b486193095c49;
    5'b00100 : xpb = 1024'h85d04f40a128b78f16fd5fa28cbf9cc58e57d9828283f9cfdef896721835e1401dcd07542866f9827d08e31df4a5dfb482b7cb0a66fd4440471b077f45cd93055e3e66ee2c2e56f9f65a28154b1acd79b97d6f0c050fccaea6436ef0e13dfe11b8de938caac3f2e7b8c611f064d159bc36d62e83e5448e15d28989839c57f285;
    5'b00101 : xpb = 1024'h22c26f1078003ddc44789da9e3abce79dcd54d7e830b3fea3851310e580157ca22c9eb0e9ae3d8f824c46c704748cb09d8521fe066b67917946a59d86b2320419e929926b38d2ec4a5fd3020ab3cadb370d90f9c9cef1e0dc7aadd310ded83a883d08ad090de353781e7a9454429938c496852fb225d2bb712584fa11cc42256;
    5'b00110 : xpb = 1024'h7061d43610c5f8f23cf953884af2477f9cc8c4ab590a267c0f8685004acf7b5c2b0f4c41d78736fc6bde35097d49c72992069c9c89227e3a9258eb8fcb4b222f5336000dea7d03d4683a3acea43a521e1c39a9c5c1549c7d9e9edd6bf4c7abd17dca143e27c17014d1c927791b51f385aad45654afc12688989690c32612b892;
    5'b00111 : xpb = 1024'hd53f405e79d7f3f6a74918fa1de7933eb4638a759916c9668df1f9c8a9af1e6300c2ffc4a0416721399be5bcfecb27ee7a0f17288dbb311dfa83de8f0a0af6b938a324671dbdb9f17dd42da045c3257d3954a565933eddcc0064bac2177316848bc0b820ddbb2649aeabecdfaaa2d55bd667acbecd9c429d86556e0a67ee863;
    5'b01000 : xpb = 1024'h5af3592b80633a5562f5476e0924f239ab39afd42f9053284014738e7d6915783851912f86a774765ab386f505edae9ea1556e2eab47b834dd96cfa050c8b159482d992da8cbb0aeda1a4d87fd59d6c27ef5e47f7d996c4c96fa4be70851599142b594efa4beed41eacc3d01d1d28d4f1ed27e257a3dbefb5ea39802afcd7e9f;
    5'b01001 : xpb = 1024'ha892be511928f56b5b75fd4c706b6b3f6b2d2701058f39ba1749c7807037390a4096f262c34ad27aa1cd4f8e3beeaabe5b09eaeacdb3bd57db856157b0f0b346fcd10014dfbb85be9c575835f6577b2d2a567ea8a1feeabc6dee4c21ef2b81ba3caf1e5d3ba2281f3aadbb35a8faed48803e817f07a1b9cce4e1d924b91c14db;
    5'b01010 : xpb = 1024'h4584de20f0007bb888f13b53c7579cf3b9aa9afd06167fd470a2621cb002af944593d61d35c7b1f04988d8e08e919613b0a43fc0cd6cf22f28d4b3b0d64640833d25324d671a5d894bfa604156795b66e1b21f3939de3c1b8f55ba621bdb075107a115a121bc6a6f03cf528a8853271892d0a5f644ba576e24b09f42398844ac;
    5'b01011 : xpb = 1024'h9324434688c636ce8171f1322e9e15f9799e1229dc15666647d7b60ea2d0d3264dd93750726b0ff490a2a179c49292336a58bc7cefd8f75226c34568366e4270f1c899349e0a32990e376aef4f76ffd18d12b9625e43ba8b6649ba9d02b52f7a019a9f0eb89fa54c53b0d0be5f7b8711f43ca94fd21e523faaeee06442d6dae8;
    5'b01100 : xpb = 1024'h301663165f9dbd1baeed2f39858a47adc81b8625dc9cac80a13050aae29c49b052d61b0ae4e7ef6a385e2acc17357d88bff31152ef922c29741297c15bc3cfad321ccb6d25690a63bdda72faaf98e00b446e59f2f6230bea87b128dd2f64b510cc8c96529eb9e79c1cd268133ed3c0e206cecdc70f36efe0eabda681c3430ab9;
    5'b01101 : xpb = 1024'h7db5c83bf8637831a76de517ecd0c0b3880efd52b29b93127865a49cd56a6d425b1b7c3e218b4d6e7f77f3654d3679a879a78e0f11fe314c72012978bbebd19ae6c032545c58df7380177da8a8968475efcef41c1a888a5a5ea52918163edd39c6861fc0359d22796cb3e64715fc20db683ad1209c9aeab270fbe7a3cc91a0f5;
    5'b01110 : xpb = 1024'h1aa7e80bcf3afe7ed4e9231f43bcf267d68c714eb322d92cd1be3f391535e3cc60185ff894082ce427337cb79fd964fdcf41e2e511b76623bf507bd1e1415ed72714648ce3b7b73e2fba85b408b864afa72a94acb267dbb9800c975842ee62d0917817041bb764c935d57d9bf5545aab7accf597d9b38853b0caadc14cfdd0c6;
    5'b01111 : xpb = 1024'h68474d316800b994cd69d8fdab036b6d967fe87b8921bfbea8f3932b0804075e685dc12bd0ab8ae86e4d4550d5da611d88f65fa134236b46bd3f0d89416960c4dbb7cb741aa78c4df1f7906201b6091a528b2ed5d6cd5a295700979329c88af98b71a071b29a9fa685b6fbcfcc7cbaa4dc38f8f1671783253708eee3564c6702;
    5'b10000 : xpb = 1024'h5396d013ed83fe1fae5170501ef9d21e4fd5c7789a905d9024c2dc747cf7de86d5aa4e643286a5e1608cea3287d4c72de90b47733dca01e0a8e5fe266beee011c0bfdaca2066418a19a986d61d7e95409e6cf666eacab88786805d356781090566397b598b4e1f64ed89324abd4f474eecb1d68a43020c676d7b500d6b896d3;
    5'b10001 : xpb = 1024'h52d8d226d79dfaf7f365cce369361627a4f0d3a45fa7ec6ad98181b93a9da17a75a006197fcbc8625d22973c5e7e4892984531335648a541087cf199c6e6efeed0af6493d8f6392863d7a31b5ad58dbeb547698f931229f84f5c060e3d5238b9505d21232f981cd39eba115882fd546e503720c231941b97fd15f622e0072d0f;
    5'b10010 : xpb = 1024'ha078374c7063b60debe682c1d07c8f2d64e44ad135a6d2fcb0b6d5ab2d6bc50c7de5674cbc6f2666a43c5fd5947f44b251f9adef78b4aa64066b8351270ef1dc8552cb7b0fe60e382614adc953d3322960a803b8b777a86826500649242c60e24a56aa90c67b57b0ee9b8f8c5a25b467b1a3241bbef8166983543744e955c34b;
    5'b10011 : xpb = 1024'h3d6a571c473b3c5b1961c0c92768c0e1b361becd362e19170a0f70476d373b9682e24b072eec05dc4bf7e927e7223007a79402c5786ddf3b53bad5aa4c647f18c5a6fdb39744e602d5b7b5d4b3f512631803a4494f56f9c747b7748950dbe6791548a1d4ac959a00b7bd26e1397dee37c4354892fc10b40ac322fd6269c1f31c;
    5'b10100 : xpb = 1024'h8b09bc41e000f77111e276a78eaf39e7735535fa0c2cffa8e144c43960055f288b27ac3a6b8f63e09311b1c11d232c2761487f819ad9e45e51a96761ac8c81067a4a649ace34bb1297f4c082acf2b6cdc3643e7273bc78371eab74c437b60ea20f422b424378d4de079ea51510a64e3125a14bec8974aedc49613e8473108958;
    5'b10101 : xpb = 1024'h27fbdc11b6d87dbe3f5db4aee59b6b9bc1d2a9f60cb445c33a9d5ed59fd0d5b290248ff4de0c43563acd3b136fc6177cb6e2d4579a9319359ef8b9bad1e20e42ba9e96d3559392dd4797c88e0d1497077abfdf030b9bc9964012e30464659438da3422862993172dd0c03c69effe880138337063c68d4c7d893004a1f37cb929;
    5'b10110 : xpb = 1024'h759b41374f9e38d437de6a8d4ce1e4a181c62122e2b32c5511d2b2c7929ef9449869f1281aafa15a81e703aca5c7139c70975113bcff1e589ce74b72320a10306f41fdba8c8367ed09d4d33c06123b722620792c300148061706e33f4b3fbc61d42dabf3c076520b20a1ba9dc726e7fa999f73bd53f1474f0f6e45c3fccb4f65;
    5'b10111 : xpb = 1024'h128d61072675bf216559a894a3ce1655d043951ee33a726f6b2b4d63d26a6fce9d66d4e28d2c80d029a28cfef869fef1c631a5e9bcb8532fea369dcb575f9d6caf962ff313e23fb7b977db4766341babdd7c19bcc7e09965386e517f77ef41f89f1fa337a690945ae9c351f2a67f21caac3198349109e4f04f3d0be17d377f36;
    5'b11000 : xpb = 1024'h602cc62cbf3b7a375dda5e730b148f5b90370c4bb93959014260a155c5389360a5ac3615c9cfded470bc55982e6afb117fe622a5df245852e8252f82b7879f5a643996da4ad214c77bb4e5f55f31c01688dcb3e5ec4617d50f6251ba5ec96a2199192ca53d73cf3839a4d0267da781c40d9d9b8e1e6ddfc1d57b4d0386861572;
    5'b11001 : xpb = 1024'hadcc2b525801354d565b1451725b0861502a83788f383f931995f547b806b6f2adf1974906733cd8b7d61e31646bf731399a9f6201905d75e613c13a17afa14818dcfdc181c1e9d73df1f0a3582f6481343d4e0f10ab9644e65651f545a3924a9312b612d4570a1589864e5a54cfe1bd6f099ee7abd1da935bb98e258fd4abae;
    5'b11010 : xpb = 1024'h4abe4b222ed8bb9a83d65258c9473a159ea7f7748fbf85ad72ee8fe3f7d22d7cb2ee7b0378f01c4e5f91a783b70ee2868f34f4380149924d336313933d052e8459312ffa0920c1a1ed94f8aeb85144baeb98ee9fa88ae7a407bdc035725317e15e04ad56ba714c6552a7e5af34281b8d819bc35ee8ea78349b8854431040db7f;
    5'b11011 : xpb = 1024'h985db047c79e76b07c570837308db31b5e9b6ea165be6c3f4a23e3d5eaa0510ebb33dc36b5937a52a6ab701ced0fdea648e970f423b597703151a54a9d2d30720dd496e1401096b1afd2035cb14ee92596f988c8ccf06613deb1c070592d400a57fe36c451548742a28963e30b507b86e307c6b8764e730621c69565198f71bb;
    5'b11100 : xpb = 1024'h354fd0179e75fcfda9d2463e8779e4cfad18e29d6645b259a37c7e722a6bc798c030bff1281059c84e66f96f3fb2c9fb9e83c5ca236ecc477ea0f7a3c282bdae4e28c919c76f6e7c5f750b681170c95f4e55295964cfb77300192eb085dcc5a122f02e08376ec9926baafb37eaa8b556f599eb2fb36710a761955b8299fba18c;
    5'b11101 : xpb = 1024'h82ef353d373bb813a252fc1ceec05dd56d0c59ca3c4498eb7ab1d2641d39eb2ac876212464b3b7cc9580c20875b3c61b5838428645dad16a7c8f895b22aabf9c02cc3000fe5f438c21b216160a6e6dc9f9b5c382893535e2d70d2eeb6cb6edca1ce9b775ce52046fbb8c796bc1d115505705ee8940cb0b78e7d39ca4a34a37c8;
    5'b11110 : xpb = 1024'h1fe1550d0e133e60cfce3a2445ac8f89bb89cdc63ccbdf05d40a6d005d0561b4cd7304ded73097423d3c4b5ac856b170add2975c45940641c9dedbb448004cd84320623985be1b56d1551e216a904e03b111641321148741f8749d2b99667360e7dbaeb9b46c46bf84ae10c0a1294f20699813007de3a91a27a262c223b66799;
    5'b11111 : xpb = 1024'h6d80ba32a6d8f976c84ef002acf3088f7b7d44f312cac597ab3fc0f24fd38546d5b8661213d3f546845613f3fe57ad906787141868000b64c7cd6d6ba8284ec5f7c3c920bcadf066939228cf638df26e5c71fe3c457a05b1cf689d6680409b89e1d538274b4f819cd48f8ef47851af19cb04165a0b47a3ebade0a3e42d04fdd5;
    endcase
end

endmodule

module compressor_array_3_2_1024_row
(
    input [1023:0] row_in_0,
    input [1023:0] row_in_1,
    input [1023:0] row_in_2,

    output [1024:0] row_out_0,
    output [1024:0] row_out_1
);











wire [2:0] col_in_0;
wire [2:0] col_in_1;
wire [2:0] col_in_2;
wire [2:0] col_in_3;
wire [2:0] col_in_4;
wire [2:0] col_in_5;
wire [2:0] col_in_6;
wire [2:0] col_in_7;
wire [2:0] col_in_8;
wire [2:0] col_in_9;
wire [2:0] col_in_10;
wire [2:0] col_in_11;
wire [2:0] col_in_12;
wire [2:0] col_in_13;
wire [2:0] col_in_14;
wire [2:0] col_in_15;
wire [2:0] col_in_16;
wire [2:0] col_in_17;
wire [2:0] col_in_18;
wire [2:0] col_in_19;
wire [2:0] col_in_20;
wire [2:0] col_in_21;
wire [2:0] col_in_22;
wire [2:0] col_in_23;
wire [2:0] col_in_24;
wire [2:0] col_in_25;
wire [2:0] col_in_26;
wire [2:0] col_in_27;
wire [2:0] col_in_28;
wire [2:0] col_in_29;
wire [2:0] col_in_30;
wire [2:0] col_in_31;
wire [2:0] col_in_32;
wire [2:0] col_in_33;
wire [2:0] col_in_34;
wire [2:0] col_in_35;
wire [2:0] col_in_36;
wire [2:0] col_in_37;
wire [2:0] col_in_38;
wire [2:0] col_in_39;
wire [2:0] col_in_40;
wire [2:0] col_in_41;
wire [2:0] col_in_42;
wire [2:0] col_in_43;
wire [2:0] col_in_44;
wire [2:0] col_in_45;
wire [2:0] col_in_46;
wire [2:0] col_in_47;
wire [2:0] col_in_48;
wire [2:0] col_in_49;
wire [2:0] col_in_50;
wire [2:0] col_in_51;
wire [2:0] col_in_52;
wire [2:0] col_in_53;
wire [2:0] col_in_54;
wire [2:0] col_in_55;
wire [2:0] col_in_56;
wire [2:0] col_in_57;
wire [2:0] col_in_58;
wire [2:0] col_in_59;
wire [2:0] col_in_60;
wire [2:0] col_in_61;
wire [2:0] col_in_62;
wire [2:0] col_in_63;
wire [2:0] col_in_64;
wire [2:0] col_in_65;
wire [2:0] col_in_66;
wire [2:0] col_in_67;
wire [2:0] col_in_68;
wire [2:0] col_in_69;
wire [2:0] col_in_70;
wire [2:0] col_in_71;
wire [2:0] col_in_72;
wire [2:0] col_in_73;
wire [2:0] col_in_74;
wire [2:0] col_in_75;
wire [2:0] col_in_76;
wire [2:0] col_in_77;
wire [2:0] col_in_78;
wire [2:0] col_in_79;
wire [2:0] col_in_80;
wire [2:0] col_in_81;
wire [2:0] col_in_82;
wire [2:0] col_in_83;
wire [2:0] col_in_84;
wire [2:0] col_in_85;
wire [2:0] col_in_86;
wire [2:0] col_in_87;
wire [2:0] col_in_88;
wire [2:0] col_in_89;
wire [2:0] col_in_90;
wire [2:0] col_in_91;
wire [2:0] col_in_92;
wire [2:0] col_in_93;
wire [2:0] col_in_94;
wire [2:0] col_in_95;
wire [2:0] col_in_96;
wire [2:0] col_in_97;
wire [2:0] col_in_98;
wire [2:0] col_in_99;
wire [2:0] col_in_100;
wire [2:0] col_in_101;
wire [2:0] col_in_102;
wire [2:0] col_in_103;
wire [2:0] col_in_104;
wire [2:0] col_in_105;
wire [2:0] col_in_106;
wire [2:0] col_in_107;
wire [2:0] col_in_108;
wire [2:0] col_in_109;
wire [2:0] col_in_110;
wire [2:0] col_in_111;
wire [2:0] col_in_112;
wire [2:0] col_in_113;
wire [2:0] col_in_114;
wire [2:0] col_in_115;
wire [2:0] col_in_116;
wire [2:0] col_in_117;
wire [2:0] col_in_118;
wire [2:0] col_in_119;
wire [2:0] col_in_120;
wire [2:0] col_in_121;
wire [2:0] col_in_122;
wire [2:0] col_in_123;
wire [2:0] col_in_124;
wire [2:0] col_in_125;
wire [2:0] col_in_126;
wire [2:0] col_in_127;
wire [2:0] col_in_128;
wire [2:0] col_in_129;
wire [2:0] col_in_130;
wire [2:0] col_in_131;
wire [2:0] col_in_132;
wire [2:0] col_in_133;
wire [2:0] col_in_134;
wire [2:0] col_in_135;
wire [2:0] col_in_136;
wire [2:0] col_in_137;
wire [2:0] col_in_138;
wire [2:0] col_in_139;
wire [2:0] col_in_140;
wire [2:0] col_in_141;
wire [2:0] col_in_142;
wire [2:0] col_in_143;
wire [2:0] col_in_144;
wire [2:0] col_in_145;
wire [2:0] col_in_146;
wire [2:0] col_in_147;
wire [2:0] col_in_148;
wire [2:0] col_in_149;
wire [2:0] col_in_150;
wire [2:0] col_in_151;
wire [2:0] col_in_152;
wire [2:0] col_in_153;
wire [2:0] col_in_154;
wire [2:0] col_in_155;
wire [2:0] col_in_156;
wire [2:0] col_in_157;
wire [2:0] col_in_158;
wire [2:0] col_in_159;
wire [2:0] col_in_160;
wire [2:0] col_in_161;
wire [2:0] col_in_162;
wire [2:0] col_in_163;
wire [2:0] col_in_164;
wire [2:0] col_in_165;
wire [2:0] col_in_166;
wire [2:0] col_in_167;
wire [2:0] col_in_168;
wire [2:0] col_in_169;
wire [2:0] col_in_170;
wire [2:0] col_in_171;
wire [2:0] col_in_172;
wire [2:0] col_in_173;
wire [2:0] col_in_174;
wire [2:0] col_in_175;
wire [2:0] col_in_176;
wire [2:0] col_in_177;
wire [2:0] col_in_178;
wire [2:0] col_in_179;
wire [2:0] col_in_180;
wire [2:0] col_in_181;
wire [2:0] col_in_182;
wire [2:0] col_in_183;
wire [2:0] col_in_184;
wire [2:0] col_in_185;
wire [2:0] col_in_186;
wire [2:0] col_in_187;
wire [2:0] col_in_188;
wire [2:0] col_in_189;
wire [2:0] col_in_190;
wire [2:0] col_in_191;
wire [2:0] col_in_192;
wire [2:0] col_in_193;
wire [2:0] col_in_194;
wire [2:0] col_in_195;
wire [2:0] col_in_196;
wire [2:0] col_in_197;
wire [2:0] col_in_198;
wire [2:0] col_in_199;
wire [2:0] col_in_200;
wire [2:0] col_in_201;
wire [2:0] col_in_202;
wire [2:0] col_in_203;
wire [2:0] col_in_204;
wire [2:0] col_in_205;
wire [2:0] col_in_206;
wire [2:0] col_in_207;
wire [2:0] col_in_208;
wire [2:0] col_in_209;
wire [2:0] col_in_210;
wire [2:0] col_in_211;
wire [2:0] col_in_212;
wire [2:0] col_in_213;
wire [2:0] col_in_214;
wire [2:0] col_in_215;
wire [2:0] col_in_216;
wire [2:0] col_in_217;
wire [2:0] col_in_218;
wire [2:0] col_in_219;
wire [2:0] col_in_220;
wire [2:0] col_in_221;
wire [2:0] col_in_222;
wire [2:0] col_in_223;
wire [2:0] col_in_224;
wire [2:0] col_in_225;
wire [2:0] col_in_226;
wire [2:0] col_in_227;
wire [2:0] col_in_228;
wire [2:0] col_in_229;
wire [2:0] col_in_230;
wire [2:0] col_in_231;
wire [2:0] col_in_232;
wire [2:0] col_in_233;
wire [2:0] col_in_234;
wire [2:0] col_in_235;
wire [2:0] col_in_236;
wire [2:0] col_in_237;
wire [2:0] col_in_238;
wire [2:0] col_in_239;
wire [2:0] col_in_240;
wire [2:0] col_in_241;
wire [2:0] col_in_242;
wire [2:0] col_in_243;
wire [2:0] col_in_244;
wire [2:0] col_in_245;
wire [2:0] col_in_246;
wire [2:0] col_in_247;
wire [2:0] col_in_248;
wire [2:0] col_in_249;
wire [2:0] col_in_250;
wire [2:0] col_in_251;
wire [2:0] col_in_252;
wire [2:0] col_in_253;
wire [2:0] col_in_254;
wire [2:0] col_in_255;
wire [2:0] col_in_256;
wire [2:0] col_in_257;
wire [2:0] col_in_258;
wire [2:0] col_in_259;
wire [2:0] col_in_260;
wire [2:0] col_in_261;
wire [2:0] col_in_262;
wire [2:0] col_in_263;
wire [2:0] col_in_264;
wire [2:0] col_in_265;
wire [2:0] col_in_266;
wire [2:0] col_in_267;
wire [2:0] col_in_268;
wire [2:0] col_in_269;
wire [2:0] col_in_270;
wire [2:0] col_in_271;
wire [2:0] col_in_272;
wire [2:0] col_in_273;
wire [2:0] col_in_274;
wire [2:0] col_in_275;
wire [2:0] col_in_276;
wire [2:0] col_in_277;
wire [2:0] col_in_278;
wire [2:0] col_in_279;
wire [2:0] col_in_280;
wire [2:0] col_in_281;
wire [2:0] col_in_282;
wire [2:0] col_in_283;
wire [2:0] col_in_284;
wire [2:0] col_in_285;
wire [2:0] col_in_286;
wire [2:0] col_in_287;
wire [2:0] col_in_288;
wire [2:0] col_in_289;
wire [2:0] col_in_290;
wire [2:0] col_in_291;
wire [2:0] col_in_292;
wire [2:0] col_in_293;
wire [2:0] col_in_294;
wire [2:0] col_in_295;
wire [2:0] col_in_296;
wire [2:0] col_in_297;
wire [2:0] col_in_298;
wire [2:0] col_in_299;
wire [2:0] col_in_300;
wire [2:0] col_in_301;
wire [2:0] col_in_302;
wire [2:0] col_in_303;
wire [2:0] col_in_304;
wire [2:0] col_in_305;
wire [2:0] col_in_306;
wire [2:0] col_in_307;
wire [2:0] col_in_308;
wire [2:0] col_in_309;
wire [2:0] col_in_310;
wire [2:0] col_in_311;
wire [2:0] col_in_312;
wire [2:0] col_in_313;
wire [2:0] col_in_314;
wire [2:0] col_in_315;
wire [2:0] col_in_316;
wire [2:0] col_in_317;
wire [2:0] col_in_318;
wire [2:0] col_in_319;
wire [2:0] col_in_320;
wire [2:0] col_in_321;
wire [2:0] col_in_322;
wire [2:0] col_in_323;
wire [2:0] col_in_324;
wire [2:0] col_in_325;
wire [2:0] col_in_326;
wire [2:0] col_in_327;
wire [2:0] col_in_328;
wire [2:0] col_in_329;
wire [2:0] col_in_330;
wire [2:0] col_in_331;
wire [2:0] col_in_332;
wire [2:0] col_in_333;
wire [2:0] col_in_334;
wire [2:0] col_in_335;
wire [2:0] col_in_336;
wire [2:0] col_in_337;
wire [2:0] col_in_338;
wire [2:0] col_in_339;
wire [2:0] col_in_340;
wire [2:0] col_in_341;
wire [2:0] col_in_342;
wire [2:0] col_in_343;
wire [2:0] col_in_344;
wire [2:0] col_in_345;
wire [2:0] col_in_346;
wire [2:0] col_in_347;
wire [2:0] col_in_348;
wire [2:0] col_in_349;
wire [2:0] col_in_350;
wire [2:0] col_in_351;
wire [2:0] col_in_352;
wire [2:0] col_in_353;
wire [2:0] col_in_354;
wire [2:0] col_in_355;
wire [2:0] col_in_356;
wire [2:0] col_in_357;
wire [2:0] col_in_358;
wire [2:0] col_in_359;
wire [2:0] col_in_360;
wire [2:0] col_in_361;
wire [2:0] col_in_362;
wire [2:0] col_in_363;
wire [2:0] col_in_364;
wire [2:0] col_in_365;
wire [2:0] col_in_366;
wire [2:0] col_in_367;
wire [2:0] col_in_368;
wire [2:0] col_in_369;
wire [2:0] col_in_370;
wire [2:0] col_in_371;
wire [2:0] col_in_372;
wire [2:0] col_in_373;
wire [2:0] col_in_374;
wire [2:0] col_in_375;
wire [2:0] col_in_376;
wire [2:0] col_in_377;
wire [2:0] col_in_378;
wire [2:0] col_in_379;
wire [2:0] col_in_380;
wire [2:0] col_in_381;
wire [2:0] col_in_382;
wire [2:0] col_in_383;
wire [2:0] col_in_384;
wire [2:0] col_in_385;
wire [2:0] col_in_386;
wire [2:0] col_in_387;
wire [2:0] col_in_388;
wire [2:0] col_in_389;
wire [2:0] col_in_390;
wire [2:0] col_in_391;
wire [2:0] col_in_392;
wire [2:0] col_in_393;
wire [2:0] col_in_394;
wire [2:0] col_in_395;
wire [2:0] col_in_396;
wire [2:0] col_in_397;
wire [2:0] col_in_398;
wire [2:0] col_in_399;
wire [2:0] col_in_400;
wire [2:0] col_in_401;
wire [2:0] col_in_402;
wire [2:0] col_in_403;
wire [2:0] col_in_404;
wire [2:0] col_in_405;
wire [2:0] col_in_406;
wire [2:0] col_in_407;
wire [2:0] col_in_408;
wire [2:0] col_in_409;
wire [2:0] col_in_410;
wire [2:0] col_in_411;
wire [2:0] col_in_412;
wire [2:0] col_in_413;
wire [2:0] col_in_414;
wire [2:0] col_in_415;
wire [2:0] col_in_416;
wire [2:0] col_in_417;
wire [2:0] col_in_418;
wire [2:0] col_in_419;
wire [2:0] col_in_420;
wire [2:0] col_in_421;
wire [2:0] col_in_422;
wire [2:0] col_in_423;
wire [2:0] col_in_424;
wire [2:0] col_in_425;
wire [2:0] col_in_426;
wire [2:0] col_in_427;
wire [2:0] col_in_428;
wire [2:0] col_in_429;
wire [2:0] col_in_430;
wire [2:0] col_in_431;
wire [2:0] col_in_432;
wire [2:0] col_in_433;
wire [2:0] col_in_434;
wire [2:0] col_in_435;
wire [2:0] col_in_436;
wire [2:0] col_in_437;
wire [2:0] col_in_438;
wire [2:0] col_in_439;
wire [2:0] col_in_440;
wire [2:0] col_in_441;
wire [2:0] col_in_442;
wire [2:0] col_in_443;
wire [2:0] col_in_444;
wire [2:0] col_in_445;
wire [2:0] col_in_446;
wire [2:0] col_in_447;
wire [2:0] col_in_448;
wire [2:0] col_in_449;
wire [2:0] col_in_450;
wire [2:0] col_in_451;
wire [2:0] col_in_452;
wire [2:0] col_in_453;
wire [2:0] col_in_454;
wire [2:0] col_in_455;
wire [2:0] col_in_456;
wire [2:0] col_in_457;
wire [2:0] col_in_458;
wire [2:0] col_in_459;
wire [2:0] col_in_460;
wire [2:0] col_in_461;
wire [2:0] col_in_462;
wire [2:0] col_in_463;
wire [2:0] col_in_464;
wire [2:0] col_in_465;
wire [2:0] col_in_466;
wire [2:0] col_in_467;
wire [2:0] col_in_468;
wire [2:0] col_in_469;
wire [2:0] col_in_470;
wire [2:0] col_in_471;
wire [2:0] col_in_472;
wire [2:0] col_in_473;
wire [2:0] col_in_474;
wire [2:0] col_in_475;
wire [2:0] col_in_476;
wire [2:0] col_in_477;
wire [2:0] col_in_478;
wire [2:0] col_in_479;
wire [2:0] col_in_480;
wire [2:0] col_in_481;
wire [2:0] col_in_482;
wire [2:0] col_in_483;
wire [2:0] col_in_484;
wire [2:0] col_in_485;
wire [2:0] col_in_486;
wire [2:0] col_in_487;
wire [2:0] col_in_488;
wire [2:0] col_in_489;
wire [2:0] col_in_490;
wire [2:0] col_in_491;
wire [2:0] col_in_492;
wire [2:0] col_in_493;
wire [2:0] col_in_494;
wire [2:0] col_in_495;
wire [2:0] col_in_496;
wire [2:0] col_in_497;
wire [2:0] col_in_498;
wire [2:0] col_in_499;
wire [2:0] col_in_500;
wire [2:0] col_in_501;
wire [2:0] col_in_502;
wire [2:0] col_in_503;
wire [2:0] col_in_504;
wire [2:0] col_in_505;
wire [2:0] col_in_506;
wire [2:0] col_in_507;
wire [2:0] col_in_508;
wire [2:0] col_in_509;
wire [2:0] col_in_510;
wire [2:0] col_in_511;
wire [2:0] col_in_512;
wire [2:0] col_in_513;
wire [2:0] col_in_514;
wire [2:0] col_in_515;
wire [2:0] col_in_516;
wire [2:0] col_in_517;
wire [2:0] col_in_518;
wire [2:0] col_in_519;
wire [2:0] col_in_520;
wire [2:0] col_in_521;
wire [2:0] col_in_522;
wire [2:0] col_in_523;
wire [2:0] col_in_524;
wire [2:0] col_in_525;
wire [2:0] col_in_526;
wire [2:0] col_in_527;
wire [2:0] col_in_528;
wire [2:0] col_in_529;
wire [2:0] col_in_530;
wire [2:0] col_in_531;
wire [2:0] col_in_532;
wire [2:0] col_in_533;
wire [2:0] col_in_534;
wire [2:0] col_in_535;
wire [2:0] col_in_536;
wire [2:0] col_in_537;
wire [2:0] col_in_538;
wire [2:0] col_in_539;
wire [2:0] col_in_540;
wire [2:0] col_in_541;
wire [2:0] col_in_542;
wire [2:0] col_in_543;
wire [2:0] col_in_544;
wire [2:0] col_in_545;
wire [2:0] col_in_546;
wire [2:0] col_in_547;
wire [2:0] col_in_548;
wire [2:0] col_in_549;
wire [2:0] col_in_550;
wire [2:0] col_in_551;
wire [2:0] col_in_552;
wire [2:0] col_in_553;
wire [2:0] col_in_554;
wire [2:0] col_in_555;
wire [2:0] col_in_556;
wire [2:0] col_in_557;
wire [2:0] col_in_558;
wire [2:0] col_in_559;
wire [2:0] col_in_560;
wire [2:0] col_in_561;
wire [2:0] col_in_562;
wire [2:0] col_in_563;
wire [2:0] col_in_564;
wire [2:0] col_in_565;
wire [2:0] col_in_566;
wire [2:0] col_in_567;
wire [2:0] col_in_568;
wire [2:0] col_in_569;
wire [2:0] col_in_570;
wire [2:0] col_in_571;
wire [2:0] col_in_572;
wire [2:0] col_in_573;
wire [2:0] col_in_574;
wire [2:0] col_in_575;
wire [2:0] col_in_576;
wire [2:0] col_in_577;
wire [2:0] col_in_578;
wire [2:0] col_in_579;
wire [2:0] col_in_580;
wire [2:0] col_in_581;
wire [2:0] col_in_582;
wire [2:0] col_in_583;
wire [2:0] col_in_584;
wire [2:0] col_in_585;
wire [2:0] col_in_586;
wire [2:0] col_in_587;
wire [2:0] col_in_588;
wire [2:0] col_in_589;
wire [2:0] col_in_590;
wire [2:0] col_in_591;
wire [2:0] col_in_592;
wire [2:0] col_in_593;
wire [2:0] col_in_594;
wire [2:0] col_in_595;
wire [2:0] col_in_596;
wire [2:0] col_in_597;
wire [2:0] col_in_598;
wire [2:0] col_in_599;
wire [2:0] col_in_600;
wire [2:0] col_in_601;
wire [2:0] col_in_602;
wire [2:0] col_in_603;
wire [2:0] col_in_604;
wire [2:0] col_in_605;
wire [2:0] col_in_606;
wire [2:0] col_in_607;
wire [2:0] col_in_608;
wire [2:0] col_in_609;
wire [2:0] col_in_610;
wire [2:0] col_in_611;
wire [2:0] col_in_612;
wire [2:0] col_in_613;
wire [2:0] col_in_614;
wire [2:0] col_in_615;
wire [2:0] col_in_616;
wire [2:0] col_in_617;
wire [2:0] col_in_618;
wire [2:0] col_in_619;
wire [2:0] col_in_620;
wire [2:0] col_in_621;
wire [2:0] col_in_622;
wire [2:0] col_in_623;
wire [2:0] col_in_624;
wire [2:0] col_in_625;
wire [2:0] col_in_626;
wire [2:0] col_in_627;
wire [2:0] col_in_628;
wire [2:0] col_in_629;
wire [2:0] col_in_630;
wire [2:0] col_in_631;
wire [2:0] col_in_632;
wire [2:0] col_in_633;
wire [2:0] col_in_634;
wire [2:0] col_in_635;
wire [2:0] col_in_636;
wire [2:0] col_in_637;
wire [2:0] col_in_638;
wire [2:0] col_in_639;
wire [2:0] col_in_640;
wire [2:0] col_in_641;
wire [2:0] col_in_642;
wire [2:0] col_in_643;
wire [2:0] col_in_644;
wire [2:0] col_in_645;
wire [2:0] col_in_646;
wire [2:0] col_in_647;
wire [2:0] col_in_648;
wire [2:0] col_in_649;
wire [2:0] col_in_650;
wire [2:0] col_in_651;
wire [2:0] col_in_652;
wire [2:0] col_in_653;
wire [2:0] col_in_654;
wire [2:0] col_in_655;
wire [2:0] col_in_656;
wire [2:0] col_in_657;
wire [2:0] col_in_658;
wire [2:0] col_in_659;
wire [2:0] col_in_660;
wire [2:0] col_in_661;
wire [2:0] col_in_662;
wire [2:0] col_in_663;
wire [2:0] col_in_664;
wire [2:0] col_in_665;
wire [2:0] col_in_666;
wire [2:0] col_in_667;
wire [2:0] col_in_668;
wire [2:0] col_in_669;
wire [2:0] col_in_670;
wire [2:0] col_in_671;
wire [2:0] col_in_672;
wire [2:0] col_in_673;
wire [2:0] col_in_674;
wire [2:0] col_in_675;
wire [2:0] col_in_676;
wire [2:0] col_in_677;
wire [2:0] col_in_678;
wire [2:0] col_in_679;
wire [2:0] col_in_680;
wire [2:0] col_in_681;
wire [2:0] col_in_682;
wire [2:0] col_in_683;
wire [2:0] col_in_684;
wire [2:0] col_in_685;
wire [2:0] col_in_686;
wire [2:0] col_in_687;
wire [2:0] col_in_688;
wire [2:0] col_in_689;
wire [2:0] col_in_690;
wire [2:0] col_in_691;
wire [2:0] col_in_692;
wire [2:0] col_in_693;
wire [2:0] col_in_694;
wire [2:0] col_in_695;
wire [2:0] col_in_696;
wire [2:0] col_in_697;
wire [2:0] col_in_698;
wire [2:0] col_in_699;
wire [2:0] col_in_700;
wire [2:0] col_in_701;
wire [2:0] col_in_702;
wire [2:0] col_in_703;
wire [2:0] col_in_704;
wire [2:0] col_in_705;
wire [2:0] col_in_706;
wire [2:0] col_in_707;
wire [2:0] col_in_708;
wire [2:0] col_in_709;
wire [2:0] col_in_710;
wire [2:0] col_in_711;
wire [2:0] col_in_712;
wire [2:0] col_in_713;
wire [2:0] col_in_714;
wire [2:0] col_in_715;
wire [2:0] col_in_716;
wire [2:0] col_in_717;
wire [2:0] col_in_718;
wire [2:0] col_in_719;
wire [2:0] col_in_720;
wire [2:0] col_in_721;
wire [2:0] col_in_722;
wire [2:0] col_in_723;
wire [2:0] col_in_724;
wire [2:0] col_in_725;
wire [2:0] col_in_726;
wire [2:0] col_in_727;
wire [2:0] col_in_728;
wire [2:0] col_in_729;
wire [2:0] col_in_730;
wire [2:0] col_in_731;
wire [2:0] col_in_732;
wire [2:0] col_in_733;
wire [2:0] col_in_734;
wire [2:0] col_in_735;
wire [2:0] col_in_736;
wire [2:0] col_in_737;
wire [2:0] col_in_738;
wire [2:0] col_in_739;
wire [2:0] col_in_740;
wire [2:0] col_in_741;
wire [2:0] col_in_742;
wire [2:0] col_in_743;
wire [2:0] col_in_744;
wire [2:0] col_in_745;
wire [2:0] col_in_746;
wire [2:0] col_in_747;
wire [2:0] col_in_748;
wire [2:0] col_in_749;
wire [2:0] col_in_750;
wire [2:0] col_in_751;
wire [2:0] col_in_752;
wire [2:0] col_in_753;
wire [2:0] col_in_754;
wire [2:0] col_in_755;
wire [2:0] col_in_756;
wire [2:0] col_in_757;
wire [2:0] col_in_758;
wire [2:0] col_in_759;
wire [2:0] col_in_760;
wire [2:0] col_in_761;
wire [2:0] col_in_762;
wire [2:0] col_in_763;
wire [2:0] col_in_764;
wire [2:0] col_in_765;
wire [2:0] col_in_766;
wire [2:0] col_in_767;
wire [2:0] col_in_768;
wire [2:0] col_in_769;
wire [2:0] col_in_770;
wire [2:0] col_in_771;
wire [2:0] col_in_772;
wire [2:0] col_in_773;
wire [2:0] col_in_774;
wire [2:0] col_in_775;
wire [2:0] col_in_776;
wire [2:0] col_in_777;
wire [2:0] col_in_778;
wire [2:0] col_in_779;
wire [2:0] col_in_780;
wire [2:0] col_in_781;
wire [2:0] col_in_782;
wire [2:0] col_in_783;
wire [2:0] col_in_784;
wire [2:0] col_in_785;
wire [2:0] col_in_786;
wire [2:0] col_in_787;
wire [2:0] col_in_788;
wire [2:0] col_in_789;
wire [2:0] col_in_790;
wire [2:0] col_in_791;
wire [2:0] col_in_792;
wire [2:0] col_in_793;
wire [2:0] col_in_794;
wire [2:0] col_in_795;
wire [2:0] col_in_796;
wire [2:0] col_in_797;
wire [2:0] col_in_798;
wire [2:0] col_in_799;
wire [2:0] col_in_800;
wire [2:0] col_in_801;
wire [2:0] col_in_802;
wire [2:0] col_in_803;
wire [2:0] col_in_804;
wire [2:0] col_in_805;
wire [2:0] col_in_806;
wire [2:0] col_in_807;
wire [2:0] col_in_808;
wire [2:0] col_in_809;
wire [2:0] col_in_810;
wire [2:0] col_in_811;
wire [2:0] col_in_812;
wire [2:0] col_in_813;
wire [2:0] col_in_814;
wire [2:0] col_in_815;
wire [2:0] col_in_816;
wire [2:0] col_in_817;
wire [2:0] col_in_818;
wire [2:0] col_in_819;
wire [2:0] col_in_820;
wire [2:0] col_in_821;
wire [2:0] col_in_822;
wire [2:0] col_in_823;
wire [2:0] col_in_824;
wire [2:0] col_in_825;
wire [2:0] col_in_826;
wire [2:0] col_in_827;
wire [2:0] col_in_828;
wire [2:0] col_in_829;
wire [2:0] col_in_830;
wire [2:0] col_in_831;
wire [2:0] col_in_832;
wire [2:0] col_in_833;
wire [2:0] col_in_834;
wire [2:0] col_in_835;
wire [2:0] col_in_836;
wire [2:0] col_in_837;
wire [2:0] col_in_838;
wire [2:0] col_in_839;
wire [2:0] col_in_840;
wire [2:0] col_in_841;
wire [2:0] col_in_842;
wire [2:0] col_in_843;
wire [2:0] col_in_844;
wire [2:0] col_in_845;
wire [2:0] col_in_846;
wire [2:0] col_in_847;
wire [2:0] col_in_848;
wire [2:0] col_in_849;
wire [2:0] col_in_850;
wire [2:0] col_in_851;
wire [2:0] col_in_852;
wire [2:0] col_in_853;
wire [2:0] col_in_854;
wire [2:0] col_in_855;
wire [2:0] col_in_856;
wire [2:0] col_in_857;
wire [2:0] col_in_858;
wire [2:0] col_in_859;
wire [2:0] col_in_860;
wire [2:0] col_in_861;
wire [2:0] col_in_862;
wire [2:0] col_in_863;
wire [2:0] col_in_864;
wire [2:0] col_in_865;
wire [2:0] col_in_866;
wire [2:0] col_in_867;
wire [2:0] col_in_868;
wire [2:0] col_in_869;
wire [2:0] col_in_870;
wire [2:0] col_in_871;
wire [2:0] col_in_872;
wire [2:0] col_in_873;
wire [2:0] col_in_874;
wire [2:0] col_in_875;
wire [2:0] col_in_876;
wire [2:0] col_in_877;
wire [2:0] col_in_878;
wire [2:0] col_in_879;
wire [2:0] col_in_880;
wire [2:0] col_in_881;
wire [2:0] col_in_882;
wire [2:0] col_in_883;
wire [2:0] col_in_884;
wire [2:0] col_in_885;
wire [2:0] col_in_886;
wire [2:0] col_in_887;
wire [2:0] col_in_888;
wire [2:0] col_in_889;
wire [2:0] col_in_890;
wire [2:0] col_in_891;
wire [2:0] col_in_892;
wire [2:0] col_in_893;
wire [2:0] col_in_894;
wire [2:0] col_in_895;
wire [2:0] col_in_896;
wire [2:0] col_in_897;
wire [2:0] col_in_898;
wire [2:0] col_in_899;
wire [2:0] col_in_900;
wire [2:0] col_in_901;
wire [2:0] col_in_902;
wire [2:0] col_in_903;
wire [2:0] col_in_904;
wire [2:0] col_in_905;
wire [2:0] col_in_906;
wire [2:0] col_in_907;
wire [2:0] col_in_908;
wire [2:0] col_in_909;
wire [2:0] col_in_910;
wire [2:0] col_in_911;
wire [2:0] col_in_912;
wire [2:0] col_in_913;
wire [2:0] col_in_914;
wire [2:0] col_in_915;
wire [2:0] col_in_916;
wire [2:0] col_in_917;
wire [2:0] col_in_918;
wire [2:0] col_in_919;
wire [2:0] col_in_920;
wire [2:0] col_in_921;
wire [2:0] col_in_922;
wire [2:0] col_in_923;
wire [2:0] col_in_924;
wire [2:0] col_in_925;
wire [2:0] col_in_926;
wire [2:0] col_in_927;
wire [2:0] col_in_928;
wire [2:0] col_in_929;
wire [2:0] col_in_930;
wire [2:0] col_in_931;
wire [2:0] col_in_932;
wire [2:0] col_in_933;
wire [2:0] col_in_934;
wire [2:0] col_in_935;
wire [2:0] col_in_936;
wire [2:0] col_in_937;
wire [2:0] col_in_938;
wire [2:0] col_in_939;
wire [2:0] col_in_940;
wire [2:0] col_in_941;
wire [2:0] col_in_942;
wire [2:0] col_in_943;
wire [2:0] col_in_944;
wire [2:0] col_in_945;
wire [2:0] col_in_946;
wire [2:0] col_in_947;
wire [2:0] col_in_948;
wire [2:0] col_in_949;
wire [2:0] col_in_950;
wire [2:0] col_in_951;
wire [2:0] col_in_952;
wire [2:0] col_in_953;
wire [2:0] col_in_954;
wire [2:0] col_in_955;
wire [2:0] col_in_956;
wire [2:0] col_in_957;
wire [2:0] col_in_958;
wire [2:0] col_in_959;
wire [2:0] col_in_960;
wire [2:0] col_in_961;
wire [2:0] col_in_962;
wire [2:0] col_in_963;
wire [2:0] col_in_964;
wire [2:0] col_in_965;
wire [2:0] col_in_966;
wire [2:0] col_in_967;
wire [2:0] col_in_968;
wire [2:0] col_in_969;
wire [2:0] col_in_970;
wire [2:0] col_in_971;
wire [2:0] col_in_972;
wire [2:0] col_in_973;
wire [2:0] col_in_974;
wire [2:0] col_in_975;
wire [2:0] col_in_976;
wire [2:0] col_in_977;
wire [2:0] col_in_978;
wire [2:0] col_in_979;
wire [2:0] col_in_980;
wire [2:0] col_in_981;
wire [2:0] col_in_982;
wire [2:0] col_in_983;
wire [2:0] col_in_984;
wire [2:0] col_in_985;
wire [2:0] col_in_986;
wire [2:0] col_in_987;
wire [2:0] col_in_988;
wire [2:0] col_in_989;
wire [2:0] col_in_990;
wire [2:0] col_in_991;
wire [2:0] col_in_992;
wire [2:0] col_in_993;
wire [2:0] col_in_994;
wire [2:0] col_in_995;
wire [2:0] col_in_996;
wire [2:0] col_in_997;
wire [2:0] col_in_998;
wire [2:0] col_in_999;
wire [2:0] col_in_1000;
wire [2:0] col_in_1001;
wire [2:0] col_in_1002;
wire [2:0] col_in_1003;
wire [2:0] col_in_1004;
wire [2:0] col_in_1005;
wire [2:0] col_in_1006;
wire [2:0] col_in_1007;
wire [2:0] col_in_1008;
wire [2:0] col_in_1009;
wire [2:0] col_in_1010;
wire [2:0] col_in_1011;
wire [2:0] col_in_1012;
wire [2:0] col_in_1013;
wire [2:0] col_in_1014;
wire [2:0] col_in_1015;
wire [2:0] col_in_1016;
wire [2:0] col_in_1017;
wire [2:0] col_in_1018;
wire [2:0] col_in_1019;
wire [2:0] col_in_1020;
wire [2:0] col_in_1021;
wire [2:0] col_in_1022;
wire [2:0] col_in_1023;


assign col_in_0 = {row_in_0[0],row_in_1[0],row_in_2[0]};
assign col_in_1 = {row_in_0[1],row_in_1[1],row_in_2[1]};
assign col_in_2 = {row_in_0[2],row_in_1[2],row_in_2[2]};
assign col_in_3 = {row_in_0[3],row_in_1[3],row_in_2[3]};
assign col_in_4 = {row_in_0[4],row_in_1[4],row_in_2[4]};
assign col_in_5 = {row_in_0[5],row_in_1[5],row_in_2[5]};
assign col_in_6 = {row_in_0[6],row_in_1[6],row_in_2[6]};
assign col_in_7 = {row_in_0[7],row_in_1[7],row_in_2[7]};
assign col_in_8 = {row_in_0[8],row_in_1[8],row_in_2[8]};
assign col_in_9 = {row_in_0[9],row_in_1[9],row_in_2[9]};
assign col_in_10 = {row_in_0[10],row_in_1[10],row_in_2[10]};
assign col_in_11 = {row_in_0[11],row_in_1[11],row_in_2[11]};
assign col_in_12 = {row_in_0[12],row_in_1[12],row_in_2[12]};
assign col_in_13 = {row_in_0[13],row_in_1[13],row_in_2[13]};
assign col_in_14 = {row_in_0[14],row_in_1[14],row_in_2[14]};
assign col_in_15 = {row_in_0[15],row_in_1[15],row_in_2[15]};
assign col_in_16 = {row_in_0[16],row_in_1[16],row_in_2[16]};
assign col_in_17 = {row_in_0[17],row_in_1[17],row_in_2[17]};
assign col_in_18 = {row_in_0[18],row_in_1[18],row_in_2[18]};
assign col_in_19 = {row_in_0[19],row_in_1[19],row_in_2[19]};
assign col_in_20 = {row_in_0[20],row_in_1[20],row_in_2[20]};
assign col_in_21 = {row_in_0[21],row_in_1[21],row_in_2[21]};
assign col_in_22 = {row_in_0[22],row_in_1[22],row_in_2[22]};
assign col_in_23 = {row_in_0[23],row_in_1[23],row_in_2[23]};
assign col_in_24 = {row_in_0[24],row_in_1[24],row_in_2[24]};
assign col_in_25 = {row_in_0[25],row_in_1[25],row_in_2[25]};
assign col_in_26 = {row_in_0[26],row_in_1[26],row_in_2[26]};
assign col_in_27 = {row_in_0[27],row_in_1[27],row_in_2[27]};
assign col_in_28 = {row_in_0[28],row_in_1[28],row_in_2[28]};
assign col_in_29 = {row_in_0[29],row_in_1[29],row_in_2[29]};
assign col_in_30 = {row_in_0[30],row_in_1[30],row_in_2[30]};
assign col_in_31 = {row_in_0[31],row_in_1[31],row_in_2[31]};
assign col_in_32 = {row_in_0[32],row_in_1[32],row_in_2[32]};
assign col_in_33 = {row_in_0[33],row_in_1[33],row_in_2[33]};
assign col_in_34 = {row_in_0[34],row_in_1[34],row_in_2[34]};
assign col_in_35 = {row_in_0[35],row_in_1[35],row_in_2[35]};
assign col_in_36 = {row_in_0[36],row_in_1[36],row_in_2[36]};
assign col_in_37 = {row_in_0[37],row_in_1[37],row_in_2[37]};
assign col_in_38 = {row_in_0[38],row_in_1[38],row_in_2[38]};
assign col_in_39 = {row_in_0[39],row_in_1[39],row_in_2[39]};
assign col_in_40 = {row_in_0[40],row_in_1[40],row_in_2[40]};
assign col_in_41 = {row_in_0[41],row_in_1[41],row_in_2[41]};
assign col_in_42 = {row_in_0[42],row_in_1[42],row_in_2[42]};
assign col_in_43 = {row_in_0[43],row_in_1[43],row_in_2[43]};
assign col_in_44 = {row_in_0[44],row_in_1[44],row_in_2[44]};
assign col_in_45 = {row_in_0[45],row_in_1[45],row_in_2[45]};
assign col_in_46 = {row_in_0[46],row_in_1[46],row_in_2[46]};
assign col_in_47 = {row_in_0[47],row_in_1[47],row_in_2[47]};
assign col_in_48 = {row_in_0[48],row_in_1[48],row_in_2[48]};
assign col_in_49 = {row_in_0[49],row_in_1[49],row_in_2[49]};
assign col_in_50 = {row_in_0[50],row_in_1[50],row_in_2[50]};
assign col_in_51 = {row_in_0[51],row_in_1[51],row_in_2[51]};
assign col_in_52 = {row_in_0[52],row_in_1[52],row_in_2[52]};
assign col_in_53 = {row_in_0[53],row_in_1[53],row_in_2[53]};
assign col_in_54 = {row_in_0[54],row_in_1[54],row_in_2[54]};
assign col_in_55 = {row_in_0[55],row_in_1[55],row_in_2[55]};
assign col_in_56 = {row_in_0[56],row_in_1[56],row_in_2[56]};
assign col_in_57 = {row_in_0[57],row_in_1[57],row_in_2[57]};
assign col_in_58 = {row_in_0[58],row_in_1[58],row_in_2[58]};
assign col_in_59 = {row_in_0[59],row_in_1[59],row_in_2[59]};
assign col_in_60 = {row_in_0[60],row_in_1[60],row_in_2[60]};
assign col_in_61 = {row_in_0[61],row_in_1[61],row_in_2[61]};
assign col_in_62 = {row_in_0[62],row_in_1[62],row_in_2[62]};
assign col_in_63 = {row_in_0[63],row_in_1[63],row_in_2[63]};
assign col_in_64 = {row_in_0[64],row_in_1[64],row_in_2[64]};
assign col_in_65 = {row_in_0[65],row_in_1[65],row_in_2[65]};
assign col_in_66 = {row_in_0[66],row_in_1[66],row_in_2[66]};
assign col_in_67 = {row_in_0[67],row_in_1[67],row_in_2[67]};
assign col_in_68 = {row_in_0[68],row_in_1[68],row_in_2[68]};
assign col_in_69 = {row_in_0[69],row_in_1[69],row_in_2[69]};
assign col_in_70 = {row_in_0[70],row_in_1[70],row_in_2[70]};
assign col_in_71 = {row_in_0[71],row_in_1[71],row_in_2[71]};
assign col_in_72 = {row_in_0[72],row_in_1[72],row_in_2[72]};
assign col_in_73 = {row_in_0[73],row_in_1[73],row_in_2[73]};
assign col_in_74 = {row_in_0[74],row_in_1[74],row_in_2[74]};
assign col_in_75 = {row_in_0[75],row_in_1[75],row_in_2[75]};
assign col_in_76 = {row_in_0[76],row_in_1[76],row_in_2[76]};
assign col_in_77 = {row_in_0[77],row_in_1[77],row_in_2[77]};
assign col_in_78 = {row_in_0[78],row_in_1[78],row_in_2[78]};
assign col_in_79 = {row_in_0[79],row_in_1[79],row_in_2[79]};
assign col_in_80 = {row_in_0[80],row_in_1[80],row_in_2[80]};
assign col_in_81 = {row_in_0[81],row_in_1[81],row_in_2[81]};
assign col_in_82 = {row_in_0[82],row_in_1[82],row_in_2[82]};
assign col_in_83 = {row_in_0[83],row_in_1[83],row_in_2[83]};
assign col_in_84 = {row_in_0[84],row_in_1[84],row_in_2[84]};
assign col_in_85 = {row_in_0[85],row_in_1[85],row_in_2[85]};
assign col_in_86 = {row_in_0[86],row_in_1[86],row_in_2[86]};
assign col_in_87 = {row_in_0[87],row_in_1[87],row_in_2[87]};
assign col_in_88 = {row_in_0[88],row_in_1[88],row_in_2[88]};
assign col_in_89 = {row_in_0[89],row_in_1[89],row_in_2[89]};
assign col_in_90 = {row_in_0[90],row_in_1[90],row_in_2[90]};
assign col_in_91 = {row_in_0[91],row_in_1[91],row_in_2[91]};
assign col_in_92 = {row_in_0[92],row_in_1[92],row_in_2[92]};
assign col_in_93 = {row_in_0[93],row_in_1[93],row_in_2[93]};
assign col_in_94 = {row_in_0[94],row_in_1[94],row_in_2[94]};
assign col_in_95 = {row_in_0[95],row_in_1[95],row_in_2[95]};
assign col_in_96 = {row_in_0[96],row_in_1[96],row_in_2[96]};
assign col_in_97 = {row_in_0[97],row_in_1[97],row_in_2[97]};
assign col_in_98 = {row_in_0[98],row_in_1[98],row_in_2[98]};
assign col_in_99 = {row_in_0[99],row_in_1[99],row_in_2[99]};
assign col_in_100 = {row_in_0[100],row_in_1[100],row_in_2[100]};
assign col_in_101 = {row_in_0[101],row_in_1[101],row_in_2[101]};
assign col_in_102 = {row_in_0[102],row_in_1[102],row_in_2[102]};
assign col_in_103 = {row_in_0[103],row_in_1[103],row_in_2[103]};
assign col_in_104 = {row_in_0[104],row_in_1[104],row_in_2[104]};
assign col_in_105 = {row_in_0[105],row_in_1[105],row_in_2[105]};
assign col_in_106 = {row_in_0[106],row_in_1[106],row_in_2[106]};
assign col_in_107 = {row_in_0[107],row_in_1[107],row_in_2[107]};
assign col_in_108 = {row_in_0[108],row_in_1[108],row_in_2[108]};
assign col_in_109 = {row_in_0[109],row_in_1[109],row_in_2[109]};
assign col_in_110 = {row_in_0[110],row_in_1[110],row_in_2[110]};
assign col_in_111 = {row_in_0[111],row_in_1[111],row_in_2[111]};
assign col_in_112 = {row_in_0[112],row_in_1[112],row_in_2[112]};
assign col_in_113 = {row_in_0[113],row_in_1[113],row_in_2[113]};
assign col_in_114 = {row_in_0[114],row_in_1[114],row_in_2[114]};
assign col_in_115 = {row_in_0[115],row_in_1[115],row_in_2[115]};
assign col_in_116 = {row_in_0[116],row_in_1[116],row_in_2[116]};
assign col_in_117 = {row_in_0[117],row_in_1[117],row_in_2[117]};
assign col_in_118 = {row_in_0[118],row_in_1[118],row_in_2[118]};
assign col_in_119 = {row_in_0[119],row_in_1[119],row_in_2[119]};
assign col_in_120 = {row_in_0[120],row_in_1[120],row_in_2[120]};
assign col_in_121 = {row_in_0[121],row_in_1[121],row_in_2[121]};
assign col_in_122 = {row_in_0[122],row_in_1[122],row_in_2[122]};
assign col_in_123 = {row_in_0[123],row_in_1[123],row_in_2[123]};
assign col_in_124 = {row_in_0[124],row_in_1[124],row_in_2[124]};
assign col_in_125 = {row_in_0[125],row_in_1[125],row_in_2[125]};
assign col_in_126 = {row_in_0[126],row_in_1[126],row_in_2[126]};
assign col_in_127 = {row_in_0[127],row_in_1[127],row_in_2[127]};
assign col_in_128 = {row_in_0[128],row_in_1[128],row_in_2[128]};
assign col_in_129 = {row_in_0[129],row_in_1[129],row_in_2[129]};
assign col_in_130 = {row_in_0[130],row_in_1[130],row_in_2[130]};
assign col_in_131 = {row_in_0[131],row_in_1[131],row_in_2[131]};
assign col_in_132 = {row_in_0[132],row_in_1[132],row_in_2[132]};
assign col_in_133 = {row_in_0[133],row_in_1[133],row_in_2[133]};
assign col_in_134 = {row_in_0[134],row_in_1[134],row_in_2[134]};
assign col_in_135 = {row_in_0[135],row_in_1[135],row_in_2[135]};
assign col_in_136 = {row_in_0[136],row_in_1[136],row_in_2[136]};
assign col_in_137 = {row_in_0[137],row_in_1[137],row_in_2[137]};
assign col_in_138 = {row_in_0[138],row_in_1[138],row_in_2[138]};
assign col_in_139 = {row_in_0[139],row_in_1[139],row_in_2[139]};
assign col_in_140 = {row_in_0[140],row_in_1[140],row_in_2[140]};
assign col_in_141 = {row_in_0[141],row_in_1[141],row_in_2[141]};
assign col_in_142 = {row_in_0[142],row_in_1[142],row_in_2[142]};
assign col_in_143 = {row_in_0[143],row_in_1[143],row_in_2[143]};
assign col_in_144 = {row_in_0[144],row_in_1[144],row_in_2[144]};
assign col_in_145 = {row_in_0[145],row_in_1[145],row_in_2[145]};
assign col_in_146 = {row_in_0[146],row_in_1[146],row_in_2[146]};
assign col_in_147 = {row_in_0[147],row_in_1[147],row_in_2[147]};
assign col_in_148 = {row_in_0[148],row_in_1[148],row_in_2[148]};
assign col_in_149 = {row_in_0[149],row_in_1[149],row_in_2[149]};
assign col_in_150 = {row_in_0[150],row_in_1[150],row_in_2[150]};
assign col_in_151 = {row_in_0[151],row_in_1[151],row_in_2[151]};
assign col_in_152 = {row_in_0[152],row_in_1[152],row_in_2[152]};
assign col_in_153 = {row_in_0[153],row_in_1[153],row_in_2[153]};
assign col_in_154 = {row_in_0[154],row_in_1[154],row_in_2[154]};
assign col_in_155 = {row_in_0[155],row_in_1[155],row_in_2[155]};
assign col_in_156 = {row_in_0[156],row_in_1[156],row_in_2[156]};
assign col_in_157 = {row_in_0[157],row_in_1[157],row_in_2[157]};
assign col_in_158 = {row_in_0[158],row_in_1[158],row_in_2[158]};
assign col_in_159 = {row_in_0[159],row_in_1[159],row_in_2[159]};
assign col_in_160 = {row_in_0[160],row_in_1[160],row_in_2[160]};
assign col_in_161 = {row_in_0[161],row_in_1[161],row_in_2[161]};
assign col_in_162 = {row_in_0[162],row_in_1[162],row_in_2[162]};
assign col_in_163 = {row_in_0[163],row_in_1[163],row_in_2[163]};
assign col_in_164 = {row_in_0[164],row_in_1[164],row_in_2[164]};
assign col_in_165 = {row_in_0[165],row_in_1[165],row_in_2[165]};
assign col_in_166 = {row_in_0[166],row_in_1[166],row_in_2[166]};
assign col_in_167 = {row_in_0[167],row_in_1[167],row_in_2[167]};
assign col_in_168 = {row_in_0[168],row_in_1[168],row_in_2[168]};
assign col_in_169 = {row_in_0[169],row_in_1[169],row_in_2[169]};
assign col_in_170 = {row_in_0[170],row_in_1[170],row_in_2[170]};
assign col_in_171 = {row_in_0[171],row_in_1[171],row_in_2[171]};
assign col_in_172 = {row_in_0[172],row_in_1[172],row_in_2[172]};
assign col_in_173 = {row_in_0[173],row_in_1[173],row_in_2[173]};
assign col_in_174 = {row_in_0[174],row_in_1[174],row_in_2[174]};
assign col_in_175 = {row_in_0[175],row_in_1[175],row_in_2[175]};
assign col_in_176 = {row_in_0[176],row_in_1[176],row_in_2[176]};
assign col_in_177 = {row_in_0[177],row_in_1[177],row_in_2[177]};
assign col_in_178 = {row_in_0[178],row_in_1[178],row_in_2[178]};
assign col_in_179 = {row_in_0[179],row_in_1[179],row_in_2[179]};
assign col_in_180 = {row_in_0[180],row_in_1[180],row_in_2[180]};
assign col_in_181 = {row_in_0[181],row_in_1[181],row_in_2[181]};
assign col_in_182 = {row_in_0[182],row_in_1[182],row_in_2[182]};
assign col_in_183 = {row_in_0[183],row_in_1[183],row_in_2[183]};
assign col_in_184 = {row_in_0[184],row_in_1[184],row_in_2[184]};
assign col_in_185 = {row_in_0[185],row_in_1[185],row_in_2[185]};
assign col_in_186 = {row_in_0[186],row_in_1[186],row_in_2[186]};
assign col_in_187 = {row_in_0[187],row_in_1[187],row_in_2[187]};
assign col_in_188 = {row_in_0[188],row_in_1[188],row_in_2[188]};
assign col_in_189 = {row_in_0[189],row_in_1[189],row_in_2[189]};
assign col_in_190 = {row_in_0[190],row_in_1[190],row_in_2[190]};
assign col_in_191 = {row_in_0[191],row_in_1[191],row_in_2[191]};
assign col_in_192 = {row_in_0[192],row_in_1[192],row_in_2[192]};
assign col_in_193 = {row_in_0[193],row_in_1[193],row_in_2[193]};
assign col_in_194 = {row_in_0[194],row_in_1[194],row_in_2[194]};
assign col_in_195 = {row_in_0[195],row_in_1[195],row_in_2[195]};
assign col_in_196 = {row_in_0[196],row_in_1[196],row_in_2[196]};
assign col_in_197 = {row_in_0[197],row_in_1[197],row_in_2[197]};
assign col_in_198 = {row_in_0[198],row_in_1[198],row_in_2[198]};
assign col_in_199 = {row_in_0[199],row_in_1[199],row_in_2[199]};
assign col_in_200 = {row_in_0[200],row_in_1[200],row_in_2[200]};
assign col_in_201 = {row_in_0[201],row_in_1[201],row_in_2[201]};
assign col_in_202 = {row_in_0[202],row_in_1[202],row_in_2[202]};
assign col_in_203 = {row_in_0[203],row_in_1[203],row_in_2[203]};
assign col_in_204 = {row_in_0[204],row_in_1[204],row_in_2[204]};
assign col_in_205 = {row_in_0[205],row_in_1[205],row_in_2[205]};
assign col_in_206 = {row_in_0[206],row_in_1[206],row_in_2[206]};
assign col_in_207 = {row_in_0[207],row_in_1[207],row_in_2[207]};
assign col_in_208 = {row_in_0[208],row_in_1[208],row_in_2[208]};
assign col_in_209 = {row_in_0[209],row_in_1[209],row_in_2[209]};
assign col_in_210 = {row_in_0[210],row_in_1[210],row_in_2[210]};
assign col_in_211 = {row_in_0[211],row_in_1[211],row_in_2[211]};
assign col_in_212 = {row_in_0[212],row_in_1[212],row_in_2[212]};
assign col_in_213 = {row_in_0[213],row_in_1[213],row_in_2[213]};
assign col_in_214 = {row_in_0[214],row_in_1[214],row_in_2[214]};
assign col_in_215 = {row_in_0[215],row_in_1[215],row_in_2[215]};
assign col_in_216 = {row_in_0[216],row_in_1[216],row_in_2[216]};
assign col_in_217 = {row_in_0[217],row_in_1[217],row_in_2[217]};
assign col_in_218 = {row_in_0[218],row_in_1[218],row_in_2[218]};
assign col_in_219 = {row_in_0[219],row_in_1[219],row_in_2[219]};
assign col_in_220 = {row_in_0[220],row_in_1[220],row_in_2[220]};
assign col_in_221 = {row_in_0[221],row_in_1[221],row_in_2[221]};
assign col_in_222 = {row_in_0[222],row_in_1[222],row_in_2[222]};
assign col_in_223 = {row_in_0[223],row_in_1[223],row_in_2[223]};
assign col_in_224 = {row_in_0[224],row_in_1[224],row_in_2[224]};
assign col_in_225 = {row_in_0[225],row_in_1[225],row_in_2[225]};
assign col_in_226 = {row_in_0[226],row_in_1[226],row_in_2[226]};
assign col_in_227 = {row_in_0[227],row_in_1[227],row_in_2[227]};
assign col_in_228 = {row_in_0[228],row_in_1[228],row_in_2[228]};
assign col_in_229 = {row_in_0[229],row_in_1[229],row_in_2[229]};
assign col_in_230 = {row_in_0[230],row_in_1[230],row_in_2[230]};
assign col_in_231 = {row_in_0[231],row_in_1[231],row_in_2[231]};
assign col_in_232 = {row_in_0[232],row_in_1[232],row_in_2[232]};
assign col_in_233 = {row_in_0[233],row_in_1[233],row_in_2[233]};
assign col_in_234 = {row_in_0[234],row_in_1[234],row_in_2[234]};
assign col_in_235 = {row_in_0[235],row_in_1[235],row_in_2[235]};
assign col_in_236 = {row_in_0[236],row_in_1[236],row_in_2[236]};
assign col_in_237 = {row_in_0[237],row_in_1[237],row_in_2[237]};
assign col_in_238 = {row_in_0[238],row_in_1[238],row_in_2[238]};
assign col_in_239 = {row_in_0[239],row_in_1[239],row_in_2[239]};
assign col_in_240 = {row_in_0[240],row_in_1[240],row_in_2[240]};
assign col_in_241 = {row_in_0[241],row_in_1[241],row_in_2[241]};
assign col_in_242 = {row_in_0[242],row_in_1[242],row_in_2[242]};
assign col_in_243 = {row_in_0[243],row_in_1[243],row_in_2[243]};
assign col_in_244 = {row_in_0[244],row_in_1[244],row_in_2[244]};
assign col_in_245 = {row_in_0[245],row_in_1[245],row_in_2[245]};
assign col_in_246 = {row_in_0[246],row_in_1[246],row_in_2[246]};
assign col_in_247 = {row_in_0[247],row_in_1[247],row_in_2[247]};
assign col_in_248 = {row_in_0[248],row_in_1[248],row_in_2[248]};
assign col_in_249 = {row_in_0[249],row_in_1[249],row_in_2[249]};
assign col_in_250 = {row_in_0[250],row_in_1[250],row_in_2[250]};
assign col_in_251 = {row_in_0[251],row_in_1[251],row_in_2[251]};
assign col_in_252 = {row_in_0[252],row_in_1[252],row_in_2[252]};
assign col_in_253 = {row_in_0[253],row_in_1[253],row_in_2[253]};
assign col_in_254 = {row_in_0[254],row_in_1[254],row_in_2[254]};
assign col_in_255 = {row_in_0[255],row_in_1[255],row_in_2[255]};
assign col_in_256 = {row_in_0[256],row_in_1[256],row_in_2[256]};
assign col_in_257 = {row_in_0[257],row_in_1[257],row_in_2[257]};
assign col_in_258 = {row_in_0[258],row_in_1[258],row_in_2[258]};
assign col_in_259 = {row_in_0[259],row_in_1[259],row_in_2[259]};
assign col_in_260 = {row_in_0[260],row_in_1[260],row_in_2[260]};
assign col_in_261 = {row_in_0[261],row_in_1[261],row_in_2[261]};
assign col_in_262 = {row_in_0[262],row_in_1[262],row_in_2[262]};
assign col_in_263 = {row_in_0[263],row_in_1[263],row_in_2[263]};
assign col_in_264 = {row_in_0[264],row_in_1[264],row_in_2[264]};
assign col_in_265 = {row_in_0[265],row_in_1[265],row_in_2[265]};
assign col_in_266 = {row_in_0[266],row_in_1[266],row_in_2[266]};
assign col_in_267 = {row_in_0[267],row_in_1[267],row_in_2[267]};
assign col_in_268 = {row_in_0[268],row_in_1[268],row_in_2[268]};
assign col_in_269 = {row_in_0[269],row_in_1[269],row_in_2[269]};
assign col_in_270 = {row_in_0[270],row_in_1[270],row_in_2[270]};
assign col_in_271 = {row_in_0[271],row_in_1[271],row_in_2[271]};
assign col_in_272 = {row_in_0[272],row_in_1[272],row_in_2[272]};
assign col_in_273 = {row_in_0[273],row_in_1[273],row_in_2[273]};
assign col_in_274 = {row_in_0[274],row_in_1[274],row_in_2[274]};
assign col_in_275 = {row_in_0[275],row_in_1[275],row_in_2[275]};
assign col_in_276 = {row_in_0[276],row_in_1[276],row_in_2[276]};
assign col_in_277 = {row_in_0[277],row_in_1[277],row_in_2[277]};
assign col_in_278 = {row_in_0[278],row_in_1[278],row_in_2[278]};
assign col_in_279 = {row_in_0[279],row_in_1[279],row_in_2[279]};
assign col_in_280 = {row_in_0[280],row_in_1[280],row_in_2[280]};
assign col_in_281 = {row_in_0[281],row_in_1[281],row_in_2[281]};
assign col_in_282 = {row_in_0[282],row_in_1[282],row_in_2[282]};
assign col_in_283 = {row_in_0[283],row_in_1[283],row_in_2[283]};
assign col_in_284 = {row_in_0[284],row_in_1[284],row_in_2[284]};
assign col_in_285 = {row_in_0[285],row_in_1[285],row_in_2[285]};
assign col_in_286 = {row_in_0[286],row_in_1[286],row_in_2[286]};
assign col_in_287 = {row_in_0[287],row_in_1[287],row_in_2[287]};
assign col_in_288 = {row_in_0[288],row_in_1[288],row_in_2[288]};
assign col_in_289 = {row_in_0[289],row_in_1[289],row_in_2[289]};
assign col_in_290 = {row_in_0[290],row_in_1[290],row_in_2[290]};
assign col_in_291 = {row_in_0[291],row_in_1[291],row_in_2[291]};
assign col_in_292 = {row_in_0[292],row_in_1[292],row_in_2[292]};
assign col_in_293 = {row_in_0[293],row_in_1[293],row_in_2[293]};
assign col_in_294 = {row_in_0[294],row_in_1[294],row_in_2[294]};
assign col_in_295 = {row_in_0[295],row_in_1[295],row_in_2[295]};
assign col_in_296 = {row_in_0[296],row_in_1[296],row_in_2[296]};
assign col_in_297 = {row_in_0[297],row_in_1[297],row_in_2[297]};
assign col_in_298 = {row_in_0[298],row_in_1[298],row_in_2[298]};
assign col_in_299 = {row_in_0[299],row_in_1[299],row_in_2[299]};
assign col_in_300 = {row_in_0[300],row_in_1[300],row_in_2[300]};
assign col_in_301 = {row_in_0[301],row_in_1[301],row_in_2[301]};
assign col_in_302 = {row_in_0[302],row_in_1[302],row_in_2[302]};
assign col_in_303 = {row_in_0[303],row_in_1[303],row_in_2[303]};
assign col_in_304 = {row_in_0[304],row_in_1[304],row_in_2[304]};
assign col_in_305 = {row_in_0[305],row_in_1[305],row_in_2[305]};
assign col_in_306 = {row_in_0[306],row_in_1[306],row_in_2[306]};
assign col_in_307 = {row_in_0[307],row_in_1[307],row_in_2[307]};
assign col_in_308 = {row_in_0[308],row_in_1[308],row_in_2[308]};
assign col_in_309 = {row_in_0[309],row_in_1[309],row_in_2[309]};
assign col_in_310 = {row_in_0[310],row_in_1[310],row_in_2[310]};
assign col_in_311 = {row_in_0[311],row_in_1[311],row_in_2[311]};
assign col_in_312 = {row_in_0[312],row_in_1[312],row_in_2[312]};
assign col_in_313 = {row_in_0[313],row_in_1[313],row_in_2[313]};
assign col_in_314 = {row_in_0[314],row_in_1[314],row_in_2[314]};
assign col_in_315 = {row_in_0[315],row_in_1[315],row_in_2[315]};
assign col_in_316 = {row_in_0[316],row_in_1[316],row_in_2[316]};
assign col_in_317 = {row_in_0[317],row_in_1[317],row_in_2[317]};
assign col_in_318 = {row_in_0[318],row_in_1[318],row_in_2[318]};
assign col_in_319 = {row_in_0[319],row_in_1[319],row_in_2[319]};
assign col_in_320 = {row_in_0[320],row_in_1[320],row_in_2[320]};
assign col_in_321 = {row_in_0[321],row_in_1[321],row_in_2[321]};
assign col_in_322 = {row_in_0[322],row_in_1[322],row_in_2[322]};
assign col_in_323 = {row_in_0[323],row_in_1[323],row_in_2[323]};
assign col_in_324 = {row_in_0[324],row_in_1[324],row_in_2[324]};
assign col_in_325 = {row_in_0[325],row_in_1[325],row_in_2[325]};
assign col_in_326 = {row_in_0[326],row_in_1[326],row_in_2[326]};
assign col_in_327 = {row_in_0[327],row_in_1[327],row_in_2[327]};
assign col_in_328 = {row_in_0[328],row_in_1[328],row_in_2[328]};
assign col_in_329 = {row_in_0[329],row_in_1[329],row_in_2[329]};
assign col_in_330 = {row_in_0[330],row_in_1[330],row_in_2[330]};
assign col_in_331 = {row_in_0[331],row_in_1[331],row_in_2[331]};
assign col_in_332 = {row_in_0[332],row_in_1[332],row_in_2[332]};
assign col_in_333 = {row_in_0[333],row_in_1[333],row_in_2[333]};
assign col_in_334 = {row_in_0[334],row_in_1[334],row_in_2[334]};
assign col_in_335 = {row_in_0[335],row_in_1[335],row_in_2[335]};
assign col_in_336 = {row_in_0[336],row_in_1[336],row_in_2[336]};
assign col_in_337 = {row_in_0[337],row_in_1[337],row_in_2[337]};
assign col_in_338 = {row_in_0[338],row_in_1[338],row_in_2[338]};
assign col_in_339 = {row_in_0[339],row_in_1[339],row_in_2[339]};
assign col_in_340 = {row_in_0[340],row_in_1[340],row_in_2[340]};
assign col_in_341 = {row_in_0[341],row_in_1[341],row_in_2[341]};
assign col_in_342 = {row_in_0[342],row_in_1[342],row_in_2[342]};
assign col_in_343 = {row_in_0[343],row_in_1[343],row_in_2[343]};
assign col_in_344 = {row_in_0[344],row_in_1[344],row_in_2[344]};
assign col_in_345 = {row_in_0[345],row_in_1[345],row_in_2[345]};
assign col_in_346 = {row_in_0[346],row_in_1[346],row_in_2[346]};
assign col_in_347 = {row_in_0[347],row_in_1[347],row_in_2[347]};
assign col_in_348 = {row_in_0[348],row_in_1[348],row_in_2[348]};
assign col_in_349 = {row_in_0[349],row_in_1[349],row_in_2[349]};
assign col_in_350 = {row_in_0[350],row_in_1[350],row_in_2[350]};
assign col_in_351 = {row_in_0[351],row_in_1[351],row_in_2[351]};
assign col_in_352 = {row_in_0[352],row_in_1[352],row_in_2[352]};
assign col_in_353 = {row_in_0[353],row_in_1[353],row_in_2[353]};
assign col_in_354 = {row_in_0[354],row_in_1[354],row_in_2[354]};
assign col_in_355 = {row_in_0[355],row_in_1[355],row_in_2[355]};
assign col_in_356 = {row_in_0[356],row_in_1[356],row_in_2[356]};
assign col_in_357 = {row_in_0[357],row_in_1[357],row_in_2[357]};
assign col_in_358 = {row_in_0[358],row_in_1[358],row_in_2[358]};
assign col_in_359 = {row_in_0[359],row_in_1[359],row_in_2[359]};
assign col_in_360 = {row_in_0[360],row_in_1[360],row_in_2[360]};
assign col_in_361 = {row_in_0[361],row_in_1[361],row_in_2[361]};
assign col_in_362 = {row_in_0[362],row_in_1[362],row_in_2[362]};
assign col_in_363 = {row_in_0[363],row_in_1[363],row_in_2[363]};
assign col_in_364 = {row_in_0[364],row_in_1[364],row_in_2[364]};
assign col_in_365 = {row_in_0[365],row_in_1[365],row_in_2[365]};
assign col_in_366 = {row_in_0[366],row_in_1[366],row_in_2[366]};
assign col_in_367 = {row_in_0[367],row_in_1[367],row_in_2[367]};
assign col_in_368 = {row_in_0[368],row_in_1[368],row_in_2[368]};
assign col_in_369 = {row_in_0[369],row_in_1[369],row_in_2[369]};
assign col_in_370 = {row_in_0[370],row_in_1[370],row_in_2[370]};
assign col_in_371 = {row_in_0[371],row_in_1[371],row_in_2[371]};
assign col_in_372 = {row_in_0[372],row_in_1[372],row_in_2[372]};
assign col_in_373 = {row_in_0[373],row_in_1[373],row_in_2[373]};
assign col_in_374 = {row_in_0[374],row_in_1[374],row_in_2[374]};
assign col_in_375 = {row_in_0[375],row_in_1[375],row_in_2[375]};
assign col_in_376 = {row_in_0[376],row_in_1[376],row_in_2[376]};
assign col_in_377 = {row_in_0[377],row_in_1[377],row_in_2[377]};
assign col_in_378 = {row_in_0[378],row_in_1[378],row_in_2[378]};
assign col_in_379 = {row_in_0[379],row_in_1[379],row_in_2[379]};
assign col_in_380 = {row_in_0[380],row_in_1[380],row_in_2[380]};
assign col_in_381 = {row_in_0[381],row_in_1[381],row_in_2[381]};
assign col_in_382 = {row_in_0[382],row_in_1[382],row_in_2[382]};
assign col_in_383 = {row_in_0[383],row_in_1[383],row_in_2[383]};
assign col_in_384 = {row_in_0[384],row_in_1[384],row_in_2[384]};
assign col_in_385 = {row_in_0[385],row_in_1[385],row_in_2[385]};
assign col_in_386 = {row_in_0[386],row_in_1[386],row_in_2[386]};
assign col_in_387 = {row_in_0[387],row_in_1[387],row_in_2[387]};
assign col_in_388 = {row_in_0[388],row_in_1[388],row_in_2[388]};
assign col_in_389 = {row_in_0[389],row_in_1[389],row_in_2[389]};
assign col_in_390 = {row_in_0[390],row_in_1[390],row_in_2[390]};
assign col_in_391 = {row_in_0[391],row_in_1[391],row_in_2[391]};
assign col_in_392 = {row_in_0[392],row_in_1[392],row_in_2[392]};
assign col_in_393 = {row_in_0[393],row_in_1[393],row_in_2[393]};
assign col_in_394 = {row_in_0[394],row_in_1[394],row_in_2[394]};
assign col_in_395 = {row_in_0[395],row_in_1[395],row_in_2[395]};
assign col_in_396 = {row_in_0[396],row_in_1[396],row_in_2[396]};
assign col_in_397 = {row_in_0[397],row_in_1[397],row_in_2[397]};
assign col_in_398 = {row_in_0[398],row_in_1[398],row_in_2[398]};
assign col_in_399 = {row_in_0[399],row_in_1[399],row_in_2[399]};
assign col_in_400 = {row_in_0[400],row_in_1[400],row_in_2[400]};
assign col_in_401 = {row_in_0[401],row_in_1[401],row_in_2[401]};
assign col_in_402 = {row_in_0[402],row_in_1[402],row_in_2[402]};
assign col_in_403 = {row_in_0[403],row_in_1[403],row_in_2[403]};
assign col_in_404 = {row_in_0[404],row_in_1[404],row_in_2[404]};
assign col_in_405 = {row_in_0[405],row_in_1[405],row_in_2[405]};
assign col_in_406 = {row_in_0[406],row_in_1[406],row_in_2[406]};
assign col_in_407 = {row_in_0[407],row_in_1[407],row_in_2[407]};
assign col_in_408 = {row_in_0[408],row_in_1[408],row_in_2[408]};
assign col_in_409 = {row_in_0[409],row_in_1[409],row_in_2[409]};
assign col_in_410 = {row_in_0[410],row_in_1[410],row_in_2[410]};
assign col_in_411 = {row_in_0[411],row_in_1[411],row_in_2[411]};
assign col_in_412 = {row_in_0[412],row_in_1[412],row_in_2[412]};
assign col_in_413 = {row_in_0[413],row_in_1[413],row_in_2[413]};
assign col_in_414 = {row_in_0[414],row_in_1[414],row_in_2[414]};
assign col_in_415 = {row_in_0[415],row_in_1[415],row_in_2[415]};
assign col_in_416 = {row_in_0[416],row_in_1[416],row_in_2[416]};
assign col_in_417 = {row_in_0[417],row_in_1[417],row_in_2[417]};
assign col_in_418 = {row_in_0[418],row_in_1[418],row_in_2[418]};
assign col_in_419 = {row_in_0[419],row_in_1[419],row_in_2[419]};
assign col_in_420 = {row_in_0[420],row_in_1[420],row_in_2[420]};
assign col_in_421 = {row_in_0[421],row_in_1[421],row_in_2[421]};
assign col_in_422 = {row_in_0[422],row_in_1[422],row_in_2[422]};
assign col_in_423 = {row_in_0[423],row_in_1[423],row_in_2[423]};
assign col_in_424 = {row_in_0[424],row_in_1[424],row_in_2[424]};
assign col_in_425 = {row_in_0[425],row_in_1[425],row_in_2[425]};
assign col_in_426 = {row_in_0[426],row_in_1[426],row_in_2[426]};
assign col_in_427 = {row_in_0[427],row_in_1[427],row_in_2[427]};
assign col_in_428 = {row_in_0[428],row_in_1[428],row_in_2[428]};
assign col_in_429 = {row_in_0[429],row_in_1[429],row_in_2[429]};
assign col_in_430 = {row_in_0[430],row_in_1[430],row_in_2[430]};
assign col_in_431 = {row_in_0[431],row_in_1[431],row_in_2[431]};
assign col_in_432 = {row_in_0[432],row_in_1[432],row_in_2[432]};
assign col_in_433 = {row_in_0[433],row_in_1[433],row_in_2[433]};
assign col_in_434 = {row_in_0[434],row_in_1[434],row_in_2[434]};
assign col_in_435 = {row_in_0[435],row_in_1[435],row_in_2[435]};
assign col_in_436 = {row_in_0[436],row_in_1[436],row_in_2[436]};
assign col_in_437 = {row_in_0[437],row_in_1[437],row_in_2[437]};
assign col_in_438 = {row_in_0[438],row_in_1[438],row_in_2[438]};
assign col_in_439 = {row_in_0[439],row_in_1[439],row_in_2[439]};
assign col_in_440 = {row_in_0[440],row_in_1[440],row_in_2[440]};
assign col_in_441 = {row_in_0[441],row_in_1[441],row_in_2[441]};
assign col_in_442 = {row_in_0[442],row_in_1[442],row_in_2[442]};
assign col_in_443 = {row_in_0[443],row_in_1[443],row_in_2[443]};
assign col_in_444 = {row_in_0[444],row_in_1[444],row_in_2[444]};
assign col_in_445 = {row_in_0[445],row_in_1[445],row_in_2[445]};
assign col_in_446 = {row_in_0[446],row_in_1[446],row_in_2[446]};
assign col_in_447 = {row_in_0[447],row_in_1[447],row_in_2[447]};
assign col_in_448 = {row_in_0[448],row_in_1[448],row_in_2[448]};
assign col_in_449 = {row_in_0[449],row_in_1[449],row_in_2[449]};
assign col_in_450 = {row_in_0[450],row_in_1[450],row_in_2[450]};
assign col_in_451 = {row_in_0[451],row_in_1[451],row_in_2[451]};
assign col_in_452 = {row_in_0[452],row_in_1[452],row_in_2[452]};
assign col_in_453 = {row_in_0[453],row_in_1[453],row_in_2[453]};
assign col_in_454 = {row_in_0[454],row_in_1[454],row_in_2[454]};
assign col_in_455 = {row_in_0[455],row_in_1[455],row_in_2[455]};
assign col_in_456 = {row_in_0[456],row_in_1[456],row_in_2[456]};
assign col_in_457 = {row_in_0[457],row_in_1[457],row_in_2[457]};
assign col_in_458 = {row_in_0[458],row_in_1[458],row_in_2[458]};
assign col_in_459 = {row_in_0[459],row_in_1[459],row_in_2[459]};
assign col_in_460 = {row_in_0[460],row_in_1[460],row_in_2[460]};
assign col_in_461 = {row_in_0[461],row_in_1[461],row_in_2[461]};
assign col_in_462 = {row_in_0[462],row_in_1[462],row_in_2[462]};
assign col_in_463 = {row_in_0[463],row_in_1[463],row_in_2[463]};
assign col_in_464 = {row_in_0[464],row_in_1[464],row_in_2[464]};
assign col_in_465 = {row_in_0[465],row_in_1[465],row_in_2[465]};
assign col_in_466 = {row_in_0[466],row_in_1[466],row_in_2[466]};
assign col_in_467 = {row_in_0[467],row_in_1[467],row_in_2[467]};
assign col_in_468 = {row_in_0[468],row_in_1[468],row_in_2[468]};
assign col_in_469 = {row_in_0[469],row_in_1[469],row_in_2[469]};
assign col_in_470 = {row_in_0[470],row_in_1[470],row_in_2[470]};
assign col_in_471 = {row_in_0[471],row_in_1[471],row_in_2[471]};
assign col_in_472 = {row_in_0[472],row_in_1[472],row_in_2[472]};
assign col_in_473 = {row_in_0[473],row_in_1[473],row_in_2[473]};
assign col_in_474 = {row_in_0[474],row_in_1[474],row_in_2[474]};
assign col_in_475 = {row_in_0[475],row_in_1[475],row_in_2[475]};
assign col_in_476 = {row_in_0[476],row_in_1[476],row_in_2[476]};
assign col_in_477 = {row_in_0[477],row_in_1[477],row_in_2[477]};
assign col_in_478 = {row_in_0[478],row_in_1[478],row_in_2[478]};
assign col_in_479 = {row_in_0[479],row_in_1[479],row_in_2[479]};
assign col_in_480 = {row_in_0[480],row_in_1[480],row_in_2[480]};
assign col_in_481 = {row_in_0[481],row_in_1[481],row_in_2[481]};
assign col_in_482 = {row_in_0[482],row_in_1[482],row_in_2[482]};
assign col_in_483 = {row_in_0[483],row_in_1[483],row_in_2[483]};
assign col_in_484 = {row_in_0[484],row_in_1[484],row_in_2[484]};
assign col_in_485 = {row_in_0[485],row_in_1[485],row_in_2[485]};
assign col_in_486 = {row_in_0[486],row_in_1[486],row_in_2[486]};
assign col_in_487 = {row_in_0[487],row_in_1[487],row_in_2[487]};
assign col_in_488 = {row_in_0[488],row_in_1[488],row_in_2[488]};
assign col_in_489 = {row_in_0[489],row_in_1[489],row_in_2[489]};
assign col_in_490 = {row_in_0[490],row_in_1[490],row_in_2[490]};
assign col_in_491 = {row_in_0[491],row_in_1[491],row_in_2[491]};
assign col_in_492 = {row_in_0[492],row_in_1[492],row_in_2[492]};
assign col_in_493 = {row_in_0[493],row_in_1[493],row_in_2[493]};
assign col_in_494 = {row_in_0[494],row_in_1[494],row_in_2[494]};
assign col_in_495 = {row_in_0[495],row_in_1[495],row_in_2[495]};
assign col_in_496 = {row_in_0[496],row_in_1[496],row_in_2[496]};
assign col_in_497 = {row_in_0[497],row_in_1[497],row_in_2[497]};
assign col_in_498 = {row_in_0[498],row_in_1[498],row_in_2[498]};
assign col_in_499 = {row_in_0[499],row_in_1[499],row_in_2[499]};
assign col_in_500 = {row_in_0[500],row_in_1[500],row_in_2[500]};
assign col_in_501 = {row_in_0[501],row_in_1[501],row_in_2[501]};
assign col_in_502 = {row_in_0[502],row_in_1[502],row_in_2[502]};
assign col_in_503 = {row_in_0[503],row_in_1[503],row_in_2[503]};
assign col_in_504 = {row_in_0[504],row_in_1[504],row_in_2[504]};
assign col_in_505 = {row_in_0[505],row_in_1[505],row_in_2[505]};
assign col_in_506 = {row_in_0[506],row_in_1[506],row_in_2[506]};
assign col_in_507 = {row_in_0[507],row_in_1[507],row_in_2[507]};
assign col_in_508 = {row_in_0[508],row_in_1[508],row_in_2[508]};
assign col_in_509 = {row_in_0[509],row_in_1[509],row_in_2[509]};
assign col_in_510 = {row_in_0[510],row_in_1[510],row_in_2[510]};
assign col_in_511 = {row_in_0[511],row_in_1[511],row_in_2[511]};
assign col_in_512 = {row_in_0[512],row_in_1[512],row_in_2[512]};
assign col_in_513 = {row_in_0[513],row_in_1[513],row_in_2[513]};
assign col_in_514 = {row_in_0[514],row_in_1[514],row_in_2[514]};
assign col_in_515 = {row_in_0[515],row_in_1[515],row_in_2[515]};
assign col_in_516 = {row_in_0[516],row_in_1[516],row_in_2[516]};
assign col_in_517 = {row_in_0[517],row_in_1[517],row_in_2[517]};
assign col_in_518 = {row_in_0[518],row_in_1[518],row_in_2[518]};
assign col_in_519 = {row_in_0[519],row_in_1[519],row_in_2[519]};
assign col_in_520 = {row_in_0[520],row_in_1[520],row_in_2[520]};
assign col_in_521 = {row_in_0[521],row_in_1[521],row_in_2[521]};
assign col_in_522 = {row_in_0[522],row_in_1[522],row_in_2[522]};
assign col_in_523 = {row_in_0[523],row_in_1[523],row_in_2[523]};
assign col_in_524 = {row_in_0[524],row_in_1[524],row_in_2[524]};
assign col_in_525 = {row_in_0[525],row_in_1[525],row_in_2[525]};
assign col_in_526 = {row_in_0[526],row_in_1[526],row_in_2[526]};
assign col_in_527 = {row_in_0[527],row_in_1[527],row_in_2[527]};
assign col_in_528 = {row_in_0[528],row_in_1[528],row_in_2[528]};
assign col_in_529 = {row_in_0[529],row_in_1[529],row_in_2[529]};
assign col_in_530 = {row_in_0[530],row_in_1[530],row_in_2[530]};
assign col_in_531 = {row_in_0[531],row_in_1[531],row_in_2[531]};
assign col_in_532 = {row_in_0[532],row_in_1[532],row_in_2[532]};
assign col_in_533 = {row_in_0[533],row_in_1[533],row_in_2[533]};
assign col_in_534 = {row_in_0[534],row_in_1[534],row_in_2[534]};
assign col_in_535 = {row_in_0[535],row_in_1[535],row_in_2[535]};
assign col_in_536 = {row_in_0[536],row_in_1[536],row_in_2[536]};
assign col_in_537 = {row_in_0[537],row_in_1[537],row_in_2[537]};
assign col_in_538 = {row_in_0[538],row_in_1[538],row_in_2[538]};
assign col_in_539 = {row_in_0[539],row_in_1[539],row_in_2[539]};
assign col_in_540 = {row_in_0[540],row_in_1[540],row_in_2[540]};
assign col_in_541 = {row_in_0[541],row_in_1[541],row_in_2[541]};
assign col_in_542 = {row_in_0[542],row_in_1[542],row_in_2[542]};
assign col_in_543 = {row_in_0[543],row_in_1[543],row_in_2[543]};
assign col_in_544 = {row_in_0[544],row_in_1[544],row_in_2[544]};
assign col_in_545 = {row_in_0[545],row_in_1[545],row_in_2[545]};
assign col_in_546 = {row_in_0[546],row_in_1[546],row_in_2[546]};
assign col_in_547 = {row_in_0[547],row_in_1[547],row_in_2[547]};
assign col_in_548 = {row_in_0[548],row_in_1[548],row_in_2[548]};
assign col_in_549 = {row_in_0[549],row_in_1[549],row_in_2[549]};
assign col_in_550 = {row_in_0[550],row_in_1[550],row_in_2[550]};
assign col_in_551 = {row_in_0[551],row_in_1[551],row_in_2[551]};
assign col_in_552 = {row_in_0[552],row_in_1[552],row_in_2[552]};
assign col_in_553 = {row_in_0[553],row_in_1[553],row_in_2[553]};
assign col_in_554 = {row_in_0[554],row_in_1[554],row_in_2[554]};
assign col_in_555 = {row_in_0[555],row_in_1[555],row_in_2[555]};
assign col_in_556 = {row_in_0[556],row_in_1[556],row_in_2[556]};
assign col_in_557 = {row_in_0[557],row_in_1[557],row_in_2[557]};
assign col_in_558 = {row_in_0[558],row_in_1[558],row_in_2[558]};
assign col_in_559 = {row_in_0[559],row_in_1[559],row_in_2[559]};
assign col_in_560 = {row_in_0[560],row_in_1[560],row_in_2[560]};
assign col_in_561 = {row_in_0[561],row_in_1[561],row_in_2[561]};
assign col_in_562 = {row_in_0[562],row_in_1[562],row_in_2[562]};
assign col_in_563 = {row_in_0[563],row_in_1[563],row_in_2[563]};
assign col_in_564 = {row_in_0[564],row_in_1[564],row_in_2[564]};
assign col_in_565 = {row_in_0[565],row_in_1[565],row_in_2[565]};
assign col_in_566 = {row_in_0[566],row_in_1[566],row_in_2[566]};
assign col_in_567 = {row_in_0[567],row_in_1[567],row_in_2[567]};
assign col_in_568 = {row_in_0[568],row_in_1[568],row_in_2[568]};
assign col_in_569 = {row_in_0[569],row_in_1[569],row_in_2[569]};
assign col_in_570 = {row_in_0[570],row_in_1[570],row_in_2[570]};
assign col_in_571 = {row_in_0[571],row_in_1[571],row_in_2[571]};
assign col_in_572 = {row_in_0[572],row_in_1[572],row_in_2[572]};
assign col_in_573 = {row_in_0[573],row_in_1[573],row_in_2[573]};
assign col_in_574 = {row_in_0[574],row_in_1[574],row_in_2[574]};
assign col_in_575 = {row_in_0[575],row_in_1[575],row_in_2[575]};
assign col_in_576 = {row_in_0[576],row_in_1[576],row_in_2[576]};
assign col_in_577 = {row_in_0[577],row_in_1[577],row_in_2[577]};
assign col_in_578 = {row_in_0[578],row_in_1[578],row_in_2[578]};
assign col_in_579 = {row_in_0[579],row_in_1[579],row_in_2[579]};
assign col_in_580 = {row_in_0[580],row_in_1[580],row_in_2[580]};
assign col_in_581 = {row_in_0[581],row_in_1[581],row_in_2[581]};
assign col_in_582 = {row_in_0[582],row_in_1[582],row_in_2[582]};
assign col_in_583 = {row_in_0[583],row_in_1[583],row_in_2[583]};
assign col_in_584 = {row_in_0[584],row_in_1[584],row_in_2[584]};
assign col_in_585 = {row_in_0[585],row_in_1[585],row_in_2[585]};
assign col_in_586 = {row_in_0[586],row_in_1[586],row_in_2[586]};
assign col_in_587 = {row_in_0[587],row_in_1[587],row_in_2[587]};
assign col_in_588 = {row_in_0[588],row_in_1[588],row_in_2[588]};
assign col_in_589 = {row_in_0[589],row_in_1[589],row_in_2[589]};
assign col_in_590 = {row_in_0[590],row_in_1[590],row_in_2[590]};
assign col_in_591 = {row_in_0[591],row_in_1[591],row_in_2[591]};
assign col_in_592 = {row_in_0[592],row_in_1[592],row_in_2[592]};
assign col_in_593 = {row_in_0[593],row_in_1[593],row_in_2[593]};
assign col_in_594 = {row_in_0[594],row_in_1[594],row_in_2[594]};
assign col_in_595 = {row_in_0[595],row_in_1[595],row_in_2[595]};
assign col_in_596 = {row_in_0[596],row_in_1[596],row_in_2[596]};
assign col_in_597 = {row_in_0[597],row_in_1[597],row_in_2[597]};
assign col_in_598 = {row_in_0[598],row_in_1[598],row_in_2[598]};
assign col_in_599 = {row_in_0[599],row_in_1[599],row_in_2[599]};
assign col_in_600 = {row_in_0[600],row_in_1[600],row_in_2[600]};
assign col_in_601 = {row_in_0[601],row_in_1[601],row_in_2[601]};
assign col_in_602 = {row_in_0[602],row_in_1[602],row_in_2[602]};
assign col_in_603 = {row_in_0[603],row_in_1[603],row_in_2[603]};
assign col_in_604 = {row_in_0[604],row_in_1[604],row_in_2[604]};
assign col_in_605 = {row_in_0[605],row_in_1[605],row_in_2[605]};
assign col_in_606 = {row_in_0[606],row_in_1[606],row_in_2[606]};
assign col_in_607 = {row_in_0[607],row_in_1[607],row_in_2[607]};
assign col_in_608 = {row_in_0[608],row_in_1[608],row_in_2[608]};
assign col_in_609 = {row_in_0[609],row_in_1[609],row_in_2[609]};
assign col_in_610 = {row_in_0[610],row_in_1[610],row_in_2[610]};
assign col_in_611 = {row_in_0[611],row_in_1[611],row_in_2[611]};
assign col_in_612 = {row_in_0[612],row_in_1[612],row_in_2[612]};
assign col_in_613 = {row_in_0[613],row_in_1[613],row_in_2[613]};
assign col_in_614 = {row_in_0[614],row_in_1[614],row_in_2[614]};
assign col_in_615 = {row_in_0[615],row_in_1[615],row_in_2[615]};
assign col_in_616 = {row_in_0[616],row_in_1[616],row_in_2[616]};
assign col_in_617 = {row_in_0[617],row_in_1[617],row_in_2[617]};
assign col_in_618 = {row_in_0[618],row_in_1[618],row_in_2[618]};
assign col_in_619 = {row_in_0[619],row_in_1[619],row_in_2[619]};
assign col_in_620 = {row_in_0[620],row_in_1[620],row_in_2[620]};
assign col_in_621 = {row_in_0[621],row_in_1[621],row_in_2[621]};
assign col_in_622 = {row_in_0[622],row_in_1[622],row_in_2[622]};
assign col_in_623 = {row_in_0[623],row_in_1[623],row_in_2[623]};
assign col_in_624 = {row_in_0[624],row_in_1[624],row_in_2[624]};
assign col_in_625 = {row_in_0[625],row_in_1[625],row_in_2[625]};
assign col_in_626 = {row_in_0[626],row_in_1[626],row_in_2[626]};
assign col_in_627 = {row_in_0[627],row_in_1[627],row_in_2[627]};
assign col_in_628 = {row_in_0[628],row_in_1[628],row_in_2[628]};
assign col_in_629 = {row_in_0[629],row_in_1[629],row_in_2[629]};
assign col_in_630 = {row_in_0[630],row_in_1[630],row_in_2[630]};
assign col_in_631 = {row_in_0[631],row_in_1[631],row_in_2[631]};
assign col_in_632 = {row_in_0[632],row_in_1[632],row_in_2[632]};
assign col_in_633 = {row_in_0[633],row_in_1[633],row_in_2[633]};
assign col_in_634 = {row_in_0[634],row_in_1[634],row_in_2[634]};
assign col_in_635 = {row_in_0[635],row_in_1[635],row_in_2[635]};
assign col_in_636 = {row_in_0[636],row_in_1[636],row_in_2[636]};
assign col_in_637 = {row_in_0[637],row_in_1[637],row_in_2[637]};
assign col_in_638 = {row_in_0[638],row_in_1[638],row_in_2[638]};
assign col_in_639 = {row_in_0[639],row_in_1[639],row_in_2[639]};
assign col_in_640 = {row_in_0[640],row_in_1[640],row_in_2[640]};
assign col_in_641 = {row_in_0[641],row_in_1[641],row_in_2[641]};
assign col_in_642 = {row_in_0[642],row_in_1[642],row_in_2[642]};
assign col_in_643 = {row_in_0[643],row_in_1[643],row_in_2[643]};
assign col_in_644 = {row_in_0[644],row_in_1[644],row_in_2[644]};
assign col_in_645 = {row_in_0[645],row_in_1[645],row_in_2[645]};
assign col_in_646 = {row_in_0[646],row_in_1[646],row_in_2[646]};
assign col_in_647 = {row_in_0[647],row_in_1[647],row_in_2[647]};
assign col_in_648 = {row_in_0[648],row_in_1[648],row_in_2[648]};
assign col_in_649 = {row_in_0[649],row_in_1[649],row_in_2[649]};
assign col_in_650 = {row_in_0[650],row_in_1[650],row_in_2[650]};
assign col_in_651 = {row_in_0[651],row_in_1[651],row_in_2[651]};
assign col_in_652 = {row_in_0[652],row_in_1[652],row_in_2[652]};
assign col_in_653 = {row_in_0[653],row_in_1[653],row_in_2[653]};
assign col_in_654 = {row_in_0[654],row_in_1[654],row_in_2[654]};
assign col_in_655 = {row_in_0[655],row_in_1[655],row_in_2[655]};
assign col_in_656 = {row_in_0[656],row_in_1[656],row_in_2[656]};
assign col_in_657 = {row_in_0[657],row_in_1[657],row_in_2[657]};
assign col_in_658 = {row_in_0[658],row_in_1[658],row_in_2[658]};
assign col_in_659 = {row_in_0[659],row_in_1[659],row_in_2[659]};
assign col_in_660 = {row_in_0[660],row_in_1[660],row_in_2[660]};
assign col_in_661 = {row_in_0[661],row_in_1[661],row_in_2[661]};
assign col_in_662 = {row_in_0[662],row_in_1[662],row_in_2[662]};
assign col_in_663 = {row_in_0[663],row_in_1[663],row_in_2[663]};
assign col_in_664 = {row_in_0[664],row_in_1[664],row_in_2[664]};
assign col_in_665 = {row_in_0[665],row_in_1[665],row_in_2[665]};
assign col_in_666 = {row_in_0[666],row_in_1[666],row_in_2[666]};
assign col_in_667 = {row_in_0[667],row_in_1[667],row_in_2[667]};
assign col_in_668 = {row_in_0[668],row_in_1[668],row_in_2[668]};
assign col_in_669 = {row_in_0[669],row_in_1[669],row_in_2[669]};
assign col_in_670 = {row_in_0[670],row_in_1[670],row_in_2[670]};
assign col_in_671 = {row_in_0[671],row_in_1[671],row_in_2[671]};
assign col_in_672 = {row_in_0[672],row_in_1[672],row_in_2[672]};
assign col_in_673 = {row_in_0[673],row_in_1[673],row_in_2[673]};
assign col_in_674 = {row_in_0[674],row_in_1[674],row_in_2[674]};
assign col_in_675 = {row_in_0[675],row_in_1[675],row_in_2[675]};
assign col_in_676 = {row_in_0[676],row_in_1[676],row_in_2[676]};
assign col_in_677 = {row_in_0[677],row_in_1[677],row_in_2[677]};
assign col_in_678 = {row_in_0[678],row_in_1[678],row_in_2[678]};
assign col_in_679 = {row_in_0[679],row_in_1[679],row_in_2[679]};
assign col_in_680 = {row_in_0[680],row_in_1[680],row_in_2[680]};
assign col_in_681 = {row_in_0[681],row_in_1[681],row_in_2[681]};
assign col_in_682 = {row_in_0[682],row_in_1[682],row_in_2[682]};
assign col_in_683 = {row_in_0[683],row_in_1[683],row_in_2[683]};
assign col_in_684 = {row_in_0[684],row_in_1[684],row_in_2[684]};
assign col_in_685 = {row_in_0[685],row_in_1[685],row_in_2[685]};
assign col_in_686 = {row_in_0[686],row_in_1[686],row_in_2[686]};
assign col_in_687 = {row_in_0[687],row_in_1[687],row_in_2[687]};
assign col_in_688 = {row_in_0[688],row_in_1[688],row_in_2[688]};
assign col_in_689 = {row_in_0[689],row_in_1[689],row_in_2[689]};
assign col_in_690 = {row_in_0[690],row_in_1[690],row_in_2[690]};
assign col_in_691 = {row_in_0[691],row_in_1[691],row_in_2[691]};
assign col_in_692 = {row_in_0[692],row_in_1[692],row_in_2[692]};
assign col_in_693 = {row_in_0[693],row_in_1[693],row_in_2[693]};
assign col_in_694 = {row_in_0[694],row_in_1[694],row_in_2[694]};
assign col_in_695 = {row_in_0[695],row_in_1[695],row_in_2[695]};
assign col_in_696 = {row_in_0[696],row_in_1[696],row_in_2[696]};
assign col_in_697 = {row_in_0[697],row_in_1[697],row_in_2[697]};
assign col_in_698 = {row_in_0[698],row_in_1[698],row_in_2[698]};
assign col_in_699 = {row_in_0[699],row_in_1[699],row_in_2[699]};
assign col_in_700 = {row_in_0[700],row_in_1[700],row_in_2[700]};
assign col_in_701 = {row_in_0[701],row_in_1[701],row_in_2[701]};
assign col_in_702 = {row_in_0[702],row_in_1[702],row_in_2[702]};
assign col_in_703 = {row_in_0[703],row_in_1[703],row_in_2[703]};
assign col_in_704 = {row_in_0[704],row_in_1[704],row_in_2[704]};
assign col_in_705 = {row_in_0[705],row_in_1[705],row_in_2[705]};
assign col_in_706 = {row_in_0[706],row_in_1[706],row_in_2[706]};
assign col_in_707 = {row_in_0[707],row_in_1[707],row_in_2[707]};
assign col_in_708 = {row_in_0[708],row_in_1[708],row_in_2[708]};
assign col_in_709 = {row_in_0[709],row_in_1[709],row_in_2[709]};
assign col_in_710 = {row_in_0[710],row_in_1[710],row_in_2[710]};
assign col_in_711 = {row_in_0[711],row_in_1[711],row_in_2[711]};
assign col_in_712 = {row_in_0[712],row_in_1[712],row_in_2[712]};
assign col_in_713 = {row_in_0[713],row_in_1[713],row_in_2[713]};
assign col_in_714 = {row_in_0[714],row_in_1[714],row_in_2[714]};
assign col_in_715 = {row_in_0[715],row_in_1[715],row_in_2[715]};
assign col_in_716 = {row_in_0[716],row_in_1[716],row_in_2[716]};
assign col_in_717 = {row_in_0[717],row_in_1[717],row_in_2[717]};
assign col_in_718 = {row_in_0[718],row_in_1[718],row_in_2[718]};
assign col_in_719 = {row_in_0[719],row_in_1[719],row_in_2[719]};
assign col_in_720 = {row_in_0[720],row_in_1[720],row_in_2[720]};
assign col_in_721 = {row_in_0[721],row_in_1[721],row_in_2[721]};
assign col_in_722 = {row_in_0[722],row_in_1[722],row_in_2[722]};
assign col_in_723 = {row_in_0[723],row_in_1[723],row_in_2[723]};
assign col_in_724 = {row_in_0[724],row_in_1[724],row_in_2[724]};
assign col_in_725 = {row_in_0[725],row_in_1[725],row_in_2[725]};
assign col_in_726 = {row_in_0[726],row_in_1[726],row_in_2[726]};
assign col_in_727 = {row_in_0[727],row_in_1[727],row_in_2[727]};
assign col_in_728 = {row_in_0[728],row_in_1[728],row_in_2[728]};
assign col_in_729 = {row_in_0[729],row_in_1[729],row_in_2[729]};
assign col_in_730 = {row_in_0[730],row_in_1[730],row_in_2[730]};
assign col_in_731 = {row_in_0[731],row_in_1[731],row_in_2[731]};
assign col_in_732 = {row_in_0[732],row_in_1[732],row_in_2[732]};
assign col_in_733 = {row_in_0[733],row_in_1[733],row_in_2[733]};
assign col_in_734 = {row_in_0[734],row_in_1[734],row_in_2[734]};
assign col_in_735 = {row_in_0[735],row_in_1[735],row_in_2[735]};
assign col_in_736 = {row_in_0[736],row_in_1[736],row_in_2[736]};
assign col_in_737 = {row_in_0[737],row_in_1[737],row_in_2[737]};
assign col_in_738 = {row_in_0[738],row_in_1[738],row_in_2[738]};
assign col_in_739 = {row_in_0[739],row_in_1[739],row_in_2[739]};
assign col_in_740 = {row_in_0[740],row_in_1[740],row_in_2[740]};
assign col_in_741 = {row_in_0[741],row_in_1[741],row_in_2[741]};
assign col_in_742 = {row_in_0[742],row_in_1[742],row_in_2[742]};
assign col_in_743 = {row_in_0[743],row_in_1[743],row_in_2[743]};
assign col_in_744 = {row_in_0[744],row_in_1[744],row_in_2[744]};
assign col_in_745 = {row_in_0[745],row_in_1[745],row_in_2[745]};
assign col_in_746 = {row_in_0[746],row_in_1[746],row_in_2[746]};
assign col_in_747 = {row_in_0[747],row_in_1[747],row_in_2[747]};
assign col_in_748 = {row_in_0[748],row_in_1[748],row_in_2[748]};
assign col_in_749 = {row_in_0[749],row_in_1[749],row_in_2[749]};
assign col_in_750 = {row_in_0[750],row_in_1[750],row_in_2[750]};
assign col_in_751 = {row_in_0[751],row_in_1[751],row_in_2[751]};
assign col_in_752 = {row_in_0[752],row_in_1[752],row_in_2[752]};
assign col_in_753 = {row_in_0[753],row_in_1[753],row_in_2[753]};
assign col_in_754 = {row_in_0[754],row_in_1[754],row_in_2[754]};
assign col_in_755 = {row_in_0[755],row_in_1[755],row_in_2[755]};
assign col_in_756 = {row_in_0[756],row_in_1[756],row_in_2[756]};
assign col_in_757 = {row_in_0[757],row_in_1[757],row_in_2[757]};
assign col_in_758 = {row_in_0[758],row_in_1[758],row_in_2[758]};
assign col_in_759 = {row_in_0[759],row_in_1[759],row_in_2[759]};
assign col_in_760 = {row_in_0[760],row_in_1[760],row_in_2[760]};
assign col_in_761 = {row_in_0[761],row_in_1[761],row_in_2[761]};
assign col_in_762 = {row_in_0[762],row_in_1[762],row_in_2[762]};
assign col_in_763 = {row_in_0[763],row_in_1[763],row_in_2[763]};
assign col_in_764 = {row_in_0[764],row_in_1[764],row_in_2[764]};
assign col_in_765 = {row_in_0[765],row_in_1[765],row_in_2[765]};
assign col_in_766 = {row_in_0[766],row_in_1[766],row_in_2[766]};
assign col_in_767 = {row_in_0[767],row_in_1[767],row_in_2[767]};
assign col_in_768 = {row_in_0[768],row_in_1[768],row_in_2[768]};
assign col_in_769 = {row_in_0[769],row_in_1[769],row_in_2[769]};
assign col_in_770 = {row_in_0[770],row_in_1[770],row_in_2[770]};
assign col_in_771 = {row_in_0[771],row_in_1[771],row_in_2[771]};
assign col_in_772 = {row_in_0[772],row_in_1[772],row_in_2[772]};
assign col_in_773 = {row_in_0[773],row_in_1[773],row_in_2[773]};
assign col_in_774 = {row_in_0[774],row_in_1[774],row_in_2[774]};
assign col_in_775 = {row_in_0[775],row_in_1[775],row_in_2[775]};
assign col_in_776 = {row_in_0[776],row_in_1[776],row_in_2[776]};
assign col_in_777 = {row_in_0[777],row_in_1[777],row_in_2[777]};
assign col_in_778 = {row_in_0[778],row_in_1[778],row_in_2[778]};
assign col_in_779 = {row_in_0[779],row_in_1[779],row_in_2[779]};
assign col_in_780 = {row_in_0[780],row_in_1[780],row_in_2[780]};
assign col_in_781 = {row_in_0[781],row_in_1[781],row_in_2[781]};
assign col_in_782 = {row_in_0[782],row_in_1[782],row_in_2[782]};
assign col_in_783 = {row_in_0[783],row_in_1[783],row_in_2[783]};
assign col_in_784 = {row_in_0[784],row_in_1[784],row_in_2[784]};
assign col_in_785 = {row_in_0[785],row_in_1[785],row_in_2[785]};
assign col_in_786 = {row_in_0[786],row_in_1[786],row_in_2[786]};
assign col_in_787 = {row_in_0[787],row_in_1[787],row_in_2[787]};
assign col_in_788 = {row_in_0[788],row_in_1[788],row_in_2[788]};
assign col_in_789 = {row_in_0[789],row_in_1[789],row_in_2[789]};
assign col_in_790 = {row_in_0[790],row_in_1[790],row_in_2[790]};
assign col_in_791 = {row_in_0[791],row_in_1[791],row_in_2[791]};
assign col_in_792 = {row_in_0[792],row_in_1[792],row_in_2[792]};
assign col_in_793 = {row_in_0[793],row_in_1[793],row_in_2[793]};
assign col_in_794 = {row_in_0[794],row_in_1[794],row_in_2[794]};
assign col_in_795 = {row_in_0[795],row_in_1[795],row_in_2[795]};
assign col_in_796 = {row_in_0[796],row_in_1[796],row_in_2[796]};
assign col_in_797 = {row_in_0[797],row_in_1[797],row_in_2[797]};
assign col_in_798 = {row_in_0[798],row_in_1[798],row_in_2[798]};
assign col_in_799 = {row_in_0[799],row_in_1[799],row_in_2[799]};
assign col_in_800 = {row_in_0[800],row_in_1[800],row_in_2[800]};
assign col_in_801 = {row_in_0[801],row_in_1[801],row_in_2[801]};
assign col_in_802 = {row_in_0[802],row_in_1[802],row_in_2[802]};
assign col_in_803 = {row_in_0[803],row_in_1[803],row_in_2[803]};
assign col_in_804 = {row_in_0[804],row_in_1[804],row_in_2[804]};
assign col_in_805 = {row_in_0[805],row_in_1[805],row_in_2[805]};
assign col_in_806 = {row_in_0[806],row_in_1[806],row_in_2[806]};
assign col_in_807 = {row_in_0[807],row_in_1[807],row_in_2[807]};
assign col_in_808 = {row_in_0[808],row_in_1[808],row_in_2[808]};
assign col_in_809 = {row_in_0[809],row_in_1[809],row_in_2[809]};
assign col_in_810 = {row_in_0[810],row_in_1[810],row_in_2[810]};
assign col_in_811 = {row_in_0[811],row_in_1[811],row_in_2[811]};
assign col_in_812 = {row_in_0[812],row_in_1[812],row_in_2[812]};
assign col_in_813 = {row_in_0[813],row_in_1[813],row_in_2[813]};
assign col_in_814 = {row_in_0[814],row_in_1[814],row_in_2[814]};
assign col_in_815 = {row_in_0[815],row_in_1[815],row_in_2[815]};
assign col_in_816 = {row_in_0[816],row_in_1[816],row_in_2[816]};
assign col_in_817 = {row_in_0[817],row_in_1[817],row_in_2[817]};
assign col_in_818 = {row_in_0[818],row_in_1[818],row_in_2[818]};
assign col_in_819 = {row_in_0[819],row_in_1[819],row_in_2[819]};
assign col_in_820 = {row_in_0[820],row_in_1[820],row_in_2[820]};
assign col_in_821 = {row_in_0[821],row_in_1[821],row_in_2[821]};
assign col_in_822 = {row_in_0[822],row_in_1[822],row_in_2[822]};
assign col_in_823 = {row_in_0[823],row_in_1[823],row_in_2[823]};
assign col_in_824 = {row_in_0[824],row_in_1[824],row_in_2[824]};
assign col_in_825 = {row_in_0[825],row_in_1[825],row_in_2[825]};
assign col_in_826 = {row_in_0[826],row_in_1[826],row_in_2[826]};
assign col_in_827 = {row_in_0[827],row_in_1[827],row_in_2[827]};
assign col_in_828 = {row_in_0[828],row_in_1[828],row_in_2[828]};
assign col_in_829 = {row_in_0[829],row_in_1[829],row_in_2[829]};
assign col_in_830 = {row_in_0[830],row_in_1[830],row_in_2[830]};
assign col_in_831 = {row_in_0[831],row_in_1[831],row_in_2[831]};
assign col_in_832 = {row_in_0[832],row_in_1[832],row_in_2[832]};
assign col_in_833 = {row_in_0[833],row_in_1[833],row_in_2[833]};
assign col_in_834 = {row_in_0[834],row_in_1[834],row_in_2[834]};
assign col_in_835 = {row_in_0[835],row_in_1[835],row_in_2[835]};
assign col_in_836 = {row_in_0[836],row_in_1[836],row_in_2[836]};
assign col_in_837 = {row_in_0[837],row_in_1[837],row_in_2[837]};
assign col_in_838 = {row_in_0[838],row_in_1[838],row_in_2[838]};
assign col_in_839 = {row_in_0[839],row_in_1[839],row_in_2[839]};
assign col_in_840 = {row_in_0[840],row_in_1[840],row_in_2[840]};
assign col_in_841 = {row_in_0[841],row_in_1[841],row_in_2[841]};
assign col_in_842 = {row_in_0[842],row_in_1[842],row_in_2[842]};
assign col_in_843 = {row_in_0[843],row_in_1[843],row_in_2[843]};
assign col_in_844 = {row_in_0[844],row_in_1[844],row_in_2[844]};
assign col_in_845 = {row_in_0[845],row_in_1[845],row_in_2[845]};
assign col_in_846 = {row_in_0[846],row_in_1[846],row_in_2[846]};
assign col_in_847 = {row_in_0[847],row_in_1[847],row_in_2[847]};
assign col_in_848 = {row_in_0[848],row_in_1[848],row_in_2[848]};
assign col_in_849 = {row_in_0[849],row_in_1[849],row_in_2[849]};
assign col_in_850 = {row_in_0[850],row_in_1[850],row_in_2[850]};
assign col_in_851 = {row_in_0[851],row_in_1[851],row_in_2[851]};
assign col_in_852 = {row_in_0[852],row_in_1[852],row_in_2[852]};
assign col_in_853 = {row_in_0[853],row_in_1[853],row_in_2[853]};
assign col_in_854 = {row_in_0[854],row_in_1[854],row_in_2[854]};
assign col_in_855 = {row_in_0[855],row_in_1[855],row_in_2[855]};
assign col_in_856 = {row_in_0[856],row_in_1[856],row_in_2[856]};
assign col_in_857 = {row_in_0[857],row_in_1[857],row_in_2[857]};
assign col_in_858 = {row_in_0[858],row_in_1[858],row_in_2[858]};
assign col_in_859 = {row_in_0[859],row_in_1[859],row_in_2[859]};
assign col_in_860 = {row_in_0[860],row_in_1[860],row_in_2[860]};
assign col_in_861 = {row_in_0[861],row_in_1[861],row_in_2[861]};
assign col_in_862 = {row_in_0[862],row_in_1[862],row_in_2[862]};
assign col_in_863 = {row_in_0[863],row_in_1[863],row_in_2[863]};
assign col_in_864 = {row_in_0[864],row_in_1[864],row_in_2[864]};
assign col_in_865 = {row_in_0[865],row_in_1[865],row_in_2[865]};
assign col_in_866 = {row_in_0[866],row_in_1[866],row_in_2[866]};
assign col_in_867 = {row_in_0[867],row_in_1[867],row_in_2[867]};
assign col_in_868 = {row_in_0[868],row_in_1[868],row_in_2[868]};
assign col_in_869 = {row_in_0[869],row_in_1[869],row_in_2[869]};
assign col_in_870 = {row_in_0[870],row_in_1[870],row_in_2[870]};
assign col_in_871 = {row_in_0[871],row_in_1[871],row_in_2[871]};
assign col_in_872 = {row_in_0[872],row_in_1[872],row_in_2[872]};
assign col_in_873 = {row_in_0[873],row_in_1[873],row_in_2[873]};
assign col_in_874 = {row_in_0[874],row_in_1[874],row_in_2[874]};
assign col_in_875 = {row_in_0[875],row_in_1[875],row_in_2[875]};
assign col_in_876 = {row_in_0[876],row_in_1[876],row_in_2[876]};
assign col_in_877 = {row_in_0[877],row_in_1[877],row_in_2[877]};
assign col_in_878 = {row_in_0[878],row_in_1[878],row_in_2[878]};
assign col_in_879 = {row_in_0[879],row_in_1[879],row_in_2[879]};
assign col_in_880 = {row_in_0[880],row_in_1[880],row_in_2[880]};
assign col_in_881 = {row_in_0[881],row_in_1[881],row_in_2[881]};
assign col_in_882 = {row_in_0[882],row_in_1[882],row_in_2[882]};
assign col_in_883 = {row_in_0[883],row_in_1[883],row_in_2[883]};
assign col_in_884 = {row_in_0[884],row_in_1[884],row_in_2[884]};
assign col_in_885 = {row_in_0[885],row_in_1[885],row_in_2[885]};
assign col_in_886 = {row_in_0[886],row_in_1[886],row_in_2[886]};
assign col_in_887 = {row_in_0[887],row_in_1[887],row_in_2[887]};
assign col_in_888 = {row_in_0[888],row_in_1[888],row_in_2[888]};
assign col_in_889 = {row_in_0[889],row_in_1[889],row_in_2[889]};
assign col_in_890 = {row_in_0[890],row_in_1[890],row_in_2[890]};
assign col_in_891 = {row_in_0[891],row_in_1[891],row_in_2[891]};
assign col_in_892 = {row_in_0[892],row_in_1[892],row_in_2[892]};
assign col_in_893 = {row_in_0[893],row_in_1[893],row_in_2[893]};
assign col_in_894 = {row_in_0[894],row_in_1[894],row_in_2[894]};
assign col_in_895 = {row_in_0[895],row_in_1[895],row_in_2[895]};
assign col_in_896 = {row_in_0[896],row_in_1[896],row_in_2[896]};
assign col_in_897 = {row_in_0[897],row_in_1[897],row_in_2[897]};
assign col_in_898 = {row_in_0[898],row_in_1[898],row_in_2[898]};
assign col_in_899 = {row_in_0[899],row_in_1[899],row_in_2[899]};
assign col_in_900 = {row_in_0[900],row_in_1[900],row_in_2[900]};
assign col_in_901 = {row_in_0[901],row_in_1[901],row_in_2[901]};
assign col_in_902 = {row_in_0[902],row_in_1[902],row_in_2[902]};
assign col_in_903 = {row_in_0[903],row_in_1[903],row_in_2[903]};
assign col_in_904 = {row_in_0[904],row_in_1[904],row_in_2[904]};
assign col_in_905 = {row_in_0[905],row_in_1[905],row_in_2[905]};
assign col_in_906 = {row_in_0[906],row_in_1[906],row_in_2[906]};
assign col_in_907 = {row_in_0[907],row_in_1[907],row_in_2[907]};
assign col_in_908 = {row_in_0[908],row_in_1[908],row_in_2[908]};
assign col_in_909 = {row_in_0[909],row_in_1[909],row_in_2[909]};
assign col_in_910 = {row_in_0[910],row_in_1[910],row_in_2[910]};
assign col_in_911 = {row_in_0[911],row_in_1[911],row_in_2[911]};
assign col_in_912 = {row_in_0[912],row_in_1[912],row_in_2[912]};
assign col_in_913 = {row_in_0[913],row_in_1[913],row_in_2[913]};
assign col_in_914 = {row_in_0[914],row_in_1[914],row_in_2[914]};
assign col_in_915 = {row_in_0[915],row_in_1[915],row_in_2[915]};
assign col_in_916 = {row_in_0[916],row_in_1[916],row_in_2[916]};
assign col_in_917 = {row_in_0[917],row_in_1[917],row_in_2[917]};
assign col_in_918 = {row_in_0[918],row_in_1[918],row_in_2[918]};
assign col_in_919 = {row_in_0[919],row_in_1[919],row_in_2[919]};
assign col_in_920 = {row_in_0[920],row_in_1[920],row_in_2[920]};
assign col_in_921 = {row_in_0[921],row_in_1[921],row_in_2[921]};
assign col_in_922 = {row_in_0[922],row_in_1[922],row_in_2[922]};
assign col_in_923 = {row_in_0[923],row_in_1[923],row_in_2[923]};
assign col_in_924 = {row_in_0[924],row_in_1[924],row_in_2[924]};
assign col_in_925 = {row_in_0[925],row_in_1[925],row_in_2[925]};
assign col_in_926 = {row_in_0[926],row_in_1[926],row_in_2[926]};
assign col_in_927 = {row_in_0[927],row_in_1[927],row_in_2[927]};
assign col_in_928 = {row_in_0[928],row_in_1[928],row_in_2[928]};
assign col_in_929 = {row_in_0[929],row_in_1[929],row_in_2[929]};
assign col_in_930 = {row_in_0[930],row_in_1[930],row_in_2[930]};
assign col_in_931 = {row_in_0[931],row_in_1[931],row_in_2[931]};
assign col_in_932 = {row_in_0[932],row_in_1[932],row_in_2[932]};
assign col_in_933 = {row_in_0[933],row_in_1[933],row_in_2[933]};
assign col_in_934 = {row_in_0[934],row_in_1[934],row_in_2[934]};
assign col_in_935 = {row_in_0[935],row_in_1[935],row_in_2[935]};
assign col_in_936 = {row_in_0[936],row_in_1[936],row_in_2[936]};
assign col_in_937 = {row_in_0[937],row_in_1[937],row_in_2[937]};
assign col_in_938 = {row_in_0[938],row_in_1[938],row_in_2[938]};
assign col_in_939 = {row_in_0[939],row_in_1[939],row_in_2[939]};
assign col_in_940 = {row_in_0[940],row_in_1[940],row_in_2[940]};
assign col_in_941 = {row_in_0[941],row_in_1[941],row_in_2[941]};
assign col_in_942 = {row_in_0[942],row_in_1[942],row_in_2[942]};
assign col_in_943 = {row_in_0[943],row_in_1[943],row_in_2[943]};
assign col_in_944 = {row_in_0[944],row_in_1[944],row_in_2[944]};
assign col_in_945 = {row_in_0[945],row_in_1[945],row_in_2[945]};
assign col_in_946 = {row_in_0[946],row_in_1[946],row_in_2[946]};
assign col_in_947 = {row_in_0[947],row_in_1[947],row_in_2[947]};
assign col_in_948 = {row_in_0[948],row_in_1[948],row_in_2[948]};
assign col_in_949 = {row_in_0[949],row_in_1[949],row_in_2[949]};
assign col_in_950 = {row_in_0[950],row_in_1[950],row_in_2[950]};
assign col_in_951 = {row_in_0[951],row_in_1[951],row_in_2[951]};
assign col_in_952 = {row_in_0[952],row_in_1[952],row_in_2[952]};
assign col_in_953 = {row_in_0[953],row_in_1[953],row_in_2[953]};
assign col_in_954 = {row_in_0[954],row_in_1[954],row_in_2[954]};
assign col_in_955 = {row_in_0[955],row_in_1[955],row_in_2[955]};
assign col_in_956 = {row_in_0[956],row_in_1[956],row_in_2[956]};
assign col_in_957 = {row_in_0[957],row_in_1[957],row_in_2[957]};
assign col_in_958 = {row_in_0[958],row_in_1[958],row_in_2[958]};
assign col_in_959 = {row_in_0[959],row_in_1[959],row_in_2[959]};
assign col_in_960 = {row_in_0[960],row_in_1[960],row_in_2[960]};
assign col_in_961 = {row_in_0[961],row_in_1[961],row_in_2[961]};
assign col_in_962 = {row_in_0[962],row_in_1[962],row_in_2[962]};
assign col_in_963 = {row_in_0[963],row_in_1[963],row_in_2[963]};
assign col_in_964 = {row_in_0[964],row_in_1[964],row_in_2[964]};
assign col_in_965 = {row_in_0[965],row_in_1[965],row_in_2[965]};
assign col_in_966 = {row_in_0[966],row_in_1[966],row_in_2[966]};
assign col_in_967 = {row_in_0[967],row_in_1[967],row_in_2[967]};
assign col_in_968 = {row_in_0[968],row_in_1[968],row_in_2[968]};
assign col_in_969 = {row_in_0[969],row_in_1[969],row_in_2[969]};
assign col_in_970 = {row_in_0[970],row_in_1[970],row_in_2[970]};
assign col_in_971 = {row_in_0[971],row_in_1[971],row_in_2[971]};
assign col_in_972 = {row_in_0[972],row_in_1[972],row_in_2[972]};
assign col_in_973 = {row_in_0[973],row_in_1[973],row_in_2[973]};
assign col_in_974 = {row_in_0[974],row_in_1[974],row_in_2[974]};
assign col_in_975 = {row_in_0[975],row_in_1[975],row_in_2[975]};
assign col_in_976 = {row_in_0[976],row_in_1[976],row_in_2[976]};
assign col_in_977 = {row_in_0[977],row_in_1[977],row_in_2[977]};
assign col_in_978 = {row_in_0[978],row_in_1[978],row_in_2[978]};
assign col_in_979 = {row_in_0[979],row_in_1[979],row_in_2[979]};
assign col_in_980 = {row_in_0[980],row_in_1[980],row_in_2[980]};
assign col_in_981 = {row_in_0[981],row_in_1[981],row_in_2[981]};
assign col_in_982 = {row_in_0[982],row_in_1[982],row_in_2[982]};
assign col_in_983 = {row_in_0[983],row_in_1[983],row_in_2[983]};
assign col_in_984 = {row_in_0[984],row_in_1[984],row_in_2[984]};
assign col_in_985 = {row_in_0[985],row_in_1[985],row_in_2[985]};
assign col_in_986 = {row_in_0[986],row_in_1[986],row_in_2[986]};
assign col_in_987 = {row_in_0[987],row_in_1[987],row_in_2[987]};
assign col_in_988 = {row_in_0[988],row_in_1[988],row_in_2[988]};
assign col_in_989 = {row_in_0[989],row_in_1[989],row_in_2[989]};
assign col_in_990 = {row_in_0[990],row_in_1[990],row_in_2[990]};
assign col_in_991 = {row_in_0[991],row_in_1[991],row_in_2[991]};
assign col_in_992 = {row_in_0[992],row_in_1[992],row_in_2[992]};
assign col_in_993 = {row_in_0[993],row_in_1[993],row_in_2[993]};
assign col_in_994 = {row_in_0[994],row_in_1[994],row_in_2[994]};
assign col_in_995 = {row_in_0[995],row_in_1[995],row_in_2[995]};
assign col_in_996 = {row_in_0[996],row_in_1[996],row_in_2[996]};
assign col_in_997 = {row_in_0[997],row_in_1[997],row_in_2[997]};
assign col_in_998 = {row_in_0[998],row_in_1[998],row_in_2[998]};
assign col_in_999 = {row_in_0[999],row_in_1[999],row_in_2[999]};
assign col_in_1000 = {row_in_0[1000],row_in_1[1000],row_in_2[1000]};
assign col_in_1001 = {row_in_0[1001],row_in_1[1001],row_in_2[1001]};
assign col_in_1002 = {row_in_0[1002],row_in_1[1002],row_in_2[1002]};
assign col_in_1003 = {row_in_0[1003],row_in_1[1003],row_in_2[1003]};
assign col_in_1004 = {row_in_0[1004],row_in_1[1004],row_in_2[1004]};
assign col_in_1005 = {row_in_0[1005],row_in_1[1005],row_in_2[1005]};
assign col_in_1006 = {row_in_0[1006],row_in_1[1006],row_in_2[1006]};
assign col_in_1007 = {row_in_0[1007],row_in_1[1007],row_in_2[1007]};
assign col_in_1008 = {row_in_0[1008],row_in_1[1008],row_in_2[1008]};
assign col_in_1009 = {row_in_0[1009],row_in_1[1009],row_in_2[1009]};
assign col_in_1010 = {row_in_0[1010],row_in_1[1010],row_in_2[1010]};
assign col_in_1011 = {row_in_0[1011],row_in_1[1011],row_in_2[1011]};
assign col_in_1012 = {row_in_0[1012],row_in_1[1012],row_in_2[1012]};
assign col_in_1013 = {row_in_0[1013],row_in_1[1013],row_in_2[1013]};
assign col_in_1014 = {row_in_0[1014],row_in_1[1014],row_in_2[1014]};
assign col_in_1015 = {row_in_0[1015],row_in_1[1015],row_in_2[1015]};
assign col_in_1016 = {row_in_0[1016],row_in_1[1016],row_in_2[1016]};
assign col_in_1017 = {row_in_0[1017],row_in_1[1017],row_in_2[1017]};
assign col_in_1018 = {row_in_0[1018],row_in_1[1018],row_in_2[1018]};
assign col_in_1019 = {row_in_0[1019],row_in_1[1019],row_in_2[1019]};
assign col_in_1020 = {row_in_0[1020],row_in_1[1020],row_in_2[1020]};
assign col_in_1021 = {row_in_0[1021],row_in_1[1021],row_in_2[1021]};
assign col_in_1022 = {row_in_0[1022],row_in_1[1022],row_in_2[1022]};
assign col_in_1023 = {row_in_0[1023],row_in_1[1023],row_in_2[1023]};
















// compressor_array_3_2_1024 Outputs
wire  [1:0]  col_out_0;
wire  [1:0]  col_out_1;
wire  [1:0]  col_out_2;
wire  [1:0]  col_out_3;
wire  [1:0]  col_out_4;
wire  [1:0]  col_out_5;
wire  [1:0]  col_out_6;
wire  [1:0]  col_out_7;
wire  [1:0]  col_out_8;
wire  [1:0]  col_out_9;
wire  [1:0]  col_out_10;
wire  [1:0]  col_out_11;
wire  [1:0]  col_out_12;
wire  [1:0]  col_out_13;
wire  [1:0]  col_out_14;
wire  [1:0]  col_out_15;
wire  [1:0]  col_out_16;
wire  [1:0]  col_out_17;
wire  [1:0]  col_out_18;
wire  [1:0]  col_out_19;
wire  [1:0]  col_out_20;
wire  [1:0]  col_out_21;
wire  [1:0]  col_out_22;
wire  [1:0]  col_out_23;
wire  [1:0]  col_out_24;
wire  [1:0]  col_out_25;
wire  [1:0]  col_out_26;
wire  [1:0]  col_out_27;
wire  [1:0]  col_out_28;
wire  [1:0]  col_out_29;
wire  [1:0]  col_out_30;
wire  [1:0]  col_out_31;
wire  [1:0]  col_out_32;
wire  [1:0]  col_out_33;
wire  [1:0]  col_out_34;
wire  [1:0]  col_out_35;
wire  [1:0]  col_out_36;
wire  [1:0]  col_out_37;
wire  [1:0]  col_out_38;
wire  [1:0]  col_out_39;
wire  [1:0]  col_out_40;
wire  [1:0]  col_out_41;
wire  [1:0]  col_out_42;
wire  [1:0]  col_out_43;
wire  [1:0]  col_out_44;
wire  [1:0]  col_out_45;
wire  [1:0]  col_out_46;
wire  [1:0]  col_out_47;
wire  [1:0]  col_out_48;
wire  [1:0]  col_out_49;
wire  [1:0]  col_out_50;
wire  [1:0]  col_out_51;
wire  [1:0]  col_out_52;
wire  [1:0]  col_out_53;
wire  [1:0]  col_out_54;
wire  [1:0]  col_out_55;
wire  [1:0]  col_out_56;
wire  [1:0]  col_out_57;
wire  [1:0]  col_out_58;
wire  [1:0]  col_out_59;
wire  [1:0]  col_out_60;
wire  [1:0]  col_out_61;
wire  [1:0]  col_out_62;
wire  [1:0]  col_out_63;
wire  [1:0]  col_out_64;
wire  [1:0]  col_out_65;
wire  [1:0]  col_out_66;
wire  [1:0]  col_out_67;
wire  [1:0]  col_out_68;
wire  [1:0]  col_out_69;
wire  [1:0]  col_out_70;
wire  [1:0]  col_out_71;
wire  [1:0]  col_out_72;
wire  [1:0]  col_out_73;
wire  [1:0]  col_out_74;
wire  [1:0]  col_out_75;
wire  [1:0]  col_out_76;
wire  [1:0]  col_out_77;
wire  [1:0]  col_out_78;
wire  [1:0]  col_out_79;
wire  [1:0]  col_out_80;
wire  [1:0]  col_out_81;
wire  [1:0]  col_out_82;
wire  [1:0]  col_out_83;
wire  [1:0]  col_out_84;
wire  [1:0]  col_out_85;
wire  [1:0]  col_out_86;
wire  [1:0]  col_out_87;
wire  [1:0]  col_out_88;
wire  [1:0]  col_out_89;
wire  [1:0]  col_out_90;
wire  [1:0]  col_out_91;
wire  [1:0]  col_out_92;
wire  [1:0]  col_out_93;
wire  [1:0]  col_out_94;
wire  [1:0]  col_out_95;
wire  [1:0]  col_out_96;
wire  [1:0]  col_out_97;
wire  [1:0]  col_out_98;
wire  [1:0]  col_out_99;
wire  [1:0]  col_out_100;
wire  [1:0]  col_out_101;
wire  [1:0]  col_out_102;
wire  [1:0]  col_out_103;
wire  [1:0]  col_out_104;
wire  [1:0]  col_out_105;
wire  [1:0]  col_out_106;
wire  [1:0]  col_out_107;
wire  [1:0]  col_out_108;
wire  [1:0]  col_out_109;
wire  [1:0]  col_out_110;
wire  [1:0]  col_out_111;
wire  [1:0]  col_out_112;
wire  [1:0]  col_out_113;
wire  [1:0]  col_out_114;
wire  [1:0]  col_out_115;
wire  [1:0]  col_out_116;
wire  [1:0]  col_out_117;
wire  [1:0]  col_out_118;
wire  [1:0]  col_out_119;
wire  [1:0]  col_out_120;
wire  [1:0]  col_out_121;
wire  [1:0]  col_out_122;
wire  [1:0]  col_out_123;
wire  [1:0]  col_out_124;
wire  [1:0]  col_out_125;
wire  [1:0]  col_out_126;
wire  [1:0]  col_out_127;
wire  [1:0]  col_out_128;
wire  [1:0]  col_out_129;
wire  [1:0]  col_out_130;
wire  [1:0]  col_out_131;
wire  [1:0]  col_out_132;
wire  [1:0]  col_out_133;
wire  [1:0]  col_out_134;
wire  [1:0]  col_out_135;
wire  [1:0]  col_out_136;
wire  [1:0]  col_out_137;
wire  [1:0]  col_out_138;
wire  [1:0]  col_out_139;
wire  [1:0]  col_out_140;
wire  [1:0]  col_out_141;
wire  [1:0]  col_out_142;
wire  [1:0]  col_out_143;
wire  [1:0]  col_out_144;
wire  [1:0]  col_out_145;
wire  [1:0]  col_out_146;
wire  [1:0]  col_out_147;
wire  [1:0]  col_out_148;
wire  [1:0]  col_out_149;
wire  [1:0]  col_out_150;
wire  [1:0]  col_out_151;
wire  [1:0]  col_out_152;
wire  [1:0]  col_out_153;
wire  [1:0]  col_out_154;
wire  [1:0]  col_out_155;
wire  [1:0]  col_out_156;
wire  [1:0]  col_out_157;
wire  [1:0]  col_out_158;
wire  [1:0]  col_out_159;
wire  [1:0]  col_out_160;
wire  [1:0]  col_out_161;
wire  [1:0]  col_out_162;
wire  [1:0]  col_out_163;
wire  [1:0]  col_out_164;
wire  [1:0]  col_out_165;
wire  [1:0]  col_out_166;
wire  [1:0]  col_out_167;
wire  [1:0]  col_out_168;
wire  [1:0]  col_out_169;
wire  [1:0]  col_out_170;
wire  [1:0]  col_out_171;
wire  [1:0]  col_out_172;
wire  [1:0]  col_out_173;
wire  [1:0]  col_out_174;
wire  [1:0]  col_out_175;
wire  [1:0]  col_out_176;
wire  [1:0]  col_out_177;
wire  [1:0]  col_out_178;
wire  [1:0]  col_out_179;
wire  [1:0]  col_out_180;
wire  [1:0]  col_out_181;
wire  [1:0]  col_out_182;
wire  [1:0]  col_out_183;
wire  [1:0]  col_out_184;
wire  [1:0]  col_out_185;
wire  [1:0]  col_out_186;
wire  [1:0]  col_out_187;
wire  [1:0]  col_out_188;
wire  [1:0]  col_out_189;
wire  [1:0]  col_out_190;
wire  [1:0]  col_out_191;
wire  [1:0]  col_out_192;
wire  [1:0]  col_out_193;
wire  [1:0]  col_out_194;
wire  [1:0]  col_out_195;
wire  [1:0]  col_out_196;
wire  [1:0]  col_out_197;
wire  [1:0]  col_out_198;
wire  [1:0]  col_out_199;
wire  [1:0]  col_out_200;
wire  [1:0]  col_out_201;
wire  [1:0]  col_out_202;
wire  [1:0]  col_out_203;
wire  [1:0]  col_out_204;
wire  [1:0]  col_out_205;
wire  [1:0]  col_out_206;
wire  [1:0]  col_out_207;
wire  [1:0]  col_out_208;
wire  [1:0]  col_out_209;
wire  [1:0]  col_out_210;
wire  [1:0]  col_out_211;
wire  [1:0]  col_out_212;
wire  [1:0]  col_out_213;
wire  [1:0]  col_out_214;
wire  [1:0]  col_out_215;
wire  [1:0]  col_out_216;
wire  [1:0]  col_out_217;
wire  [1:0]  col_out_218;
wire  [1:0]  col_out_219;
wire  [1:0]  col_out_220;
wire  [1:0]  col_out_221;
wire  [1:0]  col_out_222;
wire  [1:0]  col_out_223;
wire  [1:0]  col_out_224;
wire  [1:0]  col_out_225;
wire  [1:0]  col_out_226;
wire  [1:0]  col_out_227;
wire  [1:0]  col_out_228;
wire  [1:0]  col_out_229;
wire  [1:0]  col_out_230;
wire  [1:0]  col_out_231;
wire  [1:0]  col_out_232;
wire  [1:0]  col_out_233;
wire  [1:0]  col_out_234;
wire  [1:0]  col_out_235;
wire  [1:0]  col_out_236;
wire  [1:0]  col_out_237;
wire  [1:0]  col_out_238;
wire  [1:0]  col_out_239;
wire  [1:0]  col_out_240;
wire  [1:0]  col_out_241;
wire  [1:0]  col_out_242;
wire  [1:0]  col_out_243;
wire  [1:0]  col_out_244;
wire  [1:0]  col_out_245;
wire  [1:0]  col_out_246;
wire  [1:0]  col_out_247;
wire  [1:0]  col_out_248;
wire  [1:0]  col_out_249;
wire  [1:0]  col_out_250;
wire  [1:0]  col_out_251;
wire  [1:0]  col_out_252;
wire  [1:0]  col_out_253;
wire  [1:0]  col_out_254;
wire  [1:0]  col_out_255;
wire  [1:0]  col_out_256;
wire  [1:0]  col_out_257;
wire  [1:0]  col_out_258;
wire  [1:0]  col_out_259;
wire  [1:0]  col_out_260;
wire  [1:0]  col_out_261;
wire  [1:0]  col_out_262;
wire  [1:0]  col_out_263;
wire  [1:0]  col_out_264;
wire  [1:0]  col_out_265;
wire  [1:0]  col_out_266;
wire  [1:0]  col_out_267;
wire  [1:0]  col_out_268;
wire  [1:0]  col_out_269;
wire  [1:0]  col_out_270;
wire  [1:0]  col_out_271;
wire  [1:0]  col_out_272;
wire  [1:0]  col_out_273;
wire  [1:0]  col_out_274;
wire  [1:0]  col_out_275;
wire  [1:0]  col_out_276;
wire  [1:0]  col_out_277;
wire  [1:0]  col_out_278;
wire  [1:0]  col_out_279;
wire  [1:0]  col_out_280;
wire  [1:0]  col_out_281;
wire  [1:0]  col_out_282;
wire  [1:0]  col_out_283;
wire  [1:0]  col_out_284;
wire  [1:0]  col_out_285;
wire  [1:0]  col_out_286;
wire  [1:0]  col_out_287;
wire  [1:0]  col_out_288;
wire  [1:0]  col_out_289;
wire  [1:0]  col_out_290;
wire  [1:0]  col_out_291;
wire  [1:0]  col_out_292;
wire  [1:0]  col_out_293;
wire  [1:0]  col_out_294;
wire  [1:0]  col_out_295;
wire  [1:0]  col_out_296;
wire  [1:0]  col_out_297;
wire  [1:0]  col_out_298;
wire  [1:0]  col_out_299;
wire  [1:0]  col_out_300;
wire  [1:0]  col_out_301;
wire  [1:0]  col_out_302;
wire  [1:0]  col_out_303;
wire  [1:0]  col_out_304;
wire  [1:0]  col_out_305;
wire  [1:0]  col_out_306;
wire  [1:0]  col_out_307;
wire  [1:0]  col_out_308;
wire  [1:0]  col_out_309;
wire  [1:0]  col_out_310;
wire  [1:0]  col_out_311;
wire  [1:0]  col_out_312;
wire  [1:0]  col_out_313;
wire  [1:0]  col_out_314;
wire  [1:0]  col_out_315;
wire  [1:0]  col_out_316;
wire  [1:0]  col_out_317;
wire  [1:0]  col_out_318;
wire  [1:0]  col_out_319;
wire  [1:0]  col_out_320;
wire  [1:0]  col_out_321;
wire  [1:0]  col_out_322;
wire  [1:0]  col_out_323;
wire  [1:0]  col_out_324;
wire  [1:0]  col_out_325;
wire  [1:0]  col_out_326;
wire  [1:0]  col_out_327;
wire  [1:0]  col_out_328;
wire  [1:0]  col_out_329;
wire  [1:0]  col_out_330;
wire  [1:0]  col_out_331;
wire  [1:0]  col_out_332;
wire  [1:0]  col_out_333;
wire  [1:0]  col_out_334;
wire  [1:0]  col_out_335;
wire  [1:0]  col_out_336;
wire  [1:0]  col_out_337;
wire  [1:0]  col_out_338;
wire  [1:0]  col_out_339;
wire  [1:0]  col_out_340;
wire  [1:0]  col_out_341;
wire  [1:0]  col_out_342;
wire  [1:0]  col_out_343;
wire  [1:0]  col_out_344;
wire  [1:0]  col_out_345;
wire  [1:0]  col_out_346;
wire  [1:0]  col_out_347;
wire  [1:0]  col_out_348;
wire  [1:0]  col_out_349;
wire  [1:0]  col_out_350;
wire  [1:0]  col_out_351;
wire  [1:0]  col_out_352;
wire  [1:0]  col_out_353;
wire  [1:0]  col_out_354;
wire  [1:0]  col_out_355;
wire  [1:0]  col_out_356;
wire  [1:0]  col_out_357;
wire  [1:0]  col_out_358;
wire  [1:0]  col_out_359;
wire  [1:0]  col_out_360;
wire  [1:0]  col_out_361;
wire  [1:0]  col_out_362;
wire  [1:0]  col_out_363;
wire  [1:0]  col_out_364;
wire  [1:0]  col_out_365;
wire  [1:0]  col_out_366;
wire  [1:0]  col_out_367;
wire  [1:0]  col_out_368;
wire  [1:0]  col_out_369;
wire  [1:0]  col_out_370;
wire  [1:0]  col_out_371;
wire  [1:0]  col_out_372;
wire  [1:0]  col_out_373;
wire  [1:0]  col_out_374;
wire  [1:0]  col_out_375;
wire  [1:0]  col_out_376;
wire  [1:0]  col_out_377;
wire  [1:0]  col_out_378;
wire  [1:0]  col_out_379;
wire  [1:0]  col_out_380;
wire  [1:0]  col_out_381;
wire  [1:0]  col_out_382;
wire  [1:0]  col_out_383;
wire  [1:0]  col_out_384;
wire  [1:0]  col_out_385;
wire  [1:0]  col_out_386;
wire  [1:0]  col_out_387;
wire  [1:0]  col_out_388;
wire  [1:0]  col_out_389;
wire  [1:0]  col_out_390;
wire  [1:0]  col_out_391;
wire  [1:0]  col_out_392;
wire  [1:0]  col_out_393;
wire  [1:0]  col_out_394;
wire  [1:0]  col_out_395;
wire  [1:0]  col_out_396;
wire  [1:0]  col_out_397;
wire  [1:0]  col_out_398;
wire  [1:0]  col_out_399;
wire  [1:0]  col_out_400;
wire  [1:0]  col_out_401;
wire  [1:0]  col_out_402;
wire  [1:0]  col_out_403;
wire  [1:0]  col_out_404;
wire  [1:0]  col_out_405;
wire  [1:0]  col_out_406;
wire  [1:0]  col_out_407;
wire  [1:0]  col_out_408;
wire  [1:0]  col_out_409;
wire  [1:0]  col_out_410;
wire  [1:0]  col_out_411;
wire  [1:0]  col_out_412;
wire  [1:0]  col_out_413;
wire  [1:0]  col_out_414;
wire  [1:0]  col_out_415;
wire  [1:0]  col_out_416;
wire  [1:0]  col_out_417;
wire  [1:0]  col_out_418;
wire  [1:0]  col_out_419;
wire  [1:0]  col_out_420;
wire  [1:0]  col_out_421;
wire  [1:0]  col_out_422;
wire  [1:0]  col_out_423;
wire  [1:0]  col_out_424;
wire  [1:0]  col_out_425;
wire  [1:0]  col_out_426;
wire  [1:0]  col_out_427;
wire  [1:0]  col_out_428;
wire  [1:0]  col_out_429;
wire  [1:0]  col_out_430;
wire  [1:0]  col_out_431;
wire  [1:0]  col_out_432;
wire  [1:0]  col_out_433;
wire  [1:0]  col_out_434;
wire  [1:0]  col_out_435;
wire  [1:0]  col_out_436;
wire  [1:0]  col_out_437;
wire  [1:0]  col_out_438;
wire  [1:0]  col_out_439;
wire  [1:0]  col_out_440;
wire  [1:0]  col_out_441;
wire  [1:0]  col_out_442;
wire  [1:0]  col_out_443;
wire  [1:0]  col_out_444;
wire  [1:0]  col_out_445;
wire  [1:0]  col_out_446;
wire  [1:0]  col_out_447;
wire  [1:0]  col_out_448;
wire  [1:0]  col_out_449;
wire  [1:0]  col_out_450;
wire  [1:0]  col_out_451;
wire  [1:0]  col_out_452;
wire  [1:0]  col_out_453;
wire  [1:0]  col_out_454;
wire  [1:0]  col_out_455;
wire  [1:0]  col_out_456;
wire  [1:0]  col_out_457;
wire  [1:0]  col_out_458;
wire  [1:0]  col_out_459;
wire  [1:0]  col_out_460;
wire  [1:0]  col_out_461;
wire  [1:0]  col_out_462;
wire  [1:0]  col_out_463;
wire  [1:0]  col_out_464;
wire  [1:0]  col_out_465;
wire  [1:0]  col_out_466;
wire  [1:0]  col_out_467;
wire  [1:0]  col_out_468;
wire  [1:0]  col_out_469;
wire  [1:0]  col_out_470;
wire  [1:0]  col_out_471;
wire  [1:0]  col_out_472;
wire  [1:0]  col_out_473;
wire  [1:0]  col_out_474;
wire  [1:0]  col_out_475;
wire  [1:0]  col_out_476;
wire  [1:0]  col_out_477;
wire  [1:0]  col_out_478;
wire  [1:0]  col_out_479;
wire  [1:0]  col_out_480;
wire  [1:0]  col_out_481;
wire  [1:0]  col_out_482;
wire  [1:0]  col_out_483;
wire  [1:0]  col_out_484;
wire  [1:0]  col_out_485;
wire  [1:0]  col_out_486;
wire  [1:0]  col_out_487;
wire  [1:0]  col_out_488;
wire  [1:0]  col_out_489;
wire  [1:0]  col_out_490;
wire  [1:0]  col_out_491;
wire  [1:0]  col_out_492;
wire  [1:0]  col_out_493;
wire  [1:0]  col_out_494;
wire  [1:0]  col_out_495;
wire  [1:0]  col_out_496;
wire  [1:0]  col_out_497;
wire  [1:0]  col_out_498;
wire  [1:0]  col_out_499;
wire  [1:0]  col_out_500;
wire  [1:0]  col_out_501;
wire  [1:0]  col_out_502;
wire  [1:0]  col_out_503;
wire  [1:0]  col_out_504;
wire  [1:0]  col_out_505;
wire  [1:0]  col_out_506;
wire  [1:0]  col_out_507;
wire  [1:0]  col_out_508;
wire  [1:0]  col_out_509;
wire  [1:0]  col_out_510;
wire  [1:0]  col_out_511;
wire  [1:0]  col_out_512;
wire  [1:0]  col_out_513;
wire  [1:0]  col_out_514;
wire  [1:0]  col_out_515;
wire  [1:0]  col_out_516;
wire  [1:0]  col_out_517;
wire  [1:0]  col_out_518;
wire  [1:0]  col_out_519;
wire  [1:0]  col_out_520;
wire  [1:0]  col_out_521;
wire  [1:0]  col_out_522;
wire  [1:0]  col_out_523;
wire  [1:0]  col_out_524;
wire  [1:0]  col_out_525;
wire  [1:0]  col_out_526;
wire  [1:0]  col_out_527;
wire  [1:0]  col_out_528;
wire  [1:0]  col_out_529;
wire  [1:0]  col_out_530;
wire  [1:0]  col_out_531;
wire  [1:0]  col_out_532;
wire  [1:0]  col_out_533;
wire  [1:0]  col_out_534;
wire  [1:0]  col_out_535;
wire  [1:0]  col_out_536;
wire  [1:0]  col_out_537;
wire  [1:0]  col_out_538;
wire  [1:0]  col_out_539;
wire  [1:0]  col_out_540;
wire  [1:0]  col_out_541;
wire  [1:0]  col_out_542;
wire  [1:0]  col_out_543;
wire  [1:0]  col_out_544;
wire  [1:0]  col_out_545;
wire  [1:0]  col_out_546;
wire  [1:0]  col_out_547;
wire  [1:0]  col_out_548;
wire  [1:0]  col_out_549;
wire  [1:0]  col_out_550;
wire  [1:0]  col_out_551;
wire  [1:0]  col_out_552;
wire  [1:0]  col_out_553;
wire  [1:0]  col_out_554;
wire  [1:0]  col_out_555;
wire  [1:0]  col_out_556;
wire  [1:0]  col_out_557;
wire  [1:0]  col_out_558;
wire  [1:0]  col_out_559;
wire  [1:0]  col_out_560;
wire  [1:0]  col_out_561;
wire  [1:0]  col_out_562;
wire  [1:0]  col_out_563;
wire  [1:0]  col_out_564;
wire  [1:0]  col_out_565;
wire  [1:0]  col_out_566;
wire  [1:0]  col_out_567;
wire  [1:0]  col_out_568;
wire  [1:0]  col_out_569;
wire  [1:0]  col_out_570;
wire  [1:0]  col_out_571;
wire  [1:0]  col_out_572;
wire  [1:0]  col_out_573;
wire  [1:0]  col_out_574;
wire  [1:0]  col_out_575;
wire  [1:0]  col_out_576;
wire  [1:0]  col_out_577;
wire  [1:0]  col_out_578;
wire  [1:0]  col_out_579;
wire  [1:0]  col_out_580;
wire  [1:0]  col_out_581;
wire  [1:0]  col_out_582;
wire  [1:0]  col_out_583;
wire  [1:0]  col_out_584;
wire  [1:0]  col_out_585;
wire  [1:0]  col_out_586;
wire  [1:0]  col_out_587;
wire  [1:0]  col_out_588;
wire  [1:0]  col_out_589;
wire  [1:0]  col_out_590;
wire  [1:0]  col_out_591;
wire  [1:0]  col_out_592;
wire  [1:0]  col_out_593;
wire  [1:0]  col_out_594;
wire  [1:0]  col_out_595;
wire  [1:0]  col_out_596;
wire  [1:0]  col_out_597;
wire  [1:0]  col_out_598;
wire  [1:0]  col_out_599;
wire  [1:0]  col_out_600;
wire  [1:0]  col_out_601;
wire  [1:0]  col_out_602;
wire  [1:0]  col_out_603;
wire  [1:0]  col_out_604;
wire  [1:0]  col_out_605;
wire  [1:0]  col_out_606;
wire  [1:0]  col_out_607;
wire  [1:0]  col_out_608;
wire  [1:0]  col_out_609;
wire  [1:0]  col_out_610;
wire  [1:0]  col_out_611;
wire  [1:0]  col_out_612;
wire  [1:0]  col_out_613;
wire  [1:0]  col_out_614;
wire  [1:0]  col_out_615;
wire  [1:0]  col_out_616;
wire  [1:0]  col_out_617;
wire  [1:0]  col_out_618;
wire  [1:0]  col_out_619;
wire  [1:0]  col_out_620;
wire  [1:0]  col_out_621;
wire  [1:0]  col_out_622;
wire  [1:0]  col_out_623;
wire  [1:0]  col_out_624;
wire  [1:0]  col_out_625;
wire  [1:0]  col_out_626;
wire  [1:0]  col_out_627;
wire  [1:0]  col_out_628;
wire  [1:0]  col_out_629;
wire  [1:0]  col_out_630;
wire  [1:0]  col_out_631;
wire  [1:0]  col_out_632;
wire  [1:0]  col_out_633;
wire  [1:0]  col_out_634;
wire  [1:0]  col_out_635;
wire  [1:0]  col_out_636;
wire  [1:0]  col_out_637;
wire  [1:0]  col_out_638;
wire  [1:0]  col_out_639;
wire  [1:0]  col_out_640;
wire  [1:0]  col_out_641;
wire  [1:0]  col_out_642;
wire  [1:0]  col_out_643;
wire  [1:0]  col_out_644;
wire  [1:0]  col_out_645;
wire  [1:0]  col_out_646;
wire  [1:0]  col_out_647;
wire  [1:0]  col_out_648;
wire  [1:0]  col_out_649;
wire  [1:0]  col_out_650;
wire  [1:0]  col_out_651;
wire  [1:0]  col_out_652;
wire  [1:0]  col_out_653;
wire  [1:0]  col_out_654;
wire  [1:0]  col_out_655;
wire  [1:0]  col_out_656;
wire  [1:0]  col_out_657;
wire  [1:0]  col_out_658;
wire  [1:0]  col_out_659;
wire  [1:0]  col_out_660;
wire  [1:0]  col_out_661;
wire  [1:0]  col_out_662;
wire  [1:0]  col_out_663;
wire  [1:0]  col_out_664;
wire  [1:0]  col_out_665;
wire  [1:0]  col_out_666;
wire  [1:0]  col_out_667;
wire  [1:0]  col_out_668;
wire  [1:0]  col_out_669;
wire  [1:0]  col_out_670;
wire  [1:0]  col_out_671;
wire  [1:0]  col_out_672;
wire  [1:0]  col_out_673;
wire  [1:0]  col_out_674;
wire  [1:0]  col_out_675;
wire  [1:0]  col_out_676;
wire  [1:0]  col_out_677;
wire  [1:0]  col_out_678;
wire  [1:0]  col_out_679;
wire  [1:0]  col_out_680;
wire  [1:0]  col_out_681;
wire  [1:0]  col_out_682;
wire  [1:0]  col_out_683;
wire  [1:0]  col_out_684;
wire  [1:0]  col_out_685;
wire  [1:0]  col_out_686;
wire  [1:0]  col_out_687;
wire  [1:0]  col_out_688;
wire  [1:0]  col_out_689;
wire  [1:0]  col_out_690;
wire  [1:0]  col_out_691;
wire  [1:0]  col_out_692;
wire  [1:0]  col_out_693;
wire  [1:0]  col_out_694;
wire  [1:0]  col_out_695;
wire  [1:0]  col_out_696;
wire  [1:0]  col_out_697;
wire  [1:0]  col_out_698;
wire  [1:0]  col_out_699;
wire  [1:0]  col_out_700;
wire  [1:0]  col_out_701;
wire  [1:0]  col_out_702;
wire  [1:0]  col_out_703;
wire  [1:0]  col_out_704;
wire  [1:0]  col_out_705;
wire  [1:0]  col_out_706;
wire  [1:0]  col_out_707;
wire  [1:0]  col_out_708;
wire  [1:0]  col_out_709;
wire  [1:0]  col_out_710;
wire  [1:0]  col_out_711;
wire  [1:0]  col_out_712;
wire  [1:0]  col_out_713;
wire  [1:0]  col_out_714;
wire  [1:0]  col_out_715;
wire  [1:0]  col_out_716;
wire  [1:0]  col_out_717;
wire  [1:0]  col_out_718;
wire  [1:0]  col_out_719;
wire  [1:0]  col_out_720;
wire  [1:0]  col_out_721;
wire  [1:0]  col_out_722;
wire  [1:0]  col_out_723;
wire  [1:0]  col_out_724;
wire  [1:0]  col_out_725;
wire  [1:0]  col_out_726;
wire  [1:0]  col_out_727;
wire  [1:0]  col_out_728;
wire  [1:0]  col_out_729;
wire  [1:0]  col_out_730;
wire  [1:0]  col_out_731;
wire  [1:0]  col_out_732;
wire  [1:0]  col_out_733;
wire  [1:0]  col_out_734;
wire  [1:0]  col_out_735;
wire  [1:0]  col_out_736;
wire  [1:0]  col_out_737;
wire  [1:0]  col_out_738;
wire  [1:0]  col_out_739;
wire  [1:0]  col_out_740;
wire  [1:0]  col_out_741;
wire  [1:0]  col_out_742;
wire  [1:0]  col_out_743;
wire  [1:0]  col_out_744;
wire  [1:0]  col_out_745;
wire  [1:0]  col_out_746;
wire  [1:0]  col_out_747;
wire  [1:0]  col_out_748;
wire  [1:0]  col_out_749;
wire  [1:0]  col_out_750;
wire  [1:0]  col_out_751;
wire  [1:0]  col_out_752;
wire  [1:0]  col_out_753;
wire  [1:0]  col_out_754;
wire  [1:0]  col_out_755;
wire  [1:0]  col_out_756;
wire  [1:0]  col_out_757;
wire  [1:0]  col_out_758;
wire  [1:0]  col_out_759;
wire  [1:0]  col_out_760;
wire  [1:0]  col_out_761;
wire  [1:0]  col_out_762;
wire  [1:0]  col_out_763;
wire  [1:0]  col_out_764;
wire  [1:0]  col_out_765;
wire  [1:0]  col_out_766;
wire  [1:0]  col_out_767;
wire  [1:0]  col_out_768;
wire  [1:0]  col_out_769;
wire  [1:0]  col_out_770;
wire  [1:0]  col_out_771;
wire  [1:0]  col_out_772;
wire  [1:0]  col_out_773;
wire  [1:0]  col_out_774;
wire  [1:0]  col_out_775;
wire  [1:0]  col_out_776;
wire  [1:0]  col_out_777;
wire  [1:0]  col_out_778;
wire  [1:0]  col_out_779;
wire  [1:0]  col_out_780;
wire  [1:0]  col_out_781;
wire  [1:0]  col_out_782;
wire  [1:0]  col_out_783;
wire  [1:0]  col_out_784;
wire  [1:0]  col_out_785;
wire  [1:0]  col_out_786;
wire  [1:0]  col_out_787;
wire  [1:0]  col_out_788;
wire  [1:0]  col_out_789;
wire  [1:0]  col_out_790;
wire  [1:0]  col_out_791;
wire  [1:0]  col_out_792;
wire  [1:0]  col_out_793;
wire  [1:0]  col_out_794;
wire  [1:0]  col_out_795;
wire  [1:0]  col_out_796;
wire  [1:0]  col_out_797;
wire  [1:0]  col_out_798;
wire  [1:0]  col_out_799;
wire  [1:0]  col_out_800;
wire  [1:0]  col_out_801;
wire  [1:0]  col_out_802;
wire  [1:0]  col_out_803;
wire  [1:0]  col_out_804;
wire  [1:0]  col_out_805;
wire  [1:0]  col_out_806;
wire  [1:0]  col_out_807;
wire  [1:0]  col_out_808;
wire  [1:0]  col_out_809;
wire  [1:0]  col_out_810;
wire  [1:0]  col_out_811;
wire  [1:0]  col_out_812;
wire  [1:0]  col_out_813;
wire  [1:0]  col_out_814;
wire  [1:0]  col_out_815;
wire  [1:0]  col_out_816;
wire  [1:0]  col_out_817;
wire  [1:0]  col_out_818;
wire  [1:0]  col_out_819;
wire  [1:0]  col_out_820;
wire  [1:0]  col_out_821;
wire  [1:0]  col_out_822;
wire  [1:0]  col_out_823;
wire  [1:0]  col_out_824;
wire  [1:0]  col_out_825;
wire  [1:0]  col_out_826;
wire  [1:0]  col_out_827;
wire  [1:0]  col_out_828;
wire  [1:0]  col_out_829;
wire  [1:0]  col_out_830;
wire  [1:0]  col_out_831;
wire  [1:0]  col_out_832;
wire  [1:0]  col_out_833;
wire  [1:0]  col_out_834;
wire  [1:0]  col_out_835;
wire  [1:0]  col_out_836;
wire  [1:0]  col_out_837;
wire  [1:0]  col_out_838;
wire  [1:0]  col_out_839;
wire  [1:0]  col_out_840;
wire  [1:0]  col_out_841;
wire  [1:0]  col_out_842;
wire  [1:0]  col_out_843;
wire  [1:0]  col_out_844;
wire  [1:0]  col_out_845;
wire  [1:0]  col_out_846;
wire  [1:0]  col_out_847;
wire  [1:0]  col_out_848;
wire  [1:0]  col_out_849;
wire  [1:0]  col_out_850;
wire  [1:0]  col_out_851;
wire  [1:0]  col_out_852;
wire  [1:0]  col_out_853;
wire  [1:0]  col_out_854;
wire  [1:0]  col_out_855;
wire  [1:0]  col_out_856;
wire  [1:0]  col_out_857;
wire  [1:0]  col_out_858;
wire  [1:0]  col_out_859;
wire  [1:0]  col_out_860;
wire  [1:0]  col_out_861;
wire  [1:0]  col_out_862;
wire  [1:0]  col_out_863;
wire  [1:0]  col_out_864;
wire  [1:0]  col_out_865;
wire  [1:0]  col_out_866;
wire  [1:0]  col_out_867;
wire  [1:0]  col_out_868;
wire  [1:0]  col_out_869;
wire  [1:0]  col_out_870;
wire  [1:0]  col_out_871;
wire  [1:0]  col_out_872;
wire  [1:0]  col_out_873;
wire  [1:0]  col_out_874;
wire  [1:0]  col_out_875;
wire  [1:0]  col_out_876;
wire  [1:0]  col_out_877;
wire  [1:0]  col_out_878;
wire  [1:0]  col_out_879;
wire  [1:0]  col_out_880;
wire  [1:0]  col_out_881;
wire  [1:0]  col_out_882;
wire  [1:0]  col_out_883;
wire  [1:0]  col_out_884;
wire  [1:0]  col_out_885;
wire  [1:0]  col_out_886;
wire  [1:0]  col_out_887;
wire  [1:0]  col_out_888;
wire  [1:0]  col_out_889;
wire  [1:0]  col_out_890;
wire  [1:0]  col_out_891;
wire  [1:0]  col_out_892;
wire  [1:0]  col_out_893;
wire  [1:0]  col_out_894;
wire  [1:0]  col_out_895;
wire  [1:0]  col_out_896;
wire  [1:0]  col_out_897;
wire  [1:0]  col_out_898;
wire  [1:0]  col_out_899;
wire  [1:0]  col_out_900;
wire  [1:0]  col_out_901;
wire  [1:0]  col_out_902;
wire  [1:0]  col_out_903;
wire  [1:0]  col_out_904;
wire  [1:0]  col_out_905;
wire  [1:0]  col_out_906;
wire  [1:0]  col_out_907;
wire  [1:0]  col_out_908;
wire  [1:0]  col_out_909;
wire  [1:0]  col_out_910;
wire  [1:0]  col_out_911;
wire  [1:0]  col_out_912;
wire  [1:0]  col_out_913;
wire  [1:0]  col_out_914;
wire  [1:0]  col_out_915;
wire  [1:0]  col_out_916;
wire  [1:0]  col_out_917;
wire  [1:0]  col_out_918;
wire  [1:0]  col_out_919;
wire  [1:0]  col_out_920;
wire  [1:0]  col_out_921;
wire  [1:0]  col_out_922;
wire  [1:0]  col_out_923;
wire  [1:0]  col_out_924;
wire  [1:0]  col_out_925;
wire  [1:0]  col_out_926;
wire  [1:0]  col_out_927;
wire  [1:0]  col_out_928;
wire  [1:0]  col_out_929;
wire  [1:0]  col_out_930;
wire  [1:0]  col_out_931;
wire  [1:0]  col_out_932;
wire  [1:0]  col_out_933;
wire  [1:0]  col_out_934;
wire  [1:0]  col_out_935;
wire  [1:0]  col_out_936;
wire  [1:0]  col_out_937;
wire  [1:0]  col_out_938;
wire  [1:0]  col_out_939;
wire  [1:0]  col_out_940;
wire  [1:0]  col_out_941;
wire  [1:0]  col_out_942;
wire  [1:0]  col_out_943;
wire  [1:0]  col_out_944;
wire  [1:0]  col_out_945;
wire  [1:0]  col_out_946;
wire  [1:0]  col_out_947;
wire  [1:0]  col_out_948;
wire  [1:0]  col_out_949;
wire  [1:0]  col_out_950;
wire  [1:0]  col_out_951;
wire  [1:0]  col_out_952;
wire  [1:0]  col_out_953;
wire  [1:0]  col_out_954;
wire  [1:0]  col_out_955;
wire  [1:0]  col_out_956;
wire  [1:0]  col_out_957;
wire  [1:0]  col_out_958;
wire  [1:0]  col_out_959;
wire  [1:0]  col_out_960;
wire  [1:0]  col_out_961;
wire  [1:0]  col_out_962;
wire  [1:0]  col_out_963;
wire  [1:0]  col_out_964;
wire  [1:0]  col_out_965;
wire  [1:0]  col_out_966;
wire  [1:0]  col_out_967;
wire  [1:0]  col_out_968;
wire  [1:0]  col_out_969;
wire  [1:0]  col_out_970;
wire  [1:0]  col_out_971;
wire  [1:0]  col_out_972;
wire  [1:0]  col_out_973;
wire  [1:0]  col_out_974;
wire  [1:0]  col_out_975;
wire  [1:0]  col_out_976;
wire  [1:0]  col_out_977;
wire  [1:0]  col_out_978;
wire  [1:0]  col_out_979;
wire  [1:0]  col_out_980;
wire  [1:0]  col_out_981;
wire  [1:0]  col_out_982;
wire  [1:0]  col_out_983;
wire  [1:0]  col_out_984;
wire  [1:0]  col_out_985;
wire  [1:0]  col_out_986;
wire  [1:0]  col_out_987;
wire  [1:0]  col_out_988;
wire  [1:0]  col_out_989;
wire  [1:0]  col_out_990;
wire  [1:0]  col_out_991;
wire  [1:0]  col_out_992;
wire  [1:0]  col_out_993;
wire  [1:0]  col_out_994;
wire  [1:0]  col_out_995;
wire  [1:0]  col_out_996;
wire  [1:0]  col_out_997;
wire  [1:0]  col_out_998;
wire  [1:0]  col_out_999;
wire  [1:0]  col_out_1000;
wire  [1:0]  col_out_1001;
wire  [1:0]  col_out_1002;
wire  [1:0]  col_out_1003;
wire  [1:0]  col_out_1004;
wire  [1:0]  col_out_1005;
wire  [1:0]  col_out_1006;
wire  [1:0]  col_out_1007;
wire  [1:0]  col_out_1008;
wire  [1:0]  col_out_1009;
wire  [1:0]  col_out_1010;
wire  [1:0]  col_out_1011;
wire  [1:0]  col_out_1012;
wire  [1:0]  col_out_1013;
wire  [1:0]  col_out_1014;
wire  [1:0]  col_out_1015;
wire  [1:0]  col_out_1016;
wire  [1:0]  col_out_1017;
wire  [1:0]  col_out_1018;
wire  [1:0]  col_out_1019;
wire  [1:0]  col_out_1020;
wire  [1:0]  col_out_1021;
wire  [1:0]  col_out_1022;
wire  [1:0]  col_out_1023;
wire  [1:0]  col_out_1024;

compressor_array_3_2_1024  u_compressor_array_3_2_1024 (
    .col_in_0                ( col_in_0       ),
    .col_in_1                ( col_in_1       ),
    .col_in_2                ( col_in_2       ),
    .col_in_3                ( col_in_3       ),
    .col_in_4                ( col_in_4       ),
    .col_in_5                ( col_in_5       ),
    .col_in_6                ( col_in_6       ),
    .col_in_7                ( col_in_7       ),
    .col_in_8                ( col_in_8       ),
    .col_in_9                ( col_in_9       ),
    .col_in_10               ( col_in_10      ),
    .col_in_11               ( col_in_11      ),
    .col_in_12               ( col_in_12      ),
    .col_in_13               ( col_in_13      ),
    .col_in_14               ( col_in_14      ),
    .col_in_15               ( col_in_15      ),
    .col_in_16               ( col_in_16      ),
    .col_in_17               ( col_in_17      ),
    .col_in_18               ( col_in_18      ),
    .col_in_19               ( col_in_19      ),
    .col_in_20               ( col_in_20      ),
    .col_in_21               ( col_in_21      ),
    .col_in_22               ( col_in_22      ),
    .col_in_23               ( col_in_23      ),
    .col_in_24               ( col_in_24      ),
    .col_in_25               ( col_in_25      ),
    .col_in_26               ( col_in_26      ),
    .col_in_27               ( col_in_27      ),
    .col_in_28               ( col_in_28      ),
    .col_in_29               ( col_in_29      ),
    .col_in_30               ( col_in_30      ),
    .col_in_31               ( col_in_31      ),
    .col_in_32               ( col_in_32      ),
    .col_in_33               ( col_in_33      ),
    .col_in_34               ( col_in_34      ),
    .col_in_35               ( col_in_35      ),
    .col_in_36               ( col_in_36      ),
    .col_in_37               ( col_in_37      ),
    .col_in_38               ( col_in_38      ),
    .col_in_39               ( col_in_39      ),
    .col_in_40               ( col_in_40      ),
    .col_in_41               ( col_in_41      ),
    .col_in_42               ( col_in_42      ),
    .col_in_43               ( col_in_43      ),
    .col_in_44               ( col_in_44      ),
    .col_in_45               ( col_in_45      ),
    .col_in_46               ( col_in_46      ),
    .col_in_47               ( col_in_47      ),
    .col_in_48               ( col_in_48      ),
    .col_in_49               ( col_in_49      ),
    .col_in_50               ( col_in_50      ),
    .col_in_51               ( col_in_51      ),
    .col_in_52               ( col_in_52      ),
    .col_in_53               ( col_in_53      ),
    .col_in_54               ( col_in_54      ),
    .col_in_55               ( col_in_55      ),
    .col_in_56               ( col_in_56      ),
    .col_in_57               ( col_in_57      ),
    .col_in_58               ( col_in_58      ),
    .col_in_59               ( col_in_59      ),
    .col_in_60               ( col_in_60      ),
    .col_in_61               ( col_in_61      ),
    .col_in_62               ( col_in_62      ),
    .col_in_63               ( col_in_63      ),
    .col_in_64               ( col_in_64      ),
    .col_in_65               ( col_in_65      ),
    .col_in_66               ( col_in_66      ),
    .col_in_67               ( col_in_67      ),
    .col_in_68               ( col_in_68      ),
    .col_in_69               ( col_in_69      ),
    .col_in_70               ( col_in_70      ),
    .col_in_71               ( col_in_71      ),
    .col_in_72               ( col_in_72      ),
    .col_in_73               ( col_in_73      ),
    .col_in_74               ( col_in_74      ),
    .col_in_75               ( col_in_75      ),
    .col_in_76               ( col_in_76      ),
    .col_in_77               ( col_in_77      ),
    .col_in_78               ( col_in_78      ),
    .col_in_79               ( col_in_79      ),
    .col_in_80               ( col_in_80      ),
    .col_in_81               ( col_in_81      ),
    .col_in_82               ( col_in_82      ),
    .col_in_83               ( col_in_83      ),
    .col_in_84               ( col_in_84      ),
    .col_in_85               ( col_in_85      ),
    .col_in_86               ( col_in_86      ),
    .col_in_87               ( col_in_87      ),
    .col_in_88               ( col_in_88      ),
    .col_in_89               ( col_in_89      ),
    .col_in_90               ( col_in_90      ),
    .col_in_91               ( col_in_91      ),
    .col_in_92               ( col_in_92      ),
    .col_in_93               ( col_in_93      ),
    .col_in_94               ( col_in_94      ),
    .col_in_95               ( col_in_95      ),
    .col_in_96               ( col_in_96      ),
    .col_in_97               ( col_in_97      ),
    .col_in_98               ( col_in_98      ),
    .col_in_99               ( col_in_99      ),
    .col_in_100              ( col_in_100     ),
    .col_in_101              ( col_in_101     ),
    .col_in_102              ( col_in_102     ),
    .col_in_103              ( col_in_103     ),
    .col_in_104              ( col_in_104     ),
    .col_in_105              ( col_in_105     ),
    .col_in_106              ( col_in_106     ),
    .col_in_107              ( col_in_107     ),
    .col_in_108              ( col_in_108     ),
    .col_in_109              ( col_in_109     ),
    .col_in_110              ( col_in_110     ),
    .col_in_111              ( col_in_111     ),
    .col_in_112              ( col_in_112     ),
    .col_in_113              ( col_in_113     ),
    .col_in_114              ( col_in_114     ),
    .col_in_115              ( col_in_115     ),
    .col_in_116              ( col_in_116     ),
    .col_in_117              ( col_in_117     ),
    .col_in_118              ( col_in_118     ),
    .col_in_119              ( col_in_119     ),
    .col_in_120              ( col_in_120     ),
    .col_in_121              ( col_in_121     ),
    .col_in_122              ( col_in_122     ),
    .col_in_123              ( col_in_123     ),
    .col_in_124              ( col_in_124     ),
    .col_in_125              ( col_in_125     ),
    .col_in_126              ( col_in_126     ),
    .col_in_127              ( col_in_127     ),
    .col_in_128              ( col_in_128     ),
    .col_in_129              ( col_in_129     ),
    .col_in_130              ( col_in_130     ),
    .col_in_131              ( col_in_131     ),
    .col_in_132              ( col_in_132     ),
    .col_in_133              ( col_in_133     ),
    .col_in_134              ( col_in_134     ),
    .col_in_135              ( col_in_135     ),
    .col_in_136              ( col_in_136     ),
    .col_in_137              ( col_in_137     ),
    .col_in_138              ( col_in_138     ),
    .col_in_139              ( col_in_139     ),
    .col_in_140              ( col_in_140     ),
    .col_in_141              ( col_in_141     ),
    .col_in_142              ( col_in_142     ),
    .col_in_143              ( col_in_143     ),
    .col_in_144              ( col_in_144     ),
    .col_in_145              ( col_in_145     ),
    .col_in_146              ( col_in_146     ),
    .col_in_147              ( col_in_147     ),
    .col_in_148              ( col_in_148     ),
    .col_in_149              ( col_in_149     ),
    .col_in_150              ( col_in_150     ),
    .col_in_151              ( col_in_151     ),
    .col_in_152              ( col_in_152     ),
    .col_in_153              ( col_in_153     ),
    .col_in_154              ( col_in_154     ),
    .col_in_155              ( col_in_155     ),
    .col_in_156              ( col_in_156     ),
    .col_in_157              ( col_in_157     ),
    .col_in_158              ( col_in_158     ),
    .col_in_159              ( col_in_159     ),
    .col_in_160              ( col_in_160     ),
    .col_in_161              ( col_in_161     ),
    .col_in_162              ( col_in_162     ),
    .col_in_163              ( col_in_163     ),
    .col_in_164              ( col_in_164     ),
    .col_in_165              ( col_in_165     ),
    .col_in_166              ( col_in_166     ),
    .col_in_167              ( col_in_167     ),
    .col_in_168              ( col_in_168     ),
    .col_in_169              ( col_in_169     ),
    .col_in_170              ( col_in_170     ),
    .col_in_171              ( col_in_171     ),
    .col_in_172              ( col_in_172     ),
    .col_in_173              ( col_in_173     ),
    .col_in_174              ( col_in_174     ),
    .col_in_175              ( col_in_175     ),
    .col_in_176              ( col_in_176     ),
    .col_in_177              ( col_in_177     ),
    .col_in_178              ( col_in_178     ),
    .col_in_179              ( col_in_179     ),
    .col_in_180              ( col_in_180     ),
    .col_in_181              ( col_in_181     ),
    .col_in_182              ( col_in_182     ),
    .col_in_183              ( col_in_183     ),
    .col_in_184              ( col_in_184     ),
    .col_in_185              ( col_in_185     ),
    .col_in_186              ( col_in_186     ),
    .col_in_187              ( col_in_187     ),
    .col_in_188              ( col_in_188     ),
    .col_in_189              ( col_in_189     ),
    .col_in_190              ( col_in_190     ),
    .col_in_191              ( col_in_191     ),
    .col_in_192              ( col_in_192     ),
    .col_in_193              ( col_in_193     ),
    .col_in_194              ( col_in_194     ),
    .col_in_195              ( col_in_195     ),
    .col_in_196              ( col_in_196     ),
    .col_in_197              ( col_in_197     ),
    .col_in_198              ( col_in_198     ),
    .col_in_199              ( col_in_199     ),
    .col_in_200              ( col_in_200     ),
    .col_in_201              ( col_in_201     ),
    .col_in_202              ( col_in_202     ),
    .col_in_203              ( col_in_203     ),
    .col_in_204              ( col_in_204     ),
    .col_in_205              ( col_in_205     ),
    .col_in_206              ( col_in_206     ),
    .col_in_207              ( col_in_207     ),
    .col_in_208              ( col_in_208     ),
    .col_in_209              ( col_in_209     ),
    .col_in_210              ( col_in_210     ),
    .col_in_211              ( col_in_211     ),
    .col_in_212              ( col_in_212     ),
    .col_in_213              ( col_in_213     ),
    .col_in_214              ( col_in_214     ),
    .col_in_215              ( col_in_215     ),
    .col_in_216              ( col_in_216     ),
    .col_in_217              ( col_in_217     ),
    .col_in_218              ( col_in_218     ),
    .col_in_219              ( col_in_219     ),
    .col_in_220              ( col_in_220     ),
    .col_in_221              ( col_in_221     ),
    .col_in_222              ( col_in_222     ),
    .col_in_223              ( col_in_223     ),
    .col_in_224              ( col_in_224     ),
    .col_in_225              ( col_in_225     ),
    .col_in_226              ( col_in_226     ),
    .col_in_227              ( col_in_227     ),
    .col_in_228              ( col_in_228     ),
    .col_in_229              ( col_in_229     ),
    .col_in_230              ( col_in_230     ),
    .col_in_231              ( col_in_231     ),
    .col_in_232              ( col_in_232     ),
    .col_in_233              ( col_in_233     ),
    .col_in_234              ( col_in_234     ),
    .col_in_235              ( col_in_235     ),
    .col_in_236              ( col_in_236     ),
    .col_in_237              ( col_in_237     ),
    .col_in_238              ( col_in_238     ),
    .col_in_239              ( col_in_239     ),
    .col_in_240              ( col_in_240     ),
    .col_in_241              ( col_in_241     ),
    .col_in_242              ( col_in_242     ),
    .col_in_243              ( col_in_243     ),
    .col_in_244              ( col_in_244     ),
    .col_in_245              ( col_in_245     ),
    .col_in_246              ( col_in_246     ),
    .col_in_247              ( col_in_247     ),
    .col_in_248              ( col_in_248     ),
    .col_in_249              ( col_in_249     ),
    .col_in_250              ( col_in_250     ),
    .col_in_251              ( col_in_251     ),
    .col_in_252              ( col_in_252     ),
    .col_in_253              ( col_in_253     ),
    .col_in_254              ( col_in_254     ),
    .col_in_255              ( col_in_255     ),
    .col_in_256              ( col_in_256     ),
    .col_in_257              ( col_in_257     ),
    .col_in_258              ( col_in_258     ),
    .col_in_259              ( col_in_259     ),
    .col_in_260              ( col_in_260     ),
    .col_in_261              ( col_in_261     ),
    .col_in_262              ( col_in_262     ),
    .col_in_263              ( col_in_263     ),
    .col_in_264              ( col_in_264     ),
    .col_in_265              ( col_in_265     ),
    .col_in_266              ( col_in_266     ),
    .col_in_267              ( col_in_267     ),
    .col_in_268              ( col_in_268     ),
    .col_in_269              ( col_in_269     ),
    .col_in_270              ( col_in_270     ),
    .col_in_271              ( col_in_271     ),
    .col_in_272              ( col_in_272     ),
    .col_in_273              ( col_in_273     ),
    .col_in_274              ( col_in_274     ),
    .col_in_275              ( col_in_275     ),
    .col_in_276              ( col_in_276     ),
    .col_in_277              ( col_in_277     ),
    .col_in_278              ( col_in_278     ),
    .col_in_279              ( col_in_279     ),
    .col_in_280              ( col_in_280     ),
    .col_in_281              ( col_in_281     ),
    .col_in_282              ( col_in_282     ),
    .col_in_283              ( col_in_283     ),
    .col_in_284              ( col_in_284     ),
    .col_in_285              ( col_in_285     ),
    .col_in_286              ( col_in_286     ),
    .col_in_287              ( col_in_287     ),
    .col_in_288              ( col_in_288     ),
    .col_in_289              ( col_in_289     ),
    .col_in_290              ( col_in_290     ),
    .col_in_291              ( col_in_291     ),
    .col_in_292              ( col_in_292     ),
    .col_in_293              ( col_in_293     ),
    .col_in_294              ( col_in_294     ),
    .col_in_295              ( col_in_295     ),
    .col_in_296              ( col_in_296     ),
    .col_in_297              ( col_in_297     ),
    .col_in_298              ( col_in_298     ),
    .col_in_299              ( col_in_299     ),
    .col_in_300              ( col_in_300     ),
    .col_in_301              ( col_in_301     ),
    .col_in_302              ( col_in_302     ),
    .col_in_303              ( col_in_303     ),
    .col_in_304              ( col_in_304     ),
    .col_in_305              ( col_in_305     ),
    .col_in_306              ( col_in_306     ),
    .col_in_307              ( col_in_307     ),
    .col_in_308              ( col_in_308     ),
    .col_in_309              ( col_in_309     ),
    .col_in_310              ( col_in_310     ),
    .col_in_311              ( col_in_311     ),
    .col_in_312              ( col_in_312     ),
    .col_in_313              ( col_in_313     ),
    .col_in_314              ( col_in_314     ),
    .col_in_315              ( col_in_315     ),
    .col_in_316              ( col_in_316     ),
    .col_in_317              ( col_in_317     ),
    .col_in_318              ( col_in_318     ),
    .col_in_319              ( col_in_319     ),
    .col_in_320              ( col_in_320     ),
    .col_in_321              ( col_in_321     ),
    .col_in_322              ( col_in_322     ),
    .col_in_323              ( col_in_323     ),
    .col_in_324              ( col_in_324     ),
    .col_in_325              ( col_in_325     ),
    .col_in_326              ( col_in_326     ),
    .col_in_327              ( col_in_327     ),
    .col_in_328              ( col_in_328     ),
    .col_in_329              ( col_in_329     ),
    .col_in_330              ( col_in_330     ),
    .col_in_331              ( col_in_331     ),
    .col_in_332              ( col_in_332     ),
    .col_in_333              ( col_in_333     ),
    .col_in_334              ( col_in_334     ),
    .col_in_335              ( col_in_335     ),
    .col_in_336              ( col_in_336     ),
    .col_in_337              ( col_in_337     ),
    .col_in_338              ( col_in_338     ),
    .col_in_339              ( col_in_339     ),
    .col_in_340              ( col_in_340     ),
    .col_in_341              ( col_in_341     ),
    .col_in_342              ( col_in_342     ),
    .col_in_343              ( col_in_343     ),
    .col_in_344              ( col_in_344     ),
    .col_in_345              ( col_in_345     ),
    .col_in_346              ( col_in_346     ),
    .col_in_347              ( col_in_347     ),
    .col_in_348              ( col_in_348     ),
    .col_in_349              ( col_in_349     ),
    .col_in_350              ( col_in_350     ),
    .col_in_351              ( col_in_351     ),
    .col_in_352              ( col_in_352     ),
    .col_in_353              ( col_in_353     ),
    .col_in_354              ( col_in_354     ),
    .col_in_355              ( col_in_355     ),
    .col_in_356              ( col_in_356     ),
    .col_in_357              ( col_in_357     ),
    .col_in_358              ( col_in_358     ),
    .col_in_359              ( col_in_359     ),
    .col_in_360              ( col_in_360     ),
    .col_in_361              ( col_in_361     ),
    .col_in_362              ( col_in_362     ),
    .col_in_363              ( col_in_363     ),
    .col_in_364              ( col_in_364     ),
    .col_in_365              ( col_in_365     ),
    .col_in_366              ( col_in_366     ),
    .col_in_367              ( col_in_367     ),
    .col_in_368              ( col_in_368     ),
    .col_in_369              ( col_in_369     ),
    .col_in_370              ( col_in_370     ),
    .col_in_371              ( col_in_371     ),
    .col_in_372              ( col_in_372     ),
    .col_in_373              ( col_in_373     ),
    .col_in_374              ( col_in_374     ),
    .col_in_375              ( col_in_375     ),
    .col_in_376              ( col_in_376     ),
    .col_in_377              ( col_in_377     ),
    .col_in_378              ( col_in_378     ),
    .col_in_379              ( col_in_379     ),
    .col_in_380              ( col_in_380     ),
    .col_in_381              ( col_in_381     ),
    .col_in_382              ( col_in_382     ),
    .col_in_383              ( col_in_383     ),
    .col_in_384              ( col_in_384     ),
    .col_in_385              ( col_in_385     ),
    .col_in_386              ( col_in_386     ),
    .col_in_387              ( col_in_387     ),
    .col_in_388              ( col_in_388     ),
    .col_in_389              ( col_in_389     ),
    .col_in_390              ( col_in_390     ),
    .col_in_391              ( col_in_391     ),
    .col_in_392              ( col_in_392     ),
    .col_in_393              ( col_in_393     ),
    .col_in_394              ( col_in_394     ),
    .col_in_395              ( col_in_395     ),
    .col_in_396              ( col_in_396     ),
    .col_in_397              ( col_in_397     ),
    .col_in_398              ( col_in_398     ),
    .col_in_399              ( col_in_399     ),
    .col_in_400              ( col_in_400     ),
    .col_in_401              ( col_in_401     ),
    .col_in_402              ( col_in_402     ),
    .col_in_403              ( col_in_403     ),
    .col_in_404              ( col_in_404     ),
    .col_in_405              ( col_in_405     ),
    .col_in_406              ( col_in_406     ),
    .col_in_407              ( col_in_407     ),
    .col_in_408              ( col_in_408     ),
    .col_in_409              ( col_in_409     ),
    .col_in_410              ( col_in_410     ),
    .col_in_411              ( col_in_411     ),
    .col_in_412              ( col_in_412     ),
    .col_in_413              ( col_in_413     ),
    .col_in_414              ( col_in_414     ),
    .col_in_415              ( col_in_415     ),
    .col_in_416              ( col_in_416     ),
    .col_in_417              ( col_in_417     ),
    .col_in_418              ( col_in_418     ),
    .col_in_419              ( col_in_419     ),
    .col_in_420              ( col_in_420     ),
    .col_in_421              ( col_in_421     ),
    .col_in_422              ( col_in_422     ),
    .col_in_423              ( col_in_423     ),
    .col_in_424              ( col_in_424     ),
    .col_in_425              ( col_in_425     ),
    .col_in_426              ( col_in_426     ),
    .col_in_427              ( col_in_427     ),
    .col_in_428              ( col_in_428     ),
    .col_in_429              ( col_in_429     ),
    .col_in_430              ( col_in_430     ),
    .col_in_431              ( col_in_431     ),
    .col_in_432              ( col_in_432     ),
    .col_in_433              ( col_in_433     ),
    .col_in_434              ( col_in_434     ),
    .col_in_435              ( col_in_435     ),
    .col_in_436              ( col_in_436     ),
    .col_in_437              ( col_in_437     ),
    .col_in_438              ( col_in_438     ),
    .col_in_439              ( col_in_439     ),
    .col_in_440              ( col_in_440     ),
    .col_in_441              ( col_in_441     ),
    .col_in_442              ( col_in_442     ),
    .col_in_443              ( col_in_443     ),
    .col_in_444              ( col_in_444     ),
    .col_in_445              ( col_in_445     ),
    .col_in_446              ( col_in_446     ),
    .col_in_447              ( col_in_447     ),
    .col_in_448              ( col_in_448     ),
    .col_in_449              ( col_in_449     ),
    .col_in_450              ( col_in_450     ),
    .col_in_451              ( col_in_451     ),
    .col_in_452              ( col_in_452     ),
    .col_in_453              ( col_in_453     ),
    .col_in_454              ( col_in_454     ),
    .col_in_455              ( col_in_455     ),
    .col_in_456              ( col_in_456     ),
    .col_in_457              ( col_in_457     ),
    .col_in_458              ( col_in_458     ),
    .col_in_459              ( col_in_459     ),
    .col_in_460              ( col_in_460     ),
    .col_in_461              ( col_in_461     ),
    .col_in_462              ( col_in_462     ),
    .col_in_463              ( col_in_463     ),
    .col_in_464              ( col_in_464     ),
    .col_in_465              ( col_in_465     ),
    .col_in_466              ( col_in_466     ),
    .col_in_467              ( col_in_467     ),
    .col_in_468              ( col_in_468     ),
    .col_in_469              ( col_in_469     ),
    .col_in_470              ( col_in_470     ),
    .col_in_471              ( col_in_471     ),
    .col_in_472              ( col_in_472     ),
    .col_in_473              ( col_in_473     ),
    .col_in_474              ( col_in_474     ),
    .col_in_475              ( col_in_475     ),
    .col_in_476              ( col_in_476     ),
    .col_in_477              ( col_in_477     ),
    .col_in_478              ( col_in_478     ),
    .col_in_479              ( col_in_479     ),
    .col_in_480              ( col_in_480     ),
    .col_in_481              ( col_in_481     ),
    .col_in_482              ( col_in_482     ),
    .col_in_483              ( col_in_483     ),
    .col_in_484              ( col_in_484     ),
    .col_in_485              ( col_in_485     ),
    .col_in_486              ( col_in_486     ),
    .col_in_487              ( col_in_487     ),
    .col_in_488              ( col_in_488     ),
    .col_in_489              ( col_in_489     ),
    .col_in_490              ( col_in_490     ),
    .col_in_491              ( col_in_491     ),
    .col_in_492              ( col_in_492     ),
    .col_in_493              ( col_in_493     ),
    .col_in_494              ( col_in_494     ),
    .col_in_495              ( col_in_495     ),
    .col_in_496              ( col_in_496     ),
    .col_in_497              ( col_in_497     ),
    .col_in_498              ( col_in_498     ),
    .col_in_499              ( col_in_499     ),
    .col_in_500              ( col_in_500     ),
    .col_in_501              ( col_in_501     ),
    .col_in_502              ( col_in_502     ),
    .col_in_503              ( col_in_503     ),
    .col_in_504              ( col_in_504     ),
    .col_in_505              ( col_in_505     ),
    .col_in_506              ( col_in_506     ),
    .col_in_507              ( col_in_507     ),
    .col_in_508              ( col_in_508     ),
    .col_in_509              ( col_in_509     ),
    .col_in_510              ( col_in_510     ),
    .col_in_511              ( col_in_511     ),
    .col_in_512              ( col_in_512     ),
    .col_in_513              ( col_in_513     ),
    .col_in_514              ( col_in_514     ),
    .col_in_515              ( col_in_515     ),
    .col_in_516              ( col_in_516     ),
    .col_in_517              ( col_in_517     ),
    .col_in_518              ( col_in_518     ),
    .col_in_519              ( col_in_519     ),
    .col_in_520              ( col_in_520     ),
    .col_in_521              ( col_in_521     ),
    .col_in_522              ( col_in_522     ),
    .col_in_523              ( col_in_523     ),
    .col_in_524              ( col_in_524     ),
    .col_in_525              ( col_in_525     ),
    .col_in_526              ( col_in_526     ),
    .col_in_527              ( col_in_527     ),
    .col_in_528              ( col_in_528     ),
    .col_in_529              ( col_in_529     ),
    .col_in_530              ( col_in_530     ),
    .col_in_531              ( col_in_531     ),
    .col_in_532              ( col_in_532     ),
    .col_in_533              ( col_in_533     ),
    .col_in_534              ( col_in_534     ),
    .col_in_535              ( col_in_535     ),
    .col_in_536              ( col_in_536     ),
    .col_in_537              ( col_in_537     ),
    .col_in_538              ( col_in_538     ),
    .col_in_539              ( col_in_539     ),
    .col_in_540              ( col_in_540     ),
    .col_in_541              ( col_in_541     ),
    .col_in_542              ( col_in_542     ),
    .col_in_543              ( col_in_543     ),
    .col_in_544              ( col_in_544     ),
    .col_in_545              ( col_in_545     ),
    .col_in_546              ( col_in_546     ),
    .col_in_547              ( col_in_547     ),
    .col_in_548              ( col_in_548     ),
    .col_in_549              ( col_in_549     ),
    .col_in_550              ( col_in_550     ),
    .col_in_551              ( col_in_551     ),
    .col_in_552              ( col_in_552     ),
    .col_in_553              ( col_in_553     ),
    .col_in_554              ( col_in_554     ),
    .col_in_555              ( col_in_555     ),
    .col_in_556              ( col_in_556     ),
    .col_in_557              ( col_in_557     ),
    .col_in_558              ( col_in_558     ),
    .col_in_559              ( col_in_559     ),
    .col_in_560              ( col_in_560     ),
    .col_in_561              ( col_in_561     ),
    .col_in_562              ( col_in_562     ),
    .col_in_563              ( col_in_563     ),
    .col_in_564              ( col_in_564     ),
    .col_in_565              ( col_in_565     ),
    .col_in_566              ( col_in_566     ),
    .col_in_567              ( col_in_567     ),
    .col_in_568              ( col_in_568     ),
    .col_in_569              ( col_in_569     ),
    .col_in_570              ( col_in_570     ),
    .col_in_571              ( col_in_571     ),
    .col_in_572              ( col_in_572     ),
    .col_in_573              ( col_in_573     ),
    .col_in_574              ( col_in_574     ),
    .col_in_575              ( col_in_575     ),
    .col_in_576              ( col_in_576     ),
    .col_in_577              ( col_in_577     ),
    .col_in_578              ( col_in_578     ),
    .col_in_579              ( col_in_579     ),
    .col_in_580              ( col_in_580     ),
    .col_in_581              ( col_in_581     ),
    .col_in_582              ( col_in_582     ),
    .col_in_583              ( col_in_583     ),
    .col_in_584              ( col_in_584     ),
    .col_in_585              ( col_in_585     ),
    .col_in_586              ( col_in_586     ),
    .col_in_587              ( col_in_587     ),
    .col_in_588              ( col_in_588     ),
    .col_in_589              ( col_in_589     ),
    .col_in_590              ( col_in_590     ),
    .col_in_591              ( col_in_591     ),
    .col_in_592              ( col_in_592     ),
    .col_in_593              ( col_in_593     ),
    .col_in_594              ( col_in_594     ),
    .col_in_595              ( col_in_595     ),
    .col_in_596              ( col_in_596     ),
    .col_in_597              ( col_in_597     ),
    .col_in_598              ( col_in_598     ),
    .col_in_599              ( col_in_599     ),
    .col_in_600              ( col_in_600     ),
    .col_in_601              ( col_in_601     ),
    .col_in_602              ( col_in_602     ),
    .col_in_603              ( col_in_603     ),
    .col_in_604              ( col_in_604     ),
    .col_in_605              ( col_in_605     ),
    .col_in_606              ( col_in_606     ),
    .col_in_607              ( col_in_607     ),
    .col_in_608              ( col_in_608     ),
    .col_in_609              ( col_in_609     ),
    .col_in_610              ( col_in_610     ),
    .col_in_611              ( col_in_611     ),
    .col_in_612              ( col_in_612     ),
    .col_in_613              ( col_in_613     ),
    .col_in_614              ( col_in_614     ),
    .col_in_615              ( col_in_615     ),
    .col_in_616              ( col_in_616     ),
    .col_in_617              ( col_in_617     ),
    .col_in_618              ( col_in_618     ),
    .col_in_619              ( col_in_619     ),
    .col_in_620              ( col_in_620     ),
    .col_in_621              ( col_in_621     ),
    .col_in_622              ( col_in_622     ),
    .col_in_623              ( col_in_623     ),
    .col_in_624              ( col_in_624     ),
    .col_in_625              ( col_in_625     ),
    .col_in_626              ( col_in_626     ),
    .col_in_627              ( col_in_627     ),
    .col_in_628              ( col_in_628     ),
    .col_in_629              ( col_in_629     ),
    .col_in_630              ( col_in_630     ),
    .col_in_631              ( col_in_631     ),
    .col_in_632              ( col_in_632     ),
    .col_in_633              ( col_in_633     ),
    .col_in_634              ( col_in_634     ),
    .col_in_635              ( col_in_635     ),
    .col_in_636              ( col_in_636     ),
    .col_in_637              ( col_in_637     ),
    .col_in_638              ( col_in_638     ),
    .col_in_639              ( col_in_639     ),
    .col_in_640              ( col_in_640     ),
    .col_in_641              ( col_in_641     ),
    .col_in_642              ( col_in_642     ),
    .col_in_643              ( col_in_643     ),
    .col_in_644              ( col_in_644     ),
    .col_in_645              ( col_in_645     ),
    .col_in_646              ( col_in_646     ),
    .col_in_647              ( col_in_647     ),
    .col_in_648              ( col_in_648     ),
    .col_in_649              ( col_in_649     ),
    .col_in_650              ( col_in_650     ),
    .col_in_651              ( col_in_651     ),
    .col_in_652              ( col_in_652     ),
    .col_in_653              ( col_in_653     ),
    .col_in_654              ( col_in_654     ),
    .col_in_655              ( col_in_655     ),
    .col_in_656              ( col_in_656     ),
    .col_in_657              ( col_in_657     ),
    .col_in_658              ( col_in_658     ),
    .col_in_659              ( col_in_659     ),
    .col_in_660              ( col_in_660     ),
    .col_in_661              ( col_in_661     ),
    .col_in_662              ( col_in_662     ),
    .col_in_663              ( col_in_663     ),
    .col_in_664              ( col_in_664     ),
    .col_in_665              ( col_in_665     ),
    .col_in_666              ( col_in_666     ),
    .col_in_667              ( col_in_667     ),
    .col_in_668              ( col_in_668     ),
    .col_in_669              ( col_in_669     ),
    .col_in_670              ( col_in_670     ),
    .col_in_671              ( col_in_671     ),
    .col_in_672              ( col_in_672     ),
    .col_in_673              ( col_in_673     ),
    .col_in_674              ( col_in_674     ),
    .col_in_675              ( col_in_675     ),
    .col_in_676              ( col_in_676     ),
    .col_in_677              ( col_in_677     ),
    .col_in_678              ( col_in_678     ),
    .col_in_679              ( col_in_679     ),
    .col_in_680              ( col_in_680     ),
    .col_in_681              ( col_in_681     ),
    .col_in_682              ( col_in_682     ),
    .col_in_683              ( col_in_683     ),
    .col_in_684              ( col_in_684     ),
    .col_in_685              ( col_in_685     ),
    .col_in_686              ( col_in_686     ),
    .col_in_687              ( col_in_687     ),
    .col_in_688              ( col_in_688     ),
    .col_in_689              ( col_in_689     ),
    .col_in_690              ( col_in_690     ),
    .col_in_691              ( col_in_691     ),
    .col_in_692              ( col_in_692     ),
    .col_in_693              ( col_in_693     ),
    .col_in_694              ( col_in_694     ),
    .col_in_695              ( col_in_695     ),
    .col_in_696              ( col_in_696     ),
    .col_in_697              ( col_in_697     ),
    .col_in_698              ( col_in_698     ),
    .col_in_699              ( col_in_699     ),
    .col_in_700              ( col_in_700     ),
    .col_in_701              ( col_in_701     ),
    .col_in_702              ( col_in_702     ),
    .col_in_703              ( col_in_703     ),
    .col_in_704              ( col_in_704     ),
    .col_in_705              ( col_in_705     ),
    .col_in_706              ( col_in_706     ),
    .col_in_707              ( col_in_707     ),
    .col_in_708              ( col_in_708     ),
    .col_in_709              ( col_in_709     ),
    .col_in_710              ( col_in_710     ),
    .col_in_711              ( col_in_711     ),
    .col_in_712              ( col_in_712     ),
    .col_in_713              ( col_in_713     ),
    .col_in_714              ( col_in_714     ),
    .col_in_715              ( col_in_715     ),
    .col_in_716              ( col_in_716     ),
    .col_in_717              ( col_in_717     ),
    .col_in_718              ( col_in_718     ),
    .col_in_719              ( col_in_719     ),
    .col_in_720              ( col_in_720     ),
    .col_in_721              ( col_in_721     ),
    .col_in_722              ( col_in_722     ),
    .col_in_723              ( col_in_723     ),
    .col_in_724              ( col_in_724     ),
    .col_in_725              ( col_in_725     ),
    .col_in_726              ( col_in_726     ),
    .col_in_727              ( col_in_727     ),
    .col_in_728              ( col_in_728     ),
    .col_in_729              ( col_in_729     ),
    .col_in_730              ( col_in_730     ),
    .col_in_731              ( col_in_731     ),
    .col_in_732              ( col_in_732     ),
    .col_in_733              ( col_in_733     ),
    .col_in_734              ( col_in_734     ),
    .col_in_735              ( col_in_735     ),
    .col_in_736              ( col_in_736     ),
    .col_in_737              ( col_in_737     ),
    .col_in_738              ( col_in_738     ),
    .col_in_739              ( col_in_739     ),
    .col_in_740              ( col_in_740     ),
    .col_in_741              ( col_in_741     ),
    .col_in_742              ( col_in_742     ),
    .col_in_743              ( col_in_743     ),
    .col_in_744              ( col_in_744     ),
    .col_in_745              ( col_in_745     ),
    .col_in_746              ( col_in_746     ),
    .col_in_747              ( col_in_747     ),
    .col_in_748              ( col_in_748     ),
    .col_in_749              ( col_in_749     ),
    .col_in_750              ( col_in_750     ),
    .col_in_751              ( col_in_751     ),
    .col_in_752              ( col_in_752     ),
    .col_in_753              ( col_in_753     ),
    .col_in_754              ( col_in_754     ),
    .col_in_755              ( col_in_755     ),
    .col_in_756              ( col_in_756     ),
    .col_in_757              ( col_in_757     ),
    .col_in_758              ( col_in_758     ),
    .col_in_759              ( col_in_759     ),
    .col_in_760              ( col_in_760     ),
    .col_in_761              ( col_in_761     ),
    .col_in_762              ( col_in_762     ),
    .col_in_763              ( col_in_763     ),
    .col_in_764              ( col_in_764     ),
    .col_in_765              ( col_in_765     ),
    .col_in_766              ( col_in_766     ),
    .col_in_767              ( col_in_767     ),
    .col_in_768              ( col_in_768     ),
    .col_in_769              ( col_in_769     ),
    .col_in_770              ( col_in_770     ),
    .col_in_771              ( col_in_771     ),
    .col_in_772              ( col_in_772     ),
    .col_in_773              ( col_in_773     ),
    .col_in_774              ( col_in_774     ),
    .col_in_775              ( col_in_775     ),
    .col_in_776              ( col_in_776     ),
    .col_in_777              ( col_in_777     ),
    .col_in_778              ( col_in_778     ),
    .col_in_779              ( col_in_779     ),
    .col_in_780              ( col_in_780     ),
    .col_in_781              ( col_in_781     ),
    .col_in_782              ( col_in_782     ),
    .col_in_783              ( col_in_783     ),
    .col_in_784              ( col_in_784     ),
    .col_in_785              ( col_in_785     ),
    .col_in_786              ( col_in_786     ),
    .col_in_787              ( col_in_787     ),
    .col_in_788              ( col_in_788     ),
    .col_in_789              ( col_in_789     ),
    .col_in_790              ( col_in_790     ),
    .col_in_791              ( col_in_791     ),
    .col_in_792              ( col_in_792     ),
    .col_in_793              ( col_in_793     ),
    .col_in_794              ( col_in_794     ),
    .col_in_795              ( col_in_795     ),
    .col_in_796              ( col_in_796     ),
    .col_in_797              ( col_in_797     ),
    .col_in_798              ( col_in_798     ),
    .col_in_799              ( col_in_799     ),
    .col_in_800              ( col_in_800     ),
    .col_in_801              ( col_in_801     ),
    .col_in_802              ( col_in_802     ),
    .col_in_803              ( col_in_803     ),
    .col_in_804              ( col_in_804     ),
    .col_in_805              ( col_in_805     ),
    .col_in_806              ( col_in_806     ),
    .col_in_807              ( col_in_807     ),
    .col_in_808              ( col_in_808     ),
    .col_in_809              ( col_in_809     ),
    .col_in_810              ( col_in_810     ),
    .col_in_811              ( col_in_811     ),
    .col_in_812              ( col_in_812     ),
    .col_in_813              ( col_in_813     ),
    .col_in_814              ( col_in_814     ),
    .col_in_815              ( col_in_815     ),
    .col_in_816              ( col_in_816     ),
    .col_in_817              ( col_in_817     ),
    .col_in_818              ( col_in_818     ),
    .col_in_819              ( col_in_819     ),
    .col_in_820              ( col_in_820     ),
    .col_in_821              ( col_in_821     ),
    .col_in_822              ( col_in_822     ),
    .col_in_823              ( col_in_823     ),
    .col_in_824              ( col_in_824     ),
    .col_in_825              ( col_in_825     ),
    .col_in_826              ( col_in_826     ),
    .col_in_827              ( col_in_827     ),
    .col_in_828              ( col_in_828     ),
    .col_in_829              ( col_in_829     ),
    .col_in_830              ( col_in_830     ),
    .col_in_831              ( col_in_831     ),
    .col_in_832              ( col_in_832     ),
    .col_in_833              ( col_in_833     ),
    .col_in_834              ( col_in_834     ),
    .col_in_835              ( col_in_835     ),
    .col_in_836              ( col_in_836     ),
    .col_in_837              ( col_in_837     ),
    .col_in_838              ( col_in_838     ),
    .col_in_839              ( col_in_839     ),
    .col_in_840              ( col_in_840     ),
    .col_in_841              ( col_in_841     ),
    .col_in_842              ( col_in_842     ),
    .col_in_843              ( col_in_843     ),
    .col_in_844              ( col_in_844     ),
    .col_in_845              ( col_in_845     ),
    .col_in_846              ( col_in_846     ),
    .col_in_847              ( col_in_847     ),
    .col_in_848              ( col_in_848     ),
    .col_in_849              ( col_in_849     ),
    .col_in_850              ( col_in_850     ),
    .col_in_851              ( col_in_851     ),
    .col_in_852              ( col_in_852     ),
    .col_in_853              ( col_in_853     ),
    .col_in_854              ( col_in_854     ),
    .col_in_855              ( col_in_855     ),
    .col_in_856              ( col_in_856     ),
    .col_in_857              ( col_in_857     ),
    .col_in_858              ( col_in_858     ),
    .col_in_859              ( col_in_859     ),
    .col_in_860              ( col_in_860     ),
    .col_in_861              ( col_in_861     ),
    .col_in_862              ( col_in_862     ),
    .col_in_863              ( col_in_863     ),
    .col_in_864              ( col_in_864     ),
    .col_in_865              ( col_in_865     ),
    .col_in_866              ( col_in_866     ),
    .col_in_867              ( col_in_867     ),
    .col_in_868              ( col_in_868     ),
    .col_in_869              ( col_in_869     ),
    .col_in_870              ( col_in_870     ),
    .col_in_871              ( col_in_871     ),
    .col_in_872              ( col_in_872     ),
    .col_in_873              ( col_in_873     ),
    .col_in_874              ( col_in_874     ),
    .col_in_875              ( col_in_875     ),
    .col_in_876              ( col_in_876     ),
    .col_in_877              ( col_in_877     ),
    .col_in_878              ( col_in_878     ),
    .col_in_879              ( col_in_879     ),
    .col_in_880              ( col_in_880     ),
    .col_in_881              ( col_in_881     ),
    .col_in_882              ( col_in_882     ),
    .col_in_883              ( col_in_883     ),
    .col_in_884              ( col_in_884     ),
    .col_in_885              ( col_in_885     ),
    .col_in_886              ( col_in_886     ),
    .col_in_887              ( col_in_887     ),
    .col_in_888              ( col_in_888     ),
    .col_in_889              ( col_in_889     ),
    .col_in_890              ( col_in_890     ),
    .col_in_891              ( col_in_891     ),
    .col_in_892              ( col_in_892     ),
    .col_in_893              ( col_in_893     ),
    .col_in_894              ( col_in_894     ),
    .col_in_895              ( col_in_895     ),
    .col_in_896              ( col_in_896     ),
    .col_in_897              ( col_in_897     ),
    .col_in_898              ( col_in_898     ),
    .col_in_899              ( col_in_899     ),
    .col_in_900              ( col_in_900     ),
    .col_in_901              ( col_in_901     ),
    .col_in_902              ( col_in_902     ),
    .col_in_903              ( col_in_903     ),
    .col_in_904              ( col_in_904     ),
    .col_in_905              ( col_in_905     ),
    .col_in_906              ( col_in_906     ),
    .col_in_907              ( col_in_907     ),
    .col_in_908              ( col_in_908     ),
    .col_in_909              ( col_in_909     ),
    .col_in_910              ( col_in_910     ),
    .col_in_911              ( col_in_911     ),
    .col_in_912              ( col_in_912     ),
    .col_in_913              ( col_in_913     ),
    .col_in_914              ( col_in_914     ),
    .col_in_915              ( col_in_915     ),
    .col_in_916              ( col_in_916     ),
    .col_in_917              ( col_in_917     ),
    .col_in_918              ( col_in_918     ),
    .col_in_919              ( col_in_919     ),
    .col_in_920              ( col_in_920     ),
    .col_in_921              ( col_in_921     ),
    .col_in_922              ( col_in_922     ),
    .col_in_923              ( col_in_923     ),
    .col_in_924              ( col_in_924     ),
    .col_in_925              ( col_in_925     ),
    .col_in_926              ( col_in_926     ),
    .col_in_927              ( col_in_927     ),
    .col_in_928              ( col_in_928     ),
    .col_in_929              ( col_in_929     ),
    .col_in_930              ( col_in_930     ),
    .col_in_931              ( col_in_931     ),
    .col_in_932              ( col_in_932     ),
    .col_in_933              ( col_in_933     ),
    .col_in_934              ( col_in_934     ),
    .col_in_935              ( col_in_935     ),
    .col_in_936              ( col_in_936     ),
    .col_in_937              ( col_in_937     ),
    .col_in_938              ( col_in_938     ),
    .col_in_939              ( col_in_939     ),
    .col_in_940              ( col_in_940     ),
    .col_in_941              ( col_in_941     ),
    .col_in_942              ( col_in_942     ),
    .col_in_943              ( col_in_943     ),
    .col_in_944              ( col_in_944     ),
    .col_in_945              ( col_in_945     ),
    .col_in_946              ( col_in_946     ),
    .col_in_947              ( col_in_947     ),
    .col_in_948              ( col_in_948     ),
    .col_in_949              ( col_in_949     ),
    .col_in_950              ( col_in_950     ),
    .col_in_951              ( col_in_951     ),
    .col_in_952              ( col_in_952     ),
    .col_in_953              ( col_in_953     ),
    .col_in_954              ( col_in_954     ),
    .col_in_955              ( col_in_955     ),
    .col_in_956              ( col_in_956     ),
    .col_in_957              ( col_in_957     ),
    .col_in_958              ( col_in_958     ),
    .col_in_959              ( col_in_959     ),
    .col_in_960              ( col_in_960     ),
    .col_in_961              ( col_in_961     ),
    .col_in_962              ( col_in_962     ),
    .col_in_963              ( col_in_963     ),
    .col_in_964              ( col_in_964     ),
    .col_in_965              ( col_in_965     ),
    .col_in_966              ( col_in_966     ),
    .col_in_967              ( col_in_967     ),
    .col_in_968              ( col_in_968     ),
    .col_in_969              ( col_in_969     ),
    .col_in_970              ( col_in_970     ),
    .col_in_971              ( col_in_971     ),
    .col_in_972              ( col_in_972     ),
    .col_in_973              ( col_in_973     ),
    .col_in_974              ( col_in_974     ),
    .col_in_975              ( col_in_975     ),
    .col_in_976              ( col_in_976     ),
    .col_in_977              ( col_in_977     ),
    .col_in_978              ( col_in_978     ),
    .col_in_979              ( col_in_979     ),
    .col_in_980              ( col_in_980     ),
    .col_in_981              ( col_in_981     ),
    .col_in_982              ( col_in_982     ),
    .col_in_983              ( col_in_983     ),
    .col_in_984              ( col_in_984     ),
    .col_in_985              ( col_in_985     ),
    .col_in_986              ( col_in_986     ),
    .col_in_987              ( col_in_987     ),
    .col_in_988              ( col_in_988     ),
    .col_in_989              ( col_in_989     ),
    .col_in_990              ( col_in_990     ),
    .col_in_991              ( col_in_991     ),
    .col_in_992              ( col_in_992     ),
    .col_in_993              ( col_in_993     ),
    .col_in_994              ( col_in_994     ),
    .col_in_995              ( col_in_995     ),
    .col_in_996              ( col_in_996     ),
    .col_in_997              ( col_in_997     ),
    .col_in_998              ( col_in_998     ),
    .col_in_999              ( col_in_999     ),
    .col_in_1000             ( col_in_1000    ),
    .col_in_1001             ( col_in_1001    ),
    .col_in_1002             ( col_in_1002    ),
    .col_in_1003             ( col_in_1003    ),
    .col_in_1004             ( col_in_1004    ),
    .col_in_1005             ( col_in_1005    ),
    .col_in_1006             ( col_in_1006    ),
    .col_in_1007             ( col_in_1007    ),
    .col_in_1008             ( col_in_1008    ),
    .col_in_1009             ( col_in_1009    ),
    .col_in_1010             ( col_in_1010    ),
    .col_in_1011             ( col_in_1011    ),
    .col_in_1012             ( col_in_1012    ),
    .col_in_1013             ( col_in_1013    ),
    .col_in_1014             ( col_in_1014    ),
    .col_in_1015             ( col_in_1015    ),
    .col_in_1016             ( col_in_1016    ),
    .col_in_1017             ( col_in_1017    ),
    .col_in_1018             ( col_in_1018    ),
    .col_in_1019             ( col_in_1019    ),
    .col_in_1020             ( col_in_1020    ),
    .col_in_1021             ( col_in_1021    ),
    .col_in_1022             ( col_in_1022    ),
    .col_in_1023             ( col_in_1023    ),

    .col_out_0               ( col_out_0      ),
    .col_out_1               ( col_out_1      ),
    .col_out_2               ( col_out_2      ),
    .col_out_3               ( col_out_3      ),
    .col_out_4               ( col_out_4      ),
    .col_out_5               ( col_out_5      ),
    .col_out_6               ( col_out_6      ),
    .col_out_7               ( col_out_7      ),
    .col_out_8               ( col_out_8      ),
    .col_out_9               ( col_out_9      ),
    .col_out_10              ( col_out_10     ),
    .col_out_11              ( col_out_11     ),
    .col_out_12              ( col_out_12     ),
    .col_out_13              ( col_out_13     ),
    .col_out_14              ( col_out_14     ),
    .col_out_15              ( col_out_15     ),
    .col_out_16              ( col_out_16     ),
    .col_out_17              ( col_out_17     ),
    .col_out_18              ( col_out_18     ),
    .col_out_19              ( col_out_19     ),
    .col_out_20              ( col_out_20     ),
    .col_out_21              ( col_out_21     ),
    .col_out_22              ( col_out_22     ),
    .col_out_23              ( col_out_23     ),
    .col_out_24              ( col_out_24     ),
    .col_out_25              ( col_out_25     ),
    .col_out_26              ( col_out_26     ),
    .col_out_27              ( col_out_27     ),
    .col_out_28              ( col_out_28     ),
    .col_out_29              ( col_out_29     ),
    .col_out_30              ( col_out_30     ),
    .col_out_31              ( col_out_31     ),
    .col_out_32              ( col_out_32     ),
    .col_out_33              ( col_out_33     ),
    .col_out_34              ( col_out_34     ),
    .col_out_35              ( col_out_35     ),
    .col_out_36              ( col_out_36     ),
    .col_out_37              ( col_out_37     ),
    .col_out_38              ( col_out_38     ),
    .col_out_39              ( col_out_39     ),
    .col_out_40              ( col_out_40     ),
    .col_out_41              ( col_out_41     ),
    .col_out_42              ( col_out_42     ),
    .col_out_43              ( col_out_43     ),
    .col_out_44              ( col_out_44     ),
    .col_out_45              ( col_out_45     ),
    .col_out_46              ( col_out_46     ),
    .col_out_47              ( col_out_47     ),
    .col_out_48              ( col_out_48     ),
    .col_out_49              ( col_out_49     ),
    .col_out_50              ( col_out_50     ),
    .col_out_51              ( col_out_51     ),
    .col_out_52              ( col_out_52     ),
    .col_out_53              ( col_out_53     ),
    .col_out_54              ( col_out_54     ),
    .col_out_55              ( col_out_55     ),
    .col_out_56              ( col_out_56     ),
    .col_out_57              ( col_out_57     ),
    .col_out_58              ( col_out_58     ),
    .col_out_59              ( col_out_59     ),
    .col_out_60              ( col_out_60     ),
    .col_out_61              ( col_out_61     ),
    .col_out_62              ( col_out_62     ),
    .col_out_63              ( col_out_63     ),
    .col_out_64              ( col_out_64     ),
    .col_out_65              ( col_out_65     ),
    .col_out_66              ( col_out_66     ),
    .col_out_67              ( col_out_67     ),
    .col_out_68              ( col_out_68     ),
    .col_out_69              ( col_out_69     ),
    .col_out_70              ( col_out_70     ),
    .col_out_71              ( col_out_71     ),
    .col_out_72              ( col_out_72     ),
    .col_out_73              ( col_out_73     ),
    .col_out_74              ( col_out_74     ),
    .col_out_75              ( col_out_75     ),
    .col_out_76              ( col_out_76     ),
    .col_out_77              ( col_out_77     ),
    .col_out_78              ( col_out_78     ),
    .col_out_79              ( col_out_79     ),
    .col_out_80              ( col_out_80     ),
    .col_out_81              ( col_out_81     ),
    .col_out_82              ( col_out_82     ),
    .col_out_83              ( col_out_83     ),
    .col_out_84              ( col_out_84     ),
    .col_out_85              ( col_out_85     ),
    .col_out_86              ( col_out_86     ),
    .col_out_87              ( col_out_87     ),
    .col_out_88              ( col_out_88     ),
    .col_out_89              ( col_out_89     ),
    .col_out_90              ( col_out_90     ),
    .col_out_91              ( col_out_91     ),
    .col_out_92              ( col_out_92     ),
    .col_out_93              ( col_out_93     ),
    .col_out_94              ( col_out_94     ),
    .col_out_95              ( col_out_95     ),
    .col_out_96              ( col_out_96     ),
    .col_out_97              ( col_out_97     ),
    .col_out_98              ( col_out_98     ),
    .col_out_99              ( col_out_99     ),
    .col_out_100             ( col_out_100    ),
    .col_out_101             ( col_out_101    ),
    .col_out_102             ( col_out_102    ),
    .col_out_103             ( col_out_103    ),
    .col_out_104             ( col_out_104    ),
    .col_out_105             ( col_out_105    ),
    .col_out_106             ( col_out_106    ),
    .col_out_107             ( col_out_107    ),
    .col_out_108             ( col_out_108    ),
    .col_out_109             ( col_out_109    ),
    .col_out_110             ( col_out_110    ),
    .col_out_111             ( col_out_111    ),
    .col_out_112             ( col_out_112    ),
    .col_out_113             ( col_out_113    ),
    .col_out_114             ( col_out_114    ),
    .col_out_115             ( col_out_115    ),
    .col_out_116             ( col_out_116    ),
    .col_out_117             ( col_out_117    ),
    .col_out_118             ( col_out_118    ),
    .col_out_119             ( col_out_119    ),
    .col_out_120             ( col_out_120    ),
    .col_out_121             ( col_out_121    ),
    .col_out_122             ( col_out_122    ),
    .col_out_123             ( col_out_123    ),
    .col_out_124             ( col_out_124    ),
    .col_out_125             ( col_out_125    ),
    .col_out_126             ( col_out_126    ),
    .col_out_127             ( col_out_127    ),
    .col_out_128             ( col_out_128    ),
    .col_out_129             ( col_out_129    ),
    .col_out_130             ( col_out_130    ),
    .col_out_131             ( col_out_131    ),
    .col_out_132             ( col_out_132    ),
    .col_out_133             ( col_out_133    ),
    .col_out_134             ( col_out_134    ),
    .col_out_135             ( col_out_135    ),
    .col_out_136             ( col_out_136    ),
    .col_out_137             ( col_out_137    ),
    .col_out_138             ( col_out_138    ),
    .col_out_139             ( col_out_139    ),
    .col_out_140             ( col_out_140    ),
    .col_out_141             ( col_out_141    ),
    .col_out_142             ( col_out_142    ),
    .col_out_143             ( col_out_143    ),
    .col_out_144             ( col_out_144    ),
    .col_out_145             ( col_out_145    ),
    .col_out_146             ( col_out_146    ),
    .col_out_147             ( col_out_147    ),
    .col_out_148             ( col_out_148    ),
    .col_out_149             ( col_out_149    ),
    .col_out_150             ( col_out_150    ),
    .col_out_151             ( col_out_151    ),
    .col_out_152             ( col_out_152    ),
    .col_out_153             ( col_out_153    ),
    .col_out_154             ( col_out_154    ),
    .col_out_155             ( col_out_155    ),
    .col_out_156             ( col_out_156    ),
    .col_out_157             ( col_out_157    ),
    .col_out_158             ( col_out_158    ),
    .col_out_159             ( col_out_159    ),
    .col_out_160             ( col_out_160    ),
    .col_out_161             ( col_out_161    ),
    .col_out_162             ( col_out_162    ),
    .col_out_163             ( col_out_163    ),
    .col_out_164             ( col_out_164    ),
    .col_out_165             ( col_out_165    ),
    .col_out_166             ( col_out_166    ),
    .col_out_167             ( col_out_167    ),
    .col_out_168             ( col_out_168    ),
    .col_out_169             ( col_out_169    ),
    .col_out_170             ( col_out_170    ),
    .col_out_171             ( col_out_171    ),
    .col_out_172             ( col_out_172    ),
    .col_out_173             ( col_out_173    ),
    .col_out_174             ( col_out_174    ),
    .col_out_175             ( col_out_175    ),
    .col_out_176             ( col_out_176    ),
    .col_out_177             ( col_out_177    ),
    .col_out_178             ( col_out_178    ),
    .col_out_179             ( col_out_179    ),
    .col_out_180             ( col_out_180    ),
    .col_out_181             ( col_out_181    ),
    .col_out_182             ( col_out_182    ),
    .col_out_183             ( col_out_183    ),
    .col_out_184             ( col_out_184    ),
    .col_out_185             ( col_out_185    ),
    .col_out_186             ( col_out_186    ),
    .col_out_187             ( col_out_187    ),
    .col_out_188             ( col_out_188    ),
    .col_out_189             ( col_out_189    ),
    .col_out_190             ( col_out_190    ),
    .col_out_191             ( col_out_191    ),
    .col_out_192             ( col_out_192    ),
    .col_out_193             ( col_out_193    ),
    .col_out_194             ( col_out_194    ),
    .col_out_195             ( col_out_195    ),
    .col_out_196             ( col_out_196    ),
    .col_out_197             ( col_out_197    ),
    .col_out_198             ( col_out_198    ),
    .col_out_199             ( col_out_199    ),
    .col_out_200             ( col_out_200    ),
    .col_out_201             ( col_out_201    ),
    .col_out_202             ( col_out_202    ),
    .col_out_203             ( col_out_203    ),
    .col_out_204             ( col_out_204    ),
    .col_out_205             ( col_out_205    ),
    .col_out_206             ( col_out_206    ),
    .col_out_207             ( col_out_207    ),
    .col_out_208             ( col_out_208    ),
    .col_out_209             ( col_out_209    ),
    .col_out_210             ( col_out_210    ),
    .col_out_211             ( col_out_211    ),
    .col_out_212             ( col_out_212    ),
    .col_out_213             ( col_out_213    ),
    .col_out_214             ( col_out_214    ),
    .col_out_215             ( col_out_215    ),
    .col_out_216             ( col_out_216    ),
    .col_out_217             ( col_out_217    ),
    .col_out_218             ( col_out_218    ),
    .col_out_219             ( col_out_219    ),
    .col_out_220             ( col_out_220    ),
    .col_out_221             ( col_out_221    ),
    .col_out_222             ( col_out_222    ),
    .col_out_223             ( col_out_223    ),
    .col_out_224             ( col_out_224    ),
    .col_out_225             ( col_out_225    ),
    .col_out_226             ( col_out_226    ),
    .col_out_227             ( col_out_227    ),
    .col_out_228             ( col_out_228    ),
    .col_out_229             ( col_out_229    ),
    .col_out_230             ( col_out_230    ),
    .col_out_231             ( col_out_231    ),
    .col_out_232             ( col_out_232    ),
    .col_out_233             ( col_out_233    ),
    .col_out_234             ( col_out_234    ),
    .col_out_235             ( col_out_235    ),
    .col_out_236             ( col_out_236    ),
    .col_out_237             ( col_out_237    ),
    .col_out_238             ( col_out_238    ),
    .col_out_239             ( col_out_239    ),
    .col_out_240             ( col_out_240    ),
    .col_out_241             ( col_out_241    ),
    .col_out_242             ( col_out_242    ),
    .col_out_243             ( col_out_243    ),
    .col_out_244             ( col_out_244    ),
    .col_out_245             ( col_out_245    ),
    .col_out_246             ( col_out_246    ),
    .col_out_247             ( col_out_247    ),
    .col_out_248             ( col_out_248    ),
    .col_out_249             ( col_out_249    ),
    .col_out_250             ( col_out_250    ),
    .col_out_251             ( col_out_251    ),
    .col_out_252             ( col_out_252    ),
    .col_out_253             ( col_out_253    ),
    .col_out_254             ( col_out_254    ),
    .col_out_255             ( col_out_255    ),
    .col_out_256             ( col_out_256    ),
    .col_out_257             ( col_out_257    ),
    .col_out_258             ( col_out_258    ),
    .col_out_259             ( col_out_259    ),
    .col_out_260             ( col_out_260    ),
    .col_out_261             ( col_out_261    ),
    .col_out_262             ( col_out_262    ),
    .col_out_263             ( col_out_263    ),
    .col_out_264             ( col_out_264    ),
    .col_out_265             ( col_out_265    ),
    .col_out_266             ( col_out_266    ),
    .col_out_267             ( col_out_267    ),
    .col_out_268             ( col_out_268    ),
    .col_out_269             ( col_out_269    ),
    .col_out_270             ( col_out_270    ),
    .col_out_271             ( col_out_271    ),
    .col_out_272             ( col_out_272    ),
    .col_out_273             ( col_out_273    ),
    .col_out_274             ( col_out_274    ),
    .col_out_275             ( col_out_275    ),
    .col_out_276             ( col_out_276    ),
    .col_out_277             ( col_out_277    ),
    .col_out_278             ( col_out_278    ),
    .col_out_279             ( col_out_279    ),
    .col_out_280             ( col_out_280    ),
    .col_out_281             ( col_out_281    ),
    .col_out_282             ( col_out_282    ),
    .col_out_283             ( col_out_283    ),
    .col_out_284             ( col_out_284    ),
    .col_out_285             ( col_out_285    ),
    .col_out_286             ( col_out_286    ),
    .col_out_287             ( col_out_287    ),
    .col_out_288             ( col_out_288    ),
    .col_out_289             ( col_out_289    ),
    .col_out_290             ( col_out_290    ),
    .col_out_291             ( col_out_291    ),
    .col_out_292             ( col_out_292    ),
    .col_out_293             ( col_out_293    ),
    .col_out_294             ( col_out_294    ),
    .col_out_295             ( col_out_295    ),
    .col_out_296             ( col_out_296    ),
    .col_out_297             ( col_out_297    ),
    .col_out_298             ( col_out_298    ),
    .col_out_299             ( col_out_299    ),
    .col_out_300             ( col_out_300    ),
    .col_out_301             ( col_out_301    ),
    .col_out_302             ( col_out_302    ),
    .col_out_303             ( col_out_303    ),
    .col_out_304             ( col_out_304    ),
    .col_out_305             ( col_out_305    ),
    .col_out_306             ( col_out_306    ),
    .col_out_307             ( col_out_307    ),
    .col_out_308             ( col_out_308    ),
    .col_out_309             ( col_out_309    ),
    .col_out_310             ( col_out_310    ),
    .col_out_311             ( col_out_311    ),
    .col_out_312             ( col_out_312    ),
    .col_out_313             ( col_out_313    ),
    .col_out_314             ( col_out_314    ),
    .col_out_315             ( col_out_315    ),
    .col_out_316             ( col_out_316    ),
    .col_out_317             ( col_out_317    ),
    .col_out_318             ( col_out_318    ),
    .col_out_319             ( col_out_319    ),
    .col_out_320             ( col_out_320    ),
    .col_out_321             ( col_out_321    ),
    .col_out_322             ( col_out_322    ),
    .col_out_323             ( col_out_323    ),
    .col_out_324             ( col_out_324    ),
    .col_out_325             ( col_out_325    ),
    .col_out_326             ( col_out_326    ),
    .col_out_327             ( col_out_327    ),
    .col_out_328             ( col_out_328    ),
    .col_out_329             ( col_out_329    ),
    .col_out_330             ( col_out_330    ),
    .col_out_331             ( col_out_331    ),
    .col_out_332             ( col_out_332    ),
    .col_out_333             ( col_out_333    ),
    .col_out_334             ( col_out_334    ),
    .col_out_335             ( col_out_335    ),
    .col_out_336             ( col_out_336    ),
    .col_out_337             ( col_out_337    ),
    .col_out_338             ( col_out_338    ),
    .col_out_339             ( col_out_339    ),
    .col_out_340             ( col_out_340    ),
    .col_out_341             ( col_out_341    ),
    .col_out_342             ( col_out_342    ),
    .col_out_343             ( col_out_343    ),
    .col_out_344             ( col_out_344    ),
    .col_out_345             ( col_out_345    ),
    .col_out_346             ( col_out_346    ),
    .col_out_347             ( col_out_347    ),
    .col_out_348             ( col_out_348    ),
    .col_out_349             ( col_out_349    ),
    .col_out_350             ( col_out_350    ),
    .col_out_351             ( col_out_351    ),
    .col_out_352             ( col_out_352    ),
    .col_out_353             ( col_out_353    ),
    .col_out_354             ( col_out_354    ),
    .col_out_355             ( col_out_355    ),
    .col_out_356             ( col_out_356    ),
    .col_out_357             ( col_out_357    ),
    .col_out_358             ( col_out_358    ),
    .col_out_359             ( col_out_359    ),
    .col_out_360             ( col_out_360    ),
    .col_out_361             ( col_out_361    ),
    .col_out_362             ( col_out_362    ),
    .col_out_363             ( col_out_363    ),
    .col_out_364             ( col_out_364    ),
    .col_out_365             ( col_out_365    ),
    .col_out_366             ( col_out_366    ),
    .col_out_367             ( col_out_367    ),
    .col_out_368             ( col_out_368    ),
    .col_out_369             ( col_out_369    ),
    .col_out_370             ( col_out_370    ),
    .col_out_371             ( col_out_371    ),
    .col_out_372             ( col_out_372    ),
    .col_out_373             ( col_out_373    ),
    .col_out_374             ( col_out_374    ),
    .col_out_375             ( col_out_375    ),
    .col_out_376             ( col_out_376    ),
    .col_out_377             ( col_out_377    ),
    .col_out_378             ( col_out_378    ),
    .col_out_379             ( col_out_379    ),
    .col_out_380             ( col_out_380    ),
    .col_out_381             ( col_out_381    ),
    .col_out_382             ( col_out_382    ),
    .col_out_383             ( col_out_383    ),
    .col_out_384             ( col_out_384    ),
    .col_out_385             ( col_out_385    ),
    .col_out_386             ( col_out_386    ),
    .col_out_387             ( col_out_387    ),
    .col_out_388             ( col_out_388    ),
    .col_out_389             ( col_out_389    ),
    .col_out_390             ( col_out_390    ),
    .col_out_391             ( col_out_391    ),
    .col_out_392             ( col_out_392    ),
    .col_out_393             ( col_out_393    ),
    .col_out_394             ( col_out_394    ),
    .col_out_395             ( col_out_395    ),
    .col_out_396             ( col_out_396    ),
    .col_out_397             ( col_out_397    ),
    .col_out_398             ( col_out_398    ),
    .col_out_399             ( col_out_399    ),
    .col_out_400             ( col_out_400    ),
    .col_out_401             ( col_out_401    ),
    .col_out_402             ( col_out_402    ),
    .col_out_403             ( col_out_403    ),
    .col_out_404             ( col_out_404    ),
    .col_out_405             ( col_out_405    ),
    .col_out_406             ( col_out_406    ),
    .col_out_407             ( col_out_407    ),
    .col_out_408             ( col_out_408    ),
    .col_out_409             ( col_out_409    ),
    .col_out_410             ( col_out_410    ),
    .col_out_411             ( col_out_411    ),
    .col_out_412             ( col_out_412    ),
    .col_out_413             ( col_out_413    ),
    .col_out_414             ( col_out_414    ),
    .col_out_415             ( col_out_415    ),
    .col_out_416             ( col_out_416    ),
    .col_out_417             ( col_out_417    ),
    .col_out_418             ( col_out_418    ),
    .col_out_419             ( col_out_419    ),
    .col_out_420             ( col_out_420    ),
    .col_out_421             ( col_out_421    ),
    .col_out_422             ( col_out_422    ),
    .col_out_423             ( col_out_423    ),
    .col_out_424             ( col_out_424    ),
    .col_out_425             ( col_out_425    ),
    .col_out_426             ( col_out_426    ),
    .col_out_427             ( col_out_427    ),
    .col_out_428             ( col_out_428    ),
    .col_out_429             ( col_out_429    ),
    .col_out_430             ( col_out_430    ),
    .col_out_431             ( col_out_431    ),
    .col_out_432             ( col_out_432    ),
    .col_out_433             ( col_out_433    ),
    .col_out_434             ( col_out_434    ),
    .col_out_435             ( col_out_435    ),
    .col_out_436             ( col_out_436    ),
    .col_out_437             ( col_out_437    ),
    .col_out_438             ( col_out_438    ),
    .col_out_439             ( col_out_439    ),
    .col_out_440             ( col_out_440    ),
    .col_out_441             ( col_out_441    ),
    .col_out_442             ( col_out_442    ),
    .col_out_443             ( col_out_443    ),
    .col_out_444             ( col_out_444    ),
    .col_out_445             ( col_out_445    ),
    .col_out_446             ( col_out_446    ),
    .col_out_447             ( col_out_447    ),
    .col_out_448             ( col_out_448    ),
    .col_out_449             ( col_out_449    ),
    .col_out_450             ( col_out_450    ),
    .col_out_451             ( col_out_451    ),
    .col_out_452             ( col_out_452    ),
    .col_out_453             ( col_out_453    ),
    .col_out_454             ( col_out_454    ),
    .col_out_455             ( col_out_455    ),
    .col_out_456             ( col_out_456    ),
    .col_out_457             ( col_out_457    ),
    .col_out_458             ( col_out_458    ),
    .col_out_459             ( col_out_459    ),
    .col_out_460             ( col_out_460    ),
    .col_out_461             ( col_out_461    ),
    .col_out_462             ( col_out_462    ),
    .col_out_463             ( col_out_463    ),
    .col_out_464             ( col_out_464    ),
    .col_out_465             ( col_out_465    ),
    .col_out_466             ( col_out_466    ),
    .col_out_467             ( col_out_467    ),
    .col_out_468             ( col_out_468    ),
    .col_out_469             ( col_out_469    ),
    .col_out_470             ( col_out_470    ),
    .col_out_471             ( col_out_471    ),
    .col_out_472             ( col_out_472    ),
    .col_out_473             ( col_out_473    ),
    .col_out_474             ( col_out_474    ),
    .col_out_475             ( col_out_475    ),
    .col_out_476             ( col_out_476    ),
    .col_out_477             ( col_out_477    ),
    .col_out_478             ( col_out_478    ),
    .col_out_479             ( col_out_479    ),
    .col_out_480             ( col_out_480    ),
    .col_out_481             ( col_out_481    ),
    .col_out_482             ( col_out_482    ),
    .col_out_483             ( col_out_483    ),
    .col_out_484             ( col_out_484    ),
    .col_out_485             ( col_out_485    ),
    .col_out_486             ( col_out_486    ),
    .col_out_487             ( col_out_487    ),
    .col_out_488             ( col_out_488    ),
    .col_out_489             ( col_out_489    ),
    .col_out_490             ( col_out_490    ),
    .col_out_491             ( col_out_491    ),
    .col_out_492             ( col_out_492    ),
    .col_out_493             ( col_out_493    ),
    .col_out_494             ( col_out_494    ),
    .col_out_495             ( col_out_495    ),
    .col_out_496             ( col_out_496    ),
    .col_out_497             ( col_out_497    ),
    .col_out_498             ( col_out_498    ),
    .col_out_499             ( col_out_499    ),
    .col_out_500             ( col_out_500    ),
    .col_out_501             ( col_out_501    ),
    .col_out_502             ( col_out_502    ),
    .col_out_503             ( col_out_503    ),
    .col_out_504             ( col_out_504    ),
    .col_out_505             ( col_out_505    ),
    .col_out_506             ( col_out_506    ),
    .col_out_507             ( col_out_507    ),
    .col_out_508             ( col_out_508    ),
    .col_out_509             ( col_out_509    ),
    .col_out_510             ( col_out_510    ),
    .col_out_511             ( col_out_511    ),
    .col_out_512             ( col_out_512    ),
    .col_out_513             ( col_out_513    ),
    .col_out_514             ( col_out_514    ),
    .col_out_515             ( col_out_515    ),
    .col_out_516             ( col_out_516    ),
    .col_out_517             ( col_out_517    ),
    .col_out_518             ( col_out_518    ),
    .col_out_519             ( col_out_519    ),
    .col_out_520             ( col_out_520    ),
    .col_out_521             ( col_out_521    ),
    .col_out_522             ( col_out_522    ),
    .col_out_523             ( col_out_523    ),
    .col_out_524             ( col_out_524    ),
    .col_out_525             ( col_out_525    ),
    .col_out_526             ( col_out_526    ),
    .col_out_527             ( col_out_527    ),
    .col_out_528             ( col_out_528    ),
    .col_out_529             ( col_out_529    ),
    .col_out_530             ( col_out_530    ),
    .col_out_531             ( col_out_531    ),
    .col_out_532             ( col_out_532    ),
    .col_out_533             ( col_out_533    ),
    .col_out_534             ( col_out_534    ),
    .col_out_535             ( col_out_535    ),
    .col_out_536             ( col_out_536    ),
    .col_out_537             ( col_out_537    ),
    .col_out_538             ( col_out_538    ),
    .col_out_539             ( col_out_539    ),
    .col_out_540             ( col_out_540    ),
    .col_out_541             ( col_out_541    ),
    .col_out_542             ( col_out_542    ),
    .col_out_543             ( col_out_543    ),
    .col_out_544             ( col_out_544    ),
    .col_out_545             ( col_out_545    ),
    .col_out_546             ( col_out_546    ),
    .col_out_547             ( col_out_547    ),
    .col_out_548             ( col_out_548    ),
    .col_out_549             ( col_out_549    ),
    .col_out_550             ( col_out_550    ),
    .col_out_551             ( col_out_551    ),
    .col_out_552             ( col_out_552    ),
    .col_out_553             ( col_out_553    ),
    .col_out_554             ( col_out_554    ),
    .col_out_555             ( col_out_555    ),
    .col_out_556             ( col_out_556    ),
    .col_out_557             ( col_out_557    ),
    .col_out_558             ( col_out_558    ),
    .col_out_559             ( col_out_559    ),
    .col_out_560             ( col_out_560    ),
    .col_out_561             ( col_out_561    ),
    .col_out_562             ( col_out_562    ),
    .col_out_563             ( col_out_563    ),
    .col_out_564             ( col_out_564    ),
    .col_out_565             ( col_out_565    ),
    .col_out_566             ( col_out_566    ),
    .col_out_567             ( col_out_567    ),
    .col_out_568             ( col_out_568    ),
    .col_out_569             ( col_out_569    ),
    .col_out_570             ( col_out_570    ),
    .col_out_571             ( col_out_571    ),
    .col_out_572             ( col_out_572    ),
    .col_out_573             ( col_out_573    ),
    .col_out_574             ( col_out_574    ),
    .col_out_575             ( col_out_575    ),
    .col_out_576             ( col_out_576    ),
    .col_out_577             ( col_out_577    ),
    .col_out_578             ( col_out_578    ),
    .col_out_579             ( col_out_579    ),
    .col_out_580             ( col_out_580    ),
    .col_out_581             ( col_out_581    ),
    .col_out_582             ( col_out_582    ),
    .col_out_583             ( col_out_583    ),
    .col_out_584             ( col_out_584    ),
    .col_out_585             ( col_out_585    ),
    .col_out_586             ( col_out_586    ),
    .col_out_587             ( col_out_587    ),
    .col_out_588             ( col_out_588    ),
    .col_out_589             ( col_out_589    ),
    .col_out_590             ( col_out_590    ),
    .col_out_591             ( col_out_591    ),
    .col_out_592             ( col_out_592    ),
    .col_out_593             ( col_out_593    ),
    .col_out_594             ( col_out_594    ),
    .col_out_595             ( col_out_595    ),
    .col_out_596             ( col_out_596    ),
    .col_out_597             ( col_out_597    ),
    .col_out_598             ( col_out_598    ),
    .col_out_599             ( col_out_599    ),
    .col_out_600             ( col_out_600    ),
    .col_out_601             ( col_out_601    ),
    .col_out_602             ( col_out_602    ),
    .col_out_603             ( col_out_603    ),
    .col_out_604             ( col_out_604    ),
    .col_out_605             ( col_out_605    ),
    .col_out_606             ( col_out_606    ),
    .col_out_607             ( col_out_607    ),
    .col_out_608             ( col_out_608    ),
    .col_out_609             ( col_out_609    ),
    .col_out_610             ( col_out_610    ),
    .col_out_611             ( col_out_611    ),
    .col_out_612             ( col_out_612    ),
    .col_out_613             ( col_out_613    ),
    .col_out_614             ( col_out_614    ),
    .col_out_615             ( col_out_615    ),
    .col_out_616             ( col_out_616    ),
    .col_out_617             ( col_out_617    ),
    .col_out_618             ( col_out_618    ),
    .col_out_619             ( col_out_619    ),
    .col_out_620             ( col_out_620    ),
    .col_out_621             ( col_out_621    ),
    .col_out_622             ( col_out_622    ),
    .col_out_623             ( col_out_623    ),
    .col_out_624             ( col_out_624    ),
    .col_out_625             ( col_out_625    ),
    .col_out_626             ( col_out_626    ),
    .col_out_627             ( col_out_627    ),
    .col_out_628             ( col_out_628    ),
    .col_out_629             ( col_out_629    ),
    .col_out_630             ( col_out_630    ),
    .col_out_631             ( col_out_631    ),
    .col_out_632             ( col_out_632    ),
    .col_out_633             ( col_out_633    ),
    .col_out_634             ( col_out_634    ),
    .col_out_635             ( col_out_635    ),
    .col_out_636             ( col_out_636    ),
    .col_out_637             ( col_out_637    ),
    .col_out_638             ( col_out_638    ),
    .col_out_639             ( col_out_639    ),
    .col_out_640             ( col_out_640    ),
    .col_out_641             ( col_out_641    ),
    .col_out_642             ( col_out_642    ),
    .col_out_643             ( col_out_643    ),
    .col_out_644             ( col_out_644    ),
    .col_out_645             ( col_out_645    ),
    .col_out_646             ( col_out_646    ),
    .col_out_647             ( col_out_647    ),
    .col_out_648             ( col_out_648    ),
    .col_out_649             ( col_out_649    ),
    .col_out_650             ( col_out_650    ),
    .col_out_651             ( col_out_651    ),
    .col_out_652             ( col_out_652    ),
    .col_out_653             ( col_out_653    ),
    .col_out_654             ( col_out_654    ),
    .col_out_655             ( col_out_655    ),
    .col_out_656             ( col_out_656    ),
    .col_out_657             ( col_out_657    ),
    .col_out_658             ( col_out_658    ),
    .col_out_659             ( col_out_659    ),
    .col_out_660             ( col_out_660    ),
    .col_out_661             ( col_out_661    ),
    .col_out_662             ( col_out_662    ),
    .col_out_663             ( col_out_663    ),
    .col_out_664             ( col_out_664    ),
    .col_out_665             ( col_out_665    ),
    .col_out_666             ( col_out_666    ),
    .col_out_667             ( col_out_667    ),
    .col_out_668             ( col_out_668    ),
    .col_out_669             ( col_out_669    ),
    .col_out_670             ( col_out_670    ),
    .col_out_671             ( col_out_671    ),
    .col_out_672             ( col_out_672    ),
    .col_out_673             ( col_out_673    ),
    .col_out_674             ( col_out_674    ),
    .col_out_675             ( col_out_675    ),
    .col_out_676             ( col_out_676    ),
    .col_out_677             ( col_out_677    ),
    .col_out_678             ( col_out_678    ),
    .col_out_679             ( col_out_679    ),
    .col_out_680             ( col_out_680    ),
    .col_out_681             ( col_out_681    ),
    .col_out_682             ( col_out_682    ),
    .col_out_683             ( col_out_683    ),
    .col_out_684             ( col_out_684    ),
    .col_out_685             ( col_out_685    ),
    .col_out_686             ( col_out_686    ),
    .col_out_687             ( col_out_687    ),
    .col_out_688             ( col_out_688    ),
    .col_out_689             ( col_out_689    ),
    .col_out_690             ( col_out_690    ),
    .col_out_691             ( col_out_691    ),
    .col_out_692             ( col_out_692    ),
    .col_out_693             ( col_out_693    ),
    .col_out_694             ( col_out_694    ),
    .col_out_695             ( col_out_695    ),
    .col_out_696             ( col_out_696    ),
    .col_out_697             ( col_out_697    ),
    .col_out_698             ( col_out_698    ),
    .col_out_699             ( col_out_699    ),
    .col_out_700             ( col_out_700    ),
    .col_out_701             ( col_out_701    ),
    .col_out_702             ( col_out_702    ),
    .col_out_703             ( col_out_703    ),
    .col_out_704             ( col_out_704    ),
    .col_out_705             ( col_out_705    ),
    .col_out_706             ( col_out_706    ),
    .col_out_707             ( col_out_707    ),
    .col_out_708             ( col_out_708    ),
    .col_out_709             ( col_out_709    ),
    .col_out_710             ( col_out_710    ),
    .col_out_711             ( col_out_711    ),
    .col_out_712             ( col_out_712    ),
    .col_out_713             ( col_out_713    ),
    .col_out_714             ( col_out_714    ),
    .col_out_715             ( col_out_715    ),
    .col_out_716             ( col_out_716    ),
    .col_out_717             ( col_out_717    ),
    .col_out_718             ( col_out_718    ),
    .col_out_719             ( col_out_719    ),
    .col_out_720             ( col_out_720    ),
    .col_out_721             ( col_out_721    ),
    .col_out_722             ( col_out_722    ),
    .col_out_723             ( col_out_723    ),
    .col_out_724             ( col_out_724    ),
    .col_out_725             ( col_out_725    ),
    .col_out_726             ( col_out_726    ),
    .col_out_727             ( col_out_727    ),
    .col_out_728             ( col_out_728    ),
    .col_out_729             ( col_out_729    ),
    .col_out_730             ( col_out_730    ),
    .col_out_731             ( col_out_731    ),
    .col_out_732             ( col_out_732    ),
    .col_out_733             ( col_out_733    ),
    .col_out_734             ( col_out_734    ),
    .col_out_735             ( col_out_735    ),
    .col_out_736             ( col_out_736    ),
    .col_out_737             ( col_out_737    ),
    .col_out_738             ( col_out_738    ),
    .col_out_739             ( col_out_739    ),
    .col_out_740             ( col_out_740    ),
    .col_out_741             ( col_out_741    ),
    .col_out_742             ( col_out_742    ),
    .col_out_743             ( col_out_743    ),
    .col_out_744             ( col_out_744    ),
    .col_out_745             ( col_out_745    ),
    .col_out_746             ( col_out_746    ),
    .col_out_747             ( col_out_747    ),
    .col_out_748             ( col_out_748    ),
    .col_out_749             ( col_out_749    ),
    .col_out_750             ( col_out_750    ),
    .col_out_751             ( col_out_751    ),
    .col_out_752             ( col_out_752    ),
    .col_out_753             ( col_out_753    ),
    .col_out_754             ( col_out_754    ),
    .col_out_755             ( col_out_755    ),
    .col_out_756             ( col_out_756    ),
    .col_out_757             ( col_out_757    ),
    .col_out_758             ( col_out_758    ),
    .col_out_759             ( col_out_759    ),
    .col_out_760             ( col_out_760    ),
    .col_out_761             ( col_out_761    ),
    .col_out_762             ( col_out_762    ),
    .col_out_763             ( col_out_763    ),
    .col_out_764             ( col_out_764    ),
    .col_out_765             ( col_out_765    ),
    .col_out_766             ( col_out_766    ),
    .col_out_767             ( col_out_767    ),
    .col_out_768             ( col_out_768    ),
    .col_out_769             ( col_out_769    ),
    .col_out_770             ( col_out_770    ),
    .col_out_771             ( col_out_771    ),
    .col_out_772             ( col_out_772    ),
    .col_out_773             ( col_out_773    ),
    .col_out_774             ( col_out_774    ),
    .col_out_775             ( col_out_775    ),
    .col_out_776             ( col_out_776    ),
    .col_out_777             ( col_out_777    ),
    .col_out_778             ( col_out_778    ),
    .col_out_779             ( col_out_779    ),
    .col_out_780             ( col_out_780    ),
    .col_out_781             ( col_out_781    ),
    .col_out_782             ( col_out_782    ),
    .col_out_783             ( col_out_783    ),
    .col_out_784             ( col_out_784    ),
    .col_out_785             ( col_out_785    ),
    .col_out_786             ( col_out_786    ),
    .col_out_787             ( col_out_787    ),
    .col_out_788             ( col_out_788    ),
    .col_out_789             ( col_out_789    ),
    .col_out_790             ( col_out_790    ),
    .col_out_791             ( col_out_791    ),
    .col_out_792             ( col_out_792    ),
    .col_out_793             ( col_out_793    ),
    .col_out_794             ( col_out_794    ),
    .col_out_795             ( col_out_795    ),
    .col_out_796             ( col_out_796    ),
    .col_out_797             ( col_out_797    ),
    .col_out_798             ( col_out_798    ),
    .col_out_799             ( col_out_799    ),
    .col_out_800             ( col_out_800    ),
    .col_out_801             ( col_out_801    ),
    .col_out_802             ( col_out_802    ),
    .col_out_803             ( col_out_803    ),
    .col_out_804             ( col_out_804    ),
    .col_out_805             ( col_out_805    ),
    .col_out_806             ( col_out_806    ),
    .col_out_807             ( col_out_807    ),
    .col_out_808             ( col_out_808    ),
    .col_out_809             ( col_out_809    ),
    .col_out_810             ( col_out_810    ),
    .col_out_811             ( col_out_811    ),
    .col_out_812             ( col_out_812    ),
    .col_out_813             ( col_out_813    ),
    .col_out_814             ( col_out_814    ),
    .col_out_815             ( col_out_815    ),
    .col_out_816             ( col_out_816    ),
    .col_out_817             ( col_out_817    ),
    .col_out_818             ( col_out_818    ),
    .col_out_819             ( col_out_819    ),
    .col_out_820             ( col_out_820    ),
    .col_out_821             ( col_out_821    ),
    .col_out_822             ( col_out_822    ),
    .col_out_823             ( col_out_823    ),
    .col_out_824             ( col_out_824    ),
    .col_out_825             ( col_out_825    ),
    .col_out_826             ( col_out_826    ),
    .col_out_827             ( col_out_827    ),
    .col_out_828             ( col_out_828    ),
    .col_out_829             ( col_out_829    ),
    .col_out_830             ( col_out_830    ),
    .col_out_831             ( col_out_831    ),
    .col_out_832             ( col_out_832    ),
    .col_out_833             ( col_out_833    ),
    .col_out_834             ( col_out_834    ),
    .col_out_835             ( col_out_835    ),
    .col_out_836             ( col_out_836    ),
    .col_out_837             ( col_out_837    ),
    .col_out_838             ( col_out_838    ),
    .col_out_839             ( col_out_839    ),
    .col_out_840             ( col_out_840    ),
    .col_out_841             ( col_out_841    ),
    .col_out_842             ( col_out_842    ),
    .col_out_843             ( col_out_843    ),
    .col_out_844             ( col_out_844    ),
    .col_out_845             ( col_out_845    ),
    .col_out_846             ( col_out_846    ),
    .col_out_847             ( col_out_847    ),
    .col_out_848             ( col_out_848    ),
    .col_out_849             ( col_out_849    ),
    .col_out_850             ( col_out_850    ),
    .col_out_851             ( col_out_851    ),
    .col_out_852             ( col_out_852    ),
    .col_out_853             ( col_out_853    ),
    .col_out_854             ( col_out_854    ),
    .col_out_855             ( col_out_855    ),
    .col_out_856             ( col_out_856    ),
    .col_out_857             ( col_out_857    ),
    .col_out_858             ( col_out_858    ),
    .col_out_859             ( col_out_859    ),
    .col_out_860             ( col_out_860    ),
    .col_out_861             ( col_out_861    ),
    .col_out_862             ( col_out_862    ),
    .col_out_863             ( col_out_863    ),
    .col_out_864             ( col_out_864    ),
    .col_out_865             ( col_out_865    ),
    .col_out_866             ( col_out_866    ),
    .col_out_867             ( col_out_867    ),
    .col_out_868             ( col_out_868    ),
    .col_out_869             ( col_out_869    ),
    .col_out_870             ( col_out_870    ),
    .col_out_871             ( col_out_871    ),
    .col_out_872             ( col_out_872    ),
    .col_out_873             ( col_out_873    ),
    .col_out_874             ( col_out_874    ),
    .col_out_875             ( col_out_875    ),
    .col_out_876             ( col_out_876    ),
    .col_out_877             ( col_out_877    ),
    .col_out_878             ( col_out_878    ),
    .col_out_879             ( col_out_879    ),
    .col_out_880             ( col_out_880    ),
    .col_out_881             ( col_out_881    ),
    .col_out_882             ( col_out_882    ),
    .col_out_883             ( col_out_883    ),
    .col_out_884             ( col_out_884    ),
    .col_out_885             ( col_out_885    ),
    .col_out_886             ( col_out_886    ),
    .col_out_887             ( col_out_887    ),
    .col_out_888             ( col_out_888    ),
    .col_out_889             ( col_out_889    ),
    .col_out_890             ( col_out_890    ),
    .col_out_891             ( col_out_891    ),
    .col_out_892             ( col_out_892    ),
    .col_out_893             ( col_out_893    ),
    .col_out_894             ( col_out_894    ),
    .col_out_895             ( col_out_895    ),
    .col_out_896             ( col_out_896    ),
    .col_out_897             ( col_out_897    ),
    .col_out_898             ( col_out_898    ),
    .col_out_899             ( col_out_899    ),
    .col_out_900             ( col_out_900    ),
    .col_out_901             ( col_out_901    ),
    .col_out_902             ( col_out_902    ),
    .col_out_903             ( col_out_903    ),
    .col_out_904             ( col_out_904    ),
    .col_out_905             ( col_out_905    ),
    .col_out_906             ( col_out_906    ),
    .col_out_907             ( col_out_907    ),
    .col_out_908             ( col_out_908    ),
    .col_out_909             ( col_out_909    ),
    .col_out_910             ( col_out_910    ),
    .col_out_911             ( col_out_911    ),
    .col_out_912             ( col_out_912    ),
    .col_out_913             ( col_out_913    ),
    .col_out_914             ( col_out_914    ),
    .col_out_915             ( col_out_915    ),
    .col_out_916             ( col_out_916    ),
    .col_out_917             ( col_out_917    ),
    .col_out_918             ( col_out_918    ),
    .col_out_919             ( col_out_919    ),
    .col_out_920             ( col_out_920    ),
    .col_out_921             ( col_out_921    ),
    .col_out_922             ( col_out_922    ),
    .col_out_923             ( col_out_923    ),
    .col_out_924             ( col_out_924    ),
    .col_out_925             ( col_out_925    ),
    .col_out_926             ( col_out_926    ),
    .col_out_927             ( col_out_927    ),
    .col_out_928             ( col_out_928    ),
    .col_out_929             ( col_out_929    ),
    .col_out_930             ( col_out_930    ),
    .col_out_931             ( col_out_931    ),
    .col_out_932             ( col_out_932    ),
    .col_out_933             ( col_out_933    ),
    .col_out_934             ( col_out_934    ),
    .col_out_935             ( col_out_935    ),
    .col_out_936             ( col_out_936    ),
    .col_out_937             ( col_out_937    ),
    .col_out_938             ( col_out_938    ),
    .col_out_939             ( col_out_939    ),
    .col_out_940             ( col_out_940    ),
    .col_out_941             ( col_out_941    ),
    .col_out_942             ( col_out_942    ),
    .col_out_943             ( col_out_943    ),
    .col_out_944             ( col_out_944    ),
    .col_out_945             ( col_out_945    ),
    .col_out_946             ( col_out_946    ),
    .col_out_947             ( col_out_947    ),
    .col_out_948             ( col_out_948    ),
    .col_out_949             ( col_out_949    ),
    .col_out_950             ( col_out_950    ),
    .col_out_951             ( col_out_951    ),
    .col_out_952             ( col_out_952    ),
    .col_out_953             ( col_out_953    ),
    .col_out_954             ( col_out_954    ),
    .col_out_955             ( col_out_955    ),
    .col_out_956             ( col_out_956    ),
    .col_out_957             ( col_out_957    ),
    .col_out_958             ( col_out_958    ),
    .col_out_959             ( col_out_959    ),
    .col_out_960             ( col_out_960    ),
    .col_out_961             ( col_out_961    ),
    .col_out_962             ( col_out_962    ),
    .col_out_963             ( col_out_963    ),
    .col_out_964             ( col_out_964    ),
    .col_out_965             ( col_out_965    ),
    .col_out_966             ( col_out_966    ),
    .col_out_967             ( col_out_967    ),
    .col_out_968             ( col_out_968    ),
    .col_out_969             ( col_out_969    ),
    .col_out_970             ( col_out_970    ),
    .col_out_971             ( col_out_971    ),
    .col_out_972             ( col_out_972    ),
    .col_out_973             ( col_out_973    ),
    .col_out_974             ( col_out_974    ),
    .col_out_975             ( col_out_975    ),
    .col_out_976             ( col_out_976    ),
    .col_out_977             ( col_out_977    ),
    .col_out_978             ( col_out_978    ),
    .col_out_979             ( col_out_979    ),
    .col_out_980             ( col_out_980    ),
    .col_out_981             ( col_out_981    ),
    .col_out_982             ( col_out_982    ),
    .col_out_983             ( col_out_983    ),
    .col_out_984             ( col_out_984    ),
    .col_out_985             ( col_out_985    ),
    .col_out_986             ( col_out_986    ),
    .col_out_987             ( col_out_987    ),
    .col_out_988             ( col_out_988    ),
    .col_out_989             ( col_out_989    ),
    .col_out_990             ( col_out_990    ),
    .col_out_991             ( col_out_991    ),
    .col_out_992             ( col_out_992    ),
    .col_out_993             ( col_out_993    ),
    .col_out_994             ( col_out_994    ),
    .col_out_995             ( col_out_995    ),
    .col_out_996             ( col_out_996    ),
    .col_out_997             ( col_out_997    ),
    .col_out_998             ( col_out_998    ),
    .col_out_999             ( col_out_999    ),
    .col_out_1000            ( col_out_1000   ),
    .col_out_1001            ( col_out_1001   ),
    .col_out_1002            ( col_out_1002   ),
    .col_out_1003            ( col_out_1003   ),
    .col_out_1004            ( col_out_1004   ),
    .col_out_1005            ( col_out_1005   ),
    .col_out_1006            ( col_out_1006   ),
    .col_out_1007            ( col_out_1007   ),
    .col_out_1008            ( col_out_1008   ),
    .col_out_1009            ( col_out_1009   ),
    .col_out_1010            ( col_out_1010   ),
    .col_out_1011            ( col_out_1011   ),
    .col_out_1012            ( col_out_1012   ),
    .col_out_1013            ( col_out_1013   ),
    .col_out_1014            ( col_out_1014   ),
    .col_out_1015            ( col_out_1015   ),
    .col_out_1016            ( col_out_1016   ),
    .col_out_1017            ( col_out_1017   ),
    .col_out_1018            ( col_out_1018   ),
    .col_out_1019            ( col_out_1019   ),
    .col_out_1020            ( col_out_1020   ),
    .col_out_1021            ( col_out_1021   ),
    .col_out_1022            ( col_out_1022   ),
    .col_out_1023            ( col_out_1023   ),
    .col_out_1024            ( col_out_1024   )
);




//*****************************************************
//**************输出赋值******************************
//*****************************************************
assign row_out_0 = {col_out_1024[0], col_out_1023[0], col_out_1022[0], col_out_1021[0], col_out_1020[0], col_out_1019[0], col_out_1018[0], col_out_1017[0], col_out_1016[0], col_out_1015[0], col_out_1014[0], col_out_1013[0], col_out_1012[0], col_out_1011[0], col_out_1010[0], col_out_1009[0], col_out_1008[0], col_out_1007[0], col_out_1006[0], col_out_1005[0], col_out_1004[0], col_out_1003[0], col_out_1002[0], col_out_1001[0], col_out_1000[0], col_out_999[0], col_out_998[0], col_out_997[0], col_out_996[0], col_out_995[0], col_out_994[0], col_out_993[0], col_out_992[0], col_out_991[0], col_out_990[0], col_out_989[0], col_out_988[0], col_out_987[0], col_out_986[0], col_out_985[0], col_out_984[0], col_out_983[0], col_out_982[0], col_out_981[0], col_out_980[0], col_out_979[0], col_out_978[0], col_out_977[0], col_out_976[0], col_out_975[0], col_out_974[0], col_out_973[0], col_out_972[0], col_out_971[0], col_out_970[0], col_out_969[0], col_out_968[0], col_out_967[0], col_out_966[0], col_out_965[0], col_out_964[0], col_out_963[0], col_out_962[0], col_out_961[0], col_out_960[0], col_out_959[0], col_out_958[0], col_out_957[0], col_out_956[0], col_out_955[0], col_out_954[0], col_out_953[0], col_out_952[0], col_out_951[0], col_out_950[0], col_out_949[0], col_out_948[0], col_out_947[0], col_out_946[0], col_out_945[0], col_out_944[0], col_out_943[0], col_out_942[0], col_out_941[0], col_out_940[0], col_out_939[0], col_out_938[0], col_out_937[0], col_out_936[0], col_out_935[0], col_out_934[0], col_out_933[0], col_out_932[0], col_out_931[0], col_out_930[0], col_out_929[0], col_out_928[0], col_out_927[0], col_out_926[0], col_out_925[0], col_out_924[0], col_out_923[0], col_out_922[0], col_out_921[0], col_out_920[0], col_out_919[0], col_out_918[0], col_out_917[0], col_out_916[0], col_out_915[0], col_out_914[0], col_out_913[0], col_out_912[0], col_out_911[0], col_out_910[0], col_out_909[0], col_out_908[0], col_out_907[0], col_out_906[0], col_out_905[0], col_out_904[0], col_out_903[0], col_out_902[0], col_out_901[0], col_out_900[0], col_out_899[0], col_out_898[0], col_out_897[0], col_out_896[0], col_out_895[0], col_out_894[0], col_out_893[0], col_out_892[0], col_out_891[0], col_out_890[0], col_out_889[0], col_out_888[0], col_out_887[0], col_out_886[0], col_out_885[0], col_out_884[0], col_out_883[0], col_out_882[0], col_out_881[0], col_out_880[0], col_out_879[0], col_out_878[0], col_out_877[0], col_out_876[0], col_out_875[0], col_out_874[0], col_out_873[0], col_out_872[0], col_out_871[0], col_out_870[0], col_out_869[0], col_out_868[0], col_out_867[0], col_out_866[0], col_out_865[0], col_out_864[0], col_out_863[0], col_out_862[0], col_out_861[0], col_out_860[0], col_out_859[0], col_out_858[0], col_out_857[0], col_out_856[0], col_out_855[0], col_out_854[0], col_out_853[0], col_out_852[0], col_out_851[0], col_out_850[0], col_out_849[0], col_out_848[0], col_out_847[0], col_out_846[0], col_out_845[0], col_out_844[0], col_out_843[0], col_out_842[0], col_out_841[0], col_out_840[0], col_out_839[0], col_out_838[0], col_out_837[0], col_out_836[0], col_out_835[0], col_out_834[0], col_out_833[0], col_out_832[0], col_out_831[0], col_out_830[0], col_out_829[0], col_out_828[0], col_out_827[0], col_out_826[0], col_out_825[0], col_out_824[0], col_out_823[0], col_out_822[0], col_out_821[0], col_out_820[0], col_out_819[0], col_out_818[0], col_out_817[0], col_out_816[0], col_out_815[0], col_out_814[0], col_out_813[0], col_out_812[0], col_out_811[0], col_out_810[0], col_out_809[0], col_out_808[0], col_out_807[0], col_out_806[0], col_out_805[0], col_out_804[0], col_out_803[0], col_out_802[0], col_out_801[0], col_out_800[0], col_out_799[0], col_out_798[0], col_out_797[0], col_out_796[0], col_out_795[0], col_out_794[0], col_out_793[0], col_out_792[0], col_out_791[0], col_out_790[0], col_out_789[0], col_out_788[0], col_out_787[0], col_out_786[0], col_out_785[0], col_out_784[0], col_out_783[0], col_out_782[0], col_out_781[0], col_out_780[0], col_out_779[0], col_out_778[0], col_out_777[0], col_out_776[0], col_out_775[0], col_out_774[0], col_out_773[0], col_out_772[0], col_out_771[0], col_out_770[0], col_out_769[0], col_out_768[0], col_out_767[0], col_out_766[0], col_out_765[0], col_out_764[0], col_out_763[0], col_out_762[0], col_out_761[0], col_out_760[0], col_out_759[0], col_out_758[0], col_out_757[0], col_out_756[0], col_out_755[0], col_out_754[0], col_out_753[0], col_out_752[0], col_out_751[0], col_out_750[0], col_out_749[0], col_out_748[0], col_out_747[0], col_out_746[0], col_out_745[0], col_out_744[0], col_out_743[0], col_out_742[0], col_out_741[0], col_out_740[0], col_out_739[0], col_out_738[0], col_out_737[0], col_out_736[0], col_out_735[0], col_out_734[0], col_out_733[0], col_out_732[0], col_out_731[0], col_out_730[0], col_out_729[0], col_out_728[0], col_out_727[0], col_out_726[0], col_out_725[0], col_out_724[0], col_out_723[0], col_out_722[0], col_out_721[0], col_out_720[0], col_out_719[0], col_out_718[0], col_out_717[0], col_out_716[0], col_out_715[0], col_out_714[0], col_out_713[0], col_out_712[0], col_out_711[0], col_out_710[0], col_out_709[0], col_out_708[0], col_out_707[0], col_out_706[0], col_out_705[0], col_out_704[0], col_out_703[0], col_out_702[0], col_out_701[0], col_out_700[0], col_out_699[0], col_out_698[0], col_out_697[0], col_out_696[0], col_out_695[0], col_out_694[0], col_out_693[0], col_out_692[0], col_out_691[0], col_out_690[0], col_out_689[0], col_out_688[0], col_out_687[0], col_out_686[0], col_out_685[0], col_out_684[0], col_out_683[0], col_out_682[0], col_out_681[0], col_out_680[0], col_out_679[0], col_out_678[0], col_out_677[0], col_out_676[0], col_out_675[0], col_out_674[0], col_out_673[0], col_out_672[0], col_out_671[0], col_out_670[0], col_out_669[0], col_out_668[0], col_out_667[0], col_out_666[0], col_out_665[0], col_out_664[0], col_out_663[0], col_out_662[0], col_out_661[0], col_out_660[0], col_out_659[0], col_out_658[0], col_out_657[0], col_out_656[0], col_out_655[0], col_out_654[0], col_out_653[0], col_out_652[0], col_out_651[0], col_out_650[0], col_out_649[0], col_out_648[0], col_out_647[0], col_out_646[0], col_out_645[0], col_out_644[0], col_out_643[0], col_out_642[0], col_out_641[0], col_out_640[0], col_out_639[0], col_out_638[0], col_out_637[0], col_out_636[0], col_out_635[0], col_out_634[0], col_out_633[0], col_out_632[0], col_out_631[0], col_out_630[0], col_out_629[0], col_out_628[0], col_out_627[0], col_out_626[0], col_out_625[0], col_out_624[0], col_out_623[0], col_out_622[0], col_out_621[0], col_out_620[0], col_out_619[0], col_out_618[0], col_out_617[0], col_out_616[0], col_out_615[0], col_out_614[0], col_out_613[0], col_out_612[0], col_out_611[0], col_out_610[0], col_out_609[0], col_out_608[0], col_out_607[0], col_out_606[0], col_out_605[0], col_out_604[0], col_out_603[0], col_out_602[0], col_out_601[0], col_out_600[0], col_out_599[0], col_out_598[0], col_out_597[0], col_out_596[0], col_out_595[0], col_out_594[0], col_out_593[0], col_out_592[0], col_out_591[0], col_out_590[0], col_out_589[0], col_out_588[0], col_out_587[0], col_out_586[0], col_out_585[0], col_out_584[0], col_out_583[0], col_out_582[0], col_out_581[0], col_out_580[0], col_out_579[0], col_out_578[0], col_out_577[0], col_out_576[0], col_out_575[0], col_out_574[0], col_out_573[0], col_out_572[0], col_out_571[0], col_out_570[0], col_out_569[0], col_out_568[0], col_out_567[0], col_out_566[0], col_out_565[0], col_out_564[0], col_out_563[0], col_out_562[0], col_out_561[0], col_out_560[0], col_out_559[0], col_out_558[0], col_out_557[0], col_out_556[0], col_out_555[0], col_out_554[0], col_out_553[0], col_out_552[0], col_out_551[0], col_out_550[0], col_out_549[0], col_out_548[0], col_out_547[0], col_out_546[0], col_out_545[0], col_out_544[0], col_out_543[0], col_out_542[0], col_out_541[0], col_out_540[0], col_out_539[0], col_out_538[0], col_out_537[0], col_out_536[0], col_out_535[0], col_out_534[0], col_out_533[0], col_out_532[0], col_out_531[0], col_out_530[0], col_out_529[0], col_out_528[0], col_out_527[0], col_out_526[0], col_out_525[0], col_out_524[0], col_out_523[0], col_out_522[0], col_out_521[0], col_out_520[0], col_out_519[0], col_out_518[0], col_out_517[0], col_out_516[0], col_out_515[0], col_out_514[0], col_out_513[0], col_out_512[0], col_out_511[0], col_out_510[0], col_out_509[0], col_out_508[0], col_out_507[0], col_out_506[0], col_out_505[0], col_out_504[0], col_out_503[0], col_out_502[0], col_out_501[0], col_out_500[0], col_out_499[0], col_out_498[0], col_out_497[0], col_out_496[0], col_out_495[0], col_out_494[0], col_out_493[0], col_out_492[0], col_out_491[0], col_out_490[0], col_out_489[0], col_out_488[0], col_out_487[0], col_out_486[0], col_out_485[0], col_out_484[0], col_out_483[0], col_out_482[0], col_out_481[0], col_out_480[0], col_out_479[0], col_out_478[0], col_out_477[0], col_out_476[0], col_out_475[0], col_out_474[0], col_out_473[0], col_out_472[0], col_out_471[0], col_out_470[0], col_out_469[0], col_out_468[0], col_out_467[0], col_out_466[0], col_out_465[0], col_out_464[0], col_out_463[0], col_out_462[0], col_out_461[0], col_out_460[0], col_out_459[0], col_out_458[0], col_out_457[0], col_out_456[0], col_out_455[0], col_out_454[0], col_out_453[0], col_out_452[0], col_out_451[0], col_out_450[0], col_out_449[0], col_out_448[0], col_out_447[0], col_out_446[0], col_out_445[0], col_out_444[0], col_out_443[0], col_out_442[0], col_out_441[0], col_out_440[0], col_out_439[0], col_out_438[0], col_out_437[0], col_out_436[0], col_out_435[0], col_out_434[0], col_out_433[0], col_out_432[0], col_out_431[0], col_out_430[0], col_out_429[0], col_out_428[0], col_out_427[0], col_out_426[0], col_out_425[0], col_out_424[0], col_out_423[0], col_out_422[0], col_out_421[0], col_out_420[0], col_out_419[0], col_out_418[0], col_out_417[0], col_out_416[0], col_out_415[0], col_out_414[0], col_out_413[0], col_out_412[0], col_out_411[0], col_out_410[0], col_out_409[0], col_out_408[0], col_out_407[0], col_out_406[0], col_out_405[0], col_out_404[0], col_out_403[0], col_out_402[0], col_out_401[0], col_out_400[0], col_out_399[0], col_out_398[0], col_out_397[0], col_out_396[0], col_out_395[0], col_out_394[0], col_out_393[0], col_out_392[0], col_out_391[0], col_out_390[0], col_out_389[0], col_out_388[0], col_out_387[0], col_out_386[0], col_out_385[0], col_out_384[0], col_out_383[0], col_out_382[0], col_out_381[0], col_out_380[0], col_out_379[0], col_out_378[0], col_out_377[0], col_out_376[0], col_out_375[0], col_out_374[0], col_out_373[0], col_out_372[0], col_out_371[0], col_out_370[0], col_out_369[0], col_out_368[0], col_out_367[0], col_out_366[0], col_out_365[0], col_out_364[0], col_out_363[0], col_out_362[0], col_out_361[0], col_out_360[0], col_out_359[0], col_out_358[0], col_out_357[0], col_out_356[0], col_out_355[0], col_out_354[0], col_out_353[0], col_out_352[0], col_out_351[0], col_out_350[0], col_out_349[0], col_out_348[0], col_out_347[0], col_out_346[0], col_out_345[0], col_out_344[0], col_out_343[0], col_out_342[0], col_out_341[0], col_out_340[0], col_out_339[0], col_out_338[0], col_out_337[0], col_out_336[0], col_out_335[0], col_out_334[0], col_out_333[0], col_out_332[0], col_out_331[0], col_out_330[0], col_out_329[0], col_out_328[0], col_out_327[0], col_out_326[0], col_out_325[0], col_out_324[0], col_out_323[0], col_out_322[0], col_out_321[0], col_out_320[0], col_out_319[0], col_out_318[0], col_out_317[0], col_out_316[0], col_out_315[0], col_out_314[0], col_out_313[0], col_out_312[0], col_out_311[0], col_out_310[0], col_out_309[0], col_out_308[0], col_out_307[0], col_out_306[0], col_out_305[0], col_out_304[0], col_out_303[0], col_out_302[0], col_out_301[0], col_out_300[0], col_out_299[0], col_out_298[0], col_out_297[0], col_out_296[0], col_out_295[0], col_out_294[0], col_out_293[0], col_out_292[0], col_out_291[0], col_out_290[0], col_out_289[0], col_out_288[0], col_out_287[0], col_out_286[0], col_out_285[0], col_out_284[0], col_out_283[0], col_out_282[0], col_out_281[0], col_out_280[0], col_out_279[0], col_out_278[0], col_out_277[0], col_out_276[0], col_out_275[0], col_out_274[0], col_out_273[0], col_out_272[0], col_out_271[0], col_out_270[0], col_out_269[0], col_out_268[0], col_out_267[0], col_out_266[0], col_out_265[0], col_out_264[0], col_out_263[0], col_out_262[0], col_out_261[0], col_out_260[0], col_out_259[0], col_out_258[0], col_out_257[0], col_out_256[0], col_out_255[0], col_out_254[0], col_out_253[0], col_out_252[0], col_out_251[0], col_out_250[0], col_out_249[0], col_out_248[0], col_out_247[0], col_out_246[0], col_out_245[0], col_out_244[0], col_out_243[0], col_out_242[0], col_out_241[0], col_out_240[0], col_out_239[0], col_out_238[0], col_out_237[0], col_out_236[0], col_out_235[0], col_out_234[0], col_out_233[0], col_out_232[0], col_out_231[0], col_out_230[0], col_out_229[0], col_out_228[0], col_out_227[0], col_out_226[0], col_out_225[0], col_out_224[0], col_out_223[0], col_out_222[0], col_out_221[0], col_out_220[0], col_out_219[0], col_out_218[0], col_out_217[0], col_out_216[0], col_out_215[0], col_out_214[0], col_out_213[0], col_out_212[0], col_out_211[0], col_out_210[0], col_out_209[0], col_out_208[0], col_out_207[0], col_out_206[0], col_out_205[0], col_out_204[0], col_out_203[0], col_out_202[0], col_out_201[0], col_out_200[0], col_out_199[0], col_out_198[0], col_out_197[0], col_out_196[0], col_out_195[0], col_out_194[0], col_out_193[0], col_out_192[0], col_out_191[0], col_out_190[0], col_out_189[0], col_out_188[0], col_out_187[0], col_out_186[0], col_out_185[0], col_out_184[0], col_out_183[0], col_out_182[0], col_out_181[0], col_out_180[0], col_out_179[0], col_out_178[0], col_out_177[0], col_out_176[0], col_out_175[0], col_out_174[0], col_out_173[0], col_out_172[0], col_out_171[0], col_out_170[0], col_out_169[0], col_out_168[0], col_out_167[0], col_out_166[0], col_out_165[0], col_out_164[0], col_out_163[0], col_out_162[0], col_out_161[0], col_out_160[0], col_out_159[0], col_out_158[0], col_out_157[0], col_out_156[0], col_out_155[0], col_out_154[0], col_out_153[0], col_out_152[0], col_out_151[0], col_out_150[0], col_out_149[0], col_out_148[0], col_out_147[0], col_out_146[0], col_out_145[0], col_out_144[0], col_out_143[0], col_out_142[0], col_out_141[0], col_out_140[0], col_out_139[0], col_out_138[0], col_out_137[0], col_out_136[0], col_out_135[0], col_out_134[0], col_out_133[0], col_out_132[0], col_out_131[0], col_out_130[0], col_out_129[0], col_out_128[0], col_out_127[0], col_out_126[0], col_out_125[0], col_out_124[0], col_out_123[0], col_out_122[0], col_out_121[0], col_out_120[0], col_out_119[0], col_out_118[0], col_out_117[0], col_out_116[0], col_out_115[0], col_out_114[0], col_out_113[0], col_out_112[0], col_out_111[0], col_out_110[0], col_out_109[0], col_out_108[0], col_out_107[0], col_out_106[0], col_out_105[0], col_out_104[0], col_out_103[0], col_out_102[0], col_out_101[0], col_out_100[0], col_out_99[0], col_out_98[0], col_out_97[0], col_out_96[0], col_out_95[0], col_out_94[0], col_out_93[0], col_out_92[0], col_out_91[0], col_out_90[0], col_out_89[0], col_out_88[0], col_out_87[0], col_out_86[0], col_out_85[0], col_out_84[0], col_out_83[0], col_out_82[0], col_out_81[0], col_out_80[0], col_out_79[0], col_out_78[0], col_out_77[0], col_out_76[0], col_out_75[0], col_out_74[0], col_out_73[0], col_out_72[0], col_out_71[0], col_out_70[0], col_out_69[0], col_out_68[0], col_out_67[0], col_out_66[0], col_out_65[0], col_out_64[0], col_out_63[0], col_out_62[0], col_out_61[0], col_out_60[0], col_out_59[0], col_out_58[0], col_out_57[0], col_out_56[0], col_out_55[0], col_out_54[0], col_out_53[0], col_out_52[0], col_out_51[0], col_out_50[0], col_out_49[0], col_out_48[0], col_out_47[0], col_out_46[0], col_out_45[0], col_out_44[0], col_out_43[0], col_out_42[0], col_out_41[0], col_out_40[0], col_out_39[0], col_out_38[0], col_out_37[0], col_out_36[0], col_out_35[0], col_out_34[0], col_out_33[0], col_out_32[0], col_out_31[0], col_out_30[0], col_out_29[0], col_out_28[0], col_out_27[0], col_out_26[0], col_out_25[0], col_out_24[0], col_out_23[0], col_out_22[0], col_out_21[0], col_out_20[0], col_out_19[0], col_out_18[0], col_out_17[0], col_out_16[0], col_out_15[0], col_out_14[0], col_out_13[0], col_out_12[0], col_out_11[0], col_out_10[0], col_out_9[0], col_out_8[0], col_out_7[0], col_out_6[0], col_out_5[0], col_out_4[0], col_out_3[0], col_out_2[0], col_out_1[0], col_out_0[0]};


assign row_out_1 = {col_out_1024[1], col_out_1023[1], col_out_1022[1], col_out_1021[1], col_out_1020[1], col_out_1019[1], col_out_1018[1], col_out_1017[1], col_out_1016[1], col_out_1015[1], col_out_1014[1], col_out_1013[1], col_out_1012[1], col_out_1011[1], col_out_1010[1], col_out_1009[1], col_out_1008[1], col_out_1007[1], col_out_1006[1], col_out_1005[1], col_out_1004[1], col_out_1003[1], col_out_1002[1], col_out_1001[1], col_out_1000[1], col_out_999[1], col_out_998[1], col_out_997[1], col_out_996[1], col_out_995[1], col_out_994[1], col_out_993[1], col_out_992[1], col_out_991[1], col_out_990[1], col_out_989[1], col_out_988[1], col_out_987[1], col_out_986[1], col_out_985[1], col_out_984[1], col_out_983[1], col_out_982[1], col_out_981[1], col_out_980[1], col_out_979[1], col_out_978[1], col_out_977[1], col_out_976[1], col_out_975[1], col_out_974[1], col_out_973[1], col_out_972[1], col_out_971[1], col_out_970[1], col_out_969[1], col_out_968[1], col_out_967[1], col_out_966[1], col_out_965[1], col_out_964[1], col_out_963[1], col_out_962[1], col_out_961[1], col_out_960[1], col_out_959[1], col_out_958[1], col_out_957[1], col_out_956[1], col_out_955[1], col_out_954[1], col_out_953[1], col_out_952[1], col_out_951[1], col_out_950[1], col_out_949[1], col_out_948[1], col_out_947[1], col_out_946[1], col_out_945[1], col_out_944[1], col_out_943[1], col_out_942[1], col_out_941[1], col_out_940[1], col_out_939[1], col_out_938[1], col_out_937[1], col_out_936[1], col_out_935[1], col_out_934[1], col_out_933[1], col_out_932[1], col_out_931[1], col_out_930[1], col_out_929[1], col_out_928[1], col_out_927[1], col_out_926[1], col_out_925[1], col_out_924[1], col_out_923[1], col_out_922[1], col_out_921[1], col_out_920[1], col_out_919[1], col_out_918[1], col_out_917[1], col_out_916[1], col_out_915[1], col_out_914[1], col_out_913[1], col_out_912[1], col_out_911[1], col_out_910[1], col_out_909[1], col_out_908[1], col_out_907[1], col_out_906[1], col_out_905[1], col_out_904[1], col_out_903[1], col_out_902[1], col_out_901[1], col_out_900[1], col_out_899[1], col_out_898[1], col_out_897[1], col_out_896[1], col_out_895[1], col_out_894[1], col_out_893[1], col_out_892[1], col_out_891[1], col_out_890[1], col_out_889[1], col_out_888[1], col_out_887[1], col_out_886[1], col_out_885[1], col_out_884[1], col_out_883[1], col_out_882[1], col_out_881[1], col_out_880[1], col_out_879[1], col_out_878[1], col_out_877[1], col_out_876[1], col_out_875[1], col_out_874[1], col_out_873[1], col_out_872[1], col_out_871[1], col_out_870[1], col_out_869[1], col_out_868[1], col_out_867[1], col_out_866[1], col_out_865[1], col_out_864[1], col_out_863[1], col_out_862[1], col_out_861[1], col_out_860[1], col_out_859[1], col_out_858[1], col_out_857[1], col_out_856[1], col_out_855[1], col_out_854[1], col_out_853[1], col_out_852[1], col_out_851[1], col_out_850[1], col_out_849[1], col_out_848[1], col_out_847[1], col_out_846[1], col_out_845[1], col_out_844[1], col_out_843[1], col_out_842[1], col_out_841[1], col_out_840[1], col_out_839[1], col_out_838[1], col_out_837[1], col_out_836[1], col_out_835[1], col_out_834[1], col_out_833[1], col_out_832[1], col_out_831[1], col_out_830[1], col_out_829[1], col_out_828[1], col_out_827[1], col_out_826[1], col_out_825[1], col_out_824[1], col_out_823[1], col_out_822[1], col_out_821[1], col_out_820[1], col_out_819[1], col_out_818[1], col_out_817[1], col_out_816[1], col_out_815[1], col_out_814[1], col_out_813[1], col_out_812[1], col_out_811[1], col_out_810[1], col_out_809[1], col_out_808[1], col_out_807[1], col_out_806[1], col_out_805[1], col_out_804[1], col_out_803[1], col_out_802[1], col_out_801[1], col_out_800[1], col_out_799[1], col_out_798[1], col_out_797[1], col_out_796[1], col_out_795[1], col_out_794[1], col_out_793[1], col_out_792[1], col_out_791[1], col_out_790[1], col_out_789[1], col_out_788[1], col_out_787[1], col_out_786[1], col_out_785[1], col_out_784[1], col_out_783[1], col_out_782[1], col_out_781[1], col_out_780[1], col_out_779[1], col_out_778[1], col_out_777[1], col_out_776[1], col_out_775[1], col_out_774[1], col_out_773[1], col_out_772[1], col_out_771[1], col_out_770[1], col_out_769[1], col_out_768[1], col_out_767[1], col_out_766[1], col_out_765[1], col_out_764[1], col_out_763[1], col_out_762[1], col_out_761[1], col_out_760[1], col_out_759[1], col_out_758[1], col_out_757[1], col_out_756[1], col_out_755[1], col_out_754[1], col_out_753[1], col_out_752[1], col_out_751[1], col_out_750[1], col_out_749[1], col_out_748[1], col_out_747[1], col_out_746[1], col_out_745[1], col_out_744[1], col_out_743[1], col_out_742[1], col_out_741[1], col_out_740[1], col_out_739[1], col_out_738[1], col_out_737[1], col_out_736[1], col_out_735[1], col_out_734[1], col_out_733[1], col_out_732[1], col_out_731[1], col_out_730[1], col_out_729[1], col_out_728[1], col_out_727[1], col_out_726[1], col_out_725[1], col_out_724[1], col_out_723[1], col_out_722[1], col_out_721[1], col_out_720[1], col_out_719[1], col_out_718[1], col_out_717[1], col_out_716[1], col_out_715[1], col_out_714[1], col_out_713[1], col_out_712[1], col_out_711[1], col_out_710[1], col_out_709[1], col_out_708[1], col_out_707[1], col_out_706[1], col_out_705[1], col_out_704[1], col_out_703[1], col_out_702[1], col_out_701[1], col_out_700[1], col_out_699[1], col_out_698[1], col_out_697[1], col_out_696[1], col_out_695[1], col_out_694[1], col_out_693[1], col_out_692[1], col_out_691[1], col_out_690[1], col_out_689[1], col_out_688[1], col_out_687[1], col_out_686[1], col_out_685[1], col_out_684[1], col_out_683[1], col_out_682[1], col_out_681[1], col_out_680[1], col_out_679[1], col_out_678[1], col_out_677[1], col_out_676[1], col_out_675[1], col_out_674[1], col_out_673[1], col_out_672[1], col_out_671[1], col_out_670[1], col_out_669[1], col_out_668[1], col_out_667[1], col_out_666[1], col_out_665[1], col_out_664[1], col_out_663[1], col_out_662[1], col_out_661[1], col_out_660[1], col_out_659[1], col_out_658[1], col_out_657[1], col_out_656[1], col_out_655[1], col_out_654[1], col_out_653[1], col_out_652[1], col_out_651[1], col_out_650[1], col_out_649[1], col_out_648[1], col_out_647[1], col_out_646[1], col_out_645[1], col_out_644[1], col_out_643[1], col_out_642[1], col_out_641[1], col_out_640[1], col_out_639[1], col_out_638[1], col_out_637[1], col_out_636[1], col_out_635[1], col_out_634[1], col_out_633[1], col_out_632[1], col_out_631[1], col_out_630[1], col_out_629[1], col_out_628[1], col_out_627[1], col_out_626[1], col_out_625[1], col_out_624[1], col_out_623[1], col_out_622[1], col_out_621[1], col_out_620[1], col_out_619[1], col_out_618[1], col_out_617[1], col_out_616[1], col_out_615[1], col_out_614[1], col_out_613[1], col_out_612[1], col_out_611[1], col_out_610[1], col_out_609[1], col_out_608[1], col_out_607[1], col_out_606[1], col_out_605[1], col_out_604[1], col_out_603[1], col_out_602[1], col_out_601[1], col_out_600[1], col_out_599[1], col_out_598[1], col_out_597[1], col_out_596[1], col_out_595[1], col_out_594[1], col_out_593[1], col_out_592[1], col_out_591[1], col_out_590[1], col_out_589[1], col_out_588[1], col_out_587[1], col_out_586[1], col_out_585[1], col_out_584[1], col_out_583[1], col_out_582[1], col_out_581[1], col_out_580[1], col_out_579[1], col_out_578[1], col_out_577[1], col_out_576[1], col_out_575[1], col_out_574[1], col_out_573[1], col_out_572[1], col_out_571[1], col_out_570[1], col_out_569[1], col_out_568[1], col_out_567[1], col_out_566[1], col_out_565[1], col_out_564[1], col_out_563[1], col_out_562[1], col_out_561[1], col_out_560[1], col_out_559[1], col_out_558[1], col_out_557[1], col_out_556[1], col_out_555[1], col_out_554[1], col_out_553[1], col_out_552[1], col_out_551[1], col_out_550[1], col_out_549[1], col_out_548[1], col_out_547[1], col_out_546[1], col_out_545[1], col_out_544[1], col_out_543[1], col_out_542[1], col_out_541[1], col_out_540[1], col_out_539[1], col_out_538[1], col_out_537[1], col_out_536[1], col_out_535[1], col_out_534[1], col_out_533[1], col_out_532[1], col_out_531[1], col_out_530[1], col_out_529[1], col_out_528[1], col_out_527[1], col_out_526[1], col_out_525[1], col_out_524[1], col_out_523[1], col_out_522[1], col_out_521[1], col_out_520[1], col_out_519[1], col_out_518[1], col_out_517[1], col_out_516[1], col_out_515[1], col_out_514[1], col_out_513[1], col_out_512[1], col_out_511[1], col_out_510[1], col_out_509[1], col_out_508[1], col_out_507[1], col_out_506[1], col_out_505[1], col_out_504[1], col_out_503[1], col_out_502[1], col_out_501[1], col_out_500[1], col_out_499[1], col_out_498[1], col_out_497[1], col_out_496[1], col_out_495[1], col_out_494[1], col_out_493[1], col_out_492[1], col_out_491[1], col_out_490[1], col_out_489[1], col_out_488[1], col_out_487[1], col_out_486[1], col_out_485[1], col_out_484[1], col_out_483[1], col_out_482[1], col_out_481[1], col_out_480[1], col_out_479[1], col_out_478[1], col_out_477[1], col_out_476[1], col_out_475[1], col_out_474[1], col_out_473[1], col_out_472[1], col_out_471[1], col_out_470[1], col_out_469[1], col_out_468[1], col_out_467[1], col_out_466[1], col_out_465[1], col_out_464[1], col_out_463[1], col_out_462[1], col_out_461[1], col_out_460[1], col_out_459[1], col_out_458[1], col_out_457[1], col_out_456[1], col_out_455[1], col_out_454[1], col_out_453[1], col_out_452[1], col_out_451[1], col_out_450[1], col_out_449[1], col_out_448[1], col_out_447[1], col_out_446[1], col_out_445[1], col_out_444[1], col_out_443[1], col_out_442[1], col_out_441[1], col_out_440[1], col_out_439[1], col_out_438[1], col_out_437[1], col_out_436[1], col_out_435[1], col_out_434[1], col_out_433[1], col_out_432[1], col_out_431[1], col_out_430[1], col_out_429[1], col_out_428[1], col_out_427[1], col_out_426[1], col_out_425[1], col_out_424[1], col_out_423[1], col_out_422[1], col_out_421[1], col_out_420[1], col_out_419[1], col_out_418[1], col_out_417[1], col_out_416[1], col_out_415[1], col_out_414[1], col_out_413[1], col_out_412[1], col_out_411[1], col_out_410[1], col_out_409[1], col_out_408[1], col_out_407[1], col_out_406[1], col_out_405[1], col_out_404[1], col_out_403[1], col_out_402[1], col_out_401[1], col_out_400[1], col_out_399[1], col_out_398[1], col_out_397[1], col_out_396[1], col_out_395[1], col_out_394[1], col_out_393[1], col_out_392[1], col_out_391[1], col_out_390[1], col_out_389[1], col_out_388[1], col_out_387[1], col_out_386[1], col_out_385[1], col_out_384[1], col_out_383[1], col_out_382[1], col_out_381[1], col_out_380[1], col_out_379[1], col_out_378[1], col_out_377[1], col_out_376[1], col_out_375[1], col_out_374[1], col_out_373[1], col_out_372[1], col_out_371[1], col_out_370[1], col_out_369[1], col_out_368[1], col_out_367[1], col_out_366[1], col_out_365[1], col_out_364[1], col_out_363[1], col_out_362[1], col_out_361[1], col_out_360[1], col_out_359[1], col_out_358[1], col_out_357[1], col_out_356[1], col_out_355[1], col_out_354[1], col_out_353[1], col_out_352[1], col_out_351[1], col_out_350[1], col_out_349[1], col_out_348[1], col_out_347[1], col_out_346[1], col_out_345[1], col_out_344[1], col_out_343[1], col_out_342[1], col_out_341[1], col_out_340[1], col_out_339[1], col_out_338[1], col_out_337[1], col_out_336[1], col_out_335[1], col_out_334[1], col_out_333[1], col_out_332[1], col_out_331[1], col_out_330[1], col_out_329[1], col_out_328[1], col_out_327[1], col_out_326[1], col_out_325[1], col_out_324[1], col_out_323[1], col_out_322[1], col_out_321[1], col_out_320[1], col_out_319[1], col_out_318[1], col_out_317[1], col_out_316[1], col_out_315[1], col_out_314[1], col_out_313[1], col_out_312[1], col_out_311[1], col_out_310[1], col_out_309[1], col_out_308[1], col_out_307[1], col_out_306[1], col_out_305[1], col_out_304[1], col_out_303[1], col_out_302[1], col_out_301[1], col_out_300[1], col_out_299[1], col_out_298[1], col_out_297[1], col_out_296[1], col_out_295[1], col_out_294[1], col_out_293[1], col_out_292[1], col_out_291[1], col_out_290[1], col_out_289[1], col_out_288[1], col_out_287[1], col_out_286[1], col_out_285[1], col_out_284[1], col_out_283[1], col_out_282[1], col_out_281[1], col_out_280[1], col_out_279[1], col_out_278[1], col_out_277[1], col_out_276[1], col_out_275[1], col_out_274[1], col_out_273[1], col_out_272[1], col_out_271[1], col_out_270[1], col_out_269[1], col_out_268[1], col_out_267[1], col_out_266[1], col_out_265[1], col_out_264[1], col_out_263[1], col_out_262[1], col_out_261[1], col_out_260[1], col_out_259[1], col_out_258[1], col_out_257[1], col_out_256[1], col_out_255[1], col_out_254[1], col_out_253[1], col_out_252[1], col_out_251[1], col_out_250[1], col_out_249[1], col_out_248[1], col_out_247[1], col_out_246[1], col_out_245[1], col_out_244[1], col_out_243[1], col_out_242[1], col_out_241[1], col_out_240[1], col_out_239[1], col_out_238[1], col_out_237[1], col_out_236[1], col_out_235[1], col_out_234[1], col_out_233[1], col_out_232[1], col_out_231[1], col_out_230[1], col_out_229[1], col_out_228[1], col_out_227[1], col_out_226[1], col_out_225[1], col_out_224[1], col_out_223[1], col_out_222[1], col_out_221[1], col_out_220[1], col_out_219[1], col_out_218[1], col_out_217[1], col_out_216[1], col_out_215[1], col_out_214[1], col_out_213[1], col_out_212[1], col_out_211[1], col_out_210[1], col_out_209[1], col_out_208[1], col_out_207[1], col_out_206[1], col_out_205[1], col_out_204[1], col_out_203[1], col_out_202[1], col_out_201[1], col_out_200[1], col_out_199[1], col_out_198[1], col_out_197[1], col_out_196[1], col_out_195[1], col_out_194[1], col_out_193[1], col_out_192[1], col_out_191[1], col_out_190[1], col_out_189[1], col_out_188[1], col_out_187[1], col_out_186[1], col_out_185[1], col_out_184[1], col_out_183[1], col_out_182[1], col_out_181[1], col_out_180[1], col_out_179[1], col_out_178[1], col_out_177[1], col_out_176[1], col_out_175[1], col_out_174[1], col_out_173[1], col_out_172[1], col_out_171[1], col_out_170[1], col_out_169[1], col_out_168[1], col_out_167[1], col_out_166[1], col_out_165[1], col_out_164[1], col_out_163[1], col_out_162[1], col_out_161[1], col_out_160[1], col_out_159[1], col_out_158[1], col_out_157[1], col_out_156[1], col_out_155[1], col_out_154[1], col_out_153[1], col_out_152[1], col_out_151[1], col_out_150[1], col_out_149[1], col_out_148[1], col_out_147[1], col_out_146[1], col_out_145[1], col_out_144[1], col_out_143[1], col_out_142[1], col_out_141[1], col_out_140[1], col_out_139[1], col_out_138[1], col_out_137[1], col_out_136[1], col_out_135[1], col_out_134[1], col_out_133[1], col_out_132[1], col_out_131[1], col_out_130[1], col_out_129[1], col_out_128[1], col_out_127[1], col_out_126[1], col_out_125[1], col_out_124[1], col_out_123[1], col_out_122[1], col_out_121[1], col_out_120[1], col_out_119[1], col_out_118[1], col_out_117[1], col_out_116[1], col_out_115[1], col_out_114[1], col_out_113[1], col_out_112[1], col_out_111[1], col_out_110[1], col_out_109[1], col_out_108[1], col_out_107[1], col_out_106[1], col_out_105[1], col_out_104[1], col_out_103[1], col_out_102[1], col_out_101[1], col_out_100[1], col_out_99[1], col_out_98[1], col_out_97[1], col_out_96[1], col_out_95[1], col_out_94[1], col_out_93[1], col_out_92[1], col_out_91[1], col_out_90[1], col_out_89[1], col_out_88[1], col_out_87[1], col_out_86[1], col_out_85[1], col_out_84[1], col_out_83[1], col_out_82[1], col_out_81[1], col_out_80[1], col_out_79[1], col_out_78[1], col_out_77[1], col_out_76[1], col_out_75[1], col_out_74[1], col_out_73[1], col_out_72[1], col_out_71[1], col_out_70[1], col_out_69[1], col_out_68[1], col_out_67[1], col_out_66[1], col_out_65[1], col_out_64[1], col_out_63[1], col_out_62[1], col_out_61[1], col_out_60[1], col_out_59[1], col_out_58[1], col_out_57[1], col_out_56[1], col_out_55[1], col_out_54[1], col_out_53[1], col_out_52[1], col_out_51[1], col_out_50[1], col_out_49[1], col_out_48[1], col_out_47[1], col_out_46[1], col_out_45[1], col_out_44[1], col_out_43[1], col_out_42[1], col_out_41[1], col_out_40[1], col_out_39[1], col_out_38[1], col_out_37[1], col_out_36[1], col_out_35[1], col_out_34[1], col_out_33[1], col_out_32[1], col_out_31[1], col_out_30[1], col_out_29[1], col_out_28[1], col_out_27[1], col_out_26[1], col_out_25[1], col_out_24[1], col_out_23[1], col_out_22[1], col_out_21[1], col_out_20[1], col_out_19[1], col_out_18[1], col_out_17[1], col_out_16[1], col_out_15[1], col_out_14[1], col_out_13[1], col_out_12[1], col_out_11[1], col_out_10[1], col_out_9[1], col_out_8[1], col_out_7[1], col_out_6[1], col_out_5[1], col_out_4[1], col_out_3[1], col_out_2[1], col_out_1[1], col_out_0[1]};

//---------------------------------------------------------


endmodule
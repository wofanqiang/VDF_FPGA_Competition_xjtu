module xpb_5_355
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h2d5662df0dce901cc480418de3666da7e66d764b952ec5ef4776df00277cdf767a002c0082e929b56775811476d6decd01d7605b498c1c0dc7ac7bb8a4359a236ed4ca2717ea52fe74cdc4f5008fc34d4ab7a0570e3be2f2df81a683139249b32a8f93f4e6345b9bd00f2f848f2436c727f38357269a37c9e219eb77e8096b9c;
    5'b00010 : xpb = 1024'h5aacc5be1b9d20398900831bc6ccdb4fccdaec972a5d8bde8eedbe004ef9beecf400580105d2536aceeb0228edadbd9a03aec0b69318381b8f58f771486b3446dda9944e2fd4a5fce99b89ea011f869a956f40ae1c77c5e5bf034d0627249366551f27e9cc68b737a01e5f091e486d8e4fe706ae4d346f93c433d6efd012d738;
    5'b00011 : xpb = 1024'h8803289d296bb0564d80c4a9aa3348f7b34862e2bf8c51cdd6649d0076769e636e00840188bb7d203660833d64849c6705862111dca4542957057329eca0ce6a4c7e5e7547bef8fb5e694edf01af49e7e026e1052ab3a8d89e84f3893ab6dd197faebbdeb29d12d3702d8e8dad6ca45577da8a0573cea75da64dc267b81c42d4;
    5'b00100 : xpb = 1024'h4ac4626754c0baa46fb8e607d3f6f4e283fd5fd7f4377459ffec2aaeaf0d0d1e4b83289417e2846fe77c50af7fd6a69a3435987037d9feb6e12af845603f3dc4703f3edb0184eb4c09d11316963490436d987c3ac695ebac87a0811941e843a7b36bda9e80875e1b97cd73344c0b4f350f42e7a4a1d81f741f832db17434805;
    5'b00101 : xpb = 1024'h3202a905831a9bc70b7bcfee60a5dcf60ead4c4914723d34e775a1ab126db0485eb85e89c46751fc65ed461f6ed44936a51ab9e24d09bbf935bf2b3cfa398dffb5d8be14c802a1b3356ad62669f30c518191281abaa541ada7fbae94a7b0cdeda5c6519ece3cd17d898c06b7d3e4ebba78e7b1d170b7b9c124121e52ff4cb3a1;
    5'b00110 : xpb = 1024'h5f590be490e92be3cffc117c440c4a9df51ac294a9a103242eec80ab39ea8fbed8b88a8a47507bb1cd62c733e5ab2803a6f21a3d9695d806fd6ba6f59e6f282324ad883bdfecf4b1aa389b1b6a82cf9ecc48c871c8e124a0877d5517bb4317a0d055e593b4712d19599b363c63092281a0db35289751f18b062c09cae7561f3d;
    5'b00111 : xpb = 1024'h8caf6ec39eb7bc00947c530a2772b845db8838e03ecfc91376635fab61676f3552b8b68aca39a56734d848485c8206d0a8c97a98e021f414c51822ae42a4c24693825262f7d747b01f0660106b1292ec170068c8d71d079366fefb9aced56153fae579889aa588b529aa65c0f22d5948c8ceb87fbdec2954e845f542cf5f8ad9;
    5'b01000 : xpb = 1024'h9588c4cea9817548df71cc0fa7ede9c507fabfafe86ee8b3ffd8555d5e1a1a3c970651282fc508dfcef8a15effad4d34686b30e06fb3fd6dc255f08ac07e7b88e07e7db60309d69813a2262d2c692086db30f8758d2bd7590f41023283d0874f66d7b53d010ebc372f9ae66898169e6a1e85cf4943b03ee83f065b62e86900a;
    5'b01001 : xpb = 1024'h36aeef2bf866a77152775e4edde54c4436ed224693b5b47a87746455fd5e811a4370911305e57a4364650b2a66d1b3a0485e136950875be4a3d1dac1503d81dbfcdcb202781af067f607e757d3565555b86aafde670ea0687075b6a63bcf522820fd0f48b645475f4308ddeb18a5a0adc9dbe04bbad53bb8660a512e168ffba6;
    5'b01010 : xpb = 1024'h6405520b0635378e16f79fdcc14bb9ec1d5a989228e47a69ceeb435624db6090bd70bd1388cea3f8cbda8c3edda8926d4a3573c49a1377f26b7e5679f4731bff6bb17c29900543666ad5ac4cd3e618a303225035754a835b4ff75d294f619bdb4b8ca33d9c79a2fb13180d6fa7c9d774f1cf63a2e16f738248243ca5fe996742;
    5'b01011 : xpb = 1024'h915bb4ea1403c7aadb77e16aa4b2279403c80eddbe134059166222564c5840073770e9140bb7cdae33500d53547f713a4c0cd41fe39f9400332ad23298a8b622da864650a7ef9664dfa37141d475dbf04dd9f08c8386664e2f7903ac62f3e58e761c373282adfe96e3273cf436ee0e3c19c2e6fa0809ab4c2a3e281de6a2d2de;
    5'b01100 : xpb = 1024'he04d2735fe422fed4f2ab2177be4dea78bf81f87dca65d0dffc4800c0d27275ae28979bc47a78d4fb674f20e7f83f3ce9ca0c950a78dfc24a380e8d020bdb94d50bdbc91048ec1e41d733943c29db0ca48c974b053c1c30596e1834bc5b8caf71a438fdb81961a52c768599ce421ed9f2dc8b6ede5885e5c5e8989145c9d80f;
    5'b01101 : xpb = 1024'h3b5b35526db2b31b9972ecaf5b24bb925f2cf84412f92bc027732700e84f51ec2828c39c4763a28a62dcd0355ecf1e09eba16cf05404fbd011e48a45a64175b843e0a5f028333f1cb6a4f8893cb99e59ef4437a21377ff2338efbeb7cfedd6629c33ccf29e4dbd40fc85b51e5d6655a11ad00ec604f2bdafa80284092dd343ab;
    5'b01110 : xpb = 1024'h68b198317b8143385df32e3d3e8b293a459a6e8fa827f1af6eea06010fcc3162a228ef9cca4ccc3fca525149d5a5fcd6ed78cd4b9d9117ddd99105fe4a770fdbb2b57017401d921b2b72bd7e3d4961a739fbd7f921b3e2161871653ae3802015c6c360e7848218dccc94e4a2ec8a8c6842c3921d2b8cf5798a1c6f8115dcaf47;
    5'b01111 : xpb = 1024'h9607fb10894fd35522736fcb21f196e22c07e4db3d56b79eb660e501374910d91c291b9d4d35f5f531c7d25e4c7cdba3ef502da6e71d33eba13d81b6eeaca9ff218a3a3e5807e519a04082733dd924f484b378502fefc508f7f30bbdf71269c8f152f4dc6ab674789ca414277baec32f6ab7157452272d436c365af8fde61ae3;
    5'b10000 : xpb = 1024'h12b11899d5302ea91bee3981f4fdbd38a0ff57f5fd0ddd167ffb0aababc3434792e0ca2505f8a11bf9df142bdff5a9a68d0d661c0df67fadb84abe11580fcf711c0fcfb6c0613ad3027444c5a58d2410db661f0eb1a57aeb21e82046507a10e9ecdaf6a7a021d786e5f35ccd1302d3cd43d0b9e9287607dd07e0cb6c5d0d2014;
    5'b10001 : xpb = 1024'h40077b78e2febec5e06e7b0fd8642ae0876cce41923ca305c771e9abd34022be0ce0f62588e1cad16154954056cc88738ee4c67757829bbb7ff739c9fc4569948ae499ddd84b8dd1774209baa61ce75e261dbf65bfe15dde0169c6c9640c5a9d176a8a9c86563322b6028c51a2270a946bc43d404f103fa6e9fab6e445168bb0;
    5'b10010 : xpb = 1024'h6d5dde57f0cd4ee2a4eebc9dbbca98886dda448d276b68f50ee8c8abfabd023486e122260bcaf486c8ca1654cda3674090bc26d2a10eb7c947a3b582a07b03b7f9b96404f035e0cfec0fceafa6acaaab70d55fbcce1d40d0e0eb6d4c779ea45041fa1e916c8a8ebe8611bbd6314b415b93b7c09775aa7770cc14a25c2d1ff74c;
    5'b10011 : xpb = 1024'h9ab44136fe9bdeff696efe2b9f3106305447bad8bc9a2ee4565fa7ac2239e1ab00e14e268eb41e3c303f9769447a460d9293872dea9ad3d70f50313b44b09ddb688e2e2c082033ce60dd93a4a73c6df8bb8d0013dc5923c3c06d13cf8b30ee036c89b28652beea5a5620eb5ac06f7822bbab43ee9c44af3aae2e8dd4152962e8;
    5'b10100 : xpb = 1024'h175d5ec04a7c3a5362e9c7e2723d2c86c93f2df37c51545c1ff9cd5696b414197798fcae4776c962f856d936d7f314103050bfa311741f99265d6d95ae13c34d6313c3a470798987c31155f70ef06d15123fa6d25e0ed9a5ea622857e49895246811b451882a4d689f70340057c388c094c4e863729389d449d8fe4774506819;
    5'b10101 : xpb = 1024'h44b3c19f584aca70276a097055a39a2eafaca43f11801a4b6770ac56be30f38ff19928aeca5ff3185fcc5a4b4ec9f2dd32281ffe5b003ba6ee09e94e52495d70d1e88dcb8863dc8637df1aec0f8030625cf747296c4abc98c9e3cedaf82aded792a148466e5ea9046f7f6384e6e7bf87bcb86bba992dc19e2bf2e9bf5c59d3b5;
    5'b10110 : xpb = 1024'h720a247e66195a8cebea4afe390a07d6961a1a8aa6aee03aaee78b56e5add3066b9954af4d491ccdc741db5fc5a0d1aa33ff8059a48c57b4b5b66506f67ef79440bd57f2a04e2f84acacdfe1100ff3afa7aee7807a869f8ba965755e0bbd288abd30dc3b549304a03f8e9309760bf64ee4abef11bfc7f9680e0cd53744633f51;
    5'b10111 : xpb = 1024'h9f60875d73e7eaa9b06a8c8c1c70757e7c8790d63bdda629f65e6a570d2ab27ce59980afd03246832eb75c743c77b07735d6e0b4ee1873c27d62e0bf9ab491b7af922219b8388283217aa4d6109fb6fcf26687d788c2827e88e71be11f4f723de7c070303ac7603c0f9dc28e05302d160c9f7268e6623131f026c0af2c6caaed;
    5'b11000 : xpb = 1024'h1c09a4e6bfc845fda9e55642ef7c9bd4f17f03f0fb94cba1bff8900181a4e4eb5c512f3788f4f1a9f6ce9e41cff07e79d394192a14f1bf8494701d1a0417b729aa17b7922091d83c83ae67287853b61949192e960a783860b2dc306978b7195ee34871fb7032c34a58ed0b339c843db3e5b916ddbcb10bcb8bd131228b93b01e;
    5'b11001 : xpb = 1024'h496007c5cd96d61a6e6597d0d2e3097cd7ec7a3c90c39191076f6f01a921c461d6515b380bde1b5f5e441f5646c75d46d56b79855e7ddb925c1c98d2a84d514d18ec81b9387c2b3af87c2c1d78e3796693d0ceed18b41b53925dd6ec8c4963120dd805f056671ee628fc3ab82ba8747b0dac9a34e34b43956deb1c9a739d1bba;
    5'b11010 : xpb = 1024'h76b66aa4db65663732e5d95eb6497724be59f08825f257804ee64e01d09ea3d8505187388ec74514c5b9a06abd9e3c13d742d9e0a809f7a023c9148b4c82eb7087c14be050667e396d49f11279733cb3de886f4426effe4671df7d6f9fdbacc5386799e53c9b7a81f90b6a3cbaccab4235a01d8c09e57b5f500508125ba68756;
    5'b11011 : xpb = 1024'ha40ccd83e933f653f7661aec99afe4cca4c766d3bb211d6f965d2d01f81b834eca51b33911b06eca2d2f217f34751ae0d91a3a3bf19613adeb759043f0b88593f69616076850d137e217b6077a03000129400f9b352be139516123f2b36df67862f72dda22cfd61dc91a99c149f0e2095d93a0e3307fb329321ef38a43aff2f2;
    5'b11100 : xpb = 1024'h20b5eb0d351451a7f0e0e4a36cbc0b2319bed9ee7ad842e75ff752ac6c95b5bd410961c0ca7319f0f546634cc7ede8e376d772b1186f5f700282cc9e5a1bab05f11bab7fd0aa26f1444b7859e1b6ff1d7ff2b659b6e1971b7b56387b0cd59d995e7f2fa5583b392c1269e266e144f2a736ad455806ce8dc2cdc963fda2d6f823;
    5'b11101 : xpb = 1024'h4e0c4dec42e2e1c4b5612631502278cb002c503a100708d6a76e31ac94129533bb098dc14d5c43a65cbbe4613ec4c7b078aed30c61fb7b7dca2f4856fe5145295ff075a6e89479efb9193d4ee246c26acaaa56b0c51d7a0e5ad7defe2067e74c890ec39a3e6f94c7e27911eb7069296e5ea0c8af2d68c58cafe34f758ae063bf;
    5'b11110 : xpb = 1024'h7b62b0cb50b171e179e167bf3388e672e699c685a535cec5eee510acbb8f74aa3509b9c1d0456d5bc4316575b59ba67d7a863367ab87978b91dbc40fa286df4ccec53fce007eccee2de70243e2d685b81561f707d3595d013a59858133fa30ffb39e578f24a3f063b288416fff8d603586944c065402fd5691fd3aed72e9cf5b;
    5'b11111 : xpb = 1024'ha8b913aa5e8001fe3e61a94d16ef541acd073cd13a6494b5365beface30c5420af09e5c2532e97112ba6e68a2c72854a7c5d93c2f513b39959883fc846bc79703d9a09f518691feca2b4c738e36649056019975ee1953ff419db2c04478c7ab2de2deb840ad84bff829770f48eb196fcae87cf5d7a9d3520741726655af33af7;
    endcase
end

endmodule

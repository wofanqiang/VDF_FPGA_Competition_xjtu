module xpb_5_380
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h283c265e74be29bbe81c2e62141bdd6d3848413b093515eda09edf43fcc8f883cda05dabbb104146c200f01b92b780b1daa7f71d58da9a1f50f1ed93c9857137847c1ad4dd7f8363e482db669632b5d43e198a096938e87267e01b18a025f659125611b33eac13d751754ba0f146a71d523c1e6d26def9d42931327c914606db;
    5'b00010 : xpb = 1024'h50784cbce97c5377d0385cc42837bada70908276126a2bdb413dbe87f991f1079b40bb577620828d8401e037256f0163b54fee3ab1b5343ea1e3db27930ae26f08f835a9baff06c7c905b6cd2c656ba87c331412d271d0e4cfc03631404becb224ac23667d5827aea2ea9741e28d4e3aa4783cda4dbdf3a8526264f9228c0db6;
    5'b00011 : xpb = 1024'h78b4731b5e3a7d33b8548b263c539847a8d8c3b11b9f41c8e1dc9dcbf65ae98b68e119033130c3d44602d052b82682158ff7e5580a8fce5df2d5c8bb5c9053a68d74507e987e8a2bad889233c298217cba4c9e1c3baab95737a05149e071e30b37023519bc043b85f45fe2e2d3d3f557f6b45b47749ced7c7b939775b3d21491;
    5'b00100 : xpb = 1024'ha0f09979d2f8a6efa070b988506f75b4e12104ec24d457b6827b7d0ff323e20f368176aeec41051b0803c06e4ade02c76a9fdc75636a687d43c7b64f2615c4de11f06b5375fe0d8f920b6d9a58cad750f8662825a4e3a1c99f806c628097d964495846ccfab04f5d45d52e83c51a9c7548f079b49b7be750a4c4c9f245181b6c;
    5'b00101 : xpb = 1024'h187f7a8285c89be2bd87701354310bd0a7f342f65891cd2ca53da2fe3cea2d8b00d956e1dd2ac7d32aa67142fa3772aee12dabac99923250e41a6484b4c8c164221d5179a3ec93ae63f4465e5621c8f4427ab89681965d2b51d3f58066932d2b2ca6c65688936aa7108a9345be911d694c52b93f720f83f48786816a4d7bbbdc;
    5'b00110 : xpb = 1024'h40bba0e0fa86c59ea5a39e75684ce93de03b843161c6e31a45dc824239b3260ece79b48d983b0919eca7615e8ceef360bbd5a2c9f26ccc70350c52187e4e329ba6996c4e816c1712487721c4ec547ec88094429feacf459db9b4109906b923843efcd809c73f7e7e61ffdee6afd7c4869e8ed7ac98ee7dc8b0b7b3e6dec1c2b7;
    5'b00111 : xpb = 1024'h68f7c73f6f44ef5a8dbfccd77c68c6ab1883c56c6afbf907e67b6186367c1e929c1a1239534b4a60aea8517a1fa67412967d99e74b47668f85fe3fac47d3a3d32b1587235eeb9a762cf9fd2b8287349cbeadcca954082e1021942bb1a6df19dd5152e9bd05eb9255b3752a87a11e6ba3f0caf619bfcd779cd9e8e6637007c992;
    5'b01000 : xpb = 1024'h9133ed9de403191675dbfb399084a41850cc06a774310ef5871a40ca3345171669ba6fe50e5b8ba770a94195b25df4c471259104a42200aed6f02d401159150aaf91a1f83c6b1dda117cd89218b9ea70fcc756b2bd411682897446ca4705103663a8fb704497a62d04ea7628926512c143071486e6ac7171031a18e0014dd06d;
    5'b01001 : xpb = 1024'h8c2cea696d30e0992f2b1c494463a34179e44b1a7ee846ba9dc66b87d0b629234125017ff454e5f934bf26a61b764abe7b3603bda49ca827742db75a00c1190bfbe881e6a59a3f8e365b1561610dc1446dbe72399f3d1e43bc7cfe82d0063fd46f77af9d27ac176cf9fdaea8bdb93b546695411bd400e14e5dbd05809b170dd;
    5'b01010 : xpb = 1024'h30fef5050b9137c57b0ee026a86217a14fe685ecb1239a594a7b45fc79d45b1601b2adc3ba558fa6554ce285f46ee55dc25b5759332464a1c834c909699182c8443aa2f347d9275cc7e88cbcac4391e884f5712d032cba56a3a7eb00cd265a56594d8cad1126d54e2115268b7d223ad298a5727ee41f07e90f0d02d49af777b8;
    5'b01011 : xpb = 1024'h593b1b63804f6181632b0e88bc7df50e882ec727ba58b046eb1a2540769d5399cf530b6f7565d0ed174dd2a18726660f9d034e768bfefec11926b69d3316f3ffc8b6bdc82558aac0ac6b6823427647bcc30efb366c65a2c90b8806196d4c50af6ba39e604fd2e925728a722c6e68e1efeae190ec0afe01bd383e35512c3d7e93;
    5'b01100 : xpb = 1024'h817741c1f50d8b3d4b473cead099d27bc0770862c38dc6348bb9048473664c1d9cf3691b30761233d94ec2bd19dde6c177ab4593e4d998e06a18a430fc9c65374d32d89d02d82e2490ee4389d8a8fd910128853fd59e8b3b736821320d7247087df9b0138e7efcfcc3ffbdcd5faf890d3d1daf5931dcfb91616f67cdbd83856e;
    5'b01101 : xpb = 1024'ha9b3682069cbb4f933636b4ce4b5afe8f8bf499dccc2dc222c57e3c8702f44a16a93c6c6eb86537a9b4fb2d8ac95677352533cb13db432ffbb0a91c4c621d66ed1aef371e057b18875711ef06edbb3653f420f493ed773addb483c4aad983d61904fc1c6cd2b10d41575096e50f6302a8f59cdc658bbf5658aa09a4a4ec98c49;
    5'b01110 : xpb = 1024'h214249291c9ba9ec507a21d7e8774604bf9187a8008051984f1a09b6b9f5901d34eba6f9dc701632bdf263ad5beed75ac8e10be873dbfcd35b5d3ffa54d4d2f4e1dbd9980e4637a74759f7b46c32a50889569fba1b8a2f0f8d9bc56893939128739e41505b0e2c1de02a6e304a6cb11e92bc0d512f4f92096d6251c2572d2cb9;
    5'b01111 : xpb = 1024'h497e6f879159d3a838965039fc932371f7d9c8e309b56785efb8e8fab6be88a1028c04a5978057797ff353c8eea6580ca3890305ccb696f2ac4f2d8e1e5a442c6657f46cebc5bb0b2bdcd31b02655adcc77029c384c31781f57be08133b9878185f4530399ba3ff5319fb9d13bb3583be4f82bbe562e8bdd9693843ee8733394;
    5'b10000 : xpb = 1024'h71ba95e60617fd6420b27e9c10af00df30220a1e12ea7d739057c83eb3878124d02c6251529098c041f443e4815dd8be7e30fa2325913111fd411b21e7dfb563ead40f41c9453e6f105fae81989810b10589b3ccedfbfff45d5bfb99d3df7dda984a64b6d86653cc831505722cf9ff5937344a2b7d0d85b1bfc4b6bb79b93a6f;
    5'b10001 : xpb = 1024'h99f6bc447ad6272008ceacfe24cade4c686a4b591c1f936130f6a782b05079a89dccbffd0da0da0703f534001415597058d8f1407e6bcb314e3308b5b165269b6f502a16a6c4c1d2f4e289e82ecac68543a33dd65734e866c53c16b274057433aaa0766a171267a3d48a51131e40a67689706898a3ec7f85e8f5e9380aff414a;
    5'b10010 : xpb = 1024'h11859d4d2da61c1325e56389288c74682f3c89634fdd08d753b8cd70fa16c5246824a02ffe8a9cbf2697e4d4c36ec957cf66c077b4939504ee85b6eb401823217f7d103cd4b347f1c6cb62ac2c21b8288db7ce4733e7a3c8778f9fd05a00c7fa8deef5f3a4f582ed9f3fb5d517b7276a8cd2a8237a801c29cbb7a0b01362e1ba;
    5'b10011 : xpb = 1024'h39c1c3aba26445cf0e0191eb3ca851d56784ca9e59121ec4f457acb4f6dfbda835c4fddbb99ade05e898d4f056264a09aa0eb7950d6e2f243f77a47f099d945903f92b11b232cb55ab4e3e12c2546dfccbd158509d208c3adf6fbae8fa26be53a04507a6e3a196c4f0b5017608fdce87df0ec690a15f15fdf4e8d32ca4a8e895;
    5'b10100 : xpb = 1024'h61fdea0a17226f8af61dc04d50c42f429fcd0bd9624734b294f68bf8f3a8b62c03655b8774ab1f4caa99c50be8ddcabb84b6aeb26648c94390699212d3230590887545e68fb24eb98fd11979588723d109eae25a065974ad474fd6019a4cb4acb29b195a224daa9c422a4d16fa4475a5314ae4fdc83e0fd21e1a05a935eeef70;
    5'b10101 : xpb = 1024'h8a3a10688be09946de39eeaf64e00cafd8154d146b7c4aa035956b3cf071aeafd105b9332fbb60936c9ab5277b954b6d5f5ea5cfbf236362e15b7fa69ca876c80cf160bb6d31d21d7453f4dfeeb9d9a548046c636f925d1faf2ff11a3a72ab05c4f12b0d60f9be73939f98b7eb8b1cc28387036aef1d09a6474b3825c734f64b;
    5'b10110 : xpb = 1024'h1c8f1713eb08e39fb50a53a68a1a2cb9ee78b1e9f39c0165857912b3a37fa2b9b5d996620a5234b8f3d65fc2aeebb54d5ec7506f54b2d3681ae2ddc2b5b734e1d1e46e19b20583c463ccda3ec10cb489218fcd44c45188161837a38206dfecca83faa96eedcd9bd5e54fd79e5019db686e942f5c5b0a64a2a0cef9dcf9896bb;
    5'b10111 : xpb = 1024'h2a0517cfb36eb7f5e36cd39c7cbd8038d72fcc59a86ed603f8f6706f3700f2af68fdf711dbb56492513e5617bda63c06b0946c244e25c755d2a01b6ff4e0e485a19a61b6789fdba02abfa90a8243811cd03286ddb57e00f3c9639550c093f525ba95bc4a2d88ed94afca491ad64844d3d9256162ec8fa01e533e221a60de9d96;
    5'b11000 : xpb = 1024'h52413e2e282ce1b1cb8901fe90d95da60f780d94b1a3ebf199954fb333c9eb33369e54bd96c5a5d9133f4633505dbcb88b3c6341a700617523920903be6655bd26167c8b561f5f040f428471187636f10e4c10e71eb6e9663143b06960b9eb7eccebcdfd6c35016c013f94bbc78eebf12b617fd0136e99f27c6f5496f224a471;
    5'b11001 : xpb = 1024'h7a7d648c9ceb0b6db3a53060a4f53b1347c04ecfbad901df3a342ef73092e3b7043eb26951d5e71fd540364ee3153d6a65e45a5effdafb947483f69787ebc6f4aa929760339ee267f3c55fd7aea8ecc54c659af087efd1d89923cb8200dfe1d7df41dfb0aae1154352b4e05cb8d5930e7d9d9e3d3a4d93c6a5a08713836aab4c;
    5'b11010 : xpb = 1024'ha2b98aeb11a935299bc15ec2b91118808008900ac40e17ccdad30e3b2d5bdc3ad1df10150ce628669741266a75ccbe1c408c517c58b595b3c575e42b5171382c2f0eb235111e65cbd8483b3e44dba2998a7f24f9f128ba4b0103e69aa105d830f197f163e98d291aa42a2bfdaa1c3a2bcfd9bcaa612c8d9aced1b99014b0b227;
    5'b11011 : xpb = 1024'h1a486bf3c4792a1cb8d8154dbcd2ae9c46dace14f7cb8d42fd953429772227b69c36f047fdcfeb1eb9e3d73f25262e03b71a20b38edd5f8765c89260e02434b23f3b985b3f0cebeaaa3114024232943cd493b56acddb75acb3576fb887012bf7d4e670ed777044646edf90bfa392bb1fd33bfc3537c02a3eb19371081d145297;
    5'b11100 : xpb = 1024'h42849252393753d8a0f443afd0ee8c097f230f500100a3309e34136d73eb203a69d74df3b8e02c657be4c75ab7ddaeb591c217d0e7b7f9a6b6ba7ff4a9a9a5e9c3b7b3301c8c6f4e8eb3ef68d8654a1112ad3f7437145e1f1b378ad127272250e73c82a0b61c583bc054dc6094d9623d25781aa25e9f2412dac4a384ae5a5972;
    5'b11101 : xpb = 1024'h6ac0b8b0adf57d9489107211e50a6976b76b508b0a35b91e3ed2f2b170b418be3777ab9f73f06dac3de5b7764a952f676c6a0eee409293c607ac6d88732f17214833ce04fa0bf2b27336cacf6e97ffe550c6c97da04d46918317a5e9c74d18a9f9929453f4c86c1311ca28018620095a77b4390f857e1de703f5d6013fa0604d;
    5'b11110 : xpb = 1024'h92fcdf0f22b3a750712ca073f92646e3efb391c6136acf0bdf71d1f56d7d11420518094b2f00aef2ffe6a791dd4cb0194712060b996d2de5589e5b1c3cb48858ccafe8d9d78b761657b9a63604cab5b98ee0538709862f03eaf7c10267730f030be8a60733747fea633f73a27766b077c9f0577cac5d17bb2d27087dd0e66728;
    5'b11111 : xpb = 1024'ha8bc017d5839c438e4356fefce7dcffb685cfd0472844820233f7e3b7435cbdcf6fe97e1fea71ab228958668ca62000bd9fd542cf94f7b8f8f10951cb6784dedcdccf000579fc3529a27efa0221a75cd8f4e3f7e638ea659d4b4a204d6e62c9ef372590c1579b342df4d86470dd316bcd52970782f0b45f0fe8bff5d94a0798;
    endcase
end

endmodule

module xpb_5_770
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h7c97a7092f51e523d34b019b9aafc324afde0d15159f1271d48dba5dc3fdc1df42f88320327a70f6dab54f3dc8784099d7ba23c70affc3baa9d01ef93058bb73cbc6b07417ff23ef582afbc179c58388401fbff66c016f5a58e2fc54f5d9db100d4f9bd9a6c8000c5b5f54218dd786d65204f0e60c1c736281c3636ddbcf0ac1;
    5'b00010 : xpb = 1024'h488208bc9cb5957edb908b6025053ef7ee4616f955c6846c2b3ebb65d4f8d6b682a888c79ace635f160c5f34ad9270694b5a1fa7f34cb729a300fe9425df0236233e2c39806d4a999dbbf4e05aaf42df8c3a86544b7cb1a3fc3966af3189138deb97a5899cc7078b2ffec16423dee783553002e9c7ed8994bd174bd72ebbaf17;
    5'b00011 : xpb = 1024'h146c6a700a1945d9e3d61524af5abacb2cae20dd95edf66681efbc6de5f3eb8dc2588e6f032255c751636f2b92aca038befa1b88db99aa989c31de2f1b6548f87ab5a7fee8db7143e34cedff3b990236d8554cb22af7f3ed9f8fd1096d384c0bc9dfaf3992c60f0a049e2ea6b9e64830585b14ed83be9fc6f86b344081a8536d;
    5'b00100 : xpb = 1024'h91041179396b2afdb72116c04a0a7defdc8c2df2ab8d08d8567d76cba9f1ad6d0551118f359cc6be2c18be695b24e0d296b43f4fe6996e534601fd284bbe046c467c587300da95333b77e9c0b55e85bf18750ca896f96347f872cd5e6312271bd72f4b13398e0f165ffd82c847bdcf06aa6005d38fdb13297a2e97ae5d775e2e;
    5'b00101 : xpb = 1024'h5cee732ca6cedb58bf66a084d45ff9c31af437d6ebb47ad2ad2e77d3baecc244450117369df0b926676fce60403f10a20a543b30cee661c23f32dcc341444b2e9df3d4386948bbdd8108e2df96484516648fd3067674a5919bc937b89ec15f99b57754c32f8d1695349cf00addc52fb3ad8b17d74bac295bb5828017b0640284;
    5'b00110 : xpb = 1024'h28d8d4e014328bb3c7ac2a495eb57596595c41bb2bdbeccd03df78dbcbe7d71b84b11cde0644ab8ea2c6de57255940717df43711b73355313863bc5e36ca91f0f56b4ffdd1b6e287c699dbfe7732046db0aa996455efe7db3f1fa212da70981793bf5e73258c1e14093c5d4d73cc9060b0b629db077d3f8df0d668810350a6da;
    5'b00111 : xpb = 1024'ha5707be9438470d79af72be4f96538bb093a4ed0417aff3ed86d33398fe598fac7a99ffe38bf1c857d7c2d94edd1810b55ae5ad8c23318ebe233db5767234d64c1320071e9b606771ec4d7bff0f787f5f0ca595ac1f1573598029e67d04a7327a10efa4ccc541e20649bb16f01a4173702bb1ac11399b2f07299cbeedf1fb19b;
    5'b01000 : xpb = 1024'h715add9cb0e82132a33cb5a983bab48e47a258b481a271392f1e3441a0e0add20759a5a5a1130eedb8d33d8bd2ebb0dac94e56b9aa800c5adb64baf25ca9942718a97c3752242d216455d0ded1e1474d3ce51fb8a16c997f3b5908c20bf9aba57f5703fcc253259f393b1eb197ab77e405e62cc4cf6ac922adedb458320c55f1;
    5'b01001 : xpb = 1024'h3d453f501e4bd18dab823f6e0e103061860a6298c1c9e33385cf3549b1dbc2a94709ab4d09670155f42a4d82b805e0aa3cee529a92ccffc9d4959a8d522fdae97020f7fcba9253cba9e6c9fdb2cb06a488ffe61680e7dbc8deaf731c47a8e4235d9f0dacb8522d1e0dda8bf42db2d89109113ec88b3bdf54e9419cc184f8fa47;
    5'b01010 : xpb = 1024'h92fa1038baf81e8b3c7c9329865ac34c4726c7d01f1552ddc803651c2d6d78086b9b0f471baf3be2f815d799d201079b08e4e7b7b19f338cdc67a2847b621abc79873c223007a75ef77c31c93b4c5fbd51aac7460631e128205dd7683581ca13be7175cae51349ce279f936c3ba393e0c3c50cc470cf5872495852ad7e59e9d;
    5'b01011 : xpb = 1024'h85c7480cbb01670c8712cace33156f59745079921790679fb10df0af86d4995fc9b23414a43564b50a36acb765985113884872428619b6f377969921780edd1f935f24363aff9e6547a2bede0d7a4984153a6c6acc648d6cdae8d9cb7931f7b14936b336551934a93dd94d585191c0145e4141b2532968e9a658e898b3b4a95e;
    5'b01100 : xpb = 1024'h51b1a9c0286517678f585492bd6aeb2cb2b8837657b7d99a07bef1b797cfae37096239bc0c89571d458dbcae4ab280e2fbe86e236e66aa6270c778bc6d9523e1ead69ffba36dc50f8d33b7fcee6408db615532c8abdfcfb67e3f4425b4e1302f277ebce64b183c281278ba9ae79920c1616c53b60efa7f1be1acd10206a14db4;
    5'b01101 : xpb = 1024'h1d9c0b7395c8c7c2979dde5747c066fff1208d5a97df4b945e6ff2bfa8cac30e49123f6374dd498580e4cca52fccb0b26f886a0456b39dd169f85857631b6aa4424e1bc10bdbebb9d2c4b11bcf4dc832ad6ff9268b5b12002195ae7ff09068ad05c6c696411743a6e71827dd7da0816e649765b9cacb954e1d00b96b598df20a;
    5'b01110 : xpb = 1024'h9a33b27cc51aace66ae8dff2e2702a24a0fe9a6fad7e5e0632fdad1d6cc884ed8c0ac283a757ba7c5b9a1be2f844f14c47428dcb61b3618c13c87750937426180e14cc3523db0fa92aefacdd49134bbaed8fb91cf75c815a7a78aad4e66a43bd1316626fe7df43b342777bff0b780844b69c569fd6e808b09ec41cd9355cfccb;
    5'b01111 : xpb = 1024'h661e1430327e5d41732e69b76cc5a5f7df66a453eda5d00089aeae257dc399c4cbbac82b0fabace496f12bd9dd5f211bbae289ac4a0054fb0cf956eb88fa6cda658c47fa8c4936537080a5fc29fd0b1239aa7f7ad6d7c3a41dcf152f22197c3af15e6c1fddde4b321716e941a17f68f1b9c768a392b91ee2da1805428849a121;
    5'b10000 : xpb = 1024'h320875e39fe20d9c7b73f37bf71b21cb1dceae382dcd41fae05faf2d8ebeae9c0b6acdd277ff9f4cd2483bd0c27950eb2e82858d324d486a062a36867e80b39cbd03c3bff4b75cfdb6119f1b0ae6ca6985c545d8b65305edc1257f895dc8b4b8cfa675cfd3dd52b0ebb656843786c99ebcf27aa74e8a3515156bedabdb364577;
    5'b10001 : xpb = 1024'haea01ceccf33f2c04ebef51791cae4efcdacbb4d436c546cb4ed698b52bc707b4e6350f2aa7a1043acfd8b0e8af19185063ca9543d4d0c24affa557faed96f1088ca74340cb680ed0e3c9adc84ac4df1c5e505cf225475481a087bde53a28fc8dcf611a97aa552bd4715aaa5c55e50750ef76b8d5aa6a877972f5119b7055038;
    5'b10010 : xpb = 1024'h7a8a7ea03c97a31b57047edc1c2060c30c14c5318393c6670b9e6a9363b785528e13569a12ce02abe8549b05700bc15479dca5352599ff93a92b351aa45fb5d2e041eff97524a79753cd93fb65960d4911ffcc2d01cfb791bd5ee6388f51c846bb3e1b5970a45a3c1bb517e85b65b12212227d911677bea9d283398309f1f48e;
    5'b10011 : xpb = 1024'h4674e053a9fb53765f4a08a0a675dc964a7ccf15c3bb3861624f6b9b74b29a29cdc35c417b21f51423abaafc5525f123ed7ca1160de6f302a25c14b599e5fc9537b96bbedd92ce41995e8d1a467fcca05e1a928ae14af9db60b55092cb0100c49986250966a361baf054852af16d11cf154d8f94d248d4dc0dd721ec5cde98e4;
    5'b10100 : xpb = 1024'h125f4207175f03d1678f926530cb586988e4d8fa03e2aa5bb9006ca385adaf010d7361e8e375e77c5f02baf33a4020f3611c9cf6f633e6719b8cf4508f6c43578f30e7844600f4ebdeef863927698bf7aa3558e8c0c63c25040bbaed06b0394277ce2eb95ca26939c4f3f26d8774727c1878a1988e19eb0e492b0a55afcb3d3a;
    5'b10101 : xpb = 1024'h8ef6e91046b0e8f53ada9400cb7b1b8e38c2e60f1981bccd8d8e270149ab70e0506be50915f0587339b80a3102b8618d38d6c0be0133aa2c455d1349bfc4fecb5af797f85e0018db371a81faa12f0f7fea5518df2cc7ab7f5ceeb741fc8a1452851dca93036a69462053468f154bf9526a7d927e9a365e70caee6dc38b9a47fb;
    5'b10110 : xpb = 1024'h5ae14ac3b414995043201dc555d09761772aeff359a92ec7e43f28095aa685b7901beab07e444adb750f1a27e7d2915cac76bc9ee9809d9b3e8df2e4b54b458db26f13bdc66e3f857cab7b198218ced7366fdf3d0c42edc90045219c38394cd06365d442f96970c4f4f2b3d1ab5359ff6da8a482560774a30642562cde86ec51;
    5'b10111 : xpb = 1024'h26cbac77217849ab4b65a789e0261334b592f9d799d0a0c23af029116ba19a8ecfcbf057e6983d43b0662a1eccecc12c2016b87fd1cd910a37bed27faad18c5009e68f832edc662fc23c743863028e2e828aa59aebbe3012a39b8bf673e8854e41adddf2ef687843c9922114415abaac70d3b68611d88ad541963e96317390a7;
    5'b11000 : xpb = 1024'ha363538050ca2ecf1eb0a9257ad5d659657106ecaf6fb3340f7de36f2f9f5c6e12c473781912ae3a8b1b795c956501c5f7d0dc46dccd54c4e18ef178db2a47c3d5ad3ff746db8a1f1a676ff9dcc811b6c2aa659157bf9f6cfc7e884b69c2605e4efd79cc9630785024f17535cf324182c2d8a76c1df4fe37c359a2040d429b68;
    5'b11001 : xpb = 1024'h6f4db533be2ddf2a26f632ea052b522ca3d910d0ef97252e662ee477409a71455274791f8166a0a2c67289537a7f31956b70d827c51a4833dabfd113d0b08e862d24bbbcaf49b0c95ff86918bdb1d10e0ec52bef373ae1b69fd4f2a5a57198dc2d45837c8c2f7fcef990e2786539a22fc603b96fd9c61469fead8a6d602f3fbe;
    5'b11010 : xpb = 1024'h3b3816e72b918f852f3bbcae8f80cdffe2411ab52fbe9728bcdfe57f5195861c92247ec6e9ba930b01c9994a5f996164df10d408ad673ba2d3f0b0aec636d548849c378217b7d773a58962379e9b90655adff24d16b62400432b5cffe120d15a0b8d8d2c822e874dce304fbafb4102dcc92ecb7395972a9c3a0172d6b31be414;
    5'b11011 : xpb = 1024'h722789a98f53fe03781467319d649d320a924996fe609231390e68762909af3d1d4846e520e85733d20a94144b3913452b0cfe995b42f11cd219049bbbd1c0adc13b3478025fe1deb1a5b567f854fbca6fab8aaf6316649e681c75a1cd009d7e9d596dc782d8ecca2cfbcfd91486389cc59dd77516840ce75555b400608886a;
    5'b11100 : xpb = 1024'h83ba1fa3c84725040acc480eb4860cf7d08731ae85851b94e81ea0e5268e5cd314cd078e8488f66a17d5f87f0d2bd1ce2a6af3b0a0b3f2cc76f1af42ec15d77ea7da63bb9825220d43455717f94ad344e71a78a16232d5a43f64c3af12a9e4e7f72532b61ef58ed8fe2f111f1f1fea601e5ece5d5d84b430f718beade1d7932b;
    5'b11101 : xpb = 1024'h4fa4815735aad55f1311d1d33edb88cb0eef3b92c5ac8d8f3ecfa1ed378971aa547d0d35ecdce8d2532d0875f246019d9e0aef918900e63b70228edde19c1e40ff51df81009348b788d65036da34929c33353eff41ae17ede2bb2e094e591d65d56d3c6614f49657d2ce7e61b5274b0d2189e0611955ca63326ca71734c43781;
    5'b11110 : xpb = 1024'h1b8ee30aa30e85ba1b575b97c931049e4d57457705d3ff899580a2f548848681942d12dd5530db3a8e84186cd760316d11aaeb72714dd9aa69536e78d722650356c95b4669016f61ce674955bb1e51f37f50055d21295a37861198638a0855e3b3b546160af39dd6a76deba44b2eabba24b4f264d526e0956dc08f8087b0dbd7;
    5'b11111 : xpb = 1024'h98268a13d2606addeea25d3363e0c7c2fd35528c1b7311fb6a0e5d530c824860d72595fd87ab4c31693967aa9fd87206e9650f397c4d9d6513238d72077b207722900bba810093512692451734e3d57bbf6fc5538d2ac991def494b87fe230f3c104e1efb1bb9de302cd3fc5d906329076b9e34ae14353f7ef83f2ee637fe698;
    endcase
end

endmodule

module xpb_5_710
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h3bb79598b40ff58f855bd7e28df934378d2612b5c2ff34f13f7e357268c41a6465e77615fe5a6181278c305e45838930ad471efe59b5fa5aee14eccfcd528a752ef3c7e6cedf85946991e82056d0b4004b9863ddd095abb93bd088787d098a49547784d5bf0817053627ddce7395f9871fdfff26fd05135256d621eaecb632b3;
    5'b00010 : xpb = 1024'h776f2b31681feb1f0ab7afc51bf2686f1a4c256b85fe69e27efc6ae4d18834c8cbceec2bfcb4c3024f1860bc8b0712615a8e3dfcb36bf4b5dc29d99f9aa514ea5de78fcd9dbf0b28d323d040ada168009730c7bba12b577277a110f0fa131492a8ef09ab7e102e0a6c4fbb9ce72bf30e3fbffe4dfa0a26a4adac43d5d96c6566;
    5'b00011 : xpb = 1024'h2797b745a41abe5c50e0fd09991555535fc34f07385fe5c409de7018749a2252e6de4c930e8a5f4d74651d3ed2c8ac7a3bb3514ea6f1ec5199f87112d252aae188c2305bd0d93782a1bb5be6b9657cfeec43200e53ad61afde5076ebcf1fc49ce5efc578c4f4c821bb7b28c62f1c66c10c61e92a6c3dcc6be12eabc3d4031ae;
    5'b00100 : xpb = 1024'h3e31110d0e51a1754a69e7b3278a898cc32247a63685334d801c1c73f00dbc8994555adf2f430775fed2823232b013f8510254134425192007b473e0fa77b523477feaec8bed190c93ad9ddec2670bd03a5c95deb5d081d439b58fe739fb869322d6812d4b57638751df905ad687bff330a61db9a3c8f01914e90ca729f66461;
    5'b00101 : xpb = 1024'h79e8a6a5c2619704cfc5bf95b583bdc450485a5bf984683ebf9a51e658d1d6edfa3cd0f52d9d68f7265eb29078339d28fe4973119ddb137af5c960b0c7ca3f987673b2d35acc9ea0fd3f85ff1937bfd085f4f9bc86662d8d7586185fb70510dc774e06030a5f7a8c88076e294a1db97a50861ce0a0ce036b6bbf2e9216ac9714;
    5'b00110 : xpb = 1024'h4f2f6e8b48357cb8a1c1fa13322aaaa6bf869e0e70bfcb8813bce030e93444a5cdbc99261d14be9ae8ca3a7da59158f47766a29d4de3d8a333f0e225a4a555c3118460b7a1b26f054376b7cd72caf9fdd886401ca75ac35fbca0edd79e3f8939cbdf8af189e9904376f6518c5e38cd8218c3d254d87b98d7c25d5787a80635c;
    5'b00111 : xpb = 1024'h40aa8c8168934d5b0f77f783c11bdee1f91e7c96aa0b31a9c0ba037577575eaec2c33fa8602bad6ad618d4061fdc9ebff4bd89282e9437e52153faf2279cdfd1600c0df248faac84bdc9539d2dfd63a02920c7df9b0b57ef379a9755f6ed82dcf1357d84d7a6b0096d9742e73979865f416c3c4c4a8cccdfd2fbf7636736960f;
    5'b01000 : xpb = 1024'h7c62221a1ca342ea94d3cf664f15131986448f4c6d0a669b003838e7e01b791328aab5be5e860eebfda50464656027f0a204a826884a32400f68e7c1f4ef6a468effd5d917da3219275b3bbd84ce17a074b92bbd6ba103a8736b1fce73f70d2645ad025a96aec70ea3bf20b5ad0f7fe6614c3b734791e03229d2194e53ecc8c2;
    5'b01001 : xpb = 1024'h76c725d0ec503b14f2a2f71ccb3ffffa1f49ed15a91fb14c1d9b50495dce66f8b49ae5b92b9f1de85d2f57bc785a056eb319f3ebf4d5c4f4cde9533876f800a49a469113728ba687e53213b42c3076fcc4c9602afb08250f9af164c36d5f4dd6b1cf506a4ede586532717a528d5534432525bb7f44b96543a38c034b7c0950a;
    5'b01010 : xpb = 1024'h432407f5c2d4f940d48607545aad34372f1ab1871d9130060157ea76fea100d3f13124719114535fad5f25da0d0929879878be3d190356aa3af3820354c20a7f789830f806083ffce7e5095b9993bb7017e4f9e080462e0a357f9ec4b3df7f26bf9479dc63f5fc8b894ef5739c6b4ccb52325adef150a9a6910ee21fa476c7bd;
    5'b01011 : xpb = 1024'h7edb9d8e76e4eed059e1df36e8a6686ebc40c43ce09064f740d61fe967651b3857189a878f6eb4e0d4eb5638528cb2b845bfdd3b72b9510529086ed3221494f4a78bf8ded4e7c5915176f17bf0646f70637d5dbe50dbd9c37150273d30e90970140bfeb222fe1390bf76d3421001465272125a05ee55bcf8e7e5040a912cfa70;
    5'b01100 : xpb = 1024'h9e5edd16906af9714383f4266455554d7f0d3c1ce17f97102779c061d268894b9b79324c3a297d35d19474fb4b22b1e8eecd453a9bc7b14667e1c44b494aab862308c16f4364de0a86ed6f9ae595f3fbb10c80394eb586bf7941dbaf3c7f127397bf15e313d32086edeca318bc719b043187a4a9b0f731af84baaf0f500c6b8;
    5'b01101 : xpb = 1024'h459d836a1d16a52699941724f43e898c6516e67791172e6241f5d17885eaa2f91f9f093ac1fcf95484a577adfa35b44f3c33f3520372756f5493091481e7352d912453fdc315d3751200bf1a052a134006a92be1658104253364a63370d17b708df37633f045490da506a7ffff5d133762f879719814866d4f21ccdbe1b6f96b;
    5'b01110 : xpb = 1024'h81551902d1269ab61eefef078237bdc3f23cf92d54166353817406eaeeaebd5d85867f50c0575ad5ac31a80c3fb93d7fe97b12505d286fca42a7f5e44f39bfa2c0181be491f559097b92a73a5bfac74052418fbf3616afde6f352eabeddb05b9e26afb09af4d6012db2e85ce72f30cbe82d87898951999bfa5f7eec6ce6d2c1e;
    5'b01111 : xpb = 1024'hc5f6945c3485b7cd9464f12ffd6aaaa0ded08b2419df7cd43158307a4702ab9e82577edf48b3dc8345f9923a1deb5e632a80968942b99d9801da355e1b9d5667abcaf1cb143e158d28a8cb819efb70fa9d4fa047a262e86f5792529b0b9ed7107daedb5bd8c7e8a8a967cbdeeb8e01c53de98dd41d34fe1b65e95ad3240f866;
    5'b10000 : xpb = 1024'h4816fede7758510c5ea226f58dcfdee19b131b68049d2cbe8293b87a0d34451e4e0cee03f2e59f495bebc981e7623f16dfef2866ede194346e329025af0c5fdba9b07703802366ed3c1c74d870c06b0ff56d5de24abbda403149ada22dc377ba5c52728b7c94958fc0be5a8c624ed9a373be98043ed863340d34b7981ef72b19;
    5'b10001 : xpb = 1024'h83ce94772b68469be3fdfed81bc9131928392e1dc79c61afc211edec75f85f82b3f46419f14000ca8377f9e02ce5c8478d36476547978e8f5c477cf57c5eea50d8a43eea4f02ec81a5ae5cf8c7911f104105c1c01b5185f96d1a361aaacd0203b0c9f7613b9cac94f6e6385ad5e4d32a939e972b3bdd7686640ad9830bad5dcc;
    5'b10010 : xpb = 1024'hed8e4ba1d8a07629e545ee39967ffff43e93da2b523f62983b36a092bb9ccdf16935cb72573e3bd0ba5eaf78f0b40add6633e7d7e9ab89e99bd2a670edf00149348d2226e5174d0fca6427685860edf98992c055f6104a1f35e2c986dabe9bad639ea0d49dbcb0ca64e2f4a51aaa68864a4b76fe8972ca8747180696f812a14;
    5'b10011 : xpb = 1024'h4a907a52d199fcf223b036c627613436d10f505878232b1ac3319f7b947de7437c7ad2cd23ce453e33321b55d48ec9de83aa5d7bd850b2f987d21736dc318a89c23c9a093d30fa6566382a96dc56c2dfe4318fe32ff6b05b2f2eb510eab574042ab16ee308e3e211dc760d18c540a00f8484b696e59c3ffacb47a2545c375cc7;
    5'b10100 : xpb = 1024'h86480feb85a9f281a90c0ea8b55a686e5e35630e3b22600c02afd4edfd4201a7e26248e32228a6bf5abe4bb41a12530f30f17c7a3206ad5475e70406a98414fef13061f00c107ff9cfca12b7332776e02fc9f3c1008c5c146aff3d8967befe4d7f28f3b8c7ebf917129deae738d69996a464b5bde2a1534d221dc43f48ed8f7a;
    5'b10101 : xpb = 1024'h1152602e77cbb34863626eb432f9555479e5729328a9f485c451510ab3036f0445014180565c89b1e2ec3ccb7c37cb757a1e73926909d763b35cb1783c042ac2abd4f5282b5f084926c1f834f11c66af875d5e06449bdabcf14334072a9de604a498e664d62b178ec205e1d6b49c6cf4756ad6028f5b096f32846b25acc15bc2;
    5'b10110 : xpb = 1024'h4d09f5c72bdba8d7e8be4696c0f2898c070b8548eba9297703cf867d1bc78968aae8b79654b6eb330a786d29c1bb54a627659290c2bfd1bea1719e480956b537dac8bd0efa3e8ddd9053e05547ed1aafd2f5c1e4153186762d13bc7fa7a7704df9106b3a95332e93f82dbfa52832667b954ad5298c601cc1895a8d1099778e75;
    5'b10111 : xpb = 1024'h88c18b5fdfeb9e676e1a1e794eebbdc3943197feaea85e68434dbbef848ba3cd10d02dac53114cb432049d88073eddd6d4acb18f1c75cc198f868b17d6a93fad09bc84f5c91e1371f9e5c8759ebdceb01e8e25c1e5c7322f68e444f824b0fa974d87f010543b45992e559d739bc86002b52ad45089653013e030aefb862dc128;
    5'b11000 : xpb = 1024'h13cbdba2d20d5f2e28707e84cc8aaaa9afe1a7839c2ff2e204ef380c3a4d1129736f264987452fa6ba328e9f6964563d1dd9a8a75378f628ccfc388969295570c461182de86c9bc150ddadf35cb2be7f7621900729d6b0d7ef283b75e78fe24e72f7e2bc627a6410ddbd9463178e33608630f495361ee635f09755e1ea018d70;
    5'b11001 : xpb = 1024'h4f83713b861d54bdadcc56675a83dee13d07ba395f2f27d3446d6d7ea3112b8dd9569c5f859f9127e1bebefdaee7df6dcb20c7a5ad2ef083bb112559367bdfe5f354e014b74c2155ba6f9613b383727fc1b9f3e4fa6c5c912af8c3ee64996c97c76f679221827b1613e572318b242ce7a610f3bc3323f988476d77ccd6b7c023;
    5'b11010 : xpb = 1024'h8b3b06d43a2d4a4d33282e49e87d1318ca2dccef222e5cc483eba2f10bd545f23f3e127583f9f2a9094aef5bf46b689e7867e6a406e4eadea926122903ce6a5b2248a7fb862ba6ea24017e340a5426800d5257c2cb02084a66c94c66e1a2f6e11be6ec67e08a921b4a0d4ffffeba266ec5f0f2e330290cda9e4399b7c36df2d6;
    5'b11011 : xpb = 1024'h164557172c4f0b13ed7e8e55661bfffee5dddc740fb5f13e458d1f0dc196b34ea1dd0b12b82dd59b9178e0735690e104c194ddbc3de814ede69bbf9a964e801edced3b33a57a2f397af963b1c849164f64e5c2080f1186f2ed0d42e4a481de984156df13eec9b092f97546ef7a7ff9cc96f71327dce2c2fcaeaa409e2741bf1e;
    5'b11100 : xpb = 1024'h51fcecafe05f00a372da6637f41534367303ef29d2b5262f850b54802a5acdb307c48128b688371cb90510d19c146a356edbfcba979e0f48d4b0ac6a63a10a940be1031a7459b4cde48b4bd21f19ca4fb07e25e5dfa732ac28ddcb5d218b68e195ce63e9add1c7982f9d24bdee15f353b6d7124ed9e7d64f0580628913f7f1d1;
    5'b11101 : xpb = 1024'h8db48248946ef632f8363e1a820e686e002a01df95b45b20c48989f2931ee8176dabf73eb4e2989de091412fe197f3661c231bb8f15409a3c2c5993a30f395093ad4cb0143393a624e1d33f275ea7e4ffc1689c3b03cde6564ae53d59e94f32aea45e8bf6cd9de9d65c5028c61abecdad6b71175d6ece9a15c56847400ae2484;
    5'b11110 : xpb = 1024'h18bed28b8690b6f9b28c9e25ffad55541bda1164833bef9a862b060f48e05573d04aefdbe9167b9068bf324743bd6bcc655012d1285733b3003b46abc373aaccf5795e396287c2b1a515197033df6e1f53a9f408f44c5d0deaf24a536173dae20fb5db6b7b18fd15152cf97bdd71c038a7bd31ba83a69fc36cbd2b5a6481f0cc;
    5'b11111 : xpb = 1024'h547668243aa0ac8937e876088da6898ba900241a463b248bc5a93b81b1a46fd8363265f1e770dd11904b62a58940f4fd129731cf820d2e0dee50337b90c63542246d2620316748460ea701908ab0221f9f4257e6c4e208c726c2d2cbde7d652b642d60413a21141a4b54d74a5107b9bfc79d30e180abb315c3934d455138237f;
    endcase
end

endmodule

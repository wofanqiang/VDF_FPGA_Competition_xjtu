module xpb_5_620
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h3d929c25b044468c5c149d590a8c1c64c0ab15ebae3df57826857c8577e374bc5efa553160354758e117e8d97a1982e14525ad0a2cc5e3bbff41e2a58e82c711bda9d3577438e26cc96cf0c6c533b0408c7d276c28deaa8ffb23e3d95a2a2b1a003a0d944d37fb28f1d8b7077030344b4239f4f3add9ac68faebf8238a863b62;
    5'b00010 : xpb = 1024'h7b25384b60888d18b8293ab2151838c981562bd75c7beaf04d0af90aefc6e978bdf4aa62c06a8eb1c22fd1b2f43305c28a4b5a14598bc777fe83c54b1d058e237b53a6aee871c4d992d9e18d8a67608118fa4ed851bd551ff647c7b2b454563400741b289a6ff651e3b16e0ee06068968473e9e75bb358d1f5d7f047150c76c4;
    5'b00011 : xpb = 1024'h80a8f1b4ede9edc493860340f4a0ddcd08b3e9235423ff0f5b3bc3ab4a7b12d19a6821b5679577c03e97b458aee77d96b56df38639edae84d26689270b5e083c4ae4557ad19aa0149accfb1b6bf4c90b1727cabee15d29f3bdf19915453debbd1a6969336def8ed4eca3e3758c076b877d3fff8b941a80aaa546d6616b04bbb;
    5'b00100 : xpb = 1024'h459d2b40ff22e568a54cfd8d19d62a419136547de38035691c3938c02c8b25e978a0d74cb6ae9ed4e501641f0507fabab07c8c429064bea44c684b37ff38a795825818af21528c6e1319c0787bf2fcd13defa41816f47d2f3702fd6aae7e09d5d1e0a4278416f41640a2f53ec8f0ab03ba0df4ec671b5473a5406589a136871d;
    5'b00101 : xpb = 1024'h832fc766af672bf501619ae6246246a651e16a6991be2ae142beb545a46e9aa5d79b2c7e16e3e62dc6194cf87f217d9bf5a2394cbd2aa2604baa2ddd8dbb6ea74001ec06958b6edadc86b13f4126ad11ca6ccb843fd327bf3226e14408a834efd21ab1bbd14eef3f327bac463920df4efc47e9e014f500dca02c5dad2bbcc27f;
    5'b00110 : xpb = 1024'h10151e369dbd3db89270c0681e941bb9a1167d246a847fe1eb677875694f625a334d0436acf2aef807d2f68b15dcefb2d6adbe70c73db5d09a4cd124e16bc107895c8aaf5a33540293599f636d7e992162e4f957dc2ba53e77be3322a8a7bd77a34d2d266dbdf1da9d947c6eb180ed70efa7fff17283501554a8dacc2d609776;
    5'b00111 : xpb = 1024'h4da7ba5c4e018444ee855dc12920381e61c1931018c2755a11ecf4fae132d716924759680d27f650e8eadf648ff672941bd36b7af403998c998eb3ca6fee881947065e06ce6c366f5cc6902a32b24961ef6220c4050a4fce72e216fc02d1e891a3873ababaf5ed038f6d337621b121bc31e1f4e5205cfc7e4f94d2efb7e6d2d8;
    5'b01000 : xpb = 1024'h8b3a5681fe45cad14a99fb1a33ac5483226ca8fbc7006ad23872718059164bd2f141ae996d5d3da9ca02c83e0a0ff57560f9188520c97d4898d0966ffe714f2b04b0315e42a518dc263380f0f7e5f9a27bdf48302de8fa5e6e05fad55cfc13aba3c1484f082de82c8145ea7d91e15607741be9d8ce36a8e74a80cb13426d0e3a;
    5'b01001 : xpb = 1024'h181fad51ec9bdc94dba9209c2dde299671a1bbb69fc6bfd2e11b34b01df713874cf38652036c06740bbc71d0a0cb678c42049da92adc90b8e77339b75221a18b4e0ad007074cfe03dd066f15243de5b214577603ca4177ddb39d4cb3fcfb9c3374f3c3b9a49ceac7ec5ebaa60a416429677bffea2bc4f81ffefd48324410e331;
    5'b01010 : xpb = 1024'h55b249779ce0232137bdbdf5386a45fb324cd1a24e04b54b07a0b13595da8843abeddb8363a14dccecd45aaa1ae4ea6d872a4ab357a27474e6b51c5ce0a4689d0bb4a35e7b85e070a6735fdbe97195f2a0d49d6ff320226daec1308d5725c74d752dd14df1d4e5f0de3771ad7a719874a9b5f4ddd99ea488f9e94055ce971e93;
    5'b01011 : xpb = 1024'h9344e59d4d2469ad93d25b4e42f6625ff2f7e78dfc42aac32e262dbb0dbdfd000ae830b4c3d69525cdec438394fe6d4ecc4ff7bd84685830e5f6ff026f272faec95e76b5efbec2dd6fe050a2aea546332d51c4dc1bfeccfda9e51466b14ff2677567dee23f0ce119d01028b4eaa1ccbfebefe9d1877850f1f4d53879591d59f5;
    5'b01100 : xpb = 1024'h202a3c6d3b7a7b7124e180d03d283773422cfa48d508ffc3d6cef0ead29ec4b4669a086d59e55df00fa5ed162bb9df65ad5b7ce18e7b6ba13499a249c2d7820f12b9155eb466a80526b33ec6dafd3242c5c9f2afb8574a7cef7c6645514f7aef469a5a4cdb7be3b53b28f8dd6301dae1df4fffe2e506a02aa951b5985ac12eec;
    5'b01101 : xpb = 1024'h5dbcd892ebbec1fd80f61e2947b453d802d810348346f53bfd546d704a823970c5945d9eba1aa548f0bdd5efa5d36246f28129ebbb414f5d33db84ef515a4920d062e8b6289f8a71f0202f8da030e28352471a1be135f50ceaa04a1eab79a60946d467e128b3dede2d01afe4d3320f2d2189f4d692e04c93a43dadbbe5476a4e;
    5'b01110 : xpb = 1024'h9b4f74b89c030889dd0abb825240703cc38326203184eab423d9e9f5c265ae2d248eb2d01a4feca1d1d5bec91fece52837a6d6f5e8073319331d6794dfdd10328e0cbc0d9cd86cdeb98d2054656492c3dec441880a149f9ce5c42df805a3d123470e757575ebda071eda66ec4362437863c3e9ca40b9f8fc9f29a5df6fcda5b0;
    5'b01111 : xpb = 1024'h2834cb888a591a4d6e19e1044c72455012b838db0a4b3fb4cc82ad25874675e180408a88b05eb56c138f685bb6a8573f18b25c19f21a468981c00adc338d6292d7675ab66180520670600e7891bc7ed3773c6f5ba66d1d1c2b5b7fd6a5a359ab1840f0e0125adca289f33714bbc2519a5723ffdb9e48483553a622fe71717aa7;
    5'b10000 : xpb = 1024'h65c767ae3a9d60d9ca2e7e5d56fe61b4d3634ec6b889352cf30829aaff29ea9ddf3adfba1093fcc4f4a7513530c1da205dd809241ee02a458101ed81c21029a495112e0dd5b9347339ccff3f56f02f1403b996c7cf4bc7ac267f63afffcd84c5187afe745f92d7cb7bcbee1c2bf285e5995df4cf4c21f49e4e921b21fbf7b609;
    5'b10001 : xpb = 1024'ha35a03d3eae1a76626431bb6618a7e19940e64b266c72aa5198da630770d5f5a3e3534eb70c9441dd5bf3a0eaadb5d01a2fdb62e4ba60e018043d0275092f0b652bb016549f216e00339f0061c23df549036be33f82a723c21a3478959f7afdf18b50c08accad2f46da4a5239c22ba30db97e9c2f9fba107497e1345867df16b;
    5'b10010 : xpb = 1024'h303f5aa3d937b929b75241385bbc532ce343776d3f8d7fa5c23669603bee270e99e70ca406d80ce81778e3a14196cf1884093b5255b92171cee6736ea44343169c15a00e0e99fc07ba0cde2a487bcb6428aeec079482efbb673a9967f9f73866e9e787734939d58fd8bd754c1482c852cef7ffd45789f03ffdfa90648821c662;
    5'b10011 : xpb = 1024'h6dd1f6c9897bffb61366de9166486f91a3ee8d58edcb751de8bbe5e5b3d19bcaf8e161d5670d5440f890cc7abbb051f9c92ee85c827f052dce28561432c60a2859bf736582d2de748379cef10daf7ba4b52c1373bd619a4b625e7d4154216380ea2195079671d0b8ca962c5384b2fc9e1131f4c805639ca8f8e6888812a801c4;
    5'b10100 : xpb = 1024'hab6492ef39c046426f7b7bea70d48bf66499a3449c096a960f41626b2bb5108757dbb706c7429b99d9a8b55435c9d4db0e549566af44e8e9cd6a38b9c148d13a176946bcf70bc0e14ce6bfb7d2e32be541a93adfe64044db5d82611aae4b8e9aea5ba29be3a9cbe1bc6ee35af4e330e9536be9bbb33d4911f3d280ab9d2e3d26;
    5'b10101 : xpb = 1024'h3849e9bf28165806008aa16c6b066109b3ceb5ff74cfbf96b7ea259af095d83bb38d8ebf5d5164641b625ee6cc8546f1ef601a8ab957fc5a1c0cdc0114f9239a60c3e565bbb3a60903b9addbff3b17f4da2168b38298c25aa319b2f94e4b1722bb8e1e068018ce7d2787b3836d433f0b46cbffcd10cb984aa84efdca9ed2121d;
    5'b10110 : xpb = 1024'h75dc85e4d85a9e925c9f3ec575927d6e7479cbeb230db50ede6fa22068794cf81287e3f0bd86abbcfc7a47c0469ec9d33485c794e61de0161b4ebea6a37beaac1e6db8bd2fec8875cd269ea2c46ec835669e901fab776cea9e3d96d2a875423cbbc82b9acd50c9a619606a8add7373568905f4c0bea544b3a33af5ee29584d7f;
    5'b10111 : xpb = 1024'h2c1dcb4c6b0b055edae64476fc45281c3aedea5fbd40a0f871865502d5a14ac6e39bba9539574873e33f152dd5a3bea15914cb8f030f38669f161edf72c3d0c67c85765f4946d9d83f98cc6f0c6b444ff16bdf347cfea69e3d4e8b14874cac48cfaa70569bfcc4184793ab355d381787c660ad21c3393ec57b7730d2afc2276;
    5'b11000 : xpb = 1024'h405478da76f4f6e249c301a07a506ee68459f491aa11ff87ad9de1d5a53d8968cd3410dab3cabbe01f4bda2c5773becb5ab6f9c31cf6d7426933449385af041e25722abd68cd500a4d667d8db5fa64858b93e55f70ae94f9def8cc8aa29ef5de8d34b499b6f7c76a7651f1bac603b5c3be9fffc5ca0d405552a36b30b5825dd8;
    5'b11001 : xpb = 1024'h7de7150027393d6ea5d79ef984dc8b4b45050a7d584ff4ffd4235e5b1d20fe252c2e660c140003390063c305d18d41ac9fdca6cd49bcbafe687527391431cb2fe31bfe14dd06327716d36e547b2e14c618110ccb998d3f89da1cb063fcc920f88d6ec22e042fc293682aa8c23633ea0f00d9f4b977e6ecbe4d8f63544008993a;
    5'b11010 : xpb = 1024'hacc6bd0158f4f3236e6c47b7f0e605e943a1d3831164a007ccc218ae201c5d987e03dc4aa0ecc03421d6c986848b3c380e82bf153cfce6eb717ca8067e21d902c769cbda1ae179ecda65c78a78600d5b0893a9f35e5bd091fb402429cc8a9805ea13d98a09ec52ed34378eaae93f830f43a0acad5753bf7020be07341ac6e31;
    5'b11011 : xpb = 1024'h485f07f5c5d395be92fb61d4899a7cc354e53323df543f78a3519e1059e53a95e6da92f60a44135c23355571e26236a4c60dd8fb8095b22ab659ad25f664e4a1ea20701515e6fa0b97134d3f6cb9b1163d06620b5ec467991ad7e61bf6f2d49a5edb4b2cedd6c057c51c2ff21ec42c7c3673ffbe834ee85ffcf7d896cc32a993;
    5'b11100 : xpb = 1024'h85f1a41b7617dc4aef0fff2d942699281590490f8d9234f0c9d71a95d1c8af5245d4e8276a795ab5044d3e4b5c7bb9860b338605ad5b95e6b59b8fcb84e7abb3a7ca436c8a1fdc7860803e0631ed6156c983897787a3122915fbc9f5511cffb45f1558c13b0ebb80b6f4e6f98ef460c778adf4b2312894c8f7e3d0ba56b8e4f5;
    5'b11101 : xpb = 1024'h12d6faeb646dee0e801f24af8e586e3b64c55bca665889f1727fddc596a97706a186bfe00088237f4606e7ddf3372b9cec3f0b29b76ea957043e3312d897fe13f124e2154ec7c1a017532c2a5e454d6661fbb74b23fb8fa85b931bd3f11c883c3047d42bd77dbe1c220db72207546ee96c0e0ac38eb6e401ac604dd9585cb9ec;
    5'b11110 : xpb = 1024'h5069971114b2349adc33c20898e48aa0257071b614967f6999055a4b0e8cebc30081151160bd6ad8271ed0b76d50ae7e3164b833e4348d13038015b8671ac525aeceb56cc300a40ce0c01cf12378fda6ee78deb74cda3a3856b6ffad4b46b3563081e1c024b5b94513e66e297784a334ae47ffb73c90906aa74c45fce2e2f54e;
    5'b11111 : xpb = 1024'h8dfc3336c4f67b2738485f61a370a704e61b87a1c2d474e1bf8ad6d08670607f5f7b6a42c0f2b2310836b990e76a315f768a653e10fa70cf02c1f85df59d8c376c7888c437398679aa2d0db7e8acade77af6062375b8e4c851dae386a570de7030bbef5471edb46e05bf2530e7b4d77ff081f4aaea6a3cd3a2383e206d6930b0;
    endcase
end

endmodule

module xpb_5_480
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h5263a618b6f620c1a13a4b598a7e44dd8369b75c98eeb87a0cf29476b0829eaadced65aa925c176c87cc80266eedcd0c50f84215f60aa986cb2d9274cc11ad6ae59d34fda5e4f6ff84fae01c86caa977a0452096cc44c3ee60d7957940277ca09cc68cd5ff88a76022f60c0cbc04e6711f9296d8ba06332fa4033cf521360841;
    5'b00010 : xpb = 1024'ha4c74c316dec4183427496b314fc89bb06d36eb931dd70f419e528ed61053d55b9dacb5524b82ed90f99004cdddb9a18a1f0842bec15530d965b24e998235ad5cb3a69fb4bc9edff09f5c0390d9552ef408a412d988987dcc1af2af2804ef941398d19abff114ec045ec18197809cce23f252db1740c665f480679ea426c1082;
    5'b00011 : xpb = 1024'h467dacf462f42d7c18a96a358f20874718c722e4f55488f6a8fb040e5e852ef8937fb386ecedc7b6f807412c696b565a8ece9e5bbf6d2c48b0e978002962938f3c886a4a421de7b97c569db2fb843835ecca682bd8481eba6cfa2e71064bd34fa74c14584dd0fd92e2223d473c3e8d2a0fdde5a7ddc73c5ea59a3bdadabfb258;
    5'b00100 : xpb = 1024'h98e1530d19ea4e3db9e3b58f199ecc249c30da418e434170b5ed98850f07cda3706d19317f49df237fd3c152d8592366dfc6e071b577d5cf7c170a74f57440fa22259f47e802deb901517dcf824ee1ad8d0f88c2a48ce2a8cdd1c3ea46734ff04412a12e4d59a4f305184953f843739b2f707c8097cd6f8e499d78cffbf5ba99;
    5'b00101 : xpb = 1024'h3a97b3d00ef23a369018891193c2c9b0ae248e6d51ba5973450373a60c87bf464a120163477f78016842023263e8dfa8cca4faa188cfaf0a96a55d8b86b379b393739f96de56d87373b25b49703dc6f4394fafc0e44b7986791cc768cc7029feb1d19bda9c1953c5a14e6e81bc7833e3002934770188458da7313ac094495c6f;
    5'b00110 : xpb = 1024'h8cfb59e8c5e85af83152d46b1e410e8e318e45c9eaa911ed51f6081cbd0a5df126ff670dd9db8f6df00e8258d2d6acb51d9d3cb77eda589161d2f00052c5271e7910d494843bcf72f8ad3b65f708706bd994d057b0903d74d9f45ce20c97a69f4e9828b09ba1fb25c4447a8e787d1a541fbbcb4fbb8e78bd4b3477b5b57f64b0;
    5'b00111 : xpb = 1024'h2eb1baabbaf046f10787a7ed98650c1a4381f9f5ae2029efe10be33dba8a4f9400a44f3fa211284bd87cc3385e6668f70a7b56e7523231cc7c614316e4045fd7ea5ed4e37a8fc92d6b0e18dfe4f755b285d4f755f04ed452853f6060929480adbc57235cea61a9f8607a9fbc3cb1da9bf074834625494ebca8c839a64dd30686;
    5'b01000 : xpb = 1024'h811560c471e667b2a8c1f34722e350f7c6ebb152470ee269edfe77b46b0cee3edd91b4ea346d3fb86049435ecd5436035b7398fd483cdb53478ed58bb0160d42cffc09e12074c02cf008f8fc6bc1ff2a261a17ecbc939840e616f5d9d2bbfd4e591db032e9ea51588370abc8f8b6c10d10071a1edf4f81ec4ccb769b6f090ec7;
    5'b01001 : xpb = 1024'h22cbc18766ee53ab7ef6c6c99d074e83d8df657e0a85fa6c7d1452d5688cdfe1b7369d1bfca2d89648b7843e58e3f2454851b32d1b94b48e621d28a2415545fc414a0a3016c8b9e76269d67659b0e470d25a3eeafc522f1e9161f95858b8d75cc6dcaadf38aa002b1fa6d0f6bceb8154e0bfd215490a57ebaa5f388c075cb09d;
    5'b01010 : xpb = 1024'h752f67a01de4746d20311223278593615c491cdaa374b2e68a06e74c190f7e8c942402c68efef002d0840464c7d1bf519949f543119f5e152d4abb170d66f36726e73f2dbcadb0e6e764b692e07b8de8729f5f81c896f30cf2398ed198e053fd63a337b53832a78b429cdd0378f067c6005268ee03108b1b4e6275812892b8de;
    5'b01011 : xpb = 1024'h16e5c86312ec6065f665e5a5a1a990ed6e3cd10666ebcae9191cc26d168f702f6dc8eaf8573488e0b8f2454453617b9386280f72e4f7375047d90e2d9ea62c2098353f7cb301aaa159c5940cce6a732f1edf8680085589ea9d8492501edd2e0bd162326186f2565dded302313d25280dd10b20e46ccb611aabf63771c0e65ab4;
    5'b01100 : xpb = 1024'h69496e7bc9e2812797a030ff2c27d5caf1a68862ffda8363260f56e3c7120eda4ab650a2e990a04d40bec56ac24f489fd7205188db01e0d71306a0a26ab7d98b7dd2747a58e6a1a0dec0742955351ca6bf24a716d49a4dd8fe5c27c95f04aaac6e28bf37867afdbe01c90e3df92a0e7ef09db7bd26d1944a4ff97466e21c62f5;
    5'b01101 : xpb = 1024'haffcf3ebeea6d206dd50481a64bd357039a3c8ec3519b65b5253204c492007d245b38d4b1c6392b292d064a4ddf04e1c3fe6bb8ae59ba122d94f3b8fbf71244ef2074c94f3a9b5b512151a3432401ed6b64ce151458e4b6a9a72b47e50184badbe7b9e3d53aac909dff336bbd5ecec6c1566fb3908c6a49ad8d36577a7004cb;
    5'b01110 : xpb = 1024'h5d63755775e08de20f0f4fdb30ca18348703f3eb5c4053dfc217c67b75149f2801489e7f44225097b0f98670bcccd1ee14f6adcea4646398f8c2862dc808bfafd4bda9c6f51f925ad61c31bfc9eeab650ba9eeabe09da8a50a7ec0c12529015b78ae46b9d4c353f0c0f53f787963b537e0e9068c4a929d795190734c9ba60d0c;
    5'b01111 : xpb = 1024'hafc71b702cd6aea3b0499b34bb485d120a6dab47f52f0c59cf0a5af225973dd2de360429d67e680438c606972bba9efa65eeefe49a6f0d1fc3f018a2941a6d1aba5adec49b04895a5b1711dc50b954dcabef0f42ace26c936b56563a65507dfc1574d38fd44bfb50e3eb4b8535689ba9007b9d650498d0a8f593b041bcdc154d;
    5'b10000 : xpb = 1024'h517d7c3321de9a9c867e6eb7356c5a9e1c615f73b8a6245c5e20361323172f75b7daec5b9eb400e221344776b74a5b3c52cd0a146dc6e65ade7e6bb92559a5d42ba8df1391588314cd77ef563ea83a23582f3640eca1037116a159b8eb4d580a8333ce3c230baa23802170b2f99d5bf0d134555b6e53a6a853277232552fb723;
    5'b10001 : xpb = 1024'ha3e1224bd8d4bb5e27b8ba10bfea9f7b9fcb16d05194dcd66b12ca89d399ce2094c852063110184ea900c79d26382848a3c54c2a63d18fe1a9abfe2df16b533f11461411373d7a145272cf72c572e39af87456d7b8e5c75f7778ef322b74d4ab1ffa5b1222945183a3177cbfb5a24261f0c6ec342859d9d7f72aaf277665bf64;
    5'b10010 : xpb = 1024'h4597830ecddca756fded8d933a0e9d07b1becafc150bf4d8fa28a5aad119bfc36e6d3a37f945b12c916f087cb1c7e48a90a3665a3729691cc43a514482aa8bf8829414602d9173cec4d3acecb361c8e1a4b47dd5f8a45e3d22c3f2b0b171aeb98db955be715400563f4da1ed79d702a9c17fa42a9214afd754be71180eb9613a;
    5'b10011 : xpb = 1024'h97fb292784d2c8189f27d8ecc48ce1e535288258adfaad53071b3a21819c5e6e4b5a9fe28ba1c899193b88a320b5b196e19ba8702d3412a38f67e3b94ebc39636831495dd3766ace49ce8d093a2c725944f99e6cc4e9222b839b8829f1992b5a2a7fe29470dca7b66243adfa35dbe91ae1123b034c1ae306f8c1ae0d2fef697b;
    5'b10100 : xpb = 1024'h39b189ea79dab411755cac6f3eb0df71471c36847171c555963115427f1c501124ff881453d7617701a9c982ac456dd8ce79c2a0008bebdea9f636cfdffb721cd97f49acc9ca6488bc2f6a83281b579ff139c56b04a7b9092ee68ba877960568983edd40bf9c5688fe79d327fa10a962b1caf2f9b5d5b90656556ffdc8430b51;
    5'b10101 : xpb = 1024'h8c15300330d0d4d31696f7c8c92f244eca85ede10a607dcfa323a9b92f9eeebc01ecedbee63378e3897649a91b333ae51f7204b5f69695657523c944ac0d1f87bf1c7eaa6faf5b88412a4a9faee60117917ee601d0ec7cf78fbe2121b7bd820935056a16bf24fde9216fdf34b6158fd3d15d89d26fdbec35fa58acf2e9791392;
    5'b10110 : xpb = 1024'h2dcb90c625d8c0cbeccbcb4b435321dadc79a20ccdd795d2323984da2d1ee05edb91d5f0ae6911c171e48a88a6c2f7270c501ee5c9ee6ea08fb21c5b3d4c5841306a7ef966035542b38b28199cd4e65e3dbf0d0010ab13d53b0924a03dba5c17a2c464c30de4acbbbda604627a4a501ba21641c8d996c23557ec6ee381ccb568;
    5'b10111 : xpb = 1024'h802f36dedccee18d8e0616a4cdd166b85fe3596966c64e4c3f2c1950dda17f09b87f3b9b40c5292df9b10aaf15b0c4335d4860fbbff918275adfaed0095e05ac1607b3f70be84c4238860836239f8fd5de042d96dcefd7c39be0ba197de1d8b83f8af1990d6d541be09c106f364f368cc1a8d8a1939cf564fbefabd8a302bda9;
    5'b11000 : xpb = 1024'h21e597a1d1d6cd86643aea2747f5644471d70d952a3d664ece41f471db2170ac922423cd08fac20be21f4b8ea14080754a267b2b9350f162756e01e69a9d3e658755b446023c45fcaae6e5b0118e751c8a4454951cae6ea1472bbd9803deb2c6ad49ec455c2d02ee7cd2359cfa83f6d492619097fd57cb6459836dc93b565f7f;
    5'b11001 : xpb = 1024'h74493dba88ccee4805753580d273a921f540c4f1c32c1ec8db3488e88ba40f576f1189779b56d97869ebcbb5102e4d819b1ebd41895b9ae9409b945b66aeebd06cf2e943a8213cfc2fe1c5cc98591e942a89752be8f3328fa803531144062f674a10791b5bb5aa4e9fc841a9b688dd45b1f42770b75dfe93fd86aabe5c8c67c0;
    5'b11010 : xpb = 1024'h15ff9e7d7dd4da40dbaa09034c97a6ae0734791d86a336cb6a4a6409892400fa48b671a9638c7256525a0c949bbe09c387fcd7715cb374245b29e771f7ee2489de40e9929e7536b6a242a346864803dad6c99c2a28b1c96d534e568fca030975b7cf73c7aa7559213bfe66d77abd9d8d82acdf672118d4935b1a6caef4e00996;
    5'b11011 : xpb = 1024'h6863449634cafb027ce4545cd715eb8b8a9e307a1f91ef45773cf88039a69fa525a3d753f5e889c2da268cbb0aabd6cfd8f5198752be1dab265779e6c3ffd1f4c3de1e90445a2db6273d83630d12ad52770ebcc0f4f68d5bb425ec090a2a86165496009da9fe00815ef472e436c283fea23f763fdb1f07c2ff1da9a4161611d7;
    5'b11100 : xpb = 1024'ha19a55929d2e6fb531927df5139e9179c91e4a5e30907480652d3a137269147ff48bf85be1e22a0c294cd9a963b9311c5d333b72615f6e640e5ccfd553f0aae352c1edf3aae2770999e60dcfb019299234ee3bf34b524395f70ef8790276024c254fb49f8bdaf53fb2a9811faf7444672f82e3644d9ddc25cb16b94ae69b3ad;
    5'b11101 : xpb = 1024'h5c7d4b71e0c907bcf4537338dbb82df51ffb9c027bf7bfc213456817e7a92ff2dc362530507a3a0d4a614dc10529601e16cb75cd1c20a06d0c135f722150b8191ac953dce0931e701e9940f981cc3c10c394045600f9e827c0488500d04edcc55f1b881ff84656b41e20a41eb6fc2ab7928ac50efee010f200b4a889cf9fbbee;
    5'b11110 : xpb = 1024'haee0f18a97bf287e958dbe92663672d2a365535f14e6783c2037fc8e982bce9db9238adae2d65179d22dcde774172d2a67c3b7e3122b49f3d740f1e6ed626584006688da8678156fa39421160896e58863d924eccd3eac1621201a7a10765965fbe214f5f7cefe144116b02b73011128b21d5be7b8e64421a4b7e57ef0d5c42f;
    5'b11111 : xpb = 1024'h5097524d8cc714776bc29214e05a705eb559078ad85d903eaf4dd7af95abc04092c8730cab0bea57ba9c0ec6ffa6e96c54a1d212e583232ef1cf44fd7ea19e3d71b489297ccc0f2a15f4fe8ff685cacf10194beb0cfd42f3cc6b1df89673337469a10fa2468eace6dd4cd5593735d17082d613de22a11a21024ba76f89296605;
    endcase
end

endmodule

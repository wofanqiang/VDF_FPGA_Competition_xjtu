module xpb_5_420
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'hb645701c773797c83fa9dc102ad2d4e30f3a83faa7dfb8a4ce28490d93a9b101c7f41d920506f518401b306d1e07df5be8dcf985acf60317d79c2d006fa8b63091fd085d8c88369249029d78a45d9e61701fc76962b81da7b74a4816f8249cf41c9266751ede6e9b3edad27a778b30e0cadeb60cd259b36922be748165ef446;
    5'b00010 : xpb = 1024'h16c8ae038ee6f2f907f53b82055a5a9c61e7507f54fbf71499c50921b275362038fe83b240a0dea30803660da3c0fbeb7d1b9f30b59ec062faf385a00df516c6123fa10bb19106d2492053af148bb3cc2e03f8ed2c5703b4f6e94902df04939e83924ccea3dbcdd367db5a4f4ef1661c195bd6c19a4b366d2457ce902cbde88c;
    5'b00011 : xpb = 1024'h222d0505565a6c758befd943080787ea92daf8beff79f29ee6a78db28bafd130557dc58b60f14df48c05191475a179e13ba96ec9106e2094786d487014efa2291b5f71918a598a3b6db07d869ed18db24505f563c282858f725ded844e86dd6dc55b7335f5c9b4bd1bc90776f66a192a2609c2226770d1a3b683b5d8431cdcd2;
    5'b00100 : xpb = 1024'h2d915c071dcde5f20fea77040ab4b538c3cea0fea9f7ee29338a124364ea6c4071fd07648141bd461006cc1b4781f7d6fa373e616b3d80c5f5e70b401bea2d8c247f421763220da49240a75e291767985c07f1da58ae0769edd29205be09273d0724999d47b79ba6cfb6b49e9de2cc3832b7ad8334966cda48af9d20597bd118;
    5'b00101 : xpb = 1024'h38f5b308e5415f6e93e514c50d61e286f4c2493e5475e9b3806c96d43e2507508e7c493da1922c9794087f22196275ccb8c50df9c60ce0f77360ce1022e4b8ef2d9f129d3bea910db6d0d135b35d417e7309ee50eed98944694736872d8b710c48edc00499a5829083a461c6455b7f463f6598e401bc0810dadb84686fdac55e;
    5'b00110 : xpb = 1024'h445a0a0aacb4d8eb17dfb286100f0fd525b5f17dfef3e53dcd4f1b65175fa260aafb8b16c1e29be9180a3228eb42f3c27752dd9220dc4128f0da90e029df445236bee32314b31476db60fb0d3da31b648a0beac785050b1ee4bbdb089d0dbadb8ab6e66beb93697a37920eedecd432544c138444cee1a3476d076bb08639b9a4;
    5'b00111 : xpb = 1024'h4fbe610c742852679bda504712bc3d2356a999bda971e0c81a319ff5f09a3d70c77accefe2330b3a9c0be52fbd2371b835e0ad2a7baba15a6e5453b030d9cfb53fdeb3a8ed7b97dffff124e4c7e8f54aa10de73e1b308cf960307f8a0c9004aacc800cd33d815063eb7fbc15944ce56258c16fa59c073e7dff3352f89c98adea;
    5'b01000 : xpb = 1024'h5b22b80e3b9bcbe41fd4ee0815696a71879d41fd53efdc5267142486c9d4d880e3fa0ec902837a8c200d98368f03efadf46e7cc2d67b018bebce168037d45b1848fe842ec6441b4924814ebc522ecf30b80fe3b4b15c0ed3dba5240b7c124e7a0e49333a8f6f374d9f6d693d3bc59870656f5b06692cd9b4915f3a40b2f7a230;
    5'b01001 : xpb = 1024'h66870f10030f4560a3cf8bc9181697bfb890ea3cfe6dd7dcb3f6a917a30f7391007950a222d3e9dda40f4b3d60e46da3b2fc4c5b314a61bd6947d9503ecee67b521e54b49f0c9eb249117893dc74a916cf11e02b478790ae5719c88ceb949849501259a1e15d1e37535b1664e33e4b7e721d4667365274eb238b2188c9569676;
    5'b01010 : xpb = 1024'h71eb6611ca82bedd27ca298a1ac3c50de984927ca8ebd36700d92da87c4a0ea11cf8927b4324592f2810fe4432c4eb99718a1bf38c19c1eee6c19c2045c971de5b3e253a77d5221b6da1a26b66ba82fce613dca1ddb31288d28e6d0e5b16e21891db8009334b05210748c38c8ab6fe8c7ecb31c803781021b5b708d0dfb58abc;
    5'b01011 : xpb = 1024'h7d4fbd1391f63859abc4c74b1d70f25c1a783abc5369cef14dbbb2395584a9b13977d4546374c880ac12b14b04a5698f3017eb8be6e92220643b5ef04cc3fd41645df5c0509da5849231cc42f1005ce2fd15d91873de94634e03118fca992be7d3a4a6708538ec0abb3670b4322fb19a8b791d28d09dab5847e2f018f6147f02;
    5'b01100 : xpb = 1024'h88b414155969b1d62fbf650c201e1faa4b6be2fbfde7ca7b9a9e36ca2ebf44c155f7162d83c537d230146451d685e784eea5bb2441b88251e1b521c053be88a46d7dc646296628edb6c1f61a7b4636c91417d58f0a0a163dc977b6113a1b75b7156dccd7d726d2f46f241ddbd9a864a8982708899dc3468eda0ed7610c737348;
    5'b01101 : xpb = 1024'h94186b1720dd2b52b3ba02cd22cb4cf87c5f8b3ba865c605e780bb5b07f9dfd172765806a415a723b4161758a866657aad338abc9c87e2835f2ee4905ab91407769d96cc022eac56db521ff2058c10af2b19d205a035981844ec5a92a99dbf865736f33f2914b9de2311cb03812117b6a4d4f3ea6ae8e1c56c3abea922d2678e;
    5'b01110 : xpb = 1024'h9f7cc218e850a4cf37b4a08e25787a46ad53337b52e3c19034633febe1347ae18ef599dfc46616753817ca5f7a46e3706bc15a54f75742b4dca8a76061b39f6a7fbd6751daf72fbfffe249c98fd1ea95421bce7c366119f2c060ff1419200955990019a67b02a0c7d6ff782b2899cac4b182df4b380e7cfbfe66a5f139315bd4;
    5'b01111 : xpb = 1024'haae1191aafc41e4bbbaf3e4f2825a794de46dbbafd61bd1a8145c47cba6f15f1ab74dbb8e4b685c6bc197d664c2761662a4f29ed5226a2e65a226a3068ae2acd88dd37d7b3bfb329247273a11a17c47b591dcaf2cc8c9bcd3bd5a39588a25324dac9400dccf087b18aed2552d0127dd2be30caac0534183290928d394f90501a;
    5'b10000 : xpb = 1024'h5982ac6b54962ff74a464391a788d919dc480c9d268182d504b8fb7e0a703f9c4aba0193ae07689a0bcf1263aa9ce9184c2d19f8a4332cc26fceda234d6417f1dadd3aedcf7394d36689ad60b81da307c1acdd0d631f09701bdb61c3df9fa61ed8ad44b6e15760db81aeb9b7fbb0ab77c04d72a820e5638dc4ef97cdd0cddf5;
    5'b10001 : xpb = 1024'h10fc81c87cbcdc7bf89f01fa1d25badfceb829097ce613b79d2e1448b9e19f09e12ae1f25b30e5db24bea42d0c8a4c874350a137e51292fda476b0723bd0cce226cda434b5bfbcb65af8c4ad95c7b416931cca476c5d72717d325a9dad7c44312f53fab2c0035cf76c0898c32733bdc588b2c28b4f33f16f6e7ae0c4f36bd23b;
    5'b10010 : xpb = 1024'h1c60d8ca443055f87c999fbb1fd2e82dffabd14927640f41ea1098d9931c3a19fdaa23cb7b81552ca8c05733de6aca7d01de70d03fe1f32f21f0734242cb58452fed74ba8e88401f7f88ee85200d8dfcaa1ec6be0288f44bf8a6ff1f1cfe8e00711d211a11f143e11ff645eaceac70d39560adec1c598ca600a6c80d09cac681;
    5'b10011 : xpb = 1024'h27c52fcc0ba3cf7500943d7c2280157c309f7988d1e20acc36f31d6a6c56d52a1a2965a49bd1c47e2cc20a3ab04b4872c06c40689ab153609f6a361249c5e3a8390d45406750c388a419185caa5367e2c120c33498b47626741ba3a08c80d7cfb2e6478163df2acad3e3f312762523e1a20e994ce97f27dc92d2af552029bac7;
    5'b10100 : xpb = 1024'h332986cdd31748f1848edb3d252d42ca619321c87c60065683d5a1fb4591703a36a8a77dbc2233cfb0c3bd41822bc6687efa1000f580b3921ce3f8e250c06f0b422d15c6401946f1c8a94234349941c8d822bfab2edff800ef904821fc03219ef4af6de8b5cd11b487d1a03a1d9dd6efaebc84adb6a4c31324fe969d3688af0d;
    5'b10101 : xpb = 1024'h3e8dddcf9a8ac26e088978fe27da70189286ca0826de01e0d0b8268c1ecc0b4a5327e956dc72a32134c57048540c445e3d87df99505013c39a5dbbb257bafa6e4b4ce64c18e1ca5aed396c0bbedf1baeef24bc21c50b79db6b04eca36b856b6e3678945007baf89e3bbf4d61c51689fdbb6a700e83ca5e49b72a7de54ce7a353;
    5'b10110 : xpb = 1024'h49f234d161fe3bea8c8416bf2a879d66c37a7247d15bfd6b1d9aab1cf806a65a6fa72b2ffcc31272b8c7234f25ecc253fc15af31ab1f73f517d77e825eb585d1546cb6d1f1aa4dc411c995e34924f5950626b8985b36fbb5e6799124db07b53d7841bab759a8df87efacfa896c8f3d0bc8185b6f50eff9804956652d63469799;
    5'b10111 : xpb = 1024'h55568bd32971b567107eb4802d34cab4f46e1a877bd9f8f56a7d2fadd141416a8c266d091d1381c43cc8d655f7cd4049baa37eca05eed4269551415265b011345d8c8757ca72d12d3659bfbad36acf7b1d28b50ef1627d9061ee35a64a89ff0cba0ae11eab96c671a39aa7b11407f019d4c646d01e1594b6db824c7579a58bdf;
    5'b11000 : xpb = 1024'h60bae2d4f0e52ee3947952412fe1f8032561c2c72657f47fb75fb43eaa7bdc7aa8a5aee23d63f115c0ca895cc9adbe3f79314e6260be345812cb04226caa9c9766ac57dda33b54965ae9e9925db0a961342ab185878dff6add62da27ba0c48dbfbd40785fd84ad5b578854d8bb80a327e1743230eb3b2fed6dae33bd90048025;
    5'b11001 : xpb = 1024'h6c1f39d6b858a8601873f002328f255156556b06d0d5f00a044238cf83b6778ac524f0bb5db4606744cc3c639b8e3c3537bf1dfabb8d94899044c6f273a527fa6fcc28637c03d7ff7f7a1369e7f683474b2cadfc1db9814558d77ea9298e92ab3d9d2ded4f7294450b76020062f95635ee221d91b860cb23ffda1b05a663746b;
    5'b11010 : xpb = 1024'h778390d87fcc21dc9c6e8dc3353c529f874913467b53eb945124bd605cf1129ae1a432947e04cfb8c8cdef6a6d6eba2af64ced93165cf4bb0dbe89c27a9fb35d78ebf8e954cc5b68a40a3d41723c5d2d622eaa72b3e5031fd44c232a9910dc7a7f665454a1607b2ebf63af280a720943fad008f28586665a9206024dbcc268b1;
    5'b11011 : xpb = 1024'h82e7e7da473f9b5920692b8437e97fedb83cbb8625d1e71e9e0741f1362badaafe23746d9e553f0a4ccfa2713f4f3820b4dabd2b712c54ec8b384c92819a3ec0820bc96f2d94ded1c89a6718fc8237137930a6e94a1084fa4fc0c7ac08932649c12f7abbf34e621873515c4fb1eabc52077df45352ac01912431e995d3215cf7;
    5'b11100 : xpb = 1024'h8e4c3edc0eb314d5a463c9453a96ad3be93063c5d04fe2a8eae9c6820f6648bb1aa2b646bea5ae5bd0d15578112fb61673688cc3cbfbb51e08b20f628894ca238b2b99f5065d623aed2a90f086c810f99032a35fe03c06d4cb356c2d7815701902f8a123453c4902273f097759636f60142bdfb41fd19cc7b65dd0dde980513d;
    5'b11101 : xpb = 1024'h99b095ddd6268e52285e67063d43da8a1a240c057acdde3337cc4b12e8a0e3cb3721f81fdef61dad54d3087ee310340c31f65c5c26cb154f862bd2328f8f5586944b6a7adf25e5a411babac8110deadfa7349fd6766788af46aa10aee797b9e844c1c78a972a2febdb2cb69f00dc226e20d9cb14ecf737fe4889b825ffdf4583;
    5'b11110 : xpb = 1024'ha514ecdf9d9a07ceac5904c73ff107d84b17b445254bd9bd84aecfa3c1db7edb53a139f8ff468cfed8d4bb85b4f0b201f0842bf4819a758103a595029689e0e99d6b3b00b7ee690d364ae49f9b53c4c5be369c4d0c930a89c21eb530571a03b7868aedf1e91816d58f1a63c6a854d57c2d87b675ba1cd334dab59f6e163e39c9;
    5'b11111 : xpb = 1024'hb07943e1650d814b3053a288429e35267c0b5c84cfc9d547d19154349b1619eb70207bd21f96fc505cd66e8c86d12ff7af11fb8cdc69d5b2811f57d29d846c4ca68b0b8690b6ec765adb0e7725999eabd53898c3a2be8c643d9359b1c69c4d86c85414593b05fdbf430810ee4fcd888a3a35a1d687426e6b6ce186b62c9d2e0f;
    endcase
end

endmodule

module xpb_5_720
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h1426ace823e2e6b309fb918bcacc7a213eca870b7924e37ddc834bcf1ecbb4c32ddec2b8317ef7dacb5ff346c1021129d1220c5bf23be56b9c7799d9c9b81ce49c1267223420024b2378f198a9c8d70492d61f146955fc59e224951488896bbe4dd7caa330bc259080193073689288aaed855e138e71561c25db6791d6cc5f62;
    5'b00010 : xpb = 1024'h284d59d047c5cd6613f723179598f4427d950e16f249c6fbb906979e3d9769865bbd857062fdefb596bfe68d82042253a24418b7e477cad738ef33b3937039c93824ce446840049646f1e3315391ae0925ac3e28d2abf8b3c4492a291112d77c9baf954661784b21003260e6d1251155db0abc271ce2ac384bb6cf23ad98bec4;
    5'b00011 : xpb = 1024'h3c7406b86ba8b4191df2b4a360656e63bc5f95226b6eaa799589e36d5c631e49899c4828947ce790621fd9d44306337d73662513d6b3b042d566cd8d5d2856add43735669c6006e16a6ad4c9fd5a850db8825d3d3c01f50da66dbf3d999c433ae9875fe9923470b1804b915a39b79a00c8901a3aab540254719236b584651e26;
    5'b00100 : xpb = 1024'h509ab3a08f8b9acc27ee462f2b31e884fb2a1c2de4938df7720d2f3c7b2ed30cb77b0ae0c5fbdf6b2d7fcd1b040844a74488316fc8ef95ae71de676726e0739270499c88d080092c8de3c662a7235c124b587c51a557f167889254522225aef9375f2a8cc2f096420064c1cda24a22abb615784e39c55870976d9e475b317d88;
    5'b00101 : xpb = 1024'h64c16088b36e817f31e9d7baf5fe62a639f4a3395db871754e907b0b99fa87cfe559cd98f77ad745f8dfc061c50a55d115aa3dcbbb2b7b1a0e560140f09890770c5c03ab04a00b77b15cb7fb50ec3316de2e9b660eadedc16ab6e966aaaf1ab78536f52ff3acbbd2807df2410adcab56a39ad661c836ae8cbd4905d931fddcea;
    5'b00110 : xpb = 1024'h78e80d70d75168323be56946c0cadcc778bf2a44d6dd54f32b13c6dab8c63c931338905128f9cf20c43fb3a8860c66fae6cc4a27ad676085aacd9b1aba50ad5ba86e6acd38c00dc2d4d5a993fab50a1b7104ba7a7803ea1b4cdb7e7b33388675d30ebfd32468e163009722b4736f34019120347556a804a8e3246d6b08ca3c4c;
    5'b00111 : xpb = 1024'h8d0eba58fb344ee545e0fad28b9756e8b789b15050023871079712a9d791f156411753095a78c6fb8f9fa6ef470e7824b7ee56839fa345f1474534f48408ca404480d1ef6ce0100df84e9b2ca47de12003dad98ee159e6752f00138fbbc1f23420e68a76552506f380b05327dc01bcac7ea59288e5195ac508ffd4fcdf969bae;
    5'b01000 : xpb = 1024'ha13567411f1735984fdc8c5e5663d109f654385bc9271beee41a5e78f65da6196ef615c18bf7bed65aff9a360810894e891062df91df2b5ce3bccece4dc0e724e0933911a10012591bc78cc54e46b82496b0f8a34aafe2cf1124a8a4444b5df26ebe551985e12c8400c9839b449445576c2af09c738ab0e12edb3c8eb662fb10;
    5'b01001 : xpb = 1024'h4aeced3810be7828ed2a61310d603d9c3a8bc366cd45ef542c0f0f26226add4998c5b00f350382287014e35e5b489adf61847556168407ccf952949dca68f5808566b85258f175f2ca67bbb5f33caf835821e1f277fb2183dbcabbe12aa271e8d8e8d9305d45986fa22cd2fb556a7d90ad66fcdb1b0a9cd0e47291c044cf407;
    5'b01010 : xpb = 1024'h18d57bbba4eece3598ce379edba27dfb02734341e5f942731f443cc180f26297c76b1db924cf2ffd5261417ca6b69ad7c73a53b153a425e86c0cc323a65eac3ca468d2a759af19aa501f6d5408fca1fcc8583d3390d5ae721fe140d29b3392dcdb66583636907f177a3bfda31de93083f85bcde14021ffe9342290addb195369;
    5'b01011 : xpb = 1024'h2cfc28a3c8d1b4e8a2c9c92aa66ef81c413dca4d5f1e25f0fbc788909fbe175af549e071564e27d81dc134c367b8ac01985c600d45e00b5408845cfd7016c921407b39c98dcf1bf573985eecb2c579015b2e5c47fa2baacc0205d5e723bcfe9b293e22d9674ca4a7fa552e16867bb92ee5e12bf4ce93560559fdf83fb1e5b2cb;
    5'b01100 : xpb = 1024'h4122d58becb49b9bacc55ab6713b723d80085158d843096ed84ad45fbe89cc1e2328a32987cd1fb2e921280a28babd2b697e6c69381bf0bfa4fbf6d739cee605dc8da0ebc1ef1e40971150855c8e5005ee047b5c6381a725e42a6afbac466a597715ed7c9808ca387a6e5e89ef0e41d9d3668a085d04ac217fd95fd188b2122d;
    5'b01101 : xpb = 1024'h554982741097824eb6c0ec423c07ec5ebed2d8645167ececb4ce202edd5580e1510765e1b94c178db4811b50e9bcce553aa078c52a57d62b417390b1038702ea78a0080df60f208bba8a421e0657270a80da9a70ccd7a37fc64f001034cfd617c4edb81fc8c4efc8fa878efd57a0ca84c0ebe81beb76023da5b4c7635f7e718f;
    5'b01110 : xpb = 1024'h69702f5c347a6901c0bc7dce06d4667ffd9d5f6fca8cd06a91516bfdfc2135a47ee62899eacb0f687fe10e97aabedf7f0bc285211c93bb96ddeb2a8acd3f1fcf14b26f302a2f22d6de0333b6b01ffe0f13b0b985362d9fd9a8739524bd5941d612c582c2f98115597aa0bf70c033532fae71462f79e75859cb902ef5364ad0f1;
    5'b01111 : xpb = 1024'h7d96dc44585d4fb4cab80f59d1a0e0a13c67e67b43b1b3e86dd4b7cd1aecea67acc4eb521c4a07434b4101de6bc0f0a8dce4917d0ecfa1027a62c46496f73cb3b0c4d6525e4f2522017c254f59e8d513a686d8999f839c338a982a3945e2ad94609d4d662a3d3ae9fab9efe428c5dbda9bf6a4430858ae75f16b96870d173053;
    5'b10000 : xpb = 1024'h91bd892c7c403667d4b3a0e59c6d5ac27b326d86bcd697664a58039c39b89f2adaa3ae0a4dc8ff1e16a0f5252cc301d2ae069dd9010b866e16da5e3e60af59984cd73d74926f276d24f516e803b1ac18395cf7ae08d9988d6cbcbf4dce6c1952ae7518095af9607a7ad3205791586485897c025696ca04921746fe18e3e38fb5;
    5'b10001 : xpb = 1024'ha5e43614a0231d1adeaf32716739d4e3b9fcf49235fb7ae426db4f6b588453ee088270c27f47f6f8e200e86bedc512fc7f28aa34f3476bd9b351f8182a67767ce8e9a496c68f29b8486e0880ad7a831ccc3316c2722f94e74ee1546256f58510fc4ce2ac8bb5860afaec50caf9eaed307701606a253b5aae3d2265aabaafef17;
    5'b10010 : xpb = 1024'h95d9da70217cf051da54c2621ac07b38751786cd9a8bdea8581e1e4c44d5ba93318b601e6a070450e029c6bcb69135bec308eaac2d080f99f2a5293b94d1eb010acd70a4b1e2ebe594cf776be6795f06b043c3e4eff64307b79577c25544e3d1b1d1b260ba8b30df4459a5f6aad4fb215acdf9b6361539a1c8e52380899e80e;
    5'b10011 : xpb = 1024'h1d844a8f25fab5b827a0ddb1ec7881d4c61bff7852cda16862052db3e319106c60f778ba181f681fd9628fb28c6b2485bd529b06b50c66653ba1ec6d83053b94acbf3e2c7f3e31097cc5e90f68306cf4fdda5b52b855608a5d9dec90adddb9fb68f4e5c93c64d89e745ecad2d33fd85d03323daef1d2a9b64269b9c9df664770;
    5'b10100 : xpb = 1024'h31aaf77749dd9c6b319c6f3db744fbf604e68683cbf284e63e88798301e4c52f8ed63b72499e5ffaa4c282f94d6d35af8e74a762a7484bd0d81986474cbd587948d1a54eb35e3354a03edaa811f943f990b07a6721ab5ce43fc281a5366725b9b6ccb06c6d20fe2ef477fb463bd26107f0b79bc28043ffd26845215bb632a6d2;
    5'b10101 : xpb = 1024'h45d1a45f6dc0831e3b9800c98211761743b10d8f451768641b0bc55220b079f2bcb4fe2a7b1d57d5702276400e6f46d95f96b3be9984313c749120211675755de4e40c70e77e359fc3b7cc40bbc21afe2386997b8b01593e21e716b9bef0917804a47b0f9ddd23bf74912bb9a464e9b2de3cf9d60eb555ee8e2088ed8cff0634;
    5'b10110 : xpb = 1024'h59f8514791a369d1459392554cddf038827b949abe3c4be1f78f11213f7c2eb5ea93c0e2ac9c4fb03b826986cf71580330b8c01a8bc016a81108b9fae02d924280f673931b9e37eae730bdd9658af202b65cb88ff4575598040babce4779fd36527c45b2ce99494ff4aa5c2d0cf7725dcbc257e99d26ac0ab3fbf07f63cb6596;
    5'b10111 : xpb = 1024'h6e1efe2fb58650844f8f23e117aa6a59c1461ba637612f5fd4125cf05e47e3791872839ade1b478b06e25ccd9073692d01dacc767dfbfc13ad8053d4a9e5af271d08dab54fbe3a360aa9af720f53c9074932d7a45dad51f1e63040e2d00368f4a0541055ff556ee074c38ca07589fb08b947b5fd2b980226d9d758113a97c4f8;
    5'b11000 : xpb = 1024'h8245ab17d9693737598ab56ce276e47b0010a2b1b08612ddb095a8bf7d13983c465146530f9a3f65d242501451757a56d2fcd8d27037e17f49f7edae739dcc0bb91b41d783de3c812e22a10ab91ca00bdc08f6b8c7034e4bc854d5f7588cd4b2ee2bdaf930119470f4dcbd13de1c83b3a6cd1410ba095842ffb2bfa31164245a;
    5'b11001 : xpb = 1024'h966c57fffd4c1dea638646f8ad435e9c3edb29bd29aaf65b8d18f48e9bdf4cff7430090b411937409da2435b12778b80a41ee52e6273c6eae66f87883d55e8f0552da8f9b7fe3ecc519b92a362e577106edf15cd30594aa5aa796b0be11640713c03a59c60cdba0174f5ed8746af0c5e94527224487aae5f258e2734e83083bc;
    5'b11010 : xpb = 1024'haa9304e8212f049d6d81d884780fd8bd7da5b0c8a2cfd9d9699c405dbaab01c2a20ecbc372982f1b690236a1d3799caa7540f18a54afac5682e72162070e05d4f140101bec1e41177514843c0cae4e1501b534e199af46ff8c9e0020699fac2f89db703f9189df91f50f1dfaaf41950981d7d037d6ec047b4b698ec6befce31e;
    5'b11011 : xpb = 1024'he0c6c7a8323b687ac77f23932820b8d4afa34a3467d1cdfc842d2d72674097dcca51102d9f0a8679503eaa1b11d9d09e248d6002438c1766ebf7bdd95f3ae081903428f70ad461d85f373321d9b60e8a0865a5d767f1648b936033a37fe755ba8aba8b9117d0c94ee68678f2003f78b20834f691511fd672ad57b540ce6dc15;
    5'b11100 : xpb = 1024'h22331962a7069d3ab67383c4fd4e85ae89c4bbaebfa2005da4c61ea6453fbe40fa83d3bb0b6fa0426063dde8721fae33b36ae25c1674a6e20b3715b75fabcaecb515a9b1a4cd4868a96c64cac76437ed335c7971dfd512a29b5a984ec087e119f683735c423932256e819802889680360e08ad7ca383538350b0e2e5e3b33b77;
    5'b11101 : xpb = 1024'h3659c64acae983edc06f1550c81affcfc88f42ba38c6e3db81496a75640b7304286296733cee981d2bc3d12f3321bf5d848ceeb808b08c4da7aeaf912963e7d1512810d3d8ed4ab3cce55663712d0ef1c6329886492b0efc7d7f2d6349114cd8445b3dff72f557b5ee9ac875f12908e0fb8e0b9031f4a99f768c4a77ba7f9ad9;
    5'b11110 : xpb = 1024'h4a807332eecc6aa0ca6aa6dc92e779f10759c9c5b1ebc7595dccb64482d727c75641592b6e6d8ff7f723c475f423d08755aefb13faec71b94426496af31c04b5ed3a77f60d0d4cfef05e47fc1af5e5f65908b79ab2810b565fa3c277d19ab896923308a2a3b17d466eb3f8e959bb918be91369a3c065ffbb9c67b209914bfa3b;
    5'b11111 : xpb = 1024'h5ea7201b12af5153d46638685db3f412462450d12b10aad73a500213a1a2dc8a84201be39fec87d2c283b7bcb525e1b126d1076fed285724e09de344bcd4219a894cdf18412d4f4a13d73994c4bebcfaebded6af1bd707b041c8578c5a242454e00ad345d46da2d6eecd295cc24e1a36d698c7b74ed755d7c243199b6818599d;
    endcase
end

endmodule

module xpb_5_25
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h8344e53ae734c1f631ad6c8ab422f8b83871fe4cb59dd8d98005560613ea9ad6047531d0afce220ce17bf6589c7c5f70c8f5d51b42e166ff0b486a65568766ee776e0d23a43532282c87c74014b36573e3ff8add0ce28175356fb0afc2c713ea4de1c9938b54b3b79d54ca58d7e1ec474f9b38eab026b7ecdb925cc5a600fa7b;
    5'b00010 : xpb = 1024'h55dc85200c7b4f239855613e57ebaa1eff6df96895c4113b822df2b674d288a405a1e6289575c58b2399ad6a559aae172dd18250630ffdb265f1956c723c592b7a8ce59898d9670b46758bdd908b06b6d3fa1c218d3ed5d9b552cf64cb6385426cbc00fd65e06ee1b3e9add2b7f3b265505c92f3100212a970b53e86c31f8e8b;
    5'b00011 : xpb = 1024'h2874250531c1dc50fefd55f1fbb45b85c669f48475ea499d84568f66d5ba767206ce9a807b1d690965b7647c0eb8fcbd92ad2f85833e9465c09ac0738df14b687dabbe0d8d7d9bee6063507b0c62a7f9c3f4ad660d9b2a3e3535ee19d3fff69a8b963867406c2a0bca7e914c98057883511decfb6fdd6d6605d82047e03e229b;
    5'b00100 : xpb = 1024'habb90a4018f69e4730aac27cafd7543dfedbf2d12b882277045be56ce9a511480b43cc512aeb8b1647335ad4ab355c2e5ba304a0c61ffb64cbe32ad8e478b256f519cb3131b2ce168ceb17bb21160d6da7f438431a7dabb36aa59ec996c70a84d97801facbc0ddc367d35ba56fe764caa0b925e620042552e16a7d0d863f1d16;
    5'b00101 : xpb = 1024'h7e50aa253e3d2b749752b73053a005a4c5d7eded0bae5ad90684821d4a8cff160c7080a910932e94895111e66453aad4c07eb1d5e64e9218268c55e0002da493f838a3a6265702f9a6d8dc589cedaeb097eec9879ada0017ea88bd7e9f637bdcf8523964a64c98ed7e683f1f4ff92ae8a17a7fee7fdf800f768d5ecea35db126;
    5'b00110 : xpb = 1024'h50e84a0a6383b8a1fdfaabe3f768b70b8cd3e908ebd4933b08ad1ecdab74ece40d9d3500f63ad212cb6ec8f81d71f97b255a5f0b067d28cb813580e71be296d0fb577c1b1afb37dcc0c6a0f618c54ff387e95acc1b36547c6a6bdc33a7ffed35172c70ce80d8541794fd2299300af106a23bd9f6dfbadacc0bb0408fc07c4536;
    5'b00111 : xpb = 1024'h237fe9ef88ca45cf64a2a0979b31687253cfe424cbfacb9d0ad5bb7e0c5cdab20ec9e958dbe275910d8c8009d69048218a360c4026abbf7edbdeabee3797890dfe7654900f9f6cbfdab46593949cf13677e3ec109b92a8e0ea4efae8b09c5e8d3606a8385b640f41ab920613101cb724a2fd33ff3f963588a0d32250dd9ad946;
    5'b01000 : xpb = 1024'ha6c4cf2a6fff07c596500d224f54612a8c41e2718198a4768adb118420477588133f1b298bb0979def087662730ca792532be15b698d267de72716538e1eeffc75e461b3b3d49ee8073c2cd3a95056aa5be376eda8752a561fbeab987363727783e871cbe6b8c2f948e6d06be7fea36bf2986ce9efbced757c657f16839bd3c1;
    5'b01001 : xpb = 1024'h795c6f0f954594f2fcf801d5f31d1291533ddd8d61bedcd88d03ae34812f6356146bcf8171583b1c31262d742c2af638b8078e9089bbbd3141d0415aa9d3e23979033a28a878d3cb2129f1712527f7ed4bde083228d17eba9fa1ca4d7bffe3cfa2c2a935c1447e235f7bb3e5c8106989f359c6f24f984832118860d7a0ba67d1;
    5'b01010 : xpb = 1024'h4bf40ef4ba8c2220639ff68996e5c3f81a39d8a941e5153a8f2c4ae4e2175124159883d956ffde9a7343e485e54944df1ce33bc5a9ea53e49c796c61c588d4767c22129d9d1d08ae3b17b60ea0ff99303bd89976a92dd31f1f84e902849c5527c19ce09f9bd0394d7610975fa8222fa7f41b20faaf73a2eea6ab4298bdd8fbe1;
    5'b01011 : xpb = 1024'h1e8baed9dfd2af4dca47eb3d3aae755ee135d3c5220b4d9c9154e79542ff3ef216c538313ca78218b5619b979e67938581bee8faca18ea97f7229768e13dc6b37f40eb1291c13d9155057aac1cd73a732bd32abb298a27839f6807b78d38c67fe0771809765bf4778ca57ad98833f5c5f4dc7b030f4efdab3bce2459daf78ff1;
    5'b01100 : xpb = 1024'ha1d09414c7077143fbf557c7eed16e1719a7d211d7a92676115a3d9b56e9d9c81b3a6a01ec75a42596dd91f03ae3f2f64ab4be160cfa5197026b01ce37c52da1f6aef83635f66fb9818d41ec318a9fe70fd2b598366ca8f8d4d7b8674fffda6a2e58e19d01b0a82f29fa45326015e20d4477b3edbf75b5981760811f80f88a6c;
    5'b01101 : xpb = 1024'h746833f9ec4dfe71629d4c7b929a1f7de0a3cd2db7cf5ed81382da4bb7d1c7961c671e59d21d47a3d8fb4901f402419caf906b4b2d28e84a5d142cd5537a1fdef9cdd0ab2a9aa49c9b7b0689ad624129ffcd46dcb6c8fd5d54bad71c589c4bc24d331906dc3c6359408f28ac4027a82b45390df61f511054ac8362e09e171e7c;
    5'b01110 : xpb = 1024'h46ffd3df11948b9ec945412f3662d0e4a79fc84997f5973a15ab76fc18b9b5641d93d2b1b7c4eb221b190013ad209043146c18804d577efdb7bd57dc6f2f121bfceca9201f3ed97fb568cb272939e26cefc7d821372551c1d49df5d16138bd1a6c0d5070b6c81e8357240c2620396e4945fa67fe7f2c6b1141a644a1bb35b28c;
    5'b01111 : xpb = 1024'h199773c436db18cc2fed35e2da2b824b6e9bc365781bcf9c17d413ac79a1a3321ec087099d6c8ea05d36b725663edee97947c5b56d8615b1126682e38ae40459000b819513e30e62cf568fc4a51183afdfc26965b781a6265481148669d52e728ae787da9153d9ad6db8efa0004b346746bbc206df07c5cdd6c92662d854469c;
    5'b10000 : xpb = 1024'h9cdc58ff1e0fdac2619aa26d8e4e7b03a70dc1b22db9a87597d969b28d8c3e082335b8da4d3ab0ad3eb2ad7e02bb3e5a423d9ad0b0677cb01daeed48e16b6b4777798eb8b818408afbde5704b9c4e923c3c1f442c464279b89f0c5362c9c425cd8c9516e1ca88d650b0db9f8d82d20ae9656faf18f2e7dbab25b83287e554117;
    5'b10001 : xpb = 1024'h6f73f8e4435667efc842972132172c6a6e09bcce0ddfe0d79a020662ee742bd624626d3232e2542b80d0648fbbd98d00a7194805d09613637858184ffd205d847a98672dacbc756e15cc1ba2359c8a66b3bc858744c07c0009d3e3eb3538b3b4f7a388d7f734488f21a29d72b83ee6cc971854f9ef09d877477e64e99b73d527;
    5'b10010 : xpb = 1024'h420b98c9689cf51d2eea8bd4d5dfddd13505b7e9ee0619399c2aa3134f5c19a4258f218a1889f7a9c2ee1ba174f7dba70bf4f53af0c4aa16d301435718d54fc17db73fa2a160aa512fb9e03fb1742ba9a3b716cbc51cd06489b702a03dd5250d167dc041d1c003b9383780ec9850acea97d9af024ee53333dca146aab8926937;
    5'b10011 : xpb = 1024'h14a338ae8de3824a9592808879a88f37fc01b305ce2c519b9e533fc3b044077226bbd5e1fe319b28050bd2b32e162a4d70d0a27010f340ca2daa6e5e348a41fe80d618179604df3449a7a4dd2d4bccec93b1a810457924c9099a2155467196653557f7abac4bbee34ecc646678627308989b090aaec08df071c4286bd5b0fd47;
    5'b10100 : xpb = 1024'h97e81de975184440c73fed132dcb87f03473b15283ca2a751e5895c9c42ea2482b3107b2adffbd34e687c90bca9289be39c6778b53d4a7c938f2d8c38b11a8ecf844253b3a3a115c762f6c1d41ff326077b132ed525ba63e3f09d2050938aa4f8339c13f37a0729aec212ebf50445f4fe83641f55ee745dd4d5685317bb1f7c2;
    5'b10101 : xpb = 1024'h6a7fbdce9a5ed16e2de7e1c6d1943956fb6fac6e63f062d72081327a251690162c5dbc0a93a760b328a5801d83b0d8649ea224c074033e7c939c03caa6c69b29fb62fdb02ede463f901d30babdd6d3a367abc431d2b7faa2beecf0ba11d51ba7a213f8a9122c2dc502b612393056256de8f79bfdbec2a099e27966f298d08bd2;
    5'b10110 : xpb = 1024'h3d175db3bfa55e9b948fd67a755ceabdc26ba78a44169b3922a9cf2a85fe7de42d8a7062794f04316ac3372f3ccf270b037dd1f59431d52fee452ed1c27b8d66fe81d62523827b22aa0af55839ae74e657a6557653144f073ed00f6f1a718cffc0ee3012ecb7e8ef194af5b31067eb8be9b8f6061e9dfb56779c48b3b5ef1fe2;
    5'b10111 : xpb = 1024'hfaefd98e4ebebc8fb37cb2e19259c248967a2a6243cd39b24d26bdae6e66bb22eb724ba5ef6a7aface0ee40f5ed75b168597f2ab4606be348ee59d8de307fa401a0ae9a1826b005c3f8b9f5b586162947a0e6bad370a36bbeb32e24230dfe57dfc8677cc743a4192fdfd92cf079b1a9ea7a500e7e7956130cbf2a74d30db3f2;
    5'b11000 : xpb = 1024'h92f3e2d3cc20adbf2ce537b8cd4894dcc1d9a0f2d9daac74a4d7c1e0fad10688332c568b0ec4c9bc8e5ce4999269d522314f5445f741d2e25436c43e34b7e692790ebbbdbc5be22df0808135ca397b9d2ba07197e05324e0f422ded3e5d512422daa3110529857d0cd34a385c85b9df13a1588f92ea00dffe851873a790eae6d;
    5'b11001 : xpb = 1024'h658b82b8f1673aec938d2c6c7111464388d59c0eba00e4d6a7005e915bb8f45634590ae2f46c6d3ad07a9bab4b8823c8962b017b17706995aedfef45506cd8cf7c2d9432b10017110a6e45d346111ce01b9b02dc60af79457405fd88ee71839a4c84687a2d2412fae3c986ffa86d640f3ad6e3018e7b68bc7d7468fb962d427d;
    5'b11010 : xpb = 1024'h3823229e16adc819fa35212014d9f7aa4fd1972a9a271d38a928fb41bca0e2243585bf3ada1410b9129852bd04a6726efb06aeb0379f004909891a4c6c21cb0c7f4c6ca7a5a44bf4245c0a70c1e8be230b959420e10bcda9f3e91c3df70df4f26b5e9fe407afce24fa5e6a79887f2a2d3b983d09ee56c37912974abcb34bd68d;
    5'b11011 : xpb = 1024'habac2833bf4554760dd15d3b8a2a91116cd92467a4d559aab5197f21d88cff236b27392bfbbb43754b609cebdc4c1155fe25be557cd96fc6432455387d6bd49826b451c9a4880d73e49cf0e3dc05f65fb9025656168220e73cc3af2ffaa664a8a38d74de23b894f10f34df36890f04b3c5997124e321e35a7ba2c7dd06a6a9d;
    5'b11100 : xpb = 1024'h8dffa7be2329173d928a825e6cc5a1c94f3f90932feb2e742b56edf831736ac83b27a5636f89d644363200275a41208628d831009aaefdfb6f7aafb8de5e2437f9d952403e7db2ff6ad1964e5273c4d9df8fb0426e4aa383a93beba2c2717a34d81aa0e16d903d06ae48184c4072dc928bf4cffcfe58d622834c8943766b6518;
    5'b11101 : xpb = 1024'h609747a3486fa46af9327712108e5330163b8baf101166d62d7f8aa8925b58963c5459bb553179c2784fb739135f6f2c8db3de35badd94aeca23dabffa131674fcf82ab53321e7e284bf5aebce4b661ccf8a4186eea6f7e8291f0a57cb0deb8cf6f4d84b481bf830c4dcfbc62084a2b08cb62a055e3430df186f6b049389f928;
    5'b11110 : xpb = 1024'h332ee7886db631985fda6bc5b4570496dd3786caf0379f382fa82758f34346643d810e133ad91d40ba6d6e4acc7dbdd2f28f8b6adb0c2b6224cd05c715c808b20017032a27c61cc59ead1f894a23075fbf84d2cb6f034c4ca902290cd3aa5ce515cf0fb522a7b35adb71df40009668ce8d77840dbe0f8b9bad924cc5b0a88d38;
    5'b11111 : xpb = 1024'h5c6876d92fcbec5c6826079581fb5fda43381e6d05dd79a31d0c409542b34323eadc26b2080c0befc8b255c859c0c79576b389ffb3ac2157f7630ce317cfaef0335db9f1c6a51a8b89ae426c5faa8a2af7f640fef5fa0b128e547c1dc46ce3d34a9471efd336e84f206c2b9e0a82eec8e38de161deae65842b52e86cdc72148;
    endcase
end

endmodule

module xpb_5_265
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h62cbc9dd4e2ab0c7937011a7a7c05811533afcdb40252c10e1b2ca28874eb58a1029c9c9e24d4742ec5e44a6a057a7850f825faec3181e970dac39202e1caf491d5d0c1f0d2568dc78aaccf2ebc8a4d60550b3b475e9b3d8b33c63f01e86687016f76b0037f5714b2f9f091c92dab5c7dddb0816af5c5c663b8731a5afa696ec;
    5'b00010 : xpb = 1024'h14ea4e64da672cc65bdaab783f2668d134fff685aad2b7aa4588dafb5b9abe0c1d0b161afa740ff7395e4a065d513e3fbaea9777637d6ce26ab932e22166e9e0c66ae38f6ab9d473debb97433eb5857b169c6dd05f4d3aa0b0ec35e582e22e4dfee743d6bf21ea08d87e2b5a2de545666cdc314b0e6d5b9c309ee846d66ac76d;
    5'b00011 : xpb = 1024'h77b618422891dd8def4abd1fe6e6c0e2883af360eaf7e3bb273ba523e2e973962d34dfe4dcc1573a25bc8eacfda8e5c4ca6cf72626958b7978656c024f839929e3c7efae77df3d50576664362a7e2a511bed2184d536ee79642899d5a16896be15deaed6f7175b54081d3476c0bffb2e4ab73961bdc9b8026c2619ec86115e59;
    5'b00100 : xpb = 1024'h29d49cc9b4ce598cb7b556f07e4cd1a269ffed0b55a56f548b11b5f6b7357c183a162c35f4e81fee72bc940cbaa27c7f75d52eeec6fad9c4d57265c442cdd3c18cd5c71ed573a8e7bd772e867d6b0af62d38dba0be9a754161d86bcb05c45c9bfdce87ad7e43d411b0fc56b45bca8accd9b862961cdab738613dd08dacd58eda;
    5'b00101 : xpb = 1024'h8ca066a702f90a544b256898260d29b3bd3ae9e695ca9b656cc4801f3e8431a24a3ff5ffd73567315f1ad8b35afa240485578e9d8a12f85be31e9ee470ea830aaa32d33de29911c43621fb796933afcc32898f553484291a1514cfbb244ac50c14c5f2adb639455ce09b5fd0eea54094b7936aaccc37139e9cc502335c7c25c6;
    5'b00110 : xpb = 1024'h3ebeeb2e8f35865313900268bd733a739effe391007826fed09a90f212d03a2457214250ef5c2fe5ac1ade1317f3babf30bfc6662a7846a7402b98a66434bda25340aaae402d7d5b9c32c5c9bc20907143d549711de7afe212c4a1b088a68ae9fcb5cb843d65be1a897a820e89afd033469493e12b4812d491dcb8d483405647;
    5'b00111 : xpb = 1024'ha18ab50bdd60371aa700141065339284f23ae06c409d530fb24d5b1a9a1eefae674b0c1ad1a97728987922b9b84b624440422614ed90653e4dd7d1c692516ceb709db6cd4d52e63814dd92bca7e935474925fd2593d163bac60105a0a72cf35a13ad3684755b2f65b9198b2b1c8a85fb246f9bf7daa46f3acd63ea7a32e6ed33;
    5'b01000 : xpb = 1024'h53a93993699cb3196f6aade0fc99a344d3ffda16ab4adea916236bed6e6af830742c586be9d03fdce57928197544f8feebaa5ddd8df5b389aae4cb88859ba78319ab8e3daae751cf7aee5d0cfad615ec5a71b7417d34ea82c3b0d7960b88b937fb9d0f5afc87a82361f8ad68b7951599b370c52c39b56e70c27ba11b59ab1db4;
    5'b01001 : xpb = 1024'h5c7be1af5d92f1837d547b193ffb404b5c4d3c115f86a4279f97cc042b700b2810da4bd01f7089132792d79323e8fb9971295a62e5b01d507f1c54a78e5e21ac2b965ae087bbd66e0ff275d4dc2f6916bbd715d6698714ac160a98b6fe47f15e38ce83183b420e10ad7cfa6529fa5384271ee6098c66da6b79357bc806f4e35;
    5'b01010 : xpb = 1024'h689387f84403dfdfcb4559593bc00c1608ffd09c561d96535bac46e8ca05b63c91376e86e4444fd41ed7721fd296373ea694f554f173206c159dfe6aa7029163e01671cd15a1264359a9f450398b9b67710e2511dc822523749d0d7b8e6ae785fa845331bba9922c3a76d8c2e57a5b00204cf6774822ca0cf31a89623015e521;
    5'b01011 : xpb = 1024'h1ab20c7fd0405bde93aff329d3261cd5eac4ca46c0cb21ecbf8257bb9e51bebe9e18bad7fc6b18886bd7777f8f8fcdf951fd2d1d91d86eb772aaf82c9a4ccbfb8924493d733591dabfbabea08c787c0c8259df2dc5e5abeb724cdf70f2c6ad63e2742c0842d60ae9e355fb008084ea9eaf4e1faba733c942e832400356da15a2;
    5'b01100 : xpb = 1024'h7d7dd65d1e6b0ca6272004d17ae674e73dffc72200f04dfda13521e425a07448ae4284a1deb85fcb5835bc262fe7757e617f8ccc54f08d4e8057314cc8697b44a681555c805afab738658b93784120e287aa92e23bcf5fc425894361114d15d3f96b97087acb7c3512f5041d135fa0668d2927c2569025a923b971a90680ac8e;
    5'b01101 : xpb = 1024'h2f9c5ae4aaa788a4ef8a9ea2124c85a71fc4c0cc6b9dd997050b32b6f9ec7ccabb23d0f2f6df287fa535c185ece10c390ce7c494f555db99dd642b0ebbb3b5dc4f8f2cccddef664e9e7655e3cb2e018798f64cfe2532e68c2339155675a8dbb1e15b6fdf01f7f4f2bbd4265aae6a30051c2a50f6b5a124df18d1284a2d44dd0f;
    5'b01110 : xpb = 1024'h926824c1f8d2396c82fab049ba0cddb872ffbda7abc305a7e6bdfcdf813b3254cb4d9abcd92c6fc29194062c8d38b3be1c6a2443b86dfa30eb10642ee9d065256cec38ebeb14cf2b172122d6b6f6a65d9e4700b29b1c9a64d6757946942f4421f852dadf39ed663deb732f774144e5ccfa05590d64fd8145545859efdceb73fb;
    5'b01111 : xpb = 1024'h4486a949850eb56b4b654a1a5172ee7854c4b752167091414a940db255873ad6d82ee70df1533876de940b8c4a324a78c7d25c0c58d3487c481d5df0dd1a9fbd15fa105c48a93ac27d31ed2709e38702af92bace8480212cd4254b3bf88b09ffe042b3b5c119defb945251b4dc4f756b89068241c40e807b4970109103afa47c;
    5'b10000 : xpb = 1024'ha7527326d3396632ded55bc1f9334689a7ffb42d5695bd522c46d7dadcd5f060e858b0d7d3a07fb9caf25032ea89f1fdd754bbbb1beb671355c997110b374f0633571c7b55cea39ef5dcba19f5ac2bd8b4e36e82fa69d5058761af2c1711726ff73a1eb5f90f5046c3f15ad16f2a2b3366e18a58736adce184f74236b3563b68;
    5'b10001 : xpb = 1024'h5970f7ae5f75e231a73ff5929099574989c4add7c14348eb901ce8adb121f8e2f539fd28ebc7486e17f25592a78388b882bcf383bc50b55eb2d690d2fe81899ddc64f3ebb3630f365bed846a48990c7dc62f289ee3cd5bcd851181217b6d384ddf29f78c803bc9046cd07d0f0a34bad1f5e2b38cd27bdc177a0ef8d7da1a6be9;
    5'b10010 : xpb = 1024'hb8f7c35ebb25e306faa8f6327ff68096b89a7822bf0d484f3f2f980856e0165021b497a03ee112264f25af2647d1f732e252b4c5cb603aa0fe38a94f1cbc4358572cb5c10f77acdc1fe4eba9b85ed22d77ae2bacd30e29582c15316dfc8fe2bc719d063076841c215af9f4ca53f4a7084e3dcc1318cdb4d6f26af7900de9c6a;
    5'b10011 : xpb = 1024'h6e5b461339dd0ef8031aa10acfbfc01abec4a45d6c160095d5a5c3a90cbcb6ef12451343e63b586551509f9904d4c6f83da78afb1fce22411d8fc3b51fe8737ea2cfd77b1e1ce3aa3aa91bad874e91f8dccb966f431a966e35fdb706fe4f669bde113b633f5db30d454ea869381a003862bee4d7e0e937b3aaade11eb0853356;
    5'b10100 : xpb = 1024'h2079ca9ac6198af6cb853adb6725d0daa0899e07d6c38c2f397bd47be108bf711f265f94fe6221199e50a4f8c1ce5db2e90fc2c3c033708c7a9cbd771332ae164bddaeeb7bb14f41a0b9e5fdda3b729dee17508b2c7e1d3633ad88fc62ab2c79c6011439c68a2bcaee2dcaa6d3248fd6f1c00e0c3ffa36e99fc597bfd74963d7;
    5'b10101 : xpb = 1024'h8345947814443bbe5ef54c830ee628ebf3c49ae316e8b8401b2e9ea4685774fb2f50295ee0af685c8aaee99f62260537f8922272834b8f238848f697414f5d5f693abb0a88d6b81e1964b2f0c6041773f368043fa267d10ee6e9ecec813194e9dcf87f39fe7f9d161dccd3c365ff459ecf9b1622ef56934fdb4cc96586effac3;
    5'b10110 : xpb = 1024'h356418ffa080b7bd275fe653a64c39abd589948d819643d97f04af773ca37d7d3c3175aff8d63110d7aeeeff1f1f9bf2a3fa5a3b23b0dd6ee555f059349997f71248927ae66b23b57f757d4118f0f81904b3be5b8bcb57d6e499bee1e58d5ac7c4e8581085ac15d3c6abf6010109d53d5e9c3f574e679285d0648006adb42b44;
    5'b10111 : xpb = 1024'h982fe2dceeab6884bacff7fb4e0c91bd28c49168c1bb6fea60b7799fc3f233074c5b3f79db237853c40d33a5bf774377b37cb9e9e6c8fc05f302297962b647402fa59e99f3908c91f8204a3404b99cef0a04721001b50baf97d622d20413c337dbdfc310bda1871ef64aff1d93e48b053c77476dfdc3eeec0bebb1ac5d5ac230;
    5'b11000 : xpb = 1024'h4a4e67647ae7e483833a91cbe572a27d0a898b132c68fb83c48d8a72983e3b89593c8bcaf34a4108110d39057c70da325ee4f1b2872e4a51500f233b560081d7d8b3760a5124f8295e31148457a67d941b502c2beb1892779585f4c7686f8915c3cf9be744cdffdc9f2a215b2eef1aa3cb7870a25cd4ee220103684d841ef2b1;
    5'b11001 : xpb = 1024'had1a3141c912954b16aaa3738d32fa8e5dc487ee6c8e2794a640549b1f8cf11369665594d597884afd6b7dac1cc881b76e6751614a4668e85dbb5c5b841d3120f61082295e4a6105d6dbe177436f226a20a0dfe06102465048c258b786f5f185dac706e77cc37127cec92a77c1c9d06ba95378b90c314a883c8a99f333c5899d;
    5'b11010 : xpb = 1024'h5f38b5c9554f1149df153d4424990b4e3f898198d73bb32e0a16656df3d8f9957647a1e5edbe50ff4a6b830bd9c2187219cf8929eaabb733bac8561d77676bb89f1e5999bbdecc9d3cecabc7965c030f31ec99fc4a65cd1846722aaceb51b763c2b6dfbe03efe9e577a84cb55cd4600a3854a1ed6b4249be31a250945a89ba1e;
    5'b11011 : xpb = 1024'h11573a50e18b8d48a77fd714bbff1c0e214e7b4341e93ec76dec7640c82502178328ee3705e519b3976b886b96bbaf2cc537c0f28b11057f17d54fdf6ab1a650482c310a19733834a2fd7617e948e3b44338541833c953e04421fca24fad7d41aaa6b8948b1c62a320876ef2f7deefa8c755cb21ca5348f426ba0735814dea9f;
    5'b11100 : xpb = 1024'h7423042e2fb63e103aefe8bc63bf741f7489781e820e6ad84f9f40694f73b7a19352b800e83260f683c9cd12371356b1d4ba20a14e292416258188ff98ce559965893d292698a1111ba8430ad511888a488907cca9b307b8f75e60926e33e5b1c19e2394c311d3ee5026780f8ab9a570a530d33879afa55a624138db30f4818b;
    5'b11101 : xpb = 1024'h264188b5bbf2ba0f035a828cfb2584df564e71c8ecbbf671b375513c23bfc023a0340452005929aad0c9d271f40ced6c80225869ee8e7261828e82c18c1890310e971499842d0ca881b90d5b27fe692f59d4c1e893168e80f50e3287d28fab8fa98dfc6b4a3e4cabf9059a4d25c4350f3431fc6cd8c0a4905758ef7c57b8b20c;
    5'b11110 : xpb = 1024'h890d52930a1d6ad696ca9434a2e5dcf0a9896ea42ce1228295281b64ab0e75adb05dce1be2a670edbd281718946494f18fa4b818b1a690f8903abbe1ba353f7a2bf420b891527584fa63da4e13c70e055f25759d09004259a84a9677f11613ffc085676b8233bdf728a4a369b89eead7120d0483881d00f692e02122075f48f8;
    5'b11111 : xpb = 1024'h3b2bd71a9659e6d55f352e053a4bedb08b4e684e978eae1bf8fe2c377f5a7e2fbd3f1a6cfacd39a20a281c78515e2bac3b0cefe1520bdf43ed47b5a3ad7f7a11d501f828eee6e11c6074a49e66b3eeaa70712fb8f263c921a5fa686d5571d9dda8754042096036b4d183c5a753a97a75a10e2db7e72e002c87f7d7c32e237979;
    endcase
end

endmodule

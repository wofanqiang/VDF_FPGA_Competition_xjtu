module xpb_5_705
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h2883a3d7880c9b38689410f62003893b8d3b01485cca24c1ad843a36526eb6ace3e717231c2b3ebb3c18ff5a73e8aff5cb4ff1b24a64cd6366137d431b489dda7ae8f1c56cdeb393bf5e3fd49426988ab7bdd9b84d420739719544329ca19fe244ed641fcca437171f2b396f39d23825423ea8bab978a4fd221f13f8555737fd;
    5'b00010 : xpb = 1024'h510747af10193670d12821ec400712771a760290b99449835b08746ca4dd6d59c7ce2e4638567d767831feb4e7d15feb969fe36494c99ac6cc26fa8636913bb4f5d1e38ad9bd67277ebc7fa9284d31156f7bb3709a840e72e32a886539433fc489dac83f99486e2e3e5672de73a4704a847d517572f149fa443e27f0aaae6ffa;
    5'b00011 : xpb = 1024'h798aeb869825d1a939bc32e2600a9bb2a7b103d9165e6e45088caea2f74c2406abb545695481bc31b44afe0f5bba0fe161efd516df2e682a323a77c951d9d98f70bad550469c1abb3e1abf7dbc73c9a027398d28e7c615ac54bfcc97d5e4dfa6cec82c5f65eca5455d81ac4dad76a86fc6bbfa302c69eef7665d3be90005a7f7;
    5'b00100 : xpb = 1024'ha20e8f5e20326ce1a25043d8800e24ee34ec052173289306b610e8d949badab38f9c5c8c70acfaecf063fd69cfa2bfd72d3fc6c92993358d984df50c6d227769eba3c715b37ace4efd78ff52509a622adef766e135081ce5c65510ca72867f8913b5907f3290dc5c7cace5bce748e09508faa2eae5e293f4887c4fe1555cdff4;
    5'b00101 : xpb = 1024'h19e4eddfe650d3513fdedcf78fb766d850b10338fa7b1750e5b869b9e926e458703af636c2b1bb198d1ebd7d602d5f0294759095514532a54dc232f14d98a092f23d842c70c8849daa3d3c844be53684a2b04700f5c3f70e825dc30254fd7cd9299b62754e6c1ae61518384d294af290fc5f6cc34f0fdbc1642be8d521d1b186;
    5'b00110 : xpb = 1024'h426891b76e5d6e89a872ededafbaf013ddec048157453c12933ca3f03b959b0554220d59dedcf9d4c937bcd7d4160ef85fc582479baa0008b3d5b03468e13e6d6d2675f1dda73831699b7c58e00bcf0f5a6e20b94305fe47f3f30734f19f1cbb6e88c6951b1051fd344371bc631d2ab63e9e157e088880be864afccd7728e983;
    5'b00111 : xpb = 1024'h6aec358ef66a09c21106fee3cfbe794f6b2705c9b40f60d440c0de268e0451b23809247cfb0838900550bc3247febeee2b1573f9e60ecd6c19e92d778429dc47e80f67b74a85ebc528f9bc2d7432679a122bfa719048058165884b678e40bc9db3762ab4e7b48914536eab2b9cef62db80dcbe38c20125bba86a10c5cc802180;
    5'b01000 : xpb = 1024'h936fd9667e76a4fa799b0fd9efc2028af862071210d98595ee45185ce073085f1bf03ba01733774b4169bb8cbbe76ee3f66565ac30739acf7ffcaaba9f727a2262f8597cb7649f58e857fc0208590024c9e9d429dd8a0cbad71d8f9a2ae25c7ff8638ed4b458c02b7299e49ad6c19b00c31b66f37b79cab8ca8924be21d7597d;
    5'b01001 : xpb = 1024'hb4637e844950b6a1729a8f8ff6b447514270529982c09e01dec993d7fdf1203fc8ed54a69383777de247ba04c720e0f5d9b2f78582597e73570e89f7fe8a34b6992169374b255a7951c393403a3d47e8da2b4499e45e6e3932641d20d5959d00e4960cad033feb50b05372b18c3acfcb68030cbe4a71285a638bdb1ee4c2b0f;
    5'b01010 : xpb = 1024'h33c9dbbfcca1a6a27fbdb9ef1f6ecdb0a1620671f4f62ea1cb70d373d24dc8b0e075ec6d856376331a3d7afac05abe0528eb212aa28a654a9b8465e29b314125e47b0858e191093b547a790897ca6d0945608e01eb87ee1d04bb8604a9faf9b25336c4ea9cd835cc2a30709a5295e521f8bed9869e1fb782c857d1aa43a3630c;
    5'b01011 : xpb = 1024'h5c4d7f9754ae41dae851cae53f7256ec2e9d07ba51c0536378f50daa24bc7f5dc45d0390a18eb4ee56567a5534436dfaf43b12dcecef32ae0197e325b679df005f63fa1e4e6fbccf13d8b8dd2bf10593fd1e67ba38c9f5567650ca37469c99949824290a697c6ce3495baa098c681d473afd824157985c7fea76e5a298fa9b09;
    5'b01100 : xpb = 1024'h84d1236edcbadd1350e5dbdb5f75e027bbd80902ae8a7825267947e0772b360aa8441ab3bdb9f3a9926f79afa82c1df0bf8b048f3754001167ab6068d1c27cdada4cebe3bb4e7062d336f8b1c0179e1eb4dc4172860bfc8fe7e60e69e33e3976dd118d2a3620a3fa6886e378c63a556c7d3c2afc1111017d0c95f99aee51d306;
    5'b01101 : xpb = 1024'had54c74664c7784bb979ecd17f79696349130a4b0b549ce6d3fd8216c999ecb78c2b31d6d9e53264ce88790a1c14cde68adaf64181b8cd74cdbeddabed0b1ab55535dda9282d23f692953886543e36a96c9a1b2ad34e03c9597b529c7fdfd95921fef14a02c4db1187b21ce8000c8d91bf7ad3b6ca89a67a2eb50d9343a90b03;
    5'b01110 : xpb = 1024'h252b25c82ae5debb570885f08f22ab4d64d8086292a7213103a502f76905f65c6cc9cb812be9f2916b43391dac9f6d11f210c00da96aca8c83331b90cd8143de5bcf9abfe57ada453f5975b84f890b033052fb4a9409ddf2158404d46256d6a937e4c3401ea0199b201d6f78420e9f8db2df9d8f33b6ee470a64a687101ddc95;
    5'b01111 : xpb = 1024'h4daec99fb2f279f3bf9c96e6af263488f21309aaef7145f2b1293d2dbb74ad0950b0e2a44815314ca75c387820881d07bd60b1bff3cf97efe94698d3e8c9e1b8d6b88c8552598dd8feb7b58ce3afa38de810d502e14be52b87194906fef8768b7cd2275feb4450b23f48a8e77be0d7b2f51e4649ed2f93442c83ba7f65751492;
    5'b10000 : xpb = 1024'h76326d773aff152c2830a7dccf29bdc47f4e0af34c3b6ab45ead77640de363b63497f9c764407007e37537d29470ccfd88b0a3723e3465534f5a161704127f9351a17e4abf38416cbe15f56177d63c189fceaebb2e8dec64f8ae8d399b9a166dc1bf8b7fb7e887c95e73e256b5b30fd8375cef04a6a838414ea2ce77bacc4c8f;
    5'b10001 : xpb = 1024'h9eb6114ec30bb06490c4b8d2ef2d47000c890c3ba9058f760c31b19a60521a63187f10ea806baec31f8e372d08597cf354009524889932b6b56d935a1f5b1d6dcc8a70102c16f5007d7435360bfcd4a3578c88737bcff39e6a43d16c383bb65006acef9f848cbee07d9f1bc5ef8547fd799b97bf6020dd3e70c1e2701023848c;
    5'b10010 : xpb = 1024'h168c6fd0892a16d42e5351f1fed688ea284e0a53305813c03bd9327affbe2407f91daa94d2706eefbc48f74098e41c1ebb365ef0b04b2fce6ae1d13effd14696d3242d26e964ab4f2a3872680747a8fd1b4568933c8bcdc7264c83a41ab2b3a01c92c195a067fd6a160a6e56318759f96d006197c94e250b4c717b63dc98561e;
    5'b10011 : xpb = 1024'h3f1013a81136b20c96e762e81eda1225b5890b9b8d223881e95d6cb1522cdab4dd04c1b7ee9badaaf861f69b0ccccc14868650a2faaffd31d0f54e821b19e4714e0d1eec56435ee2e996b23c9b6e4187d303424b89cdd50097e1c7d6b7545382618025b56d0c34813535a7c56b59921eaf3f0a5282c6ca086e908f5c31ef8e1b;
    5'b10100 : xpb = 1024'h6793b77f99434d44ff7b73de3edd9b6142c40ce3e9ec5d4396e1a6e7a49b9161c0ebd8db0ac6ec66347af5f580b57c0a51d642554514ca953708cbc53662824bc8f610b1c3221276a8f4f2112f94da128ac11c03d70fdc3a09770c0953f5f364a66d89d539b06b985460e134a52bca43f17db30d3c3f6f0590afa3548746c618;
    5'b10101 : xpb = 1024'h90175b57214fe87d680f84d45ee1249ccfff0e2c46b682054465e11df70a480ea4d2effe26f22b217093f54ff49e2c001d2634078f7997f89d1c490851ab202643df02773000c60a685331e5c3bb729d427ef5bc2451e3737b0c503bf0979346eb5aedf50654a2af738c1aa3defe026933bc5bc7f5b81402b2ceb74cdc9dfe15;
    5'b10110 : xpb = 1024'h7edb9d8e76e4eed059e1df36e8a6686ebc40c43ce09064f740d61fe967651b3857189a878f6eb4e0d4eb5638528cb2b845bfdd3b72b9510529086ed3221494f4a78bf8ded4e7c5915176f17bf0646f70637d5dbe50dbd9c37150273d30e90970140bfeb222fe1390bf76d3421001465272125a05ee55bcf8e7e5040a912cfa7;
    5'b10111 : xpb = 1024'h30715db06f7aea256e322ee98e8defc278ff0d8c2ad32b1121919c34e8e508606958a0cb95222a094967b4bdf9117b214fabef8601906273b8a404304d69e729c561b1535a2d2fecd475aeec532cdf81bdf5af94324fc4d5a8aa46a66fb03079462e240aeed418502b22a6a35ad24c8a695fce5b185e00ccb09d6438fe6a07a4;
    5'b11000 : xpb = 1024'h58f50187f787855dd6c63fdfae9178fe063a0ed4879d4fd2cf15d66b3b53bf0d4d3fb7eeb14d68c48580b4186cfa2b171afbe1384bf52fd71eb7817368b28504404aa318c70be38093d3eec0e753780c75b3894c7f91cc0f1a3f8ad90c51d05b8b1b882abb784f674a4de01294a484afab9e7715d1d6a5c9d2bc783153c13fa1;
    5'b11001 : xpb = 1024'h8178a55f7f9420963f5a50d5ce9502399375101ce46774947c9a10a18dc275ba3126cf11cd78a77fc199b372e0e2db0ce64bd2ea9659fd3a84cafeb683fb22debb3394de33ea971453322e957b7a10972d716304ccd3d3488bd4cf0ba8f3703dd008ec4a881c867e69791981ce76bcd4eddd1fd08b4f4ac6f4db8c29a918779e;
    5'b11010 : xpb = 1024'ha9fc493707a0bbcea7ee61cbee988b7520b01165413199562a1e4ad7e0312c67150de634e9a3e63afdb2b2cd54cb8b02b19bc49ce0beca9deade7bf99f43c0b9361c86a3a0c94aa812906e6a0fa0a921e52f3cbd1a15da81fd6a133e4595102014f6506a54c0bd9588a452f10848f4fa301bc88b44c7efc416faa021fe6faf9b;
    5'b11011 : xpb = 1024'h21d2a7b8cdbf223e457cfaeafe41cd5f3c750f7cc8841da059c5cbb87f9d360bf5ac7fdf3ba8a6679a6d72e0e5562a2e18d18e690870c7b5a052b9de7fb9e9e23cb643ba5e1700f6bf54ab9c0aeb7d7ba8e81cdcdad1b4aab972c576280c0d702adc2260709bfc1f210fa5814a4b06f623809263adf53790f2aa3915cae4812d;
    5'b11100 : xpb = 1024'h4a564b9055cbbd76ae110be11e45569ac9b010c5254e4262074a05eed20becb8d993970257d3e522d686723b593eda23e421801b52d59519066637219b0287bcb79f357fcaf5b48a7eb2eb709f12160660a5f6952813bbe42b0809a8c4adad526fc986803d403336403adef0841d3f1b65bf3b1e676ddc8e14c94d0e203bb92a;
    5'b11101 : xpb = 1024'h72d9ef67ddd858af16a51cd73e48dfd656eb120d82186723b4ce4025247aa365bd7aae2573ff23de129f7195cd278a19af7171cd9d3a627c6c79b464b64b25973288274537d4681e3e112b453338ae911863d04d7555c31d9c9d4ddb614f4d34b4b6eaa009e46a4d5f66185fbdef7740a7fde3d920e6818b36e861067592f127;
    5'b11110 : xpb = 1024'h9b5d933f65e4f3e77f392dcd5e4c6911e4261355dee28be562527a5b76e95a12a161c548902a62994eb870f041103a0f7ac1637fe79f2fdfd28d31a7d193c371ad71190aa4b31bb1fd6f6b19c75f471bd021aa05c297ca570e32920dfdf0ed16f9a44ebfd688a1647e9151cef7c1af65ea3c8c93da5f2688590774fecaea2924;
    5'b11111 : xpb = 1024'h1333f1c12c035a571cc7c6ec6df5aafbffeb116d6635102f91f9fb3c165563b782005ef2e22f22c5eb733103d19ad93ae1f72d4c0f512cf788016f8cb209ec9ab40ad6216200d200aa33a84bc2aa1b7593da8a258353a47fca3b4445e067ea670f8a20b5f263dfee16fca45f39c3c161dda1566c438c6e5534b70df2975efab6;
    endcase
end

endmodule

module xpb_5_305
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h47301f868befce7d9048c23c1a62806967d62b9d34433850753b8a51fc2e3d7ad64d8fb264b5d4042f2613f0ac61d56dbc6b9ff41d13e138196b1c34216768c7ce8f881b5951510a4f46cc6fca63add7168d76a7fd7926b6512b4bbb97d916724169c8afd16ba032c56eb0c518c6e0633d85d40a017270731c2964f0cf231cd1;
    5'b00010 : xpb = 1024'h8e603f0d17df9cfb2091847834c500d2cfac573a688670a0ea7714a3f85c7af5ac9b1f64c96ba8085e4c27e158c3aadb78d73fe83a27c27032d6386842ced18f9d1f1036b2a2a2149e8d98df94c75bae2d1aed4ffaf24d6ca25697772fb22ce482d3915fa2d740658add618a318dc0c67b0ba81402e4e0e63852c9e19e4639a2;
    5'b00011 : xpb = 1024'h24e3193de1e136afe5d4cedd3ecd39eac60c7fa6c7520879e1d5e5a041880b687fa0319e63fafd7dee13fc8b21c76f7ed128b7f63488d35c9ba2153e2963c5a5f75f63a35c62f5d9db3a62acc64f45544fa36a5f6be547123df551380d60a0c49535c7e5c379e80ac98c2b7052847b0069b79d3bb40bf4290e0cb3cde486f008;
    5'b00100 : xpb = 1024'h6c1338c46dd1052d761d9119592fba542de2ab43fb9540ca57116ff23db648e355edc150c8b0d1821d3a107bce2944ec8d9457ea519cb494b50d31724acb2e6dc5eeebbeb5b446e42a812f1c90b2f32b6630e107695e6dc88f209cf3a539b736d69f909594e5883d8efadc356b4b5b63a73d7145b57e649c2a3618beb3aa0cd9;
    5'b00101 : xpb = 1024'h29612f537d29ee23b60db7e6337f36c2442d3b05a60d8a34e7040ee86e1d95628f2d38a634026f7ad01e525972d098fe5e5cff84bfdc5811dd90e4831602284202f3f2b5f749aa9672df8e9c23adcd188b95e16da51676e2abf56b482e82b16e901c71bb5882fe2cda9a61b8c42159d95e9666d66a577defff002aaf9eac33f;
    5'b00110 : xpb = 1024'h49c6327bc3c26d5fcba99dba7d9a73d58c18ff4d8ea410f3c3abcb40831016d0ff40633cc7f5fafbdc27f916438edefda2516fec6911a6b937442a7c52c78b4beebec746b8c5ebb3b674c5598c9e8aa89f46d4bed7ca8e247beaa2701ac141892a6b8fcb86f3d015931856e0a508f600d36f3a776817e8521c19679bc90de010;
    5'b00111 : xpb = 1024'h90f652024fb23bdd5bf25ff697fcf43ef3ef2aeac2e7494438e755927f3e544bd58df2ef2cabcf000b4e0d06eff0b46b5ebd0fe0862587f150af46b0742ef413bd4e4f6212173cbe05bb91c95702387fb5d44b66d543b4dacd15ee2bb29a57fb6bd5587b585f7048588707a5bdcfd66410f50e81698a58c53842cc8c9830fce1;
    5'b01000 : xpb = 1024'h27792c3319b3d5922135aa5ba2052d56ea4f535721b2e11d3046268ec869e4bea8930528c73b24759b15e1b0b8f4790eb70e87ee808698ddb97b23865ac3e82a178ea2cebbd7908342685b96888a2225d85cc8764636ae8068b4a7ec9048cbdb7e378f01790217ed9735d18bdec6909dffa103a91ab16c080dfcb678de71b347;
    5'b01001 : xpb = 1024'h6ea94bb9a5a3a40fb17e6c97bc67adc052257ef455f6196da581b0e0c49822397ee094db2bf0f879ca3bf5a165564e7c737a27e29d9a7a15d2e63fba7c2b50f1e61e2aea1528e18d91af280652edcffceeea3f1e43afd536b9dff3a82821e24dbfa157b14a6db8205ca48250f78d71013d26d7b31c23dc7b2a261b69ad94d018;
    5'b01010 : xpb = 1024'h52c25ea6fa53dc476c1b6fcc66fe6d84885a760b4c1b1469ce081dd0dc3b2ac51e5a714c6804def5a03ca4b2e5a131fcbcb9ff097fb8b023bb21c9062c04508405e7e56bee93552ce5bf1d38475b9a31172bc2db4a2cedc557ead6905d0562dd2038e376b105fc59b534c3718842b3b2bd2ccdacd4aefbdffe00555f3d5867e;
    5'b01011 : xpb = 1024'h4c5c4570fb950c42070a7938e0d26741b05bd2fde904e997121c0c2f09f1f027283336c72b3621f38929de3bdabbe88d88373fe4b50f6c3a551d38c48427add00eee0672183a865d1da2be434ed9677a280032d5b21bf592a6a9f9249da96ca0136d56e73c7bfff860c1fcfc314b0b9e6958a0e4cebd60311c096a46c2f8a34f;
    5'b01100 : xpb = 1024'h938c64f78784dabf97533b74fb34e7ab1831fe9b1d4821e78757968106202da1fe80c6798febf5f7b84ff22c871dbdfb44a2dfd8d2234d726e8854f8a58f1697dd7d8e8d718bd7676ce98ab3193d15513e8da97daf951c48f7d544e03582831254d71f970de7a02b2630adc14a11ec01a6de74eed02fd0a43832cf37921bc020;
    5'b01101 : xpb = 1024'h2a0f3f28518674745c9685da053d20c30e9227077c13b9c07eb6677d4f4bbe14d185d8b32a7b4b6d4817c6d65021829e9cf457e6cc845e5ed75431ce8c240aae37bde1fa1b4c2b2ca99654804ac4fef76116268d208815ee9373fea11330f6f26739561d2e8a47d064df77a76b08a63b958a6a168156e3e70decb923d85c7686;
    5'b01110 : xpb = 1024'h713f5eaedd7642f1ecdf48161f9fa12c766852a4b056f210f3f1f1cf4b79fb8fa7d368658f311f71773ddac6fc83580c595ff7dae9983f96f0bf4e02ad8b7376064d6a15749d7c36f8dd20f01528acce77a39d351e013ca4e49f4a5cab0a0d64a8a31eccfff5e8032a4e286c83cf869ed3103e2082c9545a2a161e14a77f9357;
    5'b01111 : xpb = 1024'h7c238dfa777dca6b222927b29a7da446cc87b110f2289e9eb50c2cb94a58c027ad87a9f29c074e70705af70c5871cafb1b16fe8e3f95083598b2ad89420678c608dbd821e5dcffc3589eabd46b096749a2c1a448ef4364a803e041d88b88144bb05555320988fa868fcf252a4c640d8c1bc334833f0679cffd00800edc049bd;
    5'b10000 : xpb = 1024'h4ef258663367ab24426b54b7440a5aadd49ea6ae4365c23a608c4d1d90d3c97d51260a518e7648eb362bc36171e8f21d6e1d0fdd010d31bb72f6470cb587d0542f1d459d77af210684d0b72d1114444bb0b990ec8c6d5d00d1694fd9209197b6fc6f1e02f2042fdb2e6ba317bd8d213bff4207523562d8101bf96cf1bce3668e;
    5'b10001 : xpb = 1024'h962277ecbf5779a1d2b416f35e6cdb173c74d24b77a8fa8ad5c7d76f8d0206f827739a03f32c1cef6551d7521e4ac78b2a88afd11e2112f38c616340d6ef391bfdaccdb8d1007210d417839cdb77f222c747079489e683b722949b94b86aae293dd8e6b2c36fd00df3da53dcd654019f3cc7db5c36d548833822d1e28c06835f;
    5'b10010 : xpb = 1024'h2ca5521d8959135697f761586875142f32d4fab7d6749263cd26a86bd62d976afa78ac3d8dbb7264f519abfbe74e8c2e82da27df188223dff52d4016bd842d3257ed21257ac0c5d610c44d6a0cffdbc8e9cf84a3fad97d5cbe33555596192209503b1d38e41277b332891dc2f74abbd92b73d083e7fc5bc60ddcbbced24739c5;
    5'b10011 : xpb = 1024'h73d571a41548e1d42840239482d794989aab26550ab7cab4426232bdd25bd4e5d0c63beff2714669243fbfec93b0619c3f45c7d3359605180e985c4adeeb95fa267ca940d41216e0600b19d9d76389a0005cfb4bf852a4130f5ea1112df2387b91a4e5e8b57e17e5f7f7ce8810119c3c68f9a48de96ecc392a0620bfa16a5696;
    5'b10100 : xpb = 1024'ha584bd4df4a7b88ed836df98cdfcdb0910b4ec16983628d39c103ba1b876558a3cb4e298d009bdeb40794965cb4263f97973fe12ff7160477643920c5808a1080bcfcad7dd26aa59cb7e3a708eb734622e5785b69459db8aafd5ad20ba0ac5ba4071c6ed620bf8b36a6986e3108567657a599b59a95df7bffc00aabe7ab0cfc;
    5'b10101 : xpb = 1024'h51886b5b6b3a4a067dcc3035a7424e19f8e17a5e9dc69addaefc8e0c17b5a2d37a18dddbf1b66fe2e32da8870915fbad5402dfd54d0af73c90cf5554e6e7f2d84f4c84c8d723bbafebfeb016d34f211d3972ef0366bec46efc28a68da379c2cde570e51ea78c5fbdfc15493349cf36d9952b6dbf9c084fef1be96f9cb6ce29cd;
    5'b10110 : xpb = 1024'h98b88ae1f72a18840e14f271c1a4ce8360b7a5fbd209d32e2438185e13e3e04e50666d8e566c43e71253bc77b577d11b106e7fc96a1ed874aa3a7189084f5ba01ddc0ce430750cba3b457c869db2cef4500065ab6437eb254d53f2493b52d94026daadce78f7fff0c183f9f86296173cd2b141c99d7ac0623812d48d85f1469e;
    5'b10111 : xpb = 1024'h2f3b6512c12bb238d3583cd6cbad079b5717ce6830d56b071b96e95a5d0f70c1236b7fc7f0fb995ca21b91217e7b95be68bff7d7647fe96113064e5eeee44fb6781c6050da35607f77f24653cf3ab89a7288e2bad52ae4cae8f2ac0a19014d20393ce454999aa7960032c3de838cd176c15d36f14ea1d3a50dccbe79cc31fd04;
    5'b11000 : xpb = 1024'h766b84994d1b80b663a0ff12e60f8804beedfa056518a35790d273ac593dae3bf9b90f7a55b16d60d141a5122add6b2c252b97cb8193ca992c716a93104bb87e46abe86c3386b189c73912c3999e667189165962d2a40b813a1df7c5b0da63927aa6ad046b0647c8c5a174a39c53b1d9fee30afb5014441829f6236a9b5519d5;
    5'b11001 : xpb = 1024'hcee5eca171d1a6b28e44977f017c11cb54e2271c3e43b30883144a8a2693eaeccbe21b3f040c2d6610979bbf3e12fcf7d7d0fd97bf4db85953d4768f6e0ac94a0ec3bd8dd47054f03e5dc90cb265017ab9ed67243970526d5bcb1868e88d7728d08e38a8ba8ef6e04503e89bd4a6c13ed8f0023013b575affb00d56e195d03b;
    5'b11010 : xpb = 1024'h541e7e50a30ce8e8b92d0bb40a7a41861d244e0ef8277380fd6ccefa9e977c29a30bb16654f696da902f8daca043053d39e8afcd9908bcbdaea8639d1848155c6f7bc3f436985659532ca9009589fdeec22c4d1a41102bdd26e7fd422661ede4ce72ac3a5d148fa0c9beef4ed6114c772b14d42d02adc7ce1bd97247b0b8ed0c;
    5'b11011 : xpb = 1024'h9b4e9dd72efcb7664975cdf024dcc1ef84fa79ac2c6aabd172a8594c9ac5b9a479594118b9ac6adebf55a19d4ca4daaaf6544fc1b61c9df5c8137fd139af7e243e0b4c0f8fe9a763a27375705fedabc5d8b9c3c23e895293781348fdbe3b04570fdc74ea2e802fd38f2da013eed82cda689aa837042038413802d7387fdc09dd;
    5'b11100 : xpb = 1024'h31d17807f8fe511b0eb918552ee4fb077b5aa2188b3643aa6a072a48e3f14a174c5e5352543bc0544f1d764715a89f4e4ea5c7cfb07daee230df5ca72044723a984b9f7c39a9fb28df203f3d9175956bfb4240d1af7c4c3913b202be9be97837223eab704f22d778cddc69fa0fcee71457469d5eb5474b840dbcc124c61cc043;
    5'b11101 : xpb = 1024'h7901978e84ee1f989f01da9149477b70e330cdb5bf797bfadf42b49ae01f879222abe304b8f194587e438a37c20a74bc0b1167c3cd91901a4a4a78db41abdb0266db279792fb4c332e670bad5bd9434311cfb779acf572ef64dd4e7a33c28ea963a87420208e77ab934b1abf2895c77794cc7168b6b9bbf729e62615953fdd14;
    5'b11110 : xpb = 1024'hf8471bf4eefb94d644524f6534fb488d990f6221e4513d3d6a18597294b1804f5b0f53e5380e9ce0e0b5ee18b0e395f6362dfd1c7f2a106b31655b12840cf18c11b7b043cbb9ff86b13d57a8d612ce9345834891de86c95007c083b11710289760aaaa641311f50d1f9e4a5498c81b18378669067e0cf39ffa01001db80937a;
    5'b11111 : xpb = 1024'h56b49145dadf87caf48de7326db234f2416721bf52884c244bdd0fe92579557fcbfe84f0b836bdd23d3172d237700ecd1fce7fc5e506823ecc8171e549a837e08fab031f960cf102ba5aa1ea57c4dac04ae5ab311b61934b51a753f6a94a18fbb7747356129cbf839768956a62536214c0fe3a9a69533fad1bc974f2aaa3b04b;
    endcase
end

endmodule

module xpb_5_970
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h56d9116dbc9a08d6e42d3ac9abea1b8092d18a894855a9b7e3ebe8917773e4aee040ab63dd8eed430a871832514087dafa286377d9e9cd16a47bf0d137fe556fac659213d8453d1e2f5b0343b1746758a4f8ef164212402c6efbf11bace1511c7b2ae78239720ef73624cb88cb8e9fc2464c961befcdb4985782036f24d84f4e;
    5'b00010 : xpb = 1024'hadb222db793411adc85a759357d4370125a3151290ab536fc7d7d122eee7c95dc08156c7bb1dda86150e3064a2810fb5f450c6efb3d39a2d48f7e1a26ffcaadf58cb2427b08a7a3c5eb6068762e8ceb149f1de2c84248058ddf7e23759c2a238f655cf0472e41dee6c499711971d3f848c992c37df9b6930af0406de49b09e9c;
    5'b00011 : xpb = 1024'h53ddeef373dfe5bbe1823885f3640b3046fe9c6b03895cb02de7005eb35901049d7984b2ce86493a80370950106386c68a5f02816b0a96f83cd493156d288b9d90e1818cd93eba157b7707287b8171d8fae5d3aa39b09374976741584c7950c34279245cfb8d34581bae7bbb6adbb91d840be3717f1dc098c0168f48e5a6877f;
    5'b00100 : xpb = 1024'haab700613079ee92c5af734f9f4e26b0d9d026f44bdf066811d2e8f02acce5b37dba3016ac15367d8abe218261a40ea1848765f944f4640ee15083e6a526e10d3d4713a0b183f733aad20a6c2cf5d9319fdec2c07bc2d3a106633273f95aa1dfbda40bdf34ff434f51d34744366a58dfca58798d6eeb7531179892b80a7ed6cd;
    5'b00101 : xpb = 1024'h50e2cc792b25c2a0ded736423addfadffb2bae4cbebd0fa877e2182bef3e1d5a5ab25e01bf7da531f5e6fa6dcf8685b21a95a18afc2b60d9d52d3559a252c1cb755d7105da38370cc7930b0d458e7c5950d2b83e314ee6bcbfd29194ec11506a09c76137bda859b901382bee0a28d278c1cb30c70e6dcc9928ab1b22a674bfb0;
    5'b00110 : xpb = 1024'ha7bbdde6e7bfcb77c304710be6c816608dfd38d60712b9605bce00bd66b202093af309659d0c9275006e12a020c70d8d14be0502d6152df079a9262ada51173b21c30319b27d742af6ee0e50f702e3b1f5cba754736126e92ece82b098f2a18684f248b9f71a68b0375cf776d5b7723b0817c6e2fe3b8131802d1e91cb4d0efe;
    5'b00111 : xpb = 1024'h4de7a9fee26b9f85dc2c33fe8257ea8faf58c02e79f0c2a0c1dd2ff92b2339b017eb3750b07501296b96eb8b8ea9849daacc40948d4c2abb6d85d79dd77cf7f959d9607edb31b40413af0ef20f9b86d9a6bf9cd228ed3a04e83de1d18ba95010d1159e127fc37f19e6c1dc20a975ebd3ff8a7e1c9dbdd899913fa6fc6742f7e1;
    5'b01000 : xpb = 1024'ha4c0bb6c9f05a85cc0596ec82e420610422a4ab7c2466c58a5c9188aa2971e5ef82be2b48e03ee6c761e03bddfea0c78a4f4a40c6735f7d21201c86f0f7b4d69063ef292b376f122430a1235c10fee324bb88be86aff7a315739d2ed388aa12d4c408594b9358e111ce6a7a975048b9645d714388d8b8d31e8c1aa6b8c1b472f;
    5'b01001 : xpb = 1024'h4aec878499b17c6ad98131bac9d1da3f6385d210352475990bd847c667085605d524109fa16c5d20e146dca94dcc83893b02df9e1e6cf49d05de79e20ca72e273e554ff7dc2b30fb5fcb12d6d9a89159fcac8166208b8d4d10a9320e2b414fb79863daed41dea47acc4b8c5348c3052f3d49cb722d0de499f9d432d628113012;
    5'b01010 : xpb = 1024'ha1c598f2564b8541bdae6c8475bbf5bff6575c997d7a1f50efc43057de7c3ab4b564bc037efb4a63ebcdf4db9f0d0b64352b4315f856c1b3aa5a6ab344a58396eabae20bb4706e198f26161a8b1cf8b2a1a5707c629dcd797fa52329d822a0d4138ec26f7b50b372027057dc1451a4f18396618e1cdb9932515636454ce97f60;
    5'b01011 : xpb = 1024'h47f1650a50f7594fd6d62f77114bc9ef17b2e3f1f058289155d35f93a2ed725b925ce9ee9263b91856f6cdc70cef8274cb397ea7af8dbe7e9e371c2641d1645522d13f70dd24adf2abe716bba3b59bda529965fa1829e0953914824acad94f5e5fb217c803f9c9dbb1d53c85e8101e8a7b0918c7bc5df09a6268beafe8df6843;
    5'b01100 : xpb = 1024'h9eca76780d916226bb036a40bd35e56faa846e7b38add24939bf48251a61570a729d95526ff2a65b617de5f95e300a4fc561e21f89778b9542b30cf779cfb9c4cf36d184b569eb10db4219ff552a0332f79255105a3c20c1a810736677baa07adadcff4a3d6bd8d2e7fa080eb39ebe4cc155aee3ac2ba532b9eac21f0db7b791;
    5'b01101 : xpb = 1024'h44f64290083d3634d42b2d3358c5b99ecbdff5d3ab8bdb899fce7760ded28eb14f95c33d835b150fcca6bee4cc1281605b701db140ae8860368fbe6a76fb9a83074d2ee9de1e2ae9f8031aa06dc2a65aa8864a8e0fc833dd617fd2876a714f05270054a2c614ef3c975eecb8875d37e5b8c8661d4badfc9acafd4a89a9ada074;
    5'b01110 : xpb = 1024'h9bcf53fdc4d73f0bb85867fd04afd51f5eb1805cf3e1854183ba5ff2564673602fd66ea160ea0252d72dd7171d53093b559881291a985576db0baf3baef9eff2b3b2c0fdb6636808275e1de41f370db34d7f39a451da7409d07bc3a31752a021a22b3c24ff86fe33cd83b84152ebd7a7ff14fc393b7bb133227f4df8ce85efc2;
    5'b01111 : xpb = 1024'h41fb2015bf831319d1802aefa03fa94e800d07b566bf8e81e9c98f2e1ab7ab070cce9c8c745271074256b0028b35804beba6bcbad1cf5241cee860aeac25d0b0ebc91e62df17a7e1441f1e8537cfb0dafe732f220766872589eb22c40a094eabee4e917d8830149d7ce89ceb26aa5140f687b372dafe089b3391d6636a7bd8a5;
    5'b10000 : xpb = 1024'h98d431837c1d1bf0b5ad65b94c29c4cf12de923eaf153839cdb577bf922b8fb5ed0f47f051e15e4a4cddc834dc760826e5cf2032abb91f587364517fe4242620982eb076b75ce4ff737a21c8e9441833a36c1e384978c751f8e713dfb6ea9fc8697978ffc1a22394b30d6873f238f1033cd4498ecacbbd338b13d9d28f5427f3;
    5'b10001 : xpb = 1024'h3efffd9b76c8effeced528abe7b998fe343a199721f3417a33c4a6fb569cc75cca0775db6549ccfeb806a1204a587f377bdd5bc462f01c23674102f2e15006ded0450ddbe01124d8903b226a01dcbb5b546013b5ff04da6db2567300a9a14e52b59cce584a4b39fe62724d1dc5f76a9c344700c86a4e149b9c26623d2b4a10d6;
    5'b10010 : xpb = 1024'h95d90f093362f8d5b302637593a3b47ec70ba4206a48eb3217b08f8cce10ac0baa48213f42d8ba41c28db9529b9907127605bf3c3cd9e93a0bbcf3c4194e5c4e7caa9fefb85661f6bf9625adb35122b3f95902cc41171a9a2152641c56829f6f30c7b5da83bd48f5989718a691860a5e7a9396e45a1bc933f3a865ac50226024;
    5'b10011 : xpb = 1024'h3c04db212e0ecce3cc2a26682f3388ade8672b78dd26f4727dbfbec89281e3b287404f2a564128f62db6923e097b7e230c13facdf410e604ff99a537167a3d0cb4c0fd54e10aa1cfdc57264ecbe9c5dbaa4cf849f6a32db5dac1c33d49394df97ceb0b330c665f5f47fbfd50654483f772064e1df99e209c04baee16ec184907;
    5'b10100 : xpb = 1024'h92ddec8eeaa8d5bab0576131db1da42e7b38b602257c9e2a61aba75a09f5c8616780fa8e33d01639383daa705abc05fe063c5e45cdfab31ba41596084e78927c61268f68b94fdeee0bb229927d5e2d344f45e76038b56de249bdb458f61a9f15f815f2b545d86e567e20c8d930d323b9b852e439e96bd5345c3cf18610f09855;
    5'b10101 : xpb = 1024'h3909b8a6e554a9c8c97f242476ad785d9c943d5a985aa76ac7bad695ce67000844792879473884eda366835bc89e7d0e9c4a99d78531afe697f2477b4ba4733a993ceccde2041ec728732a3395f6d05c0039dcddee4180fe032d1379e8d14da04439480dce8184c02d85ad8304919d52afc59b7388ee2c9c6d4f79f0ace68138;
    5'b10110 : xpb = 1024'h8fe2ca14a1eeb29fadac5eee229793de2f65c7e3e0b05122aba6bf2745dae4b724b9d3dd24c77230aded9b8e19df04e99672fd4f5f1b7cfd3c6e384c83a2c8aa45a27ee1ba495be557ce2d77476b37b4a532cbf43053c12a7229049595b29ebcbf642f9007f393b763aa790bd0203d14f612318f78bbe134c4d17d5fd1bed086;
    5'b10111 : xpb = 1024'h360e962c9c9a86adc6d421e0be27680d50c14f3c538e5a6311b5ee630a4c1c5e01b201c8382fe0e51916747987c17bfa2c8138e1165279c8304ae9bf80cea9687db8dc46e2fd9bbe748f2e186003dadc5626c171e5dfd4462b9863b688694d470b8784e8909caa21130f5db5a3deb6aded84e8c9183e389cd5e405ca6db4b969;
    5'b11000 : xpb = 1024'h8ce7a79a59348f84ab015caa6a11838de392d9c59be4041af5a1d6f481c0010ce1f2ad2c15bece28239d8cabd90203d526a99c58f03c46ded4c6da90b8ccfed82a1e6e5abb42d8dca3ea315c11784234fb1fb08827f214729a9454d2354a9e6386b26c6aca0eb9184934293e6f6d567033d17ee5080bed352d660939928d08b7;
    5'b11001 : xpb = 1024'h331373b253e06392c4291f9d05a157bd04ee611e0ec20d5b5bb10630463138b3beeadb1729273cdc8ec6659746e47ae5bcb7d7eaa77343a9c8a38c03b5f8df966234cbbfe3f718b5c0ab31fd2a10e55cac13a605dd7e278e5403b3f328014cedd2d5c1c352b7cf81f8990de8432bd0092b44361ea78e449d3e7891a42e82f19a;
    5'b11010 : xpb = 1024'h89ec8520107a6c69a8565a66b18b733d97bfeba75717b7133f9ceec1bda51d629f2b867b06b62a1f994d7dc9982502c0b6e03b62815d10c06d1f7cd4edf735060e9a5dd3bc3c55d3f0063540db854cb5510c951c1f9067bac2ffa50ed4e29e0a4e00a9458c29de792ebdd9710eba6fcb7190cc3a975bf93595fa9513535b40e8;
    5'b11011 : xpb = 1024'h301851380b264077c17e1d594d1b476cb91b72ffc9f5c053a5ac1dfd821655097c23b4661a1e98d4047656b5060779d14cee76f438940d8b60fc2e47eb2315c446b0bb38e4f095ad0cc735e1f41defdd02008a99d51c7ad67c6f042fc7994c949a23fe9e14d2f4e2de22be1ae278e9646903837436de509da70d1d7def5129cb;
    5'b11100 : xpb = 1024'h86f162a5c7c0494ea5ab5822f90562ed4becfd89124b6a0b8998068ef98a39b85c645fc9f7ad86170efd6ee7574801ac4716da6c127ddaa205781f1923216b33f3164d4cbd35d2cb3c223925a5925735a6f979b0172ebb02eb6af54b747a9db1154ee6204e4503da144789a3ae078926af50199026ac0535fe8f20ed14297919;
    5'b11101 : xpb = 1024'h2d1d2ebdc26c1d5cbed31b159495371c6d4884e18529734befa735cabdfb715f395c8db50b15f4cb7a2647d2c52a78bcdd2515fdc9b4d76cf954d08c204d4bf22b2caab1e5ea12a458e339c6be2afa5d57ed6f2dccbace1ea4da546c67314c3b61723b78d6ee1a43c3ac6e4d81c602bfa6c2d0c9c62e5c9e0fa1a957b01f61fc;
    5'b11110 : xpb = 1024'h83f6402b7f062633a30055df407f529d001a0f6acd7f1d03d3931e5c356f560e199d3918e8a4e20e84ad6005166b0097d74d7975a39ea4839dd0c15d584ba161d7923cc5be2f4fc2883e3d0a6f9f61b5fce65e440ecd0e4b13d6458814129d57dc9d22fb1060293af9d139d64d54a281ed0f66e5b5fc11366723acc6d4f7b14a;
    5'b11111 : xpb = 1024'h2a220c4379b1fa41bc2818d1dc0f26cc217596c3405d264439a24d97f9e08db4f6956703fc0d50c2efd638f0844d77a86d5bb5075ad5a14e91ad72d0557782200fa89a2ae6e38f9ba4ff3dab883804ddadda53c1c4592166cd45a4a906c94be228c0785399093fa4a9361e8021131c1ae4821e1f557e689e7836353170ed9a2d;
    endcase
end

endmodule

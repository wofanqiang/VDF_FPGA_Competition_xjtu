module xpb_7_0
(
    input [7:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    7'b0000000 : xpb = 1024'h0;
    7'b0000001 : xpb = 1024'h4f52baaa3e11cb3734fa8828efa5b8ae8e89fccf2a885f88822346aa4cfd52f7fcb7828735d9817160a1c0b91ca1ef359be5d819dd4d2fb44f60c0a1c52d8b4e8bb0cb51506f02baed65fd5d67243bcf0bfb06677379d2ef4a736e0545d55d6dd0f86dd64f37077279401921082fd9d6b126211dafb4a2cfb99084fb771d9995;
    7'b0000010 : xpb = 1024'h9ea575547c23966e69f51051df4b715d1d13f99e5510bf1104468d5499faa5eff96f050e6bb302e2c14381723943de6b37cbb033ba9a5f689ec181438a5b169d176196a2a0de0575dacbfabace48779e17f60ccee6f3a5de94e6dc0a8baabadba1f0dbac9e6e0ee4f2803242105fb3ad624c423b5f69459f732109f6ee3b332a;
    7'b0000011 : xpb = 1024'h3d4aeaa8f8472cdcd3ea20a3be96e2ba3a27f33caa217e22088d1aa933f54bdff2de0a1cd76605c5828702e47287bcd66f9760677534bed13d83028714b62d3a2ec32d4541bc0aebb597f5759c90ef3c2fec199dcde74bbd29cdb815175575b743e1b7593cdc1dc9e500648420bf675ac4988476bed28b3ee64213eddc766654;
    7'b0000100 : xpb = 1024'h8c9da5533658f81408e4a8ccae3c9b68c8b1f00bd4a9ddaa8ab0615380f29ed7ef958ca40d3f8736e328c39d8f29ac0c0b7d38815281ee858ce3c328d9e3b888ba73f896922b0da6a2fdf2d303b52b0b3be7200541611eac7441261a5d2ad32514da252f8c13253c5e407da528ef413175bea5946e872e0e9fd298e95393ffe9;
    7'b0000101 : xpb = 1024'h2b431aa7b27c8e8272d9b91e8d880cc5e5c5e9aa29ba9cbb8ef6eea81aed44c7e90491b278f28a19a46c450fc86d8a774348e8b50d1c4dee2ba5446c643ecf25d1d58f393309131c7dc9ed8dd1fda2a953dd2cd42854c48b09280224e8d58e00b6cb00dc2a81342150c0afe7394ef4ded80ae7cfcdf073ae12f3a2e041cf3313;
    7'b0000110 : xpb = 1024'h7a95d551f08e59b9a7d441477d2dc574744fe6795442fc44111a355267ea97bfe5bc1439aecc0b8b050e05c8e50f79acdf2ec0ceea697da27b06050e296c5a745d865a8a837815d76b2feaeb3921de785fd8333b9bce977a539b702a2eaaeb6e87c36eb279b83b93ca00c908417eceb5893108ed7da5167dcc8427dbb8eccca8;
    7'b0000111 : xpb = 1024'h193b4aa66cb1f02811c951995c7936d19163e017a953bb551560c2a701e53dafdf2b19481a7f0e6dc651873b1e53581816fa7102a503dd0b19c78651b3c7711174e7f12d24561b4d45fbe5a6076a561677ce400a82c23d58e8824c34ba55a64a29b44a5f18264a78bc80fb4a51de8262eb7d4b28dd0e5c1d3fa531d2a727ffd2;
    7'b0001000 : xpb = 1024'h688e0550aac3bb5f46c3d9c24c1eef801feddce6d3dc1add978409514ee290a7dbe29bcf50588fdf26f347f43af5474db2e0491c82510cbf692846f378f4fc600098bc7e74c51e083361e3036e8e91e583c94671f63c104832f5ba3a002b03b7faacb835675d51eb35c1146b5a0e5c399ca36c468cc2feecf935b6ce1e459967;
    7'b0001001 : xpb = 1024'h7337aa526e751cdb0b8ea142b6a60dd3d01d68528ecd9ee9bca96a5e8dd3697d551a0ddbc0b92c1e836c966743925b8eaabf9503ceb6c2807e9c837035012fd17fa532115a3237e0e2dddbe3cd709839bbf5340dd2fb626c7dc96448bd5be939c9d93e205cb60d0284146ad6a6e0fe6feefae81ec2c448c6c56c0c50c80cc91;
    7'b0001010 : xpb = 1024'h5686354f64f91d04e5b3723d1b10198bcb8bd354537539771deddd5035da898fd2092364f1e5143348d88a1f90db14ee8691d16a1a389bdc574a88d8c87d9e4ba3ab1e7266122638fb93db1ba3fb4552a7ba59a850a9891612500449d1ab1c016d9601b855026842a1815fce729de9bdb015cf9f9be0e75c25e745c0839e6626;
    7'b0001011 : xpb = 1024'ha5d8eff9a30ae83c1aadfa660ab5d23a5a15d0237dfd98ffa01123fa82d7dc87cec0a5ec27be95a4a97a4ad8ad7d04242277a983f785cb90a6ab497a8dab299a2f5be9c3b68128f3e8f9d8790b1f8121b3b5600fc4235c055cc3724f1780796f3e8e6f8ea4396fb51ac178ef7acdc394613bf0bd4b958a2bdf77cabbfabbffbb;
    7'b0001100 : xpb = 1024'h447e654e1f2e7eaa84a30ab7ea0143977729c9c1d30e5810a457b14f1cd28277c82faafa937198876abdcc4ae6c0e28f5a4359b7b2202af9456ccabe1806403746bd8066575f2e69c3c5d333d967f8bfcbab6cdeab1701e3f1aa4e59a32b344ae07f4b3b42a77e9a0d41ab318b2d7741c38832f8aafecfcb5298d4b2e8f732e5;
    7'b0001101 : xpb = 1024'h93d11ff85d4049e1b99d92e0d9a6fc4605b3c690fd96b799267af7f969cfd56fc4e72d81c94b19f8cb5f8d040362d1c4f62931d18f6d5aad94cd8b5fdd33cb85d26e4bb7a7ce3124b12bd091408c348ed7a673461e90d4d33c1dbc5ee90091b8b177b91191de860c8681c452935d511874ae54165ab3729b0c2959ae6014cc7a;
    7'b0001110 : xpb = 1024'h3276954cd963e0502392a332b8f26da322c7c02f52a776aa2ac1854e03ca7b5fbe56329034fe1cdb8ca30e763ca6b0302df4e2054a07ba16338f0ca3678ee222e9cfe25a48ac369a8bf7cb4c0ed4ac2cef9c801505847ab1d104986974ab4c94536894be304c94f17901f694a3bd04c5d6fa9651ba1cb83a7f4a63a54e4fffa4;
    7'b0001111 : xpb = 1024'h81c94ff71775ab87588d2b5ba8982651b151bcfe7d2fd632ace4cbf850c7ce57bb0db5176ad79e4ced44cf2f59489f65c9daba1f2754e9ca82efcd452cbc6d717580adab991b3955795dc8a975f8e7fbfb97867c78fe4da11b78066eba80aa02246102947f839c63f2420fb5abecde9c8820b76f69d15b0a38dae8a0c56d9939;
    7'b0010000 : xpb = 1024'h206ec54b939941f5c2823bad87e397aece65b69cd2409543b12b594ceac27447b47cba25d68aa12fae8850a1928c7dd101a66a52e1ef493321b14e88b717840e8ce2444e39f93ecb5429c36444415f9a138d934b5ff1f37fb05ee279462b64ddc651de411df1ab48e4c241f7bc4c9249ea6cf9aac93aa0a9abfbf297b3a8cc63;
    7'b0010001 : xpb = 1024'h6fc17ff5d1ab0d2cf77cc3d67789505d5cefb36bfcc8f4cc334e9ff737bfc73fb1343cad0c6422a10f2a115aaf2e6d069d8c426cbf3c78e771120f2a7c450f5d18930f9f8a684186418fc0c1ab659b691f8899b2d36bc66efad2507e8c00c24b974a4c176d28b2bb5e025b18c47c6c209b931ac878ef4379658c77932ac665f8;
    7'b0010010 : xpb = 1024'he66f54a4dcea39b6171d42856d4c1ba7a03ad0a51d9b3dd37952d4bd1ba6d2faaa341bb78172583d06d92cce8724b71d557f2a079d6d8500fd3906e06a025fa2ff4a6422b4646fc1c5bbb7c79ae1307377ea681ba5f6c4d8fb92c8917ab7d27393b27c40b96c1a050828d5ad4dc1fcdfddf5d03d8588918d8ad818a19019922;
    7'b0010011 : xpb = 1024'h5db9aff48be06ed2966c5c51467a7a69088da9d97c621365b9b873f61eb7c027a75ac442adf0a6f5310f538605143aa7713dcaba572408045f34510fcbcdb148bba571937bb549b709c1b8d9e0d24ed64379ace92dd93f3cda2c9a8e5d80da950a33959a5acdc912c9c2a67bdd0bf9a4af057e21880d2be8923e0685901f32b7;
    7'b0010100 : xpb = 1024'had0c6a9ec9f23a09cb66e47a362033179717a6a8a6ea72ee3bdbbaa06bb5131fa41246c9e3ca286691b1143f21b629dd0d23a2d4347137b8ae9511b190fb3c9747563ce4cc244c71f727b63747f68aa54f74b350a153122c24a00893a3563802db2c0370aa04d0854302bf9ce53bd37b602b9f3f37c1ceb84bce8b81073ccc4c;
    7'b0010101 : xpb = 1024'h4bb1dff34615d078355bf4cc156ba474b42ba046fbfb31ff402247f505afb90f9d814bd84f7d2b4952f495b15afa084844ef5307ef0b97214d5692f51b5653345eb7d3876d0251e7d1f3b0f2163f0243676ac01f8846b80ab986e49e2f00f2de7d1cdf1d4872df6a3582f1def59b8728c277e17a972b1457beef9577f577ff76;
    7'b0010110 : xpb = 1024'h9b049a9d84279baf6a567cf505115d2342b59d1626839187c2458e9f52ad0c079a38ce5f8556acbab396566a779bf77de0d52b21cc58c6d59cb75396e083de82ea689ed8bd7154a2bf59ae4f7d633e127365c686fbc08afa03fa52a374d6504c4e154cf397a9e6dcaec30afffdcb60ff739e029846dfb72778801a736c95990b;
    7'b0010111 : xpb = 1024'h39aa0ff2004b321dd44b8d46e45cce805fc996b47b945098c68c1bf3eca7b1f793a7d36df109af9d74d9d7dcb0dfd5e918a0db5586f3263e3b78d4da6adef52001ca357b5e4f5a189a25a90a4babb5b08b5bd355e2b430d898e12eae00810b27f00628a03617f5c1a1433d420e2b14acd5ea44d3a648fcc6eba1246a5ad0cc35;
    7'b0011000 : xpb = 1024'h88fcca9c3e5cfd550946156fd402872eee539383a61cb02148af629e39a504ef905f55f526e3310ed57b9895cd81c51eb486b36f644055f28ad9957c300c806e8d7b00ccaebe5cd3878ba667b2cff17f9756d9bd562e03c7e3549cb346566895c0fe9676854efd341a835663165aee83871065f155fd9f96a531a965d1ee65ca;
    7'b0011001 : xpb = 1024'h27a23ff0ba8093c3733b25c1b34df88c0b678d21fb2d6f324cf5eff2d39faadf89ce5b03929633f196bf1a0806c5a389ec5263a31edab55b299b16bfba67970ba4dc976f4f9c62496257a1228118691daf4ce68c3d21a9a6783b78bdd201237162ef722323bd0c190d0388a526baa230e95ca82cb566e5361852b35cc02998f4;
    7'b0011010 : xpb = 1024'h76f4fa9af8925efaa835adeaa2f3b13a99f189f125b5cebacf19369d209cfdd78685dd8ac86fb562f760dac1236792bf88383bbcfc27e50f78fbd7617f95225a308d62c0a00b65044fbd9e7fe83ca4ecbb47ecf3b09b7c95c2aee6c317d680df33e7dff972f4138b8643a1c62eea7c079a82c94a651b8805d1e3385837473289;
    7'b0011011 : xpb = 1024'h159a6fef74b5f569122abe3c823f2297b705838f7ac68dcbd35fc3f1ba97a3c77ff4e2993422b845b8a45c335cab712ac003ebf0b6c2447817bd58a509f038f747eef96340e96a7a2a89993ab6851c8ad33df9c2978f22745795c2cda3813bbad5d8bba61162227078c3d4083f4a2fb4fccf0b85c484cda54504424f258265b3;
    7'b0011100 : xpb = 1024'h64ed2a99b2c7c0a04725466571e4db46458f805ea54eed5455830a9c0794f6bf7cac652069fc39b719461cec794d60605be9c40a940f742c671e1946cf1dc445d39fc4b491586d3517ef96981da95859df39002a0b08f563a20930d2e9569928a6d1297c609929e2f203ed29477a098badf52ca374397074fe94c74a9c9fff48;
    7'b0011101 : xpb = 1024'h3929fee2eeb570eb11a56b751304ca362a379fcfa5fac6559c997f0a18f9caf761b6a2ed5af3c99da899e5eb2913ecb93b5743e4ea9d39505df9a8a5978dae2eb015b57323672aaf2bb9152ebf1cff7f72f0cf8f1fc9b4236f00cdd7501540448c20528ff0738c7e4841f6b57d9bd3910416eded3a2b61471b5d1418adb3272;
    7'b0011110 : xpb = 1024'h52e55a986cfd2245e614dee040d60551f12d76cc24e80beddbecde9aee8cefa772d2ecb60b88be0b3b2b5f17cf332e012f9b4c582bf7034955405b2c1ea6663176b226a882a57565e0218eb053160bc7032a136065766e3181637ae2bad6b17219ba72ff4e3e403a5dc4388c6009970fc1678ffc835758e42b46563d01f8cc07;
    7'b0011111 : xpb = 1024'ha2381542ab0eed7d1b0f6709307bbe007fb7739b4f706b765e1025453b8a429f6f8a6f3d41623f7c9bcd1fd0ebd51d36cb812472094432fda4a11bcde3d3f1800262f1f9d3147820cd878c0dba3a47960f2519c7d8f04120cbd6e8e800ac0edfeab2e0d59d7547acd70451ad683970e6728db11a330bfbb3e4d6db387916659c;
    7'b0100000 : xpb = 1024'h40dd8a97273283eb8504775b0fc72f5d9ccb6d39a4812a876256b299d584e88f68f9744bad15425f5d10a1432518fba2034cd4a5c3de926643629d116e2f081d19c4889c73f27d96a85386c88882bf34271b2696bfe3e6ff60bdc4f28c56c9bb8ca3bc823be35691c98483ef78992493d4d9f3559275415357f7e52f675198c6;
    7'b0100001 : xpb = 1024'h9030454165444f22b9feff83ff6ce80c2b556a08cf098a0fe479f94422823b8765b0f6d2e2eec3d0bdb261fc41baead79f32acbfa12bc21a92c35db3335c936ba57553edc461805195b98425efa6fb0333162cfe335db9eeab3132f7d22c27295d9c2a588b1a5e0442c49d1080c8fe6a860014734229e42311886a2ade6f325b;
    7'b0100010 : xpb = 1024'h2ed5ba95e167e59123f40fd5deb85969486963a7241a4920e8c08698bc7ce1775f1ffbe14ea1c6b37ef5e36e7afec942d6fe5cf35bc621833184def6bdb7aa08bcd6ea90653f85c770857ee0bdef72a14b0c39cd1a515fcd40180f025dd6e204ff8d060529886ce93544cf529128b217e84c56aea19329c284a97421ccaa6585;
    7'b0100011 : xpb = 1024'h7e2875401f79b0c858ee97fece5e1217d6f360764ea2a8a96ae3cd43097a346f5bd77e68847b4824df97a42797a0b87872e4350d3913513780e59f9882e535574887b5e1b5ae88825deb7c3e2513ae70570740348dcb32bc8a8b7d07a3ac3f72d08573db78bf745bae84e87399588bee997277cc5147cc923e39f91d43c7ff1a;
    7'b0100100 : xpb = 1024'h1ccdea949b9d4736c2e3a850ada98374f4075a14a3b367ba6f2a5a97a374da5f55468376f02e4b07a0db2599d0e496e3aaafe540f3adb0a01fa720dc0d404bf45fe94c84568c8df838b776f8f35c260e6efd4d0374bed89b1f7259122f56fa4e72764f88172d8340a1051ab5a9b83f9bfbbeba07b0b11231b15b031432033244;
    7'b0100101 : xpb = 1024'h6c20a53ed9af126df7de30799d4f3c23829156e3ce3bc742f14da141f0722d5751fe05fe2607cc79017ce652ed8686194695bd5ad0fae0546f07e17dd26dd742eb9a17d5a6fb90b3261d74565a8061dd7af8536ae838ab8a69e5c717752c57bc436ebd5e66648ab31a4533d6b1e81972ace4db256065b5016aeb880fa920cbd9;
    7'b0100110 : xpb = 1024'hac61a9355d2a8dc61d340cb7c9aad809fa55082234c8653f5942e968a6cd3474b6d0b0c91bacf5bc2c067c526ca64847e616d8e8b953fbd0dc962c15cc8ede002fbae7847d9962900e96f1128c8d97b92ee6039cf2c5168fecca32200d71297e55f990b04d299980cc56618c247cd200f311d60bfcefaa0de0c9206975bff03;
    7'b0100111 : xpb = 1024'h5a18d53d93e4741396cdc8f46c40662f2e2f4d514dd4e5dc77b77540d76a263f48248d93c79450cd2362287e436c53ba1a4745a868e26f715d2a236321f6792e8eac79c9984898e3ee4f6c6e8fed154a9ee966a142a624584940112746ac7005b65806e15409a10a86057f39ca77a6f6c0573e7e6f839d70979d17020e799898;
    7'b0101000 : xpb = 1024'ha96b8fe7d1f63f4acbc8511d5be61eddbcb94a20785d4564f9dabbeb2467793744dc101afd6dd23e8403e937600e42efb62d1dc2462f9f25ac8ae404e724047d1a5d451ae8b79b9edbb569cbf7115119aae46d08b61ff74793b37f2c8c81cd73875074b7a340a87cff45985ad2a780cd717d5f9c1f384040512d9bfd8597322d;
    7'b0101001 : xpb = 1024'h4811053c4e19d5b935bd616f3b31903ad9cd43becd6e0475fe21493fbe621f273e4b15296920d52145476aa99952215aedf8cdf600c9fe8e4b4c6548717f1b1a31bedbbd8995a114b6816486c559c8b7c2da79d79d139d26289a5b37182c884f2941506441aeb761f1c5ca9ce307347ad3c9a1d77ea185dfc44ea5f473d26557;
    7'b0101010 : xpb = 1024'h9763bfe68c2ba0f06ab7e9982ad748e96857408df7f663fe80448fea0b5f721f3b0297b09efa5692a5e92b62b5f4109089dea60fde172e429aad25ea36aca668bd6fa70eda04a3cfa3e761e42c7e0486ced5803f108d7015730dc93c5e01e5bcfa39be3a90e5bed46b05e3bdeb370e5184efc2f52e5628af7ddf2aefeaeffeec;
    7'b0101011 : xpb = 1024'h3609353b084f375ed4acf9ea0a22ba46856b3a2c4d07230f848b1d3ea55a180f34719cbf0aad5975672cacd4ef37eefbc1aa564398b18dab396ea72dc107bd05d4d13db17ae2a9457eb35c9efac67c24e6cb8d0df78115f407f4a546e9aca0989c2a99e72f53cdb95d8615fffb96c1fee73c05308dbf6e4ef10034e6d92b3216;
    7'b0101100 : xpb = 1024'h855befe54661029609a78212f9c872f513f536fb778f829806ae63e8f2576b0731291f464086dae6c7ce6d8e0bd9de315d902e5d75febd5f88cf67cf8635485460820902cb51ac006c1959fc61eab7f3f2c693756afae8e35268134c2f81fe066d2307bd7e8ad52bd6c62f2103c69bd59862264e3d74111eaa90b9e25048cbab;
    7'b0101101 : xpb = 1024'h24016539c2849904739c9264d913e45231093099cca041a90af4f13d8c5210f72a982454ac39ddc98911ef00451dbc9c955bde9130991cc82790e91310905ef177e39fa56c2fb17646e554b730332f920abca04451ee8ec1e74eef56bb2cb8e20f13e36a1cf8e410c946616314264f82faae68899cdd56be1db1c3d93e83fed5;
    7'b0101110 : xpb = 1024'h73541fe40096643ba8971a8dc8b99d00bf932d68f728a1318d1837e7d94f63ef274fa6dbe2135f3ae9b3afb961bfabd23141b6ab0de64c7c76f1a9b4d5bdea4003946af6bc9eb431344b521497576b6116b7a6abc56861b131c25d5c0102164fe00c51406c2feb8342867a841c562959abd489a74c91f98dd74248d4b5a1986a;
    7'b0101111 : xpb = 1024'h11f995387cb9faaa128c2adfa8050e5ddca727074c396042915ec53c734a09df20beabea4dc6621daaf7312b9b038a3d690d66dec880abe515b32af8601900dd1af601995d7cb9a70f174ccf659fe2ff2eadb37aac5c078fc6a939668cacd12b81fd2ced0a9dfa683506acc62cb5dd070e20cbe2abfb3f2d4a6352cba3dccb94;
    7'b0110000 : xpb = 1024'h614c4fe2bacbc5e14786b30897aac70c6b3123d676c1bfcb13820be6c0475cd71d762e71839fe38f0b98f1e4b7a5797304f33ef8a5cddb996513eb9a25468c2ba6a6cceaadebbc61fc7d4a2cccc41ece3aa8b9e21fd5da7f111ca76bd2822e9952f59ac359d501daae46c5e734e5b6ddbf46ed005bafe1fd03f3d7c71afa6529;
    7'b0110001 : xpb = 1024'hb09f0a8cf8dd91187c813b3187507fbaf9bb20a5a14a1f5395a552910d44afcf1a2db0f8b97965006c3ab29dd44768a8a0d91712831b0b4db474ac3bea74177a3257983bfe5abf1ce9e3478a33e85a9d46a3c049934fad6e5b90157118578c0723ee0899a90c094d2786df083d1590b4706d0e1e0b6484ccbd845cc29217febe;
    7'b0110010 : xpb = 1024'h4f447fe175012786e6764b83669bf11816cf1a43f65ade6499ebdfe5a73f55bf139cb607252c67e32d7e34100d8b4713d8a4c7463db56ab653362d7f74cf2e1749b92ede9f38c492c4af42450230d23b5e99cd187a43534cf076f17ba40246e2c5dee446477a18321a07114a4d754461d2b950596acdca6c30a566b9805331e8;
    7'b0110011 : xpb = 1024'h9e973a8bb312f2be1b70d3ac5641a9c6a559171320e33ded1c0f268ff43ca8b71054388e5b05e9548e1ff4c92a2d3649748a9f601b029a6aa296ee2139fcb965d569fa2fefa7c74db2153fa269550e0a6a94d37fedbd263c3aea5f80e9d7a45096d7521c96b11fa493472a6b55a51e3883df71771a826d3bea35ebb4f770cb7d;
    7'b0110100 : xpb = 1024'h3d3cafe02f36892c8565e3fe358d1b23c26d10b175f3fcfe2055b3e48e374ea709c33d9cc6b8ec374f63763b637114b4ac564f93d59cf9d341586f64c457d002eccb90d29085ccc38ce13a5d379d85a8828ae04ed4b0cc1acfd13b8b75825f2c38c82dc9351f2e8985c75cad6604d1e5e62bb3b279ebb2db5d56f5abe5abfea7;
    7'b0110101 : xpb = 1024'h8c8f6a8a6d485463ba606c272532d3d250f70d80a07c5c86a278fa8edb34a19f067ac023fc926da8b00536f4801303ea483c27adb2ea298790b9300689855b51787c5c23e0f4cf7e7a4737ba9ec1c1778e85e6b6482a9f0a1a44a990bb57bc9a09c09b9f845635fbff0775ce6e34abbc9751d4d029a055ab16e77aa75cc9983c;
    7'b0110110 : xpb = 1024'h2b34dfdee96bead224557c79047e452f6e0b071ef58d1b97a6bf87e3752f478effe9c5326845708b7148b866b956e2558007d7e16d8488f02f7ab14a13e071ee8fddf2c681d2d4f4551332756d0a3915a67bf3852f1e44e8af2b859b47027775abb1774c22c444e0f187a8107e945f69f99e170b89099b4a8a08849e4b04cb66;
    7'b0110111 : xpb = 1024'h7a879a89277db609595004a1f423fdddfc9503ee20157b2028e2ce8dc22c9a86fca147b99e1ef1fcd1ea791fd5f8d18b1bedaffb4ad1b8a47edb71ebd90dfd3d1b8ebe17d241d7af42792fd2d42e74e4b276f9eca29817d7f99ef3a08cd7d4e37ca9e52271fb4c536ac7c13186c43940aac4382938be3e1a43990999c22264fb;
    7'b0111000 : xpb = 1024'h192d0fdda3a14c77c34514f3d36f6f3b19a8fd8c75263a312d295be25c274076f6104cc809d1f4df932dfa920f3caff653b9602f056c180d1d9cf32f636913da32f054ba731fdd251d452a8da276ec82ca6d06bb898bbdb68e85cfab18828fbf1e9ac0cf10695b385d47f3739723ecee0d107a64982783b9b6ba1390b05d9825;
    7'b0111001 : xpb = 1024'h687fca87e1b317aef83f9d1cc31527e9a832fa5b9fae99b9af4ca28ca924936ef2c7cf4f3fab7650f3cfbb4b2bde9f2bef9f3848e2b947c16cfdb3d128969f28bea1200bc38edfe00aab27eb099b2851d6680d22fd0590a5d8f93db05e57ed2cef932ea55fa062aad6880c949f53c6c4be369b8247dc2689704a988c277b31ba;
    7'b0111010 : xpb = 1024'h7253fdc5dd6ae1d6234ad6ea2609946c546f3f9f4bf58cab3932fe1431f395eec36d45dab5e7933b5133cbd65227d97276ae87c9d53a72a0bbf3514b2f1b5c5d602b6ae646ce555e57722a5d7e39fefee5e19f1e3f936846de019baea02a80891840a51fe0e718fc9083ed6afb37a722082ddbda7456c28e36ba28315b664e4;
    7'b0111011 : xpb = 1024'h5677fa869be87954972f3597920651f553d0f0c91f47b85335b6768b901c8c56e8ee56e4e137faa515b4fd7681c46cccc350c0967aa0d6de5b1ff5b6781f411461b381ffb4dbe810d2dd20033f07dbbefa59205957730973b85387c02fd80576627c78284d457902424857f7b7e35448d1a8fedb56fa0ef89cfc277e8cd3fe79;
    7'b0111100 : xpb = 1024'ha5cab530d9fa448bcc29bdc081ac0aa3e25aed9849d017dbb7d9bd35dd19df4ee5a5d96c17117c167656be2f9e665c025f3698b057ee0692aa80b6583d4ccc62ed644d51054aeacbc0431d60a62c178e065426c0caecdc6302c6f5c575ad62e43374e5fe9c7c8074bb887118c0132e1f82cf1ff906aeb1c8568cac7a03f1980e;
    7'b0111101 : xpb = 1024'h44702a85561ddafa361ece1260f77c00ff6ee7369ee0d6ecbc204a8a7714853edf14de7a82c47ef9379a3fa1d7aa3a6d970248e4128865fb4942379bc7a7e30004c5e3f3a628f0419b0f181b74748f2c1e4a338fb1e0824197add1d001581dbfd565c1ab3aea8f59ae08a35ad072e1cce51b62346617f767c9adb670f22ccb38;
    7'b0111110 : xpb = 1024'h93c2e52f942fa6316b19563b509d34af8df8e405c96936753e439134c411d836dbcc6101b89e006a983c005af44c29a332e820fdefd595af98a2f83d8cd56e4e9076af44f697f2fc88751578db98cafb2a4539f7255a5530e2213fd5472d7b2da65e2f818a2196cc2748bc7bd8a2bba39641835215cc9a37833e3b6c694a64cd;
    7'b0111111 : xpb = 1024'h32685a8410533c9fd50e668d2fe8a60cab0cdda41e79f586428a1e895e0c7e26d53b66102451034d597f81cd2d90080e6ab3d131aa6ff51837647981173084eba7d845e79775f87263411033a9e14299423b46c60c4dfb0f77081bdfd2d83609484f0b2e288fa5b119c8eebde9026f50f88dc58d7535dfd6f65f4563578597f7;
    7'b1000000 : xpb = 1024'h81bb152e4e6507d70a08eeb61f8e5ebb3996da734902550ec4ad6533ab09d11ed1f2e8975a2a84beba2142864a31f7440699a94b87bd24cc86c53a22dc5e103a33891138e7e4fb2d50a70d9111057e684e364d2d7fc7cdfec17b89e518ad93771947790477c6ad23930907def1324927a9b3e6ab24ea82a6afefca5ecea3318c;
    7'b1000001 : xpb = 1024'h20608a82ca889e4573fdff07fed9d01856aad4119e13141fc8f3f2884504770ecb61eda5c5dd87a17b64c3f88375d5af3e65597f425784352586bb6666b926d74aeaa7db88c300a32b73084bdf4df606662c59fc66bb73dd566265efa4584e52bb3854b11634bc0885893a210191fcd50c0028e68453c8462310d455bcde64b6;
    7'b1000010 : xpb = 1024'h6fb3452d089a697ca8f88730ee7f88c6e534d0e0c89b73a84b1739329201ca06c819702cfbb70912dc0684b1a017c4e4da4b31991fa4b3e974e77c082be6b225d69b732cd932035e18d905a9467231d572276063da3546cca0d5d3f4ea2dabc08c30c287656bc37afec9534209c1d6abbd264a0434086b15dca1595133fbfe4b;
    7'b1000011 : xpb = 1024'he58ba8184bdffeb12ed9782cdcafa240248ca7f1dac32b94f5dc6872bfc6ff6c188753b676a0bf59d4a0623d95ba3501216e1ccda3f135213a8fd4bb641c8c2edfd09cf7a1008d3f3a5006414baa9738a1d6d32c128ecab35bcafff75d8669c2e219e3403d9d25ff14985841a218a591f728c3f9371b0b54fc2634822373175;
    7'b1000100 : xpb = 1024'h5dab752bc2cfcb2247e81fabbd70b2d290d2c74e48349241d1810d3178f9c2eebe3ff7c29d438d66fdebc6dcf5fd9285adfcb9e6b78c43066309bded7b6f541179add520ca7f0b8ee10afdc17bdee5429618739a34a2bf9a80301e04bbadc409ff1a0c0a5310d9d26a899ea52251642fd098ad5d432653850952e8439954cb0a;
    7'b1000101 : xpb = 1024'hacfe2fd600e196597ce2a7d4ad166b811f5cc41d72bcf1ca53a453dbc5f715e6baf77a49d31d0ed85e8d8796129f81bb49e2920094d972bab26a7e8f409cdf60055ea0721aee0e49ce70fb1ee3032111a2137a01a81c9289caa38c0a01832177d01279e0a247e144e3c9b7c62a813e0681bece7af2daf654c2e36d3f1072649f;
    7'b1000110 : xpb = 1024'h4ba3a52a7d052cc7e6d7b8268c61dcde3c70bdbbc7cdb0db57eae1305ff1bbd6b4667f583ed011bb1fd109084be3602681ae42344f73d223512bffd2caf7f5fd1cc03714bbcc13bfa93cf5d9b14b98afba0986d08f1038685f8a68148d2ddc537203558d40b5f029d649ea083ae0f1b3e40b10b652443bf436047735fead97c9;
    7'b1000111 : xpb = 1024'h9af65fd4bb16f7ff1bd2404f7c07958ccafaba8af2561063da0e27daacef0eceb11e01df74a9932c8072c9c168854f5c1d941a4e2cc101d7a08cc0749025814ba87102660c3b167a96a2f337186fd47ec6048d38028a0b57a9fdd619d30339c142fbc3638fecf79c4f8a03294310cb8a953131d401f8dec3ef94fc3175cb315e;
    7'b1001000 : xpb = 1024'h399bd529373a8e6d85c750a15b5306e9e80eb4294766cf74de54b52f46e9b4beaa8d06ede05c960f41b64b33a1c92dc7555fca81e75b61403f4e41b81a8097e8bfd29908ad191bf0716eedf1e6b84c1cddfa9a06e97db1363ee4b2245eadf49ce4ec9f102e5b0681420a356b53707f37f77d740f6162246362b6062864066488;
    7'b1001001 : xpb = 1024'h88ee8fd3754c59a4bac1d8ca4af8bf987698b0f871ef2efd6077fbd993e707b6a744897516361780a2580becbe6b1cfcf145a29bc4a890f48eaf0259dfae23374b836459fd881eab5ed4eb4f4ddc87ebe9f5a06e5cf7842589582029a483520ab5e50ce67d920df3bb4a4e8c5ba0590ea8a3952d1116c7331c468b23db23fe1d;
    7'b1001010 : xpb = 1024'h27940527f16ff01324b6e91c2a4430f593acaa96c6ffee0e64be892e2de1ada6a0b38e8381e91a63639b8d5ef7aefb68291152cf7f42f05d2d70839d6a0939d462e4fafc9e66242139a0e60a1c24ff8a01ebad3d43eb2a041e3efc34302e0ce657d5e8931c001cd8adca80ce6c000cbc0aefd76870800cd28f67951ac95f3147;
    7'b1001011 : xpb = 1024'h76e6bfd22f81bb4a59b1714519e9e9a42236a765f1884d96e6e1cfd87adf009e9d6b110ab7c29bd4c43d4e181450ea9dc4f72ae95c9020117cd1443f2f36c522ee95c64deed526dc2706e36783493b590de6b3a4b764fcf368b26a3976036a5428ce56696b37244b270a99ef742fe692bc15f8862034afa248f81a16407ccadc;
    7'b1001100 : xpb = 1024'h158c3526aba551b8c3a68196f9355b013f4aa10446990ca7eb285d2d14d9a68e96da161923759eb78580cf8a4d94c908fcc2db1d172a7f7a1b92c582b991dbc005f75cf08fb32c5201d2de225191b2f725dcc0739e58a2d1fd99464401ae252fcabf321609a53330198acc31848f9a401e623ac17f9df541bc19240d2eb7fe06;
    7'b1001101 : xpb = 1024'h64deefd0e9b71ceff8a109bfe8db13afcdd49dd371216c306d4ba3d761d6f986939198a0594f2028e62290436a36b83e98a8b336f477af2e6af386247ebf670e91a82841e0222f0cef38db7fb8b5eec631d7c6db11d275c1480cb4494783829d9bb79fec58dc3aa292cae5528cbf7416cf885bdf2f52981175a9a908a5d5979b;
    7'b1001110 : xpb = 1024'h384652565dab35e62961a11c826850ceae89771c6322b417192312bfbd19f768d009daec502230ba76611b5a37a96a9d074636aaf120e9709b50768091a7daba909bee481003482ca04d63a86fe666449cdd3a9f8c61b9fdcf39053d32e3d793da87b98f74a4987854b17949d1f27c431d49e1a8ebbddb0e8cab2ff9410cac5;
    7'b1001111 : xpb = 1024'h52d71fcfa3ec7e959790a23ab7cc3dbb79729440f0ba8ac9f3b577d648cef26e89b82035fadba47d0807d26ec01c85df6c5a3b848c5f3e4b5915c809ce4808fa34ba8a35d16f373db76ad397ee22a23355c8da116c3fee8f2766fe5919039ae70ea0e96f468150f9fe8b30b5a54f019ae2fabf383e708080a25b37fb0b2e645a;
    7'b1010000 : xpb = 1024'ha229da79e1fe49cccc8b2a63a771f66a07fc91101b42ea5275d8be8095cc4566866fa2bd30b525ee68a99327dcbe75150840139e69ac6dffa87688ab93759448c06b558721de39f8a4d0d0f55546de0261c3e078dfb9c17e71da6c5e5ed8f854df99574595b8586c77cb49d6ad7edb719420e055ee2523505bebbcf6824bfdef;
    7'b1010001 : xpb = 1024'h40cf4fce5e21e03b36803ab586bd67c725108aae7053a9637a1f4bd52fc6eb567fdea7cb9c6828d129ed149a16025380400bc3d22446cd68473809ef1dd0aae5d7ccec29c2bc3f6e7f9ccbb0238f55a079b9ed47c6ad675d06c14868ea83b330818a32f2342667516a4b7c18bdde8f1ef66d22914d8e68efcf0cc6ed70873119;
    7'b1010010 : xpb = 1024'h90220a789c33ab726b7ac2de76632075b39a877d9adc08ebfc42927f7cc43e4e7c962a52d241aa428a8ed55332a442b5dbf19bec0193fd1c9698ca90e2fe3634637db77b132b42296d02c90d8ab3916f85b4f3af3a273a4c5134b66e3059109e5282a0c8835d6ec3e38b9539c60e68f5a79343aefd430bbf889d4be8e7a4caae;
    7'b1010011 : xpb = 1024'h2ec77fcd185741e0d56fd33055ae91d2d0ae811befecc7fd00891fd416bee43e76052f613df4ad254bd256c56be8212113bd4c1fbc2e5c85355a4bd46d594cd17adf4e1db409479f47cec3c858fc090d9dab007e211ae02ae61b9278bc03cb79f4737c7521cb7da8d60bc77bd66e1ca309df85ea5cac515efbbe55dfd5dffdd8;
    7'b1010100 : xpb = 1024'h7e1a3a7756690d180a6a5b5945544a815f387deb1a75278582ac667e63bc373672bcb1e873ce2e96ac74177e888a1056afa32439997b8c3984bb0c763286d8200690196f04784a5a3534c125c02044dca9a606e59494b31a308f007e01d928e7c56bea4b7102851b4f4be09cde9df679bb05a7080c60f42eb54edadb4cfd976d;
    7'b1010101 : xpb = 1024'h1cbfafcbd28ca386745f6bab249fbbde7c4c77896f85e69686f2f3d2fdb6dd266c2bb6f6df8131796db798f0c1cdeec1e76ed46d5415eba2237c8db9bce1eebd1df1b011a5564fd01000bbe08e68bc7ac19c13b47b8858f8c575dc888d83e3c3675cc5f80f70940041cc12deeefdaa271d51e9436bca39ce286fe4d23b38ca97;
    7'b1010110 : xpb = 1024'h6c126a76109e6ebda959f3d41445748d0ad674589a0e461f09163a7d4ab4301e68e3397e155ab2eace5959a9de6fddf78354ac8731631b5672dd4e5b820f7a0ba9a27b62f5c5528afd66b93df58cf849cd971a1bef022be80fe94a8dd3594131385533ce5ea79b72bb0c2bfff72d83fdce780a611b7edc9de20069cdb256642c;
    7'b1010111 : xpb = 1024'hab7dfca8cc2052c134f0425f390e5ea27ea6df6ef1f05300d5cc7d1e4aed60e62523e8c810db5cd8f9cdb1c17b3bc62bb205cbaebfd7abf119ecf9f0c6a90a8c104120596a35800d832b3f8c3d56fe7e58d26ead5f5d1c6a4d026985f03fc0cda460f7afd15aa57ad8c5e42078d37ab30c44c9c7ae8223d552173c4a0919756;
    7'b1011000 : xpb = 1024'h5a0a9a74cad3d06348498c4ee3369e98b6746ac619a764b88f800e7c31ac29065f09c113b6e7373ef03e9bd53455ab98570634d4c94aaa7360ff9040d1981bf74cb4dd56e7125abbc598b1562af9abb6f1882d52496fa4b5ef43949da4d9597aab3e7d514c4cb1ca26cc77630fbd1181e1ea6dba2a9cc50d0eb1f8c017af30eb;
    7'b1011001 : xpb = 1024'ha95d551f08e59b9a7d441477d2dc574744fe6795442fc44111a355267ea97bfe5bc1439aecc0b8b050e05c8e50f79acdf2ec0ceea697da27b06050e296c5a745d865a8a837815d76b2feaeb3921de785fd8333b9bce977a539b702a2eaaeb6e87c36eb279b83b93ca00c908417eceb5893108ed7da5167dcc8427dbb8eccca80;
    7'b1011010 : xpb = 1024'h4802ca7385093208e73924c9b227c8a4621261339940835215e9e27b18a421ee553048a95873bb931223de008a3b79392ab7bd22613239904f21d2262120bde2efc73f4ad85f62ec8dcaa96e60665f2415794088a3dd1d83ce9ddead765971c41e27c6d439f1c821928cc2c6284c9f05f55cd11339baad7c3b6387b27d07fdaa;
    7'b1011011 : xpb = 1024'h9755851dc31afd401c33acf2a1cd8152f09c5e02c3c8e2da980d292565a174e651e7cb308e4d3d0472c59eb9a6dd686ec69d953c3e7f69449e8292c7e64e49317b780a9c28ce65a77b30a6cbc78a9af3217446f01756f07319114cb2bc2ecf31ef2034aa8928cf940bccdbe7307c78dca682f230e96f504bf4f40cadf425973f;
    7'b1011100 : xpb = 1024'h35fafa723f3e93ae8628bd448118f2b00db057a118d9a1eb9c53b679ff9c1ad64b56d03efa003fe73409202be02146d9fe69456ff919c8ad3d44140b70a95fce92d9a13ec9ac6b1d55fca18695d31291396a53befe4a9651adf828bd47d98a0d911110572796de78fe4d0e2940dc2c8a08cf346c48d895eb681516a4e260ca69;
    7'b1011101 : xpb = 1024'h854db51c7d505ee5bb23456d70beab5e9c3a5470436201741e76fd244c996dce480e52c62fd9c15894aae0e4fcc3360f9a4f1d89d666f8618ca4d4ad35d6eb1d1e8a6c901a1b6dd843629ee3fcf74e6045655a2671c46940f86b96c28daee77b62097e2d76cde5eb778d274a490c0660b9f55589f88d38bb21a59ba0597e63fe;
    7'b1011110 : xpb = 1024'h23f32a70f973f554251855bf500a1cbbb94e4e0e9872c08522bd8a78e69413be417d57d49b8cc43b55ee62573607147ad21acdbd910157ca2b6655f0c03201ba35ec0332baf9734e1e2e999ecb3fc5fe5d5b66f558b80f1f8d5272cd1959a25703fa59da153bf4d06a0d598c596bba0e1c4197c557f67e5a94c6a59747b99728;
    7'b1011111 : xpb = 1024'h7345e51b3785c08b5a12dde83fafd56a47d84addc2fb200da4e0d123339166b63e34da5bd16645acb690231052a903b06e00a5d76e4e877e7ac71692855f8d08c19cce840b6876090b9496fc326401cd69566d5ccc31e20ed7c5e0d25f2effc4d4f2c7b06472fc42e34d72ad619b93e4cd67b8e307ab212a4e572a92bed730bd;
    7'b1100000 : xpb = 1024'h11eb5a6fb3a956f9c407ee3a1efb46c764ec447c180bdf1ea9275e77cd8c0ca637a3df6a3d19488f77d3a4828bece21ba5cc560b28e8e6e7198897d60fbaa3a5d8fe6526ac467b7ee66091b700ac796b814c7a2bb32587ed6cacbcdcead9baa076e3a35d02e10b27d5cda4ef71fb47922fb3fb1e671466c9c1783489ad1263e7;
    7'b1100001 : xpb = 1024'h613e1519f1bb2230f90276630ea0ff75f376414b42943ea72b4aa5221a895f9e345b61f172f2ca00d875653ba88ed15141b22e250636169b68e95877d4e82ef464af3077fcb57e39d3c68f1467d0b53a8d478093269f5adcb7202ae230af180e47dc11335218129a4f0dbe107a2b2168e0da1c3c16c909997b08b985242ffd7c;
    7'b1100010 : xpb = 1024'hb090cfc42fcced682dfcfe8bfe46b82482003e1a6d1c9e2fad6debcc6786b2963112e478a8cc4b72391725f4c530c086dd98063ee383464fb84a19199a15ba42f05ffbc94d2480f4c12c8c71cef4f109994286fa9a192dcc019398e77684757c18d47f09a14f1a0cc84dd731825afb3f92003d59c67dac6934993e809b4d9711;
    7'b1100011 : xpb = 1024'h4f364518abf083d697f20edddd9229819f1437b8c22d5d40b1b47921018158862a81e987147f4e54fa5aa766fe749ef21563b6729e1da5b8570b9a5d2470d0e007c1926bee02866a9bf8872c9d3d68a7b13893c9810cd3aa967a74f2022f3057bac55ab63fbd28f1bace097392baaeecf44c7f9525e6f208a7ba48778988ca3b;
    7'b1100100 : xpb = 1024'h9e88ffc2ea024f0dccec9706cd37e2302d9e3487ecb5bcc933d7bfcb4e7eab7e27396c0e4a58cfc65afc68201b168e27b1498e8c7b6ad56ca66c5afee99e5c2e93725dbd3e718925895e848a0461a476bd339a30f486a699e0ede2f748048dc58bbdc88c8ef43064340e22949aea88c3a572a0b2d59b94d8614acd7300a663d0;
    7'b1100101 : xpb = 1024'h3d2e75176625e57c36e1a758ac83538d4ab22e2641c67bda381e4d1fe879516e20a8711cb60bd2a91c3fe992545a6c92e9153ec0360534d5452ddc4273f972cbaad3f45fdf4f8e9b642a7f44d2aa1c14d529a6ffdb7a4c7875d4bf01d3af48a12daea4392d623f49268e54d6ab4a3c7107bee2ee3504da77d46bd769eee196fa;
    7'b1100110 : xpb = 1024'h8c812fc1a437b0b36bdc2f819c290c3bd93c2af56c4edb62ba4193ca3576a4661d5ff3a3ebe5541a7ce1aa4b70fc5bc884fb16da13526489948e9ce43926fe1a3684bfb12fbe915651907ca239ce57e3e124ad674ef41f67c0482d071984a60efea7120f7c9946bb9fce6df7b37a1647b8e5040be4b97d478dfc5c6565ff308f;
    7'b1100111 : xpb = 1024'h2b26a516205b4721d5d13fd37b747d98f6502493c15f9a73be88211ecf714a5616cef8b2579856fd3e252bbdaa403a33bcc6c70dcdecc3f233501e27c38214b74de65653d09c96cc2c5c775d0816cf81f91aba3635e7c546552f0911a52f60eaa097edbc1b0755a0924ea039c3d9c9f51b3146474422c2e7011d665c543a63b9;
    7'b1101000 : xpb = 1024'h7a795fc05e6d12590acbc7fc6b1a364784da2162ebe7f9fc40ab67c91c6e9d4e13867b398d71d86e9ec6ec76c6e2296958ac9f27ab39f3a682b0dec988afa005d99721a5210b998719c274ba6f3b0b510515c09da96198359fa27716eb04be5871905b926a3e5d130b8eb95acc09a3cbcc576764f3d765b6baadeb57cb57fd4e;
    7'b1101001 : xpb = 1024'h191ed514da90a8c774c0d84e4a65a7a4a1ee1b0140f8b90d44f1f51db669433e0cf58047f924db51600a6de9002607d490784f5b65d4530f2172600d130ab6a2f0f8b847c1e99efcf48e6f753d8382ef1d0bcd6c90553e143489532176af79341381373f08ac6bf7fe0eeb9cdc6957792ea3a9a05340ab562dcef54eb9933078;
    7'b1101010 : xpb = 1024'h68718fbf18a273fea9bb60773a0b6053307817d06b811895c7153bc80366963609ad02cf2efe5cc2c0ac2ea21cc7f70a2c5e2775432182c370d320aed83841f17ca983991258a1b7e1f46cd2a4a7bebe2906d3d403cf11037efcc126bc84d6a1e479a51557e3736a774f04bde499314fdfc9cabe02f54e25e75f7a4a30b0ca0d;
    7'b1101011 : xpb = 1024'h717051394c60a6d13b070c91956d1b04d8c116ec091d7a6cb5bc91c9d613c26031c07dd9ab15fa581efb014560bd5756429d7a8fdbbe22c0f94a1f26293588e940b1a3bb336a72dbcc0678d72f0365c40fce0a2eac2b6e213e39d31482f917d866a80c1f651824f69cf36fff4f8e4fd42160cf9625e93c55a8084411eebfd37;
    7'b1101100 : xpb = 1024'h5669bfbdd2d7d5a448aaf8f208fc8a5edc160e3deb1a372f4d7f0fc6ea5e8f1dffd38a64d08ae116e29170cd72adc4ab000fafc2db0911e05ef5629427c0e3dd1fbbe58d03a5a9e8aa2664eada14722b4cf7e70a5e3c89d15e570b368e04eeeb5762ee98458889c1e30f5020fd28bed3f33c2e17121336951411093c960996cc;
    7'b1101101 : xpb = 1024'ha5bc7a6810e9a0db7da5811af8a2430d6aa00b0d15a296b7cfa25671375be215fc8b0cec06646288433331868f4fb3e09bf587dcb8564194ae562335ecee6f2bab6cb0de5414aca3978c62484138adfa58f2ed71d1b65cc0a8ca793bd3da4c59285b5c6e94bf91345c4f6942055898aaa4624f34c1c7d964cda18e380d273061;
    7'b1101110 : xpb = 1024'h4461efbc8d0d3749e79a916cd7edb46a87b404ab6ab355c8d3e8e3c5d1568805f5fa11fa7217656b0476b2f8c893924bd3c1381072f0a0fd4d17a479774985c8c2ce4780f4f2b21972585d030f81259870e8fa40b8aa029f3db155465f850734ca4c381b332da0194ecf9b8415b84c5806ae917021311f0440c2982efb62638b;
    7'b1101111 : xpb = 1024'h93b4aa66cb1f02811c951995c7936d19163e017a953bb551560c2a701e53dafdf2b19481a7f0e6dc651873b1e53581816fa7102a503dd0b19c78651b3c7711174e7f12d24561b4d45fbe5a6076a561677ce400a82c23d58e8824c34ba55a64a29b44a5f18264a78bc80fb4a51de8262eb7d4b28dd0e5c1d3fa531d2a727ffd20;
    7'b1110000 : xpb = 1024'h325a1fbb474298ef868a29e7a6dede763351fb18ea4c74625a52b7c4b84e80edec20999013a3e9bf265bf5241e795feca772c05e0ad8301a3b39e65ec6d227b465e0a974e63fba4a3a8a551b44edd90594da0d7713177b6d1d0b9f5631051f7e3d35819e20d2b670ba8fe6e72e47d9dc1a20f4c9304f07736d74272160bb304a;
    7'b1110001 : xpb = 1024'h81acda6585546426bb84b21096849724c1dbf7e814d4d3eadc75fe6f054bd3e5e8d81c17497d6b3086fdb5dd3b1b4f2243589877e8255fce8a9aa7008bffb302f19174c636aebd0527f05278ac1214d4a0d513de86914e5c677f0d5b76da7cec0e2def747009bde333d000083677b3b2cb4715e6e003aa432704ac1cd7d8c9df;
    7'b1110010 : xpb = 1024'h20524fba0177fa952579c26275d00881deeff18669e592fbe0bc8bc39f4679d5e2472125b5306e134841374f745f2d8d7b2448aba2bfbf37295c2844165ac9a008f30b68d78cc27b02bc4d337a5a8c72b8cb20ad6d84f43afc65e966028537c7b01ecb210e77ccc82650324a46d767602d9358223f6cefe29a25b613c613fd09;
    7'b1110011 : xpb = 1024'h6fa50a643f89c5cc5a744a8b6575c1306d79ee55946df28462dfd26dec43cccddefea3aceb09ef84a8e2f80891011cc3170a20c5800ceeeb78bce8e5db8854ee94a3d6ba27fbc535f0224a90e17ec841c4c62714e0fec72a46d9576b485a9535811738f75daed43a9f904b6b4f074136deb9793fef2192b253b63b0f3d31969e;
    7'b1110100 : xpb = 1024'he4a7fb8bbad5c3ac4695add44c1328d8a8de7f3e97eb19567265fc2863e72bdd86da8bb56bcf2676a26797aca44fb2e4ed5d0f93aa74e54177e6a2965e36b8bac056d5cc8d9caabcaee454bafc73fdfdcbc33e3c7f26d08dbc03375d4055011230814a3fc1ce31f92107dad5f66f4e44105bb7b4e8ad851c6d745062b6cc9c8;
    7'b1110101 : xpb = 1024'h5d9d3a62f9bf2771f963e3063466eb3c1917e4c31407111de949a66cd33bc5b5d5252b428c9673d8cac83a33e6e6ea63eabba91317f47e0866df2acb2b10f6da37b638ae1948cd66b85442a916eb7baee8b73a4b3b6c3ff82633a17b19daad7ef400827a4b53ea920b5096ce6796cebaf22bdc98fe3f7b218067ca01a28a635d;
    7'b1110110 : xpb = 1024'haceff50d37d0f2a92e5e6b2f240ca3eaa7a1e1923e8f70a66b6ced17203918add1dcadc9c26ff54a2b69faed0388d99986a1812cf541adbcb63feb6cf03e8228c36703ff69b7d021a5ba40067e0fb77df4b240b2aee612e770a70f805fb00aecc4f8f0509a8af2048490afef6fc6a891a351fdb6adf41df139f84efd19a7fcf2;
    7'b1110111 : xpb = 1024'h4b956a61b3f4891798537b8103581547c4b5db3093a02fb76fb37a6bba33be9dcb4bb2d82e22f82cecad7c5f3cccb804be6d3160afdc0d2555016cb07a9998c5dac89aa20a95d59780863ac14c582f1c0ca84d8195d9b8c6058deb8aeb5ac5c866e9cbfd38f900e97710e23180265c3f059e3ff20d5d6390ad1958f407e3301c;
    7'b1111000 : xpb = 1024'h9ae8250bf206544ecd4e03a9f2fdcdf6533fd7ffbe288f3ff1d6c11607311195c803355f63fc799e4d4f3d18596ea73a5a53097a8d293cd9a4622d523fc72414667965f35b04d8526dec381eb37c6aeb18a353e909538bb5500159903130233637e239d38830085bf050fb5288563615b6c4610fbd12066066a9ddef7f00c9b1;
    7'b1111001 : xpb = 1024'h398d9a606e29eabd374313fbd2493f537053d19e13394e50f61d4e6aa12bb785c1723a6dcfaf7c810e92be8a92b285a5921eb9ae47c39c424323ae95ca223ab17ddafc95fbe2ddc848b832d981c4e289309960b7f0473193e4e8359abcdade11d9d31580269e1740e2d12d9498b5e9c31910a34b1c7b4bffd9cae7e66d3bfcdb;
    7'b1111010 : xpb = 1024'h88e0550aac3bb5f46c3d9c24c1eef801feddce6d3dc1add978409514ee290a7dbe29bcf50588fdf26f347f43af5474db2e0491c82510cbf692846f378f4fc600098bc7e74c51e083361e3036e8e91e583c94671f63c104832f5ba3a002b03b7faacb835675d51eb35c1146b5a0e5c399ca36c468cc2feecf935b6ce1e4599670;
    7'b1111011 : xpb = 1024'h2785ca5f285f4c62d632ac76a13a695f1bf1c80b92d26cea7c8722698823b06db798c203713c00d5307800b5e898534665d041fbdfab2b5f3145f07b19aadc9d20ed5e89ed2fe5f910ea2af1b73195f6548a73ee4ab4aa61c4427faa8e5af65b4cbc5f0314432d984e9178f7b14577472c8306a42b99346f067c76d8d294c99a;
    7'b1111100 : xpb = 1024'h76d885096671179a0b2d349f90e0220daa7bc4dabd5acc72feaa6913d5210365b450448aa71582469119c16f053a427c01b61a15bcf85b1380a6b11cded867ebac9e29db3d9ee8b3fe50284f1e55d1c560857a55be2e7d510eb5edafd43053c91db4ccd9637a350ac7d19218b975511ddda927c1db4dd73ec00cfbd449b2632f;
    7'b1111101 : xpb = 1024'h157dfa5de294ae08752244f1702b936ac78fbe79126b8b8402f0f6686f1ba955adbf499912c88529525d42e13e7e20e73981ca497792ba7c1f68326069337e88c3ffc07dde7cee29d91c2309ec9e4963787b8724a522232fa39cc9ba5fdb0ea4bfa5a88601e843efba51c45ac9d504cb3ff569fd3ab71cde332e05cb37ed9659;
    7'b1111110 : xpb = 1024'h64d0b50820a6793faa1ccd1a5fd14c195619bb483cf3eb0c85143d12bc18fc4daa76cc2048a2069ab2ff039a5b20101cd567a26354dfea306ec8f3022e6109d74fb08bcf2eebf0e4c682206753c2853284768d8c189bf61eee1037bfa5b06c12909e165c511f4b623391dd7bd204dea1f11b8b1aea6bbfadecbe8ac6af0b2fee;
    7'b1111111 : xpb = 1024'h3762a5c9cca0fae1411dd6c3f1cbd76732db4e69204aa1d895aca675613a23da3e5d12eb455097d7442850c9463ee880d3352970f7a49990d8a7445b8bc207467122271cfc9f65aa14e1b22220afcd09c6c9a5aff8f9bfd82f713ca315b26ee328ef208ef8d5a4726120fbde264924f5367cd5649d5054d5fdf94bd9d466318;
    endcase
end

endmodule

module xpb_5_590
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h60306f7158291071c8ffab3a6b6460b3d251d00bdf4bb35cc9e85703aae034ba386fddfbee8d783616c7141019d7ed730f49dbae721f46d1d91fd156af283ba6a71ac97c44478398936602a23c9efb31184bbd8d798e9cc21757cb40dfdf106b89d497caa6bb08201fae14ede5e1d34a4022281305181d3662d579083dc7c4b1;
    5'b00010 : xpb = 1024'hfb3998cee63ec1ac6f9de9dc66e7a16332d9ce6e91fc64215f3f4b1a2bdbc6c6d973e7f12f471dd8e2fe8d95051ca1bba798f76c18bbd5801a0634f237e029bd9e65e49d8fe09ec143202a1e06232313c92818266970c737923048705937e44e4a19d6b9cad17b2b89c42fcd3f3806b316a7143b9e4dd3c7f3b770bf2ad22f7;
    5'b00011 : xpb = 1024'h6fe408fe468cfc8c8ff989d831d2daca057f6cf2c86b799edfdc4bb54d9df126a6071c7b0181ea13a4f6fce96a29b78ec9c36b2533ab0429dac034a5d2a63e42810127c61d458d84a79805441d012d6254de3f0fe025a935907acfc7e5728eb06e76353643681fd2d84a57eab9d553b5718c9956befcfa72e210f0143074e7a8;
    5'b00100 : xpb = 1024'h1f673319dcc7d8358df3bd3b8cdcf42c665b39cdd23f8c842be7e963457b78d8db2e7cfe25e8e3bb1c5fd1b2a0a3943774f31eed83177ab00340c69e46fc0537b3ccbc93b1fc13d828640543c0c4646279250304cd2e18e6f246090e0b26fc89c9433ad7395a2f65713885f9a7e700d662d4e28773c9ba78fe76ee17e55a45ee;
    5'b00101 : xpb = 1024'h7f97a28b34f0e8a756f36875f84154e038ad09d9b18b3fe0f5d04066f05bad93139e5afa14765bf13326e5c2ba7b81aa843cfa9bf536c181dc6097f4f62440de5ae7860ff6439770bbca07e5fd635f939170c09246bcb5a9099dd44eeb060cf55317d2a1e015378590e69ae78dc8d420a2f70a9a78e1d7af614c672023220a9f;
    5'b00110 : xpb = 1024'h2f1acca6cb2bc45054ed9bd9534b6e429988d6b4bb5f52c641dbde14e839354548c5bb7d38dd5598aa8fba8bf0f55e532f6cae6444a3380804e129ed6a7a07d38db31add8afa1dc43c9607e5a1269693b5b7848733c5255a6b690d9510ba7aceade4d842d607471829d4c8f67bda8141943f53cb2dae97b57db26523d80768e5;
    5'b00111 : xpb = 1024'h8f4b3c182354d4c21ded4713beafcef66bdaa6c09aab06230bc43518931969ff81359979276acdcec156ce9c0acd4bc63eb68a12b6c27ed9de00fb4419a2437a34cde459cf41a15ccffc0a87ddc591c4ce034214ad53c21c82c0d8d5f0998b3a37b9700d7cc24f384982dde461bc548bd4617bde32c6b4ebe087de2c15cf2d96;
    5'b01000 : xpb = 1024'h3ece6633b98fb06b1be77a7719b9e858ccb6739ba47f190857cfd2c68af6f1b1b65cf9fc4bd1c77638bfa3654147286ee9e63ddb062ef56006818d3c8df80a6f6799792763f827b050c80a878188c8c4f24a06099a5c31cde48c121c164df913928675ae72b45ecae2710bf34fce01acc5a9c50ee79374f1fceddc2fcab48bdc;
    5'b01001 : xpb = 1024'h9efed5a511b8c0dce4e725b1851e490c9f0843a783cacc6521b829ca35d7266beeccd7f83a5f3fac4f86b7755b1f15e1f9301989784e3c31dfa15e933d2046160eb442a3a83fab48e42e0d29be27c3f60a95c39713eace8ffbe3dd5cf62d097f1c5b0d79196f66eb021f20e135afd4f705cbed21ecab92285fc35538087c508d;
    5'b01010 : xpb = 1024'h4e81ffc0a7f39c85e2e15914e028626effe410828d9edf4a6dc3c7782db4ae1e23f4387b5ec63953c6ef8c3e9198f28aa45fcd51c7bab2b80821f08bb1760d0b417fd7713cf6319c64fa0d2961eafaf62edc878c00f33e415daf16a31be177587728131a0f61767d9b0d4ef023c18217f7143652a178522e7c29533bbd61aed3;
    5'b01011 : xpb = 1024'haeb26f32001cacf7abe1044f4b8cc322d235e08e6cea92a737ac1e7bd894e2d85c6416774d53b189ddb6a04eab70dffdb3a9a90039d9f989e141c1e2609e48b1e89aa0ed813db534f8600fcb9e89f627472845197a81db037506e1e3fbc087c400fcaae4b61c7e9dbabb63de09a3556237365e65a6906f64defecc43fb297384;
    5'b01100 : xpb = 1024'h5e35994d965788a0a9db37b2a696dc853311ad6976bea58c83b7bc29d0726a8a918b76fa71baab31551f7517e1eabca65ed95cc88946701009c253dad4f40fa71b6635bb15f43b88792c0fcb424d2d276b6f090e678a4ab4d6d21b2a2174f59d5bc9b085ac0e8e3053a991ecf7b50283287ea7965b5d2f6afb64ca47b00ed1ca;
    5'b01101 : xpb = 1024'hdb8c3692c926449a7d56b1601a0f5e793ed7a448092b871cfc359d7c84ff23cc6b2d77d9621a4d8cc8849e11864994f0a091090d8b2e6963242e5d34949d69c4e31ca88aaaac1dbf9f80fcae61064278fb5cd035492ba66389d547047296376b696b626a2009dc2ec97bffbe5c6afa419c6f0c71029ef7117cac84b64f43010;
    5'b01110 : xpb = 1024'h6de932da84bb74bb70d516506d05569b663f4a505fde6bce99abb0db733026f6ff22b57984af1d0ee34f5df1323c86c21952ec3f4ad22d680b62b729f8721242f54c9404eef245748d5e126d22af5f58a8018a90ce2157284ff51fb1270873e2406b4df148bba5e30c45d4e9cba882ee59e918da15420ca77aa04153a2bbf4c1;
    5'b01111 : xpb = 1024'h1d6c5cf61af650646ecf49b3c80f6ffdc71b172b69b27eb3e5b74e896b0daea9344a15fca91616b65ab832ba68b6636ac482a0079a3ea3ee33e349226cc7d938281828d283a8cbc80e2a126cc6729658cc484e85bb29c6d9b1c058f74cbce1bb9b3853923eadb575a53402f8b9ba300f4b31620aca0eccad97063f5757a15307;
    5'b10000 : xpb = 1024'h7d9ccc67731f60d637cef4ee3373d0b1996ce73748fe3210af9fa58d15ede3636cb9f3f897a38eec717f46ca828e50ddd3cc7bb60c5deac00d031a791bf014decf32f24ec7f04f60a190150f03119189e4940c1334b8639bc91824382c9bf227250ceb5ce568bd95c4e217e69f9c03598b538a1dcf26e9e3f9dbb85f956917b8;
    5'b10001 : xpb = 1024'h2d1ff683095a3c7f35c928518e7dea13fa48b41252d244f5fbab433b0dcb6b15a1e1547bbc0a8893e8e81b93b9082d867efc2f7e5bca61463583ac719045dbd401fe871c5ca6d5b4225c150ea6d4c88a08dad00821c0d34d2ae35d7e525060007fd9f0fddb5acd285dd045f58dadb07a7c9bd34e83f3a9ea1641b6634a4e75fe;
    5'b10010 : xpb = 1024'h8d5065f461834cf0fec8d38bf9e24ac7cc9a841e321df852c5939a3eb8ab9fcfda513277aa9800c9ffaf2fa3d2e01af98e460b2ccde9a8180ea37dc83f6e177aa9195098a0ee594cb5c217b0e373c3bb21268d959b4f700f423b28bf322f706c09ae88c88215d5487d7e5ae3738f83c4bcbdfb61890bc72079172f6b88163aaf;
    5'b10011 : xpb = 1024'h3cd3900ff7be2899fcc306ef54ec642a2d7650f93bf20b38119f37ecb08927820f7892facefefa717718046d0959f7a23975bef51d561e9e37240fc0b3c3de6fdbe4e56635a4dfa0368e17b08736fabb456d518a8857dfc0a406620557e3de45647b8e697807e4db166c88f261a130e5ae0644923dd88726957d2d6f3cfb98f5;
    5'b10100 : xpb = 1024'h9d03ff814fe7390bc5c2b229c050c4ddffc821051b3dbe94db878ef05b695c3c47e870f6bd8c72a78ddf187d2331e51548bf9aa38f7565701043e11762ec1a1682ffaee279ec6338c9f41a52c3d5f5ec5db90f1801e67c82bb5e2d4637c2eeb0ee5026341ec2ecfb361a9de04783042fee286ca542f0a45cf852a6777ac35da6;
    5'b10101 : xpb = 1024'h4c87299ce62214b4c3bce58d1b5ade4060a3ede02511d17a27932c9e5346e3ee7d0fd179e1f36c4f0547ed4659abc1bdf3ef4e6bdee1dbf638c4730fd741e10bb5cb43b00ea2e98c4ac01a5267992cec81ffd30ceeeeec341d29668c5d775c8a491d2bd514b4fc8dcf08cbef3594b150df70b5d5f7bd646314b8a47b2fa8bbec;
    5'b10110 : xpb = 1024'hacb7990e3e4b25268cbc90c786bf3ef432f5bdec045d84d6f17b83a1fe2718a8b57faf75d080e4851c0f01567383af3103392a1a510122c811e44466866a1cb25ce60d2c52ea6d24de261cf4a438281d9a4b909a687d88f6348131cd3d566cf5d2f1c39fbb7004adeeb6e0dd1b76849b1f92dde8fcd58199778e1d836d70809d;
    5'b10111 : xpb = 1024'h5c3ac329d48600cf8ab6c42ae1c9585693d18ac70e3197bc3d87214ff604a05aeaa70ff8f4e7de2c9377d61fa9fd8bd9ae68dde2a06d994e3a64d65efabfe3a78fb1a1f9e7a0f3785ef21cf447fb5f1dbe92548f5585f8a7964c6b13630adacf2dbec940b162144087a50eec098831bc10db2719b1a2419f93f41b872255dee3;
    5'b11000 : xpb = 1024'hbbded456ac0dc7888b0f78e3cd371b8f4ad57a21805aaa18992befdede2280d1fce707c194ed7d40ae0aae8e0776882599891aaefda0fd462e568576f15aa9cc27d36c77c5779cbdfbe1cf3ebbe961de2d91884428e6858f817a45988bf48a8888bcee1a75423d320933cfaf799dedd0223704a666f01a5b05a198ad73b3d29;
    5'b11001 : xpb = 1024'h6bee5cb6c2e9ecea51b0a2c8a837d26cc6ff27adf7515dfe537b160198c25cc7583e4e7807dc500a21a7bef8fa4f55f568e26d5961f956a63c0539ae1e3de64369980043c09efd6473241f96285d914efb24d611bc1d051b0f6f6f9a689e5914126066ac4e0f2bf3404151e8dd7bb2274245985d6b871edc132f9293150301da;
    5'b11010 : xpb = 1024'h1b7186d25924c8934faad62c0341ebcf27daf489012570e39f86b3af909fe4798d65aefb2c4349b1991093c230c9329e14122121b165cd2c6485cba69293ad389c639511555583b7f3f01f95cc20c84f1f6b9a06a92574cc713aa8e08e52c6ed6d2d6c4d44013b85d92f7ff7cb8d5f48338de18e2053dee22f959096c9e86020;
    5'b11011 : xpb = 1024'h7ba1f643b14dd90518aa81666ea64c82fa2cc494e0712440696f0ab33b801933c5d58cf71ad0c1e7afd7a7d24aa12011235bfcd0238513fe3da59cfd41bbe8df437e5e8d999d07508756223808bfc38037b7579422b4118e889274216e31d758f7020417eabc43a5f8dd94e5b16f329273b009a1256bfc18926b099f07b024d1;
    5'b11100 : xpb = 1024'h2b25205f4788b4ae16a4b4c9c9b065e55b08916fea453725b57aa861335da0e5fafced7a3f37bb8f27407c9b811afcb9ce8bb09872f18a8466262ef5b611afd47649f35b2e538da408222237ac82fa805bfe1b890fbc813fea5dad6793e6453251cf09b8e0ae533891cbc2f49f80dfb364f852d1da38bc1eaed107a2bc958317;
    5'b11101 : xpb = 1024'h8b558fd09fb1c51fdfa460043514c6992d5a617bc990ea827f62ff64de3dd5a0336ccb762dc533c53e0790ab9af2ea2cddd58c46e510d1563f46004c6539eb7b1d64bcd7729b113c9b8824d9e921f5b17449d916894b1e0201b578a873c5559ddba3a18387695b58b179d7e28562b2fda51a7ae4df50d95511a680aafa5d47c8;
    5'b11110 : xpb = 1024'h3ad8b9ec35eca0c8dd9e9367901edffb8e362e56d364fd67cb6e9d12d61b5d5268942bf9522c2d6cb5706574d16cc6d58905400f347d47dc67c69244d98fb270503051a5075197901c5424d98ce52cb198909d0b76538db36380b1ee9979c3773670a7247d5b6aeb4a6805f17374601e9662c415941d995b2e0c7eaeaf42a60e;
    5'b11111 : xpb = 1024'h9b09295d8e15b13aa69e3ea1fb8340af6087fe62b2b0b0c49556f41680fb920ca10409f540b9a5a2cc377984eb44b448984f1bbda69c8eae40e6639b88b7ee16f74b1b214b991b28afba277bc98427e2b0dc5a98efe22a757ad87d2f7958d3e2c0453eef2416730b6a161adf59563368d684ec289935b69190e1f7b6ed0a6abf;
    endcase
end

endmodule

module xpb_5_235
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h8b1a15ffa4d817436e8bddea832bf7f1bb8661f1d5a068aadfcc228b72a4f4f640d6976eb984e10902f992075f1d4a56d1c1ccf73bd40c7437e51632e238abd9eac2ec645c177d54801c80b451101aa115675688d7c0292874e10366e0e56a3b1523b4bcfe590c0ac13a086846893b1582bcaa6f8d64fe58d9a1871c35ff5d7;
    5'b00010 : xpb = 1024'h116342bff49b02e86dd17bbd50657efe3770cc3e3ab40d155bf984516e549e9ec81ad2edd7309c21205f3240ebe3a94ada38399ee77a818e86fca2c65c47157b3d585d8c8b82efaa900390168a22035422acead11af805250e9c206cdc1cad4762a476979fcb21815827410d08d12762b057954df1ac9fcb1b3430e386bfebae;
    5'b00011 : xpb = 1024'h1a14e41feee8845ca4ba399bf8983e7d5329325d580e13a009f6467a257eedee2c283c64c2c8ea31b08ecb6161d57df04754566e5b37c255ca7af4298a6aa038dc048c52d144677fd8055821cf3304fe34036039a87407b795ea30a34a2b03eb13f6b1e36fb0b242043ae1938d39bb1408835ff4ea82efb0a8ce49554a1fe185;
    5'b00100 : xpb = 1024'h22c6857fe93605d0dba2f77aa0cafdfc6ee1987c75681a2ab7f308a2dca93d3d9035a5dbae61384240be6481d7c75295b470733dcef5031d0df9458cb88e2af67ab0bb191705df552007202d144406a84559d5a235f00a4a1d3840d9b8395a8ec548ed2f3f964302b04e821a11a24ec560af2a9be3593f96366861c70d7fd75c;
    5'b00101 : xpb = 1024'h2b7826dfe3838745128bb55948fdbd7b8a99fe9b92c220b565efcacb93d38c8cf4430f5299f98652d0edfda24db9273b218c900d42b243e4517796efe6b1b5b4195ce9df5cc7572a6808e8385955085256b04b0ac36c0cdca48651102647b132769b287b0f7bd3c35c6222a0960ae276b8daf542dc2f8f7bc4027a38d0dfcd33;
    5'b00110 : xpb = 1024'h3429c83fddd108b949747337f1307cfaa65264bab01c274013ec8cf44afddbdc585078c98591d463611d96c2c3aafbe08ea8acdcb66f84ab94f5e85314d54071b80918a5a288ceffb00ab0439e6609fc6806c07350e80f6f2bd46146945607d627ed63c6df6164840875c3271a7376281106bfe9d505df61519c92aa943fc30a;
    5'b00111 : xpb = 1024'h3cdb699fd81e8a2d805d311699633c79c20acad9cd762dcac1e94f1d02282b2bbc5de240712a2273f14d2fe3399cd085fbc4c9ac2a2cc572d87439b642f8cb2f56b5476be84a46d4f80c784ee3770ba6795d35dbde641201b322717d02645e79d93f9f12af46f544b48963ad9edc09d969328a90cddc2f46df36ab1c579fb8e1;
    5'b01000 : xpb = 1024'h458d0affd26c0ba1b745eef54195fbf8ddc330f8ead034556fe61145b9527a7b206b4bb75cc27084817cc903af8ea52b68e0e67b9dea063a1bf28b19711c55ecf56176322e0bbeaa400e405a28880d508ab3ab446be014943a7081b37072b51d8a91da5e7f2c8605609d043423449d8ac15e5537c6b27f2c6cd0c38e1affaeb8;
    5'b01001 : xpb = 1024'h4e3eac5fccb98d15ee2eacd3e9c8bb77f97b9718082a3ae01de2d36e707cc9ca8478b52e485abe9511ac6224258079d0d5fd034b11a747015f70dc7c9f3fe0aa940da4f873cd367f881008656d990efa9c0a20acf95c1726c1be91e9de810bc13be415aa4f1216c60cb0a4baa7ad313c198a1fdebf88cf11fa6adbffde5fa48f;
    5'b01010 : xpb = 1024'h56f04dbfc7070e8a25176ab291fb7af71533fd372584416acbdf959727a71919e8861ea533f30ca5a1dbfb449b724e764319201a856487c8a2ef2ddfcd636b6832b9d3beb98eae54d011d070b2aa10a4ad60961586d819b9490ca2204c8f6264ed3650f61ef7a786b8c445412c15c4ed71b5ea85b85f1ef78804f471a1bf9a66;
    5'b01011 : xpb = 1024'h5fa1ef1fc1548ffe5c0028913a2e3a7630ec635642de47f579dc57bfded168694c93881c1f8b5ab6320b94651164231bb0353ce9f921c88fe66d7f42fb86f625d1660284ff50262a1813987bf7bb124ebeb70b7e14541c4bd05ab256ba9db9089e888c41eedd384764d7e5c7b07e589ec9e1b52cb1356edd159f0ce3651f903d;
    5'b01100 : xpb = 1024'h6853907fbba2117292e8e66fe260f9f54ca4c97560384e8027d919e895fbb7b8b0a0f1930b23a8c6c23b2d858755f7c11d5159b96cdf095729ebd0a629aa80e37012314b45119dff601560873ccc13f8d00d80e6a1d01ede57a8c28d28ac0fac4fdac78dbec2c90810eb864e34e6ec50220d7fd3aa0bbec2a3392555287f8614;
    5'b01101 : xpb = 1024'h710531dfb5ef92e6c9d1a44e8a93b974685d2f947d92550ad5d5dc114d26070814ae5b09f6bbf6d7526ac6a5fd47cc668a6d7688e09c4a1e6d6a220957ce0ba10ebe60118ad315d4a817289281dd15a2e163f64f2f4c2170def6d2c396ba6650012d02d98ea859c8bcff26d4b94f80017a394a7aa2e20ea830d33dc6ebdf7beb;
    5'b01110 : xpb = 1024'h79b6d33fb03d145b00ba622d32c678f3841595b39aec5b9583d29e3a0450565778bbc480e25444e7e29a5fc67339a10bf789935854598ae5b0e8736c85f1965ead6a8ed7d0948da9f018f09dc6ee174cf2ba6bb7bcc824036644e2fa04c8bcf3b27f3e255e8dea896912c75b3db813b2d26515219bb85e8dbe6d5638af3f71c2;
    5'b01111 : xpb = 1024'h8268749faa8a95cf37a3200bdaf938729fcdfbd2b846622031cf6062bb7aa5a6dcc92df7cdec92f872c9f8e6e92b75b164a5b027c816cbacf466c4cfb415211c4c16bd9e1656057f381ab8a90bff18f70410e1204a442695ed92f33072d7139763d179712e737b4a152667e1c220a7642a90dfc8948eae734c076eaa729f6799;
    5'b10000 : xpb = 1024'h8b1a15ffa4d817436e8bddea832bf7f1bb8661f1d5a068aadfcc228b72a4f4f640d6976eb984e10902f992075f1d4a56d1c1ccf73bd40c7437e51632e238abd9eac2ec645c177d54801c80b451101aa115675688d7c0292874e10366e0e56a3b1523b4bcfe590c0ac13a086846893b1582bcaa6f8d64fe58d9a1871c35ff5d70;
    5'b10001 : xpb = 1024'h93cbb75f9f2598b7a5749bc92b5eb770d73ec810f2fa6f358dc8e4b429cf4445a4e400e5a51d2f1993292b27d50f1efc3edde9c6af914d3b7b636796105c3697896f1b2aa1d8f529c81e48bf96211c4b26bdcbf1653c2bbafc2f139d4ef3c0dec675f008ce3e9ccb6d4da8eecaf1cec6dae87516863b4e3e673b9f8df95f5347;
    5'b10010 : xpb = 1024'h9c7d58bf99731a2bdc5d59a7d39176eff2f72e30105475c03bc5a6dce0f9939508f16a5c90b57d2a2358c4484b00f3a1abfa0696234e8e02bee1b8f93e7fc155281b49f0e79a6cff102010cadb321df538144159f2b82e4d837d23d3bd02178277c82b549e242d8c196149754f5a627833143fbd7f119e23f4d5b7ffbcbf491e;
    5'b10011 : xpb = 1024'ha52efa1f93c09ba0134617867bc4366f0eaf944f2dae7c4ae9c269059823e2e46cfed3d37c4dcb3ab3885d68c0f2c84719162365970bceca02600a5c6ca34c12c6c778b72d5be4d45821d8d620431f9f496ab6c2803430e00acb340a2b106e26291a66a06e09be4cc574e9fbd3c2f6298b400a6477e7ee09826fd071801f3ef5;
    5'b10100 : xpb = 1024'hade09b7f8e0e1d144a2ed56523f6f5ee2a67fa6e4b0882d597bf2b2e4f4e3233d10c3d4a67e6194b43b7f68936e49cec863240350ac90f9145de5bbf9ac6d6d06573a77d731d5ca9a023a0e1655421495ac12c2b0db0337292194440991ec4c9da6ca1ec3def4f0d71888a82582b89dae36bd50b70be3def1009e8e3437f34cc;
    5'b10101 : xpb = 1024'h5e4f789c66d69bfb6121b6cbbcf6e1bd4aa5d5c92eae8e8c7df34015375d47b31d129488957e8cd34895062c97860c78f34351e5bd3800cd8bd6dc48e17ecdc8fd0a195094dd739d58b664a11895ec27812a7fb0ea608f463dac27c4d0278db5cb74b0e5d0be74096dc4429e4c3f762ecbdc0d0194930a4573486507dfcc438;
    5'b10110 : xpb = 1024'he9698e9c0baeb33ecfad94b64022d9af062c37bb044ef7375dbf62a0aa023ca95de92bf74f036ddc4b8e9833f6a356cfc5051edcf90c0d41c3bbf27bc3b779a2e7cd05b4f0f4f0f1d8d2e55569a606c89691d639c220b86eb28d2b2bb10cf7f0e09865a2cf1780142efe4b0692c8b1444e98b77121f8089e4ce9ec2415cba0f;
    5'b10111 : xpb = 1024'h17483a49bb086ca823e3972a0c34ed1a0c1b299acd9ef5fe23d8b852c1ca7319f9ebfc36608884ee54e882a3b55c0a12696c6ebd434e019b5fba108aea5f0257cd28ff2194d0c6e4658ef6609bab62169abf92cc299e0e197276e2e9291f2622bf5bc1a5fcd708c1ef038536ed951ec59d15561e0af5d06f7268b73404bcafe6;
    5'b11000 : xpb = 1024'h1ff9dba9b555ee1c5acc5508b467ac9927d38fb9eaf8fc88d1d57a7b78f4c2695df965ad4c20d2fee5181bc42b4ddeb7d6888b8cb70b4262a33861ee18828d156bd52de7da923eb9ad90be6be0bc63c0ac160834b71a10abf9c4f31f972d7cc670adfcf1ccbc99829b1725bd71fdb276f54120c503cc20550002cfa5c81ca5bd;
    5'b11001 : xpb = 1024'h28ab7d09afa36f9091b512e75c9a6c18438bf5d9085303137fd23ca4301f11b8c206cf2437b9210f7547b4e4a13fb35d43a4a85c2ac88329e6b6b35146a617d30a815cae2053b68ef592867725cd656abd6c7d9d4496133e81130356053bd36a2200383d9ca22a43472ac643f66646284d6ceb6bfca2703a8d9ce8178b7c9b94;
    5'b11010 : xpb = 1024'h315d1e69a9f0f104c89dd0c604cd2b975f445bf825ad099e2dcefecce74961082614389b23516f2005774e0517318802b0c0c52b9e85c3f12a3504b474c9a290a92d8b7466152e643d944e826ade6714cec2f305d21215d10861138c734a2a0dd35273896c87bb03f33e66ca7aced9d9a598b612f578c0201b3700894edc916b;
    5'b11011 : xpb = 1024'h3a0ebfc9a43e7278ff868ea4acffeb167afcc21743071028dbcbc0f59e73b0578a21a2120ee9bd3095a6e7258d235ca81ddce1fb124304b86db35617a2ed2d4e47d9ba3aabd6a6398596168dafef68bee019686e5f8e18638faf23c2e15880b184a4aed53c6d4bc49f520750ff376d8afdc480b9ee4f1005a8d118fb123c8742;
    5'b11100 : xpb = 1024'h42c061299e8bf3ed366f4c835532aa9596b52836606116b389c8831e559dffa6ee2f0b88fa820b4125d680460315314d8af8feca8600457fb131a77ad110b80be685e900f1981e0ecd97de98f5006a68f16fddd6ed0a1af616fd33f94f66d75535f6ea210c52dc854b65a7d783a0013c55f04b60e7255feb366b316cd59c7d19;
    5'b11101 : xpb = 1024'h4b72028998d975616d580a61fd656a14b26d8e557dbb1d3e37c545470cc84ef6523c74ffe61a5951b6061966790705f2f8151b99f9bd8646f4aff8ddff3442c9853217c7375995e41599a6a43a116c1302c6533f7a861d889e4b442fbd752df8e749256cdc386d45f779485e080894edae1c1607dffbafd0c40549de98fc72f0;
    5'b11110 : xpb = 1024'h5423a3e99326f6d5a440c840a5982993ce25f4749b1523c8e5c2076fc3f29e45b649de76d1b2a7624635b286eef8da98653138696d7ac70e382e4a412d57cd8723de468d7d1b0db95d9b6eaf7f226dbd141cc8a80802201b259954662b83849c989b60b8ac1dfe06a38ce8e48c71289f0647e0aed8d1ffb6519f62505c5c68c7;
    5'b11111 : xpb = 1024'h5cd545498d747849db29861f4dcae912e9de5a93b86f2a5393bec9987b1ced951a5747edbd4af572d6654ba764eaaf3dd24d5538e13807d57bac9ba45b7b5844c28a7553c2dc858ea59d36bac4336f6725733e10957e22adace7649c9991db4049ed9c047c038ec74fa0896b10d9bc505e73ab55d1a84f9bdf397ac21fbc5e9e;
    endcase
end

endmodule

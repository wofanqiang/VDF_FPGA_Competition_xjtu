module xpb_5_160
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h1bf4deba50d6b45599c09d25e28d7fda4db3010a8a866f4bf5437276aa03177e70ba62db8de3952d32ac1c2394c02c060c71043b0513918e275ac7825049c45d296d201131c91503bb27701843fd34945b9529c6bf39bc536edd363f47ce8cf5fd18ed5e72c5bc64b3becd289c253727fe6fbccd0e0c5574188344ca1aa51614;
    5'b00010 : xpb = 1024'h37e9bd74a1ad68ab33813a4bc51affb49b660215150cde97ea86e4ed54062efce174c5b71bc72a5a655838472980580c18e208760a27231c4eb58f04a09388ba52da402263922a07764ee03087fa6928b72a538d7e7378a6ddba6c7e8f9d19ebfa31dabce58b78c9677d9a51384a6e4ffcdf799a1c18aae831068994354a2c28;
    5'b00011 : xpb = 1024'h53de9c2ef2841d00cd41d771a7a87f8ee919031f9f934de3dfca5763fe09467b522f2892a9aabf879804546abe40841225530cb10f3ab4aa76105686f0dd4d177c476033955b3f0b31765048cbf79dbd12bf7d543dad34fa4c97a2bdd76ba6e1f74ac81b5851352e1b3c6779d46fa577fb4f36672a25005c4989ce5e4fef423c;
    5'b00100 : xpb = 1024'h6fd37ae9435ad156670274978a35ff6936cc042a2a19bd2fd50dc9daa80c5df9c2e98b6e378e54b4cab0708e5300b01831c410ec144e46389d6b1e0941271174a5b48044c724540eec9dc0610ff4d2516e54a71afce6f14dbb74d8fd1f3a33d7f463b579cb16f192cefb34a27094dc9ff9bef334383155d0620d13286a945850;
    5'b00101 : xpb = 1024'h8bc859a3943185ac00c311bd6cc37f43847f0534b4a02c7bca513c51520f757833a3ee49c571e9e1fd5c8cb1e7c0dc1e3e3515271961d7c6c4c5e58b9170d5d1cf21a055f8ed6912a7c5307953f206e5c9e9d0e1bc20ada12a520f3c6708c0cdf17ca2d83ddcadf782ba01cb0cba13c7f82eb001463dab447a9057f285396e64;
    5'b00110 : xpb = 1024'ha7bd385de5083a019a83aee34f50ff1dd232063f3f269bc7bf94aec7fc128cf6a45e512553557f0f3008a8d57c8108244aa619621e756954ec20ad0de1ba9a2ef88ec0672ab67e1662eca09197ef3b7a257efaa87b5a69f4992f457baed74dc3ee959036b0a26a5c3678cef3a8df4aeff69e6cce544a00b893139cbc9fde8478;
    5'b00111 : xpb = 1024'h1304d1c273f0b98e693ed432218437a6ae6f0418f4356a9c36fb67e8f312f76d11d03688171295adc35685b22de3235ff2fcf5b700d62a9762dc3531f731e9daadacabc9acee95d50b7a0e074310abdd8d0f2ad6ae0df937527fe9c03c7b3827bca6eb6b729f2e336377b53d4d345beea6344ab9120af8fc6527668231a13421;
    5'b01000 : xpb = 1024'h2ef9b07cc4c76de402ff71580411b780fc2205237ebbd9e82c3eda5f9d160eeb828a9963a4f62adaf602a1d5c2a34f65ff6df9f205e9bc258a36fcb4477bae37d719cbdadeb7aad8c6a17e1f870de071e8a4549d6d47b58ac15d1fff8449c51db9bfd8c9e564ea9817368265e9599316a4a4078620174e707daaab4c4c464a35;
    5'b01001 : xpb = 1024'h4aee8f37159e22399cc00e7de69f375b49d5062e0942493421824cd647192669f344fc3f32d9c00828aebdf957637b6c0bdefe2d0afd4db3b191c43697c572950086ebec1080bfdc81c8ee37cb0b150644397e642c8171de303a563ecc185213b6d8c628582aa6fccaf54f8e857eca3ea313c4532e23a3e4962df01666eb6049;
    5'b01010 : xpb = 1024'h66e36df16674d68f3680aba3c92cb7359788073893c8b88016c5bf4cf11c3de863ff5f1ac0bd55355b5ada1cec23a772185002681010df41d8ec8bb8e80f36f229f40bfd4249d4e03cf05e500f08499a9fcea82aebbb2e319f178c7e13e6df09b3f1b386caf063617eb41cb721a40166a18381203c2ff958aeb134e08190765d;
    5'b01011 : xpb = 1024'h82d84cabb74b8ae4d04148c9abba370fe53b08431e4f27cc0c0931c39b1f5566d4b9c1f64ea0ea628e06f64080e3d37824c106a3152470d00047533b3858fb4f53612c0e7412e9e3f817ce6853057e2efb63d1f1aaf4ea850df4c2bd5bb56bffb10aa0e53db61fc63272e9dfbdc9388e9ff33ded4a3c4eccc73479aa9c358c71;
    5'b01100 : xpb = 1024'h9ecd2b6608223f3a6a01e5ef8e47b6ea32ee094da8d59718014ca43a45226ce5457424d1dc847f8fc0b3126415a3ff7e31320ade1a38025e27a21abd88a2bfac7cce4c1fa5dbfee7b33f3e809702b2c356f8fbb86a2ea6d87cd1f8fca383f8f5ae238e43b07bdc2ae631b70859ee6fb69e62faba5848a440dfb7be74b6daa285;
    5'b01101 : xpb = 1024'ha14c4ca970abec738bd0b3e607aef730f2b07275de465ec78b35d5b3c22d75bb2e60a34a041962e5400ef40c7061ab9d988e732fc98c3a09e5da2e19e1a0f5831ec3782281416a65bccabf642242326be892be69ce2361b36229d413127e3597c34e9787278a00213309d51fe4380b54df8d8a516099c84b1cb883a489d522e;
    5'b01110 : xpb = 1024'h2609a384e7e1731cd27da86443086f4d5cde0831e86ad5386df6cfd1e625eeda23a06d102e252b5b86ad0b645bc646bfe5f9eb6e01ac552ec5b86a63ee63d3b55b59579359dd2baa16f41c0e862157bb1a1e55ad5c1bf26ea4ffd38078f6704f794dd6d6e53e5c66c6ef6a7a9a68b7dd4c6895722415f1f8ca4ecd0463426842;
    5'b01111 : xpb = 1024'h41fe823f38b827726c3e458a2595ef27aa91093c72f14484633a424890290658945acfebbc08c088b9592787f08672c5f26aefa906bfe6bced1331e63ead981284c677a48ba640add21b8c26ca1e8c4f75b37f741b55aec213dd09bfc0c4fd457666c435580418cb7aae37a3368def054ad8523f3222476ce2d211ce7de77e56;
    5'b10000 : xpb = 1024'h5df360f9898edbc805fee2b008236f01f8440a46fd77b3d0587db4bf3a2c1dd7051532c749ec55b5ec0543ab85469ecbfedbf3e40bd3784b146df9688ef75c6fae3397b5bd6f55b18d42fc3f0e1bc0e3d148a93ada8f6b1582ba3fff08938a3b737fb193cac9d5302e6d04cbd2b3262d49480f0c402e9ce0fb555698988c946a;
    5'b10001 : xpb = 1024'h79e83fb3da65901d9fbf7fd5eab0eedc45f70b5187fe231c4dc12735e42f355575cf95a2d7cfeae31eb15fcf1a06cad20b4cf81f10e709d93bc8c0eadf4120ccd7a0b7c6ef386ab5486a6c575218f5782cddd30199c92768f197763e5062173170989ef23d8f9194e22bd1f46ed85d5547b7cbd94e3af25513d89b62b331aa7e;
    5'b10010 : xpb = 1024'h95dd1e6e2b3c447339801cfbcd3e6eb693aa0c5c12849268430499ac8e324cd3e689f87e65b38010515d7bf2aec6f6d817bdfc5a15fa9b676323886d2f8ae52a010dd7d821017fb90391dc6f96162a0c8872fcc85902e3bc6074ac7d9830a4276db18c50b0554df995ea9f1d0afd947d462788a65c4747c92c5be02ccdd6c092;
    5'b10011 : xpb = 1024'h124b7d2ba24c400083b424a9f71a73f6fe70a35c793613cba6b52cd8532b74a53fbdde1297096aee4ab58cf60291213c014d8aef85b5ca9d9df1091450234d5b62bc33aa3399777ac1f49e541379a6ff0032cf68bb672ff19c550c225d48e8b3bc2e785725211d0c2e98566af52a57bf5bd66911a08400cfe6fa9f25f99703b;
    5'b10100 : xpb = 1024'h1d19968d0afb7855a1fbdf7081ff2719bd9a0b405219d088afaec5442f35cec8c4b640bcb7542bdc175774f2f4e93e19cc85dce9fd6eee380139d813954bf932df98e34bd502ac7b6746b9fd8534cf044b9856bd4af02f5288a287016da31b8138dbd4e3e517ce3576a8528f4b77dca3f42d235e2814958116f2eebc7a3e864f;
    5'b10101 : xpb = 1024'h390e75475bd22cab3bbc7c96648ca6f40b4d0c4adca03fd4a4f237bad938e6473570a3984537c1094a03911689a96a1fd8f6e12502827fc628949f95e595bd900906035d06cbc17f226e2a15c9320398a72d80840a29eba5f77fbd40b571a87735f4c24257dd8a9a2a671fb7e79d13cbf29ce02b3620eaf52f76338694e39c63;
    5'b10110 : xpb = 1024'h55035401aca8e100d57d19bc471a26ce59000d556726af209a35aa31833bfdc5a62b0673d31b56367cafad3a1e699625e567e560079611544fef671835df81ed3273236e3894d682dd959a2e0d2f382d02c2aa4ac963a7f9665cf37ffd40356d330dafa0caa346fede25ece083c24af3f10c9cf8442d406947f97850af88b277;
    5'b10111 : xpb = 1024'h70f832bbfd7f95566f3db6e229a7a6a8a6b30e5ff1ad1e6c8f791ca82d3f154416e5694f60feeb63af5bc95db329c22bf1d8e99b0ca9a2e2774a2e9a8629464a5be0437f6a5deb8698bd0a46512c6cc15e57d411889d644cd53a29bf450ec26330269cff3d69036391e4ba091fe7821bef7c59c5523995dd607cbd1aca2dc88b;
    5'b11000 : xpb = 1024'h8ced11764e5649ac08fe54080c352682f4660f6a7c338db884bc8f1ed7422cc2879fcc2aeee28090e207e58147e9ee31fe49edd611bd34709ea4f61cd6730aa7854d63909c27008a53e47a5e9529a155b9ecfdd847d720a044175ffe8cdd4f592d3f8a5db02ebfc845a38731bc0cb943edec16926045eb51790001e4e4d2de9f;
    5'b11001 : xpb = 1024'ha8e1f0309f2cfe01a2bef12deec2a65d4219107506b9fd047a00019581454440f85a2f067cc615be14b401a4dcaa1a380abaf21116d0c5fec5ffbd9f26bccf04aeba83a1cdf0158e0f0bea76d926d5ea1582279f0710dcf3b2f4963dd4abdc4f2a5877bc22f47c2cf962545a5831f06bec5bd35f6e5240c5918346aeff77f4b3;
    5'b11010 : xpb = 1024'h142989952e157d8e717a167cc0f5dee61e560e4ebbc8cbd8f166bab67845aeb765cc146940832c5ca801de818e0c3573b311ce65f93187413cbb45c33c341eb063d86f0450282d4cb79957ec8448464d7d1257cd39c46c366c453a82624fc6b2f869d2f0e4f1400426613aa3fc87016a9bf1b14a2c13390963971074913aa45c;
    5'b11011 : xpb = 1024'h301e684f7eec31e40b3ab3a2a3835ec06c090f59464f3b24e6aa2d2d2248c635d6867744ce66c189daadfaa522cc6179bf82d2a0fe4518cf64160d458c7de30d8d458f1581f1425072c0c804c8457ae1d8a78193f8fe2889db2270c1aa1e53a8f582c04f57b6fc68da2007cc98ac38929a616e173a1f8e7d7c1a553eabdfba70;
    5'b11100 : xpb = 1024'h4c134709cfc2e639a4fb50c88610de9ab9bc1063d0d5aa70dbed9fa3cc4bddb44740da205c4a56b70d5a16c8b78c8d7fcbf3d6dc0358aa5d8b70d4c7dcc7a76ab6b2af26b3ba57542de8381d0c42af76343cab5ab837e4dd49ffa700f1ece09ef29badadca7cb8cd8dded4f534d16fba98d12ae4482be3f1949d9a08c684d084;
    5'b11101 : xpb = 1024'h680825c420999a8f3ebbedee689e5e75076f116e5b5c19bcd131121a764ef532b7fb3cfbea2debe4400632ec4c4cb985d864db17086c3bebb2cb9c4a2d116bc7e01fcf37e5836c57e90fa835503fe40a8fd1d5217771a130b8dcdd4039bb6d94efb49b0c3d427532419da21dd0f6a6e29740e7b156383965ad20ded2e129e698;
    5'b11110 : xpb = 1024'h83fd047e71704ee4d87c8b144b2bde4f55221278e5e28908c674849120520cb128b59fd77811811172b24f0fe10ce58be4d5df520d7fcd79da2663cc7d5b3025098cef49174c815ba437184d943d189eeb66fee836ab5d8427ba137f8189fa8aeccd886ab0083196f55c6f466d1bde0a95b0a47e64448ed9c5a4239cfbcefcac;
    5'b11111 : xpb = 1024'h9ff1e338c247033a723d283a2db95e29a2d513837068f854bbb7f707ca55242f997002b305f5163ea55e6b3375cd1191f146e38d12935f0801812b4ecda4f48232fa0f5a4915965f5f5e8865d83a4d3346fc28aef5e519d7969749bec9588780e9e675c922cdedfba91b3c6f094115329420614b7250e44dde276867167412c0;
    endcase
end

endmodule

module xpb_5_900
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h681887084361b02d0175eeadce80d4d1438873e35334ddecbf1b7cb0f64e209a5b0b7e023d0520bf38cb46649eb1dbc7049ec89fbb7ac721654682e9669ff258c1ab5de9bb52b1a8738bc55e7743acc7dee9212788bd726047fc040518ed55ac2a9482def3074b5deade84edcc210b74baa1e7e670ddd976c8658c2a65245470;
    5'b00010 : xpb = 1024'h1f83c8bac4d52b9137e665848ca76251159ae495d0f21b62005a400c3999942cb2ce7e8bafe3c2efd2384d825a05a6c3a52369595442bdf719edc674926d70000f078724c714660bd47d881a55ab955ec9cd48b684f4b7afda6b760f77b008c62621739435459e2e4efd22fca071f0c02669f0ea917055bd4a5b9d5041664275;
    5'b00011 : xpb = 1024'h879c4fc30836dbbe395c54325b283722592358792426f94ebf75bcbd2fe7b4c70dd9fc8dece8e3af0b0393e6f8b7828aa9c231f90fbd85187f34495df90d6258d0b2e50e826717b448094d78ccef4226a8b669de0db22a1022677a14909d5e7250b5f673284ce98c39dba7ea6c92fc34e10bd8d1024e2f3412c1297aa68a96e5;
    5'b00100 : xpb = 1024'h3f07917589aa57226fcccb09194ec4a22b35c92ba1e436c400b4801873332859659cfd175fc785dfa4709b04b40b4d874a46d2b2a8857bee33db8ce924dae0001e0f0e498e28cc17a8fb1034ab572abd939a916d09e96f5fb4d6ec1eef60118c4c42e7286a8b3c5c9dfa45f940e3e1804cd3e1d522e0ab7a94b73aa082cc84ea;
    5'b00101 : xpb = 1024'ha720187dcd0c074f7142b9b6e7cf99736ebe3d0ef51914b0bfcffcc9698148f3c0a87b199ccca69edd3be16952bd294e4ee59b526400430f99220fd28b7ad258dfba6c33497b7dc01c86d593229ad7857283b29492a6e1bffcd2f024084d673876d76a075d9287ba88d8cae70d04ecf50775c9bb93be84f15d1cc6cae7f0d95a;
    5'b00110 : xpb = 1024'h5e8b5a304e7f82b3a7b3308da5f626f340d0adc172d65226010ec024acccbc86186b7ba30fab48cf76a8e8870e10f44aef6a3c0bfcc839e54dc9535db74850002d16956e553d32237d78984f0102c01c5d67da238ede270f8f42622e67101a5272645abc9fd0da8aecf768f5e155d240733dd2bfb4510137df12d7f0c432c75f;
    5'b00111 : xpb = 1024'h15f69be2cff2fe17de23a764641cb47312e31e73f0938f9b424d837ff0183018702e7c2c8289eb001015efa4c964bf478feedcc5959030bb027096e8e315cda77a72bea960fee686de6a5b0adf6aa8b3484c01b28b156c5f21b1d438c5d2cd6c6df14b71e20f2d5b51160704b5a6b78bdf05dbc3d4e37d7e6108e916a074b564;
    5'b01000 : xpb = 1024'h7e0f22eb1354ae44df999612329d8944566b925743c86d8801690030e66650b2cb39fa2ebf8f0bbf48e1360968169b0e948da565510af7dc67b719d249b5c0003c1e1c931c51982f51f6206956ae557b273522da13d2debf69add83ddec023189885ce50d51678b93bf48bf281c7c30099a7c3aa45c156f5296e7541059909d4;
    5'b01001 : xpb = 1024'h357a649d94c829a9160a0ce8f0c416c4287e0309c185aafd42a7c38c29b1c44522fcfab8326dadefe24e3d27236a660b3512461ee9d2eeb21c5e5d5d75833da7897a45ce28134c92b2e7e32535163e1212194a69100a240efc1d4a483d82d6329412bf061754cb89a0132a015618a84c056fccae6653d33bab648666e1daf7d9;
    5'b01010 : xpb = 1024'h9d92eba5d829d9d6177ffb96bf44eb956c0676ed14ba88ea01c3403d1fffe4df7e0878ba6f72ceaf1b19838bc21c41d239b10ebea54db5d381a4e046dc2330004b25a3b7e365fe3b2673a883ac59ead9f1026b9098c7966f44194e4d56702bdebea741e50a5c16e78af1aeef2239b3c0c011b494d731acb273ca129146ff4c49;
    5'b01011 : xpb = 1024'h54fe2d58599d553a4df0726d7d6b79153e18e79f9277c65f43020398634b5871d5cb7943e25170dfb4868aa97d700cceda35af783e15aca9364c23d207f0ada79881ccf2ef27b29e87656b3f8ac1d370dbe6931f94fedbbed688c057b532def8ba34329a4c9a69b7ef104cfdf68a990c2bd9bd98f7c428f8f5c023b723413a4e;
    5'b01100 : xpb = 1024'hc696f0adb10d09e8460e9443b920695102b5852103503d48440c6f3a696cc042d8e79cd553013104df391c738c3d7cb7aba5031d6dda37eeaf3675d33be2b4ee5ddf62dfae96701e8572dfb6929bc07c6cabaae9136210e68f8326213f59212b5c1234f8ed8bc88532eeb0ccadb7e5797a1c69d1856a53f77b634dcff832853;
    5'b01101 : xpb = 1024'h7481f6131e7280cb85d6d7f20a12db6653b3cc356369e1c1435c43a49ce4ec9e8899f7cf923533cf86bed82bd775b3927f5918d192586aa05039ea469a5e1da7a7895417b63c18aa5be2f359e06d68cfa5b3dbd619f3936eb0f436672ce2e7bee055a62e81e007e63e0d6ffa96fc89cc5243ae8389347eb6401bc10764a77cc3;
    5'b01110 : xpb = 1024'h2bed37c59fe5fc2fbc474ec8c83968e625c63ce7e1271f36849b06ffe0306030e05cf8590513d600202bdf4992c97e8f1fddb98b2b20617604e12dd1c62b9b4ef4e57d52c1fdcd0dbcd4b615bed5516690980365162ad8be4363a8718ba59ad8dbe296e3c41e5ab6a22c0e096b4d6f17be0bb787a9c6fafcc211d22d40e96ac8;
    5'b01111 : xpb = 1024'h9405becde347ac5cbdbd3d7696ba3db7694eb0cb345bfd2343b683b0d67e80cb3b68765b4218f6bf58f725ae317b5a56247c822ae69b28976a27b0bb2ccb8da7b690db3c7d507eb630607b743618fe2e6f81248c9ee84b1e8b5fac76a492f085067719c2b725a6148d0a92f7376e7a8c78ad9f6e1aa4d4738a775e57a60dbf38;
    5'b10000 : xpb = 1024'h4b71008064bb27c0f42db44d54e0cb373b61217db2193a9884f5470c19c9f45d932b76e4b4f798eff2642ccbeccf2552c50122e47f631f6d1ecef44658990b4f03ed04778912331991523e301480e6c55a654c1b9b1f906e1dcf1e810355a39f02040a77f963f8e4f12931060bbf5fd7e475a8723b3750ba0c6d6f7d824fad3d;
    5'b10001 : xpb = 1024'h2dc4232e62ea3252a9e2b24130758b70d7392302fd6780dc6340a675d1567efeaee776e27d63b208bd133e9a822f04f6585c39e182b1642d37637d1846688f651492db294d3e77cf24400ebf2e8cf5c454973aa9756d5bdb03e908b621856b8fd90fb2d3ba24bb55547cf14e0104523503db1765bc9cd008e6380a35e919b42;
    5'b10010 : xpb = 1024'h6af4c93b299053522c1419d1e1882d8850fc0613830b55fa854f87185363888a45f9f57064db5bdfc49c7a4e46d4cc166a248c3dd3a5dd6438bcbabaeb067b4f12f48b9c5026992565cfc64a6a2c7c24243294d22014481df83a94907b05ac6528257e0c2ea9971340265402ac3150980adf995ccca7a67756c90ccdc3b5efb2;
    5'b10011 : xpb = 1024'h22600aedab03ceb6628490a89faebb08230e76c600c8936fc68e4a7396aefc1c9dbcf5f9d7b9fe105e09816c022897130aa92cf76c6dd439ed63fe4616d3f8f66050b4d75be84d88c6c18906489464bb0f16bc611c4b8d6d8aaa069ad9c85f7f23b26ec170e7e9e3a444f211808235e376a7a260ed3a22bdd8bf1df39ff7ddb7;
    5'b10100 : xpb = 1024'h8a7891f5ee657ee363fa7f566e2f8fd96696eaa953fd715c85a9c7248cfd1cb6f8c873fc14bf1ecf96d4c7d0a0da72da0f47f59727e89b5b52aa812f7d73eb4f21fc12c1173aff313a4d4e64bfd81182edffdd88a508ffcdd2a60a9ff2b5b52b4e46f1a063ef35418f2376ff4ca3415831498a475e17fc34a124aa1e051c3227;
    5'b10101 : xpb = 1024'h41e3d3a86fd8fa479a6af62d2c561d5938a95b5bd1baaed1c6e88a7fd0489049508b7485879dc1003041ceee5c2e3dd6afcc9650c0b092310751c4baa94168f66f583bfc22fcb3949b3f11209e3ffa19d8e40517a140451d65157caa5178684549d3e255a62d8811f342150e20f426a39d11934b7eaa787b231abb43e15e202c;
    5'b10110 : xpb = 1024'ha9fc5ab0b33aaa749be0e4dafad6f22a7c31cf3f24ef8cbe86040730c696b0e3ab96f287c4a2e1bf690d1552fae0199db46b5ef07c2b59526c9847a40fe15b4f310399e5de4f653d0ecad67f1583a6e1b7cd263f29fdb77dad1180af6a65bdf1746865349934d36fde2099fbed15321857b37b31ef8851f1eb80476e4682749c;
    5'b10111 : xpb = 1024'h61679c6334ae25d8d2515bb1b8fd7faa4e443ff1a2acca33c742ca8c09e224760359f311378183f0027a1c70b633e49a54efffaa14f35028213f8b2f3baed8f67e5fc320ea1119a06fbc993af3eb8f78a2b14dce2634fccd3f80f2b9c928710b6ff555e9db732640423f380ac1661763c37b8436101ace386d76589422c462a1;
    5'b11000 : xpb = 1024'h18d2de15b621a13d08c1d28877240d2a2056b0a4206a07a908818de74d2d98085b1cf39aaa6026209be7238e7187af96f574a063adbb46fdd5e6ceba677c569dcbbbec5bf5d2ce03d0ae5bf6d253780f8d95755d226c421cd1f064c427eb24256b82469f1db17910a65dd61995b6fcaf2f438d3a30ad4a7eef6c69b9ff0650a6;
    5'b11001 : xpb = 1024'h80eb651df983516a0a37c13645a4e1fb63df2487739ee595c79d0a98437bb8a2b628719ce76546dfd4b269f310398b5dfa13690369360e1f3b2d51a3ce1c48f68d674a45b1257fac443a2155499724d76c7e9684ab29b47d19ec68c940d879d19616c97e10b8c46e913c5b0761d80823e9e57520a18b23f5b7d1f5e4642aa516;
    5'b11010 : xpb = 1024'h3856a6d07af6ccce40a8380d03cb6f7b35f19539f15c230b08dbcdf386c72c350deb72265a43e9106e1f7110cb8d565a9a9809bd01fe04f4efd4952ef9e9c69ddac37380bce7340fa52be41127ff0d6e5762be13a760f9ccac5bdad39f9b2ceb91a3ba3352f7173ef55af9163628ed6f55ad7e24c21da03c39c8070a406c931b;
    5'b11011 : xpb = 1024'ha06f2dd8be587cfb421e26bad24c444c797a091d449100f7c7f74aa47d154ccf68f6f028974909cfa6eab7756a3f32219f36d25cbd78cc16551b18186089b8f69c6ed16a7839e5b818b7a96f9f42ba36364bdf3b301e6c2cf457ded8b8888297bc383d1245fe629ce0397e040249f8e4104f660b32fb79b3022d9334a590e78b;
    5'b11100 : xpb = 1024'h57da6f8b3fcbf85f788e9d919072d1cc4b8c79cfc24e3e6d09360dffc060c061c0b9f0b20a27ac004057be932592fd1e3fbb73165640c2ec09c25ba38c57369de9cafaa583fb9a1b79a96c2b7daaa2cd213006ca2c55b17c86c750e3174b35b1b7c52dc7883cb56d44581c12d69ade2f7c176f0f538df5f98423a45a81d2d590;
    5'b11101 : xpb = 1024'hf45b13dc13f73c3aeff14684e995f4c1d9eea82400b7be24a74d15b03ac33f4187cf13b7d064e30d9c4c5b0e0e6c81ae04013cfef08b9c1be699f2eb824b445372723e08fbd4e7eda9b2ee75c128b640c142e59288cf6cc1936c2ed760de8cbb3521e7cca7b083da876ba21aaebc37ae7df7813742072400619b5805e14c395;
    5'b11110 : xpb = 1024'h775e384604a123f0b07503161d1a341d61275e65934059cf09904e0bf9fa548e73886f3dba0b6ef012900c157f98a3e1e4dedc6faa8380e323b022181ec4a69df8d281ca4b1000274e26f445d356382beafd4f80b14a692c6132c6f28efb3e77dde6a15bbd82539b93553f0f770cceefa2815ff9e4fe4bb6ce7f41aac3391805;
    5'b11111 : xpb = 1024'h2ec979f886149f54e6e579ecdb40c19d3339cf1810fd97444acf11673d45c820cb4b6fc72cea1120abfd13333aec6ede85637d29434b77b8d85765a34a922445462eab0556d1b48aaf18b701b1be20c2d5e1770fad81ae7bf3a238fcedbdf191d9739210ffc0a66bf773dd1e4b5db43b0e4968fe0590c7fd507552d09f7b060a;
    endcase
end

endmodule

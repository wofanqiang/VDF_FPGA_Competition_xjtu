module xpb_5_990
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'ha02cd8d7de3a11c80fdabd1d9d6448f89c661e3eb8e4d14f5d52c7ce3c27a1b0409fa90ce80b505512fabbe37722c40e5c35632f70992a81e18092c4807de471f905a8b13b5b06edf7876188e6d3c7281c8d6bd2eb30a7cc96cdd487a49e74592d7a3f9d9c4ccf4143708ddedd30bb8665fa09953c7cbbf6856a582849996bc5;
    5'b00010 : xpb = 1024'h8fac6c59fa85eec754b002642a6e4a9fc756394c9c5202273cc8d646c54c96587df6d4a105f0221b869738800ae7775254509e78be7f84b81261e62ac62954327dbc1cb3c7251096dc74c06f34cbca1f4515de0d49db2288780f17148f1246202beced1187d0a5f5002134dec29150e37d1a344828ae1abcc465354c0a50711f;
    5'b00011 : xpb = 1024'h7f2bffdc16d1cbc6998547aab7784c46f246545a7fbf32ff1c3ee4bf4e718b00bb4e003523d4f3e1fa33b51c9eac2a964c6bd9c20c65deee434339910bd4c3f3027290b652ef1a3fc1621f5582c3cd166d9e5047a8859d44595059a1798617e72a5f9a8573547ca8bcd1dbdea7f1e640943a5efb14df79830360126fcb077679;
    5'b00100 : xpb = 1024'h6eab935e331da8c5de5a8cf144824dee1d366f68632c63d6fbb4f337d7967fa8f8a52bc941b9c5a86dd031b93270ddda4487150b5a4c392474248cf7518033b3872904b8deb923e8a64f7e3bd0bbd00d9626c282073018003a919c2e63f9e9ae28d247f95ed8535c798282de8d527b9dab5a89ae0110d849425aef938bbe7bd3;
    5'b00101 : xpb = 1024'h5e2b26e04f6985c5232fd237d18c4f9548268a76469994aedb2b01b060bb745135fc575d5f9e976ee16cae55c635911e3ca25054a832935aa505e05d972ba3740bdf78bb6a832d918b3cdd221eb3d304beaf34bc65da92bc1bd2debb4e6dbb752744f56d4a5c2a10363329de72b310fac27ab460ed42370f8155ccb74c75812d;
    5'b00110 : xpb = 1024'h4daaba626bb562c46805177e5e96513c7316a5842a06c586baa11028e9e068f9735382f17d83693555092af259fa446234bd8b9df618ed90d5e733c3dcd713349095ecbdf64d373a702a3c086cabd5fbe737a6f6c4850d77fd14214838e18d3c25b7a2e135e000c3f2e3d0de5813a657d99adf13d97395d5c050a9db0d2c8687;
    5'b00111 : xpb = 1024'h3d2a4de488013fc3acda5cc4eba052e39e06c0920d73f65e9a171ea173055da1b0aaae859b683afbc8a5a78eedbef7a62cd8c6e743ff47c706c8872a228282f5154c60c0821740e355179aeebaa3d8f30fc01931232f8833de5563d523555f03242a50552163d777af9477de3d743bb4f0bb09c6c5a4f49bff4b86fecde38be1;
    5'b01000 : xpb = 1024'h2ca9e166a44d1cc2f1afa20b78aa548ac8f6db9ff0e12736798d2d19fc2a5249ee01da19b94d0cc23c42242b8183aaea24f4023091e5a1fd37a9da90682df2b59a02d4c30de14a8c3a04f9d5089bdbea38488b6b81da02efbf96a6620dc930ca229cfdc90ce7ae2b6c451ede22d4d11207db3479b1d653623e4664228e9a913b;
    5'b01001 : xpb = 1024'h1c2974e8c098f9c23684e75205b45631f3e6f6add44e580e59033b92854f46f22b5905add731de88afdea0c815485e2e1d0f3d79dfcbfc33688b2df6add962761eb948c599ab54351ef258bb5693dee160d0fda5e0847daba0d7e8eef83d0291210fab3cf86b84df28f5c5de0835666f1efb5f2c9e07b2287d4141464f519695;
    5'b01010 : xpb = 1024'hba9086adce4d6c17b5a2c9892be57d91ed711bbb7bb88e638794a0b0e743b9a68b03141f516b04f237b1d64a90d1172152a78c32db25669996c815cf384d236a36fbcc825755dde03dfb7a1a48be1d889596fe03f2ef86782192b7be2b0d4581f8258b0e3ef5b92e5a66cdded95fbcc361b89df8a3910eebc3c1e6a10089bef;
    5'b01011 : xpb = 1024'habd5e142bb1ee8898b34e9b63022a0d1bb3d2ffa70a05a3595cc11d94a9bdd4aa94fda4edd2200a43675d948202fd580715fdbf29e4b80eb7aed14217402b6a89c75657960d064cbfb67192a8b5fa900a5e6dbb32a5fa03418e70003874f48b14cfc984e803c2ad42916fabccac6b7529c159374c6b5cce541a6769259a207b4;
    5'b01100 : xpb = 1024'h9b5574c4d76ac588d00a2efcbd2ca278e62d4b08540d8b0d75422051d3c0d1f2e6a705e2fb06d26aaa1255e4b3f488c4697b173bec31db21abce6787b9ae2669212bd97bec9a6e74e0547810d957abf7ce6f4ded890a1aeffa28429071c31a784b6f45c26bc00187e5c7a1bcb0274cafb335be27b2e72bab80a153b61a590d0e;
    5'b01101 : xpb = 1024'h8ad50846f3b6a28814df74434a36a420111d6616377abbe554b82eca5ce5c69b23fe317718eba4311daed28147b93c08619652853a183557dcafbaedff599629a5e24d7e7864781dc541d6f7274faeeef6f7c027e7b495abdb69851d5c36ec3f49e1f3365743d83ba27848bc9587e20cca55e8da9f188a71bf9c30d9db101268;
    5'b01110 : xpb = 1024'h7a549bc910027f8759b4b989d740a5c73c0d81241ae7ecbd342e3d42e60abb4361555d0b36d075f7914b4f1ddb7def4c59b18dce87fe8f8e0d910e54450505ea2a98c181042e81c6aa2f35dd7547b1e61f803262465f1067bcaac7aa46aabe064854a0aa42c7aeef5f28efbc7ae87769e176138d8b49e937fe970dfd9bc717c2;
    5'b01111 : xpb = 1024'h69d42f4b2c4e5c869e89fed0644aa76e66fd9c31fe551d9513a44bbb6f2fafeb9eac889f54b547be04e7cbba6f42a29051ccc917d5e4e9c43e7261ba8ab075aaaf4f35838ff88b6f8f1c94c3c33fb4dd4808a49ca5098b239dec0a37311e8fcd46c74e1e2e4b85a31bd996bc60490cc6f8963e40777b47fe3d91eb215c7e1d1c;
    5'b10000 : xpb = 1024'h5953c2cd489a3985e35f4416f154a91591edb73fe1c24e6cf31a5a33f854a493dc03b433729a198478844857030755d449e8046123cb43fa6f53b520d05be56b3405a9861bc295187409f3aa1137b7d4709116d703b405df7f2d4cc41b9261944539fb9219cf5c56d88a3dbc45a9a2240fb668f363aca6c47c8cc8451d352276;
    5'b10001 : xpb = 1024'h48d3564f64e616852834895d7e5eaabcbcddd24dc52f7f44d29068ac8179993c195adfc7907eeb4aec20c4f396cc091842033faa71b19e30a03508871607552bb8bc1d88a78c9ec158f752905f2fbacb99198911625e809b606e8f510606335b43aca9060553330a953ae4bc2b0a378126d693a64fde058abb87a568ddec27d0;
    5'b10010 : xpb = 1024'h3852e9d18131f3846d09cea40b68ac63e7cded5ba89cb01cb20677250a9e8de456b20b5bae63bd115fbd41902a90bc5c3a1e7af3bf97f866d1165bed5bb2c4ec3d72918b3356a86a3de4b176ad27bdc2c1a1fb4bc108fb5741afd1ddf07a0522421f5679f0d709be51eb8bbc106accde3df6be593c0f6450fa82828c9ea32d2a;
    5'b10011 : xpb = 1024'h27d27d539d7dd083b1df13ea9872ae0b12be08698c09e0f4917c859d93c3828c940936efcc488ed7d359be2cbe556fa03239b63d0d7e529d01f7af53a15e34acc229058dbf20b21322d2105cfb1fc0b9ea2a6d861fb3761322f1146adaedd6e9409203eddc5ae0720e9c32bbf5cb623b5516e90c2840c317397d5fb05f5a3284;
    5'b10100 : xpb = 1024'h175210d5b9c9ad82f6b45931257cafb23dae23776f7711cc70f294161ce87734d1606283ea2d609e46f63ac9521a22e42a54f1865b64acd332d902b9e709a46d46df79904aeabbbc07bf6f434917c3b112b2dfc07e5df0cf043256f7c561a8b03f04b161c7deb725cb4cd9bbdb2bf7986c3713bf147221dd78783cd4201137de;
    5'b10101 : xpb = 1024'h6d1a457d6158a823b899e77b286b159689e3e8552e442a45068a28ea60d6bdd0eb78e1808123264ba92b765e5ded62822702ccfa94b070963ba56202cb5142dcb95ed92d6b4c564ecacce29970fc6a83b3b51fadd086b8ae5739984afd57a773d775ed5b3628dd987fd80bbc08c8cf583573e7200a380a3b77319f7e0c83d38;
    5'b10110 : xpb = 1024'ha6fe7d2fb44f9c4a4b645b954feafa5205045cc40bc913f3adbb6a5ce2350d8d4f573724f01d82b9cd8d73495d019a367ea58fff19e4318b453ae8e4ad32f89fc49b9644120fcc52e4342fb27de38dd057c8bdcdc83913577c416e0c5473eed06af19e734faf5d1acb6e0e9a9dbd487be95148073d203c9a3cdd72202a61a8fd;
    5'b10111 : xpb = 1024'h967e10b1d09b79499039a0dbdcf4fbf92ff477d1ef3644cb8d3178d56b5a02358cae62b90e0254804129efe5f0c64d7a76c0cb4867ca8bc1761c3c4af2de686049520a469dd9d5fbc9218e98cbdb90c78051300826e38e135d82b0993ee7c09769644be73b3333ce881eb59a831dddd9007172ba29519b607bd84f43eb18ae57;
    5'b11000 : xpb = 1024'h85fda433ece75648d50ee62269fefda05ae492dfd2a375a36ca7874df47ef6ddca058e4d2be72646b4c66c82848b00be6edc0691b5b0e5f7a6fd8fb13889d820ce087e4929a3dfa4ae0eed7f19d393bea8d9a242858e08cf3ec3f326295b925e67d6f95b26b70a8244cf5c9a687e733617919d6d1582fa26bad32c67abcfb3b1;
    5'b11001 : xpb = 1024'h757d37b60933334819e42b68f708ff4785d4adedb610a67b4c1d95c67da3eb86075cb9e149cbf80d2862e91f184fb40266f741db0397402dd7dee3177e3547e152bef24bb56de94d92fc4c6567cb96b5d162147ce438838b200535b313cf64256649a6cf123ae1360180039a4ddf08932eb1c82001b458ecf9ce098b6c86b90b;
    5'b11010 : xpb = 1024'h64fccb38257f10475eb970af841300eeb0c4c8fb997dd7532b93a43f06c8e02e44b3e57567b0c9d39bff65bbac1467465f127d24517d9a6408c0367dc3e0b7a1d775664e4137f2f677e9ab4bb5c399acf9ea86b742e2fe470146783ffe4335ec64bc5442fdbeb7e9be30aa9a333f9df045d1f2d2ede5b7b338c8e6af2d3dbe65;
    5'b11011 : xpb = 1024'h547c5eba41caed46a38eb5f6111d0295dbb4e4097ceb082b0b09b2b78fedd4d6820b110985959b9a0f9be2583fd91a8a572db86d9f63f49a39a189e4098c27625c2bda50cd01fc9f5cd70a3203bb9ca42272f8f1a18d7902e287bacce8b707b3632f01b6e9428e9d7ae1519a18a0334d5cf21d85da17167977c3c3d2edf4c3bf;
    5'b11100 : xpb = 1024'h43fbf23c5e16ca45e863fb3c9e27043d06a4ff1760583902ea7fc1301912c97ebf623c9da37a6d6083385ef4d39dcdce4f48f3b6ed4a4ed06a82dd4a4f379722e0e24e5358cc064841c4691851b39f9b4afb6b2c0037f3bec3c8fd59d32ad97a61a1af2ad4c665513791f899fe00c8aa74124838c648753fb6bea0f6aeabc919;
    5'b11101 : xpb = 1024'h337b85be7a62a7452d3940832b3105e431951a2543c569dac9f5cfa8a237be26fcb96831c15f3f26f6d4db916762811247642f003b30a9069b6430b094e306e36598c255e4960ff126b1c7fe9faba2927383dd665ee26e7aa50a3fe6bd9eab4160145c9ec04a3c04f4429f99e3615e078b3272ebb279d405f5b97e1a6f62ce73;
    5'b11110 : xpb = 1024'h22fb194096ae8444720e85c9b83b078b5c85353327329ab2a96bde212b5cb2cf3a1093c5df4410ed6a71582dfb2734563f7f6a498917033ccc458416da8e76a3ea4f36587060199a0b9f26e4eda3a5899c0c4fa0bd8ce936864b8273a8127d085e870a12abce12b8b0f34699c8c1f364a2529d9e9eab32cc34b45b3e3019d3cd;
    5'b11111 : xpb = 1024'h127aacc2b2fa6143b6e3cb1045450932877550410a9fcb8a88e1ec99b481a7777767bf59fd28e2b3de0dd4ca8eebe79a379aa592d6fd5d72fd26d77d2039e6646f05aa5afc2a2342f08c85cb3b9ba880c494c1db1c3763f2678cc50092864ecf5cf9b7869751e96c6da3ed99ae2288c1b972c8518adc919273af3861f0d0d927;
    endcase
end

endmodule

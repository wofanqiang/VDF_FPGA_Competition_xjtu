module xpb_5_940
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h104fd12e4f486bca16effc333cd8b106ca5d6df5e78789713394282b281b90d54f3370fcade1d1622d1ed61d78f7b59a6f0e80985fa42b43b0e047cfa35dc0fed7c4cc77564493f7c76d0ac4ae156870fd56597d1cc0df5e4794dc8c06bf81dbcb2939726cfbc1da49ddbf98ba508c8dd08d1df0cd2a6af4fb0c723833b340c;
    5'b00010 : xpb = 1024'h209fa25c9e90d7942ddff86679b1620d94badbebcf0f12e267285056503721aa9e66e1f95bc3a2c45a3dac3af1ef6b34de1d0130bf48568761c08f9f46bb81fdaf8998eeac8927ef8eda15895c2ad0e1faacb2fa3981bebc8f29b9180d7f03b7965272e4d9f783b493bb7f3174a1191ba11a3be19a54d5e9f618e4706766818;
    5'b00011 : xpb = 1024'h30ef738aedd9435e44cff499b68a13145f1849e1b6969c539abc78817852b27fed9a52f609a57426875c82586ae720cf4d2b81c91eec81cb12a0d76eea1942fc874e656602cdbbe75647204e0a403952f8030c7756429e1ad6be95a4143e8593617bac5746f3458edd993eca2ef1a5a971a759d2677f40def12556a89b19c24;
    5'b00100 : xpb = 1024'h413f44b93d21af285bbff0ccf362c41b2975b7d79e1e25c4ce50a0aca06e43553ccdc3f2b7874588b47b5875e3ded669bc3a02617e90ad0ec3811f3e8d7703fb5f1331dd59124fdf1db42b12b855a1c3f55965f473037d791e5372301afe076f2ca4e5c9b3ef07692776fe62e9423237423477c334a9abd3ec31c8e0cecd030;
    5'b00101 : xpb = 1024'h518f15e78c6a1af272afed00303b7521f3d325cd85a5af3601e4c8d7c889d42a8c0134ef656916eae19a2e935cd68c042b4882f9de34d8527461670e30d4c4fa36d7fe54af56e3d6e52135d7666b0a34f2afbf718fc45cd765e84ebc21bd894af7ce1f3c20eac9437154bdfba392bec512c195b401d416c8e73e3b19028043c;
    5'b00110 : xpb = 1024'h61dee715dbb286bc899fe9336d142628be3093c36d2d38a73578f102f0a564ffdb34a5ec134ae84d0eb904b0d5ce419e9a5703923dd903962541aeddd43285f90e9ccacc059b77ceac8e409c148072a5f00618eeac853c35ad7d2b48287d0b26c2f758ae8de68b1dbb327d945de34b52e34eb3a4cefe81bde24aad513633848;
    5'b00111 : xpb = 1024'h722eb8442afaf286a08fe566a9ecd72f888e01b954b4c218690d192e18c0f5d52a6816e8c12cb9af3bd7dace4ec5f7390965842a9d7d2ed9d621f6ad779046f7e66197435be00bc673fb4b60c295db16ed5c726bc9461b93f51207d42f3c8d028e209220fae24cf805103d2d1833d7e0b3dbd1959c28ecb2dd571f8969e6c54;
    5'b01000 : xpb = 1024'h827e89727a435e50b77fe199e6c5883652eb6faf3c3c4b899ca1415940dc86aa799b87e56f0e8b1168f6b0ebc7bdacd3787404c2fd215a1d87023e7d1aee07f6be2663bab2249fbe3b68562570ab4387eab2cbe8e606faf23ca6e46035fc0ede5949cb9367de0ed24eedfcc5d284646e8468ef86695357a7d86391c19d9a060;
    5'b01001 : xpb = 1024'h92ce5aa0c98bca1ace6fddcd239e393d1d48dda523c3d4fad035698468f8177fc8cef8e21cf05c739615870940b5626de782855b5cc5856137e2864cbe4bc8f595eb3032086933b602d560ea1ec0abf8e809256602c7da50843bc0ec3cbb90ba24730505d4d9d0ac98cbbc5e8cd4f0fc54f60d77367dc29cd37003f9d14d46c;
    5'b01010 : xpb = 1024'ha31e2bcf18d435e4e55fda006076ea43e7a64b9b0b4b5e6c03c991af9113a855180269decad22dd5c3345d26b9ad1808569105f3bc69b0a4e8c2ce1c61a989f46daffca95eadc7adca426baeccd61469e55f7ee31f88b9aecbd09d78437b1295ef9c3e7841d59286e2a97bf747257d8a25832b6803a82d91ce7c76320500878;
    5'b01011 : xpb = 1024'hb36dfcfd681ca1aefc4fd6339d4f9b4ab203b990f2d2e7dd375db9dab92f392a6735dadb78b3ff37f053334432a4cda2c59f868c1c0ddbe899a315ec05074af34574c920b4f25ba591af76737aeb7cdae2b5d8603c49990d13657a044a3a9471bac577eaaed154612c873b9001760a17f6104958d0d29886c988e86a38b3c84;
    5'b01100 : xpb = 1024'hc3bdce2bb7650d79133fd266da284c517c612786da5a714e6af1e205e14ac9ffb6694bd82695d09a1d720961ab9c833d34ae07247bb2072c4a835dbba8650bf21d3995980b36ef9d591c81382900e54be00c31dd590a786b5afa569050fa164d85eeb15d1bcd163b7664fb28bbc696a5c69d67499dfd037bc4955aa26c67090;
    5'b01101 : xpb = 1024'hd40d9f5a06ad79432a2fce9a1700fd5846be957cc1e1fabf9e860a3109665ad5059cbcd4d477a1fc4a90df7f249438d7a3bc87bcdb56326ffb63a58b4bc2ccf0f4fe620f617b839520898bfcd7164dbcdd628b5a75cb57c9a28f331c57b998295117eacf88c8d815c042bac176172333972a853a6b276e70bfa1ccdaa01a49c;
    5'b01110 : xpb = 1024'he45d708855f5e50d411fcacd53d9ae5f111c0372a9698430d21a325c3181ebaa54d02dd18259735e77afb59c9d8bee7212cb08553afa5db3ac43ed5aef208defccc32e86b7c0178ce7f696c1852bb62ddab8e4d7928c3727ea240fa85e791a051c412441f5c499f00a207a5a3067afc167b7a32b3851d965baae3f12d3cd8a8;
    5'b01111 : xpb = 1024'hf4ad41b6a53e50d7580fc70090b25f65db79716890f10da205ae5a87599d7c7fa4039ece303b44c0a4ce8bba1683a40c81d988ed9a9e88f75d24352a927e4eeea487fafe0e04ab84af63a18633411e9ed80f3e54af4d168631b8ec3465389be0e76a5db462c05bca53fe39f2eab83c4f3844c11c057c445ab5bab14b0780cb4;
    5'b10000 : xpb = 1024'h104fd12e4f486bca16effc333cd8b106ca5d6df5e78789713394282b281b90d54f3370fcade1d1622d1ed61d78f7b59a6f0e80985fa42b43b0e047cfa35dc0fed7c4cc77564493f7c76d0ac4ae156870fd56597d1cc0df5e4794dc8c06bf81dbcb2939726cfbc1da49ddbf98ba508c8dd08d1df0cd2a6af4fb0c723833b340c0;
    5'b10001 : xpb = 1024'h1154ce41343cf286b85efbf670a63c17370344d54600020846cd6aadda9d49e2a426a80c78bfee784ff0c37f508730f415ff68a1e59e6df7ebee4c4c9d939d0ec541193ecba8dd3743e3db70f8f6bef80d2bbf14ee8ced542c0e2a54c72b79f987dbcd0993cb7df7ee7b9b9245f59556ad95efcfd9fd11a44abd395bb6ee74cc;
    5'b10010 : xpb = 1024'h1259cb541931794359cdfbb9a473c727a3a91bb4a4787a9f5a06ad308d1f02eff919df1c439e0b8e72c2b0e12816ac4dbcf050ab6b98b0ac26fc50c997c9791eb2bd6606410d2676c05aac1d43d8157f1d0124acc058fb4a1087781d87977217448e60a0ba9b3a159319778bd19a9e1f8a9ec1aee6cfb8539a6e007f3a29a8d8;
    5'b10011 : xpb = 1024'h135ec866fe25fffffb3cfb7cd8415238104ef29402f0f3366d3fefb33fa0bbfd4e0d162c0e7c28a495949e42ffa627a763e138b4f192f360620a554691ff552ea039b2cdb6716fb63cd17cc98eb96c062cd68a449225093ff500c5e648036a350140f437e16af63337b753855d3fa6e867a7938df3a25f02ea1ec7a2bd64dce4;
    5'b10100 : xpb = 1024'h1463c579e31a86bc9cabfb400c0edd487cf4c97361696bcd80793235f222750aa3004d3bd95a45bab8668ba4d735a3010ad220be778d36149d1859c38c35313e8db5ff952bd5b8f5b9484d75d99ac28d3cabefdc63f11735d97a13af086f6252bdf387cf083ab250dc552f7ee8e4afb144b0656d007505b239cf8ec640a010f0;
    5'b10101 : xpb = 1024'h1568c28cc80f0d793e1afb033fdc6858e99aa052bfe1e46493b274b8a4a42e17f7f3844ba43862d0db387906aec51e5ab1c308c7fd8778c8d8265e40866b0d4e7b324c5ca13a023535bf1e22247c19144c81557435bd252bbdf36177c8db5a707aa61b662f0a6e6e80f30b787489b87a21b9374c0d47ac61898055e9c3db44fc;
    5'b10110 : xpb = 1024'h166dbf9fad039435df89fac673a9f369564077321e5a5cfba6ebb73b5725e7254ce6bb5b6f167fe6fe0a6668865499b458b3f0d18381bb7d133462bd80a0e95e68ae9924169e4b74b235eece6f5d6f9b5c56bb0c07893321a26caf408947528e3758aefd55da2a8c2590e772002ec142fec2092b1a1a5310d9311d0d47167908;
    5'b10111 : xpb = 1024'h1772bcb291f81af280f8fa89a7777e79c2e64e117cd2d592ba24f9be09a7a032a1d9f26b39f49cfd20dc53ca5de4150dffa4d8db097bfe314e42673a7ad6c56e562ae5eb8c0294b42eacbf7aba3ec6226c2c20a3d955411786e5fd0949b34aabf40b42947ca9e6a9ca2ec36b8bd3ca0bdbcadb0a26ecf9c028e1e430ca51ad14;
    5'b11000 : xpb = 1024'h1877b9c576eca1af2267fa4cdb45098a2f8c24f0db4b4e29cd5e3c40bc29593ff6cd297b04d2ba1343ae412c35739067a695c0e48f7640e589506bb7750ca17e43a732b30166ddf3ab23902705201ca97c01863bab214f0d6b5f4ad20a1f42c9b0bdd62ba379a2c76ecc9f651778d2d4b8d3ace933bfa06f7892ab544d8ce120;
    5'b11001 : xpb = 1024'h197cb6d85be1286bc3d6fa100f12949a9c31fbd039c3c6c0e0977ec36eab124d4bc0608acfb0d72966802e8e0d030bc14d86a8ee15708399c45e70346f427d8e31237f7a76cb2733279a60d3500173308bd6ebd37ced5d034fd8989aca8b3ae76d7069c2ca495ee5136a7b5ea31ddb9d95dc7ec84092471ec8437277d0c8152c;
    5'b11010 : xpb = 1024'h1a81b3eb40d5af286545f9d342e01fab08d7d2af983c3f57f3d0c146212ccb5aa0b3979a9a8ef43f89521befe492871af47790f79b6ac64dff6c74b16978599e1e9fcc41ec2f7072a411317f9ae2c9b79bac516b4eb96af93451e6638af733052a22fd59f1191b02b80857582ec2e46672e550a74d64edce17f4399b54034938;
    5'b11011 : xpb = 1024'h1b86b0fe25ca35e506b4f99676adaabb757da98ef6b4b7ef070a03c8d3ae8467f5a6ceaa656d1155ac240951bc2202749b687901216509023a7a792e63ae35ae0c1c19096193b9b22088022be5c4203eab81b703208578ef18cb342c4b632b22e6d590f117e8d7205ca63351ba67ed2f4fee22865a37947d67a500bed73e7d44;
    5'b11100 : xpb = 1024'h1c8bae110abebca1a823f959aa7b35cbe223806e552d30861a43464b86303d754a9a05ba304b2e6bcef5f6b393b17dce4259610aa75f4bb675887dab5de411bdf99865d0d6f802f19cfed2d830a576c5bb571c9af25186e4fd4481f50bcf2340a38824883eb8933e01440f4b460cf5f82cf6f465670a3b2cb755c7e25a79b150;
    5'b11101 : xpb = 1024'h1d90ab23efb3435e4992f91cde48c0dc4ec9574db3a5a91d2d7c88ce38b1f6829f8d3cc9fb294b81f1c7e4156b40f927e94a49142d598e6ab09682285819edcde714b2984c5c4c311975a3847b86cd4ccb2c8232c41d94dae1bdcfbdcc3b1b5e603ab81f65884f5ba5e1eb44d1b1fec109ffc64473dce1dc07068f05ddb4e55c;
    5'b11110 : xpb = 1024'h1e95a836d4a7ca1aeb01f8e012164becbb6f2e2d121e21b440b5cb50eb33af8ff48073d9c60768981499d17742d07481903b311db353d11eeba486a5524fc9ddd490ff5fc1c0957095ec7430c66823d3db01e7ca95e9a2d0c6371d868ca7137c1ced4bb68c580b794a7fc73e5d570789e708982380af888b56b7562960f01968;
    5'b11111 : xpb = 1024'h1f9aa549b99c50d78c70f8a345e3d6fd2815050c70969a4b53ef0dd39db5689d4973aae990e585ae376bbed91a5fefdb372c1927394e13d326b28b224c85a5edc20d4c273724deb0126344dd11497a5aead74d6267b5b0c6aab06b4f4d130b99d99fdf4db327c796ef1da337e8fc1052c4116a028d822f3aa6681d4ce42b4d74;
    endcase
end

endmodule

module compressor_array_16_12_1033
(
    input  [15:0] col_in_0,
    input  [15:0] col_in_1,
    input  [15:0] col_in_2,
    input  [15:0] col_in_3,
    input  [15:0] col_in_4,
    input  [15:0] col_in_5,
    input  [15:0] col_in_6,
    input  [15:0] col_in_7,
    input  [15:0] col_in_8,
    input  [15:0] col_in_9,
    input  [15:0] col_in_10,
    input  [15:0] col_in_11,
    input  [15:0] col_in_12,
    input  [15:0] col_in_13,
    input  [15:0] col_in_14,
    input  [15:0] col_in_15,
    input  [15:0] col_in_16,
    input  [15:0] col_in_17,
    input  [15:0] col_in_18,
    input  [15:0] col_in_19,
    input  [15:0] col_in_20,
    input  [15:0] col_in_21,
    input  [15:0] col_in_22,
    input  [15:0] col_in_23,
    input  [15:0] col_in_24,
    input  [15:0] col_in_25,
    input  [15:0] col_in_26,
    input  [15:0] col_in_27,
    input  [15:0] col_in_28,
    input  [15:0] col_in_29,
    input  [15:0] col_in_30,
    input  [15:0] col_in_31,
    input  [15:0] col_in_32,
    input  [15:0] col_in_33,
    input  [15:0] col_in_34,
    input  [15:0] col_in_35,
    input  [15:0] col_in_36,
    input  [15:0] col_in_37,
    input  [15:0] col_in_38,
    input  [15:0] col_in_39,
    input  [15:0] col_in_40,
    input  [15:0] col_in_41,
    input  [15:0] col_in_42,
    input  [15:0] col_in_43,
    input  [15:0] col_in_44,
    input  [15:0] col_in_45,
    input  [15:0] col_in_46,
    input  [15:0] col_in_47,
    input  [15:0] col_in_48,
    input  [15:0] col_in_49,
    input  [15:0] col_in_50,
    input  [15:0] col_in_51,
    input  [15:0] col_in_52,
    input  [15:0] col_in_53,
    input  [15:0] col_in_54,
    input  [15:0] col_in_55,
    input  [15:0] col_in_56,
    input  [15:0] col_in_57,
    input  [15:0] col_in_58,
    input  [15:0] col_in_59,
    input  [15:0] col_in_60,
    input  [15:0] col_in_61,
    input  [15:0] col_in_62,
    input  [15:0] col_in_63,
    input  [15:0] col_in_64,
    input  [15:0] col_in_65,
    input  [15:0] col_in_66,
    input  [15:0] col_in_67,
    input  [15:0] col_in_68,
    input  [15:0] col_in_69,
    input  [15:0] col_in_70,
    input  [15:0] col_in_71,
    input  [15:0] col_in_72,
    input  [15:0] col_in_73,
    input  [15:0] col_in_74,
    input  [15:0] col_in_75,
    input  [15:0] col_in_76,
    input  [15:0] col_in_77,
    input  [15:0] col_in_78,
    input  [15:0] col_in_79,
    input  [15:0] col_in_80,
    input  [15:0] col_in_81,
    input  [15:0] col_in_82,
    input  [15:0] col_in_83,
    input  [15:0] col_in_84,
    input  [15:0] col_in_85,
    input  [15:0] col_in_86,
    input  [15:0] col_in_87,
    input  [15:0] col_in_88,
    input  [15:0] col_in_89,
    input  [15:0] col_in_90,
    input  [15:0] col_in_91,
    input  [15:0] col_in_92,
    input  [15:0] col_in_93,
    input  [15:0] col_in_94,
    input  [15:0] col_in_95,
    input  [15:0] col_in_96,
    input  [15:0] col_in_97,
    input  [15:0] col_in_98,
    input  [15:0] col_in_99,
    input  [15:0] col_in_100,
    input  [15:0] col_in_101,
    input  [15:0] col_in_102,
    input  [15:0] col_in_103,
    input  [15:0] col_in_104,
    input  [15:0] col_in_105,
    input  [15:0] col_in_106,
    input  [15:0] col_in_107,
    input  [15:0] col_in_108,
    input  [15:0] col_in_109,
    input  [15:0] col_in_110,
    input  [15:0] col_in_111,
    input  [15:0] col_in_112,
    input  [15:0] col_in_113,
    input  [15:0] col_in_114,
    input  [15:0] col_in_115,
    input  [15:0] col_in_116,
    input  [15:0] col_in_117,
    input  [15:0] col_in_118,
    input  [15:0] col_in_119,
    input  [15:0] col_in_120,
    input  [15:0] col_in_121,
    input  [15:0] col_in_122,
    input  [15:0] col_in_123,
    input  [15:0] col_in_124,
    input  [15:0] col_in_125,
    input  [15:0] col_in_126,
    input  [15:0] col_in_127,
    input  [15:0] col_in_128,
    input  [15:0] col_in_129,
    input  [15:0] col_in_130,
    input  [15:0] col_in_131,
    input  [15:0] col_in_132,
    input  [15:0] col_in_133,
    input  [15:0] col_in_134,
    input  [15:0] col_in_135,
    input  [15:0] col_in_136,
    input  [15:0] col_in_137,
    input  [15:0] col_in_138,
    input  [15:0] col_in_139,
    input  [15:0] col_in_140,
    input  [15:0] col_in_141,
    input  [15:0] col_in_142,
    input  [15:0] col_in_143,
    input  [15:0] col_in_144,
    input  [15:0] col_in_145,
    input  [15:0] col_in_146,
    input  [15:0] col_in_147,
    input  [15:0] col_in_148,
    input  [15:0] col_in_149,
    input  [15:0] col_in_150,
    input  [15:0] col_in_151,
    input  [15:0] col_in_152,
    input  [15:0] col_in_153,
    input  [15:0] col_in_154,
    input  [15:0] col_in_155,
    input  [15:0] col_in_156,
    input  [15:0] col_in_157,
    input  [15:0] col_in_158,
    input  [15:0] col_in_159,
    input  [15:0] col_in_160,
    input  [15:0] col_in_161,
    input  [15:0] col_in_162,
    input  [15:0] col_in_163,
    input  [15:0] col_in_164,
    input  [15:0] col_in_165,
    input  [15:0] col_in_166,
    input  [15:0] col_in_167,
    input  [15:0] col_in_168,
    input  [15:0] col_in_169,
    input  [15:0] col_in_170,
    input  [15:0] col_in_171,
    input  [15:0] col_in_172,
    input  [15:0] col_in_173,
    input  [15:0] col_in_174,
    input  [15:0] col_in_175,
    input  [15:0] col_in_176,
    input  [15:0] col_in_177,
    input  [15:0] col_in_178,
    input  [15:0] col_in_179,
    input  [15:0] col_in_180,
    input  [15:0] col_in_181,
    input  [15:0] col_in_182,
    input  [15:0] col_in_183,
    input  [15:0] col_in_184,
    input  [15:0] col_in_185,
    input  [15:0] col_in_186,
    input  [15:0] col_in_187,
    input  [15:0] col_in_188,
    input  [15:0] col_in_189,
    input  [15:0] col_in_190,
    input  [15:0] col_in_191,
    input  [15:0] col_in_192,
    input  [15:0] col_in_193,
    input  [15:0] col_in_194,
    input  [15:0] col_in_195,
    input  [15:0] col_in_196,
    input  [15:0] col_in_197,
    input  [15:0] col_in_198,
    input  [15:0] col_in_199,
    input  [15:0] col_in_200,
    input  [15:0] col_in_201,
    input  [15:0] col_in_202,
    input  [15:0] col_in_203,
    input  [15:0] col_in_204,
    input  [15:0] col_in_205,
    input  [15:0] col_in_206,
    input  [15:0] col_in_207,
    input  [15:0] col_in_208,
    input  [15:0] col_in_209,
    input  [15:0] col_in_210,
    input  [15:0] col_in_211,
    input  [15:0] col_in_212,
    input  [15:0] col_in_213,
    input  [15:0] col_in_214,
    input  [15:0] col_in_215,
    input  [15:0] col_in_216,
    input  [15:0] col_in_217,
    input  [15:0] col_in_218,
    input  [15:0] col_in_219,
    input  [15:0] col_in_220,
    input  [15:0] col_in_221,
    input  [15:0] col_in_222,
    input  [15:0] col_in_223,
    input  [15:0] col_in_224,
    input  [15:0] col_in_225,
    input  [15:0] col_in_226,
    input  [15:0] col_in_227,
    input  [15:0] col_in_228,
    input  [15:0] col_in_229,
    input  [15:0] col_in_230,
    input  [15:0] col_in_231,
    input  [15:0] col_in_232,
    input  [15:0] col_in_233,
    input  [15:0] col_in_234,
    input  [15:0] col_in_235,
    input  [15:0] col_in_236,
    input  [15:0] col_in_237,
    input  [15:0] col_in_238,
    input  [15:0] col_in_239,
    input  [15:0] col_in_240,
    input  [15:0] col_in_241,
    input  [15:0] col_in_242,
    input  [15:0] col_in_243,
    input  [15:0] col_in_244,
    input  [15:0] col_in_245,
    input  [15:0] col_in_246,
    input  [15:0] col_in_247,
    input  [15:0] col_in_248,
    input  [15:0] col_in_249,
    input  [15:0] col_in_250,
    input  [15:0] col_in_251,
    input  [15:0] col_in_252,
    input  [15:0] col_in_253,
    input  [15:0] col_in_254,
    input  [15:0] col_in_255,
    input  [15:0] col_in_256,
    input  [15:0] col_in_257,
    input  [15:0] col_in_258,
    input  [15:0] col_in_259,
    input  [15:0] col_in_260,
    input  [15:0] col_in_261,
    input  [15:0] col_in_262,
    input  [15:0] col_in_263,
    input  [15:0] col_in_264,
    input  [15:0] col_in_265,
    input  [15:0] col_in_266,
    input  [15:0] col_in_267,
    input  [15:0] col_in_268,
    input  [15:0] col_in_269,
    input  [15:0] col_in_270,
    input  [15:0] col_in_271,
    input  [15:0] col_in_272,
    input  [15:0] col_in_273,
    input  [15:0] col_in_274,
    input  [15:0] col_in_275,
    input  [15:0] col_in_276,
    input  [15:0] col_in_277,
    input  [15:0] col_in_278,
    input  [15:0] col_in_279,
    input  [15:0] col_in_280,
    input  [15:0] col_in_281,
    input  [15:0] col_in_282,
    input  [15:0] col_in_283,
    input  [15:0] col_in_284,
    input  [15:0] col_in_285,
    input  [15:0] col_in_286,
    input  [15:0] col_in_287,
    input  [15:0] col_in_288,
    input  [15:0] col_in_289,
    input  [15:0] col_in_290,
    input  [15:0] col_in_291,
    input  [15:0] col_in_292,
    input  [15:0] col_in_293,
    input  [15:0] col_in_294,
    input  [15:0] col_in_295,
    input  [15:0] col_in_296,
    input  [15:0] col_in_297,
    input  [15:0] col_in_298,
    input  [15:0] col_in_299,
    input  [15:0] col_in_300,
    input  [15:0] col_in_301,
    input  [15:0] col_in_302,
    input  [15:0] col_in_303,
    input  [15:0] col_in_304,
    input  [15:0] col_in_305,
    input  [15:0] col_in_306,
    input  [15:0] col_in_307,
    input  [15:0] col_in_308,
    input  [15:0] col_in_309,
    input  [15:0] col_in_310,
    input  [15:0] col_in_311,
    input  [15:0] col_in_312,
    input  [15:0] col_in_313,
    input  [15:0] col_in_314,
    input  [15:0] col_in_315,
    input  [15:0] col_in_316,
    input  [15:0] col_in_317,
    input  [15:0] col_in_318,
    input  [15:0] col_in_319,
    input  [15:0] col_in_320,
    input  [15:0] col_in_321,
    input  [15:0] col_in_322,
    input  [15:0] col_in_323,
    input  [15:0] col_in_324,
    input  [15:0] col_in_325,
    input  [15:0] col_in_326,
    input  [15:0] col_in_327,
    input  [15:0] col_in_328,
    input  [15:0] col_in_329,
    input  [15:0] col_in_330,
    input  [15:0] col_in_331,
    input  [15:0] col_in_332,
    input  [15:0] col_in_333,
    input  [15:0] col_in_334,
    input  [15:0] col_in_335,
    input  [15:0] col_in_336,
    input  [15:0] col_in_337,
    input  [15:0] col_in_338,
    input  [15:0] col_in_339,
    input  [15:0] col_in_340,
    input  [15:0] col_in_341,
    input  [15:0] col_in_342,
    input  [15:0] col_in_343,
    input  [15:0] col_in_344,
    input  [15:0] col_in_345,
    input  [15:0] col_in_346,
    input  [15:0] col_in_347,
    input  [15:0] col_in_348,
    input  [15:0] col_in_349,
    input  [15:0] col_in_350,
    input  [15:0] col_in_351,
    input  [15:0] col_in_352,
    input  [15:0] col_in_353,
    input  [15:0] col_in_354,
    input  [15:0] col_in_355,
    input  [15:0] col_in_356,
    input  [15:0] col_in_357,
    input  [15:0] col_in_358,
    input  [15:0] col_in_359,
    input  [15:0] col_in_360,
    input  [15:0] col_in_361,
    input  [15:0] col_in_362,
    input  [15:0] col_in_363,
    input  [15:0] col_in_364,
    input  [15:0] col_in_365,
    input  [15:0] col_in_366,
    input  [15:0] col_in_367,
    input  [15:0] col_in_368,
    input  [15:0] col_in_369,
    input  [15:0] col_in_370,
    input  [15:0] col_in_371,
    input  [15:0] col_in_372,
    input  [15:0] col_in_373,
    input  [15:0] col_in_374,
    input  [15:0] col_in_375,
    input  [15:0] col_in_376,
    input  [15:0] col_in_377,
    input  [15:0] col_in_378,
    input  [15:0] col_in_379,
    input  [15:0] col_in_380,
    input  [15:0] col_in_381,
    input  [15:0] col_in_382,
    input  [15:0] col_in_383,
    input  [15:0] col_in_384,
    input  [15:0] col_in_385,
    input  [15:0] col_in_386,
    input  [15:0] col_in_387,
    input  [15:0] col_in_388,
    input  [15:0] col_in_389,
    input  [15:0] col_in_390,
    input  [15:0] col_in_391,
    input  [15:0] col_in_392,
    input  [15:0] col_in_393,
    input  [15:0] col_in_394,
    input  [15:0] col_in_395,
    input  [15:0] col_in_396,
    input  [15:0] col_in_397,
    input  [15:0] col_in_398,
    input  [15:0] col_in_399,
    input  [15:0] col_in_400,
    input  [15:0] col_in_401,
    input  [15:0] col_in_402,
    input  [15:0] col_in_403,
    input  [15:0] col_in_404,
    input  [15:0] col_in_405,
    input  [15:0] col_in_406,
    input  [15:0] col_in_407,
    input  [15:0] col_in_408,
    input  [15:0] col_in_409,
    input  [15:0] col_in_410,
    input  [15:0] col_in_411,
    input  [15:0] col_in_412,
    input  [15:0] col_in_413,
    input  [15:0] col_in_414,
    input  [15:0] col_in_415,
    input  [15:0] col_in_416,
    input  [15:0] col_in_417,
    input  [15:0] col_in_418,
    input  [15:0] col_in_419,
    input  [15:0] col_in_420,
    input  [15:0] col_in_421,
    input  [15:0] col_in_422,
    input  [15:0] col_in_423,
    input  [15:0] col_in_424,
    input  [15:0] col_in_425,
    input  [15:0] col_in_426,
    input  [15:0] col_in_427,
    input  [15:0] col_in_428,
    input  [15:0] col_in_429,
    input  [15:0] col_in_430,
    input  [15:0] col_in_431,
    input  [15:0] col_in_432,
    input  [15:0] col_in_433,
    input  [15:0] col_in_434,
    input  [15:0] col_in_435,
    input  [15:0] col_in_436,
    input  [15:0] col_in_437,
    input  [15:0] col_in_438,
    input  [15:0] col_in_439,
    input  [15:0] col_in_440,
    input  [15:0] col_in_441,
    input  [15:0] col_in_442,
    input  [15:0] col_in_443,
    input  [15:0] col_in_444,
    input  [15:0] col_in_445,
    input  [15:0] col_in_446,
    input  [15:0] col_in_447,
    input  [15:0] col_in_448,
    input  [15:0] col_in_449,
    input  [15:0] col_in_450,
    input  [15:0] col_in_451,
    input  [15:0] col_in_452,
    input  [15:0] col_in_453,
    input  [15:0] col_in_454,
    input  [15:0] col_in_455,
    input  [15:0] col_in_456,
    input  [15:0] col_in_457,
    input  [15:0] col_in_458,
    input  [15:0] col_in_459,
    input  [15:0] col_in_460,
    input  [15:0] col_in_461,
    input  [15:0] col_in_462,
    input  [15:0] col_in_463,
    input  [15:0] col_in_464,
    input  [15:0] col_in_465,
    input  [15:0] col_in_466,
    input  [15:0] col_in_467,
    input  [15:0] col_in_468,
    input  [15:0] col_in_469,
    input  [15:0] col_in_470,
    input  [15:0] col_in_471,
    input  [15:0] col_in_472,
    input  [15:0] col_in_473,
    input  [15:0] col_in_474,
    input  [15:0] col_in_475,
    input  [15:0] col_in_476,
    input  [15:0] col_in_477,
    input  [15:0] col_in_478,
    input  [15:0] col_in_479,
    input  [15:0] col_in_480,
    input  [15:0] col_in_481,
    input  [15:0] col_in_482,
    input  [15:0] col_in_483,
    input  [15:0] col_in_484,
    input  [15:0] col_in_485,
    input  [15:0] col_in_486,
    input  [15:0] col_in_487,
    input  [15:0] col_in_488,
    input  [15:0] col_in_489,
    input  [15:0] col_in_490,
    input  [15:0] col_in_491,
    input  [15:0] col_in_492,
    input  [15:0] col_in_493,
    input  [15:0] col_in_494,
    input  [15:0] col_in_495,
    input  [15:0] col_in_496,
    input  [15:0] col_in_497,
    input  [15:0] col_in_498,
    input  [15:0] col_in_499,
    input  [15:0] col_in_500,
    input  [15:0] col_in_501,
    input  [15:0] col_in_502,
    input  [15:0] col_in_503,
    input  [15:0] col_in_504,
    input  [15:0] col_in_505,
    input  [15:0] col_in_506,
    input  [15:0] col_in_507,
    input  [15:0] col_in_508,
    input  [15:0] col_in_509,
    input  [15:0] col_in_510,
    input  [15:0] col_in_511,
    input  [15:0] col_in_512,
    input  [15:0] col_in_513,
    input  [15:0] col_in_514,
    input  [15:0] col_in_515,
    input  [15:0] col_in_516,
    input  [15:0] col_in_517,
    input  [15:0] col_in_518,
    input  [15:0] col_in_519,
    input  [15:0] col_in_520,
    input  [15:0] col_in_521,
    input  [15:0] col_in_522,
    input  [15:0] col_in_523,
    input  [15:0] col_in_524,
    input  [15:0] col_in_525,
    input  [15:0] col_in_526,
    input  [15:0] col_in_527,
    input  [15:0] col_in_528,
    input  [15:0] col_in_529,
    input  [15:0] col_in_530,
    input  [15:0] col_in_531,
    input  [15:0] col_in_532,
    input  [15:0] col_in_533,
    input  [15:0] col_in_534,
    input  [15:0] col_in_535,
    input  [15:0] col_in_536,
    input  [15:0] col_in_537,
    input  [15:0] col_in_538,
    input  [15:0] col_in_539,
    input  [15:0] col_in_540,
    input  [15:0] col_in_541,
    input  [15:0] col_in_542,
    input  [15:0] col_in_543,
    input  [15:0] col_in_544,
    input  [15:0] col_in_545,
    input  [15:0] col_in_546,
    input  [15:0] col_in_547,
    input  [15:0] col_in_548,
    input  [15:0] col_in_549,
    input  [15:0] col_in_550,
    input  [15:0] col_in_551,
    input  [15:0] col_in_552,
    input  [15:0] col_in_553,
    input  [15:0] col_in_554,
    input  [15:0] col_in_555,
    input  [15:0] col_in_556,
    input  [15:0] col_in_557,
    input  [15:0] col_in_558,
    input  [15:0] col_in_559,
    input  [15:0] col_in_560,
    input  [15:0] col_in_561,
    input  [15:0] col_in_562,
    input  [15:0] col_in_563,
    input  [15:0] col_in_564,
    input  [15:0] col_in_565,
    input  [15:0] col_in_566,
    input  [15:0] col_in_567,
    input  [15:0] col_in_568,
    input  [15:0] col_in_569,
    input  [15:0] col_in_570,
    input  [15:0] col_in_571,
    input  [15:0] col_in_572,
    input  [15:0] col_in_573,
    input  [15:0] col_in_574,
    input  [15:0] col_in_575,
    input  [15:0] col_in_576,
    input  [15:0] col_in_577,
    input  [15:0] col_in_578,
    input  [15:0] col_in_579,
    input  [15:0] col_in_580,
    input  [15:0] col_in_581,
    input  [15:0] col_in_582,
    input  [15:0] col_in_583,
    input  [15:0] col_in_584,
    input  [15:0] col_in_585,
    input  [15:0] col_in_586,
    input  [15:0] col_in_587,
    input  [15:0] col_in_588,
    input  [15:0] col_in_589,
    input  [15:0] col_in_590,
    input  [15:0] col_in_591,
    input  [15:0] col_in_592,
    input  [15:0] col_in_593,
    input  [15:0] col_in_594,
    input  [15:0] col_in_595,
    input  [15:0] col_in_596,
    input  [15:0] col_in_597,
    input  [15:0] col_in_598,
    input  [15:0] col_in_599,
    input  [15:0] col_in_600,
    input  [15:0] col_in_601,
    input  [15:0] col_in_602,
    input  [15:0] col_in_603,
    input  [15:0] col_in_604,
    input  [15:0] col_in_605,
    input  [15:0] col_in_606,
    input  [15:0] col_in_607,
    input  [15:0] col_in_608,
    input  [15:0] col_in_609,
    input  [15:0] col_in_610,
    input  [15:0] col_in_611,
    input  [15:0] col_in_612,
    input  [15:0] col_in_613,
    input  [15:0] col_in_614,
    input  [15:0] col_in_615,
    input  [15:0] col_in_616,
    input  [15:0] col_in_617,
    input  [15:0] col_in_618,
    input  [15:0] col_in_619,
    input  [15:0] col_in_620,
    input  [15:0] col_in_621,
    input  [15:0] col_in_622,
    input  [15:0] col_in_623,
    input  [15:0] col_in_624,
    input  [15:0] col_in_625,
    input  [15:0] col_in_626,
    input  [15:0] col_in_627,
    input  [15:0] col_in_628,
    input  [15:0] col_in_629,
    input  [15:0] col_in_630,
    input  [15:0] col_in_631,
    input  [15:0] col_in_632,
    input  [15:0] col_in_633,
    input  [15:0] col_in_634,
    input  [15:0] col_in_635,
    input  [15:0] col_in_636,
    input  [15:0] col_in_637,
    input  [15:0] col_in_638,
    input  [15:0] col_in_639,
    input  [15:0] col_in_640,
    input  [15:0] col_in_641,
    input  [15:0] col_in_642,
    input  [15:0] col_in_643,
    input  [15:0] col_in_644,
    input  [15:0] col_in_645,
    input  [15:0] col_in_646,
    input  [15:0] col_in_647,
    input  [15:0] col_in_648,
    input  [15:0] col_in_649,
    input  [15:0] col_in_650,
    input  [15:0] col_in_651,
    input  [15:0] col_in_652,
    input  [15:0] col_in_653,
    input  [15:0] col_in_654,
    input  [15:0] col_in_655,
    input  [15:0] col_in_656,
    input  [15:0] col_in_657,
    input  [15:0] col_in_658,
    input  [15:0] col_in_659,
    input  [15:0] col_in_660,
    input  [15:0] col_in_661,
    input  [15:0] col_in_662,
    input  [15:0] col_in_663,
    input  [15:0] col_in_664,
    input  [15:0] col_in_665,
    input  [15:0] col_in_666,
    input  [15:0] col_in_667,
    input  [15:0] col_in_668,
    input  [15:0] col_in_669,
    input  [15:0] col_in_670,
    input  [15:0] col_in_671,
    input  [15:0] col_in_672,
    input  [15:0] col_in_673,
    input  [15:0] col_in_674,
    input  [15:0] col_in_675,
    input  [15:0] col_in_676,
    input  [15:0] col_in_677,
    input  [15:0] col_in_678,
    input  [15:0] col_in_679,
    input  [15:0] col_in_680,
    input  [15:0] col_in_681,
    input  [15:0] col_in_682,
    input  [15:0] col_in_683,
    input  [15:0] col_in_684,
    input  [15:0] col_in_685,
    input  [15:0] col_in_686,
    input  [15:0] col_in_687,
    input  [15:0] col_in_688,
    input  [15:0] col_in_689,
    input  [15:0] col_in_690,
    input  [15:0] col_in_691,
    input  [15:0] col_in_692,
    input  [15:0] col_in_693,
    input  [15:0] col_in_694,
    input  [15:0] col_in_695,
    input  [15:0] col_in_696,
    input  [15:0] col_in_697,
    input  [15:0] col_in_698,
    input  [15:0] col_in_699,
    input  [15:0] col_in_700,
    input  [15:0] col_in_701,
    input  [15:0] col_in_702,
    input  [15:0] col_in_703,
    input  [15:0] col_in_704,
    input  [15:0] col_in_705,
    input  [15:0] col_in_706,
    input  [15:0] col_in_707,
    input  [15:0] col_in_708,
    input  [15:0] col_in_709,
    input  [15:0] col_in_710,
    input  [15:0] col_in_711,
    input  [15:0] col_in_712,
    input  [15:0] col_in_713,
    input  [15:0] col_in_714,
    input  [15:0] col_in_715,
    input  [15:0] col_in_716,
    input  [15:0] col_in_717,
    input  [15:0] col_in_718,
    input  [15:0] col_in_719,
    input  [15:0] col_in_720,
    input  [15:0] col_in_721,
    input  [15:0] col_in_722,
    input  [15:0] col_in_723,
    input  [15:0] col_in_724,
    input  [15:0] col_in_725,
    input  [15:0] col_in_726,
    input  [15:0] col_in_727,
    input  [15:0] col_in_728,
    input  [15:0] col_in_729,
    input  [15:0] col_in_730,
    input  [15:0] col_in_731,
    input  [15:0] col_in_732,
    input  [15:0] col_in_733,
    input  [15:0] col_in_734,
    input  [15:0] col_in_735,
    input  [15:0] col_in_736,
    input  [15:0] col_in_737,
    input  [15:0] col_in_738,
    input  [15:0] col_in_739,
    input  [15:0] col_in_740,
    input  [15:0] col_in_741,
    input  [15:0] col_in_742,
    input  [15:0] col_in_743,
    input  [15:0] col_in_744,
    input  [15:0] col_in_745,
    input  [15:0] col_in_746,
    input  [15:0] col_in_747,
    input  [15:0] col_in_748,
    input  [15:0] col_in_749,
    input  [15:0] col_in_750,
    input  [15:0] col_in_751,
    input  [15:0] col_in_752,
    input  [15:0] col_in_753,
    input  [15:0] col_in_754,
    input  [15:0] col_in_755,
    input  [15:0] col_in_756,
    input  [15:0] col_in_757,
    input  [15:0] col_in_758,
    input  [15:0] col_in_759,
    input  [15:0] col_in_760,
    input  [15:0] col_in_761,
    input  [15:0] col_in_762,
    input  [15:0] col_in_763,
    input  [15:0] col_in_764,
    input  [15:0] col_in_765,
    input  [15:0] col_in_766,
    input  [15:0] col_in_767,
    input  [15:0] col_in_768,
    input  [15:0] col_in_769,
    input  [15:0] col_in_770,
    input  [15:0] col_in_771,
    input  [15:0] col_in_772,
    input  [15:0] col_in_773,
    input  [15:0] col_in_774,
    input  [15:0] col_in_775,
    input  [15:0] col_in_776,
    input  [15:0] col_in_777,
    input  [15:0] col_in_778,
    input  [15:0] col_in_779,
    input  [15:0] col_in_780,
    input  [15:0] col_in_781,
    input  [15:0] col_in_782,
    input  [15:0] col_in_783,
    input  [15:0] col_in_784,
    input  [15:0] col_in_785,
    input  [15:0] col_in_786,
    input  [15:0] col_in_787,
    input  [15:0] col_in_788,
    input  [15:0] col_in_789,
    input  [15:0] col_in_790,
    input  [15:0] col_in_791,
    input  [15:0] col_in_792,
    input  [15:0] col_in_793,
    input  [15:0] col_in_794,
    input  [15:0] col_in_795,
    input  [15:0] col_in_796,
    input  [15:0] col_in_797,
    input  [15:0] col_in_798,
    input  [15:0] col_in_799,
    input  [15:0] col_in_800,
    input  [15:0] col_in_801,
    input  [15:0] col_in_802,
    input  [15:0] col_in_803,
    input  [15:0] col_in_804,
    input  [15:0] col_in_805,
    input  [15:0] col_in_806,
    input  [15:0] col_in_807,
    input  [15:0] col_in_808,
    input  [15:0] col_in_809,
    input  [15:0] col_in_810,
    input  [15:0] col_in_811,
    input  [15:0] col_in_812,
    input  [15:0] col_in_813,
    input  [15:0] col_in_814,
    input  [15:0] col_in_815,
    input  [15:0] col_in_816,
    input  [15:0] col_in_817,
    input  [15:0] col_in_818,
    input  [15:0] col_in_819,
    input  [15:0] col_in_820,
    input  [15:0] col_in_821,
    input  [15:0] col_in_822,
    input  [15:0] col_in_823,
    input  [15:0] col_in_824,
    input  [15:0] col_in_825,
    input  [15:0] col_in_826,
    input  [15:0] col_in_827,
    input  [15:0] col_in_828,
    input  [15:0] col_in_829,
    input  [15:0] col_in_830,
    input  [15:0] col_in_831,
    input  [15:0] col_in_832,
    input  [15:0] col_in_833,
    input  [15:0] col_in_834,
    input  [15:0] col_in_835,
    input  [15:0] col_in_836,
    input  [15:0] col_in_837,
    input  [15:0] col_in_838,
    input  [15:0] col_in_839,
    input  [15:0] col_in_840,
    input  [15:0] col_in_841,
    input  [15:0] col_in_842,
    input  [15:0] col_in_843,
    input  [15:0] col_in_844,
    input  [15:0] col_in_845,
    input  [15:0] col_in_846,
    input  [15:0] col_in_847,
    input  [15:0] col_in_848,
    input  [15:0] col_in_849,
    input  [15:0] col_in_850,
    input  [15:0] col_in_851,
    input  [15:0] col_in_852,
    input  [15:0] col_in_853,
    input  [15:0] col_in_854,
    input  [15:0] col_in_855,
    input  [15:0] col_in_856,
    input  [15:0] col_in_857,
    input  [15:0] col_in_858,
    input  [15:0] col_in_859,
    input  [15:0] col_in_860,
    input  [15:0] col_in_861,
    input  [15:0] col_in_862,
    input  [15:0] col_in_863,
    input  [15:0] col_in_864,
    input  [15:0] col_in_865,
    input  [15:0] col_in_866,
    input  [15:0] col_in_867,
    input  [15:0] col_in_868,
    input  [15:0] col_in_869,
    input  [15:0] col_in_870,
    input  [15:0] col_in_871,
    input  [15:0] col_in_872,
    input  [15:0] col_in_873,
    input  [15:0] col_in_874,
    input  [15:0] col_in_875,
    input  [15:0] col_in_876,
    input  [15:0] col_in_877,
    input  [15:0] col_in_878,
    input  [15:0] col_in_879,
    input  [15:0] col_in_880,
    input  [15:0] col_in_881,
    input  [15:0] col_in_882,
    input  [15:0] col_in_883,
    input  [15:0] col_in_884,
    input  [15:0] col_in_885,
    input  [15:0] col_in_886,
    input  [15:0] col_in_887,
    input  [15:0] col_in_888,
    input  [15:0] col_in_889,
    input  [15:0] col_in_890,
    input  [15:0] col_in_891,
    input  [15:0] col_in_892,
    input  [15:0] col_in_893,
    input  [15:0] col_in_894,
    input  [15:0] col_in_895,
    input  [15:0] col_in_896,
    input  [15:0] col_in_897,
    input  [15:0] col_in_898,
    input  [15:0] col_in_899,
    input  [15:0] col_in_900,
    input  [15:0] col_in_901,
    input  [15:0] col_in_902,
    input  [15:0] col_in_903,
    input  [15:0] col_in_904,
    input  [15:0] col_in_905,
    input  [15:0] col_in_906,
    input  [15:0] col_in_907,
    input  [15:0] col_in_908,
    input  [15:0] col_in_909,
    input  [15:0] col_in_910,
    input  [15:0] col_in_911,
    input  [15:0] col_in_912,
    input  [15:0] col_in_913,
    input  [15:0] col_in_914,
    input  [15:0] col_in_915,
    input  [15:0] col_in_916,
    input  [15:0] col_in_917,
    input  [15:0] col_in_918,
    input  [15:0] col_in_919,
    input  [15:0] col_in_920,
    input  [15:0] col_in_921,
    input  [15:0] col_in_922,
    input  [15:0] col_in_923,
    input  [15:0] col_in_924,
    input  [15:0] col_in_925,
    input  [15:0] col_in_926,
    input  [15:0] col_in_927,
    input  [15:0] col_in_928,
    input  [15:0] col_in_929,
    input  [15:0] col_in_930,
    input  [15:0] col_in_931,
    input  [15:0] col_in_932,
    input  [15:0] col_in_933,
    input  [15:0] col_in_934,
    input  [15:0] col_in_935,
    input  [15:0] col_in_936,
    input  [15:0] col_in_937,
    input  [15:0] col_in_938,
    input  [15:0] col_in_939,
    input  [15:0] col_in_940,
    input  [15:0] col_in_941,
    input  [15:0] col_in_942,
    input  [15:0] col_in_943,
    input  [15:0] col_in_944,
    input  [15:0] col_in_945,
    input  [15:0] col_in_946,
    input  [15:0] col_in_947,
    input  [15:0] col_in_948,
    input  [15:0] col_in_949,
    input  [15:0] col_in_950,
    input  [15:0] col_in_951,
    input  [15:0] col_in_952,
    input  [15:0] col_in_953,
    input  [15:0] col_in_954,
    input  [15:0] col_in_955,
    input  [15:0] col_in_956,
    input  [15:0] col_in_957,
    input  [15:0] col_in_958,
    input  [15:0] col_in_959,
    input  [15:0] col_in_960,
    input  [15:0] col_in_961,
    input  [15:0] col_in_962,
    input  [15:0] col_in_963,
    input  [15:0] col_in_964,
    input  [15:0] col_in_965,
    input  [15:0] col_in_966,
    input  [15:0] col_in_967,
    input  [15:0] col_in_968,
    input  [15:0] col_in_969,
    input  [15:0] col_in_970,
    input  [15:0] col_in_971,
    input  [15:0] col_in_972,
    input  [15:0] col_in_973,
    input  [15:0] col_in_974,
    input  [15:0] col_in_975,
    input  [15:0] col_in_976,
    input  [15:0] col_in_977,
    input  [15:0] col_in_978,
    input  [15:0] col_in_979,
    input  [15:0] col_in_980,
    input  [15:0] col_in_981,
    input  [15:0] col_in_982,
    input  [15:0] col_in_983,
    input  [15:0] col_in_984,
    input  [15:0] col_in_985,
    input  [15:0] col_in_986,
    input  [15:0] col_in_987,
    input  [15:0] col_in_988,
    input  [15:0] col_in_989,
    input  [15:0] col_in_990,
    input  [15:0] col_in_991,
    input  [15:0] col_in_992,
    input  [15:0] col_in_993,
    input  [15:0] col_in_994,
    input  [15:0] col_in_995,
    input  [15:0] col_in_996,
    input  [15:0] col_in_997,
    input  [15:0] col_in_998,
    input  [15:0] col_in_999,
    input  [15:0] col_in_1000,
    input  [15:0] col_in_1001,
    input  [15:0] col_in_1002,
    input  [15:0] col_in_1003,
    input  [15:0] col_in_1004,
    input  [15:0] col_in_1005,
    input  [15:0] col_in_1006,
    input  [15:0] col_in_1007,
    input  [15:0] col_in_1008,
    input  [15:0] col_in_1009,
    input  [15:0] col_in_1010,
    input  [15:0] col_in_1011,
    input  [15:0] col_in_1012,
    input  [15:0] col_in_1013,
    input  [15:0] col_in_1014,
    input  [15:0] col_in_1015,
    input  [15:0] col_in_1016,
    input  [15:0] col_in_1017,
    input  [15:0] col_in_1018,
    input  [15:0] col_in_1019,
    input  [15:0] col_in_1020,
    input  [15:0] col_in_1021,
    input  [15:0] col_in_1022,
    input  [15:0] col_in_1023,
    input  [15:0] col_in_1024,
    input  [15:0] col_in_1025,
    input  [15:0] col_in_1026,
    input  [15:0] col_in_1027,
    input  [15:0] col_in_1028,
    input  [15:0] col_in_1029,
    input  [15:0] col_in_1030,
    input  [15:0] col_in_1031,
    input  [15:0] col_in_1032,

    output [11:0] col_out_0,
    output [11:0] col_out_1,
    output [11:0] col_out_2,
    output [11:0] col_out_3,
    output [11:0] col_out_4,
    output [11:0] col_out_5,
    output [11:0] col_out_6,
    output [11:0] col_out_7,
    output [11:0] col_out_8,
    output [11:0] col_out_9,
    output [11:0] col_out_10,
    output [11:0] col_out_11,
    output [11:0] col_out_12,
    output [11:0] col_out_13,
    output [11:0] col_out_14,
    output [11:0] col_out_15,
    output [11:0] col_out_16,
    output [11:0] col_out_17,
    output [11:0] col_out_18,
    output [11:0] col_out_19,
    output [11:0] col_out_20,
    output [11:0] col_out_21,
    output [11:0] col_out_22,
    output [11:0] col_out_23,
    output [11:0] col_out_24,
    output [11:0] col_out_25,
    output [11:0] col_out_26,
    output [11:0] col_out_27,
    output [11:0] col_out_28,
    output [11:0] col_out_29,
    output [11:0] col_out_30,
    output [11:0] col_out_31,
    output [11:0] col_out_32,
    output [11:0] col_out_33,
    output [11:0] col_out_34,
    output [11:0] col_out_35,
    output [11:0] col_out_36,
    output [11:0] col_out_37,
    output [11:0] col_out_38,
    output [11:0] col_out_39,
    output [11:0] col_out_40,
    output [11:0] col_out_41,
    output [11:0] col_out_42,
    output [11:0] col_out_43,
    output [11:0] col_out_44,
    output [11:0] col_out_45,
    output [11:0] col_out_46,
    output [11:0] col_out_47,
    output [11:0] col_out_48,
    output [11:0] col_out_49,
    output [11:0] col_out_50,
    output [11:0] col_out_51,
    output [11:0] col_out_52,
    output [11:0] col_out_53,
    output [11:0] col_out_54,
    output [11:0] col_out_55,
    output [11:0] col_out_56,
    output [11:0] col_out_57,
    output [11:0] col_out_58,
    output [11:0] col_out_59,
    output [11:0] col_out_60,
    output [11:0] col_out_61,
    output [11:0] col_out_62,
    output [11:0] col_out_63,
    output [11:0] col_out_64,
    output [11:0] col_out_65,
    output [11:0] col_out_66,
    output [11:0] col_out_67,
    output [11:0] col_out_68,
    output [11:0] col_out_69,
    output [11:0] col_out_70,
    output [11:0] col_out_71,
    output [11:0] col_out_72,
    output [11:0] col_out_73,
    output [11:0] col_out_74,
    output [11:0] col_out_75,
    output [11:0] col_out_76,
    output [11:0] col_out_77,
    output [11:0] col_out_78,
    output [11:0] col_out_79,
    output [11:0] col_out_80,
    output [11:0] col_out_81,
    output [11:0] col_out_82,
    output [11:0] col_out_83,
    output [11:0] col_out_84,
    output [11:0] col_out_85,
    output [11:0] col_out_86,
    output [11:0] col_out_87,
    output [11:0] col_out_88,
    output [11:0] col_out_89,
    output [11:0] col_out_90,
    output [11:0] col_out_91,
    output [11:0] col_out_92,
    output [11:0] col_out_93,
    output [11:0] col_out_94,
    output [11:0] col_out_95,
    output [11:0] col_out_96,
    output [11:0] col_out_97,
    output [11:0] col_out_98,
    output [11:0] col_out_99,
    output [11:0] col_out_100,
    output [11:0] col_out_101,
    output [11:0] col_out_102,
    output [11:0] col_out_103,
    output [11:0] col_out_104,
    output [11:0] col_out_105,
    output [11:0] col_out_106,
    output [11:0] col_out_107,
    output [11:0] col_out_108,
    output [11:0] col_out_109,
    output [11:0] col_out_110,
    output [11:0] col_out_111,
    output [11:0] col_out_112,
    output [11:0] col_out_113,
    output [11:0] col_out_114,
    output [11:0] col_out_115,
    output [11:0] col_out_116,
    output [11:0] col_out_117,
    output [11:0] col_out_118,
    output [11:0] col_out_119,
    output [11:0] col_out_120,
    output [11:0] col_out_121,
    output [11:0] col_out_122,
    output [11:0] col_out_123,
    output [11:0] col_out_124,
    output [11:0] col_out_125,
    output [11:0] col_out_126,
    output [11:0] col_out_127,
    output [11:0] col_out_128,
    output [11:0] col_out_129,
    output [11:0] col_out_130,
    output [11:0] col_out_131,
    output [11:0] col_out_132,
    output [11:0] col_out_133,
    output [11:0] col_out_134,
    output [11:0] col_out_135,
    output [11:0] col_out_136,
    output [11:0] col_out_137,
    output [11:0] col_out_138,
    output [11:0] col_out_139,
    output [11:0] col_out_140,
    output [11:0] col_out_141,
    output [11:0] col_out_142,
    output [11:0] col_out_143,
    output [11:0] col_out_144,
    output [11:0] col_out_145,
    output [11:0] col_out_146,
    output [11:0] col_out_147,
    output [11:0] col_out_148,
    output [11:0] col_out_149,
    output [11:0] col_out_150,
    output [11:0] col_out_151,
    output [11:0] col_out_152,
    output [11:0] col_out_153,
    output [11:0] col_out_154,
    output [11:0] col_out_155,
    output [11:0] col_out_156,
    output [11:0] col_out_157,
    output [11:0] col_out_158,
    output [11:0] col_out_159,
    output [11:0] col_out_160,
    output [11:0] col_out_161,
    output [11:0] col_out_162,
    output [11:0] col_out_163,
    output [11:0] col_out_164,
    output [11:0] col_out_165,
    output [11:0] col_out_166,
    output [11:0] col_out_167,
    output [11:0] col_out_168,
    output [11:0] col_out_169,
    output [11:0] col_out_170,
    output [11:0] col_out_171,
    output [11:0] col_out_172,
    output [11:0] col_out_173,
    output [11:0] col_out_174,
    output [11:0] col_out_175,
    output [11:0] col_out_176,
    output [11:0] col_out_177,
    output [11:0] col_out_178,
    output [11:0] col_out_179,
    output [11:0] col_out_180,
    output [11:0] col_out_181,
    output [11:0] col_out_182,
    output [11:0] col_out_183,
    output [11:0] col_out_184,
    output [11:0] col_out_185,
    output [11:0] col_out_186,
    output [11:0] col_out_187,
    output [11:0] col_out_188,
    output [11:0] col_out_189,
    output [11:0] col_out_190,
    output [11:0] col_out_191,
    output [11:0] col_out_192,
    output [11:0] col_out_193,
    output [11:0] col_out_194,
    output [11:0] col_out_195,
    output [11:0] col_out_196,
    output [11:0] col_out_197,
    output [11:0] col_out_198,
    output [11:0] col_out_199,
    output [11:0] col_out_200,
    output [11:0] col_out_201,
    output [11:0] col_out_202,
    output [11:0] col_out_203,
    output [11:0] col_out_204,
    output [11:0] col_out_205,
    output [11:0] col_out_206,
    output [11:0] col_out_207,
    output [11:0] col_out_208,
    output [11:0] col_out_209,
    output [11:0] col_out_210,
    output [11:0] col_out_211,
    output [11:0] col_out_212,
    output [11:0] col_out_213,
    output [11:0] col_out_214,
    output [11:0] col_out_215,
    output [11:0] col_out_216,
    output [11:0] col_out_217,
    output [11:0] col_out_218,
    output [11:0] col_out_219,
    output [11:0] col_out_220,
    output [11:0] col_out_221,
    output [11:0] col_out_222,
    output [11:0] col_out_223,
    output [11:0] col_out_224,
    output [11:0] col_out_225,
    output [11:0] col_out_226,
    output [11:0] col_out_227,
    output [11:0] col_out_228,
    output [11:0] col_out_229,
    output [11:0] col_out_230,
    output [11:0] col_out_231,
    output [11:0] col_out_232,
    output [11:0] col_out_233,
    output [11:0] col_out_234,
    output [11:0] col_out_235,
    output [11:0] col_out_236,
    output [11:0] col_out_237,
    output [11:0] col_out_238,
    output [11:0] col_out_239,
    output [11:0] col_out_240,
    output [11:0] col_out_241,
    output [11:0] col_out_242,
    output [11:0] col_out_243,
    output [11:0] col_out_244,
    output [11:0] col_out_245,
    output [11:0] col_out_246,
    output [11:0] col_out_247,
    output [11:0] col_out_248,
    output [11:0] col_out_249,
    output [11:0] col_out_250,
    output [11:0] col_out_251,
    output [11:0] col_out_252,
    output [11:0] col_out_253,
    output [11:0] col_out_254,
    output [11:0] col_out_255,
    output [11:0] col_out_256,
    output [11:0] col_out_257,
    output [11:0] col_out_258,
    output [11:0] col_out_259,
    output [11:0] col_out_260,
    output [11:0] col_out_261,
    output [11:0] col_out_262,
    output [11:0] col_out_263,
    output [11:0] col_out_264,
    output [11:0] col_out_265,
    output [11:0] col_out_266,
    output [11:0] col_out_267,
    output [11:0] col_out_268,
    output [11:0] col_out_269,
    output [11:0] col_out_270,
    output [11:0] col_out_271,
    output [11:0] col_out_272,
    output [11:0] col_out_273,
    output [11:0] col_out_274,
    output [11:0] col_out_275,
    output [11:0] col_out_276,
    output [11:0] col_out_277,
    output [11:0] col_out_278,
    output [11:0] col_out_279,
    output [11:0] col_out_280,
    output [11:0] col_out_281,
    output [11:0] col_out_282,
    output [11:0] col_out_283,
    output [11:0] col_out_284,
    output [11:0] col_out_285,
    output [11:0] col_out_286,
    output [11:0] col_out_287,
    output [11:0] col_out_288,
    output [11:0] col_out_289,
    output [11:0] col_out_290,
    output [11:0] col_out_291,
    output [11:0] col_out_292,
    output [11:0] col_out_293,
    output [11:0] col_out_294,
    output [11:0] col_out_295,
    output [11:0] col_out_296,
    output [11:0] col_out_297,
    output [11:0] col_out_298,
    output [11:0] col_out_299,
    output [11:0] col_out_300,
    output [11:0] col_out_301,
    output [11:0] col_out_302,
    output [11:0] col_out_303,
    output [11:0] col_out_304,
    output [11:0] col_out_305,
    output [11:0] col_out_306,
    output [11:0] col_out_307,
    output [11:0] col_out_308,
    output [11:0] col_out_309,
    output [11:0] col_out_310,
    output [11:0] col_out_311,
    output [11:0] col_out_312,
    output [11:0] col_out_313,
    output [11:0] col_out_314,
    output [11:0] col_out_315,
    output [11:0] col_out_316,
    output [11:0] col_out_317,
    output [11:0] col_out_318,
    output [11:0] col_out_319,
    output [11:0] col_out_320,
    output [11:0] col_out_321,
    output [11:0] col_out_322,
    output [11:0] col_out_323,
    output [11:0] col_out_324,
    output [11:0] col_out_325,
    output [11:0] col_out_326,
    output [11:0] col_out_327,
    output [11:0] col_out_328,
    output [11:0] col_out_329,
    output [11:0] col_out_330,
    output [11:0] col_out_331,
    output [11:0] col_out_332,
    output [11:0] col_out_333,
    output [11:0] col_out_334,
    output [11:0] col_out_335,
    output [11:0] col_out_336,
    output [11:0] col_out_337,
    output [11:0] col_out_338,
    output [11:0] col_out_339,
    output [11:0] col_out_340,
    output [11:0] col_out_341,
    output [11:0] col_out_342,
    output [11:0] col_out_343,
    output [11:0] col_out_344,
    output [11:0] col_out_345,
    output [11:0] col_out_346,
    output [11:0] col_out_347,
    output [11:0] col_out_348,
    output [11:0] col_out_349,
    output [11:0] col_out_350,
    output [11:0] col_out_351,
    output [11:0] col_out_352,
    output [11:0] col_out_353,
    output [11:0] col_out_354,
    output [11:0] col_out_355,
    output [11:0] col_out_356,
    output [11:0] col_out_357,
    output [11:0] col_out_358,
    output [11:0] col_out_359,
    output [11:0] col_out_360,
    output [11:0] col_out_361,
    output [11:0] col_out_362,
    output [11:0] col_out_363,
    output [11:0] col_out_364,
    output [11:0] col_out_365,
    output [11:0] col_out_366,
    output [11:0] col_out_367,
    output [11:0] col_out_368,
    output [11:0] col_out_369,
    output [11:0] col_out_370,
    output [11:0] col_out_371,
    output [11:0] col_out_372,
    output [11:0] col_out_373,
    output [11:0] col_out_374,
    output [11:0] col_out_375,
    output [11:0] col_out_376,
    output [11:0] col_out_377,
    output [11:0] col_out_378,
    output [11:0] col_out_379,
    output [11:0] col_out_380,
    output [11:0] col_out_381,
    output [11:0] col_out_382,
    output [11:0] col_out_383,
    output [11:0] col_out_384,
    output [11:0] col_out_385,
    output [11:0] col_out_386,
    output [11:0] col_out_387,
    output [11:0] col_out_388,
    output [11:0] col_out_389,
    output [11:0] col_out_390,
    output [11:0] col_out_391,
    output [11:0] col_out_392,
    output [11:0] col_out_393,
    output [11:0] col_out_394,
    output [11:0] col_out_395,
    output [11:0] col_out_396,
    output [11:0] col_out_397,
    output [11:0] col_out_398,
    output [11:0] col_out_399,
    output [11:0] col_out_400,
    output [11:0] col_out_401,
    output [11:0] col_out_402,
    output [11:0] col_out_403,
    output [11:0] col_out_404,
    output [11:0] col_out_405,
    output [11:0] col_out_406,
    output [11:0] col_out_407,
    output [11:0] col_out_408,
    output [11:0] col_out_409,
    output [11:0] col_out_410,
    output [11:0] col_out_411,
    output [11:0] col_out_412,
    output [11:0] col_out_413,
    output [11:0] col_out_414,
    output [11:0] col_out_415,
    output [11:0] col_out_416,
    output [11:0] col_out_417,
    output [11:0] col_out_418,
    output [11:0] col_out_419,
    output [11:0] col_out_420,
    output [11:0] col_out_421,
    output [11:0] col_out_422,
    output [11:0] col_out_423,
    output [11:0] col_out_424,
    output [11:0] col_out_425,
    output [11:0] col_out_426,
    output [11:0] col_out_427,
    output [11:0] col_out_428,
    output [11:0] col_out_429,
    output [11:0] col_out_430,
    output [11:0] col_out_431,
    output [11:0] col_out_432,
    output [11:0] col_out_433,
    output [11:0] col_out_434,
    output [11:0] col_out_435,
    output [11:0] col_out_436,
    output [11:0] col_out_437,
    output [11:0] col_out_438,
    output [11:0] col_out_439,
    output [11:0] col_out_440,
    output [11:0] col_out_441,
    output [11:0] col_out_442,
    output [11:0] col_out_443,
    output [11:0] col_out_444,
    output [11:0] col_out_445,
    output [11:0] col_out_446,
    output [11:0] col_out_447,
    output [11:0] col_out_448,
    output [11:0] col_out_449,
    output [11:0] col_out_450,
    output [11:0] col_out_451,
    output [11:0] col_out_452,
    output [11:0] col_out_453,
    output [11:0] col_out_454,
    output [11:0] col_out_455,
    output [11:0] col_out_456,
    output [11:0] col_out_457,
    output [11:0] col_out_458,
    output [11:0] col_out_459,
    output [11:0] col_out_460,
    output [11:0] col_out_461,
    output [11:0] col_out_462,
    output [11:0] col_out_463,
    output [11:0] col_out_464,
    output [11:0] col_out_465,
    output [11:0] col_out_466,
    output [11:0] col_out_467,
    output [11:0] col_out_468,
    output [11:0] col_out_469,
    output [11:0] col_out_470,
    output [11:0] col_out_471,
    output [11:0] col_out_472,
    output [11:0] col_out_473,
    output [11:0] col_out_474,
    output [11:0] col_out_475,
    output [11:0] col_out_476,
    output [11:0] col_out_477,
    output [11:0] col_out_478,
    output [11:0] col_out_479,
    output [11:0] col_out_480,
    output [11:0] col_out_481,
    output [11:0] col_out_482,
    output [11:0] col_out_483,
    output [11:0] col_out_484,
    output [11:0] col_out_485,
    output [11:0] col_out_486,
    output [11:0] col_out_487,
    output [11:0] col_out_488,
    output [11:0] col_out_489,
    output [11:0] col_out_490,
    output [11:0] col_out_491,
    output [11:0] col_out_492,
    output [11:0] col_out_493,
    output [11:0] col_out_494,
    output [11:0] col_out_495,
    output [11:0] col_out_496,
    output [11:0] col_out_497,
    output [11:0] col_out_498,
    output [11:0] col_out_499,
    output [11:0] col_out_500,
    output [11:0] col_out_501,
    output [11:0] col_out_502,
    output [11:0] col_out_503,
    output [11:0] col_out_504,
    output [11:0] col_out_505,
    output [11:0] col_out_506,
    output [11:0] col_out_507,
    output [11:0] col_out_508,
    output [11:0] col_out_509,
    output [11:0] col_out_510,
    output [11:0] col_out_511,
    output [11:0] col_out_512,
    output [11:0] col_out_513,
    output [11:0] col_out_514,
    output [11:0] col_out_515,
    output [11:0] col_out_516,
    output [11:0] col_out_517,
    output [11:0] col_out_518,
    output [11:0] col_out_519,
    output [11:0] col_out_520,
    output [11:0] col_out_521,
    output [11:0] col_out_522,
    output [11:0] col_out_523,
    output [11:0] col_out_524,
    output [11:0] col_out_525,
    output [11:0] col_out_526,
    output [11:0] col_out_527,
    output [11:0] col_out_528,
    output [11:0] col_out_529,
    output [11:0] col_out_530,
    output [11:0] col_out_531,
    output [11:0] col_out_532,
    output [11:0] col_out_533,
    output [11:0] col_out_534,
    output [11:0] col_out_535,
    output [11:0] col_out_536,
    output [11:0] col_out_537,
    output [11:0] col_out_538,
    output [11:0] col_out_539,
    output [11:0] col_out_540,
    output [11:0] col_out_541,
    output [11:0] col_out_542,
    output [11:0] col_out_543,
    output [11:0] col_out_544,
    output [11:0] col_out_545,
    output [11:0] col_out_546,
    output [11:0] col_out_547,
    output [11:0] col_out_548,
    output [11:0] col_out_549,
    output [11:0] col_out_550,
    output [11:0] col_out_551,
    output [11:0] col_out_552,
    output [11:0] col_out_553,
    output [11:0] col_out_554,
    output [11:0] col_out_555,
    output [11:0] col_out_556,
    output [11:0] col_out_557,
    output [11:0] col_out_558,
    output [11:0] col_out_559,
    output [11:0] col_out_560,
    output [11:0] col_out_561,
    output [11:0] col_out_562,
    output [11:0] col_out_563,
    output [11:0] col_out_564,
    output [11:0] col_out_565,
    output [11:0] col_out_566,
    output [11:0] col_out_567,
    output [11:0] col_out_568,
    output [11:0] col_out_569,
    output [11:0] col_out_570,
    output [11:0] col_out_571,
    output [11:0] col_out_572,
    output [11:0] col_out_573,
    output [11:0] col_out_574,
    output [11:0] col_out_575,
    output [11:0] col_out_576,
    output [11:0] col_out_577,
    output [11:0] col_out_578,
    output [11:0] col_out_579,
    output [11:0] col_out_580,
    output [11:0] col_out_581,
    output [11:0] col_out_582,
    output [11:0] col_out_583,
    output [11:0] col_out_584,
    output [11:0] col_out_585,
    output [11:0] col_out_586,
    output [11:0] col_out_587,
    output [11:0] col_out_588,
    output [11:0] col_out_589,
    output [11:0] col_out_590,
    output [11:0] col_out_591,
    output [11:0] col_out_592,
    output [11:0] col_out_593,
    output [11:0] col_out_594,
    output [11:0] col_out_595,
    output [11:0] col_out_596,
    output [11:0] col_out_597,
    output [11:0] col_out_598,
    output [11:0] col_out_599,
    output [11:0] col_out_600,
    output [11:0] col_out_601,
    output [11:0] col_out_602,
    output [11:0] col_out_603,
    output [11:0] col_out_604,
    output [11:0] col_out_605,
    output [11:0] col_out_606,
    output [11:0] col_out_607,
    output [11:0] col_out_608,
    output [11:0] col_out_609,
    output [11:0] col_out_610,
    output [11:0] col_out_611,
    output [11:0] col_out_612,
    output [11:0] col_out_613,
    output [11:0] col_out_614,
    output [11:0] col_out_615,
    output [11:0] col_out_616,
    output [11:0] col_out_617,
    output [11:0] col_out_618,
    output [11:0] col_out_619,
    output [11:0] col_out_620,
    output [11:0] col_out_621,
    output [11:0] col_out_622,
    output [11:0] col_out_623,
    output [11:0] col_out_624,
    output [11:0] col_out_625,
    output [11:0] col_out_626,
    output [11:0] col_out_627,
    output [11:0] col_out_628,
    output [11:0] col_out_629,
    output [11:0] col_out_630,
    output [11:0] col_out_631,
    output [11:0] col_out_632,
    output [11:0] col_out_633,
    output [11:0] col_out_634,
    output [11:0] col_out_635,
    output [11:0] col_out_636,
    output [11:0] col_out_637,
    output [11:0] col_out_638,
    output [11:0] col_out_639,
    output [11:0] col_out_640,
    output [11:0] col_out_641,
    output [11:0] col_out_642,
    output [11:0] col_out_643,
    output [11:0] col_out_644,
    output [11:0] col_out_645,
    output [11:0] col_out_646,
    output [11:0] col_out_647,
    output [11:0] col_out_648,
    output [11:0] col_out_649,
    output [11:0] col_out_650,
    output [11:0] col_out_651,
    output [11:0] col_out_652,
    output [11:0] col_out_653,
    output [11:0] col_out_654,
    output [11:0] col_out_655,
    output [11:0] col_out_656,
    output [11:0] col_out_657,
    output [11:0] col_out_658,
    output [11:0] col_out_659,
    output [11:0] col_out_660,
    output [11:0] col_out_661,
    output [11:0] col_out_662,
    output [11:0] col_out_663,
    output [11:0] col_out_664,
    output [11:0] col_out_665,
    output [11:0] col_out_666,
    output [11:0] col_out_667,
    output [11:0] col_out_668,
    output [11:0] col_out_669,
    output [11:0] col_out_670,
    output [11:0] col_out_671,
    output [11:0] col_out_672,
    output [11:0] col_out_673,
    output [11:0] col_out_674,
    output [11:0] col_out_675,
    output [11:0] col_out_676,
    output [11:0] col_out_677,
    output [11:0] col_out_678,
    output [11:0] col_out_679,
    output [11:0] col_out_680,
    output [11:0] col_out_681,
    output [11:0] col_out_682,
    output [11:0] col_out_683,
    output [11:0] col_out_684,
    output [11:0] col_out_685,
    output [11:0] col_out_686,
    output [11:0] col_out_687,
    output [11:0] col_out_688,
    output [11:0] col_out_689,
    output [11:0] col_out_690,
    output [11:0] col_out_691,
    output [11:0] col_out_692,
    output [11:0] col_out_693,
    output [11:0] col_out_694,
    output [11:0] col_out_695,
    output [11:0] col_out_696,
    output [11:0] col_out_697,
    output [11:0] col_out_698,
    output [11:0] col_out_699,
    output [11:0] col_out_700,
    output [11:0] col_out_701,
    output [11:0] col_out_702,
    output [11:0] col_out_703,
    output [11:0] col_out_704,
    output [11:0] col_out_705,
    output [11:0] col_out_706,
    output [11:0] col_out_707,
    output [11:0] col_out_708,
    output [11:0] col_out_709,
    output [11:0] col_out_710,
    output [11:0] col_out_711,
    output [11:0] col_out_712,
    output [11:0] col_out_713,
    output [11:0] col_out_714,
    output [11:0] col_out_715,
    output [11:0] col_out_716,
    output [11:0] col_out_717,
    output [11:0] col_out_718,
    output [11:0] col_out_719,
    output [11:0] col_out_720,
    output [11:0] col_out_721,
    output [11:0] col_out_722,
    output [11:0] col_out_723,
    output [11:0] col_out_724,
    output [11:0] col_out_725,
    output [11:0] col_out_726,
    output [11:0] col_out_727,
    output [11:0] col_out_728,
    output [11:0] col_out_729,
    output [11:0] col_out_730,
    output [11:0] col_out_731,
    output [11:0] col_out_732,
    output [11:0] col_out_733,
    output [11:0] col_out_734,
    output [11:0] col_out_735,
    output [11:0] col_out_736,
    output [11:0] col_out_737,
    output [11:0] col_out_738,
    output [11:0] col_out_739,
    output [11:0] col_out_740,
    output [11:0] col_out_741,
    output [11:0] col_out_742,
    output [11:0] col_out_743,
    output [11:0] col_out_744,
    output [11:0] col_out_745,
    output [11:0] col_out_746,
    output [11:0] col_out_747,
    output [11:0] col_out_748,
    output [11:0] col_out_749,
    output [11:0] col_out_750,
    output [11:0] col_out_751,
    output [11:0] col_out_752,
    output [11:0] col_out_753,
    output [11:0] col_out_754,
    output [11:0] col_out_755,
    output [11:0] col_out_756,
    output [11:0] col_out_757,
    output [11:0] col_out_758,
    output [11:0] col_out_759,
    output [11:0] col_out_760,
    output [11:0] col_out_761,
    output [11:0] col_out_762,
    output [11:0] col_out_763,
    output [11:0] col_out_764,
    output [11:0] col_out_765,
    output [11:0] col_out_766,
    output [11:0] col_out_767,
    output [11:0] col_out_768,
    output [11:0] col_out_769,
    output [11:0] col_out_770,
    output [11:0] col_out_771,
    output [11:0] col_out_772,
    output [11:0] col_out_773,
    output [11:0] col_out_774,
    output [11:0] col_out_775,
    output [11:0] col_out_776,
    output [11:0] col_out_777,
    output [11:0] col_out_778,
    output [11:0] col_out_779,
    output [11:0] col_out_780,
    output [11:0] col_out_781,
    output [11:0] col_out_782,
    output [11:0] col_out_783,
    output [11:0] col_out_784,
    output [11:0] col_out_785,
    output [11:0] col_out_786,
    output [11:0] col_out_787,
    output [11:0] col_out_788,
    output [11:0] col_out_789,
    output [11:0] col_out_790,
    output [11:0] col_out_791,
    output [11:0] col_out_792,
    output [11:0] col_out_793,
    output [11:0] col_out_794,
    output [11:0] col_out_795,
    output [11:0] col_out_796,
    output [11:0] col_out_797,
    output [11:0] col_out_798,
    output [11:0] col_out_799,
    output [11:0] col_out_800,
    output [11:0] col_out_801,
    output [11:0] col_out_802,
    output [11:0] col_out_803,
    output [11:0] col_out_804,
    output [11:0] col_out_805,
    output [11:0] col_out_806,
    output [11:0] col_out_807,
    output [11:0] col_out_808,
    output [11:0] col_out_809,
    output [11:0] col_out_810,
    output [11:0] col_out_811,
    output [11:0] col_out_812,
    output [11:0] col_out_813,
    output [11:0] col_out_814,
    output [11:0] col_out_815,
    output [11:0] col_out_816,
    output [11:0] col_out_817,
    output [11:0] col_out_818,
    output [11:0] col_out_819,
    output [11:0] col_out_820,
    output [11:0] col_out_821,
    output [11:0] col_out_822,
    output [11:0] col_out_823,
    output [11:0] col_out_824,
    output [11:0] col_out_825,
    output [11:0] col_out_826,
    output [11:0] col_out_827,
    output [11:0] col_out_828,
    output [11:0] col_out_829,
    output [11:0] col_out_830,
    output [11:0] col_out_831,
    output [11:0] col_out_832,
    output [11:0] col_out_833,
    output [11:0] col_out_834,
    output [11:0] col_out_835,
    output [11:0] col_out_836,
    output [11:0] col_out_837,
    output [11:0] col_out_838,
    output [11:0] col_out_839,
    output [11:0] col_out_840,
    output [11:0] col_out_841,
    output [11:0] col_out_842,
    output [11:0] col_out_843,
    output [11:0] col_out_844,
    output [11:0] col_out_845,
    output [11:0] col_out_846,
    output [11:0] col_out_847,
    output [11:0] col_out_848,
    output [11:0] col_out_849,
    output [11:0] col_out_850,
    output [11:0] col_out_851,
    output [11:0] col_out_852,
    output [11:0] col_out_853,
    output [11:0] col_out_854,
    output [11:0] col_out_855,
    output [11:0] col_out_856,
    output [11:0] col_out_857,
    output [11:0] col_out_858,
    output [11:0] col_out_859,
    output [11:0] col_out_860,
    output [11:0] col_out_861,
    output [11:0] col_out_862,
    output [11:0] col_out_863,
    output [11:0] col_out_864,
    output [11:0] col_out_865,
    output [11:0] col_out_866,
    output [11:0] col_out_867,
    output [11:0] col_out_868,
    output [11:0] col_out_869,
    output [11:0] col_out_870,
    output [11:0] col_out_871,
    output [11:0] col_out_872,
    output [11:0] col_out_873,
    output [11:0] col_out_874,
    output [11:0] col_out_875,
    output [11:0] col_out_876,
    output [11:0] col_out_877,
    output [11:0] col_out_878,
    output [11:0] col_out_879,
    output [11:0] col_out_880,
    output [11:0] col_out_881,
    output [11:0] col_out_882,
    output [11:0] col_out_883,
    output [11:0] col_out_884,
    output [11:0] col_out_885,
    output [11:0] col_out_886,
    output [11:0] col_out_887,
    output [11:0] col_out_888,
    output [11:0] col_out_889,
    output [11:0] col_out_890,
    output [11:0] col_out_891,
    output [11:0] col_out_892,
    output [11:0] col_out_893,
    output [11:0] col_out_894,
    output [11:0] col_out_895,
    output [11:0] col_out_896,
    output [11:0] col_out_897,
    output [11:0] col_out_898,
    output [11:0] col_out_899,
    output [11:0] col_out_900,
    output [11:0] col_out_901,
    output [11:0] col_out_902,
    output [11:0] col_out_903,
    output [11:0] col_out_904,
    output [11:0] col_out_905,
    output [11:0] col_out_906,
    output [11:0] col_out_907,
    output [11:0] col_out_908,
    output [11:0] col_out_909,
    output [11:0] col_out_910,
    output [11:0] col_out_911,
    output [11:0] col_out_912,
    output [11:0] col_out_913,
    output [11:0] col_out_914,
    output [11:0] col_out_915,
    output [11:0] col_out_916,
    output [11:0] col_out_917,
    output [11:0] col_out_918,
    output [11:0] col_out_919,
    output [11:0] col_out_920,
    output [11:0] col_out_921,
    output [11:0] col_out_922,
    output [11:0] col_out_923,
    output [11:0] col_out_924,
    output [11:0] col_out_925,
    output [11:0] col_out_926,
    output [11:0] col_out_927,
    output [11:0] col_out_928,
    output [11:0] col_out_929,
    output [11:0] col_out_930,
    output [11:0] col_out_931,
    output [11:0] col_out_932,
    output [11:0] col_out_933,
    output [11:0] col_out_934,
    output [11:0] col_out_935,
    output [11:0] col_out_936,
    output [11:0] col_out_937,
    output [11:0] col_out_938,
    output [11:0] col_out_939,
    output [11:0] col_out_940,
    output [11:0] col_out_941,
    output [11:0] col_out_942,
    output [11:0] col_out_943,
    output [11:0] col_out_944,
    output [11:0] col_out_945,
    output [11:0] col_out_946,
    output [11:0] col_out_947,
    output [11:0] col_out_948,
    output [11:0] col_out_949,
    output [11:0] col_out_950,
    output [11:0] col_out_951,
    output [11:0] col_out_952,
    output [11:0] col_out_953,
    output [11:0] col_out_954,
    output [11:0] col_out_955,
    output [11:0] col_out_956,
    output [11:0] col_out_957,
    output [11:0] col_out_958,
    output [11:0] col_out_959,
    output [11:0] col_out_960,
    output [11:0] col_out_961,
    output [11:0] col_out_962,
    output [11:0] col_out_963,
    output [11:0] col_out_964,
    output [11:0] col_out_965,
    output [11:0] col_out_966,
    output [11:0] col_out_967,
    output [11:0] col_out_968,
    output [11:0] col_out_969,
    output [11:0] col_out_970,
    output [11:0] col_out_971,
    output [11:0] col_out_972,
    output [11:0] col_out_973,
    output [11:0] col_out_974,
    output [11:0] col_out_975,
    output [11:0] col_out_976,
    output [11:0] col_out_977,
    output [11:0] col_out_978,
    output [11:0] col_out_979,
    output [11:0] col_out_980,
    output [11:0] col_out_981,
    output [11:0] col_out_982,
    output [11:0] col_out_983,
    output [11:0] col_out_984,
    output [11:0] col_out_985,
    output [11:0] col_out_986,
    output [11:0] col_out_987,
    output [11:0] col_out_988,
    output [11:0] col_out_989,
    output [11:0] col_out_990,
    output [11:0] col_out_991,
    output [11:0] col_out_992,
    output [11:0] col_out_993,
    output [11:0] col_out_994,
    output [11:0] col_out_995,
    output [11:0] col_out_996,
    output [11:0] col_out_997,
    output [11:0] col_out_998,
    output [11:0] col_out_999,
    output [11:0] col_out_1000,
    output [11:0] col_out_1001,
    output [11:0] col_out_1002,
    output [11:0] col_out_1003,
    output [11:0] col_out_1004,
    output [11:0] col_out_1005,
    output [11:0] col_out_1006,
    output [11:0] col_out_1007,
    output [11:0] col_out_1008,
    output [11:0] col_out_1009,
    output [11:0] col_out_1010,
    output [11:0] col_out_1011,
    output [11:0] col_out_1012,
    output [11:0] col_out_1013,
    output [11:0] col_out_1014,
    output [11:0] col_out_1015,
    output [11:0] col_out_1016,
    output [11:0] col_out_1017,
    output [11:0] col_out_1018,
    output [11:0] col_out_1019,
    output [11:0] col_out_1020,
    output [11:0] col_out_1021,
    output [11:0] col_out_1022,
    output [11:0] col_out_1023,
    output [11:0] col_out_1024,
    output [11:0] col_out_1025,
    output [11:0] col_out_1026,
    output [11:0] col_out_1027,
    output [11:0] col_out_1028,
    output [11:0] col_out_1029,
    output [11:0] col_out_1030,
    output [11:0] col_out_1031,
    output [11:0] col_out_1032,
    output [11:0] col_out_1033
);



//--compressor_array input and output----------------------

wire [17:0] u_ca_in_0;
wire [17:0] u_ca_in_1;
wire [17:0] u_ca_in_2;
wire [17:0] u_ca_in_3;
wire [17:0] u_ca_in_4;
wire [17:0] u_ca_in_5;
wire [17:0] u_ca_in_6;
wire [17:0] u_ca_in_7;
wire [17:0] u_ca_in_8;
wire [17:0] u_ca_in_9;
wire [17:0] u_ca_in_10;
wire [17:0] u_ca_in_11;
wire [17:0] u_ca_in_12;
wire [17:0] u_ca_in_13;
wire [17:0] u_ca_in_14;
wire [17:0] u_ca_in_15;
wire [17:0] u_ca_in_16;
wire [17:0] u_ca_in_17;
wire [17:0] u_ca_in_18;
wire [17:0] u_ca_in_19;
wire [17:0] u_ca_in_20;
wire [17:0] u_ca_in_21;
wire [17:0] u_ca_in_22;
wire [17:0] u_ca_in_23;
wire [17:0] u_ca_in_24;
wire [17:0] u_ca_in_25;
wire [17:0] u_ca_in_26;
wire [17:0] u_ca_in_27;
wire [17:0] u_ca_in_28;
wire [17:0] u_ca_in_29;
wire [17:0] u_ca_in_30;
wire [17:0] u_ca_in_31;
wire [17:0] u_ca_in_32;
wire [17:0] u_ca_in_33;
wire [17:0] u_ca_in_34;
wire [17:0] u_ca_in_35;
wire [17:0] u_ca_in_36;
wire [17:0] u_ca_in_37;
wire [17:0] u_ca_in_38;
wire [17:0] u_ca_in_39;
wire [17:0] u_ca_in_40;
wire [17:0] u_ca_in_41;
wire [17:0] u_ca_in_42;
wire [17:0] u_ca_in_43;
wire [17:0] u_ca_in_44;
wire [17:0] u_ca_in_45;
wire [17:0] u_ca_in_46;
wire [17:0] u_ca_in_47;
wire [17:0] u_ca_in_48;
wire [17:0] u_ca_in_49;
wire [17:0] u_ca_in_50;
wire [17:0] u_ca_in_51;
wire [17:0] u_ca_in_52;
wire [17:0] u_ca_in_53;
wire [17:0] u_ca_in_54;
wire [17:0] u_ca_in_55;
wire [17:0] u_ca_in_56;
wire [17:0] u_ca_in_57;
wire [17:0] u_ca_in_58;
wire [17:0] u_ca_in_59;
wire [17:0] u_ca_in_60;
wire [17:0] u_ca_in_61;
wire [17:0] u_ca_in_62;
wire [17:0] u_ca_in_63;
wire [17:0] u_ca_in_64;
wire [17:0] u_ca_in_65;
wire [17:0] u_ca_in_66;
wire [17:0] u_ca_in_67;
wire [17:0] u_ca_in_68;
wire [17:0] u_ca_in_69;
wire [17:0] u_ca_in_70;
wire [17:0] u_ca_in_71;
wire [17:0] u_ca_in_72;
wire [17:0] u_ca_in_73;
wire [17:0] u_ca_in_74;
wire [17:0] u_ca_in_75;
wire [17:0] u_ca_in_76;
wire [17:0] u_ca_in_77;
wire [17:0] u_ca_in_78;
wire [17:0] u_ca_in_79;
wire [17:0] u_ca_in_80;
wire [17:0] u_ca_in_81;
wire [17:0] u_ca_in_82;
wire [17:0] u_ca_in_83;
wire [17:0] u_ca_in_84;
wire [17:0] u_ca_in_85;
wire [17:0] u_ca_in_86;
wire [17:0] u_ca_in_87;
wire [17:0] u_ca_in_88;
wire [17:0] u_ca_in_89;
wire [17:0] u_ca_in_90;
wire [17:0] u_ca_in_91;
wire [17:0] u_ca_in_92;
wire [17:0] u_ca_in_93;
wire [17:0] u_ca_in_94;
wire [17:0] u_ca_in_95;
wire [17:0] u_ca_in_96;
wire [17:0] u_ca_in_97;
wire [17:0] u_ca_in_98;
wire [17:0] u_ca_in_99;
wire [17:0] u_ca_in_100;
wire [17:0] u_ca_in_101;
wire [17:0] u_ca_in_102;
wire [17:0] u_ca_in_103;
wire [17:0] u_ca_in_104;
wire [17:0] u_ca_in_105;
wire [17:0] u_ca_in_106;
wire [17:0] u_ca_in_107;
wire [17:0] u_ca_in_108;
wire [17:0] u_ca_in_109;
wire [17:0] u_ca_in_110;
wire [17:0] u_ca_in_111;
wire [17:0] u_ca_in_112;
wire [17:0] u_ca_in_113;
wire [17:0] u_ca_in_114;
wire [17:0] u_ca_in_115;
wire [17:0] u_ca_in_116;
wire [17:0] u_ca_in_117;
wire [17:0] u_ca_in_118;
wire [17:0] u_ca_in_119;
wire [17:0] u_ca_in_120;
wire [17:0] u_ca_in_121;
wire [17:0] u_ca_in_122;
wire [17:0] u_ca_in_123;
wire [17:0] u_ca_in_124;
wire [17:0] u_ca_in_125;
wire [17:0] u_ca_in_126;
wire [17:0] u_ca_in_127;
wire [17:0] u_ca_in_128;
wire [17:0] u_ca_in_129;
wire [17:0] u_ca_in_130;
wire [17:0] u_ca_in_131;
wire [17:0] u_ca_in_132;
wire [17:0] u_ca_in_133;
wire [17:0] u_ca_in_134;
wire [17:0] u_ca_in_135;
wire [17:0] u_ca_in_136;
wire [17:0] u_ca_in_137;
wire [17:0] u_ca_in_138;
wire [17:0] u_ca_in_139;
wire [17:0] u_ca_in_140;
wire [17:0] u_ca_in_141;
wire [17:0] u_ca_in_142;
wire [17:0] u_ca_in_143;
wire [17:0] u_ca_in_144;
wire [17:0] u_ca_in_145;
wire [17:0] u_ca_in_146;
wire [17:0] u_ca_in_147;
wire [17:0] u_ca_in_148;
wire [17:0] u_ca_in_149;
wire [17:0] u_ca_in_150;
wire [17:0] u_ca_in_151;
wire [17:0] u_ca_in_152;
wire [17:0] u_ca_in_153;
wire [17:0] u_ca_in_154;
wire [17:0] u_ca_in_155;
wire [17:0] u_ca_in_156;
wire [17:0] u_ca_in_157;
wire [17:0] u_ca_in_158;
wire [17:0] u_ca_in_159;
wire [17:0] u_ca_in_160;
wire [17:0] u_ca_in_161;
wire [17:0] u_ca_in_162;
wire [17:0] u_ca_in_163;
wire [17:0] u_ca_in_164;
wire [17:0] u_ca_in_165;
wire [17:0] u_ca_in_166;
wire [17:0] u_ca_in_167;
wire [17:0] u_ca_in_168;
wire [17:0] u_ca_in_169;
wire [17:0] u_ca_in_170;
wire [17:0] u_ca_in_171;
wire [17:0] u_ca_in_172;
wire [17:0] u_ca_in_173;
wire [17:0] u_ca_in_174;
wire [17:0] u_ca_in_175;
wire [17:0] u_ca_in_176;
wire [17:0] u_ca_in_177;
wire [17:0] u_ca_in_178;
wire [17:0] u_ca_in_179;
wire [17:0] u_ca_in_180;
wire [17:0] u_ca_in_181;
wire [17:0] u_ca_in_182;
wire [17:0] u_ca_in_183;
wire [17:0] u_ca_in_184;
wire [17:0] u_ca_in_185;
wire [17:0] u_ca_in_186;
wire [17:0] u_ca_in_187;
wire [17:0] u_ca_in_188;
wire [17:0] u_ca_in_189;
wire [17:0] u_ca_in_190;
wire [17:0] u_ca_in_191;
wire [17:0] u_ca_in_192;
wire [17:0] u_ca_in_193;
wire [17:0] u_ca_in_194;
wire [17:0] u_ca_in_195;
wire [17:0] u_ca_in_196;
wire [17:0] u_ca_in_197;
wire [17:0] u_ca_in_198;
wire [17:0] u_ca_in_199;
wire [17:0] u_ca_in_200;
wire [17:0] u_ca_in_201;
wire [17:0] u_ca_in_202;
wire [17:0] u_ca_in_203;
wire [17:0] u_ca_in_204;
wire [17:0] u_ca_in_205;
wire [17:0] u_ca_in_206;
wire [17:0] u_ca_in_207;
wire [17:0] u_ca_in_208;
wire [17:0] u_ca_in_209;
wire [17:0] u_ca_in_210;
wire [17:0] u_ca_in_211;
wire [17:0] u_ca_in_212;
wire [17:0] u_ca_in_213;
wire [17:0] u_ca_in_214;
wire [17:0] u_ca_in_215;
wire [17:0] u_ca_in_216;
wire [17:0] u_ca_in_217;
wire [17:0] u_ca_in_218;
wire [17:0] u_ca_in_219;
wire [17:0] u_ca_in_220;
wire [17:0] u_ca_in_221;
wire [17:0] u_ca_in_222;
wire [17:0] u_ca_in_223;
wire [17:0] u_ca_in_224;
wire [17:0] u_ca_in_225;
wire [17:0] u_ca_in_226;
wire [17:0] u_ca_in_227;
wire [17:0] u_ca_in_228;
wire [17:0] u_ca_in_229;
wire [17:0] u_ca_in_230;
wire [17:0] u_ca_in_231;
wire [17:0] u_ca_in_232;
wire [17:0] u_ca_in_233;
wire [17:0] u_ca_in_234;
wire [17:0] u_ca_in_235;
wire [17:0] u_ca_in_236;
wire [17:0] u_ca_in_237;
wire [17:0] u_ca_in_238;
wire [17:0] u_ca_in_239;
wire [17:0] u_ca_in_240;
wire [17:0] u_ca_in_241;
wire [17:0] u_ca_in_242;
wire [17:0] u_ca_in_243;
wire [17:0] u_ca_in_244;
wire [17:0] u_ca_in_245;
wire [17:0] u_ca_in_246;
wire [17:0] u_ca_in_247;
wire [17:0] u_ca_in_248;
wire [17:0] u_ca_in_249;
wire [17:0] u_ca_in_250;
wire [17:0] u_ca_in_251;
wire [17:0] u_ca_in_252;
wire [17:0] u_ca_in_253;
wire [17:0] u_ca_in_254;
wire [17:0] u_ca_in_255;
wire [17:0] u_ca_in_256;
wire [17:0] u_ca_in_257;
wire [17:0] u_ca_in_258;
wire [17:0] u_ca_in_259;
wire [17:0] u_ca_in_260;
wire [17:0] u_ca_in_261;
wire [17:0] u_ca_in_262;
wire [17:0] u_ca_in_263;
wire [17:0] u_ca_in_264;
wire [17:0] u_ca_in_265;
wire [17:0] u_ca_in_266;
wire [17:0] u_ca_in_267;
wire [17:0] u_ca_in_268;
wire [17:0] u_ca_in_269;
wire [17:0] u_ca_in_270;
wire [17:0] u_ca_in_271;
wire [17:0] u_ca_in_272;
wire [17:0] u_ca_in_273;
wire [17:0] u_ca_in_274;
wire [17:0] u_ca_in_275;
wire [17:0] u_ca_in_276;
wire [17:0] u_ca_in_277;
wire [17:0] u_ca_in_278;
wire [17:0] u_ca_in_279;
wire [17:0] u_ca_in_280;
wire [17:0] u_ca_in_281;
wire [17:0] u_ca_in_282;
wire [17:0] u_ca_in_283;
wire [17:0] u_ca_in_284;
wire [17:0] u_ca_in_285;
wire [17:0] u_ca_in_286;
wire [17:0] u_ca_in_287;
wire [17:0] u_ca_in_288;
wire [17:0] u_ca_in_289;
wire [17:0] u_ca_in_290;
wire [17:0] u_ca_in_291;
wire [17:0] u_ca_in_292;
wire [17:0] u_ca_in_293;
wire [17:0] u_ca_in_294;
wire [17:0] u_ca_in_295;
wire [17:0] u_ca_in_296;
wire [17:0] u_ca_in_297;
wire [17:0] u_ca_in_298;
wire [17:0] u_ca_in_299;
wire [17:0] u_ca_in_300;
wire [17:0] u_ca_in_301;
wire [17:0] u_ca_in_302;
wire [17:0] u_ca_in_303;
wire [17:0] u_ca_in_304;
wire [17:0] u_ca_in_305;
wire [17:0] u_ca_in_306;
wire [17:0] u_ca_in_307;
wire [17:0] u_ca_in_308;
wire [17:0] u_ca_in_309;
wire [17:0] u_ca_in_310;
wire [17:0] u_ca_in_311;
wire [17:0] u_ca_in_312;
wire [17:0] u_ca_in_313;
wire [17:0] u_ca_in_314;
wire [17:0] u_ca_in_315;
wire [17:0] u_ca_in_316;
wire [17:0] u_ca_in_317;
wire [17:0] u_ca_in_318;
wire [17:0] u_ca_in_319;
wire [17:0] u_ca_in_320;
wire [17:0] u_ca_in_321;
wire [17:0] u_ca_in_322;
wire [17:0] u_ca_in_323;
wire [17:0] u_ca_in_324;
wire [17:0] u_ca_in_325;
wire [17:0] u_ca_in_326;
wire [17:0] u_ca_in_327;
wire [17:0] u_ca_in_328;
wire [17:0] u_ca_in_329;
wire [17:0] u_ca_in_330;
wire [17:0] u_ca_in_331;
wire [17:0] u_ca_in_332;
wire [17:0] u_ca_in_333;
wire [17:0] u_ca_in_334;
wire [17:0] u_ca_in_335;
wire [17:0] u_ca_in_336;
wire [17:0] u_ca_in_337;
wire [17:0] u_ca_in_338;
wire [17:0] u_ca_in_339;
wire [17:0] u_ca_in_340;
wire [17:0] u_ca_in_341;
wire [17:0] u_ca_in_342;
wire [17:0] u_ca_in_343;
wire [17:0] u_ca_in_344;
wire [17:0] u_ca_in_345;
wire [17:0] u_ca_in_346;
wire [17:0] u_ca_in_347;
wire [17:0] u_ca_in_348;
wire [17:0] u_ca_in_349;
wire [17:0] u_ca_in_350;
wire [17:0] u_ca_in_351;
wire [17:0] u_ca_in_352;
wire [17:0] u_ca_in_353;
wire [17:0] u_ca_in_354;
wire [17:0] u_ca_in_355;
wire [17:0] u_ca_in_356;
wire [17:0] u_ca_in_357;
wire [17:0] u_ca_in_358;
wire [17:0] u_ca_in_359;
wire [17:0] u_ca_in_360;
wire [17:0] u_ca_in_361;
wire [17:0] u_ca_in_362;
wire [17:0] u_ca_in_363;
wire [17:0] u_ca_in_364;
wire [17:0] u_ca_in_365;
wire [17:0] u_ca_in_366;
wire [17:0] u_ca_in_367;
wire [17:0] u_ca_in_368;
wire [17:0] u_ca_in_369;
wire [17:0] u_ca_in_370;
wire [17:0] u_ca_in_371;
wire [17:0] u_ca_in_372;
wire [17:0] u_ca_in_373;
wire [17:0] u_ca_in_374;
wire [17:0] u_ca_in_375;
wire [17:0] u_ca_in_376;
wire [17:0] u_ca_in_377;
wire [17:0] u_ca_in_378;
wire [17:0] u_ca_in_379;
wire [17:0] u_ca_in_380;
wire [17:0] u_ca_in_381;
wire [17:0] u_ca_in_382;
wire [17:0] u_ca_in_383;
wire [17:0] u_ca_in_384;
wire [17:0] u_ca_in_385;
wire [17:0] u_ca_in_386;
wire [17:0] u_ca_in_387;
wire [17:0] u_ca_in_388;
wire [17:0] u_ca_in_389;
wire [17:0] u_ca_in_390;
wire [17:0] u_ca_in_391;
wire [17:0] u_ca_in_392;
wire [17:0] u_ca_in_393;
wire [17:0] u_ca_in_394;
wire [17:0] u_ca_in_395;
wire [17:0] u_ca_in_396;
wire [17:0] u_ca_in_397;
wire [17:0] u_ca_in_398;
wire [17:0] u_ca_in_399;
wire [17:0] u_ca_in_400;
wire [17:0] u_ca_in_401;
wire [17:0] u_ca_in_402;
wire [17:0] u_ca_in_403;
wire [17:0] u_ca_in_404;
wire [17:0] u_ca_in_405;
wire [17:0] u_ca_in_406;
wire [17:0] u_ca_in_407;
wire [17:0] u_ca_in_408;
wire [17:0] u_ca_in_409;
wire [17:0] u_ca_in_410;
wire [17:0] u_ca_in_411;
wire [17:0] u_ca_in_412;
wire [17:0] u_ca_in_413;
wire [17:0] u_ca_in_414;
wire [17:0] u_ca_in_415;
wire [17:0] u_ca_in_416;
wire [17:0] u_ca_in_417;
wire [17:0] u_ca_in_418;
wire [17:0] u_ca_in_419;
wire [17:0] u_ca_in_420;
wire [17:0] u_ca_in_421;
wire [17:0] u_ca_in_422;
wire [17:0] u_ca_in_423;
wire [17:0] u_ca_in_424;
wire [17:0] u_ca_in_425;
wire [17:0] u_ca_in_426;
wire [17:0] u_ca_in_427;
wire [17:0] u_ca_in_428;
wire [17:0] u_ca_in_429;
wire [17:0] u_ca_in_430;
wire [17:0] u_ca_in_431;
wire [17:0] u_ca_in_432;
wire [17:0] u_ca_in_433;
wire [17:0] u_ca_in_434;
wire [17:0] u_ca_in_435;
wire [17:0] u_ca_in_436;
wire [17:0] u_ca_in_437;
wire [17:0] u_ca_in_438;
wire [17:0] u_ca_in_439;
wire [17:0] u_ca_in_440;
wire [17:0] u_ca_in_441;
wire [17:0] u_ca_in_442;
wire [17:0] u_ca_in_443;
wire [17:0] u_ca_in_444;
wire [17:0] u_ca_in_445;
wire [17:0] u_ca_in_446;
wire [17:0] u_ca_in_447;
wire [17:0] u_ca_in_448;
wire [17:0] u_ca_in_449;
wire [17:0] u_ca_in_450;
wire [17:0] u_ca_in_451;
wire [17:0] u_ca_in_452;
wire [17:0] u_ca_in_453;
wire [17:0] u_ca_in_454;
wire [17:0] u_ca_in_455;
wire [17:0] u_ca_in_456;
wire [17:0] u_ca_in_457;
wire [17:0] u_ca_in_458;
wire [17:0] u_ca_in_459;
wire [17:0] u_ca_in_460;
wire [17:0] u_ca_in_461;
wire [17:0] u_ca_in_462;
wire [17:0] u_ca_in_463;
wire [17:0] u_ca_in_464;
wire [17:0] u_ca_in_465;
wire [17:0] u_ca_in_466;
wire [17:0] u_ca_in_467;
wire [17:0] u_ca_in_468;
wire [17:0] u_ca_in_469;
wire [17:0] u_ca_in_470;
wire [17:0] u_ca_in_471;
wire [17:0] u_ca_in_472;
wire [17:0] u_ca_in_473;
wire [17:0] u_ca_in_474;
wire [17:0] u_ca_in_475;
wire [17:0] u_ca_in_476;
wire [17:0] u_ca_in_477;
wire [17:0] u_ca_in_478;
wire [17:0] u_ca_in_479;
wire [17:0] u_ca_in_480;
wire [17:0] u_ca_in_481;
wire [17:0] u_ca_in_482;
wire [17:0] u_ca_in_483;
wire [17:0] u_ca_in_484;
wire [17:0] u_ca_in_485;
wire [17:0] u_ca_in_486;
wire [17:0] u_ca_in_487;
wire [17:0] u_ca_in_488;
wire [17:0] u_ca_in_489;
wire [17:0] u_ca_in_490;
wire [17:0] u_ca_in_491;
wire [17:0] u_ca_in_492;
wire [17:0] u_ca_in_493;
wire [17:0] u_ca_in_494;
wire [17:0] u_ca_in_495;
wire [17:0] u_ca_in_496;
wire [17:0] u_ca_in_497;
wire [17:0] u_ca_in_498;
wire [17:0] u_ca_in_499;
wire [17:0] u_ca_in_500;
wire [17:0] u_ca_in_501;
wire [17:0] u_ca_in_502;
wire [17:0] u_ca_in_503;
wire [17:0] u_ca_in_504;
wire [17:0] u_ca_in_505;
wire [17:0] u_ca_in_506;
wire [17:0] u_ca_in_507;
wire [17:0] u_ca_in_508;
wire [17:0] u_ca_in_509;
wire [17:0] u_ca_in_510;
wire [17:0] u_ca_in_511;
wire [17:0] u_ca_in_512;
wire [17:0] u_ca_in_513;
wire [17:0] u_ca_in_514;
wire [17:0] u_ca_in_515;
wire [17:0] u_ca_in_516;
wire [17:0] u_ca_in_517;
wire [17:0] u_ca_in_518;
wire [17:0] u_ca_in_519;
wire [17:0] u_ca_in_520;
wire [17:0] u_ca_in_521;
wire [17:0] u_ca_in_522;
wire [17:0] u_ca_in_523;
wire [17:0] u_ca_in_524;
wire [17:0] u_ca_in_525;
wire [17:0] u_ca_in_526;
wire [17:0] u_ca_in_527;
wire [17:0] u_ca_in_528;
wire [17:0] u_ca_in_529;
wire [17:0] u_ca_in_530;
wire [17:0] u_ca_in_531;
wire [17:0] u_ca_in_532;
wire [17:0] u_ca_in_533;
wire [17:0] u_ca_in_534;
wire [17:0] u_ca_in_535;
wire [17:0] u_ca_in_536;
wire [17:0] u_ca_in_537;
wire [17:0] u_ca_in_538;
wire [17:0] u_ca_in_539;
wire [17:0] u_ca_in_540;
wire [17:0] u_ca_in_541;
wire [17:0] u_ca_in_542;
wire [17:0] u_ca_in_543;
wire [17:0] u_ca_in_544;
wire [17:0] u_ca_in_545;
wire [17:0] u_ca_in_546;
wire [17:0] u_ca_in_547;
wire [17:0] u_ca_in_548;
wire [17:0] u_ca_in_549;
wire [17:0] u_ca_in_550;
wire [17:0] u_ca_in_551;
wire [17:0] u_ca_in_552;
wire [17:0] u_ca_in_553;
wire [17:0] u_ca_in_554;
wire [17:0] u_ca_in_555;
wire [17:0] u_ca_in_556;
wire [17:0] u_ca_in_557;
wire [17:0] u_ca_in_558;
wire [17:0] u_ca_in_559;
wire [17:0] u_ca_in_560;
wire [17:0] u_ca_in_561;
wire [17:0] u_ca_in_562;
wire [17:0] u_ca_in_563;
wire [17:0] u_ca_in_564;
wire [17:0] u_ca_in_565;
wire [17:0] u_ca_in_566;
wire [17:0] u_ca_in_567;
wire [17:0] u_ca_in_568;
wire [17:0] u_ca_in_569;
wire [17:0] u_ca_in_570;
wire [17:0] u_ca_in_571;
wire [17:0] u_ca_in_572;
wire [17:0] u_ca_in_573;
wire [17:0] u_ca_in_574;
wire [17:0] u_ca_in_575;
wire [17:0] u_ca_in_576;
wire [17:0] u_ca_in_577;
wire [17:0] u_ca_in_578;
wire [17:0] u_ca_in_579;
wire [17:0] u_ca_in_580;
wire [17:0] u_ca_in_581;
wire [17:0] u_ca_in_582;
wire [17:0] u_ca_in_583;
wire [17:0] u_ca_in_584;
wire [17:0] u_ca_in_585;
wire [17:0] u_ca_in_586;
wire [17:0] u_ca_in_587;
wire [17:0] u_ca_in_588;
wire [17:0] u_ca_in_589;
wire [17:0] u_ca_in_590;
wire [17:0] u_ca_in_591;
wire [17:0] u_ca_in_592;
wire [17:0] u_ca_in_593;
wire [17:0] u_ca_in_594;
wire [17:0] u_ca_in_595;
wire [17:0] u_ca_in_596;
wire [17:0] u_ca_in_597;
wire [17:0] u_ca_in_598;
wire [17:0] u_ca_in_599;
wire [17:0] u_ca_in_600;
wire [17:0] u_ca_in_601;
wire [17:0] u_ca_in_602;
wire [17:0] u_ca_in_603;
wire [17:0] u_ca_in_604;
wire [17:0] u_ca_in_605;
wire [17:0] u_ca_in_606;
wire [17:0] u_ca_in_607;
wire [17:0] u_ca_in_608;
wire [17:0] u_ca_in_609;
wire [17:0] u_ca_in_610;
wire [17:0] u_ca_in_611;
wire [17:0] u_ca_in_612;
wire [17:0] u_ca_in_613;
wire [17:0] u_ca_in_614;
wire [17:0] u_ca_in_615;
wire [17:0] u_ca_in_616;
wire [17:0] u_ca_in_617;
wire [17:0] u_ca_in_618;
wire [17:0] u_ca_in_619;
wire [17:0] u_ca_in_620;
wire [17:0] u_ca_in_621;
wire [17:0] u_ca_in_622;
wire [17:0] u_ca_in_623;
wire [17:0] u_ca_in_624;
wire [17:0] u_ca_in_625;
wire [17:0] u_ca_in_626;
wire [17:0] u_ca_in_627;
wire [17:0] u_ca_in_628;
wire [17:0] u_ca_in_629;
wire [17:0] u_ca_in_630;
wire [17:0] u_ca_in_631;
wire [17:0] u_ca_in_632;
wire [17:0] u_ca_in_633;
wire [17:0] u_ca_in_634;
wire [17:0] u_ca_in_635;
wire [17:0] u_ca_in_636;
wire [17:0] u_ca_in_637;
wire [17:0] u_ca_in_638;
wire [17:0] u_ca_in_639;
wire [17:0] u_ca_in_640;
wire [17:0] u_ca_in_641;
wire [17:0] u_ca_in_642;
wire [17:0] u_ca_in_643;
wire [17:0] u_ca_in_644;
wire [17:0] u_ca_in_645;
wire [17:0] u_ca_in_646;
wire [17:0] u_ca_in_647;
wire [17:0] u_ca_in_648;
wire [17:0] u_ca_in_649;
wire [17:0] u_ca_in_650;
wire [17:0] u_ca_in_651;
wire [17:0] u_ca_in_652;
wire [17:0] u_ca_in_653;
wire [17:0] u_ca_in_654;
wire [17:0] u_ca_in_655;
wire [17:0] u_ca_in_656;
wire [17:0] u_ca_in_657;
wire [17:0] u_ca_in_658;
wire [17:0] u_ca_in_659;
wire [17:0] u_ca_in_660;
wire [17:0] u_ca_in_661;
wire [17:0] u_ca_in_662;
wire [17:0] u_ca_in_663;
wire [17:0] u_ca_in_664;
wire [17:0] u_ca_in_665;
wire [17:0] u_ca_in_666;
wire [17:0] u_ca_in_667;
wire [17:0] u_ca_in_668;
wire [17:0] u_ca_in_669;
wire [17:0] u_ca_in_670;
wire [17:0] u_ca_in_671;
wire [17:0] u_ca_in_672;
wire [17:0] u_ca_in_673;
wire [17:0] u_ca_in_674;
wire [17:0] u_ca_in_675;
wire [17:0] u_ca_in_676;
wire [17:0] u_ca_in_677;
wire [17:0] u_ca_in_678;
wire [17:0] u_ca_in_679;
wire [17:0] u_ca_in_680;
wire [17:0] u_ca_in_681;
wire [17:0] u_ca_in_682;
wire [17:0] u_ca_in_683;
wire [17:0] u_ca_in_684;
wire [17:0] u_ca_in_685;
wire [17:0] u_ca_in_686;
wire [17:0] u_ca_in_687;
wire [17:0] u_ca_in_688;
wire [17:0] u_ca_in_689;
wire [17:0] u_ca_in_690;
wire [17:0] u_ca_in_691;
wire [17:0] u_ca_in_692;
wire [17:0] u_ca_in_693;
wire [17:0] u_ca_in_694;
wire [17:0] u_ca_in_695;
wire [17:0] u_ca_in_696;
wire [17:0] u_ca_in_697;
wire [17:0] u_ca_in_698;
wire [17:0] u_ca_in_699;
wire [17:0] u_ca_in_700;
wire [17:0] u_ca_in_701;
wire [17:0] u_ca_in_702;
wire [17:0] u_ca_in_703;
wire [17:0] u_ca_in_704;
wire [17:0] u_ca_in_705;
wire [17:0] u_ca_in_706;
wire [17:0] u_ca_in_707;
wire [17:0] u_ca_in_708;
wire [17:0] u_ca_in_709;
wire [17:0] u_ca_in_710;
wire [17:0] u_ca_in_711;
wire [17:0] u_ca_in_712;
wire [17:0] u_ca_in_713;
wire [17:0] u_ca_in_714;
wire [17:0] u_ca_in_715;
wire [17:0] u_ca_in_716;
wire [17:0] u_ca_in_717;
wire [17:0] u_ca_in_718;
wire [17:0] u_ca_in_719;
wire [17:0] u_ca_in_720;
wire [17:0] u_ca_in_721;
wire [17:0] u_ca_in_722;
wire [17:0] u_ca_in_723;
wire [17:0] u_ca_in_724;
wire [17:0] u_ca_in_725;
wire [17:0] u_ca_in_726;
wire [17:0] u_ca_in_727;
wire [17:0] u_ca_in_728;
wire [17:0] u_ca_in_729;
wire [17:0] u_ca_in_730;
wire [17:0] u_ca_in_731;
wire [17:0] u_ca_in_732;
wire [17:0] u_ca_in_733;
wire [17:0] u_ca_in_734;
wire [17:0] u_ca_in_735;
wire [17:0] u_ca_in_736;
wire [17:0] u_ca_in_737;
wire [17:0] u_ca_in_738;
wire [17:0] u_ca_in_739;
wire [17:0] u_ca_in_740;
wire [17:0] u_ca_in_741;
wire [17:0] u_ca_in_742;
wire [17:0] u_ca_in_743;
wire [17:0] u_ca_in_744;
wire [17:0] u_ca_in_745;
wire [17:0] u_ca_in_746;
wire [17:0] u_ca_in_747;
wire [17:0] u_ca_in_748;
wire [17:0] u_ca_in_749;
wire [17:0] u_ca_in_750;
wire [17:0] u_ca_in_751;
wire [17:0] u_ca_in_752;
wire [17:0] u_ca_in_753;
wire [17:0] u_ca_in_754;
wire [17:0] u_ca_in_755;
wire [17:0] u_ca_in_756;
wire [17:0] u_ca_in_757;
wire [17:0] u_ca_in_758;
wire [17:0] u_ca_in_759;
wire [17:0] u_ca_in_760;
wire [17:0] u_ca_in_761;
wire [17:0] u_ca_in_762;
wire [17:0] u_ca_in_763;
wire [17:0] u_ca_in_764;
wire [17:0] u_ca_in_765;
wire [17:0] u_ca_in_766;
wire [17:0] u_ca_in_767;
wire [17:0] u_ca_in_768;
wire [17:0] u_ca_in_769;
wire [17:0] u_ca_in_770;
wire [17:0] u_ca_in_771;
wire [17:0] u_ca_in_772;
wire [17:0] u_ca_in_773;
wire [17:0] u_ca_in_774;
wire [17:0] u_ca_in_775;
wire [17:0] u_ca_in_776;
wire [17:0] u_ca_in_777;
wire [17:0] u_ca_in_778;
wire [17:0] u_ca_in_779;
wire [17:0] u_ca_in_780;
wire [17:0] u_ca_in_781;
wire [17:0] u_ca_in_782;
wire [17:0] u_ca_in_783;
wire [17:0] u_ca_in_784;
wire [17:0] u_ca_in_785;
wire [17:0] u_ca_in_786;
wire [17:0] u_ca_in_787;
wire [17:0] u_ca_in_788;
wire [17:0] u_ca_in_789;
wire [17:0] u_ca_in_790;
wire [17:0] u_ca_in_791;
wire [17:0] u_ca_in_792;
wire [17:0] u_ca_in_793;
wire [17:0] u_ca_in_794;
wire [17:0] u_ca_in_795;
wire [17:0] u_ca_in_796;
wire [17:0] u_ca_in_797;
wire [17:0] u_ca_in_798;
wire [17:0] u_ca_in_799;
wire [17:0] u_ca_in_800;
wire [17:0] u_ca_in_801;
wire [17:0] u_ca_in_802;
wire [17:0] u_ca_in_803;
wire [17:0] u_ca_in_804;
wire [17:0] u_ca_in_805;
wire [17:0] u_ca_in_806;
wire [17:0] u_ca_in_807;
wire [17:0] u_ca_in_808;
wire [17:0] u_ca_in_809;
wire [17:0] u_ca_in_810;
wire [17:0] u_ca_in_811;
wire [17:0] u_ca_in_812;
wire [17:0] u_ca_in_813;
wire [17:0] u_ca_in_814;
wire [17:0] u_ca_in_815;
wire [17:0] u_ca_in_816;
wire [17:0] u_ca_in_817;
wire [17:0] u_ca_in_818;
wire [17:0] u_ca_in_819;
wire [17:0] u_ca_in_820;
wire [17:0] u_ca_in_821;
wire [17:0] u_ca_in_822;
wire [17:0] u_ca_in_823;
wire [17:0] u_ca_in_824;
wire [17:0] u_ca_in_825;
wire [17:0] u_ca_in_826;
wire [17:0] u_ca_in_827;
wire [17:0] u_ca_in_828;
wire [17:0] u_ca_in_829;
wire [17:0] u_ca_in_830;
wire [17:0] u_ca_in_831;
wire [17:0] u_ca_in_832;
wire [17:0] u_ca_in_833;
wire [17:0] u_ca_in_834;
wire [17:0] u_ca_in_835;
wire [17:0] u_ca_in_836;
wire [17:0] u_ca_in_837;
wire [17:0] u_ca_in_838;
wire [17:0] u_ca_in_839;
wire [17:0] u_ca_in_840;
wire [17:0] u_ca_in_841;
wire [17:0] u_ca_in_842;
wire [17:0] u_ca_in_843;
wire [17:0] u_ca_in_844;
wire [17:0] u_ca_in_845;
wire [17:0] u_ca_in_846;
wire [17:0] u_ca_in_847;
wire [17:0] u_ca_in_848;
wire [17:0] u_ca_in_849;
wire [17:0] u_ca_in_850;
wire [17:0] u_ca_in_851;
wire [17:0] u_ca_in_852;
wire [17:0] u_ca_in_853;
wire [17:0] u_ca_in_854;
wire [17:0] u_ca_in_855;
wire [17:0] u_ca_in_856;
wire [17:0] u_ca_in_857;
wire [17:0] u_ca_in_858;
wire [17:0] u_ca_in_859;
wire [17:0] u_ca_in_860;
wire [17:0] u_ca_in_861;
wire [17:0] u_ca_in_862;
wire [17:0] u_ca_in_863;
wire [17:0] u_ca_in_864;
wire [17:0] u_ca_in_865;
wire [17:0] u_ca_in_866;
wire [17:0] u_ca_in_867;
wire [17:0] u_ca_in_868;
wire [17:0] u_ca_in_869;
wire [17:0] u_ca_in_870;
wire [17:0] u_ca_in_871;
wire [17:0] u_ca_in_872;
wire [17:0] u_ca_in_873;
wire [17:0] u_ca_in_874;
wire [17:0] u_ca_in_875;
wire [17:0] u_ca_in_876;
wire [17:0] u_ca_in_877;
wire [17:0] u_ca_in_878;
wire [17:0] u_ca_in_879;
wire [17:0] u_ca_in_880;
wire [17:0] u_ca_in_881;
wire [17:0] u_ca_in_882;
wire [17:0] u_ca_in_883;
wire [17:0] u_ca_in_884;
wire [17:0] u_ca_in_885;
wire [17:0] u_ca_in_886;
wire [17:0] u_ca_in_887;
wire [17:0] u_ca_in_888;
wire [17:0] u_ca_in_889;
wire [17:0] u_ca_in_890;
wire [17:0] u_ca_in_891;
wire [17:0] u_ca_in_892;
wire [17:0] u_ca_in_893;
wire [17:0] u_ca_in_894;
wire [17:0] u_ca_in_895;
wire [17:0] u_ca_in_896;
wire [17:0] u_ca_in_897;
wire [17:0] u_ca_in_898;
wire [17:0] u_ca_in_899;
wire [17:0] u_ca_in_900;
wire [17:0] u_ca_in_901;
wire [17:0] u_ca_in_902;
wire [17:0] u_ca_in_903;
wire [17:0] u_ca_in_904;
wire [17:0] u_ca_in_905;
wire [17:0] u_ca_in_906;
wire [17:0] u_ca_in_907;
wire [17:0] u_ca_in_908;
wire [17:0] u_ca_in_909;
wire [17:0] u_ca_in_910;
wire [17:0] u_ca_in_911;
wire [17:0] u_ca_in_912;
wire [17:0] u_ca_in_913;
wire [17:0] u_ca_in_914;
wire [17:0] u_ca_in_915;
wire [17:0] u_ca_in_916;
wire [17:0] u_ca_in_917;
wire [17:0] u_ca_in_918;
wire [17:0] u_ca_in_919;
wire [17:0] u_ca_in_920;
wire [17:0] u_ca_in_921;
wire [17:0] u_ca_in_922;
wire [17:0] u_ca_in_923;
wire [17:0] u_ca_in_924;
wire [17:0] u_ca_in_925;
wire [17:0] u_ca_in_926;
wire [17:0] u_ca_in_927;
wire [17:0] u_ca_in_928;
wire [17:0] u_ca_in_929;
wire [17:0] u_ca_in_930;
wire [17:0] u_ca_in_931;
wire [17:0] u_ca_in_932;
wire [17:0] u_ca_in_933;
wire [17:0] u_ca_in_934;
wire [17:0] u_ca_in_935;
wire [17:0] u_ca_in_936;
wire [17:0] u_ca_in_937;
wire [17:0] u_ca_in_938;
wire [17:0] u_ca_in_939;
wire [17:0] u_ca_in_940;
wire [17:0] u_ca_in_941;
wire [17:0] u_ca_in_942;
wire [17:0] u_ca_in_943;
wire [17:0] u_ca_in_944;
wire [17:0] u_ca_in_945;
wire [17:0] u_ca_in_946;
wire [17:0] u_ca_in_947;
wire [17:0] u_ca_in_948;
wire [17:0] u_ca_in_949;
wire [17:0] u_ca_in_950;
wire [17:0] u_ca_in_951;
wire [17:0] u_ca_in_952;
wire [17:0] u_ca_in_953;
wire [17:0] u_ca_in_954;
wire [17:0] u_ca_in_955;
wire [17:0] u_ca_in_956;
wire [17:0] u_ca_in_957;
wire [17:0] u_ca_in_958;
wire [17:0] u_ca_in_959;
wire [17:0] u_ca_in_960;
wire [17:0] u_ca_in_961;
wire [17:0] u_ca_in_962;
wire [17:0] u_ca_in_963;
wire [17:0] u_ca_in_964;
wire [17:0] u_ca_in_965;
wire [17:0] u_ca_in_966;
wire [17:0] u_ca_in_967;
wire [17:0] u_ca_in_968;
wire [17:0] u_ca_in_969;
wire [17:0] u_ca_in_970;
wire [17:0] u_ca_in_971;
wire [17:0] u_ca_in_972;
wire [17:0] u_ca_in_973;
wire [17:0] u_ca_in_974;
wire [17:0] u_ca_in_975;
wire [17:0] u_ca_in_976;
wire [17:0] u_ca_in_977;
wire [17:0] u_ca_in_978;
wire [17:0] u_ca_in_979;
wire [17:0] u_ca_in_980;
wire [17:0] u_ca_in_981;
wire [17:0] u_ca_in_982;
wire [17:0] u_ca_in_983;
wire [17:0] u_ca_in_984;
wire [17:0] u_ca_in_985;
wire [17:0] u_ca_in_986;
wire [17:0] u_ca_in_987;
wire [17:0] u_ca_in_988;
wire [17:0] u_ca_in_989;
wire [17:0] u_ca_in_990;
wire [17:0] u_ca_in_991;
wire [17:0] u_ca_in_992;
wire [17:0] u_ca_in_993;
wire [17:0] u_ca_in_994;
wire [17:0] u_ca_in_995;
wire [17:0] u_ca_in_996;
wire [17:0] u_ca_in_997;
wire [17:0] u_ca_in_998;
wire [17:0] u_ca_in_999;
wire [17:0] u_ca_in_1000;
wire [17:0] u_ca_in_1001;
wire [17:0] u_ca_in_1002;
wire [17:0] u_ca_in_1003;
wire [17:0] u_ca_in_1004;
wire [17:0] u_ca_in_1005;
wire [17:0] u_ca_in_1006;
wire [17:0] u_ca_in_1007;
wire [17:0] u_ca_in_1008;
wire [17:0] u_ca_in_1009;
wire [17:0] u_ca_in_1010;
wire [17:0] u_ca_in_1011;
wire [17:0] u_ca_in_1012;
wire [17:0] u_ca_in_1013;
wire [17:0] u_ca_in_1014;
wire [17:0] u_ca_in_1015;
wire [17:0] u_ca_in_1016;
wire [17:0] u_ca_in_1017;
wire [17:0] u_ca_in_1018;
wire [17:0] u_ca_in_1019;
wire [17:0] u_ca_in_1020;
wire [17:0] u_ca_in_1021;
wire [17:0] u_ca_in_1022;
wire [17:0] u_ca_in_1023;
wire [17:0] u_ca_in_1024;
wire [17:0] u_ca_in_1025;
wire [17:0] u_ca_in_1026;
wire [17:0] u_ca_in_1027;
wire [17:0] u_ca_in_1028;
wire [17:0] u_ca_in_1029;
wire [17:0] u_ca_in_1030;
wire [17:0] u_ca_in_1031;
wire [17:0] u_ca_in_1032;
wire [11:0] u_ca_out_0;
wire [11:0] u_ca_out_1;
wire [11:0] u_ca_out_2;
wire [11:0] u_ca_out_3;
wire [11:0] u_ca_out_4;
wire [11:0] u_ca_out_5;
wire [11:0] u_ca_out_6;
wire [11:0] u_ca_out_7;
wire [11:0] u_ca_out_8;
wire [11:0] u_ca_out_9;
wire [11:0] u_ca_out_10;
wire [11:0] u_ca_out_11;
wire [11:0] u_ca_out_12;
wire [11:0] u_ca_out_13;
wire [11:0] u_ca_out_14;
wire [11:0] u_ca_out_15;
wire [11:0] u_ca_out_16;
wire [11:0] u_ca_out_17;
wire [11:0] u_ca_out_18;
wire [11:0] u_ca_out_19;
wire [11:0] u_ca_out_20;
wire [11:0] u_ca_out_21;
wire [11:0] u_ca_out_22;
wire [11:0] u_ca_out_23;
wire [11:0] u_ca_out_24;
wire [11:0] u_ca_out_25;
wire [11:0] u_ca_out_26;
wire [11:0] u_ca_out_27;
wire [11:0] u_ca_out_28;
wire [11:0] u_ca_out_29;
wire [11:0] u_ca_out_30;
wire [11:0] u_ca_out_31;
wire [11:0] u_ca_out_32;
wire [11:0] u_ca_out_33;
wire [11:0] u_ca_out_34;
wire [11:0] u_ca_out_35;
wire [11:0] u_ca_out_36;
wire [11:0] u_ca_out_37;
wire [11:0] u_ca_out_38;
wire [11:0] u_ca_out_39;
wire [11:0] u_ca_out_40;
wire [11:0] u_ca_out_41;
wire [11:0] u_ca_out_42;
wire [11:0] u_ca_out_43;
wire [11:0] u_ca_out_44;
wire [11:0] u_ca_out_45;
wire [11:0] u_ca_out_46;
wire [11:0] u_ca_out_47;
wire [11:0] u_ca_out_48;
wire [11:0] u_ca_out_49;
wire [11:0] u_ca_out_50;
wire [11:0] u_ca_out_51;
wire [11:0] u_ca_out_52;
wire [11:0] u_ca_out_53;
wire [11:0] u_ca_out_54;
wire [11:0] u_ca_out_55;
wire [11:0] u_ca_out_56;
wire [11:0] u_ca_out_57;
wire [11:0] u_ca_out_58;
wire [11:0] u_ca_out_59;
wire [11:0] u_ca_out_60;
wire [11:0] u_ca_out_61;
wire [11:0] u_ca_out_62;
wire [11:0] u_ca_out_63;
wire [11:0] u_ca_out_64;
wire [11:0] u_ca_out_65;
wire [11:0] u_ca_out_66;
wire [11:0] u_ca_out_67;
wire [11:0] u_ca_out_68;
wire [11:0] u_ca_out_69;
wire [11:0] u_ca_out_70;
wire [11:0] u_ca_out_71;
wire [11:0] u_ca_out_72;
wire [11:0] u_ca_out_73;
wire [11:0] u_ca_out_74;
wire [11:0] u_ca_out_75;
wire [11:0] u_ca_out_76;
wire [11:0] u_ca_out_77;
wire [11:0] u_ca_out_78;
wire [11:0] u_ca_out_79;
wire [11:0] u_ca_out_80;
wire [11:0] u_ca_out_81;
wire [11:0] u_ca_out_82;
wire [11:0] u_ca_out_83;
wire [11:0] u_ca_out_84;
wire [11:0] u_ca_out_85;
wire [11:0] u_ca_out_86;
wire [11:0] u_ca_out_87;
wire [11:0] u_ca_out_88;
wire [11:0] u_ca_out_89;
wire [11:0] u_ca_out_90;
wire [11:0] u_ca_out_91;
wire [11:0] u_ca_out_92;
wire [11:0] u_ca_out_93;
wire [11:0] u_ca_out_94;
wire [11:0] u_ca_out_95;
wire [11:0] u_ca_out_96;
wire [11:0] u_ca_out_97;
wire [11:0] u_ca_out_98;
wire [11:0] u_ca_out_99;
wire [11:0] u_ca_out_100;
wire [11:0] u_ca_out_101;
wire [11:0] u_ca_out_102;
wire [11:0] u_ca_out_103;
wire [11:0] u_ca_out_104;
wire [11:0] u_ca_out_105;
wire [11:0] u_ca_out_106;
wire [11:0] u_ca_out_107;
wire [11:0] u_ca_out_108;
wire [11:0] u_ca_out_109;
wire [11:0] u_ca_out_110;
wire [11:0] u_ca_out_111;
wire [11:0] u_ca_out_112;
wire [11:0] u_ca_out_113;
wire [11:0] u_ca_out_114;
wire [11:0] u_ca_out_115;
wire [11:0] u_ca_out_116;
wire [11:0] u_ca_out_117;
wire [11:0] u_ca_out_118;
wire [11:0] u_ca_out_119;
wire [11:0] u_ca_out_120;
wire [11:0] u_ca_out_121;
wire [11:0] u_ca_out_122;
wire [11:0] u_ca_out_123;
wire [11:0] u_ca_out_124;
wire [11:0] u_ca_out_125;
wire [11:0] u_ca_out_126;
wire [11:0] u_ca_out_127;
wire [11:0] u_ca_out_128;
wire [11:0] u_ca_out_129;
wire [11:0] u_ca_out_130;
wire [11:0] u_ca_out_131;
wire [11:0] u_ca_out_132;
wire [11:0] u_ca_out_133;
wire [11:0] u_ca_out_134;
wire [11:0] u_ca_out_135;
wire [11:0] u_ca_out_136;
wire [11:0] u_ca_out_137;
wire [11:0] u_ca_out_138;
wire [11:0] u_ca_out_139;
wire [11:0] u_ca_out_140;
wire [11:0] u_ca_out_141;
wire [11:0] u_ca_out_142;
wire [11:0] u_ca_out_143;
wire [11:0] u_ca_out_144;
wire [11:0] u_ca_out_145;
wire [11:0] u_ca_out_146;
wire [11:0] u_ca_out_147;
wire [11:0] u_ca_out_148;
wire [11:0] u_ca_out_149;
wire [11:0] u_ca_out_150;
wire [11:0] u_ca_out_151;
wire [11:0] u_ca_out_152;
wire [11:0] u_ca_out_153;
wire [11:0] u_ca_out_154;
wire [11:0] u_ca_out_155;
wire [11:0] u_ca_out_156;
wire [11:0] u_ca_out_157;
wire [11:0] u_ca_out_158;
wire [11:0] u_ca_out_159;
wire [11:0] u_ca_out_160;
wire [11:0] u_ca_out_161;
wire [11:0] u_ca_out_162;
wire [11:0] u_ca_out_163;
wire [11:0] u_ca_out_164;
wire [11:0] u_ca_out_165;
wire [11:0] u_ca_out_166;
wire [11:0] u_ca_out_167;
wire [11:0] u_ca_out_168;
wire [11:0] u_ca_out_169;
wire [11:0] u_ca_out_170;
wire [11:0] u_ca_out_171;
wire [11:0] u_ca_out_172;
wire [11:0] u_ca_out_173;
wire [11:0] u_ca_out_174;
wire [11:0] u_ca_out_175;
wire [11:0] u_ca_out_176;
wire [11:0] u_ca_out_177;
wire [11:0] u_ca_out_178;
wire [11:0] u_ca_out_179;
wire [11:0] u_ca_out_180;
wire [11:0] u_ca_out_181;
wire [11:0] u_ca_out_182;
wire [11:0] u_ca_out_183;
wire [11:0] u_ca_out_184;
wire [11:0] u_ca_out_185;
wire [11:0] u_ca_out_186;
wire [11:0] u_ca_out_187;
wire [11:0] u_ca_out_188;
wire [11:0] u_ca_out_189;
wire [11:0] u_ca_out_190;
wire [11:0] u_ca_out_191;
wire [11:0] u_ca_out_192;
wire [11:0] u_ca_out_193;
wire [11:0] u_ca_out_194;
wire [11:0] u_ca_out_195;
wire [11:0] u_ca_out_196;
wire [11:0] u_ca_out_197;
wire [11:0] u_ca_out_198;
wire [11:0] u_ca_out_199;
wire [11:0] u_ca_out_200;
wire [11:0] u_ca_out_201;
wire [11:0] u_ca_out_202;
wire [11:0] u_ca_out_203;
wire [11:0] u_ca_out_204;
wire [11:0] u_ca_out_205;
wire [11:0] u_ca_out_206;
wire [11:0] u_ca_out_207;
wire [11:0] u_ca_out_208;
wire [11:0] u_ca_out_209;
wire [11:0] u_ca_out_210;
wire [11:0] u_ca_out_211;
wire [11:0] u_ca_out_212;
wire [11:0] u_ca_out_213;
wire [11:0] u_ca_out_214;
wire [11:0] u_ca_out_215;
wire [11:0] u_ca_out_216;
wire [11:0] u_ca_out_217;
wire [11:0] u_ca_out_218;
wire [11:0] u_ca_out_219;
wire [11:0] u_ca_out_220;
wire [11:0] u_ca_out_221;
wire [11:0] u_ca_out_222;
wire [11:0] u_ca_out_223;
wire [11:0] u_ca_out_224;
wire [11:0] u_ca_out_225;
wire [11:0] u_ca_out_226;
wire [11:0] u_ca_out_227;
wire [11:0] u_ca_out_228;
wire [11:0] u_ca_out_229;
wire [11:0] u_ca_out_230;
wire [11:0] u_ca_out_231;
wire [11:0] u_ca_out_232;
wire [11:0] u_ca_out_233;
wire [11:0] u_ca_out_234;
wire [11:0] u_ca_out_235;
wire [11:0] u_ca_out_236;
wire [11:0] u_ca_out_237;
wire [11:0] u_ca_out_238;
wire [11:0] u_ca_out_239;
wire [11:0] u_ca_out_240;
wire [11:0] u_ca_out_241;
wire [11:0] u_ca_out_242;
wire [11:0] u_ca_out_243;
wire [11:0] u_ca_out_244;
wire [11:0] u_ca_out_245;
wire [11:0] u_ca_out_246;
wire [11:0] u_ca_out_247;
wire [11:0] u_ca_out_248;
wire [11:0] u_ca_out_249;
wire [11:0] u_ca_out_250;
wire [11:0] u_ca_out_251;
wire [11:0] u_ca_out_252;
wire [11:0] u_ca_out_253;
wire [11:0] u_ca_out_254;
wire [11:0] u_ca_out_255;
wire [11:0] u_ca_out_256;
wire [11:0] u_ca_out_257;
wire [11:0] u_ca_out_258;
wire [11:0] u_ca_out_259;
wire [11:0] u_ca_out_260;
wire [11:0] u_ca_out_261;
wire [11:0] u_ca_out_262;
wire [11:0] u_ca_out_263;
wire [11:0] u_ca_out_264;
wire [11:0] u_ca_out_265;
wire [11:0] u_ca_out_266;
wire [11:0] u_ca_out_267;
wire [11:0] u_ca_out_268;
wire [11:0] u_ca_out_269;
wire [11:0] u_ca_out_270;
wire [11:0] u_ca_out_271;
wire [11:0] u_ca_out_272;
wire [11:0] u_ca_out_273;
wire [11:0] u_ca_out_274;
wire [11:0] u_ca_out_275;
wire [11:0] u_ca_out_276;
wire [11:0] u_ca_out_277;
wire [11:0] u_ca_out_278;
wire [11:0] u_ca_out_279;
wire [11:0] u_ca_out_280;
wire [11:0] u_ca_out_281;
wire [11:0] u_ca_out_282;
wire [11:0] u_ca_out_283;
wire [11:0] u_ca_out_284;
wire [11:0] u_ca_out_285;
wire [11:0] u_ca_out_286;
wire [11:0] u_ca_out_287;
wire [11:0] u_ca_out_288;
wire [11:0] u_ca_out_289;
wire [11:0] u_ca_out_290;
wire [11:0] u_ca_out_291;
wire [11:0] u_ca_out_292;
wire [11:0] u_ca_out_293;
wire [11:0] u_ca_out_294;
wire [11:0] u_ca_out_295;
wire [11:0] u_ca_out_296;
wire [11:0] u_ca_out_297;
wire [11:0] u_ca_out_298;
wire [11:0] u_ca_out_299;
wire [11:0] u_ca_out_300;
wire [11:0] u_ca_out_301;
wire [11:0] u_ca_out_302;
wire [11:0] u_ca_out_303;
wire [11:0] u_ca_out_304;
wire [11:0] u_ca_out_305;
wire [11:0] u_ca_out_306;
wire [11:0] u_ca_out_307;
wire [11:0] u_ca_out_308;
wire [11:0] u_ca_out_309;
wire [11:0] u_ca_out_310;
wire [11:0] u_ca_out_311;
wire [11:0] u_ca_out_312;
wire [11:0] u_ca_out_313;
wire [11:0] u_ca_out_314;
wire [11:0] u_ca_out_315;
wire [11:0] u_ca_out_316;
wire [11:0] u_ca_out_317;
wire [11:0] u_ca_out_318;
wire [11:0] u_ca_out_319;
wire [11:0] u_ca_out_320;
wire [11:0] u_ca_out_321;
wire [11:0] u_ca_out_322;
wire [11:0] u_ca_out_323;
wire [11:0] u_ca_out_324;
wire [11:0] u_ca_out_325;
wire [11:0] u_ca_out_326;
wire [11:0] u_ca_out_327;
wire [11:0] u_ca_out_328;
wire [11:0] u_ca_out_329;
wire [11:0] u_ca_out_330;
wire [11:0] u_ca_out_331;
wire [11:0] u_ca_out_332;
wire [11:0] u_ca_out_333;
wire [11:0] u_ca_out_334;
wire [11:0] u_ca_out_335;
wire [11:0] u_ca_out_336;
wire [11:0] u_ca_out_337;
wire [11:0] u_ca_out_338;
wire [11:0] u_ca_out_339;
wire [11:0] u_ca_out_340;
wire [11:0] u_ca_out_341;
wire [11:0] u_ca_out_342;
wire [11:0] u_ca_out_343;
wire [11:0] u_ca_out_344;
wire [11:0] u_ca_out_345;
wire [11:0] u_ca_out_346;
wire [11:0] u_ca_out_347;
wire [11:0] u_ca_out_348;
wire [11:0] u_ca_out_349;
wire [11:0] u_ca_out_350;
wire [11:0] u_ca_out_351;
wire [11:0] u_ca_out_352;
wire [11:0] u_ca_out_353;
wire [11:0] u_ca_out_354;
wire [11:0] u_ca_out_355;
wire [11:0] u_ca_out_356;
wire [11:0] u_ca_out_357;
wire [11:0] u_ca_out_358;
wire [11:0] u_ca_out_359;
wire [11:0] u_ca_out_360;
wire [11:0] u_ca_out_361;
wire [11:0] u_ca_out_362;
wire [11:0] u_ca_out_363;
wire [11:0] u_ca_out_364;
wire [11:0] u_ca_out_365;
wire [11:0] u_ca_out_366;
wire [11:0] u_ca_out_367;
wire [11:0] u_ca_out_368;
wire [11:0] u_ca_out_369;
wire [11:0] u_ca_out_370;
wire [11:0] u_ca_out_371;
wire [11:0] u_ca_out_372;
wire [11:0] u_ca_out_373;
wire [11:0] u_ca_out_374;
wire [11:0] u_ca_out_375;
wire [11:0] u_ca_out_376;
wire [11:0] u_ca_out_377;
wire [11:0] u_ca_out_378;
wire [11:0] u_ca_out_379;
wire [11:0] u_ca_out_380;
wire [11:0] u_ca_out_381;
wire [11:0] u_ca_out_382;
wire [11:0] u_ca_out_383;
wire [11:0] u_ca_out_384;
wire [11:0] u_ca_out_385;
wire [11:0] u_ca_out_386;
wire [11:0] u_ca_out_387;
wire [11:0] u_ca_out_388;
wire [11:0] u_ca_out_389;
wire [11:0] u_ca_out_390;
wire [11:0] u_ca_out_391;
wire [11:0] u_ca_out_392;
wire [11:0] u_ca_out_393;
wire [11:0] u_ca_out_394;
wire [11:0] u_ca_out_395;
wire [11:0] u_ca_out_396;
wire [11:0] u_ca_out_397;
wire [11:0] u_ca_out_398;
wire [11:0] u_ca_out_399;
wire [11:0] u_ca_out_400;
wire [11:0] u_ca_out_401;
wire [11:0] u_ca_out_402;
wire [11:0] u_ca_out_403;
wire [11:0] u_ca_out_404;
wire [11:0] u_ca_out_405;
wire [11:0] u_ca_out_406;
wire [11:0] u_ca_out_407;
wire [11:0] u_ca_out_408;
wire [11:0] u_ca_out_409;
wire [11:0] u_ca_out_410;
wire [11:0] u_ca_out_411;
wire [11:0] u_ca_out_412;
wire [11:0] u_ca_out_413;
wire [11:0] u_ca_out_414;
wire [11:0] u_ca_out_415;
wire [11:0] u_ca_out_416;
wire [11:0] u_ca_out_417;
wire [11:0] u_ca_out_418;
wire [11:0] u_ca_out_419;
wire [11:0] u_ca_out_420;
wire [11:0] u_ca_out_421;
wire [11:0] u_ca_out_422;
wire [11:0] u_ca_out_423;
wire [11:0] u_ca_out_424;
wire [11:0] u_ca_out_425;
wire [11:0] u_ca_out_426;
wire [11:0] u_ca_out_427;
wire [11:0] u_ca_out_428;
wire [11:0] u_ca_out_429;
wire [11:0] u_ca_out_430;
wire [11:0] u_ca_out_431;
wire [11:0] u_ca_out_432;
wire [11:0] u_ca_out_433;
wire [11:0] u_ca_out_434;
wire [11:0] u_ca_out_435;
wire [11:0] u_ca_out_436;
wire [11:0] u_ca_out_437;
wire [11:0] u_ca_out_438;
wire [11:0] u_ca_out_439;
wire [11:0] u_ca_out_440;
wire [11:0] u_ca_out_441;
wire [11:0] u_ca_out_442;
wire [11:0] u_ca_out_443;
wire [11:0] u_ca_out_444;
wire [11:0] u_ca_out_445;
wire [11:0] u_ca_out_446;
wire [11:0] u_ca_out_447;
wire [11:0] u_ca_out_448;
wire [11:0] u_ca_out_449;
wire [11:0] u_ca_out_450;
wire [11:0] u_ca_out_451;
wire [11:0] u_ca_out_452;
wire [11:0] u_ca_out_453;
wire [11:0] u_ca_out_454;
wire [11:0] u_ca_out_455;
wire [11:0] u_ca_out_456;
wire [11:0] u_ca_out_457;
wire [11:0] u_ca_out_458;
wire [11:0] u_ca_out_459;
wire [11:0] u_ca_out_460;
wire [11:0] u_ca_out_461;
wire [11:0] u_ca_out_462;
wire [11:0] u_ca_out_463;
wire [11:0] u_ca_out_464;
wire [11:0] u_ca_out_465;
wire [11:0] u_ca_out_466;
wire [11:0] u_ca_out_467;
wire [11:0] u_ca_out_468;
wire [11:0] u_ca_out_469;
wire [11:0] u_ca_out_470;
wire [11:0] u_ca_out_471;
wire [11:0] u_ca_out_472;
wire [11:0] u_ca_out_473;
wire [11:0] u_ca_out_474;
wire [11:0] u_ca_out_475;
wire [11:0] u_ca_out_476;
wire [11:0] u_ca_out_477;
wire [11:0] u_ca_out_478;
wire [11:0] u_ca_out_479;
wire [11:0] u_ca_out_480;
wire [11:0] u_ca_out_481;
wire [11:0] u_ca_out_482;
wire [11:0] u_ca_out_483;
wire [11:0] u_ca_out_484;
wire [11:0] u_ca_out_485;
wire [11:0] u_ca_out_486;
wire [11:0] u_ca_out_487;
wire [11:0] u_ca_out_488;
wire [11:0] u_ca_out_489;
wire [11:0] u_ca_out_490;
wire [11:0] u_ca_out_491;
wire [11:0] u_ca_out_492;
wire [11:0] u_ca_out_493;
wire [11:0] u_ca_out_494;
wire [11:0] u_ca_out_495;
wire [11:0] u_ca_out_496;
wire [11:0] u_ca_out_497;
wire [11:0] u_ca_out_498;
wire [11:0] u_ca_out_499;
wire [11:0] u_ca_out_500;
wire [11:0] u_ca_out_501;
wire [11:0] u_ca_out_502;
wire [11:0] u_ca_out_503;
wire [11:0] u_ca_out_504;
wire [11:0] u_ca_out_505;
wire [11:0] u_ca_out_506;
wire [11:0] u_ca_out_507;
wire [11:0] u_ca_out_508;
wire [11:0] u_ca_out_509;
wire [11:0] u_ca_out_510;
wire [11:0] u_ca_out_511;
wire [11:0] u_ca_out_512;
wire [11:0] u_ca_out_513;
wire [11:0] u_ca_out_514;
wire [11:0] u_ca_out_515;
wire [11:0] u_ca_out_516;
wire [11:0] u_ca_out_517;
wire [11:0] u_ca_out_518;
wire [11:0] u_ca_out_519;
wire [11:0] u_ca_out_520;
wire [11:0] u_ca_out_521;
wire [11:0] u_ca_out_522;
wire [11:0] u_ca_out_523;
wire [11:0] u_ca_out_524;
wire [11:0] u_ca_out_525;
wire [11:0] u_ca_out_526;
wire [11:0] u_ca_out_527;
wire [11:0] u_ca_out_528;
wire [11:0] u_ca_out_529;
wire [11:0] u_ca_out_530;
wire [11:0] u_ca_out_531;
wire [11:0] u_ca_out_532;
wire [11:0] u_ca_out_533;
wire [11:0] u_ca_out_534;
wire [11:0] u_ca_out_535;
wire [11:0] u_ca_out_536;
wire [11:0] u_ca_out_537;
wire [11:0] u_ca_out_538;
wire [11:0] u_ca_out_539;
wire [11:0] u_ca_out_540;
wire [11:0] u_ca_out_541;
wire [11:0] u_ca_out_542;
wire [11:0] u_ca_out_543;
wire [11:0] u_ca_out_544;
wire [11:0] u_ca_out_545;
wire [11:0] u_ca_out_546;
wire [11:0] u_ca_out_547;
wire [11:0] u_ca_out_548;
wire [11:0] u_ca_out_549;
wire [11:0] u_ca_out_550;
wire [11:0] u_ca_out_551;
wire [11:0] u_ca_out_552;
wire [11:0] u_ca_out_553;
wire [11:0] u_ca_out_554;
wire [11:0] u_ca_out_555;
wire [11:0] u_ca_out_556;
wire [11:0] u_ca_out_557;
wire [11:0] u_ca_out_558;
wire [11:0] u_ca_out_559;
wire [11:0] u_ca_out_560;
wire [11:0] u_ca_out_561;
wire [11:0] u_ca_out_562;
wire [11:0] u_ca_out_563;
wire [11:0] u_ca_out_564;
wire [11:0] u_ca_out_565;
wire [11:0] u_ca_out_566;
wire [11:0] u_ca_out_567;
wire [11:0] u_ca_out_568;
wire [11:0] u_ca_out_569;
wire [11:0] u_ca_out_570;
wire [11:0] u_ca_out_571;
wire [11:0] u_ca_out_572;
wire [11:0] u_ca_out_573;
wire [11:0] u_ca_out_574;
wire [11:0] u_ca_out_575;
wire [11:0] u_ca_out_576;
wire [11:0] u_ca_out_577;
wire [11:0] u_ca_out_578;
wire [11:0] u_ca_out_579;
wire [11:0] u_ca_out_580;
wire [11:0] u_ca_out_581;
wire [11:0] u_ca_out_582;
wire [11:0] u_ca_out_583;
wire [11:0] u_ca_out_584;
wire [11:0] u_ca_out_585;
wire [11:0] u_ca_out_586;
wire [11:0] u_ca_out_587;
wire [11:0] u_ca_out_588;
wire [11:0] u_ca_out_589;
wire [11:0] u_ca_out_590;
wire [11:0] u_ca_out_591;
wire [11:0] u_ca_out_592;
wire [11:0] u_ca_out_593;
wire [11:0] u_ca_out_594;
wire [11:0] u_ca_out_595;
wire [11:0] u_ca_out_596;
wire [11:0] u_ca_out_597;
wire [11:0] u_ca_out_598;
wire [11:0] u_ca_out_599;
wire [11:0] u_ca_out_600;
wire [11:0] u_ca_out_601;
wire [11:0] u_ca_out_602;
wire [11:0] u_ca_out_603;
wire [11:0] u_ca_out_604;
wire [11:0] u_ca_out_605;
wire [11:0] u_ca_out_606;
wire [11:0] u_ca_out_607;
wire [11:0] u_ca_out_608;
wire [11:0] u_ca_out_609;
wire [11:0] u_ca_out_610;
wire [11:0] u_ca_out_611;
wire [11:0] u_ca_out_612;
wire [11:0] u_ca_out_613;
wire [11:0] u_ca_out_614;
wire [11:0] u_ca_out_615;
wire [11:0] u_ca_out_616;
wire [11:0] u_ca_out_617;
wire [11:0] u_ca_out_618;
wire [11:0] u_ca_out_619;
wire [11:0] u_ca_out_620;
wire [11:0] u_ca_out_621;
wire [11:0] u_ca_out_622;
wire [11:0] u_ca_out_623;
wire [11:0] u_ca_out_624;
wire [11:0] u_ca_out_625;
wire [11:0] u_ca_out_626;
wire [11:0] u_ca_out_627;
wire [11:0] u_ca_out_628;
wire [11:0] u_ca_out_629;
wire [11:0] u_ca_out_630;
wire [11:0] u_ca_out_631;
wire [11:0] u_ca_out_632;
wire [11:0] u_ca_out_633;
wire [11:0] u_ca_out_634;
wire [11:0] u_ca_out_635;
wire [11:0] u_ca_out_636;
wire [11:0] u_ca_out_637;
wire [11:0] u_ca_out_638;
wire [11:0] u_ca_out_639;
wire [11:0] u_ca_out_640;
wire [11:0] u_ca_out_641;
wire [11:0] u_ca_out_642;
wire [11:0] u_ca_out_643;
wire [11:0] u_ca_out_644;
wire [11:0] u_ca_out_645;
wire [11:0] u_ca_out_646;
wire [11:0] u_ca_out_647;
wire [11:0] u_ca_out_648;
wire [11:0] u_ca_out_649;
wire [11:0] u_ca_out_650;
wire [11:0] u_ca_out_651;
wire [11:0] u_ca_out_652;
wire [11:0] u_ca_out_653;
wire [11:0] u_ca_out_654;
wire [11:0] u_ca_out_655;
wire [11:0] u_ca_out_656;
wire [11:0] u_ca_out_657;
wire [11:0] u_ca_out_658;
wire [11:0] u_ca_out_659;
wire [11:0] u_ca_out_660;
wire [11:0] u_ca_out_661;
wire [11:0] u_ca_out_662;
wire [11:0] u_ca_out_663;
wire [11:0] u_ca_out_664;
wire [11:0] u_ca_out_665;
wire [11:0] u_ca_out_666;
wire [11:0] u_ca_out_667;
wire [11:0] u_ca_out_668;
wire [11:0] u_ca_out_669;
wire [11:0] u_ca_out_670;
wire [11:0] u_ca_out_671;
wire [11:0] u_ca_out_672;
wire [11:0] u_ca_out_673;
wire [11:0] u_ca_out_674;
wire [11:0] u_ca_out_675;
wire [11:0] u_ca_out_676;
wire [11:0] u_ca_out_677;
wire [11:0] u_ca_out_678;
wire [11:0] u_ca_out_679;
wire [11:0] u_ca_out_680;
wire [11:0] u_ca_out_681;
wire [11:0] u_ca_out_682;
wire [11:0] u_ca_out_683;
wire [11:0] u_ca_out_684;
wire [11:0] u_ca_out_685;
wire [11:0] u_ca_out_686;
wire [11:0] u_ca_out_687;
wire [11:0] u_ca_out_688;
wire [11:0] u_ca_out_689;
wire [11:0] u_ca_out_690;
wire [11:0] u_ca_out_691;
wire [11:0] u_ca_out_692;
wire [11:0] u_ca_out_693;
wire [11:0] u_ca_out_694;
wire [11:0] u_ca_out_695;
wire [11:0] u_ca_out_696;
wire [11:0] u_ca_out_697;
wire [11:0] u_ca_out_698;
wire [11:0] u_ca_out_699;
wire [11:0] u_ca_out_700;
wire [11:0] u_ca_out_701;
wire [11:0] u_ca_out_702;
wire [11:0] u_ca_out_703;
wire [11:0] u_ca_out_704;
wire [11:0] u_ca_out_705;
wire [11:0] u_ca_out_706;
wire [11:0] u_ca_out_707;
wire [11:0] u_ca_out_708;
wire [11:0] u_ca_out_709;
wire [11:0] u_ca_out_710;
wire [11:0] u_ca_out_711;
wire [11:0] u_ca_out_712;
wire [11:0] u_ca_out_713;
wire [11:0] u_ca_out_714;
wire [11:0] u_ca_out_715;
wire [11:0] u_ca_out_716;
wire [11:0] u_ca_out_717;
wire [11:0] u_ca_out_718;
wire [11:0] u_ca_out_719;
wire [11:0] u_ca_out_720;
wire [11:0] u_ca_out_721;
wire [11:0] u_ca_out_722;
wire [11:0] u_ca_out_723;
wire [11:0] u_ca_out_724;
wire [11:0] u_ca_out_725;
wire [11:0] u_ca_out_726;
wire [11:0] u_ca_out_727;
wire [11:0] u_ca_out_728;
wire [11:0] u_ca_out_729;
wire [11:0] u_ca_out_730;
wire [11:0] u_ca_out_731;
wire [11:0] u_ca_out_732;
wire [11:0] u_ca_out_733;
wire [11:0] u_ca_out_734;
wire [11:0] u_ca_out_735;
wire [11:0] u_ca_out_736;
wire [11:0] u_ca_out_737;
wire [11:0] u_ca_out_738;
wire [11:0] u_ca_out_739;
wire [11:0] u_ca_out_740;
wire [11:0] u_ca_out_741;
wire [11:0] u_ca_out_742;
wire [11:0] u_ca_out_743;
wire [11:0] u_ca_out_744;
wire [11:0] u_ca_out_745;
wire [11:0] u_ca_out_746;
wire [11:0] u_ca_out_747;
wire [11:0] u_ca_out_748;
wire [11:0] u_ca_out_749;
wire [11:0] u_ca_out_750;
wire [11:0] u_ca_out_751;
wire [11:0] u_ca_out_752;
wire [11:0] u_ca_out_753;
wire [11:0] u_ca_out_754;
wire [11:0] u_ca_out_755;
wire [11:0] u_ca_out_756;
wire [11:0] u_ca_out_757;
wire [11:0] u_ca_out_758;
wire [11:0] u_ca_out_759;
wire [11:0] u_ca_out_760;
wire [11:0] u_ca_out_761;
wire [11:0] u_ca_out_762;
wire [11:0] u_ca_out_763;
wire [11:0] u_ca_out_764;
wire [11:0] u_ca_out_765;
wire [11:0] u_ca_out_766;
wire [11:0] u_ca_out_767;
wire [11:0] u_ca_out_768;
wire [11:0] u_ca_out_769;
wire [11:0] u_ca_out_770;
wire [11:0] u_ca_out_771;
wire [11:0] u_ca_out_772;
wire [11:0] u_ca_out_773;
wire [11:0] u_ca_out_774;
wire [11:0] u_ca_out_775;
wire [11:0] u_ca_out_776;
wire [11:0] u_ca_out_777;
wire [11:0] u_ca_out_778;
wire [11:0] u_ca_out_779;
wire [11:0] u_ca_out_780;
wire [11:0] u_ca_out_781;
wire [11:0] u_ca_out_782;
wire [11:0] u_ca_out_783;
wire [11:0] u_ca_out_784;
wire [11:0] u_ca_out_785;
wire [11:0] u_ca_out_786;
wire [11:0] u_ca_out_787;
wire [11:0] u_ca_out_788;
wire [11:0] u_ca_out_789;
wire [11:0] u_ca_out_790;
wire [11:0] u_ca_out_791;
wire [11:0] u_ca_out_792;
wire [11:0] u_ca_out_793;
wire [11:0] u_ca_out_794;
wire [11:0] u_ca_out_795;
wire [11:0] u_ca_out_796;
wire [11:0] u_ca_out_797;
wire [11:0] u_ca_out_798;
wire [11:0] u_ca_out_799;
wire [11:0] u_ca_out_800;
wire [11:0] u_ca_out_801;
wire [11:0] u_ca_out_802;
wire [11:0] u_ca_out_803;
wire [11:0] u_ca_out_804;
wire [11:0] u_ca_out_805;
wire [11:0] u_ca_out_806;
wire [11:0] u_ca_out_807;
wire [11:0] u_ca_out_808;
wire [11:0] u_ca_out_809;
wire [11:0] u_ca_out_810;
wire [11:0] u_ca_out_811;
wire [11:0] u_ca_out_812;
wire [11:0] u_ca_out_813;
wire [11:0] u_ca_out_814;
wire [11:0] u_ca_out_815;
wire [11:0] u_ca_out_816;
wire [11:0] u_ca_out_817;
wire [11:0] u_ca_out_818;
wire [11:0] u_ca_out_819;
wire [11:0] u_ca_out_820;
wire [11:0] u_ca_out_821;
wire [11:0] u_ca_out_822;
wire [11:0] u_ca_out_823;
wire [11:0] u_ca_out_824;
wire [11:0] u_ca_out_825;
wire [11:0] u_ca_out_826;
wire [11:0] u_ca_out_827;
wire [11:0] u_ca_out_828;
wire [11:0] u_ca_out_829;
wire [11:0] u_ca_out_830;
wire [11:0] u_ca_out_831;
wire [11:0] u_ca_out_832;
wire [11:0] u_ca_out_833;
wire [11:0] u_ca_out_834;
wire [11:0] u_ca_out_835;
wire [11:0] u_ca_out_836;
wire [11:0] u_ca_out_837;
wire [11:0] u_ca_out_838;
wire [11:0] u_ca_out_839;
wire [11:0] u_ca_out_840;
wire [11:0] u_ca_out_841;
wire [11:0] u_ca_out_842;
wire [11:0] u_ca_out_843;
wire [11:0] u_ca_out_844;
wire [11:0] u_ca_out_845;
wire [11:0] u_ca_out_846;
wire [11:0] u_ca_out_847;
wire [11:0] u_ca_out_848;
wire [11:0] u_ca_out_849;
wire [11:0] u_ca_out_850;
wire [11:0] u_ca_out_851;
wire [11:0] u_ca_out_852;
wire [11:0] u_ca_out_853;
wire [11:0] u_ca_out_854;
wire [11:0] u_ca_out_855;
wire [11:0] u_ca_out_856;
wire [11:0] u_ca_out_857;
wire [11:0] u_ca_out_858;
wire [11:0] u_ca_out_859;
wire [11:0] u_ca_out_860;
wire [11:0] u_ca_out_861;
wire [11:0] u_ca_out_862;
wire [11:0] u_ca_out_863;
wire [11:0] u_ca_out_864;
wire [11:0] u_ca_out_865;
wire [11:0] u_ca_out_866;
wire [11:0] u_ca_out_867;
wire [11:0] u_ca_out_868;
wire [11:0] u_ca_out_869;
wire [11:0] u_ca_out_870;
wire [11:0] u_ca_out_871;
wire [11:0] u_ca_out_872;
wire [11:0] u_ca_out_873;
wire [11:0] u_ca_out_874;
wire [11:0] u_ca_out_875;
wire [11:0] u_ca_out_876;
wire [11:0] u_ca_out_877;
wire [11:0] u_ca_out_878;
wire [11:0] u_ca_out_879;
wire [11:0] u_ca_out_880;
wire [11:0] u_ca_out_881;
wire [11:0] u_ca_out_882;
wire [11:0] u_ca_out_883;
wire [11:0] u_ca_out_884;
wire [11:0] u_ca_out_885;
wire [11:0] u_ca_out_886;
wire [11:0] u_ca_out_887;
wire [11:0] u_ca_out_888;
wire [11:0] u_ca_out_889;
wire [11:0] u_ca_out_890;
wire [11:0] u_ca_out_891;
wire [11:0] u_ca_out_892;
wire [11:0] u_ca_out_893;
wire [11:0] u_ca_out_894;
wire [11:0] u_ca_out_895;
wire [11:0] u_ca_out_896;
wire [11:0] u_ca_out_897;
wire [11:0] u_ca_out_898;
wire [11:0] u_ca_out_899;
wire [11:0] u_ca_out_900;
wire [11:0] u_ca_out_901;
wire [11:0] u_ca_out_902;
wire [11:0] u_ca_out_903;
wire [11:0] u_ca_out_904;
wire [11:0] u_ca_out_905;
wire [11:0] u_ca_out_906;
wire [11:0] u_ca_out_907;
wire [11:0] u_ca_out_908;
wire [11:0] u_ca_out_909;
wire [11:0] u_ca_out_910;
wire [11:0] u_ca_out_911;
wire [11:0] u_ca_out_912;
wire [11:0] u_ca_out_913;
wire [11:0] u_ca_out_914;
wire [11:0] u_ca_out_915;
wire [11:0] u_ca_out_916;
wire [11:0] u_ca_out_917;
wire [11:0] u_ca_out_918;
wire [11:0] u_ca_out_919;
wire [11:0] u_ca_out_920;
wire [11:0] u_ca_out_921;
wire [11:0] u_ca_out_922;
wire [11:0] u_ca_out_923;
wire [11:0] u_ca_out_924;
wire [11:0] u_ca_out_925;
wire [11:0] u_ca_out_926;
wire [11:0] u_ca_out_927;
wire [11:0] u_ca_out_928;
wire [11:0] u_ca_out_929;
wire [11:0] u_ca_out_930;
wire [11:0] u_ca_out_931;
wire [11:0] u_ca_out_932;
wire [11:0] u_ca_out_933;
wire [11:0] u_ca_out_934;
wire [11:0] u_ca_out_935;
wire [11:0] u_ca_out_936;
wire [11:0] u_ca_out_937;
wire [11:0] u_ca_out_938;
wire [11:0] u_ca_out_939;
wire [11:0] u_ca_out_940;
wire [11:0] u_ca_out_941;
wire [11:0] u_ca_out_942;
wire [11:0] u_ca_out_943;
wire [11:0] u_ca_out_944;
wire [11:0] u_ca_out_945;
wire [11:0] u_ca_out_946;
wire [11:0] u_ca_out_947;
wire [11:0] u_ca_out_948;
wire [11:0] u_ca_out_949;
wire [11:0] u_ca_out_950;
wire [11:0] u_ca_out_951;
wire [11:0] u_ca_out_952;
wire [11:0] u_ca_out_953;
wire [11:0] u_ca_out_954;
wire [11:0] u_ca_out_955;
wire [11:0] u_ca_out_956;
wire [11:0] u_ca_out_957;
wire [11:0] u_ca_out_958;
wire [11:0] u_ca_out_959;
wire [11:0] u_ca_out_960;
wire [11:0] u_ca_out_961;
wire [11:0] u_ca_out_962;
wire [11:0] u_ca_out_963;
wire [11:0] u_ca_out_964;
wire [11:0] u_ca_out_965;
wire [11:0] u_ca_out_966;
wire [11:0] u_ca_out_967;
wire [11:0] u_ca_out_968;
wire [11:0] u_ca_out_969;
wire [11:0] u_ca_out_970;
wire [11:0] u_ca_out_971;
wire [11:0] u_ca_out_972;
wire [11:0] u_ca_out_973;
wire [11:0] u_ca_out_974;
wire [11:0] u_ca_out_975;
wire [11:0] u_ca_out_976;
wire [11:0] u_ca_out_977;
wire [11:0] u_ca_out_978;
wire [11:0] u_ca_out_979;
wire [11:0] u_ca_out_980;
wire [11:0] u_ca_out_981;
wire [11:0] u_ca_out_982;
wire [11:0] u_ca_out_983;
wire [11:0] u_ca_out_984;
wire [11:0] u_ca_out_985;
wire [11:0] u_ca_out_986;
wire [11:0] u_ca_out_987;
wire [11:0] u_ca_out_988;
wire [11:0] u_ca_out_989;
wire [11:0] u_ca_out_990;
wire [11:0] u_ca_out_991;
wire [11:0] u_ca_out_992;
wire [11:0] u_ca_out_993;
wire [11:0] u_ca_out_994;
wire [11:0] u_ca_out_995;
wire [11:0] u_ca_out_996;
wire [11:0] u_ca_out_997;
wire [11:0] u_ca_out_998;
wire [11:0] u_ca_out_999;
wire [11:0] u_ca_out_1000;
wire [11:0] u_ca_out_1001;
wire [11:0] u_ca_out_1002;
wire [11:0] u_ca_out_1003;
wire [11:0] u_ca_out_1004;
wire [11:0] u_ca_out_1005;
wire [11:0] u_ca_out_1006;
wire [11:0] u_ca_out_1007;
wire [11:0] u_ca_out_1008;
wire [11:0] u_ca_out_1009;
wire [11:0] u_ca_out_1010;
wire [11:0] u_ca_out_1011;
wire [11:0] u_ca_out_1012;
wire [11:0] u_ca_out_1013;
wire [11:0] u_ca_out_1014;
wire [11:0] u_ca_out_1015;
wire [11:0] u_ca_out_1016;
wire [11:0] u_ca_out_1017;
wire [11:0] u_ca_out_1018;
wire [11:0] u_ca_out_1019;
wire [11:0] u_ca_out_1020;
wire [11:0] u_ca_out_1021;
wire [11:0] u_ca_out_1022;
wire [11:0] u_ca_out_1023;
wire [11:0] u_ca_out_1024;
wire [11:0] u_ca_out_1025;
wire [11:0] u_ca_out_1026;
wire [11:0] u_ca_out_1027;
wire [11:0] u_ca_out_1028;
wire [11:0] u_ca_out_1029;
wire [11:0] u_ca_out_1030;
wire [11:0] u_ca_out_1031;
wire [11:0] u_ca_out_1032;

assign u_ca_in_0 = {{2{1'b0}}, col_in_0};
assign u_ca_in_1 = {{2{1'b0}}, col_in_1};
assign u_ca_in_2 = {{2{1'b0}}, col_in_2};
assign u_ca_in_3 = {{2{1'b0}}, col_in_3};
assign u_ca_in_4 = {{2{1'b0}}, col_in_4};
assign u_ca_in_5 = {{2{1'b0}}, col_in_5};
assign u_ca_in_6 = {{2{1'b0}}, col_in_6};
assign u_ca_in_7 = {{2{1'b0}}, col_in_7};
assign u_ca_in_8 = {{2{1'b0}}, col_in_8};
assign u_ca_in_9 = {{2{1'b0}}, col_in_9};
assign u_ca_in_10 = {{2{1'b0}}, col_in_10};
assign u_ca_in_11 = {{2{1'b0}}, col_in_11};
assign u_ca_in_12 = {{2{1'b0}}, col_in_12};
assign u_ca_in_13 = {{2{1'b0}}, col_in_13};
assign u_ca_in_14 = {{2{1'b0}}, col_in_14};
assign u_ca_in_15 = {{2{1'b0}}, col_in_15};
assign u_ca_in_16 = {{2{1'b0}}, col_in_16};
assign u_ca_in_17 = {{2{1'b0}}, col_in_17};
assign u_ca_in_18 = {{2{1'b0}}, col_in_18};
assign u_ca_in_19 = {{2{1'b0}}, col_in_19};
assign u_ca_in_20 = {{2{1'b0}}, col_in_20};
assign u_ca_in_21 = {{2{1'b0}}, col_in_21};
assign u_ca_in_22 = {{2{1'b0}}, col_in_22};
assign u_ca_in_23 = {{2{1'b0}}, col_in_23};
assign u_ca_in_24 = {{2{1'b0}}, col_in_24};
assign u_ca_in_25 = {{2{1'b0}}, col_in_25};
assign u_ca_in_26 = {{2{1'b0}}, col_in_26};
assign u_ca_in_27 = {{2{1'b0}}, col_in_27};
assign u_ca_in_28 = {{2{1'b0}}, col_in_28};
assign u_ca_in_29 = {{2{1'b0}}, col_in_29};
assign u_ca_in_30 = {{2{1'b0}}, col_in_30};
assign u_ca_in_31 = {{2{1'b0}}, col_in_31};
assign u_ca_in_32 = {{2{1'b0}}, col_in_32};
assign u_ca_in_33 = {{2{1'b0}}, col_in_33};
assign u_ca_in_34 = {{2{1'b0}}, col_in_34};
assign u_ca_in_35 = {{2{1'b0}}, col_in_35};
assign u_ca_in_36 = {{2{1'b0}}, col_in_36};
assign u_ca_in_37 = {{2{1'b0}}, col_in_37};
assign u_ca_in_38 = {{2{1'b0}}, col_in_38};
assign u_ca_in_39 = {{2{1'b0}}, col_in_39};
assign u_ca_in_40 = {{2{1'b0}}, col_in_40};
assign u_ca_in_41 = {{2{1'b0}}, col_in_41};
assign u_ca_in_42 = {{2{1'b0}}, col_in_42};
assign u_ca_in_43 = {{2{1'b0}}, col_in_43};
assign u_ca_in_44 = {{2{1'b0}}, col_in_44};
assign u_ca_in_45 = {{2{1'b0}}, col_in_45};
assign u_ca_in_46 = {{2{1'b0}}, col_in_46};
assign u_ca_in_47 = {{2{1'b0}}, col_in_47};
assign u_ca_in_48 = {{2{1'b0}}, col_in_48};
assign u_ca_in_49 = {{2{1'b0}}, col_in_49};
assign u_ca_in_50 = {{2{1'b0}}, col_in_50};
assign u_ca_in_51 = {{2{1'b0}}, col_in_51};
assign u_ca_in_52 = {{2{1'b0}}, col_in_52};
assign u_ca_in_53 = {{2{1'b0}}, col_in_53};
assign u_ca_in_54 = {{2{1'b0}}, col_in_54};
assign u_ca_in_55 = {{2{1'b0}}, col_in_55};
assign u_ca_in_56 = {{2{1'b0}}, col_in_56};
assign u_ca_in_57 = {{2{1'b0}}, col_in_57};
assign u_ca_in_58 = {{2{1'b0}}, col_in_58};
assign u_ca_in_59 = {{2{1'b0}}, col_in_59};
assign u_ca_in_60 = {{2{1'b0}}, col_in_60};
assign u_ca_in_61 = {{2{1'b0}}, col_in_61};
assign u_ca_in_62 = {{2{1'b0}}, col_in_62};
assign u_ca_in_63 = {{2{1'b0}}, col_in_63};
assign u_ca_in_64 = {{2{1'b0}}, col_in_64};
assign u_ca_in_65 = {{2{1'b0}}, col_in_65};
assign u_ca_in_66 = {{2{1'b0}}, col_in_66};
assign u_ca_in_67 = {{2{1'b0}}, col_in_67};
assign u_ca_in_68 = {{2{1'b0}}, col_in_68};
assign u_ca_in_69 = {{2{1'b0}}, col_in_69};
assign u_ca_in_70 = {{2{1'b0}}, col_in_70};
assign u_ca_in_71 = {{2{1'b0}}, col_in_71};
assign u_ca_in_72 = {{2{1'b0}}, col_in_72};
assign u_ca_in_73 = {{2{1'b0}}, col_in_73};
assign u_ca_in_74 = {{2{1'b0}}, col_in_74};
assign u_ca_in_75 = {{2{1'b0}}, col_in_75};
assign u_ca_in_76 = {{2{1'b0}}, col_in_76};
assign u_ca_in_77 = {{2{1'b0}}, col_in_77};
assign u_ca_in_78 = {{2{1'b0}}, col_in_78};
assign u_ca_in_79 = {{2{1'b0}}, col_in_79};
assign u_ca_in_80 = {{2{1'b0}}, col_in_80};
assign u_ca_in_81 = {{2{1'b0}}, col_in_81};
assign u_ca_in_82 = {{2{1'b0}}, col_in_82};
assign u_ca_in_83 = {{2{1'b0}}, col_in_83};
assign u_ca_in_84 = {{2{1'b0}}, col_in_84};
assign u_ca_in_85 = {{2{1'b0}}, col_in_85};
assign u_ca_in_86 = {{2{1'b0}}, col_in_86};
assign u_ca_in_87 = {{2{1'b0}}, col_in_87};
assign u_ca_in_88 = {{2{1'b0}}, col_in_88};
assign u_ca_in_89 = {{2{1'b0}}, col_in_89};
assign u_ca_in_90 = {{2{1'b0}}, col_in_90};
assign u_ca_in_91 = {{2{1'b0}}, col_in_91};
assign u_ca_in_92 = {{2{1'b0}}, col_in_92};
assign u_ca_in_93 = {{2{1'b0}}, col_in_93};
assign u_ca_in_94 = {{2{1'b0}}, col_in_94};
assign u_ca_in_95 = {{2{1'b0}}, col_in_95};
assign u_ca_in_96 = {{2{1'b0}}, col_in_96};
assign u_ca_in_97 = {{2{1'b0}}, col_in_97};
assign u_ca_in_98 = {{2{1'b0}}, col_in_98};
assign u_ca_in_99 = {{2{1'b0}}, col_in_99};
assign u_ca_in_100 = {{2{1'b0}}, col_in_100};
assign u_ca_in_101 = {{2{1'b0}}, col_in_101};
assign u_ca_in_102 = {{2{1'b0}}, col_in_102};
assign u_ca_in_103 = {{2{1'b0}}, col_in_103};
assign u_ca_in_104 = {{2{1'b0}}, col_in_104};
assign u_ca_in_105 = {{2{1'b0}}, col_in_105};
assign u_ca_in_106 = {{2{1'b0}}, col_in_106};
assign u_ca_in_107 = {{2{1'b0}}, col_in_107};
assign u_ca_in_108 = {{2{1'b0}}, col_in_108};
assign u_ca_in_109 = {{2{1'b0}}, col_in_109};
assign u_ca_in_110 = {{2{1'b0}}, col_in_110};
assign u_ca_in_111 = {{2{1'b0}}, col_in_111};
assign u_ca_in_112 = {{2{1'b0}}, col_in_112};
assign u_ca_in_113 = {{2{1'b0}}, col_in_113};
assign u_ca_in_114 = {{2{1'b0}}, col_in_114};
assign u_ca_in_115 = {{2{1'b0}}, col_in_115};
assign u_ca_in_116 = {{2{1'b0}}, col_in_116};
assign u_ca_in_117 = {{2{1'b0}}, col_in_117};
assign u_ca_in_118 = {{2{1'b0}}, col_in_118};
assign u_ca_in_119 = {{2{1'b0}}, col_in_119};
assign u_ca_in_120 = {{2{1'b0}}, col_in_120};
assign u_ca_in_121 = {{2{1'b0}}, col_in_121};
assign u_ca_in_122 = {{2{1'b0}}, col_in_122};
assign u_ca_in_123 = {{2{1'b0}}, col_in_123};
assign u_ca_in_124 = {{2{1'b0}}, col_in_124};
assign u_ca_in_125 = {{2{1'b0}}, col_in_125};
assign u_ca_in_126 = {{2{1'b0}}, col_in_126};
assign u_ca_in_127 = {{2{1'b0}}, col_in_127};
assign u_ca_in_128 = {{2{1'b0}}, col_in_128};
assign u_ca_in_129 = {{2{1'b0}}, col_in_129};
assign u_ca_in_130 = {{2{1'b0}}, col_in_130};
assign u_ca_in_131 = {{2{1'b0}}, col_in_131};
assign u_ca_in_132 = {{2{1'b0}}, col_in_132};
assign u_ca_in_133 = {{2{1'b0}}, col_in_133};
assign u_ca_in_134 = {{2{1'b0}}, col_in_134};
assign u_ca_in_135 = {{2{1'b0}}, col_in_135};
assign u_ca_in_136 = {{2{1'b0}}, col_in_136};
assign u_ca_in_137 = {{2{1'b0}}, col_in_137};
assign u_ca_in_138 = {{2{1'b0}}, col_in_138};
assign u_ca_in_139 = {{2{1'b0}}, col_in_139};
assign u_ca_in_140 = {{2{1'b0}}, col_in_140};
assign u_ca_in_141 = {{2{1'b0}}, col_in_141};
assign u_ca_in_142 = {{2{1'b0}}, col_in_142};
assign u_ca_in_143 = {{2{1'b0}}, col_in_143};
assign u_ca_in_144 = {{2{1'b0}}, col_in_144};
assign u_ca_in_145 = {{2{1'b0}}, col_in_145};
assign u_ca_in_146 = {{2{1'b0}}, col_in_146};
assign u_ca_in_147 = {{2{1'b0}}, col_in_147};
assign u_ca_in_148 = {{2{1'b0}}, col_in_148};
assign u_ca_in_149 = {{2{1'b0}}, col_in_149};
assign u_ca_in_150 = {{2{1'b0}}, col_in_150};
assign u_ca_in_151 = {{2{1'b0}}, col_in_151};
assign u_ca_in_152 = {{2{1'b0}}, col_in_152};
assign u_ca_in_153 = {{2{1'b0}}, col_in_153};
assign u_ca_in_154 = {{2{1'b0}}, col_in_154};
assign u_ca_in_155 = {{2{1'b0}}, col_in_155};
assign u_ca_in_156 = {{2{1'b0}}, col_in_156};
assign u_ca_in_157 = {{2{1'b0}}, col_in_157};
assign u_ca_in_158 = {{2{1'b0}}, col_in_158};
assign u_ca_in_159 = {{2{1'b0}}, col_in_159};
assign u_ca_in_160 = {{2{1'b0}}, col_in_160};
assign u_ca_in_161 = {{2{1'b0}}, col_in_161};
assign u_ca_in_162 = {{2{1'b0}}, col_in_162};
assign u_ca_in_163 = {{2{1'b0}}, col_in_163};
assign u_ca_in_164 = {{2{1'b0}}, col_in_164};
assign u_ca_in_165 = {{2{1'b0}}, col_in_165};
assign u_ca_in_166 = {{2{1'b0}}, col_in_166};
assign u_ca_in_167 = {{2{1'b0}}, col_in_167};
assign u_ca_in_168 = {{2{1'b0}}, col_in_168};
assign u_ca_in_169 = {{2{1'b0}}, col_in_169};
assign u_ca_in_170 = {{2{1'b0}}, col_in_170};
assign u_ca_in_171 = {{2{1'b0}}, col_in_171};
assign u_ca_in_172 = {{2{1'b0}}, col_in_172};
assign u_ca_in_173 = {{2{1'b0}}, col_in_173};
assign u_ca_in_174 = {{2{1'b0}}, col_in_174};
assign u_ca_in_175 = {{2{1'b0}}, col_in_175};
assign u_ca_in_176 = {{2{1'b0}}, col_in_176};
assign u_ca_in_177 = {{2{1'b0}}, col_in_177};
assign u_ca_in_178 = {{2{1'b0}}, col_in_178};
assign u_ca_in_179 = {{2{1'b0}}, col_in_179};
assign u_ca_in_180 = {{2{1'b0}}, col_in_180};
assign u_ca_in_181 = {{2{1'b0}}, col_in_181};
assign u_ca_in_182 = {{2{1'b0}}, col_in_182};
assign u_ca_in_183 = {{2{1'b0}}, col_in_183};
assign u_ca_in_184 = {{2{1'b0}}, col_in_184};
assign u_ca_in_185 = {{2{1'b0}}, col_in_185};
assign u_ca_in_186 = {{2{1'b0}}, col_in_186};
assign u_ca_in_187 = {{2{1'b0}}, col_in_187};
assign u_ca_in_188 = {{2{1'b0}}, col_in_188};
assign u_ca_in_189 = {{2{1'b0}}, col_in_189};
assign u_ca_in_190 = {{2{1'b0}}, col_in_190};
assign u_ca_in_191 = {{2{1'b0}}, col_in_191};
assign u_ca_in_192 = {{2{1'b0}}, col_in_192};
assign u_ca_in_193 = {{2{1'b0}}, col_in_193};
assign u_ca_in_194 = {{2{1'b0}}, col_in_194};
assign u_ca_in_195 = {{2{1'b0}}, col_in_195};
assign u_ca_in_196 = {{2{1'b0}}, col_in_196};
assign u_ca_in_197 = {{2{1'b0}}, col_in_197};
assign u_ca_in_198 = {{2{1'b0}}, col_in_198};
assign u_ca_in_199 = {{2{1'b0}}, col_in_199};
assign u_ca_in_200 = {{2{1'b0}}, col_in_200};
assign u_ca_in_201 = {{2{1'b0}}, col_in_201};
assign u_ca_in_202 = {{2{1'b0}}, col_in_202};
assign u_ca_in_203 = {{2{1'b0}}, col_in_203};
assign u_ca_in_204 = {{2{1'b0}}, col_in_204};
assign u_ca_in_205 = {{2{1'b0}}, col_in_205};
assign u_ca_in_206 = {{2{1'b0}}, col_in_206};
assign u_ca_in_207 = {{2{1'b0}}, col_in_207};
assign u_ca_in_208 = {{2{1'b0}}, col_in_208};
assign u_ca_in_209 = {{2{1'b0}}, col_in_209};
assign u_ca_in_210 = {{2{1'b0}}, col_in_210};
assign u_ca_in_211 = {{2{1'b0}}, col_in_211};
assign u_ca_in_212 = {{2{1'b0}}, col_in_212};
assign u_ca_in_213 = {{2{1'b0}}, col_in_213};
assign u_ca_in_214 = {{2{1'b0}}, col_in_214};
assign u_ca_in_215 = {{2{1'b0}}, col_in_215};
assign u_ca_in_216 = {{2{1'b0}}, col_in_216};
assign u_ca_in_217 = {{2{1'b0}}, col_in_217};
assign u_ca_in_218 = {{2{1'b0}}, col_in_218};
assign u_ca_in_219 = {{2{1'b0}}, col_in_219};
assign u_ca_in_220 = {{2{1'b0}}, col_in_220};
assign u_ca_in_221 = {{2{1'b0}}, col_in_221};
assign u_ca_in_222 = {{2{1'b0}}, col_in_222};
assign u_ca_in_223 = {{2{1'b0}}, col_in_223};
assign u_ca_in_224 = {{2{1'b0}}, col_in_224};
assign u_ca_in_225 = {{2{1'b0}}, col_in_225};
assign u_ca_in_226 = {{2{1'b0}}, col_in_226};
assign u_ca_in_227 = {{2{1'b0}}, col_in_227};
assign u_ca_in_228 = {{2{1'b0}}, col_in_228};
assign u_ca_in_229 = {{2{1'b0}}, col_in_229};
assign u_ca_in_230 = {{2{1'b0}}, col_in_230};
assign u_ca_in_231 = {{2{1'b0}}, col_in_231};
assign u_ca_in_232 = {{2{1'b0}}, col_in_232};
assign u_ca_in_233 = {{2{1'b0}}, col_in_233};
assign u_ca_in_234 = {{2{1'b0}}, col_in_234};
assign u_ca_in_235 = {{2{1'b0}}, col_in_235};
assign u_ca_in_236 = {{2{1'b0}}, col_in_236};
assign u_ca_in_237 = {{2{1'b0}}, col_in_237};
assign u_ca_in_238 = {{2{1'b0}}, col_in_238};
assign u_ca_in_239 = {{2{1'b0}}, col_in_239};
assign u_ca_in_240 = {{2{1'b0}}, col_in_240};
assign u_ca_in_241 = {{2{1'b0}}, col_in_241};
assign u_ca_in_242 = {{2{1'b0}}, col_in_242};
assign u_ca_in_243 = {{2{1'b0}}, col_in_243};
assign u_ca_in_244 = {{2{1'b0}}, col_in_244};
assign u_ca_in_245 = {{2{1'b0}}, col_in_245};
assign u_ca_in_246 = {{2{1'b0}}, col_in_246};
assign u_ca_in_247 = {{2{1'b0}}, col_in_247};
assign u_ca_in_248 = {{2{1'b0}}, col_in_248};
assign u_ca_in_249 = {{2{1'b0}}, col_in_249};
assign u_ca_in_250 = {{2{1'b0}}, col_in_250};
assign u_ca_in_251 = {{2{1'b0}}, col_in_251};
assign u_ca_in_252 = {{2{1'b0}}, col_in_252};
assign u_ca_in_253 = {{2{1'b0}}, col_in_253};
assign u_ca_in_254 = {{2{1'b0}}, col_in_254};
assign u_ca_in_255 = {{2{1'b0}}, col_in_255};
assign u_ca_in_256 = {{2{1'b0}}, col_in_256};
assign u_ca_in_257 = {{2{1'b0}}, col_in_257};
assign u_ca_in_258 = {{2{1'b0}}, col_in_258};
assign u_ca_in_259 = {{2{1'b0}}, col_in_259};
assign u_ca_in_260 = {{2{1'b0}}, col_in_260};
assign u_ca_in_261 = {{2{1'b0}}, col_in_261};
assign u_ca_in_262 = {{2{1'b0}}, col_in_262};
assign u_ca_in_263 = {{2{1'b0}}, col_in_263};
assign u_ca_in_264 = {{2{1'b0}}, col_in_264};
assign u_ca_in_265 = {{2{1'b0}}, col_in_265};
assign u_ca_in_266 = {{2{1'b0}}, col_in_266};
assign u_ca_in_267 = {{2{1'b0}}, col_in_267};
assign u_ca_in_268 = {{2{1'b0}}, col_in_268};
assign u_ca_in_269 = {{2{1'b0}}, col_in_269};
assign u_ca_in_270 = {{2{1'b0}}, col_in_270};
assign u_ca_in_271 = {{2{1'b0}}, col_in_271};
assign u_ca_in_272 = {{2{1'b0}}, col_in_272};
assign u_ca_in_273 = {{2{1'b0}}, col_in_273};
assign u_ca_in_274 = {{2{1'b0}}, col_in_274};
assign u_ca_in_275 = {{2{1'b0}}, col_in_275};
assign u_ca_in_276 = {{2{1'b0}}, col_in_276};
assign u_ca_in_277 = {{2{1'b0}}, col_in_277};
assign u_ca_in_278 = {{2{1'b0}}, col_in_278};
assign u_ca_in_279 = {{2{1'b0}}, col_in_279};
assign u_ca_in_280 = {{2{1'b0}}, col_in_280};
assign u_ca_in_281 = {{2{1'b0}}, col_in_281};
assign u_ca_in_282 = {{2{1'b0}}, col_in_282};
assign u_ca_in_283 = {{2{1'b0}}, col_in_283};
assign u_ca_in_284 = {{2{1'b0}}, col_in_284};
assign u_ca_in_285 = {{2{1'b0}}, col_in_285};
assign u_ca_in_286 = {{2{1'b0}}, col_in_286};
assign u_ca_in_287 = {{2{1'b0}}, col_in_287};
assign u_ca_in_288 = {{2{1'b0}}, col_in_288};
assign u_ca_in_289 = {{2{1'b0}}, col_in_289};
assign u_ca_in_290 = {{2{1'b0}}, col_in_290};
assign u_ca_in_291 = {{2{1'b0}}, col_in_291};
assign u_ca_in_292 = {{2{1'b0}}, col_in_292};
assign u_ca_in_293 = {{2{1'b0}}, col_in_293};
assign u_ca_in_294 = {{2{1'b0}}, col_in_294};
assign u_ca_in_295 = {{2{1'b0}}, col_in_295};
assign u_ca_in_296 = {{2{1'b0}}, col_in_296};
assign u_ca_in_297 = {{2{1'b0}}, col_in_297};
assign u_ca_in_298 = {{2{1'b0}}, col_in_298};
assign u_ca_in_299 = {{2{1'b0}}, col_in_299};
assign u_ca_in_300 = {{2{1'b0}}, col_in_300};
assign u_ca_in_301 = {{2{1'b0}}, col_in_301};
assign u_ca_in_302 = {{2{1'b0}}, col_in_302};
assign u_ca_in_303 = {{2{1'b0}}, col_in_303};
assign u_ca_in_304 = {{2{1'b0}}, col_in_304};
assign u_ca_in_305 = {{2{1'b0}}, col_in_305};
assign u_ca_in_306 = {{2{1'b0}}, col_in_306};
assign u_ca_in_307 = {{2{1'b0}}, col_in_307};
assign u_ca_in_308 = {{2{1'b0}}, col_in_308};
assign u_ca_in_309 = {{2{1'b0}}, col_in_309};
assign u_ca_in_310 = {{2{1'b0}}, col_in_310};
assign u_ca_in_311 = {{2{1'b0}}, col_in_311};
assign u_ca_in_312 = {{2{1'b0}}, col_in_312};
assign u_ca_in_313 = {{2{1'b0}}, col_in_313};
assign u_ca_in_314 = {{2{1'b0}}, col_in_314};
assign u_ca_in_315 = {{2{1'b0}}, col_in_315};
assign u_ca_in_316 = {{2{1'b0}}, col_in_316};
assign u_ca_in_317 = {{2{1'b0}}, col_in_317};
assign u_ca_in_318 = {{2{1'b0}}, col_in_318};
assign u_ca_in_319 = {{2{1'b0}}, col_in_319};
assign u_ca_in_320 = {{2{1'b0}}, col_in_320};
assign u_ca_in_321 = {{2{1'b0}}, col_in_321};
assign u_ca_in_322 = {{2{1'b0}}, col_in_322};
assign u_ca_in_323 = {{2{1'b0}}, col_in_323};
assign u_ca_in_324 = {{2{1'b0}}, col_in_324};
assign u_ca_in_325 = {{2{1'b0}}, col_in_325};
assign u_ca_in_326 = {{2{1'b0}}, col_in_326};
assign u_ca_in_327 = {{2{1'b0}}, col_in_327};
assign u_ca_in_328 = {{2{1'b0}}, col_in_328};
assign u_ca_in_329 = {{2{1'b0}}, col_in_329};
assign u_ca_in_330 = {{2{1'b0}}, col_in_330};
assign u_ca_in_331 = {{2{1'b0}}, col_in_331};
assign u_ca_in_332 = {{2{1'b0}}, col_in_332};
assign u_ca_in_333 = {{2{1'b0}}, col_in_333};
assign u_ca_in_334 = {{2{1'b0}}, col_in_334};
assign u_ca_in_335 = {{2{1'b0}}, col_in_335};
assign u_ca_in_336 = {{2{1'b0}}, col_in_336};
assign u_ca_in_337 = {{2{1'b0}}, col_in_337};
assign u_ca_in_338 = {{2{1'b0}}, col_in_338};
assign u_ca_in_339 = {{2{1'b0}}, col_in_339};
assign u_ca_in_340 = {{2{1'b0}}, col_in_340};
assign u_ca_in_341 = {{2{1'b0}}, col_in_341};
assign u_ca_in_342 = {{2{1'b0}}, col_in_342};
assign u_ca_in_343 = {{2{1'b0}}, col_in_343};
assign u_ca_in_344 = {{2{1'b0}}, col_in_344};
assign u_ca_in_345 = {{2{1'b0}}, col_in_345};
assign u_ca_in_346 = {{2{1'b0}}, col_in_346};
assign u_ca_in_347 = {{2{1'b0}}, col_in_347};
assign u_ca_in_348 = {{2{1'b0}}, col_in_348};
assign u_ca_in_349 = {{2{1'b0}}, col_in_349};
assign u_ca_in_350 = {{2{1'b0}}, col_in_350};
assign u_ca_in_351 = {{2{1'b0}}, col_in_351};
assign u_ca_in_352 = {{2{1'b0}}, col_in_352};
assign u_ca_in_353 = {{2{1'b0}}, col_in_353};
assign u_ca_in_354 = {{2{1'b0}}, col_in_354};
assign u_ca_in_355 = {{2{1'b0}}, col_in_355};
assign u_ca_in_356 = {{2{1'b0}}, col_in_356};
assign u_ca_in_357 = {{2{1'b0}}, col_in_357};
assign u_ca_in_358 = {{2{1'b0}}, col_in_358};
assign u_ca_in_359 = {{2{1'b0}}, col_in_359};
assign u_ca_in_360 = {{2{1'b0}}, col_in_360};
assign u_ca_in_361 = {{2{1'b0}}, col_in_361};
assign u_ca_in_362 = {{2{1'b0}}, col_in_362};
assign u_ca_in_363 = {{2{1'b0}}, col_in_363};
assign u_ca_in_364 = {{2{1'b0}}, col_in_364};
assign u_ca_in_365 = {{2{1'b0}}, col_in_365};
assign u_ca_in_366 = {{2{1'b0}}, col_in_366};
assign u_ca_in_367 = {{2{1'b0}}, col_in_367};
assign u_ca_in_368 = {{2{1'b0}}, col_in_368};
assign u_ca_in_369 = {{2{1'b0}}, col_in_369};
assign u_ca_in_370 = {{2{1'b0}}, col_in_370};
assign u_ca_in_371 = {{2{1'b0}}, col_in_371};
assign u_ca_in_372 = {{2{1'b0}}, col_in_372};
assign u_ca_in_373 = {{2{1'b0}}, col_in_373};
assign u_ca_in_374 = {{2{1'b0}}, col_in_374};
assign u_ca_in_375 = {{2{1'b0}}, col_in_375};
assign u_ca_in_376 = {{2{1'b0}}, col_in_376};
assign u_ca_in_377 = {{2{1'b0}}, col_in_377};
assign u_ca_in_378 = {{2{1'b0}}, col_in_378};
assign u_ca_in_379 = {{2{1'b0}}, col_in_379};
assign u_ca_in_380 = {{2{1'b0}}, col_in_380};
assign u_ca_in_381 = {{2{1'b0}}, col_in_381};
assign u_ca_in_382 = {{2{1'b0}}, col_in_382};
assign u_ca_in_383 = {{2{1'b0}}, col_in_383};
assign u_ca_in_384 = {{2{1'b0}}, col_in_384};
assign u_ca_in_385 = {{2{1'b0}}, col_in_385};
assign u_ca_in_386 = {{2{1'b0}}, col_in_386};
assign u_ca_in_387 = {{2{1'b0}}, col_in_387};
assign u_ca_in_388 = {{2{1'b0}}, col_in_388};
assign u_ca_in_389 = {{2{1'b0}}, col_in_389};
assign u_ca_in_390 = {{2{1'b0}}, col_in_390};
assign u_ca_in_391 = {{2{1'b0}}, col_in_391};
assign u_ca_in_392 = {{2{1'b0}}, col_in_392};
assign u_ca_in_393 = {{2{1'b0}}, col_in_393};
assign u_ca_in_394 = {{2{1'b0}}, col_in_394};
assign u_ca_in_395 = {{2{1'b0}}, col_in_395};
assign u_ca_in_396 = {{2{1'b0}}, col_in_396};
assign u_ca_in_397 = {{2{1'b0}}, col_in_397};
assign u_ca_in_398 = {{2{1'b0}}, col_in_398};
assign u_ca_in_399 = {{2{1'b0}}, col_in_399};
assign u_ca_in_400 = {{2{1'b0}}, col_in_400};
assign u_ca_in_401 = {{2{1'b0}}, col_in_401};
assign u_ca_in_402 = {{2{1'b0}}, col_in_402};
assign u_ca_in_403 = {{2{1'b0}}, col_in_403};
assign u_ca_in_404 = {{2{1'b0}}, col_in_404};
assign u_ca_in_405 = {{2{1'b0}}, col_in_405};
assign u_ca_in_406 = {{2{1'b0}}, col_in_406};
assign u_ca_in_407 = {{2{1'b0}}, col_in_407};
assign u_ca_in_408 = {{2{1'b0}}, col_in_408};
assign u_ca_in_409 = {{2{1'b0}}, col_in_409};
assign u_ca_in_410 = {{2{1'b0}}, col_in_410};
assign u_ca_in_411 = {{2{1'b0}}, col_in_411};
assign u_ca_in_412 = {{2{1'b0}}, col_in_412};
assign u_ca_in_413 = {{2{1'b0}}, col_in_413};
assign u_ca_in_414 = {{2{1'b0}}, col_in_414};
assign u_ca_in_415 = {{2{1'b0}}, col_in_415};
assign u_ca_in_416 = {{2{1'b0}}, col_in_416};
assign u_ca_in_417 = {{2{1'b0}}, col_in_417};
assign u_ca_in_418 = {{2{1'b0}}, col_in_418};
assign u_ca_in_419 = {{2{1'b0}}, col_in_419};
assign u_ca_in_420 = {{2{1'b0}}, col_in_420};
assign u_ca_in_421 = {{2{1'b0}}, col_in_421};
assign u_ca_in_422 = {{2{1'b0}}, col_in_422};
assign u_ca_in_423 = {{2{1'b0}}, col_in_423};
assign u_ca_in_424 = {{2{1'b0}}, col_in_424};
assign u_ca_in_425 = {{2{1'b0}}, col_in_425};
assign u_ca_in_426 = {{2{1'b0}}, col_in_426};
assign u_ca_in_427 = {{2{1'b0}}, col_in_427};
assign u_ca_in_428 = {{2{1'b0}}, col_in_428};
assign u_ca_in_429 = {{2{1'b0}}, col_in_429};
assign u_ca_in_430 = {{2{1'b0}}, col_in_430};
assign u_ca_in_431 = {{2{1'b0}}, col_in_431};
assign u_ca_in_432 = {{2{1'b0}}, col_in_432};
assign u_ca_in_433 = {{2{1'b0}}, col_in_433};
assign u_ca_in_434 = {{2{1'b0}}, col_in_434};
assign u_ca_in_435 = {{2{1'b0}}, col_in_435};
assign u_ca_in_436 = {{2{1'b0}}, col_in_436};
assign u_ca_in_437 = {{2{1'b0}}, col_in_437};
assign u_ca_in_438 = {{2{1'b0}}, col_in_438};
assign u_ca_in_439 = {{2{1'b0}}, col_in_439};
assign u_ca_in_440 = {{2{1'b0}}, col_in_440};
assign u_ca_in_441 = {{2{1'b0}}, col_in_441};
assign u_ca_in_442 = {{2{1'b0}}, col_in_442};
assign u_ca_in_443 = {{2{1'b0}}, col_in_443};
assign u_ca_in_444 = {{2{1'b0}}, col_in_444};
assign u_ca_in_445 = {{2{1'b0}}, col_in_445};
assign u_ca_in_446 = {{2{1'b0}}, col_in_446};
assign u_ca_in_447 = {{2{1'b0}}, col_in_447};
assign u_ca_in_448 = {{2{1'b0}}, col_in_448};
assign u_ca_in_449 = {{2{1'b0}}, col_in_449};
assign u_ca_in_450 = {{2{1'b0}}, col_in_450};
assign u_ca_in_451 = {{2{1'b0}}, col_in_451};
assign u_ca_in_452 = {{2{1'b0}}, col_in_452};
assign u_ca_in_453 = {{2{1'b0}}, col_in_453};
assign u_ca_in_454 = {{2{1'b0}}, col_in_454};
assign u_ca_in_455 = {{2{1'b0}}, col_in_455};
assign u_ca_in_456 = {{2{1'b0}}, col_in_456};
assign u_ca_in_457 = {{2{1'b0}}, col_in_457};
assign u_ca_in_458 = {{2{1'b0}}, col_in_458};
assign u_ca_in_459 = {{2{1'b0}}, col_in_459};
assign u_ca_in_460 = {{2{1'b0}}, col_in_460};
assign u_ca_in_461 = {{2{1'b0}}, col_in_461};
assign u_ca_in_462 = {{2{1'b0}}, col_in_462};
assign u_ca_in_463 = {{2{1'b0}}, col_in_463};
assign u_ca_in_464 = {{2{1'b0}}, col_in_464};
assign u_ca_in_465 = {{2{1'b0}}, col_in_465};
assign u_ca_in_466 = {{2{1'b0}}, col_in_466};
assign u_ca_in_467 = {{2{1'b0}}, col_in_467};
assign u_ca_in_468 = {{2{1'b0}}, col_in_468};
assign u_ca_in_469 = {{2{1'b0}}, col_in_469};
assign u_ca_in_470 = {{2{1'b0}}, col_in_470};
assign u_ca_in_471 = {{2{1'b0}}, col_in_471};
assign u_ca_in_472 = {{2{1'b0}}, col_in_472};
assign u_ca_in_473 = {{2{1'b0}}, col_in_473};
assign u_ca_in_474 = {{2{1'b0}}, col_in_474};
assign u_ca_in_475 = {{2{1'b0}}, col_in_475};
assign u_ca_in_476 = {{2{1'b0}}, col_in_476};
assign u_ca_in_477 = {{2{1'b0}}, col_in_477};
assign u_ca_in_478 = {{2{1'b0}}, col_in_478};
assign u_ca_in_479 = {{2{1'b0}}, col_in_479};
assign u_ca_in_480 = {{2{1'b0}}, col_in_480};
assign u_ca_in_481 = {{2{1'b0}}, col_in_481};
assign u_ca_in_482 = {{2{1'b0}}, col_in_482};
assign u_ca_in_483 = {{2{1'b0}}, col_in_483};
assign u_ca_in_484 = {{2{1'b0}}, col_in_484};
assign u_ca_in_485 = {{2{1'b0}}, col_in_485};
assign u_ca_in_486 = {{2{1'b0}}, col_in_486};
assign u_ca_in_487 = {{2{1'b0}}, col_in_487};
assign u_ca_in_488 = {{2{1'b0}}, col_in_488};
assign u_ca_in_489 = {{2{1'b0}}, col_in_489};
assign u_ca_in_490 = {{2{1'b0}}, col_in_490};
assign u_ca_in_491 = {{2{1'b0}}, col_in_491};
assign u_ca_in_492 = {{2{1'b0}}, col_in_492};
assign u_ca_in_493 = {{2{1'b0}}, col_in_493};
assign u_ca_in_494 = {{2{1'b0}}, col_in_494};
assign u_ca_in_495 = {{2{1'b0}}, col_in_495};
assign u_ca_in_496 = {{2{1'b0}}, col_in_496};
assign u_ca_in_497 = {{2{1'b0}}, col_in_497};
assign u_ca_in_498 = {{2{1'b0}}, col_in_498};
assign u_ca_in_499 = {{2{1'b0}}, col_in_499};
assign u_ca_in_500 = {{2{1'b0}}, col_in_500};
assign u_ca_in_501 = {{2{1'b0}}, col_in_501};
assign u_ca_in_502 = {{2{1'b0}}, col_in_502};
assign u_ca_in_503 = {{2{1'b0}}, col_in_503};
assign u_ca_in_504 = {{2{1'b0}}, col_in_504};
assign u_ca_in_505 = {{2{1'b0}}, col_in_505};
assign u_ca_in_506 = {{2{1'b0}}, col_in_506};
assign u_ca_in_507 = {{2{1'b0}}, col_in_507};
assign u_ca_in_508 = {{2{1'b0}}, col_in_508};
assign u_ca_in_509 = {{2{1'b0}}, col_in_509};
assign u_ca_in_510 = {{2{1'b0}}, col_in_510};
assign u_ca_in_511 = {{2{1'b0}}, col_in_511};
assign u_ca_in_512 = {{2{1'b0}}, col_in_512};
assign u_ca_in_513 = {{2{1'b0}}, col_in_513};
assign u_ca_in_514 = {{2{1'b0}}, col_in_514};
assign u_ca_in_515 = {{2{1'b0}}, col_in_515};
assign u_ca_in_516 = {{2{1'b0}}, col_in_516};
assign u_ca_in_517 = {{2{1'b0}}, col_in_517};
assign u_ca_in_518 = {{2{1'b0}}, col_in_518};
assign u_ca_in_519 = {{2{1'b0}}, col_in_519};
assign u_ca_in_520 = {{2{1'b0}}, col_in_520};
assign u_ca_in_521 = {{2{1'b0}}, col_in_521};
assign u_ca_in_522 = {{2{1'b0}}, col_in_522};
assign u_ca_in_523 = {{2{1'b0}}, col_in_523};
assign u_ca_in_524 = {{2{1'b0}}, col_in_524};
assign u_ca_in_525 = {{2{1'b0}}, col_in_525};
assign u_ca_in_526 = {{2{1'b0}}, col_in_526};
assign u_ca_in_527 = {{2{1'b0}}, col_in_527};
assign u_ca_in_528 = {{2{1'b0}}, col_in_528};
assign u_ca_in_529 = {{2{1'b0}}, col_in_529};
assign u_ca_in_530 = {{2{1'b0}}, col_in_530};
assign u_ca_in_531 = {{2{1'b0}}, col_in_531};
assign u_ca_in_532 = {{2{1'b0}}, col_in_532};
assign u_ca_in_533 = {{2{1'b0}}, col_in_533};
assign u_ca_in_534 = {{2{1'b0}}, col_in_534};
assign u_ca_in_535 = {{2{1'b0}}, col_in_535};
assign u_ca_in_536 = {{2{1'b0}}, col_in_536};
assign u_ca_in_537 = {{2{1'b0}}, col_in_537};
assign u_ca_in_538 = {{2{1'b0}}, col_in_538};
assign u_ca_in_539 = {{2{1'b0}}, col_in_539};
assign u_ca_in_540 = {{2{1'b0}}, col_in_540};
assign u_ca_in_541 = {{2{1'b0}}, col_in_541};
assign u_ca_in_542 = {{2{1'b0}}, col_in_542};
assign u_ca_in_543 = {{2{1'b0}}, col_in_543};
assign u_ca_in_544 = {{2{1'b0}}, col_in_544};
assign u_ca_in_545 = {{2{1'b0}}, col_in_545};
assign u_ca_in_546 = {{2{1'b0}}, col_in_546};
assign u_ca_in_547 = {{2{1'b0}}, col_in_547};
assign u_ca_in_548 = {{2{1'b0}}, col_in_548};
assign u_ca_in_549 = {{2{1'b0}}, col_in_549};
assign u_ca_in_550 = {{2{1'b0}}, col_in_550};
assign u_ca_in_551 = {{2{1'b0}}, col_in_551};
assign u_ca_in_552 = {{2{1'b0}}, col_in_552};
assign u_ca_in_553 = {{2{1'b0}}, col_in_553};
assign u_ca_in_554 = {{2{1'b0}}, col_in_554};
assign u_ca_in_555 = {{2{1'b0}}, col_in_555};
assign u_ca_in_556 = {{2{1'b0}}, col_in_556};
assign u_ca_in_557 = {{2{1'b0}}, col_in_557};
assign u_ca_in_558 = {{2{1'b0}}, col_in_558};
assign u_ca_in_559 = {{2{1'b0}}, col_in_559};
assign u_ca_in_560 = {{2{1'b0}}, col_in_560};
assign u_ca_in_561 = {{2{1'b0}}, col_in_561};
assign u_ca_in_562 = {{2{1'b0}}, col_in_562};
assign u_ca_in_563 = {{2{1'b0}}, col_in_563};
assign u_ca_in_564 = {{2{1'b0}}, col_in_564};
assign u_ca_in_565 = {{2{1'b0}}, col_in_565};
assign u_ca_in_566 = {{2{1'b0}}, col_in_566};
assign u_ca_in_567 = {{2{1'b0}}, col_in_567};
assign u_ca_in_568 = {{2{1'b0}}, col_in_568};
assign u_ca_in_569 = {{2{1'b0}}, col_in_569};
assign u_ca_in_570 = {{2{1'b0}}, col_in_570};
assign u_ca_in_571 = {{2{1'b0}}, col_in_571};
assign u_ca_in_572 = {{2{1'b0}}, col_in_572};
assign u_ca_in_573 = {{2{1'b0}}, col_in_573};
assign u_ca_in_574 = {{2{1'b0}}, col_in_574};
assign u_ca_in_575 = {{2{1'b0}}, col_in_575};
assign u_ca_in_576 = {{2{1'b0}}, col_in_576};
assign u_ca_in_577 = {{2{1'b0}}, col_in_577};
assign u_ca_in_578 = {{2{1'b0}}, col_in_578};
assign u_ca_in_579 = {{2{1'b0}}, col_in_579};
assign u_ca_in_580 = {{2{1'b0}}, col_in_580};
assign u_ca_in_581 = {{2{1'b0}}, col_in_581};
assign u_ca_in_582 = {{2{1'b0}}, col_in_582};
assign u_ca_in_583 = {{2{1'b0}}, col_in_583};
assign u_ca_in_584 = {{2{1'b0}}, col_in_584};
assign u_ca_in_585 = {{2{1'b0}}, col_in_585};
assign u_ca_in_586 = {{2{1'b0}}, col_in_586};
assign u_ca_in_587 = {{2{1'b0}}, col_in_587};
assign u_ca_in_588 = {{2{1'b0}}, col_in_588};
assign u_ca_in_589 = {{2{1'b0}}, col_in_589};
assign u_ca_in_590 = {{2{1'b0}}, col_in_590};
assign u_ca_in_591 = {{2{1'b0}}, col_in_591};
assign u_ca_in_592 = {{2{1'b0}}, col_in_592};
assign u_ca_in_593 = {{2{1'b0}}, col_in_593};
assign u_ca_in_594 = {{2{1'b0}}, col_in_594};
assign u_ca_in_595 = {{2{1'b0}}, col_in_595};
assign u_ca_in_596 = {{2{1'b0}}, col_in_596};
assign u_ca_in_597 = {{2{1'b0}}, col_in_597};
assign u_ca_in_598 = {{2{1'b0}}, col_in_598};
assign u_ca_in_599 = {{2{1'b0}}, col_in_599};
assign u_ca_in_600 = {{2{1'b0}}, col_in_600};
assign u_ca_in_601 = {{2{1'b0}}, col_in_601};
assign u_ca_in_602 = {{2{1'b0}}, col_in_602};
assign u_ca_in_603 = {{2{1'b0}}, col_in_603};
assign u_ca_in_604 = {{2{1'b0}}, col_in_604};
assign u_ca_in_605 = {{2{1'b0}}, col_in_605};
assign u_ca_in_606 = {{2{1'b0}}, col_in_606};
assign u_ca_in_607 = {{2{1'b0}}, col_in_607};
assign u_ca_in_608 = {{2{1'b0}}, col_in_608};
assign u_ca_in_609 = {{2{1'b0}}, col_in_609};
assign u_ca_in_610 = {{2{1'b0}}, col_in_610};
assign u_ca_in_611 = {{2{1'b0}}, col_in_611};
assign u_ca_in_612 = {{2{1'b0}}, col_in_612};
assign u_ca_in_613 = {{2{1'b0}}, col_in_613};
assign u_ca_in_614 = {{2{1'b0}}, col_in_614};
assign u_ca_in_615 = {{2{1'b0}}, col_in_615};
assign u_ca_in_616 = {{2{1'b0}}, col_in_616};
assign u_ca_in_617 = {{2{1'b0}}, col_in_617};
assign u_ca_in_618 = {{2{1'b0}}, col_in_618};
assign u_ca_in_619 = {{2{1'b0}}, col_in_619};
assign u_ca_in_620 = {{2{1'b0}}, col_in_620};
assign u_ca_in_621 = {{2{1'b0}}, col_in_621};
assign u_ca_in_622 = {{2{1'b0}}, col_in_622};
assign u_ca_in_623 = {{2{1'b0}}, col_in_623};
assign u_ca_in_624 = {{2{1'b0}}, col_in_624};
assign u_ca_in_625 = {{2{1'b0}}, col_in_625};
assign u_ca_in_626 = {{2{1'b0}}, col_in_626};
assign u_ca_in_627 = {{2{1'b0}}, col_in_627};
assign u_ca_in_628 = {{2{1'b0}}, col_in_628};
assign u_ca_in_629 = {{2{1'b0}}, col_in_629};
assign u_ca_in_630 = {{2{1'b0}}, col_in_630};
assign u_ca_in_631 = {{2{1'b0}}, col_in_631};
assign u_ca_in_632 = {{2{1'b0}}, col_in_632};
assign u_ca_in_633 = {{2{1'b0}}, col_in_633};
assign u_ca_in_634 = {{2{1'b0}}, col_in_634};
assign u_ca_in_635 = {{2{1'b0}}, col_in_635};
assign u_ca_in_636 = {{2{1'b0}}, col_in_636};
assign u_ca_in_637 = {{2{1'b0}}, col_in_637};
assign u_ca_in_638 = {{2{1'b0}}, col_in_638};
assign u_ca_in_639 = {{2{1'b0}}, col_in_639};
assign u_ca_in_640 = {{2{1'b0}}, col_in_640};
assign u_ca_in_641 = {{2{1'b0}}, col_in_641};
assign u_ca_in_642 = {{2{1'b0}}, col_in_642};
assign u_ca_in_643 = {{2{1'b0}}, col_in_643};
assign u_ca_in_644 = {{2{1'b0}}, col_in_644};
assign u_ca_in_645 = {{2{1'b0}}, col_in_645};
assign u_ca_in_646 = {{2{1'b0}}, col_in_646};
assign u_ca_in_647 = {{2{1'b0}}, col_in_647};
assign u_ca_in_648 = {{2{1'b0}}, col_in_648};
assign u_ca_in_649 = {{2{1'b0}}, col_in_649};
assign u_ca_in_650 = {{2{1'b0}}, col_in_650};
assign u_ca_in_651 = {{2{1'b0}}, col_in_651};
assign u_ca_in_652 = {{2{1'b0}}, col_in_652};
assign u_ca_in_653 = {{2{1'b0}}, col_in_653};
assign u_ca_in_654 = {{2{1'b0}}, col_in_654};
assign u_ca_in_655 = {{2{1'b0}}, col_in_655};
assign u_ca_in_656 = {{2{1'b0}}, col_in_656};
assign u_ca_in_657 = {{2{1'b0}}, col_in_657};
assign u_ca_in_658 = {{2{1'b0}}, col_in_658};
assign u_ca_in_659 = {{2{1'b0}}, col_in_659};
assign u_ca_in_660 = {{2{1'b0}}, col_in_660};
assign u_ca_in_661 = {{2{1'b0}}, col_in_661};
assign u_ca_in_662 = {{2{1'b0}}, col_in_662};
assign u_ca_in_663 = {{2{1'b0}}, col_in_663};
assign u_ca_in_664 = {{2{1'b0}}, col_in_664};
assign u_ca_in_665 = {{2{1'b0}}, col_in_665};
assign u_ca_in_666 = {{2{1'b0}}, col_in_666};
assign u_ca_in_667 = {{2{1'b0}}, col_in_667};
assign u_ca_in_668 = {{2{1'b0}}, col_in_668};
assign u_ca_in_669 = {{2{1'b0}}, col_in_669};
assign u_ca_in_670 = {{2{1'b0}}, col_in_670};
assign u_ca_in_671 = {{2{1'b0}}, col_in_671};
assign u_ca_in_672 = {{2{1'b0}}, col_in_672};
assign u_ca_in_673 = {{2{1'b0}}, col_in_673};
assign u_ca_in_674 = {{2{1'b0}}, col_in_674};
assign u_ca_in_675 = {{2{1'b0}}, col_in_675};
assign u_ca_in_676 = {{2{1'b0}}, col_in_676};
assign u_ca_in_677 = {{2{1'b0}}, col_in_677};
assign u_ca_in_678 = {{2{1'b0}}, col_in_678};
assign u_ca_in_679 = {{2{1'b0}}, col_in_679};
assign u_ca_in_680 = {{2{1'b0}}, col_in_680};
assign u_ca_in_681 = {{2{1'b0}}, col_in_681};
assign u_ca_in_682 = {{2{1'b0}}, col_in_682};
assign u_ca_in_683 = {{2{1'b0}}, col_in_683};
assign u_ca_in_684 = {{2{1'b0}}, col_in_684};
assign u_ca_in_685 = {{2{1'b0}}, col_in_685};
assign u_ca_in_686 = {{2{1'b0}}, col_in_686};
assign u_ca_in_687 = {{2{1'b0}}, col_in_687};
assign u_ca_in_688 = {{2{1'b0}}, col_in_688};
assign u_ca_in_689 = {{2{1'b0}}, col_in_689};
assign u_ca_in_690 = {{2{1'b0}}, col_in_690};
assign u_ca_in_691 = {{2{1'b0}}, col_in_691};
assign u_ca_in_692 = {{2{1'b0}}, col_in_692};
assign u_ca_in_693 = {{2{1'b0}}, col_in_693};
assign u_ca_in_694 = {{2{1'b0}}, col_in_694};
assign u_ca_in_695 = {{2{1'b0}}, col_in_695};
assign u_ca_in_696 = {{2{1'b0}}, col_in_696};
assign u_ca_in_697 = {{2{1'b0}}, col_in_697};
assign u_ca_in_698 = {{2{1'b0}}, col_in_698};
assign u_ca_in_699 = {{2{1'b0}}, col_in_699};
assign u_ca_in_700 = {{2{1'b0}}, col_in_700};
assign u_ca_in_701 = {{2{1'b0}}, col_in_701};
assign u_ca_in_702 = {{2{1'b0}}, col_in_702};
assign u_ca_in_703 = {{2{1'b0}}, col_in_703};
assign u_ca_in_704 = {{2{1'b0}}, col_in_704};
assign u_ca_in_705 = {{2{1'b0}}, col_in_705};
assign u_ca_in_706 = {{2{1'b0}}, col_in_706};
assign u_ca_in_707 = {{2{1'b0}}, col_in_707};
assign u_ca_in_708 = {{2{1'b0}}, col_in_708};
assign u_ca_in_709 = {{2{1'b0}}, col_in_709};
assign u_ca_in_710 = {{2{1'b0}}, col_in_710};
assign u_ca_in_711 = {{2{1'b0}}, col_in_711};
assign u_ca_in_712 = {{2{1'b0}}, col_in_712};
assign u_ca_in_713 = {{2{1'b0}}, col_in_713};
assign u_ca_in_714 = {{2{1'b0}}, col_in_714};
assign u_ca_in_715 = {{2{1'b0}}, col_in_715};
assign u_ca_in_716 = {{2{1'b0}}, col_in_716};
assign u_ca_in_717 = {{2{1'b0}}, col_in_717};
assign u_ca_in_718 = {{2{1'b0}}, col_in_718};
assign u_ca_in_719 = {{2{1'b0}}, col_in_719};
assign u_ca_in_720 = {{2{1'b0}}, col_in_720};
assign u_ca_in_721 = {{2{1'b0}}, col_in_721};
assign u_ca_in_722 = {{2{1'b0}}, col_in_722};
assign u_ca_in_723 = {{2{1'b0}}, col_in_723};
assign u_ca_in_724 = {{2{1'b0}}, col_in_724};
assign u_ca_in_725 = {{2{1'b0}}, col_in_725};
assign u_ca_in_726 = {{2{1'b0}}, col_in_726};
assign u_ca_in_727 = {{2{1'b0}}, col_in_727};
assign u_ca_in_728 = {{2{1'b0}}, col_in_728};
assign u_ca_in_729 = {{2{1'b0}}, col_in_729};
assign u_ca_in_730 = {{2{1'b0}}, col_in_730};
assign u_ca_in_731 = {{2{1'b0}}, col_in_731};
assign u_ca_in_732 = {{2{1'b0}}, col_in_732};
assign u_ca_in_733 = {{2{1'b0}}, col_in_733};
assign u_ca_in_734 = {{2{1'b0}}, col_in_734};
assign u_ca_in_735 = {{2{1'b0}}, col_in_735};
assign u_ca_in_736 = {{2{1'b0}}, col_in_736};
assign u_ca_in_737 = {{2{1'b0}}, col_in_737};
assign u_ca_in_738 = {{2{1'b0}}, col_in_738};
assign u_ca_in_739 = {{2{1'b0}}, col_in_739};
assign u_ca_in_740 = {{2{1'b0}}, col_in_740};
assign u_ca_in_741 = {{2{1'b0}}, col_in_741};
assign u_ca_in_742 = {{2{1'b0}}, col_in_742};
assign u_ca_in_743 = {{2{1'b0}}, col_in_743};
assign u_ca_in_744 = {{2{1'b0}}, col_in_744};
assign u_ca_in_745 = {{2{1'b0}}, col_in_745};
assign u_ca_in_746 = {{2{1'b0}}, col_in_746};
assign u_ca_in_747 = {{2{1'b0}}, col_in_747};
assign u_ca_in_748 = {{2{1'b0}}, col_in_748};
assign u_ca_in_749 = {{2{1'b0}}, col_in_749};
assign u_ca_in_750 = {{2{1'b0}}, col_in_750};
assign u_ca_in_751 = {{2{1'b0}}, col_in_751};
assign u_ca_in_752 = {{2{1'b0}}, col_in_752};
assign u_ca_in_753 = {{2{1'b0}}, col_in_753};
assign u_ca_in_754 = {{2{1'b0}}, col_in_754};
assign u_ca_in_755 = {{2{1'b0}}, col_in_755};
assign u_ca_in_756 = {{2{1'b0}}, col_in_756};
assign u_ca_in_757 = {{2{1'b0}}, col_in_757};
assign u_ca_in_758 = {{2{1'b0}}, col_in_758};
assign u_ca_in_759 = {{2{1'b0}}, col_in_759};
assign u_ca_in_760 = {{2{1'b0}}, col_in_760};
assign u_ca_in_761 = {{2{1'b0}}, col_in_761};
assign u_ca_in_762 = {{2{1'b0}}, col_in_762};
assign u_ca_in_763 = {{2{1'b0}}, col_in_763};
assign u_ca_in_764 = {{2{1'b0}}, col_in_764};
assign u_ca_in_765 = {{2{1'b0}}, col_in_765};
assign u_ca_in_766 = {{2{1'b0}}, col_in_766};
assign u_ca_in_767 = {{2{1'b0}}, col_in_767};
assign u_ca_in_768 = {{2{1'b0}}, col_in_768};
assign u_ca_in_769 = {{2{1'b0}}, col_in_769};
assign u_ca_in_770 = {{2{1'b0}}, col_in_770};
assign u_ca_in_771 = {{2{1'b0}}, col_in_771};
assign u_ca_in_772 = {{2{1'b0}}, col_in_772};
assign u_ca_in_773 = {{2{1'b0}}, col_in_773};
assign u_ca_in_774 = {{2{1'b0}}, col_in_774};
assign u_ca_in_775 = {{2{1'b0}}, col_in_775};
assign u_ca_in_776 = {{2{1'b0}}, col_in_776};
assign u_ca_in_777 = {{2{1'b0}}, col_in_777};
assign u_ca_in_778 = {{2{1'b0}}, col_in_778};
assign u_ca_in_779 = {{2{1'b0}}, col_in_779};
assign u_ca_in_780 = {{2{1'b0}}, col_in_780};
assign u_ca_in_781 = {{2{1'b0}}, col_in_781};
assign u_ca_in_782 = {{2{1'b0}}, col_in_782};
assign u_ca_in_783 = {{2{1'b0}}, col_in_783};
assign u_ca_in_784 = {{2{1'b0}}, col_in_784};
assign u_ca_in_785 = {{2{1'b0}}, col_in_785};
assign u_ca_in_786 = {{2{1'b0}}, col_in_786};
assign u_ca_in_787 = {{2{1'b0}}, col_in_787};
assign u_ca_in_788 = {{2{1'b0}}, col_in_788};
assign u_ca_in_789 = {{2{1'b0}}, col_in_789};
assign u_ca_in_790 = {{2{1'b0}}, col_in_790};
assign u_ca_in_791 = {{2{1'b0}}, col_in_791};
assign u_ca_in_792 = {{2{1'b0}}, col_in_792};
assign u_ca_in_793 = {{2{1'b0}}, col_in_793};
assign u_ca_in_794 = {{2{1'b0}}, col_in_794};
assign u_ca_in_795 = {{2{1'b0}}, col_in_795};
assign u_ca_in_796 = {{2{1'b0}}, col_in_796};
assign u_ca_in_797 = {{2{1'b0}}, col_in_797};
assign u_ca_in_798 = {{2{1'b0}}, col_in_798};
assign u_ca_in_799 = {{2{1'b0}}, col_in_799};
assign u_ca_in_800 = {{2{1'b0}}, col_in_800};
assign u_ca_in_801 = {{2{1'b0}}, col_in_801};
assign u_ca_in_802 = {{2{1'b0}}, col_in_802};
assign u_ca_in_803 = {{2{1'b0}}, col_in_803};
assign u_ca_in_804 = {{2{1'b0}}, col_in_804};
assign u_ca_in_805 = {{2{1'b0}}, col_in_805};
assign u_ca_in_806 = {{2{1'b0}}, col_in_806};
assign u_ca_in_807 = {{2{1'b0}}, col_in_807};
assign u_ca_in_808 = {{2{1'b0}}, col_in_808};
assign u_ca_in_809 = {{2{1'b0}}, col_in_809};
assign u_ca_in_810 = {{2{1'b0}}, col_in_810};
assign u_ca_in_811 = {{2{1'b0}}, col_in_811};
assign u_ca_in_812 = {{2{1'b0}}, col_in_812};
assign u_ca_in_813 = {{2{1'b0}}, col_in_813};
assign u_ca_in_814 = {{2{1'b0}}, col_in_814};
assign u_ca_in_815 = {{2{1'b0}}, col_in_815};
assign u_ca_in_816 = {{2{1'b0}}, col_in_816};
assign u_ca_in_817 = {{2{1'b0}}, col_in_817};
assign u_ca_in_818 = {{2{1'b0}}, col_in_818};
assign u_ca_in_819 = {{2{1'b0}}, col_in_819};
assign u_ca_in_820 = {{2{1'b0}}, col_in_820};
assign u_ca_in_821 = {{2{1'b0}}, col_in_821};
assign u_ca_in_822 = {{2{1'b0}}, col_in_822};
assign u_ca_in_823 = {{2{1'b0}}, col_in_823};
assign u_ca_in_824 = {{2{1'b0}}, col_in_824};
assign u_ca_in_825 = {{2{1'b0}}, col_in_825};
assign u_ca_in_826 = {{2{1'b0}}, col_in_826};
assign u_ca_in_827 = {{2{1'b0}}, col_in_827};
assign u_ca_in_828 = {{2{1'b0}}, col_in_828};
assign u_ca_in_829 = {{2{1'b0}}, col_in_829};
assign u_ca_in_830 = {{2{1'b0}}, col_in_830};
assign u_ca_in_831 = {{2{1'b0}}, col_in_831};
assign u_ca_in_832 = {{2{1'b0}}, col_in_832};
assign u_ca_in_833 = {{2{1'b0}}, col_in_833};
assign u_ca_in_834 = {{2{1'b0}}, col_in_834};
assign u_ca_in_835 = {{2{1'b0}}, col_in_835};
assign u_ca_in_836 = {{2{1'b0}}, col_in_836};
assign u_ca_in_837 = {{2{1'b0}}, col_in_837};
assign u_ca_in_838 = {{2{1'b0}}, col_in_838};
assign u_ca_in_839 = {{2{1'b0}}, col_in_839};
assign u_ca_in_840 = {{2{1'b0}}, col_in_840};
assign u_ca_in_841 = {{2{1'b0}}, col_in_841};
assign u_ca_in_842 = {{2{1'b0}}, col_in_842};
assign u_ca_in_843 = {{2{1'b0}}, col_in_843};
assign u_ca_in_844 = {{2{1'b0}}, col_in_844};
assign u_ca_in_845 = {{2{1'b0}}, col_in_845};
assign u_ca_in_846 = {{2{1'b0}}, col_in_846};
assign u_ca_in_847 = {{2{1'b0}}, col_in_847};
assign u_ca_in_848 = {{2{1'b0}}, col_in_848};
assign u_ca_in_849 = {{2{1'b0}}, col_in_849};
assign u_ca_in_850 = {{2{1'b0}}, col_in_850};
assign u_ca_in_851 = {{2{1'b0}}, col_in_851};
assign u_ca_in_852 = {{2{1'b0}}, col_in_852};
assign u_ca_in_853 = {{2{1'b0}}, col_in_853};
assign u_ca_in_854 = {{2{1'b0}}, col_in_854};
assign u_ca_in_855 = {{2{1'b0}}, col_in_855};
assign u_ca_in_856 = {{2{1'b0}}, col_in_856};
assign u_ca_in_857 = {{2{1'b0}}, col_in_857};
assign u_ca_in_858 = {{2{1'b0}}, col_in_858};
assign u_ca_in_859 = {{2{1'b0}}, col_in_859};
assign u_ca_in_860 = {{2{1'b0}}, col_in_860};
assign u_ca_in_861 = {{2{1'b0}}, col_in_861};
assign u_ca_in_862 = {{2{1'b0}}, col_in_862};
assign u_ca_in_863 = {{2{1'b0}}, col_in_863};
assign u_ca_in_864 = {{2{1'b0}}, col_in_864};
assign u_ca_in_865 = {{2{1'b0}}, col_in_865};
assign u_ca_in_866 = {{2{1'b0}}, col_in_866};
assign u_ca_in_867 = {{2{1'b0}}, col_in_867};
assign u_ca_in_868 = {{2{1'b0}}, col_in_868};
assign u_ca_in_869 = {{2{1'b0}}, col_in_869};
assign u_ca_in_870 = {{2{1'b0}}, col_in_870};
assign u_ca_in_871 = {{2{1'b0}}, col_in_871};
assign u_ca_in_872 = {{2{1'b0}}, col_in_872};
assign u_ca_in_873 = {{2{1'b0}}, col_in_873};
assign u_ca_in_874 = {{2{1'b0}}, col_in_874};
assign u_ca_in_875 = {{2{1'b0}}, col_in_875};
assign u_ca_in_876 = {{2{1'b0}}, col_in_876};
assign u_ca_in_877 = {{2{1'b0}}, col_in_877};
assign u_ca_in_878 = {{2{1'b0}}, col_in_878};
assign u_ca_in_879 = {{2{1'b0}}, col_in_879};
assign u_ca_in_880 = {{2{1'b0}}, col_in_880};
assign u_ca_in_881 = {{2{1'b0}}, col_in_881};
assign u_ca_in_882 = {{2{1'b0}}, col_in_882};
assign u_ca_in_883 = {{2{1'b0}}, col_in_883};
assign u_ca_in_884 = {{2{1'b0}}, col_in_884};
assign u_ca_in_885 = {{2{1'b0}}, col_in_885};
assign u_ca_in_886 = {{2{1'b0}}, col_in_886};
assign u_ca_in_887 = {{2{1'b0}}, col_in_887};
assign u_ca_in_888 = {{2{1'b0}}, col_in_888};
assign u_ca_in_889 = {{2{1'b0}}, col_in_889};
assign u_ca_in_890 = {{2{1'b0}}, col_in_890};
assign u_ca_in_891 = {{2{1'b0}}, col_in_891};
assign u_ca_in_892 = {{2{1'b0}}, col_in_892};
assign u_ca_in_893 = {{2{1'b0}}, col_in_893};
assign u_ca_in_894 = {{2{1'b0}}, col_in_894};
assign u_ca_in_895 = {{2{1'b0}}, col_in_895};
assign u_ca_in_896 = {{2{1'b0}}, col_in_896};
assign u_ca_in_897 = {{2{1'b0}}, col_in_897};
assign u_ca_in_898 = {{2{1'b0}}, col_in_898};
assign u_ca_in_899 = {{2{1'b0}}, col_in_899};
assign u_ca_in_900 = {{2{1'b0}}, col_in_900};
assign u_ca_in_901 = {{2{1'b0}}, col_in_901};
assign u_ca_in_902 = {{2{1'b0}}, col_in_902};
assign u_ca_in_903 = {{2{1'b0}}, col_in_903};
assign u_ca_in_904 = {{2{1'b0}}, col_in_904};
assign u_ca_in_905 = {{2{1'b0}}, col_in_905};
assign u_ca_in_906 = {{2{1'b0}}, col_in_906};
assign u_ca_in_907 = {{2{1'b0}}, col_in_907};
assign u_ca_in_908 = {{2{1'b0}}, col_in_908};
assign u_ca_in_909 = {{2{1'b0}}, col_in_909};
assign u_ca_in_910 = {{2{1'b0}}, col_in_910};
assign u_ca_in_911 = {{2{1'b0}}, col_in_911};
assign u_ca_in_912 = {{2{1'b0}}, col_in_912};
assign u_ca_in_913 = {{2{1'b0}}, col_in_913};
assign u_ca_in_914 = {{2{1'b0}}, col_in_914};
assign u_ca_in_915 = {{2{1'b0}}, col_in_915};
assign u_ca_in_916 = {{2{1'b0}}, col_in_916};
assign u_ca_in_917 = {{2{1'b0}}, col_in_917};
assign u_ca_in_918 = {{2{1'b0}}, col_in_918};
assign u_ca_in_919 = {{2{1'b0}}, col_in_919};
assign u_ca_in_920 = {{2{1'b0}}, col_in_920};
assign u_ca_in_921 = {{2{1'b0}}, col_in_921};
assign u_ca_in_922 = {{2{1'b0}}, col_in_922};
assign u_ca_in_923 = {{2{1'b0}}, col_in_923};
assign u_ca_in_924 = {{2{1'b0}}, col_in_924};
assign u_ca_in_925 = {{2{1'b0}}, col_in_925};
assign u_ca_in_926 = {{2{1'b0}}, col_in_926};
assign u_ca_in_927 = {{2{1'b0}}, col_in_927};
assign u_ca_in_928 = {{2{1'b0}}, col_in_928};
assign u_ca_in_929 = {{2{1'b0}}, col_in_929};
assign u_ca_in_930 = {{2{1'b0}}, col_in_930};
assign u_ca_in_931 = {{2{1'b0}}, col_in_931};
assign u_ca_in_932 = {{2{1'b0}}, col_in_932};
assign u_ca_in_933 = {{2{1'b0}}, col_in_933};
assign u_ca_in_934 = {{2{1'b0}}, col_in_934};
assign u_ca_in_935 = {{2{1'b0}}, col_in_935};
assign u_ca_in_936 = {{2{1'b0}}, col_in_936};
assign u_ca_in_937 = {{2{1'b0}}, col_in_937};
assign u_ca_in_938 = {{2{1'b0}}, col_in_938};
assign u_ca_in_939 = {{2{1'b0}}, col_in_939};
assign u_ca_in_940 = {{2{1'b0}}, col_in_940};
assign u_ca_in_941 = {{2{1'b0}}, col_in_941};
assign u_ca_in_942 = {{2{1'b0}}, col_in_942};
assign u_ca_in_943 = {{2{1'b0}}, col_in_943};
assign u_ca_in_944 = {{2{1'b0}}, col_in_944};
assign u_ca_in_945 = {{2{1'b0}}, col_in_945};
assign u_ca_in_946 = {{2{1'b0}}, col_in_946};
assign u_ca_in_947 = {{2{1'b0}}, col_in_947};
assign u_ca_in_948 = {{2{1'b0}}, col_in_948};
assign u_ca_in_949 = {{2{1'b0}}, col_in_949};
assign u_ca_in_950 = {{2{1'b0}}, col_in_950};
assign u_ca_in_951 = {{2{1'b0}}, col_in_951};
assign u_ca_in_952 = {{2{1'b0}}, col_in_952};
assign u_ca_in_953 = {{2{1'b0}}, col_in_953};
assign u_ca_in_954 = {{2{1'b0}}, col_in_954};
assign u_ca_in_955 = {{2{1'b0}}, col_in_955};
assign u_ca_in_956 = {{2{1'b0}}, col_in_956};
assign u_ca_in_957 = {{2{1'b0}}, col_in_957};
assign u_ca_in_958 = {{2{1'b0}}, col_in_958};
assign u_ca_in_959 = {{2{1'b0}}, col_in_959};
assign u_ca_in_960 = {{2{1'b0}}, col_in_960};
assign u_ca_in_961 = {{2{1'b0}}, col_in_961};
assign u_ca_in_962 = {{2{1'b0}}, col_in_962};
assign u_ca_in_963 = {{2{1'b0}}, col_in_963};
assign u_ca_in_964 = {{2{1'b0}}, col_in_964};
assign u_ca_in_965 = {{2{1'b0}}, col_in_965};
assign u_ca_in_966 = {{2{1'b0}}, col_in_966};
assign u_ca_in_967 = {{2{1'b0}}, col_in_967};
assign u_ca_in_968 = {{2{1'b0}}, col_in_968};
assign u_ca_in_969 = {{2{1'b0}}, col_in_969};
assign u_ca_in_970 = {{2{1'b0}}, col_in_970};
assign u_ca_in_971 = {{2{1'b0}}, col_in_971};
assign u_ca_in_972 = {{2{1'b0}}, col_in_972};
assign u_ca_in_973 = {{2{1'b0}}, col_in_973};
assign u_ca_in_974 = {{2{1'b0}}, col_in_974};
assign u_ca_in_975 = {{2{1'b0}}, col_in_975};
assign u_ca_in_976 = {{2{1'b0}}, col_in_976};
assign u_ca_in_977 = {{2{1'b0}}, col_in_977};
assign u_ca_in_978 = {{2{1'b0}}, col_in_978};
assign u_ca_in_979 = {{2{1'b0}}, col_in_979};
assign u_ca_in_980 = {{2{1'b0}}, col_in_980};
assign u_ca_in_981 = {{2{1'b0}}, col_in_981};
assign u_ca_in_982 = {{2{1'b0}}, col_in_982};
assign u_ca_in_983 = {{2{1'b0}}, col_in_983};
assign u_ca_in_984 = {{2{1'b0}}, col_in_984};
assign u_ca_in_985 = {{2{1'b0}}, col_in_985};
assign u_ca_in_986 = {{2{1'b0}}, col_in_986};
assign u_ca_in_987 = {{2{1'b0}}, col_in_987};
assign u_ca_in_988 = {{2{1'b0}}, col_in_988};
assign u_ca_in_989 = {{2{1'b0}}, col_in_989};
assign u_ca_in_990 = {{2{1'b0}}, col_in_990};
assign u_ca_in_991 = {{2{1'b0}}, col_in_991};
assign u_ca_in_992 = {{2{1'b0}}, col_in_992};
assign u_ca_in_993 = {{2{1'b0}}, col_in_993};
assign u_ca_in_994 = {{2{1'b0}}, col_in_994};
assign u_ca_in_995 = {{2{1'b0}}, col_in_995};
assign u_ca_in_996 = {{2{1'b0}}, col_in_996};
assign u_ca_in_997 = {{2{1'b0}}, col_in_997};
assign u_ca_in_998 = {{2{1'b0}}, col_in_998};
assign u_ca_in_999 = {{2{1'b0}}, col_in_999};
assign u_ca_in_1000 = {{2{1'b0}}, col_in_1000};
assign u_ca_in_1001 = {{2{1'b0}}, col_in_1001};
assign u_ca_in_1002 = {{2{1'b0}}, col_in_1002};
assign u_ca_in_1003 = {{2{1'b0}}, col_in_1003};
assign u_ca_in_1004 = {{2{1'b0}}, col_in_1004};
assign u_ca_in_1005 = {{2{1'b0}}, col_in_1005};
assign u_ca_in_1006 = {{2{1'b0}}, col_in_1006};
assign u_ca_in_1007 = {{2{1'b0}}, col_in_1007};
assign u_ca_in_1008 = {{2{1'b0}}, col_in_1008};
assign u_ca_in_1009 = {{2{1'b0}}, col_in_1009};
assign u_ca_in_1010 = {{2{1'b0}}, col_in_1010};
assign u_ca_in_1011 = {{2{1'b0}}, col_in_1011};
assign u_ca_in_1012 = {{2{1'b0}}, col_in_1012};
assign u_ca_in_1013 = {{2{1'b0}}, col_in_1013};
assign u_ca_in_1014 = {{2{1'b0}}, col_in_1014};
assign u_ca_in_1015 = {{2{1'b0}}, col_in_1015};
assign u_ca_in_1016 = {{2{1'b0}}, col_in_1016};
assign u_ca_in_1017 = {{2{1'b0}}, col_in_1017};
assign u_ca_in_1018 = {{2{1'b0}}, col_in_1018};
assign u_ca_in_1019 = {{2{1'b0}}, col_in_1019};
assign u_ca_in_1020 = {{2{1'b0}}, col_in_1020};
assign u_ca_in_1021 = {{2{1'b0}}, col_in_1021};
assign u_ca_in_1022 = {{2{1'b0}}, col_in_1022};
assign u_ca_in_1023 = {{2{1'b0}}, col_in_1023};
assign u_ca_in_1024 = {{2{1'b0}}, col_in_1024};
assign u_ca_in_1025 = {{2{1'b0}}, col_in_1025};
assign u_ca_in_1026 = {{2{1'b0}}, col_in_1026};
assign u_ca_in_1027 = {{2{1'b0}}, col_in_1027};
assign u_ca_in_1028 = {{2{1'b0}}, col_in_1028};
assign u_ca_in_1029 = {{2{1'b0}}, col_in_1029};
assign u_ca_in_1030 = {{2{1'b0}}, col_in_1030};
assign u_ca_in_1031 = {{2{1'b0}}, col_in_1031};
assign u_ca_in_1032 = {{2{1'b0}}, col_in_1032};

//---------------------------------------------------------



//--compressor_array---------------------------------------
compressor_18_12 u_ca_18_12_0(.d_in(u_ca_in_0), .d_out(u_ca_out_0));
compressor_18_12 u_ca_18_12_1(.d_in(u_ca_in_1), .d_out(u_ca_out_1));
compressor_18_12 u_ca_18_12_2(.d_in(u_ca_in_2), .d_out(u_ca_out_2));
compressor_18_12 u_ca_18_12_3(.d_in(u_ca_in_3), .d_out(u_ca_out_3));
compressor_18_12 u_ca_18_12_4(.d_in(u_ca_in_4), .d_out(u_ca_out_4));
compressor_18_12 u_ca_18_12_5(.d_in(u_ca_in_5), .d_out(u_ca_out_5));
compressor_18_12 u_ca_18_12_6(.d_in(u_ca_in_6), .d_out(u_ca_out_6));
compressor_18_12 u_ca_18_12_7(.d_in(u_ca_in_7), .d_out(u_ca_out_7));
compressor_18_12 u_ca_18_12_8(.d_in(u_ca_in_8), .d_out(u_ca_out_8));
compressor_18_12 u_ca_18_12_9(.d_in(u_ca_in_9), .d_out(u_ca_out_9));
compressor_18_12 u_ca_18_12_10(.d_in(u_ca_in_10), .d_out(u_ca_out_10));
compressor_18_12 u_ca_18_12_11(.d_in(u_ca_in_11), .d_out(u_ca_out_11));
compressor_18_12 u_ca_18_12_12(.d_in(u_ca_in_12), .d_out(u_ca_out_12));
compressor_18_12 u_ca_18_12_13(.d_in(u_ca_in_13), .d_out(u_ca_out_13));
compressor_18_12 u_ca_18_12_14(.d_in(u_ca_in_14), .d_out(u_ca_out_14));
compressor_18_12 u_ca_18_12_15(.d_in(u_ca_in_15), .d_out(u_ca_out_15));
compressor_18_12 u_ca_18_12_16(.d_in(u_ca_in_16), .d_out(u_ca_out_16));
compressor_18_12 u_ca_18_12_17(.d_in(u_ca_in_17), .d_out(u_ca_out_17));
compressor_18_12 u_ca_18_12_18(.d_in(u_ca_in_18), .d_out(u_ca_out_18));
compressor_18_12 u_ca_18_12_19(.d_in(u_ca_in_19), .d_out(u_ca_out_19));
compressor_18_12 u_ca_18_12_20(.d_in(u_ca_in_20), .d_out(u_ca_out_20));
compressor_18_12 u_ca_18_12_21(.d_in(u_ca_in_21), .d_out(u_ca_out_21));
compressor_18_12 u_ca_18_12_22(.d_in(u_ca_in_22), .d_out(u_ca_out_22));
compressor_18_12 u_ca_18_12_23(.d_in(u_ca_in_23), .d_out(u_ca_out_23));
compressor_18_12 u_ca_18_12_24(.d_in(u_ca_in_24), .d_out(u_ca_out_24));
compressor_18_12 u_ca_18_12_25(.d_in(u_ca_in_25), .d_out(u_ca_out_25));
compressor_18_12 u_ca_18_12_26(.d_in(u_ca_in_26), .d_out(u_ca_out_26));
compressor_18_12 u_ca_18_12_27(.d_in(u_ca_in_27), .d_out(u_ca_out_27));
compressor_18_12 u_ca_18_12_28(.d_in(u_ca_in_28), .d_out(u_ca_out_28));
compressor_18_12 u_ca_18_12_29(.d_in(u_ca_in_29), .d_out(u_ca_out_29));
compressor_18_12 u_ca_18_12_30(.d_in(u_ca_in_30), .d_out(u_ca_out_30));
compressor_18_12 u_ca_18_12_31(.d_in(u_ca_in_31), .d_out(u_ca_out_31));
compressor_18_12 u_ca_18_12_32(.d_in(u_ca_in_32), .d_out(u_ca_out_32));
compressor_18_12 u_ca_18_12_33(.d_in(u_ca_in_33), .d_out(u_ca_out_33));
compressor_18_12 u_ca_18_12_34(.d_in(u_ca_in_34), .d_out(u_ca_out_34));
compressor_18_12 u_ca_18_12_35(.d_in(u_ca_in_35), .d_out(u_ca_out_35));
compressor_18_12 u_ca_18_12_36(.d_in(u_ca_in_36), .d_out(u_ca_out_36));
compressor_18_12 u_ca_18_12_37(.d_in(u_ca_in_37), .d_out(u_ca_out_37));
compressor_18_12 u_ca_18_12_38(.d_in(u_ca_in_38), .d_out(u_ca_out_38));
compressor_18_12 u_ca_18_12_39(.d_in(u_ca_in_39), .d_out(u_ca_out_39));
compressor_18_12 u_ca_18_12_40(.d_in(u_ca_in_40), .d_out(u_ca_out_40));
compressor_18_12 u_ca_18_12_41(.d_in(u_ca_in_41), .d_out(u_ca_out_41));
compressor_18_12 u_ca_18_12_42(.d_in(u_ca_in_42), .d_out(u_ca_out_42));
compressor_18_12 u_ca_18_12_43(.d_in(u_ca_in_43), .d_out(u_ca_out_43));
compressor_18_12 u_ca_18_12_44(.d_in(u_ca_in_44), .d_out(u_ca_out_44));
compressor_18_12 u_ca_18_12_45(.d_in(u_ca_in_45), .d_out(u_ca_out_45));
compressor_18_12 u_ca_18_12_46(.d_in(u_ca_in_46), .d_out(u_ca_out_46));
compressor_18_12 u_ca_18_12_47(.d_in(u_ca_in_47), .d_out(u_ca_out_47));
compressor_18_12 u_ca_18_12_48(.d_in(u_ca_in_48), .d_out(u_ca_out_48));
compressor_18_12 u_ca_18_12_49(.d_in(u_ca_in_49), .d_out(u_ca_out_49));
compressor_18_12 u_ca_18_12_50(.d_in(u_ca_in_50), .d_out(u_ca_out_50));
compressor_18_12 u_ca_18_12_51(.d_in(u_ca_in_51), .d_out(u_ca_out_51));
compressor_18_12 u_ca_18_12_52(.d_in(u_ca_in_52), .d_out(u_ca_out_52));
compressor_18_12 u_ca_18_12_53(.d_in(u_ca_in_53), .d_out(u_ca_out_53));
compressor_18_12 u_ca_18_12_54(.d_in(u_ca_in_54), .d_out(u_ca_out_54));
compressor_18_12 u_ca_18_12_55(.d_in(u_ca_in_55), .d_out(u_ca_out_55));
compressor_18_12 u_ca_18_12_56(.d_in(u_ca_in_56), .d_out(u_ca_out_56));
compressor_18_12 u_ca_18_12_57(.d_in(u_ca_in_57), .d_out(u_ca_out_57));
compressor_18_12 u_ca_18_12_58(.d_in(u_ca_in_58), .d_out(u_ca_out_58));
compressor_18_12 u_ca_18_12_59(.d_in(u_ca_in_59), .d_out(u_ca_out_59));
compressor_18_12 u_ca_18_12_60(.d_in(u_ca_in_60), .d_out(u_ca_out_60));
compressor_18_12 u_ca_18_12_61(.d_in(u_ca_in_61), .d_out(u_ca_out_61));
compressor_18_12 u_ca_18_12_62(.d_in(u_ca_in_62), .d_out(u_ca_out_62));
compressor_18_12 u_ca_18_12_63(.d_in(u_ca_in_63), .d_out(u_ca_out_63));
compressor_18_12 u_ca_18_12_64(.d_in(u_ca_in_64), .d_out(u_ca_out_64));
compressor_18_12 u_ca_18_12_65(.d_in(u_ca_in_65), .d_out(u_ca_out_65));
compressor_18_12 u_ca_18_12_66(.d_in(u_ca_in_66), .d_out(u_ca_out_66));
compressor_18_12 u_ca_18_12_67(.d_in(u_ca_in_67), .d_out(u_ca_out_67));
compressor_18_12 u_ca_18_12_68(.d_in(u_ca_in_68), .d_out(u_ca_out_68));
compressor_18_12 u_ca_18_12_69(.d_in(u_ca_in_69), .d_out(u_ca_out_69));
compressor_18_12 u_ca_18_12_70(.d_in(u_ca_in_70), .d_out(u_ca_out_70));
compressor_18_12 u_ca_18_12_71(.d_in(u_ca_in_71), .d_out(u_ca_out_71));
compressor_18_12 u_ca_18_12_72(.d_in(u_ca_in_72), .d_out(u_ca_out_72));
compressor_18_12 u_ca_18_12_73(.d_in(u_ca_in_73), .d_out(u_ca_out_73));
compressor_18_12 u_ca_18_12_74(.d_in(u_ca_in_74), .d_out(u_ca_out_74));
compressor_18_12 u_ca_18_12_75(.d_in(u_ca_in_75), .d_out(u_ca_out_75));
compressor_18_12 u_ca_18_12_76(.d_in(u_ca_in_76), .d_out(u_ca_out_76));
compressor_18_12 u_ca_18_12_77(.d_in(u_ca_in_77), .d_out(u_ca_out_77));
compressor_18_12 u_ca_18_12_78(.d_in(u_ca_in_78), .d_out(u_ca_out_78));
compressor_18_12 u_ca_18_12_79(.d_in(u_ca_in_79), .d_out(u_ca_out_79));
compressor_18_12 u_ca_18_12_80(.d_in(u_ca_in_80), .d_out(u_ca_out_80));
compressor_18_12 u_ca_18_12_81(.d_in(u_ca_in_81), .d_out(u_ca_out_81));
compressor_18_12 u_ca_18_12_82(.d_in(u_ca_in_82), .d_out(u_ca_out_82));
compressor_18_12 u_ca_18_12_83(.d_in(u_ca_in_83), .d_out(u_ca_out_83));
compressor_18_12 u_ca_18_12_84(.d_in(u_ca_in_84), .d_out(u_ca_out_84));
compressor_18_12 u_ca_18_12_85(.d_in(u_ca_in_85), .d_out(u_ca_out_85));
compressor_18_12 u_ca_18_12_86(.d_in(u_ca_in_86), .d_out(u_ca_out_86));
compressor_18_12 u_ca_18_12_87(.d_in(u_ca_in_87), .d_out(u_ca_out_87));
compressor_18_12 u_ca_18_12_88(.d_in(u_ca_in_88), .d_out(u_ca_out_88));
compressor_18_12 u_ca_18_12_89(.d_in(u_ca_in_89), .d_out(u_ca_out_89));
compressor_18_12 u_ca_18_12_90(.d_in(u_ca_in_90), .d_out(u_ca_out_90));
compressor_18_12 u_ca_18_12_91(.d_in(u_ca_in_91), .d_out(u_ca_out_91));
compressor_18_12 u_ca_18_12_92(.d_in(u_ca_in_92), .d_out(u_ca_out_92));
compressor_18_12 u_ca_18_12_93(.d_in(u_ca_in_93), .d_out(u_ca_out_93));
compressor_18_12 u_ca_18_12_94(.d_in(u_ca_in_94), .d_out(u_ca_out_94));
compressor_18_12 u_ca_18_12_95(.d_in(u_ca_in_95), .d_out(u_ca_out_95));
compressor_18_12 u_ca_18_12_96(.d_in(u_ca_in_96), .d_out(u_ca_out_96));
compressor_18_12 u_ca_18_12_97(.d_in(u_ca_in_97), .d_out(u_ca_out_97));
compressor_18_12 u_ca_18_12_98(.d_in(u_ca_in_98), .d_out(u_ca_out_98));
compressor_18_12 u_ca_18_12_99(.d_in(u_ca_in_99), .d_out(u_ca_out_99));
compressor_18_12 u_ca_18_12_100(.d_in(u_ca_in_100), .d_out(u_ca_out_100));
compressor_18_12 u_ca_18_12_101(.d_in(u_ca_in_101), .d_out(u_ca_out_101));
compressor_18_12 u_ca_18_12_102(.d_in(u_ca_in_102), .d_out(u_ca_out_102));
compressor_18_12 u_ca_18_12_103(.d_in(u_ca_in_103), .d_out(u_ca_out_103));
compressor_18_12 u_ca_18_12_104(.d_in(u_ca_in_104), .d_out(u_ca_out_104));
compressor_18_12 u_ca_18_12_105(.d_in(u_ca_in_105), .d_out(u_ca_out_105));
compressor_18_12 u_ca_18_12_106(.d_in(u_ca_in_106), .d_out(u_ca_out_106));
compressor_18_12 u_ca_18_12_107(.d_in(u_ca_in_107), .d_out(u_ca_out_107));
compressor_18_12 u_ca_18_12_108(.d_in(u_ca_in_108), .d_out(u_ca_out_108));
compressor_18_12 u_ca_18_12_109(.d_in(u_ca_in_109), .d_out(u_ca_out_109));
compressor_18_12 u_ca_18_12_110(.d_in(u_ca_in_110), .d_out(u_ca_out_110));
compressor_18_12 u_ca_18_12_111(.d_in(u_ca_in_111), .d_out(u_ca_out_111));
compressor_18_12 u_ca_18_12_112(.d_in(u_ca_in_112), .d_out(u_ca_out_112));
compressor_18_12 u_ca_18_12_113(.d_in(u_ca_in_113), .d_out(u_ca_out_113));
compressor_18_12 u_ca_18_12_114(.d_in(u_ca_in_114), .d_out(u_ca_out_114));
compressor_18_12 u_ca_18_12_115(.d_in(u_ca_in_115), .d_out(u_ca_out_115));
compressor_18_12 u_ca_18_12_116(.d_in(u_ca_in_116), .d_out(u_ca_out_116));
compressor_18_12 u_ca_18_12_117(.d_in(u_ca_in_117), .d_out(u_ca_out_117));
compressor_18_12 u_ca_18_12_118(.d_in(u_ca_in_118), .d_out(u_ca_out_118));
compressor_18_12 u_ca_18_12_119(.d_in(u_ca_in_119), .d_out(u_ca_out_119));
compressor_18_12 u_ca_18_12_120(.d_in(u_ca_in_120), .d_out(u_ca_out_120));
compressor_18_12 u_ca_18_12_121(.d_in(u_ca_in_121), .d_out(u_ca_out_121));
compressor_18_12 u_ca_18_12_122(.d_in(u_ca_in_122), .d_out(u_ca_out_122));
compressor_18_12 u_ca_18_12_123(.d_in(u_ca_in_123), .d_out(u_ca_out_123));
compressor_18_12 u_ca_18_12_124(.d_in(u_ca_in_124), .d_out(u_ca_out_124));
compressor_18_12 u_ca_18_12_125(.d_in(u_ca_in_125), .d_out(u_ca_out_125));
compressor_18_12 u_ca_18_12_126(.d_in(u_ca_in_126), .d_out(u_ca_out_126));
compressor_18_12 u_ca_18_12_127(.d_in(u_ca_in_127), .d_out(u_ca_out_127));
compressor_18_12 u_ca_18_12_128(.d_in(u_ca_in_128), .d_out(u_ca_out_128));
compressor_18_12 u_ca_18_12_129(.d_in(u_ca_in_129), .d_out(u_ca_out_129));
compressor_18_12 u_ca_18_12_130(.d_in(u_ca_in_130), .d_out(u_ca_out_130));
compressor_18_12 u_ca_18_12_131(.d_in(u_ca_in_131), .d_out(u_ca_out_131));
compressor_18_12 u_ca_18_12_132(.d_in(u_ca_in_132), .d_out(u_ca_out_132));
compressor_18_12 u_ca_18_12_133(.d_in(u_ca_in_133), .d_out(u_ca_out_133));
compressor_18_12 u_ca_18_12_134(.d_in(u_ca_in_134), .d_out(u_ca_out_134));
compressor_18_12 u_ca_18_12_135(.d_in(u_ca_in_135), .d_out(u_ca_out_135));
compressor_18_12 u_ca_18_12_136(.d_in(u_ca_in_136), .d_out(u_ca_out_136));
compressor_18_12 u_ca_18_12_137(.d_in(u_ca_in_137), .d_out(u_ca_out_137));
compressor_18_12 u_ca_18_12_138(.d_in(u_ca_in_138), .d_out(u_ca_out_138));
compressor_18_12 u_ca_18_12_139(.d_in(u_ca_in_139), .d_out(u_ca_out_139));
compressor_18_12 u_ca_18_12_140(.d_in(u_ca_in_140), .d_out(u_ca_out_140));
compressor_18_12 u_ca_18_12_141(.d_in(u_ca_in_141), .d_out(u_ca_out_141));
compressor_18_12 u_ca_18_12_142(.d_in(u_ca_in_142), .d_out(u_ca_out_142));
compressor_18_12 u_ca_18_12_143(.d_in(u_ca_in_143), .d_out(u_ca_out_143));
compressor_18_12 u_ca_18_12_144(.d_in(u_ca_in_144), .d_out(u_ca_out_144));
compressor_18_12 u_ca_18_12_145(.d_in(u_ca_in_145), .d_out(u_ca_out_145));
compressor_18_12 u_ca_18_12_146(.d_in(u_ca_in_146), .d_out(u_ca_out_146));
compressor_18_12 u_ca_18_12_147(.d_in(u_ca_in_147), .d_out(u_ca_out_147));
compressor_18_12 u_ca_18_12_148(.d_in(u_ca_in_148), .d_out(u_ca_out_148));
compressor_18_12 u_ca_18_12_149(.d_in(u_ca_in_149), .d_out(u_ca_out_149));
compressor_18_12 u_ca_18_12_150(.d_in(u_ca_in_150), .d_out(u_ca_out_150));
compressor_18_12 u_ca_18_12_151(.d_in(u_ca_in_151), .d_out(u_ca_out_151));
compressor_18_12 u_ca_18_12_152(.d_in(u_ca_in_152), .d_out(u_ca_out_152));
compressor_18_12 u_ca_18_12_153(.d_in(u_ca_in_153), .d_out(u_ca_out_153));
compressor_18_12 u_ca_18_12_154(.d_in(u_ca_in_154), .d_out(u_ca_out_154));
compressor_18_12 u_ca_18_12_155(.d_in(u_ca_in_155), .d_out(u_ca_out_155));
compressor_18_12 u_ca_18_12_156(.d_in(u_ca_in_156), .d_out(u_ca_out_156));
compressor_18_12 u_ca_18_12_157(.d_in(u_ca_in_157), .d_out(u_ca_out_157));
compressor_18_12 u_ca_18_12_158(.d_in(u_ca_in_158), .d_out(u_ca_out_158));
compressor_18_12 u_ca_18_12_159(.d_in(u_ca_in_159), .d_out(u_ca_out_159));
compressor_18_12 u_ca_18_12_160(.d_in(u_ca_in_160), .d_out(u_ca_out_160));
compressor_18_12 u_ca_18_12_161(.d_in(u_ca_in_161), .d_out(u_ca_out_161));
compressor_18_12 u_ca_18_12_162(.d_in(u_ca_in_162), .d_out(u_ca_out_162));
compressor_18_12 u_ca_18_12_163(.d_in(u_ca_in_163), .d_out(u_ca_out_163));
compressor_18_12 u_ca_18_12_164(.d_in(u_ca_in_164), .d_out(u_ca_out_164));
compressor_18_12 u_ca_18_12_165(.d_in(u_ca_in_165), .d_out(u_ca_out_165));
compressor_18_12 u_ca_18_12_166(.d_in(u_ca_in_166), .d_out(u_ca_out_166));
compressor_18_12 u_ca_18_12_167(.d_in(u_ca_in_167), .d_out(u_ca_out_167));
compressor_18_12 u_ca_18_12_168(.d_in(u_ca_in_168), .d_out(u_ca_out_168));
compressor_18_12 u_ca_18_12_169(.d_in(u_ca_in_169), .d_out(u_ca_out_169));
compressor_18_12 u_ca_18_12_170(.d_in(u_ca_in_170), .d_out(u_ca_out_170));
compressor_18_12 u_ca_18_12_171(.d_in(u_ca_in_171), .d_out(u_ca_out_171));
compressor_18_12 u_ca_18_12_172(.d_in(u_ca_in_172), .d_out(u_ca_out_172));
compressor_18_12 u_ca_18_12_173(.d_in(u_ca_in_173), .d_out(u_ca_out_173));
compressor_18_12 u_ca_18_12_174(.d_in(u_ca_in_174), .d_out(u_ca_out_174));
compressor_18_12 u_ca_18_12_175(.d_in(u_ca_in_175), .d_out(u_ca_out_175));
compressor_18_12 u_ca_18_12_176(.d_in(u_ca_in_176), .d_out(u_ca_out_176));
compressor_18_12 u_ca_18_12_177(.d_in(u_ca_in_177), .d_out(u_ca_out_177));
compressor_18_12 u_ca_18_12_178(.d_in(u_ca_in_178), .d_out(u_ca_out_178));
compressor_18_12 u_ca_18_12_179(.d_in(u_ca_in_179), .d_out(u_ca_out_179));
compressor_18_12 u_ca_18_12_180(.d_in(u_ca_in_180), .d_out(u_ca_out_180));
compressor_18_12 u_ca_18_12_181(.d_in(u_ca_in_181), .d_out(u_ca_out_181));
compressor_18_12 u_ca_18_12_182(.d_in(u_ca_in_182), .d_out(u_ca_out_182));
compressor_18_12 u_ca_18_12_183(.d_in(u_ca_in_183), .d_out(u_ca_out_183));
compressor_18_12 u_ca_18_12_184(.d_in(u_ca_in_184), .d_out(u_ca_out_184));
compressor_18_12 u_ca_18_12_185(.d_in(u_ca_in_185), .d_out(u_ca_out_185));
compressor_18_12 u_ca_18_12_186(.d_in(u_ca_in_186), .d_out(u_ca_out_186));
compressor_18_12 u_ca_18_12_187(.d_in(u_ca_in_187), .d_out(u_ca_out_187));
compressor_18_12 u_ca_18_12_188(.d_in(u_ca_in_188), .d_out(u_ca_out_188));
compressor_18_12 u_ca_18_12_189(.d_in(u_ca_in_189), .d_out(u_ca_out_189));
compressor_18_12 u_ca_18_12_190(.d_in(u_ca_in_190), .d_out(u_ca_out_190));
compressor_18_12 u_ca_18_12_191(.d_in(u_ca_in_191), .d_out(u_ca_out_191));
compressor_18_12 u_ca_18_12_192(.d_in(u_ca_in_192), .d_out(u_ca_out_192));
compressor_18_12 u_ca_18_12_193(.d_in(u_ca_in_193), .d_out(u_ca_out_193));
compressor_18_12 u_ca_18_12_194(.d_in(u_ca_in_194), .d_out(u_ca_out_194));
compressor_18_12 u_ca_18_12_195(.d_in(u_ca_in_195), .d_out(u_ca_out_195));
compressor_18_12 u_ca_18_12_196(.d_in(u_ca_in_196), .d_out(u_ca_out_196));
compressor_18_12 u_ca_18_12_197(.d_in(u_ca_in_197), .d_out(u_ca_out_197));
compressor_18_12 u_ca_18_12_198(.d_in(u_ca_in_198), .d_out(u_ca_out_198));
compressor_18_12 u_ca_18_12_199(.d_in(u_ca_in_199), .d_out(u_ca_out_199));
compressor_18_12 u_ca_18_12_200(.d_in(u_ca_in_200), .d_out(u_ca_out_200));
compressor_18_12 u_ca_18_12_201(.d_in(u_ca_in_201), .d_out(u_ca_out_201));
compressor_18_12 u_ca_18_12_202(.d_in(u_ca_in_202), .d_out(u_ca_out_202));
compressor_18_12 u_ca_18_12_203(.d_in(u_ca_in_203), .d_out(u_ca_out_203));
compressor_18_12 u_ca_18_12_204(.d_in(u_ca_in_204), .d_out(u_ca_out_204));
compressor_18_12 u_ca_18_12_205(.d_in(u_ca_in_205), .d_out(u_ca_out_205));
compressor_18_12 u_ca_18_12_206(.d_in(u_ca_in_206), .d_out(u_ca_out_206));
compressor_18_12 u_ca_18_12_207(.d_in(u_ca_in_207), .d_out(u_ca_out_207));
compressor_18_12 u_ca_18_12_208(.d_in(u_ca_in_208), .d_out(u_ca_out_208));
compressor_18_12 u_ca_18_12_209(.d_in(u_ca_in_209), .d_out(u_ca_out_209));
compressor_18_12 u_ca_18_12_210(.d_in(u_ca_in_210), .d_out(u_ca_out_210));
compressor_18_12 u_ca_18_12_211(.d_in(u_ca_in_211), .d_out(u_ca_out_211));
compressor_18_12 u_ca_18_12_212(.d_in(u_ca_in_212), .d_out(u_ca_out_212));
compressor_18_12 u_ca_18_12_213(.d_in(u_ca_in_213), .d_out(u_ca_out_213));
compressor_18_12 u_ca_18_12_214(.d_in(u_ca_in_214), .d_out(u_ca_out_214));
compressor_18_12 u_ca_18_12_215(.d_in(u_ca_in_215), .d_out(u_ca_out_215));
compressor_18_12 u_ca_18_12_216(.d_in(u_ca_in_216), .d_out(u_ca_out_216));
compressor_18_12 u_ca_18_12_217(.d_in(u_ca_in_217), .d_out(u_ca_out_217));
compressor_18_12 u_ca_18_12_218(.d_in(u_ca_in_218), .d_out(u_ca_out_218));
compressor_18_12 u_ca_18_12_219(.d_in(u_ca_in_219), .d_out(u_ca_out_219));
compressor_18_12 u_ca_18_12_220(.d_in(u_ca_in_220), .d_out(u_ca_out_220));
compressor_18_12 u_ca_18_12_221(.d_in(u_ca_in_221), .d_out(u_ca_out_221));
compressor_18_12 u_ca_18_12_222(.d_in(u_ca_in_222), .d_out(u_ca_out_222));
compressor_18_12 u_ca_18_12_223(.d_in(u_ca_in_223), .d_out(u_ca_out_223));
compressor_18_12 u_ca_18_12_224(.d_in(u_ca_in_224), .d_out(u_ca_out_224));
compressor_18_12 u_ca_18_12_225(.d_in(u_ca_in_225), .d_out(u_ca_out_225));
compressor_18_12 u_ca_18_12_226(.d_in(u_ca_in_226), .d_out(u_ca_out_226));
compressor_18_12 u_ca_18_12_227(.d_in(u_ca_in_227), .d_out(u_ca_out_227));
compressor_18_12 u_ca_18_12_228(.d_in(u_ca_in_228), .d_out(u_ca_out_228));
compressor_18_12 u_ca_18_12_229(.d_in(u_ca_in_229), .d_out(u_ca_out_229));
compressor_18_12 u_ca_18_12_230(.d_in(u_ca_in_230), .d_out(u_ca_out_230));
compressor_18_12 u_ca_18_12_231(.d_in(u_ca_in_231), .d_out(u_ca_out_231));
compressor_18_12 u_ca_18_12_232(.d_in(u_ca_in_232), .d_out(u_ca_out_232));
compressor_18_12 u_ca_18_12_233(.d_in(u_ca_in_233), .d_out(u_ca_out_233));
compressor_18_12 u_ca_18_12_234(.d_in(u_ca_in_234), .d_out(u_ca_out_234));
compressor_18_12 u_ca_18_12_235(.d_in(u_ca_in_235), .d_out(u_ca_out_235));
compressor_18_12 u_ca_18_12_236(.d_in(u_ca_in_236), .d_out(u_ca_out_236));
compressor_18_12 u_ca_18_12_237(.d_in(u_ca_in_237), .d_out(u_ca_out_237));
compressor_18_12 u_ca_18_12_238(.d_in(u_ca_in_238), .d_out(u_ca_out_238));
compressor_18_12 u_ca_18_12_239(.d_in(u_ca_in_239), .d_out(u_ca_out_239));
compressor_18_12 u_ca_18_12_240(.d_in(u_ca_in_240), .d_out(u_ca_out_240));
compressor_18_12 u_ca_18_12_241(.d_in(u_ca_in_241), .d_out(u_ca_out_241));
compressor_18_12 u_ca_18_12_242(.d_in(u_ca_in_242), .d_out(u_ca_out_242));
compressor_18_12 u_ca_18_12_243(.d_in(u_ca_in_243), .d_out(u_ca_out_243));
compressor_18_12 u_ca_18_12_244(.d_in(u_ca_in_244), .d_out(u_ca_out_244));
compressor_18_12 u_ca_18_12_245(.d_in(u_ca_in_245), .d_out(u_ca_out_245));
compressor_18_12 u_ca_18_12_246(.d_in(u_ca_in_246), .d_out(u_ca_out_246));
compressor_18_12 u_ca_18_12_247(.d_in(u_ca_in_247), .d_out(u_ca_out_247));
compressor_18_12 u_ca_18_12_248(.d_in(u_ca_in_248), .d_out(u_ca_out_248));
compressor_18_12 u_ca_18_12_249(.d_in(u_ca_in_249), .d_out(u_ca_out_249));
compressor_18_12 u_ca_18_12_250(.d_in(u_ca_in_250), .d_out(u_ca_out_250));
compressor_18_12 u_ca_18_12_251(.d_in(u_ca_in_251), .d_out(u_ca_out_251));
compressor_18_12 u_ca_18_12_252(.d_in(u_ca_in_252), .d_out(u_ca_out_252));
compressor_18_12 u_ca_18_12_253(.d_in(u_ca_in_253), .d_out(u_ca_out_253));
compressor_18_12 u_ca_18_12_254(.d_in(u_ca_in_254), .d_out(u_ca_out_254));
compressor_18_12 u_ca_18_12_255(.d_in(u_ca_in_255), .d_out(u_ca_out_255));
compressor_18_12 u_ca_18_12_256(.d_in(u_ca_in_256), .d_out(u_ca_out_256));
compressor_18_12 u_ca_18_12_257(.d_in(u_ca_in_257), .d_out(u_ca_out_257));
compressor_18_12 u_ca_18_12_258(.d_in(u_ca_in_258), .d_out(u_ca_out_258));
compressor_18_12 u_ca_18_12_259(.d_in(u_ca_in_259), .d_out(u_ca_out_259));
compressor_18_12 u_ca_18_12_260(.d_in(u_ca_in_260), .d_out(u_ca_out_260));
compressor_18_12 u_ca_18_12_261(.d_in(u_ca_in_261), .d_out(u_ca_out_261));
compressor_18_12 u_ca_18_12_262(.d_in(u_ca_in_262), .d_out(u_ca_out_262));
compressor_18_12 u_ca_18_12_263(.d_in(u_ca_in_263), .d_out(u_ca_out_263));
compressor_18_12 u_ca_18_12_264(.d_in(u_ca_in_264), .d_out(u_ca_out_264));
compressor_18_12 u_ca_18_12_265(.d_in(u_ca_in_265), .d_out(u_ca_out_265));
compressor_18_12 u_ca_18_12_266(.d_in(u_ca_in_266), .d_out(u_ca_out_266));
compressor_18_12 u_ca_18_12_267(.d_in(u_ca_in_267), .d_out(u_ca_out_267));
compressor_18_12 u_ca_18_12_268(.d_in(u_ca_in_268), .d_out(u_ca_out_268));
compressor_18_12 u_ca_18_12_269(.d_in(u_ca_in_269), .d_out(u_ca_out_269));
compressor_18_12 u_ca_18_12_270(.d_in(u_ca_in_270), .d_out(u_ca_out_270));
compressor_18_12 u_ca_18_12_271(.d_in(u_ca_in_271), .d_out(u_ca_out_271));
compressor_18_12 u_ca_18_12_272(.d_in(u_ca_in_272), .d_out(u_ca_out_272));
compressor_18_12 u_ca_18_12_273(.d_in(u_ca_in_273), .d_out(u_ca_out_273));
compressor_18_12 u_ca_18_12_274(.d_in(u_ca_in_274), .d_out(u_ca_out_274));
compressor_18_12 u_ca_18_12_275(.d_in(u_ca_in_275), .d_out(u_ca_out_275));
compressor_18_12 u_ca_18_12_276(.d_in(u_ca_in_276), .d_out(u_ca_out_276));
compressor_18_12 u_ca_18_12_277(.d_in(u_ca_in_277), .d_out(u_ca_out_277));
compressor_18_12 u_ca_18_12_278(.d_in(u_ca_in_278), .d_out(u_ca_out_278));
compressor_18_12 u_ca_18_12_279(.d_in(u_ca_in_279), .d_out(u_ca_out_279));
compressor_18_12 u_ca_18_12_280(.d_in(u_ca_in_280), .d_out(u_ca_out_280));
compressor_18_12 u_ca_18_12_281(.d_in(u_ca_in_281), .d_out(u_ca_out_281));
compressor_18_12 u_ca_18_12_282(.d_in(u_ca_in_282), .d_out(u_ca_out_282));
compressor_18_12 u_ca_18_12_283(.d_in(u_ca_in_283), .d_out(u_ca_out_283));
compressor_18_12 u_ca_18_12_284(.d_in(u_ca_in_284), .d_out(u_ca_out_284));
compressor_18_12 u_ca_18_12_285(.d_in(u_ca_in_285), .d_out(u_ca_out_285));
compressor_18_12 u_ca_18_12_286(.d_in(u_ca_in_286), .d_out(u_ca_out_286));
compressor_18_12 u_ca_18_12_287(.d_in(u_ca_in_287), .d_out(u_ca_out_287));
compressor_18_12 u_ca_18_12_288(.d_in(u_ca_in_288), .d_out(u_ca_out_288));
compressor_18_12 u_ca_18_12_289(.d_in(u_ca_in_289), .d_out(u_ca_out_289));
compressor_18_12 u_ca_18_12_290(.d_in(u_ca_in_290), .d_out(u_ca_out_290));
compressor_18_12 u_ca_18_12_291(.d_in(u_ca_in_291), .d_out(u_ca_out_291));
compressor_18_12 u_ca_18_12_292(.d_in(u_ca_in_292), .d_out(u_ca_out_292));
compressor_18_12 u_ca_18_12_293(.d_in(u_ca_in_293), .d_out(u_ca_out_293));
compressor_18_12 u_ca_18_12_294(.d_in(u_ca_in_294), .d_out(u_ca_out_294));
compressor_18_12 u_ca_18_12_295(.d_in(u_ca_in_295), .d_out(u_ca_out_295));
compressor_18_12 u_ca_18_12_296(.d_in(u_ca_in_296), .d_out(u_ca_out_296));
compressor_18_12 u_ca_18_12_297(.d_in(u_ca_in_297), .d_out(u_ca_out_297));
compressor_18_12 u_ca_18_12_298(.d_in(u_ca_in_298), .d_out(u_ca_out_298));
compressor_18_12 u_ca_18_12_299(.d_in(u_ca_in_299), .d_out(u_ca_out_299));
compressor_18_12 u_ca_18_12_300(.d_in(u_ca_in_300), .d_out(u_ca_out_300));
compressor_18_12 u_ca_18_12_301(.d_in(u_ca_in_301), .d_out(u_ca_out_301));
compressor_18_12 u_ca_18_12_302(.d_in(u_ca_in_302), .d_out(u_ca_out_302));
compressor_18_12 u_ca_18_12_303(.d_in(u_ca_in_303), .d_out(u_ca_out_303));
compressor_18_12 u_ca_18_12_304(.d_in(u_ca_in_304), .d_out(u_ca_out_304));
compressor_18_12 u_ca_18_12_305(.d_in(u_ca_in_305), .d_out(u_ca_out_305));
compressor_18_12 u_ca_18_12_306(.d_in(u_ca_in_306), .d_out(u_ca_out_306));
compressor_18_12 u_ca_18_12_307(.d_in(u_ca_in_307), .d_out(u_ca_out_307));
compressor_18_12 u_ca_18_12_308(.d_in(u_ca_in_308), .d_out(u_ca_out_308));
compressor_18_12 u_ca_18_12_309(.d_in(u_ca_in_309), .d_out(u_ca_out_309));
compressor_18_12 u_ca_18_12_310(.d_in(u_ca_in_310), .d_out(u_ca_out_310));
compressor_18_12 u_ca_18_12_311(.d_in(u_ca_in_311), .d_out(u_ca_out_311));
compressor_18_12 u_ca_18_12_312(.d_in(u_ca_in_312), .d_out(u_ca_out_312));
compressor_18_12 u_ca_18_12_313(.d_in(u_ca_in_313), .d_out(u_ca_out_313));
compressor_18_12 u_ca_18_12_314(.d_in(u_ca_in_314), .d_out(u_ca_out_314));
compressor_18_12 u_ca_18_12_315(.d_in(u_ca_in_315), .d_out(u_ca_out_315));
compressor_18_12 u_ca_18_12_316(.d_in(u_ca_in_316), .d_out(u_ca_out_316));
compressor_18_12 u_ca_18_12_317(.d_in(u_ca_in_317), .d_out(u_ca_out_317));
compressor_18_12 u_ca_18_12_318(.d_in(u_ca_in_318), .d_out(u_ca_out_318));
compressor_18_12 u_ca_18_12_319(.d_in(u_ca_in_319), .d_out(u_ca_out_319));
compressor_18_12 u_ca_18_12_320(.d_in(u_ca_in_320), .d_out(u_ca_out_320));
compressor_18_12 u_ca_18_12_321(.d_in(u_ca_in_321), .d_out(u_ca_out_321));
compressor_18_12 u_ca_18_12_322(.d_in(u_ca_in_322), .d_out(u_ca_out_322));
compressor_18_12 u_ca_18_12_323(.d_in(u_ca_in_323), .d_out(u_ca_out_323));
compressor_18_12 u_ca_18_12_324(.d_in(u_ca_in_324), .d_out(u_ca_out_324));
compressor_18_12 u_ca_18_12_325(.d_in(u_ca_in_325), .d_out(u_ca_out_325));
compressor_18_12 u_ca_18_12_326(.d_in(u_ca_in_326), .d_out(u_ca_out_326));
compressor_18_12 u_ca_18_12_327(.d_in(u_ca_in_327), .d_out(u_ca_out_327));
compressor_18_12 u_ca_18_12_328(.d_in(u_ca_in_328), .d_out(u_ca_out_328));
compressor_18_12 u_ca_18_12_329(.d_in(u_ca_in_329), .d_out(u_ca_out_329));
compressor_18_12 u_ca_18_12_330(.d_in(u_ca_in_330), .d_out(u_ca_out_330));
compressor_18_12 u_ca_18_12_331(.d_in(u_ca_in_331), .d_out(u_ca_out_331));
compressor_18_12 u_ca_18_12_332(.d_in(u_ca_in_332), .d_out(u_ca_out_332));
compressor_18_12 u_ca_18_12_333(.d_in(u_ca_in_333), .d_out(u_ca_out_333));
compressor_18_12 u_ca_18_12_334(.d_in(u_ca_in_334), .d_out(u_ca_out_334));
compressor_18_12 u_ca_18_12_335(.d_in(u_ca_in_335), .d_out(u_ca_out_335));
compressor_18_12 u_ca_18_12_336(.d_in(u_ca_in_336), .d_out(u_ca_out_336));
compressor_18_12 u_ca_18_12_337(.d_in(u_ca_in_337), .d_out(u_ca_out_337));
compressor_18_12 u_ca_18_12_338(.d_in(u_ca_in_338), .d_out(u_ca_out_338));
compressor_18_12 u_ca_18_12_339(.d_in(u_ca_in_339), .d_out(u_ca_out_339));
compressor_18_12 u_ca_18_12_340(.d_in(u_ca_in_340), .d_out(u_ca_out_340));
compressor_18_12 u_ca_18_12_341(.d_in(u_ca_in_341), .d_out(u_ca_out_341));
compressor_18_12 u_ca_18_12_342(.d_in(u_ca_in_342), .d_out(u_ca_out_342));
compressor_18_12 u_ca_18_12_343(.d_in(u_ca_in_343), .d_out(u_ca_out_343));
compressor_18_12 u_ca_18_12_344(.d_in(u_ca_in_344), .d_out(u_ca_out_344));
compressor_18_12 u_ca_18_12_345(.d_in(u_ca_in_345), .d_out(u_ca_out_345));
compressor_18_12 u_ca_18_12_346(.d_in(u_ca_in_346), .d_out(u_ca_out_346));
compressor_18_12 u_ca_18_12_347(.d_in(u_ca_in_347), .d_out(u_ca_out_347));
compressor_18_12 u_ca_18_12_348(.d_in(u_ca_in_348), .d_out(u_ca_out_348));
compressor_18_12 u_ca_18_12_349(.d_in(u_ca_in_349), .d_out(u_ca_out_349));
compressor_18_12 u_ca_18_12_350(.d_in(u_ca_in_350), .d_out(u_ca_out_350));
compressor_18_12 u_ca_18_12_351(.d_in(u_ca_in_351), .d_out(u_ca_out_351));
compressor_18_12 u_ca_18_12_352(.d_in(u_ca_in_352), .d_out(u_ca_out_352));
compressor_18_12 u_ca_18_12_353(.d_in(u_ca_in_353), .d_out(u_ca_out_353));
compressor_18_12 u_ca_18_12_354(.d_in(u_ca_in_354), .d_out(u_ca_out_354));
compressor_18_12 u_ca_18_12_355(.d_in(u_ca_in_355), .d_out(u_ca_out_355));
compressor_18_12 u_ca_18_12_356(.d_in(u_ca_in_356), .d_out(u_ca_out_356));
compressor_18_12 u_ca_18_12_357(.d_in(u_ca_in_357), .d_out(u_ca_out_357));
compressor_18_12 u_ca_18_12_358(.d_in(u_ca_in_358), .d_out(u_ca_out_358));
compressor_18_12 u_ca_18_12_359(.d_in(u_ca_in_359), .d_out(u_ca_out_359));
compressor_18_12 u_ca_18_12_360(.d_in(u_ca_in_360), .d_out(u_ca_out_360));
compressor_18_12 u_ca_18_12_361(.d_in(u_ca_in_361), .d_out(u_ca_out_361));
compressor_18_12 u_ca_18_12_362(.d_in(u_ca_in_362), .d_out(u_ca_out_362));
compressor_18_12 u_ca_18_12_363(.d_in(u_ca_in_363), .d_out(u_ca_out_363));
compressor_18_12 u_ca_18_12_364(.d_in(u_ca_in_364), .d_out(u_ca_out_364));
compressor_18_12 u_ca_18_12_365(.d_in(u_ca_in_365), .d_out(u_ca_out_365));
compressor_18_12 u_ca_18_12_366(.d_in(u_ca_in_366), .d_out(u_ca_out_366));
compressor_18_12 u_ca_18_12_367(.d_in(u_ca_in_367), .d_out(u_ca_out_367));
compressor_18_12 u_ca_18_12_368(.d_in(u_ca_in_368), .d_out(u_ca_out_368));
compressor_18_12 u_ca_18_12_369(.d_in(u_ca_in_369), .d_out(u_ca_out_369));
compressor_18_12 u_ca_18_12_370(.d_in(u_ca_in_370), .d_out(u_ca_out_370));
compressor_18_12 u_ca_18_12_371(.d_in(u_ca_in_371), .d_out(u_ca_out_371));
compressor_18_12 u_ca_18_12_372(.d_in(u_ca_in_372), .d_out(u_ca_out_372));
compressor_18_12 u_ca_18_12_373(.d_in(u_ca_in_373), .d_out(u_ca_out_373));
compressor_18_12 u_ca_18_12_374(.d_in(u_ca_in_374), .d_out(u_ca_out_374));
compressor_18_12 u_ca_18_12_375(.d_in(u_ca_in_375), .d_out(u_ca_out_375));
compressor_18_12 u_ca_18_12_376(.d_in(u_ca_in_376), .d_out(u_ca_out_376));
compressor_18_12 u_ca_18_12_377(.d_in(u_ca_in_377), .d_out(u_ca_out_377));
compressor_18_12 u_ca_18_12_378(.d_in(u_ca_in_378), .d_out(u_ca_out_378));
compressor_18_12 u_ca_18_12_379(.d_in(u_ca_in_379), .d_out(u_ca_out_379));
compressor_18_12 u_ca_18_12_380(.d_in(u_ca_in_380), .d_out(u_ca_out_380));
compressor_18_12 u_ca_18_12_381(.d_in(u_ca_in_381), .d_out(u_ca_out_381));
compressor_18_12 u_ca_18_12_382(.d_in(u_ca_in_382), .d_out(u_ca_out_382));
compressor_18_12 u_ca_18_12_383(.d_in(u_ca_in_383), .d_out(u_ca_out_383));
compressor_18_12 u_ca_18_12_384(.d_in(u_ca_in_384), .d_out(u_ca_out_384));
compressor_18_12 u_ca_18_12_385(.d_in(u_ca_in_385), .d_out(u_ca_out_385));
compressor_18_12 u_ca_18_12_386(.d_in(u_ca_in_386), .d_out(u_ca_out_386));
compressor_18_12 u_ca_18_12_387(.d_in(u_ca_in_387), .d_out(u_ca_out_387));
compressor_18_12 u_ca_18_12_388(.d_in(u_ca_in_388), .d_out(u_ca_out_388));
compressor_18_12 u_ca_18_12_389(.d_in(u_ca_in_389), .d_out(u_ca_out_389));
compressor_18_12 u_ca_18_12_390(.d_in(u_ca_in_390), .d_out(u_ca_out_390));
compressor_18_12 u_ca_18_12_391(.d_in(u_ca_in_391), .d_out(u_ca_out_391));
compressor_18_12 u_ca_18_12_392(.d_in(u_ca_in_392), .d_out(u_ca_out_392));
compressor_18_12 u_ca_18_12_393(.d_in(u_ca_in_393), .d_out(u_ca_out_393));
compressor_18_12 u_ca_18_12_394(.d_in(u_ca_in_394), .d_out(u_ca_out_394));
compressor_18_12 u_ca_18_12_395(.d_in(u_ca_in_395), .d_out(u_ca_out_395));
compressor_18_12 u_ca_18_12_396(.d_in(u_ca_in_396), .d_out(u_ca_out_396));
compressor_18_12 u_ca_18_12_397(.d_in(u_ca_in_397), .d_out(u_ca_out_397));
compressor_18_12 u_ca_18_12_398(.d_in(u_ca_in_398), .d_out(u_ca_out_398));
compressor_18_12 u_ca_18_12_399(.d_in(u_ca_in_399), .d_out(u_ca_out_399));
compressor_18_12 u_ca_18_12_400(.d_in(u_ca_in_400), .d_out(u_ca_out_400));
compressor_18_12 u_ca_18_12_401(.d_in(u_ca_in_401), .d_out(u_ca_out_401));
compressor_18_12 u_ca_18_12_402(.d_in(u_ca_in_402), .d_out(u_ca_out_402));
compressor_18_12 u_ca_18_12_403(.d_in(u_ca_in_403), .d_out(u_ca_out_403));
compressor_18_12 u_ca_18_12_404(.d_in(u_ca_in_404), .d_out(u_ca_out_404));
compressor_18_12 u_ca_18_12_405(.d_in(u_ca_in_405), .d_out(u_ca_out_405));
compressor_18_12 u_ca_18_12_406(.d_in(u_ca_in_406), .d_out(u_ca_out_406));
compressor_18_12 u_ca_18_12_407(.d_in(u_ca_in_407), .d_out(u_ca_out_407));
compressor_18_12 u_ca_18_12_408(.d_in(u_ca_in_408), .d_out(u_ca_out_408));
compressor_18_12 u_ca_18_12_409(.d_in(u_ca_in_409), .d_out(u_ca_out_409));
compressor_18_12 u_ca_18_12_410(.d_in(u_ca_in_410), .d_out(u_ca_out_410));
compressor_18_12 u_ca_18_12_411(.d_in(u_ca_in_411), .d_out(u_ca_out_411));
compressor_18_12 u_ca_18_12_412(.d_in(u_ca_in_412), .d_out(u_ca_out_412));
compressor_18_12 u_ca_18_12_413(.d_in(u_ca_in_413), .d_out(u_ca_out_413));
compressor_18_12 u_ca_18_12_414(.d_in(u_ca_in_414), .d_out(u_ca_out_414));
compressor_18_12 u_ca_18_12_415(.d_in(u_ca_in_415), .d_out(u_ca_out_415));
compressor_18_12 u_ca_18_12_416(.d_in(u_ca_in_416), .d_out(u_ca_out_416));
compressor_18_12 u_ca_18_12_417(.d_in(u_ca_in_417), .d_out(u_ca_out_417));
compressor_18_12 u_ca_18_12_418(.d_in(u_ca_in_418), .d_out(u_ca_out_418));
compressor_18_12 u_ca_18_12_419(.d_in(u_ca_in_419), .d_out(u_ca_out_419));
compressor_18_12 u_ca_18_12_420(.d_in(u_ca_in_420), .d_out(u_ca_out_420));
compressor_18_12 u_ca_18_12_421(.d_in(u_ca_in_421), .d_out(u_ca_out_421));
compressor_18_12 u_ca_18_12_422(.d_in(u_ca_in_422), .d_out(u_ca_out_422));
compressor_18_12 u_ca_18_12_423(.d_in(u_ca_in_423), .d_out(u_ca_out_423));
compressor_18_12 u_ca_18_12_424(.d_in(u_ca_in_424), .d_out(u_ca_out_424));
compressor_18_12 u_ca_18_12_425(.d_in(u_ca_in_425), .d_out(u_ca_out_425));
compressor_18_12 u_ca_18_12_426(.d_in(u_ca_in_426), .d_out(u_ca_out_426));
compressor_18_12 u_ca_18_12_427(.d_in(u_ca_in_427), .d_out(u_ca_out_427));
compressor_18_12 u_ca_18_12_428(.d_in(u_ca_in_428), .d_out(u_ca_out_428));
compressor_18_12 u_ca_18_12_429(.d_in(u_ca_in_429), .d_out(u_ca_out_429));
compressor_18_12 u_ca_18_12_430(.d_in(u_ca_in_430), .d_out(u_ca_out_430));
compressor_18_12 u_ca_18_12_431(.d_in(u_ca_in_431), .d_out(u_ca_out_431));
compressor_18_12 u_ca_18_12_432(.d_in(u_ca_in_432), .d_out(u_ca_out_432));
compressor_18_12 u_ca_18_12_433(.d_in(u_ca_in_433), .d_out(u_ca_out_433));
compressor_18_12 u_ca_18_12_434(.d_in(u_ca_in_434), .d_out(u_ca_out_434));
compressor_18_12 u_ca_18_12_435(.d_in(u_ca_in_435), .d_out(u_ca_out_435));
compressor_18_12 u_ca_18_12_436(.d_in(u_ca_in_436), .d_out(u_ca_out_436));
compressor_18_12 u_ca_18_12_437(.d_in(u_ca_in_437), .d_out(u_ca_out_437));
compressor_18_12 u_ca_18_12_438(.d_in(u_ca_in_438), .d_out(u_ca_out_438));
compressor_18_12 u_ca_18_12_439(.d_in(u_ca_in_439), .d_out(u_ca_out_439));
compressor_18_12 u_ca_18_12_440(.d_in(u_ca_in_440), .d_out(u_ca_out_440));
compressor_18_12 u_ca_18_12_441(.d_in(u_ca_in_441), .d_out(u_ca_out_441));
compressor_18_12 u_ca_18_12_442(.d_in(u_ca_in_442), .d_out(u_ca_out_442));
compressor_18_12 u_ca_18_12_443(.d_in(u_ca_in_443), .d_out(u_ca_out_443));
compressor_18_12 u_ca_18_12_444(.d_in(u_ca_in_444), .d_out(u_ca_out_444));
compressor_18_12 u_ca_18_12_445(.d_in(u_ca_in_445), .d_out(u_ca_out_445));
compressor_18_12 u_ca_18_12_446(.d_in(u_ca_in_446), .d_out(u_ca_out_446));
compressor_18_12 u_ca_18_12_447(.d_in(u_ca_in_447), .d_out(u_ca_out_447));
compressor_18_12 u_ca_18_12_448(.d_in(u_ca_in_448), .d_out(u_ca_out_448));
compressor_18_12 u_ca_18_12_449(.d_in(u_ca_in_449), .d_out(u_ca_out_449));
compressor_18_12 u_ca_18_12_450(.d_in(u_ca_in_450), .d_out(u_ca_out_450));
compressor_18_12 u_ca_18_12_451(.d_in(u_ca_in_451), .d_out(u_ca_out_451));
compressor_18_12 u_ca_18_12_452(.d_in(u_ca_in_452), .d_out(u_ca_out_452));
compressor_18_12 u_ca_18_12_453(.d_in(u_ca_in_453), .d_out(u_ca_out_453));
compressor_18_12 u_ca_18_12_454(.d_in(u_ca_in_454), .d_out(u_ca_out_454));
compressor_18_12 u_ca_18_12_455(.d_in(u_ca_in_455), .d_out(u_ca_out_455));
compressor_18_12 u_ca_18_12_456(.d_in(u_ca_in_456), .d_out(u_ca_out_456));
compressor_18_12 u_ca_18_12_457(.d_in(u_ca_in_457), .d_out(u_ca_out_457));
compressor_18_12 u_ca_18_12_458(.d_in(u_ca_in_458), .d_out(u_ca_out_458));
compressor_18_12 u_ca_18_12_459(.d_in(u_ca_in_459), .d_out(u_ca_out_459));
compressor_18_12 u_ca_18_12_460(.d_in(u_ca_in_460), .d_out(u_ca_out_460));
compressor_18_12 u_ca_18_12_461(.d_in(u_ca_in_461), .d_out(u_ca_out_461));
compressor_18_12 u_ca_18_12_462(.d_in(u_ca_in_462), .d_out(u_ca_out_462));
compressor_18_12 u_ca_18_12_463(.d_in(u_ca_in_463), .d_out(u_ca_out_463));
compressor_18_12 u_ca_18_12_464(.d_in(u_ca_in_464), .d_out(u_ca_out_464));
compressor_18_12 u_ca_18_12_465(.d_in(u_ca_in_465), .d_out(u_ca_out_465));
compressor_18_12 u_ca_18_12_466(.d_in(u_ca_in_466), .d_out(u_ca_out_466));
compressor_18_12 u_ca_18_12_467(.d_in(u_ca_in_467), .d_out(u_ca_out_467));
compressor_18_12 u_ca_18_12_468(.d_in(u_ca_in_468), .d_out(u_ca_out_468));
compressor_18_12 u_ca_18_12_469(.d_in(u_ca_in_469), .d_out(u_ca_out_469));
compressor_18_12 u_ca_18_12_470(.d_in(u_ca_in_470), .d_out(u_ca_out_470));
compressor_18_12 u_ca_18_12_471(.d_in(u_ca_in_471), .d_out(u_ca_out_471));
compressor_18_12 u_ca_18_12_472(.d_in(u_ca_in_472), .d_out(u_ca_out_472));
compressor_18_12 u_ca_18_12_473(.d_in(u_ca_in_473), .d_out(u_ca_out_473));
compressor_18_12 u_ca_18_12_474(.d_in(u_ca_in_474), .d_out(u_ca_out_474));
compressor_18_12 u_ca_18_12_475(.d_in(u_ca_in_475), .d_out(u_ca_out_475));
compressor_18_12 u_ca_18_12_476(.d_in(u_ca_in_476), .d_out(u_ca_out_476));
compressor_18_12 u_ca_18_12_477(.d_in(u_ca_in_477), .d_out(u_ca_out_477));
compressor_18_12 u_ca_18_12_478(.d_in(u_ca_in_478), .d_out(u_ca_out_478));
compressor_18_12 u_ca_18_12_479(.d_in(u_ca_in_479), .d_out(u_ca_out_479));
compressor_18_12 u_ca_18_12_480(.d_in(u_ca_in_480), .d_out(u_ca_out_480));
compressor_18_12 u_ca_18_12_481(.d_in(u_ca_in_481), .d_out(u_ca_out_481));
compressor_18_12 u_ca_18_12_482(.d_in(u_ca_in_482), .d_out(u_ca_out_482));
compressor_18_12 u_ca_18_12_483(.d_in(u_ca_in_483), .d_out(u_ca_out_483));
compressor_18_12 u_ca_18_12_484(.d_in(u_ca_in_484), .d_out(u_ca_out_484));
compressor_18_12 u_ca_18_12_485(.d_in(u_ca_in_485), .d_out(u_ca_out_485));
compressor_18_12 u_ca_18_12_486(.d_in(u_ca_in_486), .d_out(u_ca_out_486));
compressor_18_12 u_ca_18_12_487(.d_in(u_ca_in_487), .d_out(u_ca_out_487));
compressor_18_12 u_ca_18_12_488(.d_in(u_ca_in_488), .d_out(u_ca_out_488));
compressor_18_12 u_ca_18_12_489(.d_in(u_ca_in_489), .d_out(u_ca_out_489));
compressor_18_12 u_ca_18_12_490(.d_in(u_ca_in_490), .d_out(u_ca_out_490));
compressor_18_12 u_ca_18_12_491(.d_in(u_ca_in_491), .d_out(u_ca_out_491));
compressor_18_12 u_ca_18_12_492(.d_in(u_ca_in_492), .d_out(u_ca_out_492));
compressor_18_12 u_ca_18_12_493(.d_in(u_ca_in_493), .d_out(u_ca_out_493));
compressor_18_12 u_ca_18_12_494(.d_in(u_ca_in_494), .d_out(u_ca_out_494));
compressor_18_12 u_ca_18_12_495(.d_in(u_ca_in_495), .d_out(u_ca_out_495));
compressor_18_12 u_ca_18_12_496(.d_in(u_ca_in_496), .d_out(u_ca_out_496));
compressor_18_12 u_ca_18_12_497(.d_in(u_ca_in_497), .d_out(u_ca_out_497));
compressor_18_12 u_ca_18_12_498(.d_in(u_ca_in_498), .d_out(u_ca_out_498));
compressor_18_12 u_ca_18_12_499(.d_in(u_ca_in_499), .d_out(u_ca_out_499));
compressor_18_12 u_ca_18_12_500(.d_in(u_ca_in_500), .d_out(u_ca_out_500));
compressor_18_12 u_ca_18_12_501(.d_in(u_ca_in_501), .d_out(u_ca_out_501));
compressor_18_12 u_ca_18_12_502(.d_in(u_ca_in_502), .d_out(u_ca_out_502));
compressor_18_12 u_ca_18_12_503(.d_in(u_ca_in_503), .d_out(u_ca_out_503));
compressor_18_12 u_ca_18_12_504(.d_in(u_ca_in_504), .d_out(u_ca_out_504));
compressor_18_12 u_ca_18_12_505(.d_in(u_ca_in_505), .d_out(u_ca_out_505));
compressor_18_12 u_ca_18_12_506(.d_in(u_ca_in_506), .d_out(u_ca_out_506));
compressor_18_12 u_ca_18_12_507(.d_in(u_ca_in_507), .d_out(u_ca_out_507));
compressor_18_12 u_ca_18_12_508(.d_in(u_ca_in_508), .d_out(u_ca_out_508));
compressor_18_12 u_ca_18_12_509(.d_in(u_ca_in_509), .d_out(u_ca_out_509));
compressor_18_12 u_ca_18_12_510(.d_in(u_ca_in_510), .d_out(u_ca_out_510));
compressor_18_12 u_ca_18_12_511(.d_in(u_ca_in_511), .d_out(u_ca_out_511));
compressor_18_12 u_ca_18_12_512(.d_in(u_ca_in_512), .d_out(u_ca_out_512));
compressor_18_12 u_ca_18_12_513(.d_in(u_ca_in_513), .d_out(u_ca_out_513));
compressor_18_12 u_ca_18_12_514(.d_in(u_ca_in_514), .d_out(u_ca_out_514));
compressor_18_12 u_ca_18_12_515(.d_in(u_ca_in_515), .d_out(u_ca_out_515));
compressor_18_12 u_ca_18_12_516(.d_in(u_ca_in_516), .d_out(u_ca_out_516));
compressor_18_12 u_ca_18_12_517(.d_in(u_ca_in_517), .d_out(u_ca_out_517));
compressor_18_12 u_ca_18_12_518(.d_in(u_ca_in_518), .d_out(u_ca_out_518));
compressor_18_12 u_ca_18_12_519(.d_in(u_ca_in_519), .d_out(u_ca_out_519));
compressor_18_12 u_ca_18_12_520(.d_in(u_ca_in_520), .d_out(u_ca_out_520));
compressor_18_12 u_ca_18_12_521(.d_in(u_ca_in_521), .d_out(u_ca_out_521));
compressor_18_12 u_ca_18_12_522(.d_in(u_ca_in_522), .d_out(u_ca_out_522));
compressor_18_12 u_ca_18_12_523(.d_in(u_ca_in_523), .d_out(u_ca_out_523));
compressor_18_12 u_ca_18_12_524(.d_in(u_ca_in_524), .d_out(u_ca_out_524));
compressor_18_12 u_ca_18_12_525(.d_in(u_ca_in_525), .d_out(u_ca_out_525));
compressor_18_12 u_ca_18_12_526(.d_in(u_ca_in_526), .d_out(u_ca_out_526));
compressor_18_12 u_ca_18_12_527(.d_in(u_ca_in_527), .d_out(u_ca_out_527));
compressor_18_12 u_ca_18_12_528(.d_in(u_ca_in_528), .d_out(u_ca_out_528));
compressor_18_12 u_ca_18_12_529(.d_in(u_ca_in_529), .d_out(u_ca_out_529));
compressor_18_12 u_ca_18_12_530(.d_in(u_ca_in_530), .d_out(u_ca_out_530));
compressor_18_12 u_ca_18_12_531(.d_in(u_ca_in_531), .d_out(u_ca_out_531));
compressor_18_12 u_ca_18_12_532(.d_in(u_ca_in_532), .d_out(u_ca_out_532));
compressor_18_12 u_ca_18_12_533(.d_in(u_ca_in_533), .d_out(u_ca_out_533));
compressor_18_12 u_ca_18_12_534(.d_in(u_ca_in_534), .d_out(u_ca_out_534));
compressor_18_12 u_ca_18_12_535(.d_in(u_ca_in_535), .d_out(u_ca_out_535));
compressor_18_12 u_ca_18_12_536(.d_in(u_ca_in_536), .d_out(u_ca_out_536));
compressor_18_12 u_ca_18_12_537(.d_in(u_ca_in_537), .d_out(u_ca_out_537));
compressor_18_12 u_ca_18_12_538(.d_in(u_ca_in_538), .d_out(u_ca_out_538));
compressor_18_12 u_ca_18_12_539(.d_in(u_ca_in_539), .d_out(u_ca_out_539));
compressor_18_12 u_ca_18_12_540(.d_in(u_ca_in_540), .d_out(u_ca_out_540));
compressor_18_12 u_ca_18_12_541(.d_in(u_ca_in_541), .d_out(u_ca_out_541));
compressor_18_12 u_ca_18_12_542(.d_in(u_ca_in_542), .d_out(u_ca_out_542));
compressor_18_12 u_ca_18_12_543(.d_in(u_ca_in_543), .d_out(u_ca_out_543));
compressor_18_12 u_ca_18_12_544(.d_in(u_ca_in_544), .d_out(u_ca_out_544));
compressor_18_12 u_ca_18_12_545(.d_in(u_ca_in_545), .d_out(u_ca_out_545));
compressor_18_12 u_ca_18_12_546(.d_in(u_ca_in_546), .d_out(u_ca_out_546));
compressor_18_12 u_ca_18_12_547(.d_in(u_ca_in_547), .d_out(u_ca_out_547));
compressor_18_12 u_ca_18_12_548(.d_in(u_ca_in_548), .d_out(u_ca_out_548));
compressor_18_12 u_ca_18_12_549(.d_in(u_ca_in_549), .d_out(u_ca_out_549));
compressor_18_12 u_ca_18_12_550(.d_in(u_ca_in_550), .d_out(u_ca_out_550));
compressor_18_12 u_ca_18_12_551(.d_in(u_ca_in_551), .d_out(u_ca_out_551));
compressor_18_12 u_ca_18_12_552(.d_in(u_ca_in_552), .d_out(u_ca_out_552));
compressor_18_12 u_ca_18_12_553(.d_in(u_ca_in_553), .d_out(u_ca_out_553));
compressor_18_12 u_ca_18_12_554(.d_in(u_ca_in_554), .d_out(u_ca_out_554));
compressor_18_12 u_ca_18_12_555(.d_in(u_ca_in_555), .d_out(u_ca_out_555));
compressor_18_12 u_ca_18_12_556(.d_in(u_ca_in_556), .d_out(u_ca_out_556));
compressor_18_12 u_ca_18_12_557(.d_in(u_ca_in_557), .d_out(u_ca_out_557));
compressor_18_12 u_ca_18_12_558(.d_in(u_ca_in_558), .d_out(u_ca_out_558));
compressor_18_12 u_ca_18_12_559(.d_in(u_ca_in_559), .d_out(u_ca_out_559));
compressor_18_12 u_ca_18_12_560(.d_in(u_ca_in_560), .d_out(u_ca_out_560));
compressor_18_12 u_ca_18_12_561(.d_in(u_ca_in_561), .d_out(u_ca_out_561));
compressor_18_12 u_ca_18_12_562(.d_in(u_ca_in_562), .d_out(u_ca_out_562));
compressor_18_12 u_ca_18_12_563(.d_in(u_ca_in_563), .d_out(u_ca_out_563));
compressor_18_12 u_ca_18_12_564(.d_in(u_ca_in_564), .d_out(u_ca_out_564));
compressor_18_12 u_ca_18_12_565(.d_in(u_ca_in_565), .d_out(u_ca_out_565));
compressor_18_12 u_ca_18_12_566(.d_in(u_ca_in_566), .d_out(u_ca_out_566));
compressor_18_12 u_ca_18_12_567(.d_in(u_ca_in_567), .d_out(u_ca_out_567));
compressor_18_12 u_ca_18_12_568(.d_in(u_ca_in_568), .d_out(u_ca_out_568));
compressor_18_12 u_ca_18_12_569(.d_in(u_ca_in_569), .d_out(u_ca_out_569));
compressor_18_12 u_ca_18_12_570(.d_in(u_ca_in_570), .d_out(u_ca_out_570));
compressor_18_12 u_ca_18_12_571(.d_in(u_ca_in_571), .d_out(u_ca_out_571));
compressor_18_12 u_ca_18_12_572(.d_in(u_ca_in_572), .d_out(u_ca_out_572));
compressor_18_12 u_ca_18_12_573(.d_in(u_ca_in_573), .d_out(u_ca_out_573));
compressor_18_12 u_ca_18_12_574(.d_in(u_ca_in_574), .d_out(u_ca_out_574));
compressor_18_12 u_ca_18_12_575(.d_in(u_ca_in_575), .d_out(u_ca_out_575));
compressor_18_12 u_ca_18_12_576(.d_in(u_ca_in_576), .d_out(u_ca_out_576));
compressor_18_12 u_ca_18_12_577(.d_in(u_ca_in_577), .d_out(u_ca_out_577));
compressor_18_12 u_ca_18_12_578(.d_in(u_ca_in_578), .d_out(u_ca_out_578));
compressor_18_12 u_ca_18_12_579(.d_in(u_ca_in_579), .d_out(u_ca_out_579));
compressor_18_12 u_ca_18_12_580(.d_in(u_ca_in_580), .d_out(u_ca_out_580));
compressor_18_12 u_ca_18_12_581(.d_in(u_ca_in_581), .d_out(u_ca_out_581));
compressor_18_12 u_ca_18_12_582(.d_in(u_ca_in_582), .d_out(u_ca_out_582));
compressor_18_12 u_ca_18_12_583(.d_in(u_ca_in_583), .d_out(u_ca_out_583));
compressor_18_12 u_ca_18_12_584(.d_in(u_ca_in_584), .d_out(u_ca_out_584));
compressor_18_12 u_ca_18_12_585(.d_in(u_ca_in_585), .d_out(u_ca_out_585));
compressor_18_12 u_ca_18_12_586(.d_in(u_ca_in_586), .d_out(u_ca_out_586));
compressor_18_12 u_ca_18_12_587(.d_in(u_ca_in_587), .d_out(u_ca_out_587));
compressor_18_12 u_ca_18_12_588(.d_in(u_ca_in_588), .d_out(u_ca_out_588));
compressor_18_12 u_ca_18_12_589(.d_in(u_ca_in_589), .d_out(u_ca_out_589));
compressor_18_12 u_ca_18_12_590(.d_in(u_ca_in_590), .d_out(u_ca_out_590));
compressor_18_12 u_ca_18_12_591(.d_in(u_ca_in_591), .d_out(u_ca_out_591));
compressor_18_12 u_ca_18_12_592(.d_in(u_ca_in_592), .d_out(u_ca_out_592));
compressor_18_12 u_ca_18_12_593(.d_in(u_ca_in_593), .d_out(u_ca_out_593));
compressor_18_12 u_ca_18_12_594(.d_in(u_ca_in_594), .d_out(u_ca_out_594));
compressor_18_12 u_ca_18_12_595(.d_in(u_ca_in_595), .d_out(u_ca_out_595));
compressor_18_12 u_ca_18_12_596(.d_in(u_ca_in_596), .d_out(u_ca_out_596));
compressor_18_12 u_ca_18_12_597(.d_in(u_ca_in_597), .d_out(u_ca_out_597));
compressor_18_12 u_ca_18_12_598(.d_in(u_ca_in_598), .d_out(u_ca_out_598));
compressor_18_12 u_ca_18_12_599(.d_in(u_ca_in_599), .d_out(u_ca_out_599));
compressor_18_12 u_ca_18_12_600(.d_in(u_ca_in_600), .d_out(u_ca_out_600));
compressor_18_12 u_ca_18_12_601(.d_in(u_ca_in_601), .d_out(u_ca_out_601));
compressor_18_12 u_ca_18_12_602(.d_in(u_ca_in_602), .d_out(u_ca_out_602));
compressor_18_12 u_ca_18_12_603(.d_in(u_ca_in_603), .d_out(u_ca_out_603));
compressor_18_12 u_ca_18_12_604(.d_in(u_ca_in_604), .d_out(u_ca_out_604));
compressor_18_12 u_ca_18_12_605(.d_in(u_ca_in_605), .d_out(u_ca_out_605));
compressor_18_12 u_ca_18_12_606(.d_in(u_ca_in_606), .d_out(u_ca_out_606));
compressor_18_12 u_ca_18_12_607(.d_in(u_ca_in_607), .d_out(u_ca_out_607));
compressor_18_12 u_ca_18_12_608(.d_in(u_ca_in_608), .d_out(u_ca_out_608));
compressor_18_12 u_ca_18_12_609(.d_in(u_ca_in_609), .d_out(u_ca_out_609));
compressor_18_12 u_ca_18_12_610(.d_in(u_ca_in_610), .d_out(u_ca_out_610));
compressor_18_12 u_ca_18_12_611(.d_in(u_ca_in_611), .d_out(u_ca_out_611));
compressor_18_12 u_ca_18_12_612(.d_in(u_ca_in_612), .d_out(u_ca_out_612));
compressor_18_12 u_ca_18_12_613(.d_in(u_ca_in_613), .d_out(u_ca_out_613));
compressor_18_12 u_ca_18_12_614(.d_in(u_ca_in_614), .d_out(u_ca_out_614));
compressor_18_12 u_ca_18_12_615(.d_in(u_ca_in_615), .d_out(u_ca_out_615));
compressor_18_12 u_ca_18_12_616(.d_in(u_ca_in_616), .d_out(u_ca_out_616));
compressor_18_12 u_ca_18_12_617(.d_in(u_ca_in_617), .d_out(u_ca_out_617));
compressor_18_12 u_ca_18_12_618(.d_in(u_ca_in_618), .d_out(u_ca_out_618));
compressor_18_12 u_ca_18_12_619(.d_in(u_ca_in_619), .d_out(u_ca_out_619));
compressor_18_12 u_ca_18_12_620(.d_in(u_ca_in_620), .d_out(u_ca_out_620));
compressor_18_12 u_ca_18_12_621(.d_in(u_ca_in_621), .d_out(u_ca_out_621));
compressor_18_12 u_ca_18_12_622(.d_in(u_ca_in_622), .d_out(u_ca_out_622));
compressor_18_12 u_ca_18_12_623(.d_in(u_ca_in_623), .d_out(u_ca_out_623));
compressor_18_12 u_ca_18_12_624(.d_in(u_ca_in_624), .d_out(u_ca_out_624));
compressor_18_12 u_ca_18_12_625(.d_in(u_ca_in_625), .d_out(u_ca_out_625));
compressor_18_12 u_ca_18_12_626(.d_in(u_ca_in_626), .d_out(u_ca_out_626));
compressor_18_12 u_ca_18_12_627(.d_in(u_ca_in_627), .d_out(u_ca_out_627));
compressor_18_12 u_ca_18_12_628(.d_in(u_ca_in_628), .d_out(u_ca_out_628));
compressor_18_12 u_ca_18_12_629(.d_in(u_ca_in_629), .d_out(u_ca_out_629));
compressor_18_12 u_ca_18_12_630(.d_in(u_ca_in_630), .d_out(u_ca_out_630));
compressor_18_12 u_ca_18_12_631(.d_in(u_ca_in_631), .d_out(u_ca_out_631));
compressor_18_12 u_ca_18_12_632(.d_in(u_ca_in_632), .d_out(u_ca_out_632));
compressor_18_12 u_ca_18_12_633(.d_in(u_ca_in_633), .d_out(u_ca_out_633));
compressor_18_12 u_ca_18_12_634(.d_in(u_ca_in_634), .d_out(u_ca_out_634));
compressor_18_12 u_ca_18_12_635(.d_in(u_ca_in_635), .d_out(u_ca_out_635));
compressor_18_12 u_ca_18_12_636(.d_in(u_ca_in_636), .d_out(u_ca_out_636));
compressor_18_12 u_ca_18_12_637(.d_in(u_ca_in_637), .d_out(u_ca_out_637));
compressor_18_12 u_ca_18_12_638(.d_in(u_ca_in_638), .d_out(u_ca_out_638));
compressor_18_12 u_ca_18_12_639(.d_in(u_ca_in_639), .d_out(u_ca_out_639));
compressor_18_12 u_ca_18_12_640(.d_in(u_ca_in_640), .d_out(u_ca_out_640));
compressor_18_12 u_ca_18_12_641(.d_in(u_ca_in_641), .d_out(u_ca_out_641));
compressor_18_12 u_ca_18_12_642(.d_in(u_ca_in_642), .d_out(u_ca_out_642));
compressor_18_12 u_ca_18_12_643(.d_in(u_ca_in_643), .d_out(u_ca_out_643));
compressor_18_12 u_ca_18_12_644(.d_in(u_ca_in_644), .d_out(u_ca_out_644));
compressor_18_12 u_ca_18_12_645(.d_in(u_ca_in_645), .d_out(u_ca_out_645));
compressor_18_12 u_ca_18_12_646(.d_in(u_ca_in_646), .d_out(u_ca_out_646));
compressor_18_12 u_ca_18_12_647(.d_in(u_ca_in_647), .d_out(u_ca_out_647));
compressor_18_12 u_ca_18_12_648(.d_in(u_ca_in_648), .d_out(u_ca_out_648));
compressor_18_12 u_ca_18_12_649(.d_in(u_ca_in_649), .d_out(u_ca_out_649));
compressor_18_12 u_ca_18_12_650(.d_in(u_ca_in_650), .d_out(u_ca_out_650));
compressor_18_12 u_ca_18_12_651(.d_in(u_ca_in_651), .d_out(u_ca_out_651));
compressor_18_12 u_ca_18_12_652(.d_in(u_ca_in_652), .d_out(u_ca_out_652));
compressor_18_12 u_ca_18_12_653(.d_in(u_ca_in_653), .d_out(u_ca_out_653));
compressor_18_12 u_ca_18_12_654(.d_in(u_ca_in_654), .d_out(u_ca_out_654));
compressor_18_12 u_ca_18_12_655(.d_in(u_ca_in_655), .d_out(u_ca_out_655));
compressor_18_12 u_ca_18_12_656(.d_in(u_ca_in_656), .d_out(u_ca_out_656));
compressor_18_12 u_ca_18_12_657(.d_in(u_ca_in_657), .d_out(u_ca_out_657));
compressor_18_12 u_ca_18_12_658(.d_in(u_ca_in_658), .d_out(u_ca_out_658));
compressor_18_12 u_ca_18_12_659(.d_in(u_ca_in_659), .d_out(u_ca_out_659));
compressor_18_12 u_ca_18_12_660(.d_in(u_ca_in_660), .d_out(u_ca_out_660));
compressor_18_12 u_ca_18_12_661(.d_in(u_ca_in_661), .d_out(u_ca_out_661));
compressor_18_12 u_ca_18_12_662(.d_in(u_ca_in_662), .d_out(u_ca_out_662));
compressor_18_12 u_ca_18_12_663(.d_in(u_ca_in_663), .d_out(u_ca_out_663));
compressor_18_12 u_ca_18_12_664(.d_in(u_ca_in_664), .d_out(u_ca_out_664));
compressor_18_12 u_ca_18_12_665(.d_in(u_ca_in_665), .d_out(u_ca_out_665));
compressor_18_12 u_ca_18_12_666(.d_in(u_ca_in_666), .d_out(u_ca_out_666));
compressor_18_12 u_ca_18_12_667(.d_in(u_ca_in_667), .d_out(u_ca_out_667));
compressor_18_12 u_ca_18_12_668(.d_in(u_ca_in_668), .d_out(u_ca_out_668));
compressor_18_12 u_ca_18_12_669(.d_in(u_ca_in_669), .d_out(u_ca_out_669));
compressor_18_12 u_ca_18_12_670(.d_in(u_ca_in_670), .d_out(u_ca_out_670));
compressor_18_12 u_ca_18_12_671(.d_in(u_ca_in_671), .d_out(u_ca_out_671));
compressor_18_12 u_ca_18_12_672(.d_in(u_ca_in_672), .d_out(u_ca_out_672));
compressor_18_12 u_ca_18_12_673(.d_in(u_ca_in_673), .d_out(u_ca_out_673));
compressor_18_12 u_ca_18_12_674(.d_in(u_ca_in_674), .d_out(u_ca_out_674));
compressor_18_12 u_ca_18_12_675(.d_in(u_ca_in_675), .d_out(u_ca_out_675));
compressor_18_12 u_ca_18_12_676(.d_in(u_ca_in_676), .d_out(u_ca_out_676));
compressor_18_12 u_ca_18_12_677(.d_in(u_ca_in_677), .d_out(u_ca_out_677));
compressor_18_12 u_ca_18_12_678(.d_in(u_ca_in_678), .d_out(u_ca_out_678));
compressor_18_12 u_ca_18_12_679(.d_in(u_ca_in_679), .d_out(u_ca_out_679));
compressor_18_12 u_ca_18_12_680(.d_in(u_ca_in_680), .d_out(u_ca_out_680));
compressor_18_12 u_ca_18_12_681(.d_in(u_ca_in_681), .d_out(u_ca_out_681));
compressor_18_12 u_ca_18_12_682(.d_in(u_ca_in_682), .d_out(u_ca_out_682));
compressor_18_12 u_ca_18_12_683(.d_in(u_ca_in_683), .d_out(u_ca_out_683));
compressor_18_12 u_ca_18_12_684(.d_in(u_ca_in_684), .d_out(u_ca_out_684));
compressor_18_12 u_ca_18_12_685(.d_in(u_ca_in_685), .d_out(u_ca_out_685));
compressor_18_12 u_ca_18_12_686(.d_in(u_ca_in_686), .d_out(u_ca_out_686));
compressor_18_12 u_ca_18_12_687(.d_in(u_ca_in_687), .d_out(u_ca_out_687));
compressor_18_12 u_ca_18_12_688(.d_in(u_ca_in_688), .d_out(u_ca_out_688));
compressor_18_12 u_ca_18_12_689(.d_in(u_ca_in_689), .d_out(u_ca_out_689));
compressor_18_12 u_ca_18_12_690(.d_in(u_ca_in_690), .d_out(u_ca_out_690));
compressor_18_12 u_ca_18_12_691(.d_in(u_ca_in_691), .d_out(u_ca_out_691));
compressor_18_12 u_ca_18_12_692(.d_in(u_ca_in_692), .d_out(u_ca_out_692));
compressor_18_12 u_ca_18_12_693(.d_in(u_ca_in_693), .d_out(u_ca_out_693));
compressor_18_12 u_ca_18_12_694(.d_in(u_ca_in_694), .d_out(u_ca_out_694));
compressor_18_12 u_ca_18_12_695(.d_in(u_ca_in_695), .d_out(u_ca_out_695));
compressor_18_12 u_ca_18_12_696(.d_in(u_ca_in_696), .d_out(u_ca_out_696));
compressor_18_12 u_ca_18_12_697(.d_in(u_ca_in_697), .d_out(u_ca_out_697));
compressor_18_12 u_ca_18_12_698(.d_in(u_ca_in_698), .d_out(u_ca_out_698));
compressor_18_12 u_ca_18_12_699(.d_in(u_ca_in_699), .d_out(u_ca_out_699));
compressor_18_12 u_ca_18_12_700(.d_in(u_ca_in_700), .d_out(u_ca_out_700));
compressor_18_12 u_ca_18_12_701(.d_in(u_ca_in_701), .d_out(u_ca_out_701));
compressor_18_12 u_ca_18_12_702(.d_in(u_ca_in_702), .d_out(u_ca_out_702));
compressor_18_12 u_ca_18_12_703(.d_in(u_ca_in_703), .d_out(u_ca_out_703));
compressor_18_12 u_ca_18_12_704(.d_in(u_ca_in_704), .d_out(u_ca_out_704));
compressor_18_12 u_ca_18_12_705(.d_in(u_ca_in_705), .d_out(u_ca_out_705));
compressor_18_12 u_ca_18_12_706(.d_in(u_ca_in_706), .d_out(u_ca_out_706));
compressor_18_12 u_ca_18_12_707(.d_in(u_ca_in_707), .d_out(u_ca_out_707));
compressor_18_12 u_ca_18_12_708(.d_in(u_ca_in_708), .d_out(u_ca_out_708));
compressor_18_12 u_ca_18_12_709(.d_in(u_ca_in_709), .d_out(u_ca_out_709));
compressor_18_12 u_ca_18_12_710(.d_in(u_ca_in_710), .d_out(u_ca_out_710));
compressor_18_12 u_ca_18_12_711(.d_in(u_ca_in_711), .d_out(u_ca_out_711));
compressor_18_12 u_ca_18_12_712(.d_in(u_ca_in_712), .d_out(u_ca_out_712));
compressor_18_12 u_ca_18_12_713(.d_in(u_ca_in_713), .d_out(u_ca_out_713));
compressor_18_12 u_ca_18_12_714(.d_in(u_ca_in_714), .d_out(u_ca_out_714));
compressor_18_12 u_ca_18_12_715(.d_in(u_ca_in_715), .d_out(u_ca_out_715));
compressor_18_12 u_ca_18_12_716(.d_in(u_ca_in_716), .d_out(u_ca_out_716));
compressor_18_12 u_ca_18_12_717(.d_in(u_ca_in_717), .d_out(u_ca_out_717));
compressor_18_12 u_ca_18_12_718(.d_in(u_ca_in_718), .d_out(u_ca_out_718));
compressor_18_12 u_ca_18_12_719(.d_in(u_ca_in_719), .d_out(u_ca_out_719));
compressor_18_12 u_ca_18_12_720(.d_in(u_ca_in_720), .d_out(u_ca_out_720));
compressor_18_12 u_ca_18_12_721(.d_in(u_ca_in_721), .d_out(u_ca_out_721));
compressor_18_12 u_ca_18_12_722(.d_in(u_ca_in_722), .d_out(u_ca_out_722));
compressor_18_12 u_ca_18_12_723(.d_in(u_ca_in_723), .d_out(u_ca_out_723));
compressor_18_12 u_ca_18_12_724(.d_in(u_ca_in_724), .d_out(u_ca_out_724));
compressor_18_12 u_ca_18_12_725(.d_in(u_ca_in_725), .d_out(u_ca_out_725));
compressor_18_12 u_ca_18_12_726(.d_in(u_ca_in_726), .d_out(u_ca_out_726));
compressor_18_12 u_ca_18_12_727(.d_in(u_ca_in_727), .d_out(u_ca_out_727));
compressor_18_12 u_ca_18_12_728(.d_in(u_ca_in_728), .d_out(u_ca_out_728));
compressor_18_12 u_ca_18_12_729(.d_in(u_ca_in_729), .d_out(u_ca_out_729));
compressor_18_12 u_ca_18_12_730(.d_in(u_ca_in_730), .d_out(u_ca_out_730));
compressor_18_12 u_ca_18_12_731(.d_in(u_ca_in_731), .d_out(u_ca_out_731));
compressor_18_12 u_ca_18_12_732(.d_in(u_ca_in_732), .d_out(u_ca_out_732));
compressor_18_12 u_ca_18_12_733(.d_in(u_ca_in_733), .d_out(u_ca_out_733));
compressor_18_12 u_ca_18_12_734(.d_in(u_ca_in_734), .d_out(u_ca_out_734));
compressor_18_12 u_ca_18_12_735(.d_in(u_ca_in_735), .d_out(u_ca_out_735));
compressor_18_12 u_ca_18_12_736(.d_in(u_ca_in_736), .d_out(u_ca_out_736));
compressor_18_12 u_ca_18_12_737(.d_in(u_ca_in_737), .d_out(u_ca_out_737));
compressor_18_12 u_ca_18_12_738(.d_in(u_ca_in_738), .d_out(u_ca_out_738));
compressor_18_12 u_ca_18_12_739(.d_in(u_ca_in_739), .d_out(u_ca_out_739));
compressor_18_12 u_ca_18_12_740(.d_in(u_ca_in_740), .d_out(u_ca_out_740));
compressor_18_12 u_ca_18_12_741(.d_in(u_ca_in_741), .d_out(u_ca_out_741));
compressor_18_12 u_ca_18_12_742(.d_in(u_ca_in_742), .d_out(u_ca_out_742));
compressor_18_12 u_ca_18_12_743(.d_in(u_ca_in_743), .d_out(u_ca_out_743));
compressor_18_12 u_ca_18_12_744(.d_in(u_ca_in_744), .d_out(u_ca_out_744));
compressor_18_12 u_ca_18_12_745(.d_in(u_ca_in_745), .d_out(u_ca_out_745));
compressor_18_12 u_ca_18_12_746(.d_in(u_ca_in_746), .d_out(u_ca_out_746));
compressor_18_12 u_ca_18_12_747(.d_in(u_ca_in_747), .d_out(u_ca_out_747));
compressor_18_12 u_ca_18_12_748(.d_in(u_ca_in_748), .d_out(u_ca_out_748));
compressor_18_12 u_ca_18_12_749(.d_in(u_ca_in_749), .d_out(u_ca_out_749));
compressor_18_12 u_ca_18_12_750(.d_in(u_ca_in_750), .d_out(u_ca_out_750));
compressor_18_12 u_ca_18_12_751(.d_in(u_ca_in_751), .d_out(u_ca_out_751));
compressor_18_12 u_ca_18_12_752(.d_in(u_ca_in_752), .d_out(u_ca_out_752));
compressor_18_12 u_ca_18_12_753(.d_in(u_ca_in_753), .d_out(u_ca_out_753));
compressor_18_12 u_ca_18_12_754(.d_in(u_ca_in_754), .d_out(u_ca_out_754));
compressor_18_12 u_ca_18_12_755(.d_in(u_ca_in_755), .d_out(u_ca_out_755));
compressor_18_12 u_ca_18_12_756(.d_in(u_ca_in_756), .d_out(u_ca_out_756));
compressor_18_12 u_ca_18_12_757(.d_in(u_ca_in_757), .d_out(u_ca_out_757));
compressor_18_12 u_ca_18_12_758(.d_in(u_ca_in_758), .d_out(u_ca_out_758));
compressor_18_12 u_ca_18_12_759(.d_in(u_ca_in_759), .d_out(u_ca_out_759));
compressor_18_12 u_ca_18_12_760(.d_in(u_ca_in_760), .d_out(u_ca_out_760));
compressor_18_12 u_ca_18_12_761(.d_in(u_ca_in_761), .d_out(u_ca_out_761));
compressor_18_12 u_ca_18_12_762(.d_in(u_ca_in_762), .d_out(u_ca_out_762));
compressor_18_12 u_ca_18_12_763(.d_in(u_ca_in_763), .d_out(u_ca_out_763));
compressor_18_12 u_ca_18_12_764(.d_in(u_ca_in_764), .d_out(u_ca_out_764));
compressor_18_12 u_ca_18_12_765(.d_in(u_ca_in_765), .d_out(u_ca_out_765));
compressor_18_12 u_ca_18_12_766(.d_in(u_ca_in_766), .d_out(u_ca_out_766));
compressor_18_12 u_ca_18_12_767(.d_in(u_ca_in_767), .d_out(u_ca_out_767));
compressor_18_12 u_ca_18_12_768(.d_in(u_ca_in_768), .d_out(u_ca_out_768));
compressor_18_12 u_ca_18_12_769(.d_in(u_ca_in_769), .d_out(u_ca_out_769));
compressor_18_12 u_ca_18_12_770(.d_in(u_ca_in_770), .d_out(u_ca_out_770));
compressor_18_12 u_ca_18_12_771(.d_in(u_ca_in_771), .d_out(u_ca_out_771));
compressor_18_12 u_ca_18_12_772(.d_in(u_ca_in_772), .d_out(u_ca_out_772));
compressor_18_12 u_ca_18_12_773(.d_in(u_ca_in_773), .d_out(u_ca_out_773));
compressor_18_12 u_ca_18_12_774(.d_in(u_ca_in_774), .d_out(u_ca_out_774));
compressor_18_12 u_ca_18_12_775(.d_in(u_ca_in_775), .d_out(u_ca_out_775));
compressor_18_12 u_ca_18_12_776(.d_in(u_ca_in_776), .d_out(u_ca_out_776));
compressor_18_12 u_ca_18_12_777(.d_in(u_ca_in_777), .d_out(u_ca_out_777));
compressor_18_12 u_ca_18_12_778(.d_in(u_ca_in_778), .d_out(u_ca_out_778));
compressor_18_12 u_ca_18_12_779(.d_in(u_ca_in_779), .d_out(u_ca_out_779));
compressor_18_12 u_ca_18_12_780(.d_in(u_ca_in_780), .d_out(u_ca_out_780));
compressor_18_12 u_ca_18_12_781(.d_in(u_ca_in_781), .d_out(u_ca_out_781));
compressor_18_12 u_ca_18_12_782(.d_in(u_ca_in_782), .d_out(u_ca_out_782));
compressor_18_12 u_ca_18_12_783(.d_in(u_ca_in_783), .d_out(u_ca_out_783));
compressor_18_12 u_ca_18_12_784(.d_in(u_ca_in_784), .d_out(u_ca_out_784));
compressor_18_12 u_ca_18_12_785(.d_in(u_ca_in_785), .d_out(u_ca_out_785));
compressor_18_12 u_ca_18_12_786(.d_in(u_ca_in_786), .d_out(u_ca_out_786));
compressor_18_12 u_ca_18_12_787(.d_in(u_ca_in_787), .d_out(u_ca_out_787));
compressor_18_12 u_ca_18_12_788(.d_in(u_ca_in_788), .d_out(u_ca_out_788));
compressor_18_12 u_ca_18_12_789(.d_in(u_ca_in_789), .d_out(u_ca_out_789));
compressor_18_12 u_ca_18_12_790(.d_in(u_ca_in_790), .d_out(u_ca_out_790));
compressor_18_12 u_ca_18_12_791(.d_in(u_ca_in_791), .d_out(u_ca_out_791));
compressor_18_12 u_ca_18_12_792(.d_in(u_ca_in_792), .d_out(u_ca_out_792));
compressor_18_12 u_ca_18_12_793(.d_in(u_ca_in_793), .d_out(u_ca_out_793));
compressor_18_12 u_ca_18_12_794(.d_in(u_ca_in_794), .d_out(u_ca_out_794));
compressor_18_12 u_ca_18_12_795(.d_in(u_ca_in_795), .d_out(u_ca_out_795));
compressor_18_12 u_ca_18_12_796(.d_in(u_ca_in_796), .d_out(u_ca_out_796));
compressor_18_12 u_ca_18_12_797(.d_in(u_ca_in_797), .d_out(u_ca_out_797));
compressor_18_12 u_ca_18_12_798(.d_in(u_ca_in_798), .d_out(u_ca_out_798));
compressor_18_12 u_ca_18_12_799(.d_in(u_ca_in_799), .d_out(u_ca_out_799));
compressor_18_12 u_ca_18_12_800(.d_in(u_ca_in_800), .d_out(u_ca_out_800));
compressor_18_12 u_ca_18_12_801(.d_in(u_ca_in_801), .d_out(u_ca_out_801));
compressor_18_12 u_ca_18_12_802(.d_in(u_ca_in_802), .d_out(u_ca_out_802));
compressor_18_12 u_ca_18_12_803(.d_in(u_ca_in_803), .d_out(u_ca_out_803));
compressor_18_12 u_ca_18_12_804(.d_in(u_ca_in_804), .d_out(u_ca_out_804));
compressor_18_12 u_ca_18_12_805(.d_in(u_ca_in_805), .d_out(u_ca_out_805));
compressor_18_12 u_ca_18_12_806(.d_in(u_ca_in_806), .d_out(u_ca_out_806));
compressor_18_12 u_ca_18_12_807(.d_in(u_ca_in_807), .d_out(u_ca_out_807));
compressor_18_12 u_ca_18_12_808(.d_in(u_ca_in_808), .d_out(u_ca_out_808));
compressor_18_12 u_ca_18_12_809(.d_in(u_ca_in_809), .d_out(u_ca_out_809));
compressor_18_12 u_ca_18_12_810(.d_in(u_ca_in_810), .d_out(u_ca_out_810));
compressor_18_12 u_ca_18_12_811(.d_in(u_ca_in_811), .d_out(u_ca_out_811));
compressor_18_12 u_ca_18_12_812(.d_in(u_ca_in_812), .d_out(u_ca_out_812));
compressor_18_12 u_ca_18_12_813(.d_in(u_ca_in_813), .d_out(u_ca_out_813));
compressor_18_12 u_ca_18_12_814(.d_in(u_ca_in_814), .d_out(u_ca_out_814));
compressor_18_12 u_ca_18_12_815(.d_in(u_ca_in_815), .d_out(u_ca_out_815));
compressor_18_12 u_ca_18_12_816(.d_in(u_ca_in_816), .d_out(u_ca_out_816));
compressor_18_12 u_ca_18_12_817(.d_in(u_ca_in_817), .d_out(u_ca_out_817));
compressor_18_12 u_ca_18_12_818(.d_in(u_ca_in_818), .d_out(u_ca_out_818));
compressor_18_12 u_ca_18_12_819(.d_in(u_ca_in_819), .d_out(u_ca_out_819));
compressor_18_12 u_ca_18_12_820(.d_in(u_ca_in_820), .d_out(u_ca_out_820));
compressor_18_12 u_ca_18_12_821(.d_in(u_ca_in_821), .d_out(u_ca_out_821));
compressor_18_12 u_ca_18_12_822(.d_in(u_ca_in_822), .d_out(u_ca_out_822));
compressor_18_12 u_ca_18_12_823(.d_in(u_ca_in_823), .d_out(u_ca_out_823));
compressor_18_12 u_ca_18_12_824(.d_in(u_ca_in_824), .d_out(u_ca_out_824));
compressor_18_12 u_ca_18_12_825(.d_in(u_ca_in_825), .d_out(u_ca_out_825));
compressor_18_12 u_ca_18_12_826(.d_in(u_ca_in_826), .d_out(u_ca_out_826));
compressor_18_12 u_ca_18_12_827(.d_in(u_ca_in_827), .d_out(u_ca_out_827));
compressor_18_12 u_ca_18_12_828(.d_in(u_ca_in_828), .d_out(u_ca_out_828));
compressor_18_12 u_ca_18_12_829(.d_in(u_ca_in_829), .d_out(u_ca_out_829));
compressor_18_12 u_ca_18_12_830(.d_in(u_ca_in_830), .d_out(u_ca_out_830));
compressor_18_12 u_ca_18_12_831(.d_in(u_ca_in_831), .d_out(u_ca_out_831));
compressor_18_12 u_ca_18_12_832(.d_in(u_ca_in_832), .d_out(u_ca_out_832));
compressor_18_12 u_ca_18_12_833(.d_in(u_ca_in_833), .d_out(u_ca_out_833));
compressor_18_12 u_ca_18_12_834(.d_in(u_ca_in_834), .d_out(u_ca_out_834));
compressor_18_12 u_ca_18_12_835(.d_in(u_ca_in_835), .d_out(u_ca_out_835));
compressor_18_12 u_ca_18_12_836(.d_in(u_ca_in_836), .d_out(u_ca_out_836));
compressor_18_12 u_ca_18_12_837(.d_in(u_ca_in_837), .d_out(u_ca_out_837));
compressor_18_12 u_ca_18_12_838(.d_in(u_ca_in_838), .d_out(u_ca_out_838));
compressor_18_12 u_ca_18_12_839(.d_in(u_ca_in_839), .d_out(u_ca_out_839));
compressor_18_12 u_ca_18_12_840(.d_in(u_ca_in_840), .d_out(u_ca_out_840));
compressor_18_12 u_ca_18_12_841(.d_in(u_ca_in_841), .d_out(u_ca_out_841));
compressor_18_12 u_ca_18_12_842(.d_in(u_ca_in_842), .d_out(u_ca_out_842));
compressor_18_12 u_ca_18_12_843(.d_in(u_ca_in_843), .d_out(u_ca_out_843));
compressor_18_12 u_ca_18_12_844(.d_in(u_ca_in_844), .d_out(u_ca_out_844));
compressor_18_12 u_ca_18_12_845(.d_in(u_ca_in_845), .d_out(u_ca_out_845));
compressor_18_12 u_ca_18_12_846(.d_in(u_ca_in_846), .d_out(u_ca_out_846));
compressor_18_12 u_ca_18_12_847(.d_in(u_ca_in_847), .d_out(u_ca_out_847));
compressor_18_12 u_ca_18_12_848(.d_in(u_ca_in_848), .d_out(u_ca_out_848));
compressor_18_12 u_ca_18_12_849(.d_in(u_ca_in_849), .d_out(u_ca_out_849));
compressor_18_12 u_ca_18_12_850(.d_in(u_ca_in_850), .d_out(u_ca_out_850));
compressor_18_12 u_ca_18_12_851(.d_in(u_ca_in_851), .d_out(u_ca_out_851));
compressor_18_12 u_ca_18_12_852(.d_in(u_ca_in_852), .d_out(u_ca_out_852));
compressor_18_12 u_ca_18_12_853(.d_in(u_ca_in_853), .d_out(u_ca_out_853));
compressor_18_12 u_ca_18_12_854(.d_in(u_ca_in_854), .d_out(u_ca_out_854));
compressor_18_12 u_ca_18_12_855(.d_in(u_ca_in_855), .d_out(u_ca_out_855));
compressor_18_12 u_ca_18_12_856(.d_in(u_ca_in_856), .d_out(u_ca_out_856));
compressor_18_12 u_ca_18_12_857(.d_in(u_ca_in_857), .d_out(u_ca_out_857));
compressor_18_12 u_ca_18_12_858(.d_in(u_ca_in_858), .d_out(u_ca_out_858));
compressor_18_12 u_ca_18_12_859(.d_in(u_ca_in_859), .d_out(u_ca_out_859));
compressor_18_12 u_ca_18_12_860(.d_in(u_ca_in_860), .d_out(u_ca_out_860));
compressor_18_12 u_ca_18_12_861(.d_in(u_ca_in_861), .d_out(u_ca_out_861));
compressor_18_12 u_ca_18_12_862(.d_in(u_ca_in_862), .d_out(u_ca_out_862));
compressor_18_12 u_ca_18_12_863(.d_in(u_ca_in_863), .d_out(u_ca_out_863));
compressor_18_12 u_ca_18_12_864(.d_in(u_ca_in_864), .d_out(u_ca_out_864));
compressor_18_12 u_ca_18_12_865(.d_in(u_ca_in_865), .d_out(u_ca_out_865));
compressor_18_12 u_ca_18_12_866(.d_in(u_ca_in_866), .d_out(u_ca_out_866));
compressor_18_12 u_ca_18_12_867(.d_in(u_ca_in_867), .d_out(u_ca_out_867));
compressor_18_12 u_ca_18_12_868(.d_in(u_ca_in_868), .d_out(u_ca_out_868));
compressor_18_12 u_ca_18_12_869(.d_in(u_ca_in_869), .d_out(u_ca_out_869));
compressor_18_12 u_ca_18_12_870(.d_in(u_ca_in_870), .d_out(u_ca_out_870));
compressor_18_12 u_ca_18_12_871(.d_in(u_ca_in_871), .d_out(u_ca_out_871));
compressor_18_12 u_ca_18_12_872(.d_in(u_ca_in_872), .d_out(u_ca_out_872));
compressor_18_12 u_ca_18_12_873(.d_in(u_ca_in_873), .d_out(u_ca_out_873));
compressor_18_12 u_ca_18_12_874(.d_in(u_ca_in_874), .d_out(u_ca_out_874));
compressor_18_12 u_ca_18_12_875(.d_in(u_ca_in_875), .d_out(u_ca_out_875));
compressor_18_12 u_ca_18_12_876(.d_in(u_ca_in_876), .d_out(u_ca_out_876));
compressor_18_12 u_ca_18_12_877(.d_in(u_ca_in_877), .d_out(u_ca_out_877));
compressor_18_12 u_ca_18_12_878(.d_in(u_ca_in_878), .d_out(u_ca_out_878));
compressor_18_12 u_ca_18_12_879(.d_in(u_ca_in_879), .d_out(u_ca_out_879));
compressor_18_12 u_ca_18_12_880(.d_in(u_ca_in_880), .d_out(u_ca_out_880));
compressor_18_12 u_ca_18_12_881(.d_in(u_ca_in_881), .d_out(u_ca_out_881));
compressor_18_12 u_ca_18_12_882(.d_in(u_ca_in_882), .d_out(u_ca_out_882));
compressor_18_12 u_ca_18_12_883(.d_in(u_ca_in_883), .d_out(u_ca_out_883));
compressor_18_12 u_ca_18_12_884(.d_in(u_ca_in_884), .d_out(u_ca_out_884));
compressor_18_12 u_ca_18_12_885(.d_in(u_ca_in_885), .d_out(u_ca_out_885));
compressor_18_12 u_ca_18_12_886(.d_in(u_ca_in_886), .d_out(u_ca_out_886));
compressor_18_12 u_ca_18_12_887(.d_in(u_ca_in_887), .d_out(u_ca_out_887));
compressor_18_12 u_ca_18_12_888(.d_in(u_ca_in_888), .d_out(u_ca_out_888));
compressor_18_12 u_ca_18_12_889(.d_in(u_ca_in_889), .d_out(u_ca_out_889));
compressor_18_12 u_ca_18_12_890(.d_in(u_ca_in_890), .d_out(u_ca_out_890));
compressor_18_12 u_ca_18_12_891(.d_in(u_ca_in_891), .d_out(u_ca_out_891));
compressor_18_12 u_ca_18_12_892(.d_in(u_ca_in_892), .d_out(u_ca_out_892));
compressor_18_12 u_ca_18_12_893(.d_in(u_ca_in_893), .d_out(u_ca_out_893));
compressor_18_12 u_ca_18_12_894(.d_in(u_ca_in_894), .d_out(u_ca_out_894));
compressor_18_12 u_ca_18_12_895(.d_in(u_ca_in_895), .d_out(u_ca_out_895));
compressor_18_12 u_ca_18_12_896(.d_in(u_ca_in_896), .d_out(u_ca_out_896));
compressor_18_12 u_ca_18_12_897(.d_in(u_ca_in_897), .d_out(u_ca_out_897));
compressor_18_12 u_ca_18_12_898(.d_in(u_ca_in_898), .d_out(u_ca_out_898));
compressor_18_12 u_ca_18_12_899(.d_in(u_ca_in_899), .d_out(u_ca_out_899));
compressor_18_12 u_ca_18_12_900(.d_in(u_ca_in_900), .d_out(u_ca_out_900));
compressor_18_12 u_ca_18_12_901(.d_in(u_ca_in_901), .d_out(u_ca_out_901));
compressor_18_12 u_ca_18_12_902(.d_in(u_ca_in_902), .d_out(u_ca_out_902));
compressor_18_12 u_ca_18_12_903(.d_in(u_ca_in_903), .d_out(u_ca_out_903));
compressor_18_12 u_ca_18_12_904(.d_in(u_ca_in_904), .d_out(u_ca_out_904));
compressor_18_12 u_ca_18_12_905(.d_in(u_ca_in_905), .d_out(u_ca_out_905));
compressor_18_12 u_ca_18_12_906(.d_in(u_ca_in_906), .d_out(u_ca_out_906));
compressor_18_12 u_ca_18_12_907(.d_in(u_ca_in_907), .d_out(u_ca_out_907));
compressor_18_12 u_ca_18_12_908(.d_in(u_ca_in_908), .d_out(u_ca_out_908));
compressor_18_12 u_ca_18_12_909(.d_in(u_ca_in_909), .d_out(u_ca_out_909));
compressor_18_12 u_ca_18_12_910(.d_in(u_ca_in_910), .d_out(u_ca_out_910));
compressor_18_12 u_ca_18_12_911(.d_in(u_ca_in_911), .d_out(u_ca_out_911));
compressor_18_12 u_ca_18_12_912(.d_in(u_ca_in_912), .d_out(u_ca_out_912));
compressor_18_12 u_ca_18_12_913(.d_in(u_ca_in_913), .d_out(u_ca_out_913));
compressor_18_12 u_ca_18_12_914(.d_in(u_ca_in_914), .d_out(u_ca_out_914));
compressor_18_12 u_ca_18_12_915(.d_in(u_ca_in_915), .d_out(u_ca_out_915));
compressor_18_12 u_ca_18_12_916(.d_in(u_ca_in_916), .d_out(u_ca_out_916));
compressor_18_12 u_ca_18_12_917(.d_in(u_ca_in_917), .d_out(u_ca_out_917));
compressor_18_12 u_ca_18_12_918(.d_in(u_ca_in_918), .d_out(u_ca_out_918));
compressor_18_12 u_ca_18_12_919(.d_in(u_ca_in_919), .d_out(u_ca_out_919));
compressor_18_12 u_ca_18_12_920(.d_in(u_ca_in_920), .d_out(u_ca_out_920));
compressor_18_12 u_ca_18_12_921(.d_in(u_ca_in_921), .d_out(u_ca_out_921));
compressor_18_12 u_ca_18_12_922(.d_in(u_ca_in_922), .d_out(u_ca_out_922));
compressor_18_12 u_ca_18_12_923(.d_in(u_ca_in_923), .d_out(u_ca_out_923));
compressor_18_12 u_ca_18_12_924(.d_in(u_ca_in_924), .d_out(u_ca_out_924));
compressor_18_12 u_ca_18_12_925(.d_in(u_ca_in_925), .d_out(u_ca_out_925));
compressor_18_12 u_ca_18_12_926(.d_in(u_ca_in_926), .d_out(u_ca_out_926));
compressor_18_12 u_ca_18_12_927(.d_in(u_ca_in_927), .d_out(u_ca_out_927));
compressor_18_12 u_ca_18_12_928(.d_in(u_ca_in_928), .d_out(u_ca_out_928));
compressor_18_12 u_ca_18_12_929(.d_in(u_ca_in_929), .d_out(u_ca_out_929));
compressor_18_12 u_ca_18_12_930(.d_in(u_ca_in_930), .d_out(u_ca_out_930));
compressor_18_12 u_ca_18_12_931(.d_in(u_ca_in_931), .d_out(u_ca_out_931));
compressor_18_12 u_ca_18_12_932(.d_in(u_ca_in_932), .d_out(u_ca_out_932));
compressor_18_12 u_ca_18_12_933(.d_in(u_ca_in_933), .d_out(u_ca_out_933));
compressor_18_12 u_ca_18_12_934(.d_in(u_ca_in_934), .d_out(u_ca_out_934));
compressor_18_12 u_ca_18_12_935(.d_in(u_ca_in_935), .d_out(u_ca_out_935));
compressor_18_12 u_ca_18_12_936(.d_in(u_ca_in_936), .d_out(u_ca_out_936));
compressor_18_12 u_ca_18_12_937(.d_in(u_ca_in_937), .d_out(u_ca_out_937));
compressor_18_12 u_ca_18_12_938(.d_in(u_ca_in_938), .d_out(u_ca_out_938));
compressor_18_12 u_ca_18_12_939(.d_in(u_ca_in_939), .d_out(u_ca_out_939));
compressor_18_12 u_ca_18_12_940(.d_in(u_ca_in_940), .d_out(u_ca_out_940));
compressor_18_12 u_ca_18_12_941(.d_in(u_ca_in_941), .d_out(u_ca_out_941));
compressor_18_12 u_ca_18_12_942(.d_in(u_ca_in_942), .d_out(u_ca_out_942));
compressor_18_12 u_ca_18_12_943(.d_in(u_ca_in_943), .d_out(u_ca_out_943));
compressor_18_12 u_ca_18_12_944(.d_in(u_ca_in_944), .d_out(u_ca_out_944));
compressor_18_12 u_ca_18_12_945(.d_in(u_ca_in_945), .d_out(u_ca_out_945));
compressor_18_12 u_ca_18_12_946(.d_in(u_ca_in_946), .d_out(u_ca_out_946));
compressor_18_12 u_ca_18_12_947(.d_in(u_ca_in_947), .d_out(u_ca_out_947));
compressor_18_12 u_ca_18_12_948(.d_in(u_ca_in_948), .d_out(u_ca_out_948));
compressor_18_12 u_ca_18_12_949(.d_in(u_ca_in_949), .d_out(u_ca_out_949));
compressor_18_12 u_ca_18_12_950(.d_in(u_ca_in_950), .d_out(u_ca_out_950));
compressor_18_12 u_ca_18_12_951(.d_in(u_ca_in_951), .d_out(u_ca_out_951));
compressor_18_12 u_ca_18_12_952(.d_in(u_ca_in_952), .d_out(u_ca_out_952));
compressor_18_12 u_ca_18_12_953(.d_in(u_ca_in_953), .d_out(u_ca_out_953));
compressor_18_12 u_ca_18_12_954(.d_in(u_ca_in_954), .d_out(u_ca_out_954));
compressor_18_12 u_ca_18_12_955(.d_in(u_ca_in_955), .d_out(u_ca_out_955));
compressor_18_12 u_ca_18_12_956(.d_in(u_ca_in_956), .d_out(u_ca_out_956));
compressor_18_12 u_ca_18_12_957(.d_in(u_ca_in_957), .d_out(u_ca_out_957));
compressor_18_12 u_ca_18_12_958(.d_in(u_ca_in_958), .d_out(u_ca_out_958));
compressor_18_12 u_ca_18_12_959(.d_in(u_ca_in_959), .d_out(u_ca_out_959));
compressor_18_12 u_ca_18_12_960(.d_in(u_ca_in_960), .d_out(u_ca_out_960));
compressor_18_12 u_ca_18_12_961(.d_in(u_ca_in_961), .d_out(u_ca_out_961));
compressor_18_12 u_ca_18_12_962(.d_in(u_ca_in_962), .d_out(u_ca_out_962));
compressor_18_12 u_ca_18_12_963(.d_in(u_ca_in_963), .d_out(u_ca_out_963));
compressor_18_12 u_ca_18_12_964(.d_in(u_ca_in_964), .d_out(u_ca_out_964));
compressor_18_12 u_ca_18_12_965(.d_in(u_ca_in_965), .d_out(u_ca_out_965));
compressor_18_12 u_ca_18_12_966(.d_in(u_ca_in_966), .d_out(u_ca_out_966));
compressor_18_12 u_ca_18_12_967(.d_in(u_ca_in_967), .d_out(u_ca_out_967));
compressor_18_12 u_ca_18_12_968(.d_in(u_ca_in_968), .d_out(u_ca_out_968));
compressor_18_12 u_ca_18_12_969(.d_in(u_ca_in_969), .d_out(u_ca_out_969));
compressor_18_12 u_ca_18_12_970(.d_in(u_ca_in_970), .d_out(u_ca_out_970));
compressor_18_12 u_ca_18_12_971(.d_in(u_ca_in_971), .d_out(u_ca_out_971));
compressor_18_12 u_ca_18_12_972(.d_in(u_ca_in_972), .d_out(u_ca_out_972));
compressor_18_12 u_ca_18_12_973(.d_in(u_ca_in_973), .d_out(u_ca_out_973));
compressor_18_12 u_ca_18_12_974(.d_in(u_ca_in_974), .d_out(u_ca_out_974));
compressor_18_12 u_ca_18_12_975(.d_in(u_ca_in_975), .d_out(u_ca_out_975));
compressor_18_12 u_ca_18_12_976(.d_in(u_ca_in_976), .d_out(u_ca_out_976));
compressor_18_12 u_ca_18_12_977(.d_in(u_ca_in_977), .d_out(u_ca_out_977));
compressor_18_12 u_ca_18_12_978(.d_in(u_ca_in_978), .d_out(u_ca_out_978));
compressor_18_12 u_ca_18_12_979(.d_in(u_ca_in_979), .d_out(u_ca_out_979));
compressor_18_12 u_ca_18_12_980(.d_in(u_ca_in_980), .d_out(u_ca_out_980));
compressor_18_12 u_ca_18_12_981(.d_in(u_ca_in_981), .d_out(u_ca_out_981));
compressor_18_12 u_ca_18_12_982(.d_in(u_ca_in_982), .d_out(u_ca_out_982));
compressor_18_12 u_ca_18_12_983(.d_in(u_ca_in_983), .d_out(u_ca_out_983));
compressor_18_12 u_ca_18_12_984(.d_in(u_ca_in_984), .d_out(u_ca_out_984));
compressor_18_12 u_ca_18_12_985(.d_in(u_ca_in_985), .d_out(u_ca_out_985));
compressor_18_12 u_ca_18_12_986(.d_in(u_ca_in_986), .d_out(u_ca_out_986));
compressor_18_12 u_ca_18_12_987(.d_in(u_ca_in_987), .d_out(u_ca_out_987));
compressor_18_12 u_ca_18_12_988(.d_in(u_ca_in_988), .d_out(u_ca_out_988));
compressor_18_12 u_ca_18_12_989(.d_in(u_ca_in_989), .d_out(u_ca_out_989));
compressor_18_12 u_ca_18_12_990(.d_in(u_ca_in_990), .d_out(u_ca_out_990));
compressor_18_12 u_ca_18_12_991(.d_in(u_ca_in_991), .d_out(u_ca_out_991));
compressor_18_12 u_ca_18_12_992(.d_in(u_ca_in_992), .d_out(u_ca_out_992));
compressor_18_12 u_ca_18_12_993(.d_in(u_ca_in_993), .d_out(u_ca_out_993));
compressor_18_12 u_ca_18_12_994(.d_in(u_ca_in_994), .d_out(u_ca_out_994));
compressor_18_12 u_ca_18_12_995(.d_in(u_ca_in_995), .d_out(u_ca_out_995));
compressor_18_12 u_ca_18_12_996(.d_in(u_ca_in_996), .d_out(u_ca_out_996));
compressor_18_12 u_ca_18_12_997(.d_in(u_ca_in_997), .d_out(u_ca_out_997));
compressor_18_12 u_ca_18_12_998(.d_in(u_ca_in_998), .d_out(u_ca_out_998));
compressor_18_12 u_ca_18_12_999(.d_in(u_ca_in_999), .d_out(u_ca_out_999));
compressor_18_12 u_ca_18_12_1000(.d_in(u_ca_in_1000), .d_out(u_ca_out_1000));
compressor_18_12 u_ca_18_12_1001(.d_in(u_ca_in_1001), .d_out(u_ca_out_1001));
compressor_18_12 u_ca_18_12_1002(.d_in(u_ca_in_1002), .d_out(u_ca_out_1002));
compressor_18_12 u_ca_18_12_1003(.d_in(u_ca_in_1003), .d_out(u_ca_out_1003));
compressor_18_12 u_ca_18_12_1004(.d_in(u_ca_in_1004), .d_out(u_ca_out_1004));
compressor_18_12 u_ca_18_12_1005(.d_in(u_ca_in_1005), .d_out(u_ca_out_1005));
compressor_18_12 u_ca_18_12_1006(.d_in(u_ca_in_1006), .d_out(u_ca_out_1006));
compressor_18_12 u_ca_18_12_1007(.d_in(u_ca_in_1007), .d_out(u_ca_out_1007));
compressor_18_12 u_ca_18_12_1008(.d_in(u_ca_in_1008), .d_out(u_ca_out_1008));
compressor_18_12 u_ca_18_12_1009(.d_in(u_ca_in_1009), .d_out(u_ca_out_1009));
compressor_18_12 u_ca_18_12_1010(.d_in(u_ca_in_1010), .d_out(u_ca_out_1010));
compressor_18_12 u_ca_18_12_1011(.d_in(u_ca_in_1011), .d_out(u_ca_out_1011));
compressor_18_12 u_ca_18_12_1012(.d_in(u_ca_in_1012), .d_out(u_ca_out_1012));
compressor_18_12 u_ca_18_12_1013(.d_in(u_ca_in_1013), .d_out(u_ca_out_1013));
compressor_18_12 u_ca_18_12_1014(.d_in(u_ca_in_1014), .d_out(u_ca_out_1014));
compressor_18_12 u_ca_18_12_1015(.d_in(u_ca_in_1015), .d_out(u_ca_out_1015));
compressor_18_12 u_ca_18_12_1016(.d_in(u_ca_in_1016), .d_out(u_ca_out_1016));
compressor_18_12 u_ca_18_12_1017(.d_in(u_ca_in_1017), .d_out(u_ca_out_1017));
compressor_18_12 u_ca_18_12_1018(.d_in(u_ca_in_1018), .d_out(u_ca_out_1018));
compressor_18_12 u_ca_18_12_1019(.d_in(u_ca_in_1019), .d_out(u_ca_out_1019));
compressor_18_12 u_ca_18_12_1020(.d_in(u_ca_in_1020), .d_out(u_ca_out_1020));
compressor_18_12 u_ca_18_12_1021(.d_in(u_ca_in_1021), .d_out(u_ca_out_1021));
compressor_18_12 u_ca_18_12_1022(.d_in(u_ca_in_1022), .d_out(u_ca_out_1022));
compressor_18_12 u_ca_18_12_1023(.d_in(u_ca_in_1023), .d_out(u_ca_out_1023));
compressor_18_12 u_ca_18_12_1024(.d_in(u_ca_in_1024), .d_out(u_ca_out_1024));
compressor_18_12 u_ca_18_12_1025(.d_in(u_ca_in_1025), .d_out(u_ca_out_1025));
compressor_18_12 u_ca_18_12_1026(.d_in(u_ca_in_1026), .d_out(u_ca_out_1026));
compressor_18_12 u_ca_18_12_1027(.d_in(u_ca_in_1027), .d_out(u_ca_out_1027));
compressor_18_12 u_ca_18_12_1028(.d_in(u_ca_in_1028), .d_out(u_ca_out_1028));
compressor_18_12 u_ca_18_12_1029(.d_in(u_ca_in_1029), .d_out(u_ca_out_1029));
compressor_18_12 u_ca_18_12_1030(.d_in(u_ca_in_1030), .d_out(u_ca_out_1030));
compressor_18_12 u_ca_18_12_1031(.d_in(u_ca_in_1031), .d_out(u_ca_out_1031));
compressor_18_12 u_ca_18_12_1032(.d_in(u_ca_in_1032), .d_out(u_ca_out_1032));

//---------------------------------------------------------



//--output-------------------------------------------------

assign col_out_0 = {{6{1'b0}}, u_ca_out_0[5:0]};
assign col_out_1 = {u_ca_out_1[5:0], u_ca_out_0[11:6]};
assign col_out_2 = {u_ca_out_2[5:0], u_ca_out_1[11:6]};
assign col_out_3 = {u_ca_out_3[5:0], u_ca_out_2[11:6]};
assign col_out_4 = {u_ca_out_4[5:0], u_ca_out_3[11:6]};
assign col_out_5 = {u_ca_out_5[5:0], u_ca_out_4[11:6]};
assign col_out_6 = {u_ca_out_6[5:0], u_ca_out_5[11:6]};
assign col_out_7 = {u_ca_out_7[5:0], u_ca_out_6[11:6]};
assign col_out_8 = {u_ca_out_8[5:0], u_ca_out_7[11:6]};
assign col_out_9 = {u_ca_out_9[5:0], u_ca_out_8[11:6]};
assign col_out_10 = {u_ca_out_10[5:0], u_ca_out_9[11:6]};
assign col_out_11 = {u_ca_out_11[5:0], u_ca_out_10[11:6]};
assign col_out_12 = {u_ca_out_12[5:0], u_ca_out_11[11:6]};
assign col_out_13 = {u_ca_out_13[5:0], u_ca_out_12[11:6]};
assign col_out_14 = {u_ca_out_14[5:0], u_ca_out_13[11:6]};
assign col_out_15 = {u_ca_out_15[5:0], u_ca_out_14[11:6]};
assign col_out_16 = {u_ca_out_16[5:0], u_ca_out_15[11:6]};
assign col_out_17 = {u_ca_out_17[5:0], u_ca_out_16[11:6]};
assign col_out_18 = {u_ca_out_18[5:0], u_ca_out_17[11:6]};
assign col_out_19 = {u_ca_out_19[5:0], u_ca_out_18[11:6]};
assign col_out_20 = {u_ca_out_20[5:0], u_ca_out_19[11:6]};
assign col_out_21 = {u_ca_out_21[5:0], u_ca_out_20[11:6]};
assign col_out_22 = {u_ca_out_22[5:0], u_ca_out_21[11:6]};
assign col_out_23 = {u_ca_out_23[5:0], u_ca_out_22[11:6]};
assign col_out_24 = {u_ca_out_24[5:0], u_ca_out_23[11:6]};
assign col_out_25 = {u_ca_out_25[5:0], u_ca_out_24[11:6]};
assign col_out_26 = {u_ca_out_26[5:0], u_ca_out_25[11:6]};
assign col_out_27 = {u_ca_out_27[5:0], u_ca_out_26[11:6]};
assign col_out_28 = {u_ca_out_28[5:0], u_ca_out_27[11:6]};
assign col_out_29 = {u_ca_out_29[5:0], u_ca_out_28[11:6]};
assign col_out_30 = {u_ca_out_30[5:0], u_ca_out_29[11:6]};
assign col_out_31 = {u_ca_out_31[5:0], u_ca_out_30[11:6]};
assign col_out_32 = {u_ca_out_32[5:0], u_ca_out_31[11:6]};
assign col_out_33 = {u_ca_out_33[5:0], u_ca_out_32[11:6]};
assign col_out_34 = {u_ca_out_34[5:0], u_ca_out_33[11:6]};
assign col_out_35 = {u_ca_out_35[5:0], u_ca_out_34[11:6]};
assign col_out_36 = {u_ca_out_36[5:0], u_ca_out_35[11:6]};
assign col_out_37 = {u_ca_out_37[5:0], u_ca_out_36[11:6]};
assign col_out_38 = {u_ca_out_38[5:0], u_ca_out_37[11:6]};
assign col_out_39 = {u_ca_out_39[5:0], u_ca_out_38[11:6]};
assign col_out_40 = {u_ca_out_40[5:0], u_ca_out_39[11:6]};
assign col_out_41 = {u_ca_out_41[5:0], u_ca_out_40[11:6]};
assign col_out_42 = {u_ca_out_42[5:0], u_ca_out_41[11:6]};
assign col_out_43 = {u_ca_out_43[5:0], u_ca_out_42[11:6]};
assign col_out_44 = {u_ca_out_44[5:0], u_ca_out_43[11:6]};
assign col_out_45 = {u_ca_out_45[5:0], u_ca_out_44[11:6]};
assign col_out_46 = {u_ca_out_46[5:0], u_ca_out_45[11:6]};
assign col_out_47 = {u_ca_out_47[5:0], u_ca_out_46[11:6]};
assign col_out_48 = {u_ca_out_48[5:0], u_ca_out_47[11:6]};
assign col_out_49 = {u_ca_out_49[5:0], u_ca_out_48[11:6]};
assign col_out_50 = {u_ca_out_50[5:0], u_ca_out_49[11:6]};
assign col_out_51 = {u_ca_out_51[5:0], u_ca_out_50[11:6]};
assign col_out_52 = {u_ca_out_52[5:0], u_ca_out_51[11:6]};
assign col_out_53 = {u_ca_out_53[5:0], u_ca_out_52[11:6]};
assign col_out_54 = {u_ca_out_54[5:0], u_ca_out_53[11:6]};
assign col_out_55 = {u_ca_out_55[5:0], u_ca_out_54[11:6]};
assign col_out_56 = {u_ca_out_56[5:0], u_ca_out_55[11:6]};
assign col_out_57 = {u_ca_out_57[5:0], u_ca_out_56[11:6]};
assign col_out_58 = {u_ca_out_58[5:0], u_ca_out_57[11:6]};
assign col_out_59 = {u_ca_out_59[5:0], u_ca_out_58[11:6]};
assign col_out_60 = {u_ca_out_60[5:0], u_ca_out_59[11:6]};
assign col_out_61 = {u_ca_out_61[5:0], u_ca_out_60[11:6]};
assign col_out_62 = {u_ca_out_62[5:0], u_ca_out_61[11:6]};
assign col_out_63 = {u_ca_out_63[5:0], u_ca_out_62[11:6]};
assign col_out_64 = {u_ca_out_64[5:0], u_ca_out_63[11:6]};
assign col_out_65 = {u_ca_out_65[5:0], u_ca_out_64[11:6]};
assign col_out_66 = {u_ca_out_66[5:0], u_ca_out_65[11:6]};
assign col_out_67 = {u_ca_out_67[5:0], u_ca_out_66[11:6]};
assign col_out_68 = {u_ca_out_68[5:0], u_ca_out_67[11:6]};
assign col_out_69 = {u_ca_out_69[5:0], u_ca_out_68[11:6]};
assign col_out_70 = {u_ca_out_70[5:0], u_ca_out_69[11:6]};
assign col_out_71 = {u_ca_out_71[5:0], u_ca_out_70[11:6]};
assign col_out_72 = {u_ca_out_72[5:0], u_ca_out_71[11:6]};
assign col_out_73 = {u_ca_out_73[5:0], u_ca_out_72[11:6]};
assign col_out_74 = {u_ca_out_74[5:0], u_ca_out_73[11:6]};
assign col_out_75 = {u_ca_out_75[5:0], u_ca_out_74[11:6]};
assign col_out_76 = {u_ca_out_76[5:0], u_ca_out_75[11:6]};
assign col_out_77 = {u_ca_out_77[5:0], u_ca_out_76[11:6]};
assign col_out_78 = {u_ca_out_78[5:0], u_ca_out_77[11:6]};
assign col_out_79 = {u_ca_out_79[5:0], u_ca_out_78[11:6]};
assign col_out_80 = {u_ca_out_80[5:0], u_ca_out_79[11:6]};
assign col_out_81 = {u_ca_out_81[5:0], u_ca_out_80[11:6]};
assign col_out_82 = {u_ca_out_82[5:0], u_ca_out_81[11:6]};
assign col_out_83 = {u_ca_out_83[5:0], u_ca_out_82[11:6]};
assign col_out_84 = {u_ca_out_84[5:0], u_ca_out_83[11:6]};
assign col_out_85 = {u_ca_out_85[5:0], u_ca_out_84[11:6]};
assign col_out_86 = {u_ca_out_86[5:0], u_ca_out_85[11:6]};
assign col_out_87 = {u_ca_out_87[5:0], u_ca_out_86[11:6]};
assign col_out_88 = {u_ca_out_88[5:0], u_ca_out_87[11:6]};
assign col_out_89 = {u_ca_out_89[5:0], u_ca_out_88[11:6]};
assign col_out_90 = {u_ca_out_90[5:0], u_ca_out_89[11:6]};
assign col_out_91 = {u_ca_out_91[5:0], u_ca_out_90[11:6]};
assign col_out_92 = {u_ca_out_92[5:0], u_ca_out_91[11:6]};
assign col_out_93 = {u_ca_out_93[5:0], u_ca_out_92[11:6]};
assign col_out_94 = {u_ca_out_94[5:0], u_ca_out_93[11:6]};
assign col_out_95 = {u_ca_out_95[5:0], u_ca_out_94[11:6]};
assign col_out_96 = {u_ca_out_96[5:0], u_ca_out_95[11:6]};
assign col_out_97 = {u_ca_out_97[5:0], u_ca_out_96[11:6]};
assign col_out_98 = {u_ca_out_98[5:0], u_ca_out_97[11:6]};
assign col_out_99 = {u_ca_out_99[5:0], u_ca_out_98[11:6]};
assign col_out_100 = {u_ca_out_100[5:0], u_ca_out_99[11:6]};
assign col_out_101 = {u_ca_out_101[5:0], u_ca_out_100[11:6]};
assign col_out_102 = {u_ca_out_102[5:0], u_ca_out_101[11:6]};
assign col_out_103 = {u_ca_out_103[5:0], u_ca_out_102[11:6]};
assign col_out_104 = {u_ca_out_104[5:0], u_ca_out_103[11:6]};
assign col_out_105 = {u_ca_out_105[5:0], u_ca_out_104[11:6]};
assign col_out_106 = {u_ca_out_106[5:0], u_ca_out_105[11:6]};
assign col_out_107 = {u_ca_out_107[5:0], u_ca_out_106[11:6]};
assign col_out_108 = {u_ca_out_108[5:0], u_ca_out_107[11:6]};
assign col_out_109 = {u_ca_out_109[5:0], u_ca_out_108[11:6]};
assign col_out_110 = {u_ca_out_110[5:0], u_ca_out_109[11:6]};
assign col_out_111 = {u_ca_out_111[5:0], u_ca_out_110[11:6]};
assign col_out_112 = {u_ca_out_112[5:0], u_ca_out_111[11:6]};
assign col_out_113 = {u_ca_out_113[5:0], u_ca_out_112[11:6]};
assign col_out_114 = {u_ca_out_114[5:0], u_ca_out_113[11:6]};
assign col_out_115 = {u_ca_out_115[5:0], u_ca_out_114[11:6]};
assign col_out_116 = {u_ca_out_116[5:0], u_ca_out_115[11:6]};
assign col_out_117 = {u_ca_out_117[5:0], u_ca_out_116[11:6]};
assign col_out_118 = {u_ca_out_118[5:0], u_ca_out_117[11:6]};
assign col_out_119 = {u_ca_out_119[5:0], u_ca_out_118[11:6]};
assign col_out_120 = {u_ca_out_120[5:0], u_ca_out_119[11:6]};
assign col_out_121 = {u_ca_out_121[5:0], u_ca_out_120[11:6]};
assign col_out_122 = {u_ca_out_122[5:0], u_ca_out_121[11:6]};
assign col_out_123 = {u_ca_out_123[5:0], u_ca_out_122[11:6]};
assign col_out_124 = {u_ca_out_124[5:0], u_ca_out_123[11:6]};
assign col_out_125 = {u_ca_out_125[5:0], u_ca_out_124[11:6]};
assign col_out_126 = {u_ca_out_126[5:0], u_ca_out_125[11:6]};
assign col_out_127 = {u_ca_out_127[5:0], u_ca_out_126[11:6]};
assign col_out_128 = {u_ca_out_128[5:0], u_ca_out_127[11:6]};
assign col_out_129 = {u_ca_out_129[5:0], u_ca_out_128[11:6]};
assign col_out_130 = {u_ca_out_130[5:0], u_ca_out_129[11:6]};
assign col_out_131 = {u_ca_out_131[5:0], u_ca_out_130[11:6]};
assign col_out_132 = {u_ca_out_132[5:0], u_ca_out_131[11:6]};
assign col_out_133 = {u_ca_out_133[5:0], u_ca_out_132[11:6]};
assign col_out_134 = {u_ca_out_134[5:0], u_ca_out_133[11:6]};
assign col_out_135 = {u_ca_out_135[5:0], u_ca_out_134[11:6]};
assign col_out_136 = {u_ca_out_136[5:0], u_ca_out_135[11:6]};
assign col_out_137 = {u_ca_out_137[5:0], u_ca_out_136[11:6]};
assign col_out_138 = {u_ca_out_138[5:0], u_ca_out_137[11:6]};
assign col_out_139 = {u_ca_out_139[5:0], u_ca_out_138[11:6]};
assign col_out_140 = {u_ca_out_140[5:0], u_ca_out_139[11:6]};
assign col_out_141 = {u_ca_out_141[5:0], u_ca_out_140[11:6]};
assign col_out_142 = {u_ca_out_142[5:0], u_ca_out_141[11:6]};
assign col_out_143 = {u_ca_out_143[5:0], u_ca_out_142[11:6]};
assign col_out_144 = {u_ca_out_144[5:0], u_ca_out_143[11:6]};
assign col_out_145 = {u_ca_out_145[5:0], u_ca_out_144[11:6]};
assign col_out_146 = {u_ca_out_146[5:0], u_ca_out_145[11:6]};
assign col_out_147 = {u_ca_out_147[5:0], u_ca_out_146[11:6]};
assign col_out_148 = {u_ca_out_148[5:0], u_ca_out_147[11:6]};
assign col_out_149 = {u_ca_out_149[5:0], u_ca_out_148[11:6]};
assign col_out_150 = {u_ca_out_150[5:0], u_ca_out_149[11:6]};
assign col_out_151 = {u_ca_out_151[5:0], u_ca_out_150[11:6]};
assign col_out_152 = {u_ca_out_152[5:0], u_ca_out_151[11:6]};
assign col_out_153 = {u_ca_out_153[5:0], u_ca_out_152[11:6]};
assign col_out_154 = {u_ca_out_154[5:0], u_ca_out_153[11:6]};
assign col_out_155 = {u_ca_out_155[5:0], u_ca_out_154[11:6]};
assign col_out_156 = {u_ca_out_156[5:0], u_ca_out_155[11:6]};
assign col_out_157 = {u_ca_out_157[5:0], u_ca_out_156[11:6]};
assign col_out_158 = {u_ca_out_158[5:0], u_ca_out_157[11:6]};
assign col_out_159 = {u_ca_out_159[5:0], u_ca_out_158[11:6]};
assign col_out_160 = {u_ca_out_160[5:0], u_ca_out_159[11:6]};
assign col_out_161 = {u_ca_out_161[5:0], u_ca_out_160[11:6]};
assign col_out_162 = {u_ca_out_162[5:0], u_ca_out_161[11:6]};
assign col_out_163 = {u_ca_out_163[5:0], u_ca_out_162[11:6]};
assign col_out_164 = {u_ca_out_164[5:0], u_ca_out_163[11:6]};
assign col_out_165 = {u_ca_out_165[5:0], u_ca_out_164[11:6]};
assign col_out_166 = {u_ca_out_166[5:0], u_ca_out_165[11:6]};
assign col_out_167 = {u_ca_out_167[5:0], u_ca_out_166[11:6]};
assign col_out_168 = {u_ca_out_168[5:0], u_ca_out_167[11:6]};
assign col_out_169 = {u_ca_out_169[5:0], u_ca_out_168[11:6]};
assign col_out_170 = {u_ca_out_170[5:0], u_ca_out_169[11:6]};
assign col_out_171 = {u_ca_out_171[5:0], u_ca_out_170[11:6]};
assign col_out_172 = {u_ca_out_172[5:0], u_ca_out_171[11:6]};
assign col_out_173 = {u_ca_out_173[5:0], u_ca_out_172[11:6]};
assign col_out_174 = {u_ca_out_174[5:0], u_ca_out_173[11:6]};
assign col_out_175 = {u_ca_out_175[5:0], u_ca_out_174[11:6]};
assign col_out_176 = {u_ca_out_176[5:0], u_ca_out_175[11:6]};
assign col_out_177 = {u_ca_out_177[5:0], u_ca_out_176[11:6]};
assign col_out_178 = {u_ca_out_178[5:0], u_ca_out_177[11:6]};
assign col_out_179 = {u_ca_out_179[5:0], u_ca_out_178[11:6]};
assign col_out_180 = {u_ca_out_180[5:0], u_ca_out_179[11:6]};
assign col_out_181 = {u_ca_out_181[5:0], u_ca_out_180[11:6]};
assign col_out_182 = {u_ca_out_182[5:0], u_ca_out_181[11:6]};
assign col_out_183 = {u_ca_out_183[5:0], u_ca_out_182[11:6]};
assign col_out_184 = {u_ca_out_184[5:0], u_ca_out_183[11:6]};
assign col_out_185 = {u_ca_out_185[5:0], u_ca_out_184[11:6]};
assign col_out_186 = {u_ca_out_186[5:0], u_ca_out_185[11:6]};
assign col_out_187 = {u_ca_out_187[5:0], u_ca_out_186[11:6]};
assign col_out_188 = {u_ca_out_188[5:0], u_ca_out_187[11:6]};
assign col_out_189 = {u_ca_out_189[5:0], u_ca_out_188[11:6]};
assign col_out_190 = {u_ca_out_190[5:0], u_ca_out_189[11:6]};
assign col_out_191 = {u_ca_out_191[5:0], u_ca_out_190[11:6]};
assign col_out_192 = {u_ca_out_192[5:0], u_ca_out_191[11:6]};
assign col_out_193 = {u_ca_out_193[5:0], u_ca_out_192[11:6]};
assign col_out_194 = {u_ca_out_194[5:0], u_ca_out_193[11:6]};
assign col_out_195 = {u_ca_out_195[5:0], u_ca_out_194[11:6]};
assign col_out_196 = {u_ca_out_196[5:0], u_ca_out_195[11:6]};
assign col_out_197 = {u_ca_out_197[5:0], u_ca_out_196[11:6]};
assign col_out_198 = {u_ca_out_198[5:0], u_ca_out_197[11:6]};
assign col_out_199 = {u_ca_out_199[5:0], u_ca_out_198[11:6]};
assign col_out_200 = {u_ca_out_200[5:0], u_ca_out_199[11:6]};
assign col_out_201 = {u_ca_out_201[5:0], u_ca_out_200[11:6]};
assign col_out_202 = {u_ca_out_202[5:0], u_ca_out_201[11:6]};
assign col_out_203 = {u_ca_out_203[5:0], u_ca_out_202[11:6]};
assign col_out_204 = {u_ca_out_204[5:0], u_ca_out_203[11:6]};
assign col_out_205 = {u_ca_out_205[5:0], u_ca_out_204[11:6]};
assign col_out_206 = {u_ca_out_206[5:0], u_ca_out_205[11:6]};
assign col_out_207 = {u_ca_out_207[5:0], u_ca_out_206[11:6]};
assign col_out_208 = {u_ca_out_208[5:0], u_ca_out_207[11:6]};
assign col_out_209 = {u_ca_out_209[5:0], u_ca_out_208[11:6]};
assign col_out_210 = {u_ca_out_210[5:0], u_ca_out_209[11:6]};
assign col_out_211 = {u_ca_out_211[5:0], u_ca_out_210[11:6]};
assign col_out_212 = {u_ca_out_212[5:0], u_ca_out_211[11:6]};
assign col_out_213 = {u_ca_out_213[5:0], u_ca_out_212[11:6]};
assign col_out_214 = {u_ca_out_214[5:0], u_ca_out_213[11:6]};
assign col_out_215 = {u_ca_out_215[5:0], u_ca_out_214[11:6]};
assign col_out_216 = {u_ca_out_216[5:0], u_ca_out_215[11:6]};
assign col_out_217 = {u_ca_out_217[5:0], u_ca_out_216[11:6]};
assign col_out_218 = {u_ca_out_218[5:0], u_ca_out_217[11:6]};
assign col_out_219 = {u_ca_out_219[5:0], u_ca_out_218[11:6]};
assign col_out_220 = {u_ca_out_220[5:0], u_ca_out_219[11:6]};
assign col_out_221 = {u_ca_out_221[5:0], u_ca_out_220[11:6]};
assign col_out_222 = {u_ca_out_222[5:0], u_ca_out_221[11:6]};
assign col_out_223 = {u_ca_out_223[5:0], u_ca_out_222[11:6]};
assign col_out_224 = {u_ca_out_224[5:0], u_ca_out_223[11:6]};
assign col_out_225 = {u_ca_out_225[5:0], u_ca_out_224[11:6]};
assign col_out_226 = {u_ca_out_226[5:0], u_ca_out_225[11:6]};
assign col_out_227 = {u_ca_out_227[5:0], u_ca_out_226[11:6]};
assign col_out_228 = {u_ca_out_228[5:0], u_ca_out_227[11:6]};
assign col_out_229 = {u_ca_out_229[5:0], u_ca_out_228[11:6]};
assign col_out_230 = {u_ca_out_230[5:0], u_ca_out_229[11:6]};
assign col_out_231 = {u_ca_out_231[5:0], u_ca_out_230[11:6]};
assign col_out_232 = {u_ca_out_232[5:0], u_ca_out_231[11:6]};
assign col_out_233 = {u_ca_out_233[5:0], u_ca_out_232[11:6]};
assign col_out_234 = {u_ca_out_234[5:0], u_ca_out_233[11:6]};
assign col_out_235 = {u_ca_out_235[5:0], u_ca_out_234[11:6]};
assign col_out_236 = {u_ca_out_236[5:0], u_ca_out_235[11:6]};
assign col_out_237 = {u_ca_out_237[5:0], u_ca_out_236[11:6]};
assign col_out_238 = {u_ca_out_238[5:0], u_ca_out_237[11:6]};
assign col_out_239 = {u_ca_out_239[5:0], u_ca_out_238[11:6]};
assign col_out_240 = {u_ca_out_240[5:0], u_ca_out_239[11:6]};
assign col_out_241 = {u_ca_out_241[5:0], u_ca_out_240[11:6]};
assign col_out_242 = {u_ca_out_242[5:0], u_ca_out_241[11:6]};
assign col_out_243 = {u_ca_out_243[5:0], u_ca_out_242[11:6]};
assign col_out_244 = {u_ca_out_244[5:0], u_ca_out_243[11:6]};
assign col_out_245 = {u_ca_out_245[5:0], u_ca_out_244[11:6]};
assign col_out_246 = {u_ca_out_246[5:0], u_ca_out_245[11:6]};
assign col_out_247 = {u_ca_out_247[5:0], u_ca_out_246[11:6]};
assign col_out_248 = {u_ca_out_248[5:0], u_ca_out_247[11:6]};
assign col_out_249 = {u_ca_out_249[5:0], u_ca_out_248[11:6]};
assign col_out_250 = {u_ca_out_250[5:0], u_ca_out_249[11:6]};
assign col_out_251 = {u_ca_out_251[5:0], u_ca_out_250[11:6]};
assign col_out_252 = {u_ca_out_252[5:0], u_ca_out_251[11:6]};
assign col_out_253 = {u_ca_out_253[5:0], u_ca_out_252[11:6]};
assign col_out_254 = {u_ca_out_254[5:0], u_ca_out_253[11:6]};
assign col_out_255 = {u_ca_out_255[5:0], u_ca_out_254[11:6]};
assign col_out_256 = {u_ca_out_256[5:0], u_ca_out_255[11:6]};
assign col_out_257 = {u_ca_out_257[5:0], u_ca_out_256[11:6]};
assign col_out_258 = {u_ca_out_258[5:0], u_ca_out_257[11:6]};
assign col_out_259 = {u_ca_out_259[5:0], u_ca_out_258[11:6]};
assign col_out_260 = {u_ca_out_260[5:0], u_ca_out_259[11:6]};
assign col_out_261 = {u_ca_out_261[5:0], u_ca_out_260[11:6]};
assign col_out_262 = {u_ca_out_262[5:0], u_ca_out_261[11:6]};
assign col_out_263 = {u_ca_out_263[5:0], u_ca_out_262[11:6]};
assign col_out_264 = {u_ca_out_264[5:0], u_ca_out_263[11:6]};
assign col_out_265 = {u_ca_out_265[5:0], u_ca_out_264[11:6]};
assign col_out_266 = {u_ca_out_266[5:0], u_ca_out_265[11:6]};
assign col_out_267 = {u_ca_out_267[5:0], u_ca_out_266[11:6]};
assign col_out_268 = {u_ca_out_268[5:0], u_ca_out_267[11:6]};
assign col_out_269 = {u_ca_out_269[5:0], u_ca_out_268[11:6]};
assign col_out_270 = {u_ca_out_270[5:0], u_ca_out_269[11:6]};
assign col_out_271 = {u_ca_out_271[5:0], u_ca_out_270[11:6]};
assign col_out_272 = {u_ca_out_272[5:0], u_ca_out_271[11:6]};
assign col_out_273 = {u_ca_out_273[5:0], u_ca_out_272[11:6]};
assign col_out_274 = {u_ca_out_274[5:0], u_ca_out_273[11:6]};
assign col_out_275 = {u_ca_out_275[5:0], u_ca_out_274[11:6]};
assign col_out_276 = {u_ca_out_276[5:0], u_ca_out_275[11:6]};
assign col_out_277 = {u_ca_out_277[5:0], u_ca_out_276[11:6]};
assign col_out_278 = {u_ca_out_278[5:0], u_ca_out_277[11:6]};
assign col_out_279 = {u_ca_out_279[5:0], u_ca_out_278[11:6]};
assign col_out_280 = {u_ca_out_280[5:0], u_ca_out_279[11:6]};
assign col_out_281 = {u_ca_out_281[5:0], u_ca_out_280[11:6]};
assign col_out_282 = {u_ca_out_282[5:0], u_ca_out_281[11:6]};
assign col_out_283 = {u_ca_out_283[5:0], u_ca_out_282[11:6]};
assign col_out_284 = {u_ca_out_284[5:0], u_ca_out_283[11:6]};
assign col_out_285 = {u_ca_out_285[5:0], u_ca_out_284[11:6]};
assign col_out_286 = {u_ca_out_286[5:0], u_ca_out_285[11:6]};
assign col_out_287 = {u_ca_out_287[5:0], u_ca_out_286[11:6]};
assign col_out_288 = {u_ca_out_288[5:0], u_ca_out_287[11:6]};
assign col_out_289 = {u_ca_out_289[5:0], u_ca_out_288[11:6]};
assign col_out_290 = {u_ca_out_290[5:0], u_ca_out_289[11:6]};
assign col_out_291 = {u_ca_out_291[5:0], u_ca_out_290[11:6]};
assign col_out_292 = {u_ca_out_292[5:0], u_ca_out_291[11:6]};
assign col_out_293 = {u_ca_out_293[5:0], u_ca_out_292[11:6]};
assign col_out_294 = {u_ca_out_294[5:0], u_ca_out_293[11:6]};
assign col_out_295 = {u_ca_out_295[5:0], u_ca_out_294[11:6]};
assign col_out_296 = {u_ca_out_296[5:0], u_ca_out_295[11:6]};
assign col_out_297 = {u_ca_out_297[5:0], u_ca_out_296[11:6]};
assign col_out_298 = {u_ca_out_298[5:0], u_ca_out_297[11:6]};
assign col_out_299 = {u_ca_out_299[5:0], u_ca_out_298[11:6]};
assign col_out_300 = {u_ca_out_300[5:0], u_ca_out_299[11:6]};
assign col_out_301 = {u_ca_out_301[5:0], u_ca_out_300[11:6]};
assign col_out_302 = {u_ca_out_302[5:0], u_ca_out_301[11:6]};
assign col_out_303 = {u_ca_out_303[5:0], u_ca_out_302[11:6]};
assign col_out_304 = {u_ca_out_304[5:0], u_ca_out_303[11:6]};
assign col_out_305 = {u_ca_out_305[5:0], u_ca_out_304[11:6]};
assign col_out_306 = {u_ca_out_306[5:0], u_ca_out_305[11:6]};
assign col_out_307 = {u_ca_out_307[5:0], u_ca_out_306[11:6]};
assign col_out_308 = {u_ca_out_308[5:0], u_ca_out_307[11:6]};
assign col_out_309 = {u_ca_out_309[5:0], u_ca_out_308[11:6]};
assign col_out_310 = {u_ca_out_310[5:0], u_ca_out_309[11:6]};
assign col_out_311 = {u_ca_out_311[5:0], u_ca_out_310[11:6]};
assign col_out_312 = {u_ca_out_312[5:0], u_ca_out_311[11:6]};
assign col_out_313 = {u_ca_out_313[5:0], u_ca_out_312[11:6]};
assign col_out_314 = {u_ca_out_314[5:0], u_ca_out_313[11:6]};
assign col_out_315 = {u_ca_out_315[5:0], u_ca_out_314[11:6]};
assign col_out_316 = {u_ca_out_316[5:0], u_ca_out_315[11:6]};
assign col_out_317 = {u_ca_out_317[5:0], u_ca_out_316[11:6]};
assign col_out_318 = {u_ca_out_318[5:0], u_ca_out_317[11:6]};
assign col_out_319 = {u_ca_out_319[5:0], u_ca_out_318[11:6]};
assign col_out_320 = {u_ca_out_320[5:0], u_ca_out_319[11:6]};
assign col_out_321 = {u_ca_out_321[5:0], u_ca_out_320[11:6]};
assign col_out_322 = {u_ca_out_322[5:0], u_ca_out_321[11:6]};
assign col_out_323 = {u_ca_out_323[5:0], u_ca_out_322[11:6]};
assign col_out_324 = {u_ca_out_324[5:0], u_ca_out_323[11:6]};
assign col_out_325 = {u_ca_out_325[5:0], u_ca_out_324[11:6]};
assign col_out_326 = {u_ca_out_326[5:0], u_ca_out_325[11:6]};
assign col_out_327 = {u_ca_out_327[5:0], u_ca_out_326[11:6]};
assign col_out_328 = {u_ca_out_328[5:0], u_ca_out_327[11:6]};
assign col_out_329 = {u_ca_out_329[5:0], u_ca_out_328[11:6]};
assign col_out_330 = {u_ca_out_330[5:0], u_ca_out_329[11:6]};
assign col_out_331 = {u_ca_out_331[5:0], u_ca_out_330[11:6]};
assign col_out_332 = {u_ca_out_332[5:0], u_ca_out_331[11:6]};
assign col_out_333 = {u_ca_out_333[5:0], u_ca_out_332[11:6]};
assign col_out_334 = {u_ca_out_334[5:0], u_ca_out_333[11:6]};
assign col_out_335 = {u_ca_out_335[5:0], u_ca_out_334[11:6]};
assign col_out_336 = {u_ca_out_336[5:0], u_ca_out_335[11:6]};
assign col_out_337 = {u_ca_out_337[5:0], u_ca_out_336[11:6]};
assign col_out_338 = {u_ca_out_338[5:0], u_ca_out_337[11:6]};
assign col_out_339 = {u_ca_out_339[5:0], u_ca_out_338[11:6]};
assign col_out_340 = {u_ca_out_340[5:0], u_ca_out_339[11:6]};
assign col_out_341 = {u_ca_out_341[5:0], u_ca_out_340[11:6]};
assign col_out_342 = {u_ca_out_342[5:0], u_ca_out_341[11:6]};
assign col_out_343 = {u_ca_out_343[5:0], u_ca_out_342[11:6]};
assign col_out_344 = {u_ca_out_344[5:0], u_ca_out_343[11:6]};
assign col_out_345 = {u_ca_out_345[5:0], u_ca_out_344[11:6]};
assign col_out_346 = {u_ca_out_346[5:0], u_ca_out_345[11:6]};
assign col_out_347 = {u_ca_out_347[5:0], u_ca_out_346[11:6]};
assign col_out_348 = {u_ca_out_348[5:0], u_ca_out_347[11:6]};
assign col_out_349 = {u_ca_out_349[5:0], u_ca_out_348[11:6]};
assign col_out_350 = {u_ca_out_350[5:0], u_ca_out_349[11:6]};
assign col_out_351 = {u_ca_out_351[5:0], u_ca_out_350[11:6]};
assign col_out_352 = {u_ca_out_352[5:0], u_ca_out_351[11:6]};
assign col_out_353 = {u_ca_out_353[5:0], u_ca_out_352[11:6]};
assign col_out_354 = {u_ca_out_354[5:0], u_ca_out_353[11:6]};
assign col_out_355 = {u_ca_out_355[5:0], u_ca_out_354[11:6]};
assign col_out_356 = {u_ca_out_356[5:0], u_ca_out_355[11:6]};
assign col_out_357 = {u_ca_out_357[5:0], u_ca_out_356[11:6]};
assign col_out_358 = {u_ca_out_358[5:0], u_ca_out_357[11:6]};
assign col_out_359 = {u_ca_out_359[5:0], u_ca_out_358[11:6]};
assign col_out_360 = {u_ca_out_360[5:0], u_ca_out_359[11:6]};
assign col_out_361 = {u_ca_out_361[5:0], u_ca_out_360[11:6]};
assign col_out_362 = {u_ca_out_362[5:0], u_ca_out_361[11:6]};
assign col_out_363 = {u_ca_out_363[5:0], u_ca_out_362[11:6]};
assign col_out_364 = {u_ca_out_364[5:0], u_ca_out_363[11:6]};
assign col_out_365 = {u_ca_out_365[5:0], u_ca_out_364[11:6]};
assign col_out_366 = {u_ca_out_366[5:0], u_ca_out_365[11:6]};
assign col_out_367 = {u_ca_out_367[5:0], u_ca_out_366[11:6]};
assign col_out_368 = {u_ca_out_368[5:0], u_ca_out_367[11:6]};
assign col_out_369 = {u_ca_out_369[5:0], u_ca_out_368[11:6]};
assign col_out_370 = {u_ca_out_370[5:0], u_ca_out_369[11:6]};
assign col_out_371 = {u_ca_out_371[5:0], u_ca_out_370[11:6]};
assign col_out_372 = {u_ca_out_372[5:0], u_ca_out_371[11:6]};
assign col_out_373 = {u_ca_out_373[5:0], u_ca_out_372[11:6]};
assign col_out_374 = {u_ca_out_374[5:0], u_ca_out_373[11:6]};
assign col_out_375 = {u_ca_out_375[5:0], u_ca_out_374[11:6]};
assign col_out_376 = {u_ca_out_376[5:0], u_ca_out_375[11:6]};
assign col_out_377 = {u_ca_out_377[5:0], u_ca_out_376[11:6]};
assign col_out_378 = {u_ca_out_378[5:0], u_ca_out_377[11:6]};
assign col_out_379 = {u_ca_out_379[5:0], u_ca_out_378[11:6]};
assign col_out_380 = {u_ca_out_380[5:0], u_ca_out_379[11:6]};
assign col_out_381 = {u_ca_out_381[5:0], u_ca_out_380[11:6]};
assign col_out_382 = {u_ca_out_382[5:0], u_ca_out_381[11:6]};
assign col_out_383 = {u_ca_out_383[5:0], u_ca_out_382[11:6]};
assign col_out_384 = {u_ca_out_384[5:0], u_ca_out_383[11:6]};
assign col_out_385 = {u_ca_out_385[5:0], u_ca_out_384[11:6]};
assign col_out_386 = {u_ca_out_386[5:0], u_ca_out_385[11:6]};
assign col_out_387 = {u_ca_out_387[5:0], u_ca_out_386[11:6]};
assign col_out_388 = {u_ca_out_388[5:0], u_ca_out_387[11:6]};
assign col_out_389 = {u_ca_out_389[5:0], u_ca_out_388[11:6]};
assign col_out_390 = {u_ca_out_390[5:0], u_ca_out_389[11:6]};
assign col_out_391 = {u_ca_out_391[5:0], u_ca_out_390[11:6]};
assign col_out_392 = {u_ca_out_392[5:0], u_ca_out_391[11:6]};
assign col_out_393 = {u_ca_out_393[5:0], u_ca_out_392[11:6]};
assign col_out_394 = {u_ca_out_394[5:0], u_ca_out_393[11:6]};
assign col_out_395 = {u_ca_out_395[5:0], u_ca_out_394[11:6]};
assign col_out_396 = {u_ca_out_396[5:0], u_ca_out_395[11:6]};
assign col_out_397 = {u_ca_out_397[5:0], u_ca_out_396[11:6]};
assign col_out_398 = {u_ca_out_398[5:0], u_ca_out_397[11:6]};
assign col_out_399 = {u_ca_out_399[5:0], u_ca_out_398[11:6]};
assign col_out_400 = {u_ca_out_400[5:0], u_ca_out_399[11:6]};
assign col_out_401 = {u_ca_out_401[5:0], u_ca_out_400[11:6]};
assign col_out_402 = {u_ca_out_402[5:0], u_ca_out_401[11:6]};
assign col_out_403 = {u_ca_out_403[5:0], u_ca_out_402[11:6]};
assign col_out_404 = {u_ca_out_404[5:0], u_ca_out_403[11:6]};
assign col_out_405 = {u_ca_out_405[5:0], u_ca_out_404[11:6]};
assign col_out_406 = {u_ca_out_406[5:0], u_ca_out_405[11:6]};
assign col_out_407 = {u_ca_out_407[5:0], u_ca_out_406[11:6]};
assign col_out_408 = {u_ca_out_408[5:0], u_ca_out_407[11:6]};
assign col_out_409 = {u_ca_out_409[5:0], u_ca_out_408[11:6]};
assign col_out_410 = {u_ca_out_410[5:0], u_ca_out_409[11:6]};
assign col_out_411 = {u_ca_out_411[5:0], u_ca_out_410[11:6]};
assign col_out_412 = {u_ca_out_412[5:0], u_ca_out_411[11:6]};
assign col_out_413 = {u_ca_out_413[5:0], u_ca_out_412[11:6]};
assign col_out_414 = {u_ca_out_414[5:0], u_ca_out_413[11:6]};
assign col_out_415 = {u_ca_out_415[5:0], u_ca_out_414[11:6]};
assign col_out_416 = {u_ca_out_416[5:0], u_ca_out_415[11:6]};
assign col_out_417 = {u_ca_out_417[5:0], u_ca_out_416[11:6]};
assign col_out_418 = {u_ca_out_418[5:0], u_ca_out_417[11:6]};
assign col_out_419 = {u_ca_out_419[5:0], u_ca_out_418[11:6]};
assign col_out_420 = {u_ca_out_420[5:0], u_ca_out_419[11:6]};
assign col_out_421 = {u_ca_out_421[5:0], u_ca_out_420[11:6]};
assign col_out_422 = {u_ca_out_422[5:0], u_ca_out_421[11:6]};
assign col_out_423 = {u_ca_out_423[5:0], u_ca_out_422[11:6]};
assign col_out_424 = {u_ca_out_424[5:0], u_ca_out_423[11:6]};
assign col_out_425 = {u_ca_out_425[5:0], u_ca_out_424[11:6]};
assign col_out_426 = {u_ca_out_426[5:0], u_ca_out_425[11:6]};
assign col_out_427 = {u_ca_out_427[5:0], u_ca_out_426[11:6]};
assign col_out_428 = {u_ca_out_428[5:0], u_ca_out_427[11:6]};
assign col_out_429 = {u_ca_out_429[5:0], u_ca_out_428[11:6]};
assign col_out_430 = {u_ca_out_430[5:0], u_ca_out_429[11:6]};
assign col_out_431 = {u_ca_out_431[5:0], u_ca_out_430[11:6]};
assign col_out_432 = {u_ca_out_432[5:0], u_ca_out_431[11:6]};
assign col_out_433 = {u_ca_out_433[5:0], u_ca_out_432[11:6]};
assign col_out_434 = {u_ca_out_434[5:0], u_ca_out_433[11:6]};
assign col_out_435 = {u_ca_out_435[5:0], u_ca_out_434[11:6]};
assign col_out_436 = {u_ca_out_436[5:0], u_ca_out_435[11:6]};
assign col_out_437 = {u_ca_out_437[5:0], u_ca_out_436[11:6]};
assign col_out_438 = {u_ca_out_438[5:0], u_ca_out_437[11:6]};
assign col_out_439 = {u_ca_out_439[5:0], u_ca_out_438[11:6]};
assign col_out_440 = {u_ca_out_440[5:0], u_ca_out_439[11:6]};
assign col_out_441 = {u_ca_out_441[5:0], u_ca_out_440[11:6]};
assign col_out_442 = {u_ca_out_442[5:0], u_ca_out_441[11:6]};
assign col_out_443 = {u_ca_out_443[5:0], u_ca_out_442[11:6]};
assign col_out_444 = {u_ca_out_444[5:0], u_ca_out_443[11:6]};
assign col_out_445 = {u_ca_out_445[5:0], u_ca_out_444[11:6]};
assign col_out_446 = {u_ca_out_446[5:0], u_ca_out_445[11:6]};
assign col_out_447 = {u_ca_out_447[5:0], u_ca_out_446[11:6]};
assign col_out_448 = {u_ca_out_448[5:0], u_ca_out_447[11:6]};
assign col_out_449 = {u_ca_out_449[5:0], u_ca_out_448[11:6]};
assign col_out_450 = {u_ca_out_450[5:0], u_ca_out_449[11:6]};
assign col_out_451 = {u_ca_out_451[5:0], u_ca_out_450[11:6]};
assign col_out_452 = {u_ca_out_452[5:0], u_ca_out_451[11:6]};
assign col_out_453 = {u_ca_out_453[5:0], u_ca_out_452[11:6]};
assign col_out_454 = {u_ca_out_454[5:0], u_ca_out_453[11:6]};
assign col_out_455 = {u_ca_out_455[5:0], u_ca_out_454[11:6]};
assign col_out_456 = {u_ca_out_456[5:0], u_ca_out_455[11:6]};
assign col_out_457 = {u_ca_out_457[5:0], u_ca_out_456[11:6]};
assign col_out_458 = {u_ca_out_458[5:0], u_ca_out_457[11:6]};
assign col_out_459 = {u_ca_out_459[5:0], u_ca_out_458[11:6]};
assign col_out_460 = {u_ca_out_460[5:0], u_ca_out_459[11:6]};
assign col_out_461 = {u_ca_out_461[5:0], u_ca_out_460[11:6]};
assign col_out_462 = {u_ca_out_462[5:0], u_ca_out_461[11:6]};
assign col_out_463 = {u_ca_out_463[5:0], u_ca_out_462[11:6]};
assign col_out_464 = {u_ca_out_464[5:0], u_ca_out_463[11:6]};
assign col_out_465 = {u_ca_out_465[5:0], u_ca_out_464[11:6]};
assign col_out_466 = {u_ca_out_466[5:0], u_ca_out_465[11:6]};
assign col_out_467 = {u_ca_out_467[5:0], u_ca_out_466[11:6]};
assign col_out_468 = {u_ca_out_468[5:0], u_ca_out_467[11:6]};
assign col_out_469 = {u_ca_out_469[5:0], u_ca_out_468[11:6]};
assign col_out_470 = {u_ca_out_470[5:0], u_ca_out_469[11:6]};
assign col_out_471 = {u_ca_out_471[5:0], u_ca_out_470[11:6]};
assign col_out_472 = {u_ca_out_472[5:0], u_ca_out_471[11:6]};
assign col_out_473 = {u_ca_out_473[5:0], u_ca_out_472[11:6]};
assign col_out_474 = {u_ca_out_474[5:0], u_ca_out_473[11:6]};
assign col_out_475 = {u_ca_out_475[5:0], u_ca_out_474[11:6]};
assign col_out_476 = {u_ca_out_476[5:0], u_ca_out_475[11:6]};
assign col_out_477 = {u_ca_out_477[5:0], u_ca_out_476[11:6]};
assign col_out_478 = {u_ca_out_478[5:0], u_ca_out_477[11:6]};
assign col_out_479 = {u_ca_out_479[5:0], u_ca_out_478[11:6]};
assign col_out_480 = {u_ca_out_480[5:0], u_ca_out_479[11:6]};
assign col_out_481 = {u_ca_out_481[5:0], u_ca_out_480[11:6]};
assign col_out_482 = {u_ca_out_482[5:0], u_ca_out_481[11:6]};
assign col_out_483 = {u_ca_out_483[5:0], u_ca_out_482[11:6]};
assign col_out_484 = {u_ca_out_484[5:0], u_ca_out_483[11:6]};
assign col_out_485 = {u_ca_out_485[5:0], u_ca_out_484[11:6]};
assign col_out_486 = {u_ca_out_486[5:0], u_ca_out_485[11:6]};
assign col_out_487 = {u_ca_out_487[5:0], u_ca_out_486[11:6]};
assign col_out_488 = {u_ca_out_488[5:0], u_ca_out_487[11:6]};
assign col_out_489 = {u_ca_out_489[5:0], u_ca_out_488[11:6]};
assign col_out_490 = {u_ca_out_490[5:0], u_ca_out_489[11:6]};
assign col_out_491 = {u_ca_out_491[5:0], u_ca_out_490[11:6]};
assign col_out_492 = {u_ca_out_492[5:0], u_ca_out_491[11:6]};
assign col_out_493 = {u_ca_out_493[5:0], u_ca_out_492[11:6]};
assign col_out_494 = {u_ca_out_494[5:0], u_ca_out_493[11:6]};
assign col_out_495 = {u_ca_out_495[5:0], u_ca_out_494[11:6]};
assign col_out_496 = {u_ca_out_496[5:0], u_ca_out_495[11:6]};
assign col_out_497 = {u_ca_out_497[5:0], u_ca_out_496[11:6]};
assign col_out_498 = {u_ca_out_498[5:0], u_ca_out_497[11:6]};
assign col_out_499 = {u_ca_out_499[5:0], u_ca_out_498[11:6]};
assign col_out_500 = {u_ca_out_500[5:0], u_ca_out_499[11:6]};
assign col_out_501 = {u_ca_out_501[5:0], u_ca_out_500[11:6]};
assign col_out_502 = {u_ca_out_502[5:0], u_ca_out_501[11:6]};
assign col_out_503 = {u_ca_out_503[5:0], u_ca_out_502[11:6]};
assign col_out_504 = {u_ca_out_504[5:0], u_ca_out_503[11:6]};
assign col_out_505 = {u_ca_out_505[5:0], u_ca_out_504[11:6]};
assign col_out_506 = {u_ca_out_506[5:0], u_ca_out_505[11:6]};
assign col_out_507 = {u_ca_out_507[5:0], u_ca_out_506[11:6]};
assign col_out_508 = {u_ca_out_508[5:0], u_ca_out_507[11:6]};
assign col_out_509 = {u_ca_out_509[5:0], u_ca_out_508[11:6]};
assign col_out_510 = {u_ca_out_510[5:0], u_ca_out_509[11:6]};
assign col_out_511 = {u_ca_out_511[5:0], u_ca_out_510[11:6]};
assign col_out_512 = {u_ca_out_512[5:0], u_ca_out_511[11:6]};
assign col_out_513 = {u_ca_out_513[5:0], u_ca_out_512[11:6]};
assign col_out_514 = {u_ca_out_514[5:0], u_ca_out_513[11:6]};
assign col_out_515 = {u_ca_out_515[5:0], u_ca_out_514[11:6]};
assign col_out_516 = {u_ca_out_516[5:0], u_ca_out_515[11:6]};
assign col_out_517 = {u_ca_out_517[5:0], u_ca_out_516[11:6]};
assign col_out_518 = {u_ca_out_518[5:0], u_ca_out_517[11:6]};
assign col_out_519 = {u_ca_out_519[5:0], u_ca_out_518[11:6]};
assign col_out_520 = {u_ca_out_520[5:0], u_ca_out_519[11:6]};
assign col_out_521 = {u_ca_out_521[5:0], u_ca_out_520[11:6]};
assign col_out_522 = {u_ca_out_522[5:0], u_ca_out_521[11:6]};
assign col_out_523 = {u_ca_out_523[5:0], u_ca_out_522[11:6]};
assign col_out_524 = {u_ca_out_524[5:0], u_ca_out_523[11:6]};
assign col_out_525 = {u_ca_out_525[5:0], u_ca_out_524[11:6]};
assign col_out_526 = {u_ca_out_526[5:0], u_ca_out_525[11:6]};
assign col_out_527 = {u_ca_out_527[5:0], u_ca_out_526[11:6]};
assign col_out_528 = {u_ca_out_528[5:0], u_ca_out_527[11:6]};
assign col_out_529 = {u_ca_out_529[5:0], u_ca_out_528[11:6]};
assign col_out_530 = {u_ca_out_530[5:0], u_ca_out_529[11:6]};
assign col_out_531 = {u_ca_out_531[5:0], u_ca_out_530[11:6]};
assign col_out_532 = {u_ca_out_532[5:0], u_ca_out_531[11:6]};
assign col_out_533 = {u_ca_out_533[5:0], u_ca_out_532[11:6]};
assign col_out_534 = {u_ca_out_534[5:0], u_ca_out_533[11:6]};
assign col_out_535 = {u_ca_out_535[5:0], u_ca_out_534[11:6]};
assign col_out_536 = {u_ca_out_536[5:0], u_ca_out_535[11:6]};
assign col_out_537 = {u_ca_out_537[5:0], u_ca_out_536[11:6]};
assign col_out_538 = {u_ca_out_538[5:0], u_ca_out_537[11:6]};
assign col_out_539 = {u_ca_out_539[5:0], u_ca_out_538[11:6]};
assign col_out_540 = {u_ca_out_540[5:0], u_ca_out_539[11:6]};
assign col_out_541 = {u_ca_out_541[5:0], u_ca_out_540[11:6]};
assign col_out_542 = {u_ca_out_542[5:0], u_ca_out_541[11:6]};
assign col_out_543 = {u_ca_out_543[5:0], u_ca_out_542[11:6]};
assign col_out_544 = {u_ca_out_544[5:0], u_ca_out_543[11:6]};
assign col_out_545 = {u_ca_out_545[5:0], u_ca_out_544[11:6]};
assign col_out_546 = {u_ca_out_546[5:0], u_ca_out_545[11:6]};
assign col_out_547 = {u_ca_out_547[5:0], u_ca_out_546[11:6]};
assign col_out_548 = {u_ca_out_548[5:0], u_ca_out_547[11:6]};
assign col_out_549 = {u_ca_out_549[5:0], u_ca_out_548[11:6]};
assign col_out_550 = {u_ca_out_550[5:0], u_ca_out_549[11:6]};
assign col_out_551 = {u_ca_out_551[5:0], u_ca_out_550[11:6]};
assign col_out_552 = {u_ca_out_552[5:0], u_ca_out_551[11:6]};
assign col_out_553 = {u_ca_out_553[5:0], u_ca_out_552[11:6]};
assign col_out_554 = {u_ca_out_554[5:0], u_ca_out_553[11:6]};
assign col_out_555 = {u_ca_out_555[5:0], u_ca_out_554[11:6]};
assign col_out_556 = {u_ca_out_556[5:0], u_ca_out_555[11:6]};
assign col_out_557 = {u_ca_out_557[5:0], u_ca_out_556[11:6]};
assign col_out_558 = {u_ca_out_558[5:0], u_ca_out_557[11:6]};
assign col_out_559 = {u_ca_out_559[5:0], u_ca_out_558[11:6]};
assign col_out_560 = {u_ca_out_560[5:0], u_ca_out_559[11:6]};
assign col_out_561 = {u_ca_out_561[5:0], u_ca_out_560[11:6]};
assign col_out_562 = {u_ca_out_562[5:0], u_ca_out_561[11:6]};
assign col_out_563 = {u_ca_out_563[5:0], u_ca_out_562[11:6]};
assign col_out_564 = {u_ca_out_564[5:0], u_ca_out_563[11:6]};
assign col_out_565 = {u_ca_out_565[5:0], u_ca_out_564[11:6]};
assign col_out_566 = {u_ca_out_566[5:0], u_ca_out_565[11:6]};
assign col_out_567 = {u_ca_out_567[5:0], u_ca_out_566[11:6]};
assign col_out_568 = {u_ca_out_568[5:0], u_ca_out_567[11:6]};
assign col_out_569 = {u_ca_out_569[5:0], u_ca_out_568[11:6]};
assign col_out_570 = {u_ca_out_570[5:0], u_ca_out_569[11:6]};
assign col_out_571 = {u_ca_out_571[5:0], u_ca_out_570[11:6]};
assign col_out_572 = {u_ca_out_572[5:0], u_ca_out_571[11:6]};
assign col_out_573 = {u_ca_out_573[5:0], u_ca_out_572[11:6]};
assign col_out_574 = {u_ca_out_574[5:0], u_ca_out_573[11:6]};
assign col_out_575 = {u_ca_out_575[5:0], u_ca_out_574[11:6]};
assign col_out_576 = {u_ca_out_576[5:0], u_ca_out_575[11:6]};
assign col_out_577 = {u_ca_out_577[5:0], u_ca_out_576[11:6]};
assign col_out_578 = {u_ca_out_578[5:0], u_ca_out_577[11:6]};
assign col_out_579 = {u_ca_out_579[5:0], u_ca_out_578[11:6]};
assign col_out_580 = {u_ca_out_580[5:0], u_ca_out_579[11:6]};
assign col_out_581 = {u_ca_out_581[5:0], u_ca_out_580[11:6]};
assign col_out_582 = {u_ca_out_582[5:0], u_ca_out_581[11:6]};
assign col_out_583 = {u_ca_out_583[5:0], u_ca_out_582[11:6]};
assign col_out_584 = {u_ca_out_584[5:0], u_ca_out_583[11:6]};
assign col_out_585 = {u_ca_out_585[5:0], u_ca_out_584[11:6]};
assign col_out_586 = {u_ca_out_586[5:0], u_ca_out_585[11:6]};
assign col_out_587 = {u_ca_out_587[5:0], u_ca_out_586[11:6]};
assign col_out_588 = {u_ca_out_588[5:0], u_ca_out_587[11:6]};
assign col_out_589 = {u_ca_out_589[5:0], u_ca_out_588[11:6]};
assign col_out_590 = {u_ca_out_590[5:0], u_ca_out_589[11:6]};
assign col_out_591 = {u_ca_out_591[5:0], u_ca_out_590[11:6]};
assign col_out_592 = {u_ca_out_592[5:0], u_ca_out_591[11:6]};
assign col_out_593 = {u_ca_out_593[5:0], u_ca_out_592[11:6]};
assign col_out_594 = {u_ca_out_594[5:0], u_ca_out_593[11:6]};
assign col_out_595 = {u_ca_out_595[5:0], u_ca_out_594[11:6]};
assign col_out_596 = {u_ca_out_596[5:0], u_ca_out_595[11:6]};
assign col_out_597 = {u_ca_out_597[5:0], u_ca_out_596[11:6]};
assign col_out_598 = {u_ca_out_598[5:0], u_ca_out_597[11:6]};
assign col_out_599 = {u_ca_out_599[5:0], u_ca_out_598[11:6]};
assign col_out_600 = {u_ca_out_600[5:0], u_ca_out_599[11:6]};
assign col_out_601 = {u_ca_out_601[5:0], u_ca_out_600[11:6]};
assign col_out_602 = {u_ca_out_602[5:0], u_ca_out_601[11:6]};
assign col_out_603 = {u_ca_out_603[5:0], u_ca_out_602[11:6]};
assign col_out_604 = {u_ca_out_604[5:0], u_ca_out_603[11:6]};
assign col_out_605 = {u_ca_out_605[5:0], u_ca_out_604[11:6]};
assign col_out_606 = {u_ca_out_606[5:0], u_ca_out_605[11:6]};
assign col_out_607 = {u_ca_out_607[5:0], u_ca_out_606[11:6]};
assign col_out_608 = {u_ca_out_608[5:0], u_ca_out_607[11:6]};
assign col_out_609 = {u_ca_out_609[5:0], u_ca_out_608[11:6]};
assign col_out_610 = {u_ca_out_610[5:0], u_ca_out_609[11:6]};
assign col_out_611 = {u_ca_out_611[5:0], u_ca_out_610[11:6]};
assign col_out_612 = {u_ca_out_612[5:0], u_ca_out_611[11:6]};
assign col_out_613 = {u_ca_out_613[5:0], u_ca_out_612[11:6]};
assign col_out_614 = {u_ca_out_614[5:0], u_ca_out_613[11:6]};
assign col_out_615 = {u_ca_out_615[5:0], u_ca_out_614[11:6]};
assign col_out_616 = {u_ca_out_616[5:0], u_ca_out_615[11:6]};
assign col_out_617 = {u_ca_out_617[5:0], u_ca_out_616[11:6]};
assign col_out_618 = {u_ca_out_618[5:0], u_ca_out_617[11:6]};
assign col_out_619 = {u_ca_out_619[5:0], u_ca_out_618[11:6]};
assign col_out_620 = {u_ca_out_620[5:0], u_ca_out_619[11:6]};
assign col_out_621 = {u_ca_out_621[5:0], u_ca_out_620[11:6]};
assign col_out_622 = {u_ca_out_622[5:0], u_ca_out_621[11:6]};
assign col_out_623 = {u_ca_out_623[5:0], u_ca_out_622[11:6]};
assign col_out_624 = {u_ca_out_624[5:0], u_ca_out_623[11:6]};
assign col_out_625 = {u_ca_out_625[5:0], u_ca_out_624[11:6]};
assign col_out_626 = {u_ca_out_626[5:0], u_ca_out_625[11:6]};
assign col_out_627 = {u_ca_out_627[5:0], u_ca_out_626[11:6]};
assign col_out_628 = {u_ca_out_628[5:0], u_ca_out_627[11:6]};
assign col_out_629 = {u_ca_out_629[5:0], u_ca_out_628[11:6]};
assign col_out_630 = {u_ca_out_630[5:0], u_ca_out_629[11:6]};
assign col_out_631 = {u_ca_out_631[5:0], u_ca_out_630[11:6]};
assign col_out_632 = {u_ca_out_632[5:0], u_ca_out_631[11:6]};
assign col_out_633 = {u_ca_out_633[5:0], u_ca_out_632[11:6]};
assign col_out_634 = {u_ca_out_634[5:0], u_ca_out_633[11:6]};
assign col_out_635 = {u_ca_out_635[5:0], u_ca_out_634[11:6]};
assign col_out_636 = {u_ca_out_636[5:0], u_ca_out_635[11:6]};
assign col_out_637 = {u_ca_out_637[5:0], u_ca_out_636[11:6]};
assign col_out_638 = {u_ca_out_638[5:0], u_ca_out_637[11:6]};
assign col_out_639 = {u_ca_out_639[5:0], u_ca_out_638[11:6]};
assign col_out_640 = {u_ca_out_640[5:0], u_ca_out_639[11:6]};
assign col_out_641 = {u_ca_out_641[5:0], u_ca_out_640[11:6]};
assign col_out_642 = {u_ca_out_642[5:0], u_ca_out_641[11:6]};
assign col_out_643 = {u_ca_out_643[5:0], u_ca_out_642[11:6]};
assign col_out_644 = {u_ca_out_644[5:0], u_ca_out_643[11:6]};
assign col_out_645 = {u_ca_out_645[5:0], u_ca_out_644[11:6]};
assign col_out_646 = {u_ca_out_646[5:0], u_ca_out_645[11:6]};
assign col_out_647 = {u_ca_out_647[5:0], u_ca_out_646[11:6]};
assign col_out_648 = {u_ca_out_648[5:0], u_ca_out_647[11:6]};
assign col_out_649 = {u_ca_out_649[5:0], u_ca_out_648[11:6]};
assign col_out_650 = {u_ca_out_650[5:0], u_ca_out_649[11:6]};
assign col_out_651 = {u_ca_out_651[5:0], u_ca_out_650[11:6]};
assign col_out_652 = {u_ca_out_652[5:0], u_ca_out_651[11:6]};
assign col_out_653 = {u_ca_out_653[5:0], u_ca_out_652[11:6]};
assign col_out_654 = {u_ca_out_654[5:0], u_ca_out_653[11:6]};
assign col_out_655 = {u_ca_out_655[5:0], u_ca_out_654[11:6]};
assign col_out_656 = {u_ca_out_656[5:0], u_ca_out_655[11:6]};
assign col_out_657 = {u_ca_out_657[5:0], u_ca_out_656[11:6]};
assign col_out_658 = {u_ca_out_658[5:0], u_ca_out_657[11:6]};
assign col_out_659 = {u_ca_out_659[5:0], u_ca_out_658[11:6]};
assign col_out_660 = {u_ca_out_660[5:0], u_ca_out_659[11:6]};
assign col_out_661 = {u_ca_out_661[5:0], u_ca_out_660[11:6]};
assign col_out_662 = {u_ca_out_662[5:0], u_ca_out_661[11:6]};
assign col_out_663 = {u_ca_out_663[5:0], u_ca_out_662[11:6]};
assign col_out_664 = {u_ca_out_664[5:0], u_ca_out_663[11:6]};
assign col_out_665 = {u_ca_out_665[5:0], u_ca_out_664[11:6]};
assign col_out_666 = {u_ca_out_666[5:0], u_ca_out_665[11:6]};
assign col_out_667 = {u_ca_out_667[5:0], u_ca_out_666[11:6]};
assign col_out_668 = {u_ca_out_668[5:0], u_ca_out_667[11:6]};
assign col_out_669 = {u_ca_out_669[5:0], u_ca_out_668[11:6]};
assign col_out_670 = {u_ca_out_670[5:0], u_ca_out_669[11:6]};
assign col_out_671 = {u_ca_out_671[5:0], u_ca_out_670[11:6]};
assign col_out_672 = {u_ca_out_672[5:0], u_ca_out_671[11:6]};
assign col_out_673 = {u_ca_out_673[5:0], u_ca_out_672[11:6]};
assign col_out_674 = {u_ca_out_674[5:0], u_ca_out_673[11:6]};
assign col_out_675 = {u_ca_out_675[5:0], u_ca_out_674[11:6]};
assign col_out_676 = {u_ca_out_676[5:0], u_ca_out_675[11:6]};
assign col_out_677 = {u_ca_out_677[5:0], u_ca_out_676[11:6]};
assign col_out_678 = {u_ca_out_678[5:0], u_ca_out_677[11:6]};
assign col_out_679 = {u_ca_out_679[5:0], u_ca_out_678[11:6]};
assign col_out_680 = {u_ca_out_680[5:0], u_ca_out_679[11:6]};
assign col_out_681 = {u_ca_out_681[5:0], u_ca_out_680[11:6]};
assign col_out_682 = {u_ca_out_682[5:0], u_ca_out_681[11:6]};
assign col_out_683 = {u_ca_out_683[5:0], u_ca_out_682[11:6]};
assign col_out_684 = {u_ca_out_684[5:0], u_ca_out_683[11:6]};
assign col_out_685 = {u_ca_out_685[5:0], u_ca_out_684[11:6]};
assign col_out_686 = {u_ca_out_686[5:0], u_ca_out_685[11:6]};
assign col_out_687 = {u_ca_out_687[5:0], u_ca_out_686[11:6]};
assign col_out_688 = {u_ca_out_688[5:0], u_ca_out_687[11:6]};
assign col_out_689 = {u_ca_out_689[5:0], u_ca_out_688[11:6]};
assign col_out_690 = {u_ca_out_690[5:0], u_ca_out_689[11:6]};
assign col_out_691 = {u_ca_out_691[5:0], u_ca_out_690[11:6]};
assign col_out_692 = {u_ca_out_692[5:0], u_ca_out_691[11:6]};
assign col_out_693 = {u_ca_out_693[5:0], u_ca_out_692[11:6]};
assign col_out_694 = {u_ca_out_694[5:0], u_ca_out_693[11:6]};
assign col_out_695 = {u_ca_out_695[5:0], u_ca_out_694[11:6]};
assign col_out_696 = {u_ca_out_696[5:0], u_ca_out_695[11:6]};
assign col_out_697 = {u_ca_out_697[5:0], u_ca_out_696[11:6]};
assign col_out_698 = {u_ca_out_698[5:0], u_ca_out_697[11:6]};
assign col_out_699 = {u_ca_out_699[5:0], u_ca_out_698[11:6]};
assign col_out_700 = {u_ca_out_700[5:0], u_ca_out_699[11:6]};
assign col_out_701 = {u_ca_out_701[5:0], u_ca_out_700[11:6]};
assign col_out_702 = {u_ca_out_702[5:0], u_ca_out_701[11:6]};
assign col_out_703 = {u_ca_out_703[5:0], u_ca_out_702[11:6]};
assign col_out_704 = {u_ca_out_704[5:0], u_ca_out_703[11:6]};
assign col_out_705 = {u_ca_out_705[5:0], u_ca_out_704[11:6]};
assign col_out_706 = {u_ca_out_706[5:0], u_ca_out_705[11:6]};
assign col_out_707 = {u_ca_out_707[5:0], u_ca_out_706[11:6]};
assign col_out_708 = {u_ca_out_708[5:0], u_ca_out_707[11:6]};
assign col_out_709 = {u_ca_out_709[5:0], u_ca_out_708[11:6]};
assign col_out_710 = {u_ca_out_710[5:0], u_ca_out_709[11:6]};
assign col_out_711 = {u_ca_out_711[5:0], u_ca_out_710[11:6]};
assign col_out_712 = {u_ca_out_712[5:0], u_ca_out_711[11:6]};
assign col_out_713 = {u_ca_out_713[5:0], u_ca_out_712[11:6]};
assign col_out_714 = {u_ca_out_714[5:0], u_ca_out_713[11:6]};
assign col_out_715 = {u_ca_out_715[5:0], u_ca_out_714[11:6]};
assign col_out_716 = {u_ca_out_716[5:0], u_ca_out_715[11:6]};
assign col_out_717 = {u_ca_out_717[5:0], u_ca_out_716[11:6]};
assign col_out_718 = {u_ca_out_718[5:0], u_ca_out_717[11:6]};
assign col_out_719 = {u_ca_out_719[5:0], u_ca_out_718[11:6]};
assign col_out_720 = {u_ca_out_720[5:0], u_ca_out_719[11:6]};
assign col_out_721 = {u_ca_out_721[5:0], u_ca_out_720[11:6]};
assign col_out_722 = {u_ca_out_722[5:0], u_ca_out_721[11:6]};
assign col_out_723 = {u_ca_out_723[5:0], u_ca_out_722[11:6]};
assign col_out_724 = {u_ca_out_724[5:0], u_ca_out_723[11:6]};
assign col_out_725 = {u_ca_out_725[5:0], u_ca_out_724[11:6]};
assign col_out_726 = {u_ca_out_726[5:0], u_ca_out_725[11:6]};
assign col_out_727 = {u_ca_out_727[5:0], u_ca_out_726[11:6]};
assign col_out_728 = {u_ca_out_728[5:0], u_ca_out_727[11:6]};
assign col_out_729 = {u_ca_out_729[5:0], u_ca_out_728[11:6]};
assign col_out_730 = {u_ca_out_730[5:0], u_ca_out_729[11:6]};
assign col_out_731 = {u_ca_out_731[5:0], u_ca_out_730[11:6]};
assign col_out_732 = {u_ca_out_732[5:0], u_ca_out_731[11:6]};
assign col_out_733 = {u_ca_out_733[5:0], u_ca_out_732[11:6]};
assign col_out_734 = {u_ca_out_734[5:0], u_ca_out_733[11:6]};
assign col_out_735 = {u_ca_out_735[5:0], u_ca_out_734[11:6]};
assign col_out_736 = {u_ca_out_736[5:0], u_ca_out_735[11:6]};
assign col_out_737 = {u_ca_out_737[5:0], u_ca_out_736[11:6]};
assign col_out_738 = {u_ca_out_738[5:0], u_ca_out_737[11:6]};
assign col_out_739 = {u_ca_out_739[5:0], u_ca_out_738[11:6]};
assign col_out_740 = {u_ca_out_740[5:0], u_ca_out_739[11:6]};
assign col_out_741 = {u_ca_out_741[5:0], u_ca_out_740[11:6]};
assign col_out_742 = {u_ca_out_742[5:0], u_ca_out_741[11:6]};
assign col_out_743 = {u_ca_out_743[5:0], u_ca_out_742[11:6]};
assign col_out_744 = {u_ca_out_744[5:0], u_ca_out_743[11:6]};
assign col_out_745 = {u_ca_out_745[5:0], u_ca_out_744[11:6]};
assign col_out_746 = {u_ca_out_746[5:0], u_ca_out_745[11:6]};
assign col_out_747 = {u_ca_out_747[5:0], u_ca_out_746[11:6]};
assign col_out_748 = {u_ca_out_748[5:0], u_ca_out_747[11:6]};
assign col_out_749 = {u_ca_out_749[5:0], u_ca_out_748[11:6]};
assign col_out_750 = {u_ca_out_750[5:0], u_ca_out_749[11:6]};
assign col_out_751 = {u_ca_out_751[5:0], u_ca_out_750[11:6]};
assign col_out_752 = {u_ca_out_752[5:0], u_ca_out_751[11:6]};
assign col_out_753 = {u_ca_out_753[5:0], u_ca_out_752[11:6]};
assign col_out_754 = {u_ca_out_754[5:0], u_ca_out_753[11:6]};
assign col_out_755 = {u_ca_out_755[5:0], u_ca_out_754[11:6]};
assign col_out_756 = {u_ca_out_756[5:0], u_ca_out_755[11:6]};
assign col_out_757 = {u_ca_out_757[5:0], u_ca_out_756[11:6]};
assign col_out_758 = {u_ca_out_758[5:0], u_ca_out_757[11:6]};
assign col_out_759 = {u_ca_out_759[5:0], u_ca_out_758[11:6]};
assign col_out_760 = {u_ca_out_760[5:0], u_ca_out_759[11:6]};
assign col_out_761 = {u_ca_out_761[5:0], u_ca_out_760[11:6]};
assign col_out_762 = {u_ca_out_762[5:0], u_ca_out_761[11:6]};
assign col_out_763 = {u_ca_out_763[5:0], u_ca_out_762[11:6]};
assign col_out_764 = {u_ca_out_764[5:0], u_ca_out_763[11:6]};
assign col_out_765 = {u_ca_out_765[5:0], u_ca_out_764[11:6]};
assign col_out_766 = {u_ca_out_766[5:0], u_ca_out_765[11:6]};
assign col_out_767 = {u_ca_out_767[5:0], u_ca_out_766[11:6]};
assign col_out_768 = {u_ca_out_768[5:0], u_ca_out_767[11:6]};
assign col_out_769 = {u_ca_out_769[5:0], u_ca_out_768[11:6]};
assign col_out_770 = {u_ca_out_770[5:0], u_ca_out_769[11:6]};
assign col_out_771 = {u_ca_out_771[5:0], u_ca_out_770[11:6]};
assign col_out_772 = {u_ca_out_772[5:0], u_ca_out_771[11:6]};
assign col_out_773 = {u_ca_out_773[5:0], u_ca_out_772[11:6]};
assign col_out_774 = {u_ca_out_774[5:0], u_ca_out_773[11:6]};
assign col_out_775 = {u_ca_out_775[5:0], u_ca_out_774[11:6]};
assign col_out_776 = {u_ca_out_776[5:0], u_ca_out_775[11:6]};
assign col_out_777 = {u_ca_out_777[5:0], u_ca_out_776[11:6]};
assign col_out_778 = {u_ca_out_778[5:0], u_ca_out_777[11:6]};
assign col_out_779 = {u_ca_out_779[5:0], u_ca_out_778[11:6]};
assign col_out_780 = {u_ca_out_780[5:0], u_ca_out_779[11:6]};
assign col_out_781 = {u_ca_out_781[5:0], u_ca_out_780[11:6]};
assign col_out_782 = {u_ca_out_782[5:0], u_ca_out_781[11:6]};
assign col_out_783 = {u_ca_out_783[5:0], u_ca_out_782[11:6]};
assign col_out_784 = {u_ca_out_784[5:0], u_ca_out_783[11:6]};
assign col_out_785 = {u_ca_out_785[5:0], u_ca_out_784[11:6]};
assign col_out_786 = {u_ca_out_786[5:0], u_ca_out_785[11:6]};
assign col_out_787 = {u_ca_out_787[5:0], u_ca_out_786[11:6]};
assign col_out_788 = {u_ca_out_788[5:0], u_ca_out_787[11:6]};
assign col_out_789 = {u_ca_out_789[5:0], u_ca_out_788[11:6]};
assign col_out_790 = {u_ca_out_790[5:0], u_ca_out_789[11:6]};
assign col_out_791 = {u_ca_out_791[5:0], u_ca_out_790[11:6]};
assign col_out_792 = {u_ca_out_792[5:0], u_ca_out_791[11:6]};
assign col_out_793 = {u_ca_out_793[5:0], u_ca_out_792[11:6]};
assign col_out_794 = {u_ca_out_794[5:0], u_ca_out_793[11:6]};
assign col_out_795 = {u_ca_out_795[5:0], u_ca_out_794[11:6]};
assign col_out_796 = {u_ca_out_796[5:0], u_ca_out_795[11:6]};
assign col_out_797 = {u_ca_out_797[5:0], u_ca_out_796[11:6]};
assign col_out_798 = {u_ca_out_798[5:0], u_ca_out_797[11:6]};
assign col_out_799 = {u_ca_out_799[5:0], u_ca_out_798[11:6]};
assign col_out_800 = {u_ca_out_800[5:0], u_ca_out_799[11:6]};
assign col_out_801 = {u_ca_out_801[5:0], u_ca_out_800[11:6]};
assign col_out_802 = {u_ca_out_802[5:0], u_ca_out_801[11:6]};
assign col_out_803 = {u_ca_out_803[5:0], u_ca_out_802[11:6]};
assign col_out_804 = {u_ca_out_804[5:0], u_ca_out_803[11:6]};
assign col_out_805 = {u_ca_out_805[5:0], u_ca_out_804[11:6]};
assign col_out_806 = {u_ca_out_806[5:0], u_ca_out_805[11:6]};
assign col_out_807 = {u_ca_out_807[5:0], u_ca_out_806[11:6]};
assign col_out_808 = {u_ca_out_808[5:0], u_ca_out_807[11:6]};
assign col_out_809 = {u_ca_out_809[5:0], u_ca_out_808[11:6]};
assign col_out_810 = {u_ca_out_810[5:0], u_ca_out_809[11:6]};
assign col_out_811 = {u_ca_out_811[5:0], u_ca_out_810[11:6]};
assign col_out_812 = {u_ca_out_812[5:0], u_ca_out_811[11:6]};
assign col_out_813 = {u_ca_out_813[5:0], u_ca_out_812[11:6]};
assign col_out_814 = {u_ca_out_814[5:0], u_ca_out_813[11:6]};
assign col_out_815 = {u_ca_out_815[5:0], u_ca_out_814[11:6]};
assign col_out_816 = {u_ca_out_816[5:0], u_ca_out_815[11:6]};
assign col_out_817 = {u_ca_out_817[5:0], u_ca_out_816[11:6]};
assign col_out_818 = {u_ca_out_818[5:0], u_ca_out_817[11:6]};
assign col_out_819 = {u_ca_out_819[5:0], u_ca_out_818[11:6]};
assign col_out_820 = {u_ca_out_820[5:0], u_ca_out_819[11:6]};
assign col_out_821 = {u_ca_out_821[5:0], u_ca_out_820[11:6]};
assign col_out_822 = {u_ca_out_822[5:0], u_ca_out_821[11:6]};
assign col_out_823 = {u_ca_out_823[5:0], u_ca_out_822[11:6]};
assign col_out_824 = {u_ca_out_824[5:0], u_ca_out_823[11:6]};
assign col_out_825 = {u_ca_out_825[5:0], u_ca_out_824[11:6]};
assign col_out_826 = {u_ca_out_826[5:0], u_ca_out_825[11:6]};
assign col_out_827 = {u_ca_out_827[5:0], u_ca_out_826[11:6]};
assign col_out_828 = {u_ca_out_828[5:0], u_ca_out_827[11:6]};
assign col_out_829 = {u_ca_out_829[5:0], u_ca_out_828[11:6]};
assign col_out_830 = {u_ca_out_830[5:0], u_ca_out_829[11:6]};
assign col_out_831 = {u_ca_out_831[5:0], u_ca_out_830[11:6]};
assign col_out_832 = {u_ca_out_832[5:0], u_ca_out_831[11:6]};
assign col_out_833 = {u_ca_out_833[5:0], u_ca_out_832[11:6]};
assign col_out_834 = {u_ca_out_834[5:0], u_ca_out_833[11:6]};
assign col_out_835 = {u_ca_out_835[5:0], u_ca_out_834[11:6]};
assign col_out_836 = {u_ca_out_836[5:0], u_ca_out_835[11:6]};
assign col_out_837 = {u_ca_out_837[5:0], u_ca_out_836[11:6]};
assign col_out_838 = {u_ca_out_838[5:0], u_ca_out_837[11:6]};
assign col_out_839 = {u_ca_out_839[5:0], u_ca_out_838[11:6]};
assign col_out_840 = {u_ca_out_840[5:0], u_ca_out_839[11:6]};
assign col_out_841 = {u_ca_out_841[5:0], u_ca_out_840[11:6]};
assign col_out_842 = {u_ca_out_842[5:0], u_ca_out_841[11:6]};
assign col_out_843 = {u_ca_out_843[5:0], u_ca_out_842[11:6]};
assign col_out_844 = {u_ca_out_844[5:0], u_ca_out_843[11:6]};
assign col_out_845 = {u_ca_out_845[5:0], u_ca_out_844[11:6]};
assign col_out_846 = {u_ca_out_846[5:0], u_ca_out_845[11:6]};
assign col_out_847 = {u_ca_out_847[5:0], u_ca_out_846[11:6]};
assign col_out_848 = {u_ca_out_848[5:0], u_ca_out_847[11:6]};
assign col_out_849 = {u_ca_out_849[5:0], u_ca_out_848[11:6]};
assign col_out_850 = {u_ca_out_850[5:0], u_ca_out_849[11:6]};
assign col_out_851 = {u_ca_out_851[5:0], u_ca_out_850[11:6]};
assign col_out_852 = {u_ca_out_852[5:0], u_ca_out_851[11:6]};
assign col_out_853 = {u_ca_out_853[5:0], u_ca_out_852[11:6]};
assign col_out_854 = {u_ca_out_854[5:0], u_ca_out_853[11:6]};
assign col_out_855 = {u_ca_out_855[5:0], u_ca_out_854[11:6]};
assign col_out_856 = {u_ca_out_856[5:0], u_ca_out_855[11:6]};
assign col_out_857 = {u_ca_out_857[5:0], u_ca_out_856[11:6]};
assign col_out_858 = {u_ca_out_858[5:0], u_ca_out_857[11:6]};
assign col_out_859 = {u_ca_out_859[5:0], u_ca_out_858[11:6]};
assign col_out_860 = {u_ca_out_860[5:0], u_ca_out_859[11:6]};
assign col_out_861 = {u_ca_out_861[5:0], u_ca_out_860[11:6]};
assign col_out_862 = {u_ca_out_862[5:0], u_ca_out_861[11:6]};
assign col_out_863 = {u_ca_out_863[5:0], u_ca_out_862[11:6]};
assign col_out_864 = {u_ca_out_864[5:0], u_ca_out_863[11:6]};
assign col_out_865 = {u_ca_out_865[5:0], u_ca_out_864[11:6]};
assign col_out_866 = {u_ca_out_866[5:0], u_ca_out_865[11:6]};
assign col_out_867 = {u_ca_out_867[5:0], u_ca_out_866[11:6]};
assign col_out_868 = {u_ca_out_868[5:0], u_ca_out_867[11:6]};
assign col_out_869 = {u_ca_out_869[5:0], u_ca_out_868[11:6]};
assign col_out_870 = {u_ca_out_870[5:0], u_ca_out_869[11:6]};
assign col_out_871 = {u_ca_out_871[5:0], u_ca_out_870[11:6]};
assign col_out_872 = {u_ca_out_872[5:0], u_ca_out_871[11:6]};
assign col_out_873 = {u_ca_out_873[5:0], u_ca_out_872[11:6]};
assign col_out_874 = {u_ca_out_874[5:0], u_ca_out_873[11:6]};
assign col_out_875 = {u_ca_out_875[5:0], u_ca_out_874[11:6]};
assign col_out_876 = {u_ca_out_876[5:0], u_ca_out_875[11:6]};
assign col_out_877 = {u_ca_out_877[5:0], u_ca_out_876[11:6]};
assign col_out_878 = {u_ca_out_878[5:0], u_ca_out_877[11:6]};
assign col_out_879 = {u_ca_out_879[5:0], u_ca_out_878[11:6]};
assign col_out_880 = {u_ca_out_880[5:0], u_ca_out_879[11:6]};
assign col_out_881 = {u_ca_out_881[5:0], u_ca_out_880[11:6]};
assign col_out_882 = {u_ca_out_882[5:0], u_ca_out_881[11:6]};
assign col_out_883 = {u_ca_out_883[5:0], u_ca_out_882[11:6]};
assign col_out_884 = {u_ca_out_884[5:0], u_ca_out_883[11:6]};
assign col_out_885 = {u_ca_out_885[5:0], u_ca_out_884[11:6]};
assign col_out_886 = {u_ca_out_886[5:0], u_ca_out_885[11:6]};
assign col_out_887 = {u_ca_out_887[5:0], u_ca_out_886[11:6]};
assign col_out_888 = {u_ca_out_888[5:0], u_ca_out_887[11:6]};
assign col_out_889 = {u_ca_out_889[5:0], u_ca_out_888[11:6]};
assign col_out_890 = {u_ca_out_890[5:0], u_ca_out_889[11:6]};
assign col_out_891 = {u_ca_out_891[5:0], u_ca_out_890[11:6]};
assign col_out_892 = {u_ca_out_892[5:0], u_ca_out_891[11:6]};
assign col_out_893 = {u_ca_out_893[5:0], u_ca_out_892[11:6]};
assign col_out_894 = {u_ca_out_894[5:0], u_ca_out_893[11:6]};
assign col_out_895 = {u_ca_out_895[5:0], u_ca_out_894[11:6]};
assign col_out_896 = {u_ca_out_896[5:0], u_ca_out_895[11:6]};
assign col_out_897 = {u_ca_out_897[5:0], u_ca_out_896[11:6]};
assign col_out_898 = {u_ca_out_898[5:0], u_ca_out_897[11:6]};
assign col_out_899 = {u_ca_out_899[5:0], u_ca_out_898[11:6]};
assign col_out_900 = {u_ca_out_900[5:0], u_ca_out_899[11:6]};
assign col_out_901 = {u_ca_out_901[5:0], u_ca_out_900[11:6]};
assign col_out_902 = {u_ca_out_902[5:0], u_ca_out_901[11:6]};
assign col_out_903 = {u_ca_out_903[5:0], u_ca_out_902[11:6]};
assign col_out_904 = {u_ca_out_904[5:0], u_ca_out_903[11:6]};
assign col_out_905 = {u_ca_out_905[5:0], u_ca_out_904[11:6]};
assign col_out_906 = {u_ca_out_906[5:0], u_ca_out_905[11:6]};
assign col_out_907 = {u_ca_out_907[5:0], u_ca_out_906[11:6]};
assign col_out_908 = {u_ca_out_908[5:0], u_ca_out_907[11:6]};
assign col_out_909 = {u_ca_out_909[5:0], u_ca_out_908[11:6]};
assign col_out_910 = {u_ca_out_910[5:0], u_ca_out_909[11:6]};
assign col_out_911 = {u_ca_out_911[5:0], u_ca_out_910[11:6]};
assign col_out_912 = {u_ca_out_912[5:0], u_ca_out_911[11:6]};
assign col_out_913 = {u_ca_out_913[5:0], u_ca_out_912[11:6]};
assign col_out_914 = {u_ca_out_914[5:0], u_ca_out_913[11:6]};
assign col_out_915 = {u_ca_out_915[5:0], u_ca_out_914[11:6]};
assign col_out_916 = {u_ca_out_916[5:0], u_ca_out_915[11:6]};
assign col_out_917 = {u_ca_out_917[5:0], u_ca_out_916[11:6]};
assign col_out_918 = {u_ca_out_918[5:0], u_ca_out_917[11:6]};
assign col_out_919 = {u_ca_out_919[5:0], u_ca_out_918[11:6]};
assign col_out_920 = {u_ca_out_920[5:0], u_ca_out_919[11:6]};
assign col_out_921 = {u_ca_out_921[5:0], u_ca_out_920[11:6]};
assign col_out_922 = {u_ca_out_922[5:0], u_ca_out_921[11:6]};
assign col_out_923 = {u_ca_out_923[5:0], u_ca_out_922[11:6]};
assign col_out_924 = {u_ca_out_924[5:0], u_ca_out_923[11:6]};
assign col_out_925 = {u_ca_out_925[5:0], u_ca_out_924[11:6]};
assign col_out_926 = {u_ca_out_926[5:0], u_ca_out_925[11:6]};
assign col_out_927 = {u_ca_out_927[5:0], u_ca_out_926[11:6]};
assign col_out_928 = {u_ca_out_928[5:0], u_ca_out_927[11:6]};
assign col_out_929 = {u_ca_out_929[5:0], u_ca_out_928[11:6]};
assign col_out_930 = {u_ca_out_930[5:0], u_ca_out_929[11:6]};
assign col_out_931 = {u_ca_out_931[5:0], u_ca_out_930[11:6]};
assign col_out_932 = {u_ca_out_932[5:0], u_ca_out_931[11:6]};
assign col_out_933 = {u_ca_out_933[5:0], u_ca_out_932[11:6]};
assign col_out_934 = {u_ca_out_934[5:0], u_ca_out_933[11:6]};
assign col_out_935 = {u_ca_out_935[5:0], u_ca_out_934[11:6]};
assign col_out_936 = {u_ca_out_936[5:0], u_ca_out_935[11:6]};
assign col_out_937 = {u_ca_out_937[5:0], u_ca_out_936[11:6]};
assign col_out_938 = {u_ca_out_938[5:0], u_ca_out_937[11:6]};
assign col_out_939 = {u_ca_out_939[5:0], u_ca_out_938[11:6]};
assign col_out_940 = {u_ca_out_940[5:0], u_ca_out_939[11:6]};
assign col_out_941 = {u_ca_out_941[5:0], u_ca_out_940[11:6]};
assign col_out_942 = {u_ca_out_942[5:0], u_ca_out_941[11:6]};
assign col_out_943 = {u_ca_out_943[5:0], u_ca_out_942[11:6]};
assign col_out_944 = {u_ca_out_944[5:0], u_ca_out_943[11:6]};
assign col_out_945 = {u_ca_out_945[5:0], u_ca_out_944[11:6]};
assign col_out_946 = {u_ca_out_946[5:0], u_ca_out_945[11:6]};
assign col_out_947 = {u_ca_out_947[5:0], u_ca_out_946[11:6]};
assign col_out_948 = {u_ca_out_948[5:0], u_ca_out_947[11:6]};
assign col_out_949 = {u_ca_out_949[5:0], u_ca_out_948[11:6]};
assign col_out_950 = {u_ca_out_950[5:0], u_ca_out_949[11:6]};
assign col_out_951 = {u_ca_out_951[5:0], u_ca_out_950[11:6]};
assign col_out_952 = {u_ca_out_952[5:0], u_ca_out_951[11:6]};
assign col_out_953 = {u_ca_out_953[5:0], u_ca_out_952[11:6]};
assign col_out_954 = {u_ca_out_954[5:0], u_ca_out_953[11:6]};
assign col_out_955 = {u_ca_out_955[5:0], u_ca_out_954[11:6]};
assign col_out_956 = {u_ca_out_956[5:0], u_ca_out_955[11:6]};
assign col_out_957 = {u_ca_out_957[5:0], u_ca_out_956[11:6]};
assign col_out_958 = {u_ca_out_958[5:0], u_ca_out_957[11:6]};
assign col_out_959 = {u_ca_out_959[5:0], u_ca_out_958[11:6]};
assign col_out_960 = {u_ca_out_960[5:0], u_ca_out_959[11:6]};
assign col_out_961 = {u_ca_out_961[5:0], u_ca_out_960[11:6]};
assign col_out_962 = {u_ca_out_962[5:0], u_ca_out_961[11:6]};
assign col_out_963 = {u_ca_out_963[5:0], u_ca_out_962[11:6]};
assign col_out_964 = {u_ca_out_964[5:0], u_ca_out_963[11:6]};
assign col_out_965 = {u_ca_out_965[5:0], u_ca_out_964[11:6]};
assign col_out_966 = {u_ca_out_966[5:0], u_ca_out_965[11:6]};
assign col_out_967 = {u_ca_out_967[5:0], u_ca_out_966[11:6]};
assign col_out_968 = {u_ca_out_968[5:0], u_ca_out_967[11:6]};
assign col_out_969 = {u_ca_out_969[5:0], u_ca_out_968[11:6]};
assign col_out_970 = {u_ca_out_970[5:0], u_ca_out_969[11:6]};
assign col_out_971 = {u_ca_out_971[5:0], u_ca_out_970[11:6]};
assign col_out_972 = {u_ca_out_972[5:0], u_ca_out_971[11:6]};
assign col_out_973 = {u_ca_out_973[5:0], u_ca_out_972[11:6]};
assign col_out_974 = {u_ca_out_974[5:0], u_ca_out_973[11:6]};
assign col_out_975 = {u_ca_out_975[5:0], u_ca_out_974[11:6]};
assign col_out_976 = {u_ca_out_976[5:0], u_ca_out_975[11:6]};
assign col_out_977 = {u_ca_out_977[5:0], u_ca_out_976[11:6]};
assign col_out_978 = {u_ca_out_978[5:0], u_ca_out_977[11:6]};
assign col_out_979 = {u_ca_out_979[5:0], u_ca_out_978[11:6]};
assign col_out_980 = {u_ca_out_980[5:0], u_ca_out_979[11:6]};
assign col_out_981 = {u_ca_out_981[5:0], u_ca_out_980[11:6]};
assign col_out_982 = {u_ca_out_982[5:0], u_ca_out_981[11:6]};
assign col_out_983 = {u_ca_out_983[5:0], u_ca_out_982[11:6]};
assign col_out_984 = {u_ca_out_984[5:0], u_ca_out_983[11:6]};
assign col_out_985 = {u_ca_out_985[5:0], u_ca_out_984[11:6]};
assign col_out_986 = {u_ca_out_986[5:0], u_ca_out_985[11:6]};
assign col_out_987 = {u_ca_out_987[5:0], u_ca_out_986[11:6]};
assign col_out_988 = {u_ca_out_988[5:0], u_ca_out_987[11:6]};
assign col_out_989 = {u_ca_out_989[5:0], u_ca_out_988[11:6]};
assign col_out_990 = {u_ca_out_990[5:0], u_ca_out_989[11:6]};
assign col_out_991 = {u_ca_out_991[5:0], u_ca_out_990[11:6]};
assign col_out_992 = {u_ca_out_992[5:0], u_ca_out_991[11:6]};
assign col_out_993 = {u_ca_out_993[5:0], u_ca_out_992[11:6]};
assign col_out_994 = {u_ca_out_994[5:0], u_ca_out_993[11:6]};
assign col_out_995 = {u_ca_out_995[5:0], u_ca_out_994[11:6]};
assign col_out_996 = {u_ca_out_996[5:0], u_ca_out_995[11:6]};
assign col_out_997 = {u_ca_out_997[5:0], u_ca_out_996[11:6]};
assign col_out_998 = {u_ca_out_998[5:0], u_ca_out_997[11:6]};
assign col_out_999 = {u_ca_out_999[5:0], u_ca_out_998[11:6]};
assign col_out_1000 = {u_ca_out_1000[5:0], u_ca_out_999[11:6]};
assign col_out_1001 = {u_ca_out_1001[5:0], u_ca_out_1000[11:6]};
assign col_out_1002 = {u_ca_out_1002[5:0], u_ca_out_1001[11:6]};
assign col_out_1003 = {u_ca_out_1003[5:0], u_ca_out_1002[11:6]};
assign col_out_1004 = {u_ca_out_1004[5:0], u_ca_out_1003[11:6]};
assign col_out_1005 = {u_ca_out_1005[5:0], u_ca_out_1004[11:6]};
assign col_out_1006 = {u_ca_out_1006[5:0], u_ca_out_1005[11:6]};
assign col_out_1007 = {u_ca_out_1007[5:0], u_ca_out_1006[11:6]};
assign col_out_1008 = {u_ca_out_1008[5:0], u_ca_out_1007[11:6]};
assign col_out_1009 = {u_ca_out_1009[5:0], u_ca_out_1008[11:6]};
assign col_out_1010 = {u_ca_out_1010[5:0], u_ca_out_1009[11:6]};
assign col_out_1011 = {u_ca_out_1011[5:0], u_ca_out_1010[11:6]};
assign col_out_1012 = {u_ca_out_1012[5:0], u_ca_out_1011[11:6]};
assign col_out_1013 = {u_ca_out_1013[5:0], u_ca_out_1012[11:6]};
assign col_out_1014 = {u_ca_out_1014[5:0], u_ca_out_1013[11:6]};
assign col_out_1015 = {u_ca_out_1015[5:0], u_ca_out_1014[11:6]};
assign col_out_1016 = {u_ca_out_1016[5:0], u_ca_out_1015[11:6]};
assign col_out_1017 = {u_ca_out_1017[5:0], u_ca_out_1016[11:6]};
assign col_out_1018 = {u_ca_out_1018[5:0], u_ca_out_1017[11:6]};
assign col_out_1019 = {u_ca_out_1019[5:0], u_ca_out_1018[11:6]};
assign col_out_1020 = {u_ca_out_1020[5:0], u_ca_out_1019[11:6]};
assign col_out_1021 = {u_ca_out_1021[5:0], u_ca_out_1020[11:6]};
assign col_out_1022 = {u_ca_out_1022[5:0], u_ca_out_1021[11:6]};
assign col_out_1023 = {u_ca_out_1023[5:0], u_ca_out_1022[11:6]};
assign col_out_1024 = {u_ca_out_1024[5:0], u_ca_out_1023[11:6]};
assign col_out_1025 = {u_ca_out_1025[5:0], u_ca_out_1024[11:6]};
assign col_out_1026 = {u_ca_out_1026[5:0], u_ca_out_1025[11:6]};
assign col_out_1027 = {u_ca_out_1027[5:0], u_ca_out_1026[11:6]};
assign col_out_1028 = {u_ca_out_1028[5:0], u_ca_out_1027[11:6]};
assign col_out_1029 = {u_ca_out_1029[5:0], u_ca_out_1028[11:6]};
assign col_out_1030 = {u_ca_out_1030[5:0], u_ca_out_1029[11:6]};
assign col_out_1031 = {u_ca_out_1031[5:0], u_ca_out_1030[11:6]};
assign col_out_1032 = {u_ca_out_1032[5:0], u_ca_out_1031[11:6]};
assign col_out_1033 = {{6{1'b0}}, u_ca_out_1032[11:6]};

//---------------------------------------------------------


endmodule
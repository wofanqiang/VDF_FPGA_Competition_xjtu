module xpb_5_505
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h4c9d68f8c6db0250c4c8193e694c78e09584eac1e2ccbd07d9a780423ae84c303910ec0e0caa864ff83357e58305b242b992e0cfc43ff81037f19651848e6025ea26b2e30c7e975d6a4d0796f0e861f3ee504462f6b34a22506f5eb5444d7a782ff42d1e32ebdbc866045cd8792acbabb8df4a494cbfa40452ff8abe17ab4e43;
    5'b00010 : xpb = 1024'h993ad1f18db604a18990327cd298f1c12b09d583c5997a0fb34f008475d098607221d81c19550c9ff066afcb060b64857325c19f887ff0206fe32ca3091cc04bd44d65c618fd2ebad49a0f2de1d0c3e7dca088c5ed669444a0debd6a889af4f05fe85a3c65d7b790cc08b9b0f255975771be9492997f4808a5ff157c2f569c86;
    5'b00011 : xpb = 1024'h352af59492a2d2298352d3e42b8b23504f18bd14d2ee96a00f19c770fdb63788a7ea46b15bd91461493bc869a5b305fdc89e7a892a0d17e4f735839652d8abc04a24e3fa75eac8d32c4d142239dd61aad6ebd3905793b1563bc18a2512bdccd660d4f530e7fa9acbab4d2faa73b03cd9dbc3fff995f38edcb28f2535be1f845e;
    5'b00100 : xpb = 1024'h81c85e8d597dd47a481aed2294d79c30e49da7d6b5bb53a7e8c147b3389e83b8e0fb32bf68839ab1416f204f28b8b84082315b58ee4d0ff52f2719e7d7670be6344b96dd82696030969a1bb92ac5c39ec53c17f34e46fb788c30e8da570b474e90c9224f1ae6769411518c82ecdb088594a34a42e2b332e1058eaff3d5cad2a1;
    5'b00101 : xpb = 1024'h1db882305e6aa20241dd8e89edc9cdc008ac8f67c3107038448c0e9fc08422e116c3a154ab07a2729a4438edc86059b8d7aa14428fda37b9b67970db2122f75aaa231511df56fa48ee4d20ad82d26161bf8762bdb874188a2713b594e12e1f3491b5bd439d0959cef096027c6e35ae07fea8b5a9df2779b5121ebfad6493ba79;
    5'b00110 : xpb = 1024'h6a55eb292545a45306a5a7c8571646a09e317a29a5dd2d401e338ee1fb6c6f114fd48d62b7b228c2927790d34b660bfb913cf512541a2fc9ee6b072ca5b157809449c7f4ebd591a6589a284473bac355add7a720af2762ac7783144a257b99acc1a9ea61cff53597569a5f54e76079b3b787fff32be71db9651e4a6b7c3f08bc;
    5'b00111 : xpb = 1024'h6460ecc2a3271db0068492fb008782fc24061bab33249d079fe55ce83520e39859cfbf7fa363083eb4ca971eb0dad73e6b5adfbf5a7578e75bd5e1fef6d42f50a21462948c32bbeb04d2d38cbc76118a822f1eb19547fbe1265e104af9e7192c2968556521818d235ded54e68bb1f36218d6b5a285b648d71ae5a250b07f094;
    5'b01000 : xpb = 1024'h52e377c4f10d742bc530626e1954f11057c54c7c95ff06d853a5d610be3a5a69beade80606e0b6d3e38001576e135fb6a0488ecbb9e74f9eadaef47173fba31af447f90c5541c31c1a9a34cfbcafc30c9673364e1007c9e062d53fb9f3ebec0af28ab2748503f49a9be33226e1e5eae1da6cb5a3751b0891c4ade4e322b33ed7;
    5'b01001 : xpb = 1024'h9f80e0bdb7e8767c89f87bac82a169f0ed4a373e78cbc3e02d4d5652f922a699f7bed414138b3d23dbb3593cf11911f959db6f9b7e2747aee5a08ac2f88a0340de6eabef61c05a7984e73c66ad98250084c37ab106bb1402b3449e6f38396683227edf92b7efd06301e78eff5b10b68d934bffecc1daac9617ad6fa13a5e8d1a;
    5'b01010 : xpb = 1024'h3b710460bcd5440483bb1d13db939b8011591ecf8620e07089181d3f810845c22d8742a9560f44e5348871db90c0b371af5428851fb46f736cf2e1b64245eeb554462a23beadf491dc9a415b05a4c2c37f0ec57b70e831144e276b29c25c3e69236b7a873a12b39de12c04f8dc6b5c0ffd516b53be4ef36a243d7f5ac92774f2;
    5'b01011 : xpb = 1024'h880e6d5983b046554883365244e01460a6de099168ed9d7862bf9d81bbf091f266982eb762b9cb352cbbc9c113c665b468e70954e3f46783a4e47807c6d44edb3e6cdd06cb2c8bef46e748f1f68d24b76d5f09de679b7b369e96c9df06a9b8e1535fa7a56cfe8f66473061d1559627bbb630b59d0b0e976e773d0a18e0d2c335;
    5'b01100 : xpb = 1024'h23fe90fc889d13dd4245d7b99dd245efcaecf1227642ba08be8a646e43d6311a9c609d4ca53dd2f68590e25fb36e072cbe5fc23e85818f482c36cefb10903a4fb4445b3b281a26079e9a4de64e99c27a67aa54a8d1c898483979969990cc90c7544c4299ef2172a12674d7cad6f0cd3e203621040782de4283cd19d26f9bab0d;
    5'b01101 : xpb = 1024'h709bf9f54f78162e070df0f8071ebed06071dbe4590f77109831e4b07ebe7d4ad571895ab1e859467dc43a453673b96f77f2a30e49c187586428654c951e9a759e6b0e1e3498bd6508e7557d3f82246e55fa990bc87be26a89e8f54ed51a0b3f84406fb8220d4e698c7934a3501b98e9d9156b4d54428246d6cca4908746f950;
    5'b01110 : xpb = 1024'hc8c1d985464e3b600d0925f6010f05f8480c375666493a0f3fcab9d06a41c730b39f7eff46c6107d69952e3d61b5ae7cd6b5bf7eb4eaf1ceb7abc3fdeda85ea14428c529186577d609a5a71978ec2315045e3d632a8ff7c24cbc2095f3ce325852d0aaca43031a46bbdaa9cd1763e6c431ad6b450b6c91ae35cb44a160fe128;
    5'b01111 : xpb = 1024'h592986911b3fe606c598ab9dc95d69401a05ae37493150a8cda42bdf418c68a3444ae3fe0116e757ceccaac959210d2a86fe3cc7af8ea72d236c52916368e60ffe693f359e04eedacae76208887724253e962839295c499e753b20bea38a5d9db52137cad71c0d6cd1c207754aa10a17fbfa20fd9d766d1f365c3f082dbb2f6b;
    5'b10000 : xpb = 1024'ha5c6ef89e21ae8578a60c4dc32a9e220af8a98f92bfe0db0a74bac217c74b4d37d5bd00c0dc16da7c70002aedc26bf6d40911d9773ce9f3d5b5de8e2e7f74635e88ff218aa8386383534699f795f86192ce66c9c200f93c0c5aa7f73e7d7d815e51564e90a07e93537c6644dc3cbd5c3b4d96b46ea361123895bc9c645667dae;
    5'b10001 : xpb = 1024'h41b7132ce707b5df842366438b9c13afd399808a39532a410316730e045a53fbb3243ea1504575691fd51b4d7bce60e59609d681155bc701e2b03fd631b331aa5e67704d077120508ce76e93d16c23dc2731b7668a3cb0d2608d4c2e71faaffbe601ffdd8c2acc70170ada4745267b461eded6ade6aa57f795ebd97fd42f6586;
    5'b10010 : xpb = 1024'h8e547c25ade2b83048eb7f81f4e88c90691e6b4c1c1fe748dcbdf3503f42a02bec352aaf5ceffbb918087332fed413284f9cb750d99bbf121aa1d627b64191d0488e233013efb7adf734762ac25485d01581fbc980effaf4b0fcaae3b6482a7415f62cfbbf16a8387d0f371fbe5146f1d7be20f73369fbfbe8eb643debdab3c9;
    5'b10011 : xpb = 1024'h2a449fc8b2cf85b842ae20e94ddabe1f8d2d52dd297503d93888ba3cc7283f5421fd99449f74037a70dd8bd19e7bb4a0a515703a7b28e6d6a1f42d1afffd7d44be65a16470dd51c64ee77b1f1a6123930fcd4693eb1d18064bdf779e406b025a16e2c7f041398b735c53ad193fabec7441c38c5e2fde42cff57b73f77aa39ba1;
    5'b10100 : xpb = 1024'h76e208c179aa880907763a27b727370022b23d9f0c41c0e112303a7f02108b845b0e8552ac1e89ca6910e3b7218166e35ea8510a3f68dee6d9e5c36c848bdd6aa88c54477d5be923b93482b60b498586fe1d8af6e1d062289c4ed65384b87cd246d6f50e7425673bc25809f1b8d6b81ffaa2d6a77c9de6d4487afeb5924ee9e4;
    5'b10101 : xpb = 1024'h12d22c647e9755910138db8f1019688f46c125301996dd716dfb016b89f62aac90d6f3e7eea2918bc1e5fc55c129085bb42109f3e0f606ab61381a5fce47c8df1e63d27bda49833c10e787aa63562349f868d5c14bfd7f3a3731a30e0edb54b847c39002f6484a76a19c7feb3a315da264a8420e79122da8550b0e6f2117d1bc;
    5'b10110 : xpb = 1024'h5f6f955d457257e1c600f4cd7965e16fdc460ff1fc639a7947a281adc4de76dcc9e7dff5fb4d17dbba19543b442eba9e6db3eac3a535febb9929b0b152d62905088a855ee6c81a997b348f41543e853de6b91a2442b0c95c87a101c35328cf3077b7bd212934263f07a0dcc3b35c294e1d878c57c5d1d1aca80a992d38c31fff;
    5'b10111 : xpb = 1024'hac0cfe560c4d5a328ac90e0be2b25a5071cafab3df305781214a01efffc6c30d02f8cc0407f79e2bb24cac20c7346ce12746cb936975f6cbd11b4702d764892af2b13841f346b1f6e58196d84526e731d5095e873964137ed8106078977649a8a7abea3f5c2002076da5399c2c86f4f9d666d6a1129175b0fb0a23eb506e6e42;
    5'b11000 : xpb = 1024'h47fd21f9113a27ba848baf733ba48bdf95d9e244ec8574117d14c8dc87ac623538c13a994a7ba5ed0b21c4bf66dc0e597cbf847d0b031e90586d9df62120749f6888b67650344c0f3d349bcc9d3384f4cf54a951a391309072f32d332199218ea8988533de42e5424ce9af95ade19a7c406c42080f05bc85079a33a4df37561a;
    5'b11001 : xpb = 1024'h949a8af1d8152a0b4953c8b1a4f104c02b5ecd06cf52311956bc491ec294ae6571d226a757262c3d03551ca4e9e1c09c3652654ccf4316a0905f3447a5aed4c552af69595cb2e36ca781a3638e1be6e8bda4edb49a447ab2c3628be865e69c06d88cb252112ec10ab2ee0c6e270c6627f94b8c515bc560895a99be62f6e2a45d;
    5'b11010 : xpb = 1024'h308aae94dd01f79343166a18fde3364f4f6db497dca74da9b287100b4a7a4d8da79a953c99aa33fe5c2a3543898962148bcb1e3670d03e6517b18b3aef6ac039c886e78db9a07d84ff34a857e62884abb7f0387f047197c45e4558a2f00973ecd9794d469351a44592328267a8670baa6350f7b85839a75d6729ce1c85ab8c35;
    5'b11011 : xpb = 1024'h7d28178da3dcf9e407de8357672faf2fe4f29f59bf740ab18c2e904d856299bde0ab814aa654ba4e545d8d290c8f1457455dff06351036754fa3218c73f9205fb2ad9a70c61f14e26981afeed710e69fa6407ce1fb24e1e6aeb4b7583456ee65096d7a64c63d800df836df402191d7561c304201a4f94b61ba2958da9d56da78;
    5'b11100 : xpb = 1024'h19183b30a8c9c76c01a124bec021e0bf090186eaccc92741e7f9573a0d4838e61673efdfe8d8c20fad32a5c7ac36b5cf9ad6b7efd69d5e39d6f5787fbdb50bd4288518a5230caefac134b4e32f1d8462a08bc7ac6551fef849978412be79c64b0a5a155948606348d77b5539a2ec7cd88635ad68a16d9235c6b968942c1fc250;
    5'b11101 : xpb = 1024'h65b5a4296fa4c9bcc6693dfd296e599f9e8671acaf95e449c1a0d77c483085164f84dbedf583485fa565fdad2f3c6812546998bf9add564a0ee70ed142436bfa12abcb882f8b46582b81bc7a2005e6568edc0c0f5c05491a9a06e2c802c740c33a4e42777b4c3f113d7fb2121c1748843f14f7b1ee2d363a19b8f35243cb1093;
    5'b11110 : xpb = 1024'h1a5c7cc74919744c02bdf6482608b2ec295593dbceb00da1d6b9e68d016243e854d4a8338075020fe3b164bcee4098aa9e251a93c6a7e0e963965c48bff576e888349bc8c78e0708334c16e78128419892756d9c632662c34e9af828cea18a93b3add6bfd6f224c1cc4280b9d71ee06a91a6318eaa17d0e2649030bd293f86b;
    5'b11111 : xpb = 1024'h4e4330c53b6c999584f3f8a2ebad040f581a43ff9fb7bde1f7131eab0afe706ebe5e369144b1d670f66e6e3151e9bbcd6375327900aa761ece2afc16108db79472a9fc9f98f777cded81c90568fae60d77779b3cbce5b04e85590e37d13793216b2f0a8a305afe1482c884e4169cb9b261f9ad623761211279488dc9ea3f46ae;
    endcase
end

endmodule

module xpb_5_810
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h68a1bb3bcfba5151431cec300048119e0d1c2257d30314beba4be73898e1f1f0f9439adc2acc0c63aa7684fc69ef610e6182ac6bd1a39165814b93227bddf8a62fc34afedc4a5fc19a6a46bed364f0a63d9e69ad3d859dc1d8dff6f8b4bfc09e5978e70465ab8d7caef30b4cac9698fa4a8fe86dbb243737bdb4d5af8e6ab074;
    5'b00010 : xpb = 1024'h20963121dd866dd9bb346088f035dbeaa8c2417ed08e8905f6bb151b7ec136d9ef3eb83f8b719a38b58ecab1f080b1525eeb30f18094527f51f7e6e6bce97c9aeb37614f0903c23e223a8adb0dee1d1b8737d9c1ee850e72fc335bf6af54deaa83ea3bdf1a8e226bd7262fba615d0bcb4645f1f925fd113f34fa305a93f2fa7d;
    5'b00011 : xpb = 1024'h8937ec5dad40bf2afe514cb8f07ded88b5de63d6a3919dc4b106fc5417a328cae882531bb63da69c60054fae5a701260c06ddd5d5237e3e4d3437a0938c775411afaac4de54e21ffbca4d199e1530dc1c4d6436f2c0aac34d51352ef64149f48dd6322e38039afe886193b070df3a4c590d5da66e1214876f2af060a225daaf1;
    5'b00100 : xpb = 1024'h412c6243bb0cdbb37668c111e06bb7d5518482fda11d120bed762a36fd826db3de7d707f16e334716b1d9563e10162a4bdd661e30128a4fea3efcdcd79d2f935d66ec29e1207847c447515b61bdc3a370e6fb383dd0a1ce5f866b7ed5ea9bd5507d477be351c44d7ae4c5f74c2ba17968c8be3f24bfa227e69f460b527e5f4fa;
    5'b00101 : xpb = 1024'ha9ce1d7f8ac72d04b985ad41e0b3c9735ea0a555742026caa7c2116f96645fa4d7c10b5b41af40d515941a604af0c3b31f590e4ed2cc3664253b60eff5b0f1dc06320d9cee51e43ddedf5c74ef412add4c0e1d311a8fbaa7d146aee613697df3614d5ec29ac7d2545d3f6ac16f50b090d71bcc60071e59b627a93664b650a56e;
    5'b00110 : xpb = 1024'h61c293659893498d319d219ad0a193bffa46c47c71ab9b11e4313f527c43a48dcdbc28bea254ceaa20ac6015d18213f71cc192d481bcf77df5e7b4b436bc75d0c1a623ed1b0b46ba66afa09129ca575295a78d45cb8f2b58f49a13e40dfe9bff8bbeb39d4faa674385728f2f24172361d2d1d5eb71f733bd9eee910fbbd8ef77;
    5'b00111 : xpb = 1024'h19b7094ba65f6615a9b495f3c08f5e0c95ece3a36f370f5920a06d356222e976c3b7462202fa5c7f2bc4a5cb5813643b1a2a175a30adb897c694087877c7f9c57d1a3a3d47c4a936ee7fe4ad645383c7df40fd5a7c8e9c0a17ed78e20893ba0bb6300878048cfc32ada5b39cd8dd9632ce87df76dcd00dc51633ebbac1613980;
    5'b01000 : xpb = 1024'h8258c4877619b766ecd18223c0d76faaa30905fb423a2417daec546dfb04db67bcfae0fe2dc668e2d63b2ac7c202c5497bacc3c6025149fd47df9b9af3a5f26bacdd853c240f08f888ea2b6c37b8746e1cdf6707ba1439cbf0cd6fdabd537aaa0fa8ef7c6a3889af5c98bee985742f2d1917c7e497f444fcd3e8c16a4fcbe9f4;
    5'b01001 : xpb = 1024'h3a4d3a6d83e5d3ef64e8f67cb0c539f73eaf25223fc5985f175b8250e0e42050b2f5fe618e6bf6b7e153707d4894158d7915484bb1420b17188bef5f34b1766068519b8c50c86b7510ba6f887241a0e36678d71c6b13aa7d1420d4d8b7e898b63a1a44571f1b1e9e84cbe3573a3aa1fe14cdd17002cd1f044b2e1c15555433fd;
    5'b01010 : xpb = 1024'ha2eef5a953a02540a805e2acb10d4b954bcb477a12c8ad1dd1a7698979c61241ac39993db938031b8bc9f579b283769bda97f4b782e59c7c99d78281b08f6f069814e68b2d12cb36ab24b64745a69189a41740c9a899483eed00cbd16ca8595493932b5b84c6ac1b33beeea3e6d13af85f5db9ddbdf1563c08e2f1c4e3bee471;
    5'b01011 : xpb = 1024'h5ae36b8f616c41c9201d5705a0fb15e1e77166a1105421650e16976c5fa5572aa234b6a119dd90f096e23b2f3914c6dfd800793d31d65d966a83d645f19af2fb5388fcdb59cc2db332f4fa63802fbdfeedb0b0de5998b8f0105430cf673d7760be04803639a9410a5bf213119b97adc95b13c36928ca304380284c6fe9472e7a;
    5'b01100 : xpb = 1024'h12d7e1756f385e519834cb5e90e8e02e831785c80ddf95ac4a85c54f45849c13982fd4047a831ec5a1fa80e4bfa61723d568fdc2e0c71eb03b302a0a32a676f00efd132b8685902fbac53e7fbab8ea74374a20f30a9829a133a795cd61d2956ce875d510ee8bd5f98425377f505e209a56c9ccf493a30a4af76da71aeecf7883;
    5'b01101 : xpb = 1024'h7b799cb13ef2afa2db51b78e9130f1cc9033a81fe0e2aa6b04d1ac87de668e0491736ee0a54f2b294c7105e12995783236ebaa2eb26ab015bc7bbd2cae846f963ec05e2a62cfeff1552f853e8e1ddb1a74e88aa0481dc7630c878cc61692560b41eebc1554376376331842cbfcf4b994a159b5624ec74182b5227cca7d3a28f7;
    5'b01110 : xpb = 1024'h336e12974cbecc2b53692be7811ebc192bd9c746de6e1eb24140da6ac445d2ed876e8c4405f4b8fe57894b96b026c87634542eb4615b712f8d2810f0ef8ff38afa34747a8f89526ddcffc95ac8a7078fbe81fab4f91d38142fdaf1c4112774176c6010f00919f8655b4b6739b1bb2c659d0fbeedb9a01b8a2c67d77582c27300;
    5'b01111 : xpb = 1024'h9c0fcdd31c791d7c968618178166cdb738f5e99eb1713370fb8cc1a35d27c4de80b2272030c0c56201ffd0931a16298495d6db2032ff02950e73a4136b6dec3129f7bf796bd3b22f776a10199c0bf835fc20646236a2d5d608bae8bcc5e734b5c5d8f7f46ec585e20a3e72865e51c55fe79fa75b74c452c1ea1cad25112d2374;
    5'b10000 : xpb = 1024'h540443b92a453a050e9d8c7071549803d49c08c5aefca7b837fbef86430709c776ad4483916653370d181648a0a779c8933f5fa5e1efc3aedf1ff7d7ac797025e56bd5c9988d14abff3a5435d69524ab45b9d476e7a246872c0e4dbac07c52c1f04a4ccf23a81ad1327196f413183830e355b0e6df9d2cc9616207d016b56d7d;
    5'b10001 : xpb = 1024'hbf8b99f3811568d86b500c961426250704227ecac881bff746b1d6928e64eb06ca861e6f20be10c18305bfe2738ca0c90a7e42b90e084c8afcc4b9bed84f41aa0dfec19c5467728870a9852111e51208f53448b98a1b7384f61b2b8bb1170ce1abba1a9d88aafc05aa4bb61c7deab01df0bba724a7606d0d8a7627b1c3db786;
    5'b10010 : xpb = 1024'h749a74db07cba7dec9d1ecf9618a73ee7d5e4a447f8b30be2eb704a1c1c840a165ebfcc31cd7ed6fc2a6e0fa91282b1af22a90976284162e3117debe6962ecc0d0a33718a190d6ea2174df10e48341c6ccf1ae38d62754fa2841a9b16fd1316c743488ae3e363d3d0997c6ae747543fc299ba2e0059a3e08965c382aaaa867fa;
    5'b10011 : xpb = 1024'h2c8eeac11597c46741e9615251783e3b1904696b7d16a5056b263284a7a7858a5be71a267d7d7b44cdbf26b017b97b5eef93151d1174d74801c43282aa6e70b58c174d68ce4a3966a945232d1f0c6e3c168b1e4d8726c5ab4b950eaf6a664f789ea5dd88f318d22c31caeb1c293bb6cd2551ac6b707318100da192d5b030b203;
    5'b10100 : xpb = 1024'h9530a5fce55215b885064d8251c04fd926208bc35019b9c4257219bd4089777b552ab502a84987a87835abac81a8dc6d5115c188e31868ad830fc5a5264c695bbbda9867aa94992843af69ebf2715ee2542987fac4ac636d247505a81f261016f81ec48d58c45fa8e0bdf668d5d24fc76fe194d92b974f47cb5668853e9b6277;
    5'b10101 : xpb = 1024'h4d251be2f31e3240fd1dc1db41ae1a25c1c6aaea4da52e0b61e147a02668bc644b25d26608ef157d834df162083a2cb14e7e460e920929c753bc19696757ed50774eaeb7d74dfba4cb7fae082cfa8b579dc2f80f75abd41e47c86aa619bb2e23229019680da6f49808f11ad68a98c2986b979e649670294f429bc3304423ac80;
    5'b10110 : xpb = 1024'h51991c900ea4ec975353634319be4725d6cca114b30a2529e5075830c48014d4120efc96994a3528e6637178ecb7cf54be6ca9440f9eae124686d2da863714532c2c50804075e21534ff2246783b7cce75c682426ab44cf6b1bcfa414504c2f4d016e42c289898731243f443f5f3569674da7f001490356b9e11ddb49abf689;
    5'b10111 : xpb = 1024'h6dbb4d04d0a4a01ab852226431e3f6106a88ec691e33b711589c5cbba529f33e3a648aa59460afb638dcbc13f8bade03ad697700129d7c46a5b40050244169eb62861006e051bde2edba38e33ae8a87324fad1d16430e29143fbc69cc9100ccda67a554728351703e0174a90ebf5ce63b1dd905dbc6d3a8e7795f38ad816a6fd;
    5'b11000 : xpb = 1024'h25afc2eade70bca3306996bd21d1c05d062f0b901bbf2b58950b8a9e8b093827305fa808f5063d8b43f501c97f4c2e47aad1fb85c18e3d6076605414654cede01dfa26570d0b205f758a7cff7571d4e86e9441e615305342674f2b9ac3a52ad9d0ebaa21dd17abf3084a6efea0bc4134ad9399e927461495eedb4e35dd9ef106;
    5'b11001 : xpb = 1024'h8e517e26ae2b0df4738682ed2219d1fb134b2de7eec240174f5771d723eb2a1829a342e51fd249eeee6b86c5e93b8f560c54a7f19331cec5f7abe736e12ae6864dbd7155e95580210ff4c3be48d6c58eac32ab9352b5f104402f22937864eb782a64912642c3396fb73d7a4b4d52da2ef8238256e26a4bcdac9023e56c09a17a;
    5'b11010 : xpb = 1024'h4645f40cbbf72a7ceb9df74612079c47aef14d0eec4db45e8bc69fba09ca6f011f9e60488077d7c3f983cc7b6fccdf9a09bd2c7742228fdfc8583afb22366a7b093187a6160ee29d97c507da835ff203f5cc1ba803b561b56382879172fa098454d5e600f7a5ce5edf709eb902194cfff3d98be24d4325d523d57e907191eb83;
    5'b11011 : xpb = 1024'haee7af488bb17bce2ebae376124fade5bc0d6f66bf50c91d461286f2a2ac60f218e1fb24ab43e427a3fa5177d9bc40a86b3fd8e313c6214549a3ce1d9e14632138f4d2a4f259425f322f4e9956c4e2aa336a8555413aff773c627e8a27b9ca22ae4ecd055d515bdb8e63aa05aeafe5fa3e69745008675d0ce18a543ffffc9bf7;
    5'b11100 : xpb = 1024'h66dc252e997d9856a6d257cf023d783257b38e8dbcdc3d648281b4d5888ba5db0edd18880be971fcaf12972d604d90ec68a85d68c2b6e25f1a5021e1df1fe715f468e8f51f12a4dbb9ff92b5914e0f1f7d03f569f23a70285fb5e388224ee82ed8c021e01233f0cab696ce73637658cb3a1f7ddb7340371458cfaeeb0584e600;
    5'b11101 : xpb = 1024'h1ed09b14a749b4df1ee9cc27f22b427ef359adb4ba67b1abbef0e2b86e6aeac404d835eb6c8effd1ba2adce2e6dee1306610e1ee71a7a378eafc75a6202b6b0aafdcff454bcc075841cfd6d1cbd73b94c69d657ea339e0d9830948861ce4063b033176bac71685b9dec9f2e1183ccb9c35d58766de19111bd01509960b0d3009;
    5'b11110 : xpb = 1024'h87725650770406306206b857f273541d0075d00c8d6ac66a793cc9f1074cdcb4fe1bd0c7975b0c3564a161df50ce423ec7938e5a434b34de6c4808c89c0963b0dfa04a4428166719dc3a1d909f3c2c3b043bcf2be0bf7e9b5be93f7ed1a3c6d95caa5dbf2cc213368dbcfe2dc4d3649680656fd4993d48538dc9df459977e07d;
    5'b11111 : xpb = 1024'h3f66cc3684d022b8da1e2cb0e2611e699c1bef338af63ab1b5abf7d3ed2c219df416ee2af8009a0a6fb9a794d75f9282c4fc12dff23bf5f83cf45c8cdd14e7a59b14609454cfc996640a61acd9c558b04dd53f4091beef4c7f3ca47ccc38e4e5871bb299e1a4a825b5f0229b7999d7677c1b79600416225b050f39f09f002a86;
    endcase
end

endmodule

module xpb_5_750
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h962bad4fd9be8ec5ffbcc4f81e2fa2a8705b6c7e0a294f6013b389d7288558f1e336d8f7d3be0562791a336251e84dfb67e946107ecf76ea4ad554c3a5dd39ddcaca299cebb0a55ab08999b3335aa6bd1f5870c78ee3f844da5276b80912f9940fdeef67adf11b4a5ca6e9160e6ade561da325a1a1b38070e61b6c5f31df3350;
    5'b00010 : xpb = 1024'h7baa1549f18ee8c3347412192c04fdff6f40d5cb3edafe48a98a5a589e0804dbc3253476dd558c3652d6277dc0728b2c6bb8643adaec1d88e50b6a2910e7ff0a21451e8b27d04d704e7930c3cdd989494aabe7f69141c378ff185b7557fb5095f0b64ca5ab193e07328deb4d25059682ec6c6c60f31ba3b185c75db9dadc0035;
    5'b00011 : xpb = 1024'h61287d44095f42c0692b5f3a39da59566e263f18738cad313f612ada138ab0c5a3138ff5e6ed130a2c921b992efcc85d6f8782653708c4277f417f8e7bf2c43677c0137963eff585ec68c7d468586bd575ff5f25939f8ead23de4032a6e3a797d18da9e3a84160c40874ed843ba04eafbb35b3204483c6f225734f1483d8cd1a;
    5'b00100 : xpb = 1024'h46a6e53e212f9cbd9de2ac5b47afb4ad6d0ba865a83e5c19d537fb5b890d5caf8301eb74f08499de064e0fb49d87058e7356a08f93256ac6197794f3e6fd8962ce3b0867a00f9d9b8a585ee502d74e61a152d65495fd59e148a424eff5cbfe99b2650721a5698380de5befbb523b06dc89fef9df95ebea32c51f406f2cd599ff;
    5'b00101 : xpb = 1024'h2c254d3838fff6bad299f97c558510046bf111b2dcf00b026b0ecbdcfe90089962f046f3fa1c20b1e00a03d00c1142bf7725beb9ef421164b3adaa5952084e8f24b5fd55dc2f45b12847f5f59d5630edcca64d83985b25156d6a09ad44b4559b933c645fa291a63db442f1f268d5bf0958c8409ee7540d7364cb31c9d5d266e4;
    5'b00110 : xpb = 1024'h11a3b53250d050b80751469d635a6b5b6ad67b0011a1b9eb00e59c5e7412b48342dea27303b3a785b9c5f7eb7a9b7ff07af4dce44b5eb8034de3bfbebd1313bb7b30f244184eedc6c6378d0637d51379f7f9c4b29ab8f049922fee6a939cac9d7413c19d9fb9c8fa8a29f4297f7077362791875e38bc30b4047723247ecf33c9;
    5'b00111 : xpb = 1024'ha7cf62822a8edf7e070e0b95818a0e03db31e77e1bcb094b149926359c980d7526157b6ad771ace832e02b4dcc83cdebe2de22f4ca2e2eed98b9148262f04d9945fb1be103ff932176c126b96b2fba371752357a299ce88e6c8265229cafa63183f2b1054daae444e6d0dd3f8ddb558c4534acffda6fb124ea928f83b0ae6719;
    5'b01000 : xpb = 1024'h8d4dca7c425f397b3bc558b68f5f695ada1750cb507cb833aa6ff6b7121ab95f0603d6e9e10933bc0c9c1f693b0e0b1ce6ad411f264ad58c32ef29e7cdfb12c59c7610cf401f3b3714b0bdca05ae9cc342a5aca92bfab3c2914849dfeb97fd3364ca0e434ad30701bcb7df76a4760db913fdf3bf2bd7d4658a3e80de59ab33fe;
    5'b01001 : xpb = 1024'h72cc32765a2f9378707ca5d79d34c4b1d8fcba18852e671c4046c738879d6548e5f23268eaa0ba8fe6581384a998484dea7c5f4982677c2acd253f4d3905d7f1f2f105bd7c3ee34cb2a054daa02d7f4f6df923d82e587ef6b60e2e9d3a80543545a16b8147fb29be929ee1adbb10c5e5e2c73a7e7d3ff7a629ea723902a800e3;
    5'b01010 : xpb = 1024'h584a9a7071ffed75a533f2f8ab0a2008d7e22365b9e01604d61d97b9fd201132c5e08de7f4384163c01407a01822857eee4b7d73de8422c9675b54b2a4109d1e496bfaabb85e8b62508febeb3aac61db994c9b0730b64a2adad4135a8968ab372678c8bf45234c7b6885e3e4d1ab7e12b190813dcea81ae6c9966393aba4cdc8;
    5'b01011 : xpb = 1024'h3dc9026a89d04772d9eb4019b8df7b5fd6c78cb2ee91c4ed6bf4683b72a2bd1ca5cee966fdcfc83799cffbbb86acc2aff21a9b9e3aa0c96801916a180f1b624a9fe6ef99f47e3377ee7f82fbd52b4467c4a012363314155eff99f817d8510239075025fd424b6f383e6ce61be846363f8059c7fd20103e27694254ee54a19aad;
    5'b01100 : xpb = 1024'h23476a64a1a0a1700ea28d3ac6b4d6b6d5acf600234373d601cb38bce825690685bd44e607674f0b738befd6f536ffe0f5e9b9c896bd70069bc77f7d7a262776f661e488309ddb8d8c6f1a0c6faa26f3eff389653571e093245fdcd52739593ae827833b3f7391f51453e852fee0ee6c4f230ebc7178616808ee4648fd9e6792;
    5'b01101 : xpb = 1024'h8c5d25eb970fb6d4359da5bd48a320dd4925f4d57f522be97a2093e5da814f065aba06510fed5df4d47e3f263c13d11f9b8d7f2f2da16a535fd94e2e530eca34cdcd9766cbd83a32a5eb11d0a2909801b47009437cfabc74925c1927621b03cc8fee0793c9bb4b1ea3aea8a157ba6991dec557bc2e084a8a89a37a3a69b3477;
    5'b01110 : xpb = 1024'h9ef17fae932f8a3343169f53f2b9d4b644edcbcb621e721eab559315862d6de248e2795ce4bcdb41c6621754b5a98b0d61a21e0371a98d8f80d2e9a68b0e268117a70313586e28fddae84ad03d83b03d3a9f715bc6b3a40c2378384a7f34a9d0d8ddcfe0ea8ccffc46e1d3a023e684ef3b8f7b1d649405198eb5a402d87a67c7;
    5'b01111 : xpb = 1024'h846fe7a8aaffe43077cdec75008f300d43d3351896d02107412c6396fbb019cc28d0d4dbee546215a01e0b702433c83e65713c2dcdc6342e1b08ff0bf618ebad6e21f801948dd11378d7e1e0d80292c965f2e88ac9116f40483e1d07ce1d00d2b9b52d1ee7b4f2b91cc8d5d73a813d1c0a58c1dcb5fc285a2e61955d817734ac;
    5'b10000 : xpb = 1024'h69ee4fa2c2d03e2dac8539960e648b6442b89e65cb81cfefd70334187132c5b608bf305af7ebe8e979d9ff8b92be056f69405a5829e2daccb53f14716123b0d9c49cecefd0ad792916c778f17281755591465fb9cb6f3a746d0401c51d0557d49a8c8a5ce4dd1575f2afd80e511bf548d922089c07644b9ace0d86b82a740191;
    5'b10001 : xpb = 1024'h4f6cb79cdaa0982ae13c86b71c39e6bb419e07b300337ed86cda0499e6b5719fe8ad8bda01836fbd5395f3a7014842a06d0f788285ff816b4f7529d6cc2e76061b17e1de0ccd213eb4b710020d0057e1bc99d6e8cdcd05a891c9e6826bedaed67b63e79ae2053832c896da4567b6ad75a7eb4f5b58cc6edb6db97812d370ce76;
    5'b10010 : xpb = 1024'h34eb1f96f270f22815f3d3d82a0f42124083710034e52dc102b0d51b5c381d89c89be7590b1af6912d51e7c26fd27fd170de96ace21c2809e9ab3f3c37393b327192d6cc48ecc95452a6a712a77f3a6de7ed4e17d02ad0dcb68fcb3fbad605d85c3b44d8df2d5aef9e7ddc7c7e5165a276b4961aaa34921c0d65696d7c6d9b5b;
    5'b10011 : xpb = 1024'h1a6987910a414c254aab20f937e49d693f68da4d6996dca99887a59cd1bac973a88a42d814b27d65070ddbddde5cbd0274adb4d73e38cea883e154a1a244005ec80dcbba850c7169f0963e2341fe1cfa1340c546d2889c10db55affd09be5cda3d12a216dc557dac7464deb394ec1dcf457ddcd9fb9cb55cad115ac8256a6840;
    5'b10100 : xpb = 1024'hb09534e0e3ffdaeb4a67e5f156144011afc446cb73c02c09ac3b2f73fa4022658bc11bcfe87082c780280f4030450afddc96fae7bd084592ceb6a96548213a3c92d7f55770bd16c4a11fd7d67558c3b73299360e616c9455b5a826b512d1566e4cf1917e8a4698f6d10bc7c9a356fc256321027b9d5035cd932cc72757499b90;
    5'b10101 : xpb = 1024'h96139cdafbd034e87f1f331263e99b68aea9b018a871daf24211fff56fc2ce4f6baf774ef208099b59e4035b9ecf482ee06619121924ec3168ecbecab32bff68e952ea45acdcbeda3f0f6ee70fd7a6435decad3d63ca5f89da6e0b7261b9ad702dc8eebc876ebbb3a6f2ca00b9f1b45231ea493aeeb8590e32d8b88200466875;
    5'b10110 : xpb = 1024'h7b9204d513a08ee5b3d6803371bef6bfad8f1965dd2389dad7e8d076e5457a394b9dd2cdfb9f906f339ff7770d59855fe435373c754192d00322d4301e36c4953fcddf33e8fc66efdcff05f7aa5688cf8940246c66282abdff33f02fb0a204720ea04bfa8496de707cd9cc37d08c6c7f00b38ffa40207c4ed284a9dca943355a;
    5'b10111 : xpb = 1024'h61106ccf2b70e8e2e88dcd547f945216ac7482b311d538c36dbfa0f85ac826232b8c2e4d053717430d5beb927be3c290e8045566d15e396e9d58e995894189c19648d422251c0f057aee9d0844d56b5bb4939b9b6885f5f223f9d4ecff8a5b73ef77a93881bf012d52c0ce6ee72724abcf7cd6b991889f8f72309b375240023f;
    5'b11000 : xpb = 1024'h468ed4c9434142e01d451a758d69ad6dab59ec004686e7ac03967179d04ad20d0b7a89cc0ece9e16e717dfadea6dffc1ebd373912d7ae00d378efefaf44c4eedecc3c910613bb71b18de3418df544de7dfe712ca6ae3c12648bfb9aa4e72b275d04f06767ee723ea28a7d0a5fdc1dcd89e461d78e2f0c2d011dc8c91fb3ccf24;
    5'b11001 : xpb = 1024'h2c0d3cc35b119cdd51fc67969b3f08c4aa3f554d7b389694996d41fb45cd7df6eb68e54b186624eac0d3d3c958f83cf2efa291bb899786abd1c514605f57141a433ebdfe9d5b5f30b6cdcb2979d330740b3a89f96d418c5a6d859e679d5b0977b12663b47c0f46a6fe8ed2dd145c95056d0f64383458e610b1887deca4399c09;
    5'b11010 : xpb = 1024'h118ba4bd72e1f6da86b3b4b7a914641ba924be9aafea457d2f44127cbb5029e0cb5740ca21fdabbe9a8fc7e4c7827a23f371afe5e5b42d4a6bfb29c5ca61d94699b9b2ecd97b074654bd623a14521300368e01286f9f578e924b8324ec43607991fdc0f279376963d475d5142af74d323bd8aaf785c1095151346f474d3668ee;
    5'b11011 : xpb = 1024'ha7b7520d4ca085a0867079afc74406c419802b18ba1394dd42f79c53e3d582d2ae8e19c1f5bbb12113a9fb47196ac81f5b5af5f66483a434b6d07e89703f13246483dc89c52baca10546fbed47acb9bd55e671effe834fd36c9df9dcf5565a0da1dcb05a272884ae311cbe2a39622b88597bd099277489c2374fdba67f159c3e;
    5'b11100 : xpb = 1024'h8d35ba076470df9dbb27c6d0d519621b18659465eec543c5d8ce6cd559582ebc8e7c7540ff5337f4ed65ef6287f505505f2a1420c0a04ad3510693eedb49d850bafed178014b54b6a33692fde22b9c498139e91f00e11b079163de9a443eb10f82b40d982450a76b0703c0614ffce3b52845175878dcad02d6fbcd0128126923;
    5'b11101 : xpb = 1024'h72b422017c41399aefdf13f1e2eebd72174afdb32376f2ae6ea53d56cedadaa66e6ad0c008eabec8c721e37df67f428162f9324b1cbcf171eb3ca95446549d7d1179c6663d6afccc41262a0e7caa7ed5ac8d604e033ee63bb629c35793270811638b6ad62178ca27dceac29866979be1f70e5e17ca44d04376a7be5bd10f3608;
    5'b11110 : xpb = 1024'h583289fb9411939824966112f0c418c9163067005828a197047c0dd8445d86904e592c3f1282459ca0ddd79965097fb266c8507578d998108572beb9b15f62a967f4bb54798aa4e1df15c11f17296161d7e0d77d059cb16fdaefa814e20f5f134462c8141ea0ece4b2d1c4cf7d32540ec5d7a4d71bacf3841653afb67a0c02ed;
    5'b11111 : xpb = 1024'h3db0f1f5abe1ed95594dae33fe9974201515d04d8cda507f9a52de59b9e0327a2e4787be1c19cc707a99cbb4d393bce36a976e9fd4f63eaf1fa8d41f1c6a27d5be6fb042b5aa4cf77d05582fb1a843ee03344eac07fa7ca3ffb58cd230f7b615253a25521bc90fa188b8c70693cd0c3b94a0eb966d1516c4b5ffa1112308cfd2;
    endcase
end

endmodule

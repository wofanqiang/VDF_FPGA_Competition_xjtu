module xpb_5_805
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h195ab68496bb9923a379965c620d89771e97a178d9470cb4e58df6647b27653088332c85fa9b3034f13f7c10bfbb3d21bf8f5a6022e37694a21e4484db393e5b600800edccd472a6af26928a49b6a00b506d92807b7cf290257891f71ceb525738acb97d59467b7d964f9536445eb98cfc2fbb1fb7e28d5fc6bb960e0d8fa251;
    5'b00010 : xpb = 1024'h32b56d092d77324746f32cb8c41b12ee3d2f42f1b28e1969cb1becc8f64eca611066590bf5366069e27ef8217f767a437f1eb4c045c6ed29443c8909b6727cb6c01001db99a8e54d5e4d2514936d4016a0db2500f6f9e5204af123ee39d6a4ae715972fab28cf6fb2c9f2a6c88bd7319f85f763f6fc51abf8d772c1c1b1f44a2;
    5'b00011 : xpb = 1024'h4c10238dc432cb6aea6cc31526289c655bc6e46a8bd5261eb0a9e32d71762f9198998591efd1909ed3be74323f31b7653eae0f2068aa63bde65acd8e91abbb12201802c9667d57f40d73b79edd23e021f148b7817276d7b07069b5e556c1f705aa062c780bd37278c2eebfa2cd1c2ca6f48f315f27a7a81f5432c22a28aee6f3;
    5'b00100 : xpb = 1024'h656ada125aee648e8de65971883625dc7a5e85e3651c32d39637d991ec9d94c220ccb217ea6cc0d3c4fdf042feecf486fe3d69808b8dda52887912136ce4f96d802003b73351ca9abc9a4a2926da802d41b64a01edf3ca4095e247dc73ad495ce2b2e5f56519edf6593e54d9117ae633f0beec7edf8a357f1aee5838363e8944;
    5'b00101 : xpb = 1024'h7ec59096f1a9fdb2315fefcdea43af5398f6275c3e633f887bc5cff667c4f9f2a8ffde9de507f108b63d6c53bea831a8bdccc3e0ae7150e72a975698481e37c8e02804a500263d416bc0dcb3709120389223dc826970bcd0bb5ad9d390989bb41b5f9f72be606973ef8dea0f55d99fc0eceea79e976cc2dee1a9ee4643ce2b95;
    5'b00110 : xpb = 1024'h9820471b886596d5d4d9862a4c5138cab78dc8d517aa4c3d6153c65ae2ec5f2331330b23dfa3213da77ce8647e636eca7d5c1e40d154c77bccb59b1d2357762440300592ccfaafe81ae76f3dba47c043e2916f02e4edaf60e0d36bcaad83ee0b540c58f017a6e4f185dd7f459a38594de91e62be4f4f503ea8658454515dcde6;
    5'b00111 : xpb = 1024'hcdb84a5d32fb30ad4da4af9e047af064af671d1b79b87ac9050369ab11174bb61dba311017d2e3f95e252e5ac09b21d8d150bad1856dc4be34a043c3be3fce2be8d1d1ea3e2549b773ff256b229c1e3efa07ead3e474e050bf6bc710449dd05db18043c02467e1956d2d9ce6c6ecb196743efbb6e6806e28b19f5dd60b09cc;
    5'b01000 : xpb = 1024'h1a286ecef3ee945450c73b0c0012046783470895f4c0c52fae92f9ce26387c7c3e50e6b70ab30318ea9da13f1a7bd8439860ab1af468e4596052e4c89ef77e298bf0d2bfb71297f0669a91afb4d93c298f679a6b4f6167707637fdbe2d2ff027965e39c1196ae35f2bbcc2d32b25a63e92a3fa1b6ec90dcdef6d356be39aac1d;
    5'b01001 : xpb = 1024'h338325538aaa2d77f440d168621f8ddea1deaa0ece07d1e49420f032a15fe1acc684133d054e334ddbdd1d4fda37156557f0057b174c5aee0271294d7a30bc84ebf8d3ad83e70a9715c12439fe8fdc34dfd52cebcade5a009bb08fb54a1b427ecf0af33e72b15edcc20c58096f845fcb8ed3b53b26ab9b2db628cb79f12a4e6e;
    5'b01010 : xpb = 1024'h4cdddbd82165c69b97ba67c4c42d1755c0764b87a74ede9979aee6971c8746dd4eb73fc2ffe96382cd1c996099f25287177f5fdb3a2fd182a48f6dd25569fae04c00d49b50bb7d3dc4e7b6c448467c403042bf6c465b4c90c12921ac670694d607b7acbbcbf7da5a585bed3fb3e319588b03705ade8e288d7ce46187feb9f0bf;
    5'b01011 : xpb = 1024'h6638925cb8215fbf3b33fe21263aa0ccdf0ded008095eb4e5f3cdcfb97aeac0dd6ea6c48fa8493b7be5c157159ad8fa8d70eba3b5d13481746adb25730a3393bac08d5891d8fefe4740e494e91fd1c4b80b051ecc1d83f20e6a1b3a383f1e72d40646639253e55d7eeab8275f841d2e587332b7a9670b5ed439ff7960c499310;
    5'b01100 : xpb = 1024'h7f9348e14edcf8e2dead947d88482a43fda58e7959dcf80344cad36012d6113e5f1d98cef51fc3ecaf9b91821968ccca969e149b7ff6beabe8cbf6dc0bdc77970c10d676ea64628b2334dbd8dbb3bc56d11de46d3d5531b10c1a459aa0dd398479111fb67e84d15584fb17ac3ca08c728362e69a4e53434d0a5b8da419d93561;
    5'b01101 : xpb = 1024'h98edff65e598920682272ad9ea55b3bb1c3d2ff2332404b82a58c9c48dfd766ee750c554efbaf421a0db0d92d92409ec562d6efba2da35408aea3b60e715b5f26c18d764b738d531d25b6e63256a5c62218b76edb8d224413192d791bdc88bdbb1bdd933d7cb4cd31b4aace280ff45ff7f92a1ba0635d0acd11723b22768d7b2;
    5'b01110 : xpb = 1024'h19b7094ba65f6615a9b495f3c08f5e0c95ece3a36f370f5920a06d356222e976c3b7462202fa5c7f2bc4a5cb5813643b1a2a175a30adb897c694087877c7f9c57d1a3a3d47c4a936ee7fe4ad645383c7df40fd5a7c8e9c0a17ed78e20893ba0bb6300878048cfc32ada5b39cd8dd9632ce87df76dcd00dc51633ebbac161398;
    5'b01111 : xpb = 1024'h1af6271951218f84fe14dfbb9e167f57e7f66fb3103a7daa7797fd37d14993c7f46ea0e81acad5fce3fbc66d753c73657131fbd5c5ee521e1e87850c62b5bdf7b7d9a491a150bd3a1e0e90d51ffbd847ce61a2562345dc50c6f769853d748df7f40fba04d98f4b40c129f07011ec92f02918391725af8e3c181ed4c9b9a5b5e9;
    5'b10000 : xpb = 1024'h3450dd9de7dd28a8a18e7618002408cf068e112be9818a5f5d25f39c4c70f8f87ca1cd6e15660631d53b427e34f7b08730c15635e8d1c8b2c0a5c9913deefc5317e1a57f6e252fe0cd35235f69b278531ecf34d69ec2cee0ec6ffb7c5a5fe04f2cbc738232d5c6be577985a6564b4c7d2547f436dd921b9bdeda6ad7c735583a;
    5'b10001 : xpb = 1024'h4dab94227e98c1cc45080c74623192462525b2a4c2c8971442b3ea00c7985e2904d4f9f410013666c67abe8ef4b2eda8f050b0960bb53f4762c40e1619283aae77e9a66d3af9a2877c5bb5e9b369185e6f3cc7571a3fc17111e88d73774b32a665692cff8c1c423bedc91adc9aaa060a2177af569574a8fba59600e5d4c4fa8b;
    5'b10010 : xpb = 1024'h67064aa715545aefe881a2d0c43f1bbd43bd541d9c0fa3c92841e06542bfc3598d08267a0a9c669bb7ba3a9fb46e2acaafe00af62e98b5dc04e2529af4617909d7f1a75b07ce152e2b824873fd1fb869bfaa59d795bcb40137611f6a943684fd9e15e67ce562bdb98418b012df08bf971da76a764d57365b6c5196f3e2549cdc;
    5'b10011 : xpb = 1024'h8061012bac0ff4138bfb392d264ca5346254f5967556b07e0dcfd6c9bde7288a153b5300053796d0a8f9b6b0742967ec6f6f6556517c2c70a700971fcf9ab76537f9a848d4a287d4daa8dafe46d658751017ec581139a6915cd9b161b121d754d6c29ffa3ea939371a6845492367792419d725960539c3bb330d2d01efe43f2d;
    5'b10100 : xpb = 1024'h99bbb7b042cb8d372f74cf89885a2eab80ec970f4e9dbd32f35dcd2e390e8dba9d6e7f85ffd2c7059a3932c133e4a50e2efebfb6745fa305491edba4aad3f5c09801a936a176fa7b89cf6d88908cf88060857ed88cb6992182524358ce0d29ac0f6f597797efb4b4b0b7da7f67c632b11606e0b5bd1c511af9c8c30ffd73e17e;
    5'b10101 : xpb = 1024'h26928df1798f19207e8ee0eda0d70d12e0e3557526d29705b0f0a3d013345e322592e93304778abec1a6f8b1041d1658a73f2307490494e3a9de0cb4b3abf6a83ba7575beba6fdd265bfd704167d45abcee17c07bad5ea0f23e435530cdd971191480cb406d37a4c04788d6b454c614c35cbcf324b3814a7a14de1982211d64;
    5'b10110 : xpb = 1024'h1bc3df63ae548ab5ab62846b3c1afa484ca5d6d02bb43625409d00a17c5aab13aa8c5b192ae2a8e0dd59eb9bcffd0e874a034c909773bfe2dcbc25502673fdc5e3c276638b8ee283d5828ffa8b1e74660d5baa40f72a513117b6d54c4db92bc851c13a4899b3b32256971e0cf8b37fa1bf8c7812dc960eaa40d074278fb0bfb5;
    5'b10111 : xpb = 1024'h351e95e8451023d94edc1ac79e2883bf6b3d784904fb42da262af705f782104432bf879f257dd915ce9967ac8fb84ba90992a6f0ba5736777eda69d501ad3c2143ca77515863552a84a92284d4d514715dc93cc172a743c13d2f67436aa47e1f8a6df3c5f2fa2e9fece6b3433d12392ebbbc333294789c0a078c0a359d406206;
    5'b11000 : xpb = 1024'h4e794c6cdbcbbcfcf255b12400360d3689d519c1de424f8f0bb8ed6a72a97574baf2b4252019094abfd8e3bd4f7388cac9220150dd3aad0c20f8ae59dce67a7ca3d2783f2537c7d133cfb50f1e8bb47cae36cf41ee24365162a7f93a878fd076c31aad434c40aa1d833648798170f2bbb7ebee524c5b2969ce47a043aad00457;
    5'b11001 : xpb = 1024'h67d402f17287562095cf4780624396ada86cbb3ab7895c43f146e3ceedd0daa54325e0ab1ab4397fb1185fce0f2ec5ec88b15bb1001e23a0c316f2deb81fb8d803da792cf20c3a77e2f6479968425487fea461c269a128e188208b31a47b22cdfbc766c0a587259b1985ddafc5cfac48b41ba972043db6c995033651b85fa6a8;
    5'b11010 : xpb = 1024'h812eb9760942ef443948dddcc4512024c7045cb390d068f8d6d4da3368f83fd5cb590d31154f69b4a257dbdeceea030e4840b61123019a35653537639358f73363e27a1abee0ad1e921cda23b1f8f4934f11f442e51e1b71ad991d28c16675253474203dfecda118afd572e60a2e65d5b04b6491bc2044295bbecc5fc5ef48f9;
    5'b11011 : xpb = 1024'h9a896ffa9ffe8867dcc27439265ea99be59bfe2c6a1775adbc62d097e41fa506538c39b70fea99e9939757ef8ea5403007d0107145e510ca07537be86e92358ec3ea7b088bb51fc541436cadfbaf949e9f7f86c3609b0e01d311af1fde51c77c6d20d9bb58141c964625081c4e8d1f62ac7b1fb17402d189227a626dd37eeb4a;
    5'b11100 : xpb = 1024'h336e12974cbecc2b53692be7811ebc192bd9c746de6e1eb24140da6ac445d2ed876e8c4405f4b8fe57894b96b026c87634542eb4615b712f8d2810f0ef8ff38afa34747a8f89526ddcffc95ac8a7078fbe81fab4f91d38142fdaf1c4112774176c6010f00919f8655b4b6739b1bb2c659d0fbeedb9a01b8a2c67d77582c2730;
    5'b11101 : xpb = 1024'h1c9197ae0b8785e658b0291ada1f7538b1553ded472deea009a2040b276bc25f60aa154a3afa7bc4d6b810ca2abda9a922d49d4b68f92da79af0c593ea323d940fab483575cd07cd8cf68f1ff64110844c55b22bcb0ec611687641135dfdc998af72ba8c59d81b03ec044ba9df7a6c535600b70e937c8f186982138565bbc981;
    5'b11110 : xpb = 1024'h35ec4e32a2431f09fc29bf773c2cfeafcfecdf662074fb54ef2ffa6fa293278fe8dd41d03595abf9c7f78cdaea78e6cae263f7ab8bdca43c3d0f0a18c56b7bef6fb3492342a17a743c1d21aa3ff7b08f9cc344ac468bb8a18deed30a7ae91befe81f7409b31e96818253e0e023d925e05230722e4b5f1c78303da993734b6bd2;
    5'b11111 : xpb = 1024'h4f4704b738feb82d9fa355d39e3a8826ee8480def9bc0809d4bdf0d41dba8cc071106e563030dc2eb93708ebaa3423eca1f3520baec01ad0df2d4e9da0a4ba4acfbb4a110f75ed1aeb43b43489ae509aed30d72cc208ab31b367650197d46e4720cc2d870c6511ff18a376166837df6d4e602d4e0341a9d7f6f93fa180db0e23;
    endcase
end

endmodule

module xpb_5_830
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h9eb4b6a138236332dec7c8a9ea01f62bee99423a5905e5be2dd4a67b50079b3d97f95525ad20b3078129a7210ac4954d7f94ce87c3ea210efdf19978c4705320fbb857489e7c5ab5dfdd0ced038c0e7046d6812fa8b12df989800a5d749b74b52f2a187b49bfc5d1ede72438d94b56bace8e3976966520a39ccc9aade4d1366c;
    5'b00010 : xpb = 1024'h8cbc27ecae58919cf28a197cc3a9a5066bbc8143dc942b04ddcc93a0ed0c89732caa2cd2901ae78062f50efb322b19d09b0f7529652171d24b43f3934e0e3190832179e28d67b826ad2017376e3c58af99a808c6c4dc2ee25d7382c02f0c46d82f4c9ecce2b69316550e6192bac6874c4e42940adc7ee416f329ba5740c0066d;
    5'b00011 : xpb = 1024'h7ac39938248dc007064c6a4f9d5153e0e8dfc04d6022704b8dc480c68a1177a8c15b047f73151bf944c076d559919e53b68a1bcb0658c29598964dadd7ac10000a8a9c7c7c5315977a632181d8eca2eeec79905de1072fcb3166fb22e97d18fb2f6f251e7bad605abc359eec9c41b7ddcdf6ee9f2298a78a4986da009caed66e;
    5'b00100 : xpb = 1024'h68cb0a839ac2ee711a0ebb2276f902bb6602ff56e3b0b5923dbc6dec271665de560bdc2c560f5072268bdeaf80f822d6d204c26ca7901358e5e8a7c86149ee6f91f3bf166b3e730847a62bcc439ced2e3f4b17f4fd3230b4055a7385a3edeb1e2f91ab7014a42d9f235cdc467dbce86f4dab493368b26afd9fe3f9a9f89da66f;
    5'b00101 : xpb = 1024'h56d27bcf10f81cdb2dd10bf550a0b195e3263e60673efad8edb45b11c41b5413eabcb3d9390984eb08574689a85ea759ed7f690e48c7641c333b01e2eae7ccdf195ce1b05a29d07914e93616ae4d376d921c9f8c195d319cd94debe85e5ebd412fb431c1ad9afae38a8419a05f381900cd5fa3c7aecc2e70f6411953548c7670;
    5'b00110 : xpb = 1024'h44d9ed1a872d4b4541935cc82a48607060497d69eacd401f9dac4837612042497f6d8b861c03b963ea22ae63cfc52bdd08fa0fafe9feb4df808d5bfd7485ab4ea0c6044a49152de9e22c406118fd81ace4ee272335883285ad41644b18cf8f642fd6b8134691c827f1ab56fa40b349924d13fe5bf4e5f1e44c9e38fcb07b4671;
    5'b00111 : xpb = 1024'h32e15e65fd6279af5555ad9b03f00f4add6cbc736e5b85664da4355cfe25307f141e6332fefdeddccbee163df72bb0602474b6518b3605a2cddfb617fe2389be282f26e438008b5aaf6f4aab83adcbec37bfaeba51b3336e8134dcadd34061872ff93e64df88956c58d29454222e7a23ccc858f03affb557a2fb58a60c6a1672;
    5'b01000 : xpb = 1024'h20e8cfb17397a8196917fe6ddd97be255a8ffb7cf1e9caacfd9c22829b2a1eb4a8cf3adfe1f82255adb97e181e9234e33fef5cf32c6d56661b32103287c1682daf98497e26ebe8cb7cb254f5ee5e162b8a9136516dde3457552855108db133aa301bc4b6787f62b0bff9d1ae03a9aab54c7cb384811978caf958784f6858e673;
    5'b01001 : xpb = 1024'hef040fce9ccd6837cda4f40b73f6cffd7b33a8675780ff3ad940fa8382f0cea3d80128cc4f256ce8f84e5f245f8b9665b6a0394cda4a72968846a4d115f469d37016c1815d7463c49f55f40590e606add62bde88a093540291bcd73482205cd303e4b0811762ff527210f07e524db46cc310e18c7333c3e4fb597f8c447b674;
    5'b01010 : xpb = 1024'hada4f79e21f039b65ba217eaa141632bc64c7cc0ce7df5b1db68b6238836a827d57967b2721309d610ae8d1350bd4eb3dafed21c918ec838667603c5d5cf99be32b9c360b453a0f229d26c2d5c9a6edb24393f1832ba6339b29bd7d0bcbd7a825f6863835b35f5c715083340be7032019abf478f5d985ce1ec8232a6a918ece0;
    5'b01011 : xpb = 1024'h9bac68e9982568206f6468bd7ae91206436fbbca520c3af88b60a349253b965d6a2a3f5f550d3e4ef279f4ed7823d336f67978be32c618fbb3c85de05f6d782dba22e5faa33efe62f7157677c74ab91a770ac6af4ee56422868f5033772e4ca55f8ae9d4f42cc30b7c2f709a9feb62931a73a223a3b2205542df52500507bce1;
    5'b01100 : xpb = 1024'h89b3da350e5a968a8326b9905490c0e0c092fad3d59a803f3b58906ec2408492fedb170c380772c7d4455cc79f8a57ba11f41f5fd3fd69bf011ab7fae90b569d418c0894922a5bd3c45880c231fb0359c9dc4e466b10650b5a82c896319f1ec85fad70268d23904fe356adf4816693249a27fcb7e9cbe3c8993c71f960f68ce2;
    5'b01101 : xpb = 1024'h77bb4b80848fc4f496e90a632e386fbb3db639dd5928c585eb507d945f4572c8938beeb91b01a740b610c4a1c6f0dc3d2d6ec6017534ba824e6d121572a9350cc8f52b2e8115b944919b8b0c9cab4d991cadd5dd873b65f42e7640f8ec0ff0eb5fcff678261a5d944a7deb4e62e1c3b619dc574c2fe5a73bef9991a2bce55ce3;
    5'b01110 : xpb = 1024'h65c2bccbfac4f35eaaab5b3607e01e95bad978e6dcb70acc9b486ab9fc4a60fe283cc665fdfbdbb997dc2c7bee5760c048e96ca3166c0b459bbf6c2ffc47137c505e4dc8700116b55ede9557075b97d86f7f5d74a36666dd0269b95ba680c30e5ff27cc9bf112ad8b1a528a8445cf4479990b1e075ff6aaf45f6b14c18d42ce4;
    5'b01111 : xpb = 1024'h53ca2e1770fa21c8be6dac08e187cd7037fcb7f0604550134b4057df994f4f33bced9e12e0f6103279a7945615bde54364641344b7a35c08e911c64a85e4f1ebd7c770625eec74262c219fa1720be217c250e50bbf9167c5d65d31be60f195316015031b5807f81d18cc660225d824d919450c74bc192e229c53d0f574c2fce5;
    5'b10000 : xpb = 1024'h41d19f62e72f5032d22ffcdbbb2f7c4ab51ff6f9e3d39559fb38450536543d69519e75bfc3f044ab5b72fc303d2469c67fdeb9e658daaccc366420650f82d05b5f3092fc4dd7d196f964a9ebdcbc2c5715226ca2dbbc68aeaa50aa211b6267546037896cf0fec5617ff3a35c0753556a98f967090232f195f2b0f09ed0b1cce6;
    5'b10001 : xpb = 1024'h2fd910ae5d647e9ce5f24dae94d72b25324336036761daa0ab30322ad3592b9ee64f4d6ca6ea79243d3e640a648aee499b596087fa11fd8f83b67a7f9920aecae699b5963cc32f07c6a7b436476c769667f3f439f7e769977e442283d5d33977605a0fbe89f592a5e71ae0b5e8ce85fc18adc19d484cb509490e10482ca09ce7;
    5'b10010 : xpb = 1024'h1de081f9d399ad06f9b49e816e7ed9ffaf66750ceaf01fe75b281f50705e19d47b00251989e4ad9d1f09cbe48bf172ccb6d407299b494e52d108d49a22be8d3a6e02d8302bae8c7893eabe80b21cc0d5bac57bd114126a8052379ae690440b9a607c961022ec5fea4e421e0fca49b68d98621c318e66787c9f6b2ff1888f6ce8;
    5'b10011 : xpb = 1024'hbe7f34549cedb710d76ef54482688da2c89b4166e7e652e0b200c760d63080a0fb0fcc66cdee21600d533beb357f74fd24eadcb3c809f161e5b2eb4ac5c6ba9f56bfaca1a99e9e9612dc8cb1ccd0b150d970368303d6b69262b13494ab4ddbd609f1c61bbe32d2eb5695b69abc4e71f181676c5d4803beff5c84f9ae47e3ce9;
    5'b10100 : xpb = 1024'haa9ca9e681f23ea3ec3eb7fe32287f061b22f650c7844aec38f4b2f15d6aa347a7aa51ec19ff951d81fedadfbe1c8c9d51e37c53006ac0251c4cc82d70ccbecaf1245212b916449f410ad5b820591985546d8497d8ee9962afab1da6bf5052728fc934dd05a2f300a3507fa285103dd9e6a4b03c6ae55c939294ea48c94f7355;
    5'b10101 : xpb = 1024'h98a41b31f8276d0e000108d10bd02de09846355a4b129032e8eca016fa6f917d3c5b2998fcf9c99663ca42b9e58311206d5e22f4a1a210e8699f2247fa6a9d3a788d74aca801a2100e4de0028b0963c4a73f0c2ef5199a4b839e960979c124958febbb2e9e99c0450a77bcfc668b6e6b66590ad0b0ff2006e8f209f2253e4356;
    5'b10110 : xpb = 1024'h86ab8c7d6e5c9b7813c359a3e577dcbb15697463cea0d57998e48d3c97747fb2d10c0145dff3fe0f4595aa940ce995a388d8c99642d961abb6f17c6284087ba9fff6974696ecff80db90ea4cf5b9ae03fa1093c611449b3457920e6c3431f6b8900e418037908d89719efa5648069efce60d6564f718e37a3f4f299b812d1357;
    5'b10111 : xpb = 1024'h74b2fdc8e491c9e22785aa76bf1f8b95928cb36d522f1ac048dc7a6234796de865bcd8f2c2ee32882761126e34501a26a4537037e410b26f0443d67d0da65a19875fb9e085d85cf1a8d3f4976069f8434ce21b5d2d6f9c1d2b8586ceeea2c8db9030c7d1d0875acdd8c637b02981cf8e65c1bff93d32a6ed95ac4944dd1be358;
    5'b11000 : xpb = 1024'h62ba6f145ac6f84c3b47fb4998c73a700faff276d5bd6006f8d46787d17e5c1dfa6db09fa5e86701092c7a485bb69ea9bfce16d98548033251963097974438890ec8dc7a74c3ba627616fee1cb1a42829fb3a2f4499a9d05ff78ff31a9139afe90534e23697e28123fed750a0afd001fe5761a8d834c6a60ec0968ee390ab359;
    5'b11001 : xpb = 1024'h50c1e05fd0fc26b64f0a4c1c726ee94a8cd33180594ba54da8cc54ad6e834a538f1e884c88e29b79eaf7e222831d232cdb48bd7b267f53f59ee88ab220e216f89631ff1463af17d3435a092c35ca8cc1f2852a8b65c59deed36c779463846d219075d4750274f556a714b263ec7830b1652a7521c9662dd44266889794f9835a;
    5'b11010 : xpb = 1024'h3ec951ab4731552062cc9cef4c16982509f67089dcd9ea9458c441d30b88388923cf5ff96bdccff2ccc349fcaa83a7aff6c3641cc7b6a4b8ec3ae4ccaa7ff5681d9b21ae529a7544109d1376a07ad7014556b22281f09ed7a75feff71df53f4490985ac69b6bc29b0e3befbdcdf36142e4decfb60f7ff14798c3a840f0e8535b;
    5'b11011 : xpb = 1024'h2cd0c2f6bd66838a768eedc225be46ff8719af9360682fdb08bc2ef8a88d26beb88037a64ed7046bae8eb1d6d1ea2c33123e0abe68edf57c398d3ee7341dd3d7a50444484185d2b4dde01dc10b2b2140982839b99e1b9fc07b536859d866116790bae11834628fdf75632d17af6e91d464932a4a5599b4baef20c7ea4cd7235c;
    5'b11100 : xpb = 1024'h1ad83442339bb1f48a513e94ff65f5da043cee9ce3f67521b8b41c1e459214f44d310f5331d138e4905a19b0f950b0b62db8b1600a25463f86df9901bdbbb2472c6d66e230713025ab23280b75db6b7feaf9c150ba46a0a94f46e0bc92d6e38a90dd6769cd595d23dc8a6a7190e9c265e44784de9bb3782e457de793a8c5f35d;
    5'b11101 : xpb = 1024'h8dfa58da9d0e05e9e138f67d90da4b481602da66784ba6868ac0943e2970329e1e1e70014cb6d5d7225818b20b7353949335801ab5c9702d431f31c475990b6b3d6897c1f5c8d9678663255e08bb5bf3dcb48e7d671a192233a591f4d47b5ad90ffedbb66502a6843b1a7cb7264f2f763fbdf72e1cd3ba19bdb073d04b4c35e;
    5'b11110 : xpb = 1024'ha7945c2ee1f443917cdb5811c30f9ae06ff96fe0c08aa0269680afbf329e9e6779db3c25c1ec2064f34f28ac2b7bca86c8c826896f46b811d2238c950bc9e3d7af8ee0c4bdd8e84c58433f42e417c42f84a1ca177f22cf8bacba637cc1e32a62c02a0636b00ff03a3198cc044bb049b2328a18e978325c4538a7a1eae985f9ca;
    5'b11111 : xpb = 1024'h959bcd7a582971fb909da8e49cb749baed1caeea4418e56d46789ce4cfa38c9d0e8c13d2a4e654ddd51a908652e24f09e442cd2b107e08d51f75e6af9567c24736f8035eacc445bd2586498d4ec80e6ed77351ae9b4dd07480addbdf7c53fc85c04c8c884906bd7e98c0095e2d2b7a43b23e737dbe4c1fb88f04c1944574c9cb;
    endcase
end

endmodule

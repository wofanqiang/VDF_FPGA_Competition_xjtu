`timescale 1ns/1ns
/*******************************************************************************
    Institute:   Xi'an Jiaotong University
    Department:  Microelectronic
    Author :     Li Xiaocong

    Unless you get the permission of the Author, you can't modify,
    distribute or use for commercial purposes.
*******************************************************************************/
module msq_product_period4
(
	input wire [1023:0] al,
	input wire [1:0] sel,
	output wire [127:0] col_0,
	output wire [127:0] col_1,
	output wire [127:0] col_2,
	output wire [127:0] col_3,
	output wire [127:0] col_4,
	output wire [127:0] col_5,
	output wire [127:0] col_6,
	output wire [127:0] col_7,
	output wire [127:0] col_8,
	output wire [127:0] col_9,
	output wire [127:0] col_10,
	output wire [127:0] col_11,
	output wire [127:0] col_12,
	output wire [127:0] col_13,
	output wire [127:0] col_14,
	output wire [127:0] col_15,
	output wire [127:0] col_16,
	output wire [127:0] col_17,
	output wire [127:0] col_18,
	output wire [127:0] col_19,
	output wire [127:0] col_20,
	output wire [127:0] col_21,
	output wire [127:0] col_22,
	output wire [127:0] col_23,
	output wire [127:0] col_24,
	output wire [127:0] col_25,
	output wire [127:0] col_26,
	output wire [127:0] col_27,
	output wire [127:0] col_28,
	output wire [127:0] col_29,
	output wire [127:0] col_30,
	output wire [127:0] col_31,
	output wire [127:0] col_32,
	output wire [127:0] col_33,
	output wire [127:0] col_34,
	output wire [127:0] col_35,
	output wire [127:0] col_36,
	output wire [127:0] col_37,
	output wire [127:0] col_38,
	output wire [127:0] col_39,
	output wire [127:0] col_40,
	output wire [127:0] col_41,
	output wire [127:0] col_42,
	output wire [127:0] col_43,
	output wire [127:0] col_44,
	output wire [127:0] col_45,
	output wire [127:0] col_46,
	output wire [127:0] col_47,
	output wire [127:0] col_48,
	output wire [127:0] col_49,
	output wire [127:0] col_50,
	output wire [127:0] col_51,
	output wire [127:0] col_52,
	output wire [127:0] col_53,
	output wire [127:0] col_54,
	output wire [127:0] col_55,
	output wire [127:0] col_56,
	output wire [127:0] col_57,
	output wire [127:0] col_58,
	output wire [127:0] col_59,
	output wire [127:0] col_60,
	output wire [127:0] col_61,
	output wire [127:0] col_62,
	output wire [127:0] col_63,
	output wire [127:0] col_64,
	output wire [127:0] col_65,
	output wire [127:0] col_66,
	output wire [127:0] col_67,
	output wire [127:0] col_68,
	output wire [127:0] col_69,
	output wire [127:0] col_70,
	output wire [127:0] col_71,
	output wire [127:0] col_72,
	output wire [127:0] col_73,
	output wire [127:0] col_74,
	output wire [127:0] col_75,
	output wire [127:0] col_76,
	output wire [127:0] col_77,
	output wire [127:0] col_78,
	output wire [127:0] col_79,
	output wire [127:0] col_80,
	output wire [127:0] col_81,
	output wire [127:0] col_82,
	output wire [127:0] col_83,
	output wire [127:0] col_84,
	output wire [127:0] col_85,
	output wire [127:0] col_86,
	output wire [127:0] col_87,
	output wire [127:0] col_88,
	output wire [127:0] col_89,
	output wire [127:0] col_90,
	output wire [127:0] col_91,
	output wire [127:0] col_92,
	output wire [127:0] col_93,
	output wire [127:0] col_94,
	output wire [127:0] col_95,
	output wire [127:0] col_96,
	output wire [127:0] col_97,
	output wire [127:0] col_98,
	output wire [127:0] col_99,
	output wire [127:0] col_100,
	output wire [127:0] col_101,
	output wire [127:0] col_102,
	output wire [127:0] col_103,
	output wire [127:0] col_104,
	output wire [127:0] col_105,
	output wire [127:0] col_106,
	output wire [127:0] col_107,
	output wire [127:0] col_108,
	output wire [127:0] col_109,
	output wire [127:0] col_110,
	output wire [127:0] col_111,
	output wire [127:0] col_112,
	output wire [127:0] col_113,
	output wire [127:0] col_114,
	output wire [127:0] col_115,
	output wire [127:0] col_116,
	output wire [127:0] col_117,
	output wire [127:0] col_118,
	output wire [127:0] col_119,
	output wire [127:0] col_120,
	output wire [127:0] col_121,
	output wire [127:0] col_122,
	output wire [127:0] col_123,
	output wire [127:0] col_124,
	output wire [127:0] col_125,
	output wire [127:0] col_126,
	output wire [127:0] col_127,
	output wire [127:0] col_128,
	output wire [127:0] col_129,
	output wire [127:0] col_130,
	output wire [127:0] col_131,
	output wire [127:0] col_132,
	output wire [127:0] col_133,
	output wire [127:0] col_134,
	output wire [127:0] col_135,
	output wire [127:0] col_136,
	output wire [127:0] col_137,
	output wire [127:0] col_138,
	output wire [127:0] col_139,
	output wire [127:0] col_140,
	output wire [127:0] col_141,
	output wire [127:0] col_142,
	output wire [127:0] col_143,
	output wire [127:0] col_144,
	output wire [127:0] col_145,
	output wire [127:0] col_146,
	output wire [127:0] col_147,
	output wire [127:0] col_148,
	output wire [127:0] col_149,
	output wire [127:0] col_150,
	output wire [127:0] col_151,
	output wire [127:0] col_152,
	output wire [127:0] col_153,
	output wire [127:0] col_154,
	output wire [127:0] col_155,
	output wire [127:0] col_156,
	output wire [127:0] col_157,
	output wire [127:0] col_158,
	output wire [127:0] col_159,
	output wire [127:0] col_160,
	output wire [127:0] col_161,
	output wire [127:0] col_162,
	output wire [127:0] col_163,
	output wire [127:0] col_164,
	output wire [127:0] col_165,
	output wire [127:0] col_166,
	output wire [127:0] col_167,
	output wire [127:0] col_168,
	output wire [127:0] col_169,
	output wire [127:0] col_170,
	output wire [127:0] col_171,
	output wire [127:0] col_172,
	output wire [127:0] col_173,
	output wire [127:0] col_174,
	output wire [127:0] col_175,
	output wire [127:0] col_176,
	output wire [127:0] col_177,
	output wire [127:0] col_178,
	output wire [127:0] col_179,
	output wire [127:0] col_180,
	output wire [127:0] col_181,
	output wire [127:0] col_182,
	output wire [127:0] col_183,
	output wire [127:0] col_184,
	output wire [127:0] col_185,
	output wire [127:0] col_186,
	output wire [127:0] col_187,
	output wire [127:0] col_188,
	output wire [127:0] col_189,
	output wire [127:0] col_190,
	output wire [127:0] col_191,
	output wire [127:0] col_192,
	output wire [127:0] col_193,
	output wire [127:0] col_194,
	output wire [127:0] col_195,
	output wire [127:0] col_196,
	output wire [127:0] col_197,
	output wire [127:0] col_198,
	output wire [127:0] col_199,
	output wire [127:0] col_200,
	output wire [127:0] col_201,
	output wire [127:0] col_202,
	output wire [127:0] col_203,
	output wire [127:0] col_204,
	output wire [127:0] col_205,
	output wire [127:0] col_206,
	output wire [127:0] col_207,
	output wire [127:0] col_208,
	output wire [127:0] col_209,
	output wire [127:0] col_210,
	output wire [127:0] col_211,
	output wire [127:0] col_212,
	output wire [127:0] col_213,
	output wire [127:0] col_214,
	output wire [127:0] col_215,
	output wire [127:0] col_216,
	output wire [127:0] col_217,
	output wire [127:0] col_218,
	output wire [127:0] col_219,
	output wire [127:0] col_220,
	output wire [127:0] col_221,
	output wire [127:0] col_222,
	output wire [127:0] col_223,
	output wire [127:0] col_224,
	output wire [127:0] col_225,
	output wire [127:0] col_226,
	output wire [127:0] col_227,
	output wire [127:0] col_228,
	output wire [127:0] col_229,
	output wire [127:0] col_230,
	output wire [127:0] col_231,
	output wire [127:0] col_232,
	output wire [127:0] col_233,
	output wire [127:0] col_234,
	output wire [127:0] col_235,
	output wire [127:0] col_236,
	output wire [127:0] col_237,
	output wire [127:0] col_238,
	output wire [127:0] col_239,
	output wire [127:0] col_240,
	output wire [127:0] col_241,
	output wire [127:0] col_242,
	output wire [127:0] col_243,
	output wire [127:0] col_244,
	output wire [127:0] col_245,
	output wire [127:0] col_246,
	output wire [127:0] col_247,
	output wire [127:0] col_248,
	output wire [127:0] col_249,
	output wire [127:0] col_250,
	output wire [127:0] col_251,
	output wire [127:0] col_252,
	output wire [127:0] col_253,
	output wire [127:0] col_254,
	output wire [127:0] col_255,
	output wire [127:0] col_256,
	output wire [127:0] col_257,
	output wire [127:0] col_258,
	output wire [127:0] col_259,
	output wire [127:0] col_260,
	output wire [127:0] col_261,
	output wire [127:0] col_262,
	output wire [127:0] col_263,
	output wire [127:0] col_264,
	output wire [127:0] col_265,
	output wire [127:0] col_266,
	output wire [127:0] col_267,
	output wire [127:0] col_268,
	output wire [127:0] col_269,
	output wire [127:0] col_270,
	output wire [127:0] col_271,
	output wire [127:0] col_272,
	output wire [127:0] col_273,
	output wire [127:0] col_274,
	output wire [127:0] col_275,
	output wire [127:0] col_276,
	output wire [127:0] col_277,
	output wire [127:0] col_278,
	output wire [127:0] col_279,
	output wire [127:0] col_280,
	output wire [127:0] col_281,
	output wire [127:0] col_282,
	output wire [127:0] col_283,
	output wire [127:0] col_284,
	output wire [127:0] col_285,
	output wire [127:0] col_286,
	output wire [127:0] col_287,
	output wire [127:0] col_288,
	output wire [127:0] col_289,
	output wire [127:0] col_290,
	output wire [127:0] col_291,
	output wire [127:0] col_292,
	output wire [127:0] col_293,
	output wire [127:0] col_294,
	output wire [127:0] col_295,
	output wire [127:0] col_296,
	output wire [127:0] col_297,
	output wire [127:0] col_298,
	output wire [127:0] col_299,
	output wire [127:0] col_300,
	output wire [127:0] col_301,
	output wire [127:0] col_302,
	output wire [127:0] col_303,
	output wire [127:0] col_304,
	output wire [127:0] col_305,
	output wire [127:0] col_306,
	output wire [127:0] col_307,
	output wire [127:0] col_308,
	output wire [127:0] col_309,
	output wire [127:0] col_310,
	output wire [127:0] col_311,
	output wire [127:0] col_312,
	output wire [127:0] col_313,
	output wire [127:0] col_314,
	output wire [127:0] col_315,
	output wire [127:0] col_316,
	output wire [127:0] col_317,
	output wire [127:0] col_318,
	output wire [127:0] col_319,
	output wire [127:0] col_320,
	output wire [127:0] col_321,
	output wire [127:0] col_322,
	output wire [127:0] col_323,
	output wire [127:0] col_324,
	output wire [127:0] col_325,
	output wire [127:0] col_326,
	output wire [127:0] col_327,
	output wire [127:0] col_328,
	output wire [127:0] col_329,
	output wire [127:0] col_330,
	output wire [127:0] col_331,
	output wire [127:0] col_332,
	output wire [127:0] col_333,
	output wire [127:0] col_334,
	output wire [127:0] col_335,
	output wire [127:0] col_336,
	output wire [127:0] col_337,
	output wire [127:0] col_338,
	output wire [127:0] col_339,
	output wire [127:0] col_340,
	output wire [127:0] col_341,
	output wire [127:0] col_342,
	output wire [127:0] col_343,
	output wire [127:0] col_344,
	output wire [127:0] col_345,
	output wire [127:0] col_346,
	output wire [127:0] col_347,
	output wire [127:0] col_348,
	output wire [127:0] col_349,
	output wire [127:0] col_350,
	output wire [127:0] col_351,
	output wire [127:0] col_352,
	output wire [127:0] col_353,
	output wire [127:0] col_354,
	output wire [127:0] col_355,
	output wire [127:0] col_356,
	output wire [127:0] col_357,
	output wire [127:0] col_358,
	output wire [127:0] col_359,
	output wire [127:0] col_360,
	output wire [127:0] col_361,
	output wire [127:0] col_362,
	output wire [127:0] col_363,
	output wire [127:0] col_364,
	output wire [127:0] col_365,
	output wire [127:0] col_366,
	output wire [127:0] col_367,
	output wire [127:0] col_368,
	output wire [127:0] col_369,
	output wire [127:0] col_370,
	output wire [127:0] col_371,
	output wire [127:0] col_372,
	output wire [127:0] col_373,
	output wire [127:0] col_374,
	output wire [127:0] col_375,
	output wire [127:0] col_376,
	output wire [127:0] col_377,
	output wire [127:0] col_378,
	output wire [127:0] col_379,
	output wire [127:0] col_380,
	output wire [127:0] col_381,
	output wire [127:0] col_382,
	output wire [127:0] col_383,
	output wire [127:0] col_384,
	output wire [127:0] col_385,
	output wire [127:0] col_386,
	output wire [127:0] col_387,
	output wire [127:0] col_388,
	output wire [127:0] col_389,
	output wire [127:0] col_390,
	output wire [127:0] col_391,
	output wire [127:0] col_392,
	output wire [127:0] col_393,
	output wire [127:0] col_394,
	output wire [127:0] col_395,
	output wire [127:0] col_396,
	output wire [127:0] col_397,
	output wire [127:0] col_398,
	output wire [127:0] col_399,
	output wire [127:0] col_400,
	output wire [127:0] col_401,
	output wire [127:0] col_402,
	output wire [127:0] col_403,
	output wire [127:0] col_404,
	output wire [127:0] col_405,
	output wire [127:0] col_406,
	output wire [127:0] col_407,
	output wire [127:0] col_408,
	output wire [127:0] col_409,
	output wire [127:0] col_410,
	output wire [127:0] col_411,
	output wire [127:0] col_412,
	output wire [127:0] col_413,
	output wire [127:0] col_414,
	output wire [127:0] col_415,
	output wire [127:0] col_416,
	output wire [127:0] col_417,
	output wire [127:0] col_418,
	output wire [127:0] col_419,
	output wire [127:0] col_420,
	output wire [127:0] col_421,
	output wire [127:0] col_422,
	output wire [127:0] col_423,
	output wire [127:0] col_424,
	output wire [127:0] col_425,
	output wire [127:0] col_426,
	output wire [127:0] col_427,
	output wire [127:0] col_428,
	output wire [127:0] col_429,
	output wire [127:0] col_430,
	output wire [127:0] col_431,
	output wire [127:0] col_432,
	output wire [127:0] col_433,
	output wire [127:0] col_434,
	output wire [127:0] col_435,
	output wire [127:0] col_436,
	output wire [127:0] col_437,
	output wire [127:0] col_438,
	output wire [127:0] col_439,
	output wire [127:0] col_440,
	output wire [127:0] col_441,
	output wire [127:0] col_442,
	output wire [127:0] col_443,
	output wire [127:0] col_444,
	output wire [127:0] col_445,
	output wire [127:0] col_446,
	output wire [127:0] col_447,
	output wire [127:0] col_448,
	output wire [127:0] col_449,
	output wire [127:0] col_450,
	output wire [127:0] col_451,
	output wire [127:0] col_452,
	output wire [127:0] col_453,
	output wire [127:0] col_454,
	output wire [127:0] col_455,
	output wire [127:0] col_456,
	output wire [127:0] col_457,
	output wire [127:0] col_458,
	output wire [127:0] col_459,
	output wire [127:0] col_460,
	output wire [127:0] col_461,
	output wire [127:0] col_462,
	output wire [127:0] col_463,
	output wire [127:0] col_464,
	output wire [127:0] col_465,
	output wire [127:0] col_466,
	output wire [127:0] col_467,
	output wire [127:0] col_468,
	output wire [127:0] col_469,
	output wire [127:0] col_470,
	output wire [127:0] col_471,
	output wire [127:0] col_472,
	output wire [127:0] col_473,
	output wire [127:0] col_474,
	output wire [127:0] col_475,
	output wire [127:0] col_476,
	output wire [127:0] col_477,
	output wire [127:0] col_478,
	output wire [127:0] col_479,
	output wire [127:0] col_480,
	output wire [127:0] col_481,
	output wire [127:0] col_482,
	output wire [127:0] col_483,
	output wire [127:0] col_484,
	output wire [127:0] col_485,
	output wire [127:0] col_486,
	output wire [127:0] col_487,
	output wire [127:0] col_488,
	output wire [127:0] col_489,
	output wire [127:0] col_490,
	output wire [127:0] col_491,
	output wire [127:0] col_492,
	output wire [127:0] col_493,
	output wire [127:0] col_494,
	output wire [127:0] col_495,
	output wire [127:0] col_496,
	output wire [127:0] col_497,
	output wire [127:0] col_498,
	output wire [127:0] col_499,
	output wire [127:0] col_500,
	output wire [127:0] col_501,
	output wire [127:0] col_502,
	output wire [127:0] col_503,
	output wire [127:0] col_504,
	output wire [127:0] col_505,
	output wire [127:0] col_506,
	output wire [127:0] col_507,
	output wire [127:0] col_508,
	output wire [127:0] col_509,
	output wire [127:0] col_510,
	output wire [127:0] col_511,
	output wire [127:0] col_512,
	output wire [127:0] col_513,
	output wire [127:0] col_514,
	output wire [127:0] col_515,
	output wire [127:0] col_516,
	output wire [127:0] col_517,
	output wire [127:0] col_518,
	output wire [127:0] col_519,
	output wire [127:0] col_520,
	output wire [127:0] col_521,
	output wire [127:0] col_522,
	output wire [127:0] col_523,
	output wire [127:0] col_524,
	output wire [127:0] col_525,
	output wire [127:0] col_526,
	output wire [127:0] col_527,
	output wire [127:0] col_528,
	output wire [127:0] col_529,
	output wire [127:0] col_530,
	output wire [127:0] col_531,
	output wire [127:0] col_532,
	output wire [127:0] col_533,
	output wire [127:0] col_534,
	output wire [127:0] col_535,
	output wire [127:0] col_536,
	output wire [127:0] col_537,
	output wire [127:0] col_538,
	output wire [127:0] col_539,
	output wire [127:0] col_540,
	output wire [127:0] col_541,
	output wire [127:0] col_542,
	output wire [127:0] col_543,
	output wire [127:0] col_544,
	output wire [127:0] col_545,
	output wire [127:0] col_546,
	output wire [127:0] col_547,
	output wire [127:0] col_548,
	output wire [127:0] col_549,
	output wire [127:0] col_550,
	output wire [127:0] col_551,
	output wire [127:0] col_552,
	output wire [127:0] col_553,
	output wire [127:0] col_554,
	output wire [127:0] col_555,
	output wire [127:0] col_556,
	output wire [127:0] col_557,
	output wire [127:0] col_558,
	output wire [127:0] col_559,
	output wire [127:0] col_560,
	output wire [127:0] col_561,
	output wire [127:0] col_562,
	output wire [127:0] col_563,
	output wire [127:0] col_564,
	output wire [127:0] col_565,
	output wire [127:0] col_566,
	output wire [127:0] col_567,
	output wire [127:0] col_568,
	output wire [127:0] col_569,
	output wire [127:0] col_570,
	output wire [127:0] col_571,
	output wire [127:0] col_572,
	output wire [127:0] col_573,
	output wire [127:0] col_574,
	output wire [127:0] col_575,
	output wire [127:0] col_576,
	output wire [127:0] col_577,
	output wire [127:0] col_578,
	output wire [127:0] col_579,
	output wire [127:0] col_580,
	output wire [127:0] col_581,
	output wire [127:0] col_582,
	output wire [127:0] col_583,
	output wire [127:0] col_584,
	output wire [127:0] col_585,
	output wire [127:0] col_586,
	output wire [127:0] col_587,
	output wire [127:0] col_588,
	output wire [127:0] col_589,
	output wire [127:0] col_590,
	output wire [127:0] col_591,
	output wire [127:0] col_592,
	output wire [127:0] col_593,
	output wire [127:0] col_594,
	output wire [127:0] col_595,
	output wire [127:0] col_596,
	output wire [127:0] col_597,
	output wire [127:0] col_598,
	output wire [127:0] col_599,
	output wire [127:0] col_600,
	output wire [127:0] col_601,
	output wire [127:0] col_602,
	output wire [127:0] col_603,
	output wire [127:0] col_604,
	output wire [127:0] col_605,
	output wire [127:0] col_606,
	output wire [127:0] col_607,
	output wire [127:0] col_608,
	output wire [127:0] col_609,
	output wire [127:0] col_610,
	output wire [127:0] col_611,
	output wire [127:0] col_612,
	output wire [127:0] col_613,
	output wire [127:0] col_614,
	output wire [127:0] col_615,
	output wire [127:0] col_616,
	output wire [127:0] col_617,
	output wire [127:0] col_618,
	output wire [127:0] col_619,
	output wire [127:0] col_620,
	output wire [127:0] col_621,
	output wire [127:0] col_622,
	output wire [127:0] col_623,
	output wire [127:0] col_624,
	output wire [127:0] col_625,
	output wire [127:0] col_626,
	output wire [127:0] col_627,
	output wire [127:0] col_628,
	output wire [127:0] col_629,
	output wire [127:0] col_630,
	output wire [127:0] col_631,
	output wire [127:0] col_632,
	output wire [127:0] col_633,
	output wire [127:0] col_634,
	output wire [127:0] col_635,
	output wire [127:0] col_636,
	output wire [127:0] col_637,
	output wire [127:0] col_638,
	output wire [127:0] col_639,
	output wire [127:0] col_640,
	output wire [127:0] col_641,
	output wire [127:0] col_642,
	output wire [127:0] col_643,
	output wire [127:0] col_644,
	output wire [127:0] col_645,
	output wire [127:0] col_646,
	output wire [127:0] col_647,
	output wire [127:0] col_648,
	output wire [127:0] col_649,
	output wire [127:0] col_650,
	output wire [127:0] col_651,
	output wire [127:0] col_652,
	output wire [127:0] col_653,
	output wire [127:0] col_654,
	output wire [127:0] col_655,
	output wire [127:0] col_656,
	output wire [127:0] col_657,
	output wire [127:0] col_658,
	output wire [127:0] col_659,
	output wire [127:0] col_660,
	output wire [127:0] col_661,
	output wire [127:0] col_662,
	output wire [127:0] col_663,
	output wire [127:0] col_664,
	output wire [127:0] col_665,
	output wire [127:0] col_666,
	output wire [127:0] col_667,
	output wire [127:0] col_668,
	output wire [127:0] col_669,
	output wire [127:0] col_670,
	output wire [127:0] col_671,
	output wire [127:0] col_672,
	output wire [127:0] col_673,
	output wire [127:0] col_674,
	output wire [127:0] col_675,
	output wire [127:0] col_676,
	output wire [127:0] col_677,
	output wire [127:0] col_678,
	output wire [127:0] col_679,
	output wire [127:0] col_680,
	output wire [127:0] col_681,
	output wire [127:0] col_682,
	output wire [127:0] col_683,
	output wire [127:0] col_684,
	output wire [127:0] col_685,
	output wire [127:0] col_686,
	output wire [127:0] col_687,
	output wire [127:0] col_688,
	output wire [127:0] col_689,
	output wire [127:0] col_690,
	output wire [127:0] col_691,
	output wire [127:0] col_692,
	output wire [127:0] col_693,
	output wire [127:0] col_694,
	output wire [127:0] col_695,
	output wire [127:0] col_696,
	output wire [127:0] col_697,
	output wire [127:0] col_698,
	output wire [127:0] col_699,
	output wire [127:0] col_700,
	output wire [127:0] col_701,
	output wire [127:0] col_702,
	output wire [127:0] col_703,
	output wire [127:0] col_704,
	output wire [127:0] col_705,
	output wire [127:0] col_706,
	output wire [127:0] col_707,
	output wire [127:0] col_708,
	output wire [127:0] col_709,
	output wire [127:0] col_710,
	output wire [127:0] col_711,
	output wire [127:0] col_712,
	output wire [127:0] col_713,
	output wire [127:0] col_714,
	output wire [127:0] col_715,
	output wire [127:0] col_716,
	output wire [127:0] col_717,
	output wire [127:0] col_718,
	output wire [127:0] col_719,
	output wire [127:0] col_720,
	output wire [127:0] col_721,
	output wire [127:0] col_722,
	output wire [127:0] col_723,
	output wire [127:0] col_724,
	output wire [127:0] col_725,
	output wire [127:0] col_726,
	output wire [127:0] col_727,
	output wire [127:0] col_728,
	output wire [127:0] col_729,
	output wire [127:0] col_730,
	output wire [127:0] col_731,
	output wire [127:0] col_732,
	output wire [127:0] col_733,
	output wire [127:0] col_734,
	output wire [127:0] col_735,
	output wire [127:0] col_736,
	output wire [127:0] col_737,
	output wire [127:0] col_738,
	output wire [127:0] col_739,
	output wire [127:0] col_740,
	output wire [127:0] col_741,
	output wire [127:0] col_742,
	output wire [127:0] col_743,
	output wire [127:0] col_744,
	output wire [127:0] col_745,
	output wire [127:0] col_746,
	output wire [127:0] col_747,
	output wire [127:0] col_748,
	output wire [127:0] col_749,
	output wire [127:0] col_750,
	output wire [127:0] col_751,
	output wire [127:0] col_752,
	output wire [127:0] col_753,
	output wire [127:0] col_754,
	output wire [127:0] col_755,
	output wire [127:0] col_756,
	output wire [127:0] col_757,
	output wire [127:0] col_758,
	output wire [127:0] col_759,
	output wire [127:0] col_760,
	output wire [127:0] col_761,
	output wire [127:0] col_762,
	output wire [127:0] col_763,
	output wire [127:0] col_764,
	output wire [127:0] col_765,
	output wire [127:0] col_766,
	output wire [127:0] col_767,
	output wire [127:0] col_768,
	output wire [127:0] col_769,
	output wire [127:0] col_770,
	output wire [127:0] col_771,
	output wire [127:0] col_772,
	output wire [127:0] col_773,
	output wire [127:0] col_774,
	output wire [127:0] col_775,
	output wire [127:0] col_776,
	output wire [127:0] col_777,
	output wire [127:0] col_778,
	output wire [127:0] col_779,
	output wire [127:0] col_780,
	output wire [127:0] col_781,
	output wire [127:0] col_782,
	output wire [127:0] col_783,
	output wire [127:0] col_784,
	output wire [127:0] col_785,
	output wire [127:0] col_786,
	output wire [127:0] col_787,
	output wire [127:0] col_788,
	output wire [127:0] col_789,
	output wire [127:0] col_790,
	output wire [127:0] col_791,
	output wire [127:0] col_792,
	output wire [127:0] col_793,
	output wire [127:0] col_794,
	output wire [127:0] col_795,
	output wire [127:0] col_796,
	output wire [127:0] col_797,
	output wire [127:0] col_798,
	output wire [127:0] col_799,
	output wire [127:0] col_800,
	output wire [127:0] col_801,
	output wire [127:0] col_802,
	output wire [127:0] col_803,
	output wire [127:0] col_804,
	output wire [127:0] col_805,
	output wire [127:0] col_806,
	output wire [127:0] col_807,
	output wire [127:0] col_808,
	output wire [127:0] col_809,
	output wire [127:0] col_810,
	output wire [127:0] col_811,
	output wire [127:0] col_812,
	output wire [127:0] col_813,
	output wire [127:0] col_814,
	output wire [127:0] col_815,
	output wire [127:0] col_816,
	output wire [127:0] col_817,
	output wire [127:0] col_818,
	output wire [127:0] col_819,
	output wire [127:0] col_820,
	output wire [127:0] col_821,
	output wire [127:0] col_822,
	output wire [127:0] col_823,
	output wire [127:0] col_824,
	output wire [127:0] col_825,
	output wire [127:0] col_826,
	output wire [127:0] col_827,
	output wire [127:0] col_828,
	output wire [127:0] col_829,
	output wire [127:0] col_830,
	output wire [127:0] col_831,
	output wire [127:0] col_832,
	output wire [127:0] col_833,
	output wire [127:0] col_834,
	output wire [127:0] col_835,
	output wire [127:0] col_836,
	output wire [127:0] col_837,
	output wire [127:0] col_838,
	output wire [127:0] col_839,
	output wire [127:0] col_840,
	output wire [127:0] col_841,
	output wire [127:0] col_842,
	output wire [127:0] col_843,
	output wire [127:0] col_844,
	output wire [127:0] col_845,
	output wire [127:0] col_846,
	output wire [127:0] col_847,
	output wire [127:0] col_848,
	output wire [127:0] col_849,
	output wire [127:0] col_850,
	output wire [127:0] col_851,
	output wire [127:0] col_852,
	output wire [127:0] col_853,
	output wire [127:0] col_854,
	output wire [127:0] col_855,
	output wire [127:0] col_856,
	output wire [127:0] col_857,
	output wire [127:0] col_858,
	output wire [127:0] col_859,
	output wire [127:0] col_860,
	output wire [127:0] col_861,
	output wire [127:0] col_862,
	output wire [127:0] col_863,
	output wire [127:0] col_864,
	output wire [127:0] col_865,
	output wire [127:0] col_866,
	output wire [127:0] col_867,
	output wire [127:0] col_868,
	output wire [127:0] col_869,
	output wire [127:0] col_870,
	output wire [127:0] col_871,
	output wire [127:0] col_872,
	output wire [127:0] col_873,
	output wire [127:0] col_874,
	output wire [127:0] col_875,
	output wire [127:0] col_876,
	output wire [127:0] col_877,
	output wire [127:0] col_878,
	output wire [127:0] col_879,
	output wire [127:0] col_880,
	output wire [127:0] col_881,
	output wire [127:0] col_882,
	output wire [127:0] col_883,
	output wire [127:0] col_884,
	output wire [127:0] col_885,
	output wire [127:0] col_886,
	output wire [127:0] col_887,
	output wire [127:0] col_888,
	output wire [127:0] col_889,
	output wire [127:0] col_890,
	output wire [127:0] col_891,
	output wire [127:0] col_892,
	output wire [127:0] col_893,
	output wire [127:0] col_894,
	output wire [127:0] col_895,
	output wire [127:0] col_896,
	output wire [127:0] col_897,
	output wire [127:0] col_898,
	output wire [127:0] col_899,
	output wire [127:0] col_900,
	output wire [127:0] col_901,
	output wire [127:0] col_902,
	output wire [127:0] col_903,
	output wire [127:0] col_904,
	output wire [127:0] col_905,
	output wire [127:0] col_906,
	output wire [127:0] col_907,
	output wire [127:0] col_908,
	output wire [127:0] col_909,
	output wire [127:0] col_910,
	output wire [127:0] col_911,
	output wire [127:0] col_912,
	output wire [127:0] col_913,
	output wire [127:0] col_914,
	output wire [127:0] col_915,
	output wire [127:0] col_916,
	output wire [127:0] col_917,
	output wire [127:0] col_918,
	output wire [127:0] col_919,
	output wire [127:0] col_920,
	output wire [127:0] col_921,
	output wire [127:0] col_922,
	output wire [127:0] col_923,
	output wire [127:0] col_924,
	output wire [127:0] col_925,
	output wire [127:0] col_926,
	output wire [127:0] col_927,
	output wire [127:0] col_928,
	output wire [127:0] col_929,
	output wire [127:0] col_930,
	output wire [127:0] col_931,
	output wire [127:0] col_932,
	output wire [127:0] col_933,
	output wire [127:0] col_934,
	output wire [127:0] col_935,
	output wire [127:0] col_936,
	output wire [127:0] col_937,
	output wire [127:0] col_938,
	output wire [127:0] col_939,
	output wire [127:0] col_940,
	output wire [127:0] col_941,
	output wire [127:0] col_942,
	output wire [127:0] col_943,
	output wire [127:0] col_944,
	output wire [127:0] col_945,
	output wire [127:0] col_946,
	output wire [127:0] col_947,
	output wire [127:0] col_948,
	output wire [127:0] col_949,
	output wire [127:0] col_950,
	output wire [127:0] col_951,
	output wire [127:0] col_952,
	output wire [127:0] col_953,
	output wire [127:0] col_954,
	output wire [127:0] col_955,
	output wire [127:0] col_956,
	output wire [127:0] col_957,
	output wire [127:0] col_958,
	output wire [127:0] col_959,
	output wire [127:0] col_960,
	output wire [127:0] col_961,
	output wire [127:0] col_962,
	output wire [127:0] col_963,
	output wire [127:0] col_964,
	output wire [127:0] col_965,
	output wire [127:0] col_966,
	output wire [127:0] col_967,
	output wire [127:0] col_968,
	output wire [127:0] col_969,
	output wire [127:0] col_970,
	output wire [127:0] col_971,
	output wire [127:0] col_972,
	output wire [127:0] col_973,
	output wire [127:0] col_974,
	output wire [127:0] col_975,
	output wire [127:0] col_976,
	output wire [127:0] col_977,
	output wire [127:0] col_978,
	output wire [127:0] col_979,
	output wire [127:0] col_980,
	output wire [127:0] col_981,
	output wire [127:0] col_982,
	output wire [127:0] col_983,
	output wire [127:0] col_984,
	output wire [127:0] col_985,
	output wire [127:0] col_986,
	output wire [127:0] col_987,
	output wire [127:0] col_988,
	output wire [127:0] col_989,
	output wire [127:0] col_990,
	output wire [127:0] col_991,
	output wire [127:0] col_992,
	output wire [127:0] col_993,
	output wire [127:0] col_994,
	output wire [127:0] col_995,
	output wire [127:0] col_996,
	output wire [127:0] col_997,
	output wire [127:0] col_998,
	output wire [127:0] col_999,
	output wire [127:0] col_1000,
	output wire [127:0] col_1001,
	output wire [127:0] col_1002,
	output wire [127:0] col_1003,
	output wire [127:0] col_1004,
	output wire [127:0] col_1005,
	output wire [127:0] col_1006,
	output wire [127:0] col_1007,
	output wire [127:0] col_1008,
	output wire [127:0] col_1009,
	output wire [127:0] col_1010,
	output wire [127:0] col_1011,
	output wire [127:0] col_1012,
	output wire [127:0] col_1013,
	output wire [127:0] col_1014,
	output wire [127:0] col_1015,
	output wire [127:0] col_1016,
	output wire [127:0] col_1017,
	output wire [127:0] col_1018,
	output wire [127:0] col_1019,
	output wire [127:0] col_1020,
	output wire [127:0] col_1021,
	output wire [127:0] col_1022,
	output wire [127:0] col_1023,
	output wire [127:0] col_1024,
	output wire [127:0] col_1025,
	output wire [127:0] col_1026,
	output wire [127:0] col_1027,
	output wire [127:0] col_1028,
	output wire [127:0] col_1029,
	output wire [127:0] col_1030,
	output wire [127:0] col_1031,
	output wire [127:0] col_1032,
	output wire [127:0] col_1033,
	output wire [127:0] col_1034,
	output wire [127:0] col_1035,
	output wire [127:0] col_1036,
	output wire [127:0] col_1037,
	output wire [127:0] col_1038,
	output wire [127:0] col_1039,
	output wire [127:0] col_1040,
	output wire [127:0] col_1041,
	output wire [127:0] col_1042,
	output wire [127:0] col_1043,
	output wire [127:0] col_1044,
	output wire [127:0] col_1045,
	output wire [127:0] col_1046,
	output wire [127:0] col_1047,
	output wire [127:0] col_1048,
	output wire [127:0] col_1049,
	output wire [127:0] col_1050,
	output wire [127:0] col_1051,
	output wire [127:0] col_1052,
	output wire [127:0] col_1053,
	output wire [127:0] col_1054,
	output wire [127:0] col_1055,
	output wire [127:0] col_1056,
	output wire [127:0] col_1057,
	output wire [127:0] col_1058,
	output wire [127:0] col_1059,
	output wire [127:0] col_1060,
	output wire [127:0] col_1061,
	output wire [127:0] col_1062,
	output wire [127:0] col_1063,
	output wire [127:0] col_1064,
	output wire [127:0] col_1065,
	output wire [127:0] col_1066,
	output wire [127:0] col_1067,
	output wire [127:0] col_1068,
	output wire [127:0] col_1069,
	output wire [127:0] col_1070,
	output wire [127:0] col_1071,
	output wire [127:0] col_1072,
	output wire [127:0] col_1073,
	output wire [127:0] col_1074,
	output wire [127:0] col_1075,
	output wire [127:0] col_1076,
	output wire [127:0] col_1077,
	output wire [127:0] col_1078,
	output wire [127:0] col_1079,
	output wire [127:0] col_1080,
	output wire [127:0] col_1081,
	output wire [127:0] col_1082,
	output wire [127:0] col_1083,
	output wire [127:0] col_1084,
	output wire [127:0] col_1085,
	output wire [127:0] col_1086,
	output wire [127:0] col_1087,
	output wire [127:0] col_1088,
	output wire [127:0] col_1089,
	output wire [127:0] col_1090,
	output wire [127:0] col_1091,
	output wire [127:0] col_1092,
	output wire [127:0] col_1093,
	output wire [127:0] col_1094,
	output wire [127:0] col_1095,
	output wire [127:0] col_1096,
	output wire [127:0] col_1097,
	output wire [127:0] col_1098,
	output wire [127:0] col_1099,
	output wire [127:0] col_1100,
	output wire [127:0] col_1101,
	output wire [127:0] col_1102,
	output wire [127:0] col_1103,
	output wire [127:0] col_1104,
	output wire [127:0] col_1105,
	output wire [127:0] col_1106,
	output wire [127:0] col_1107,
	output wire [127:0] col_1108,
	output wire [127:0] col_1109,
	output wire [127:0] col_1110,
	output wire [127:0] col_1111,
	output wire [127:0] col_1112,
	output wire [127:0] col_1113,
	output wire [127:0] col_1114,
	output wire [127:0] col_1115,
	output wire [127:0] col_1116,
	output wire [127:0] col_1117,
	output wire [127:0] col_1118,
	output wire [127:0] col_1119,
	output wire [127:0] col_1120,
	output wire [127:0] col_1121,
	output wire [127:0] col_1122,
	output wire [127:0] col_1123,
	output wire [127:0] col_1124,
	output wire [127:0] col_1125,
	output wire [127:0] col_1126,
	output wire [127:0] col_1127,
	output wire [127:0] col_1128,
	output wire [127:0] col_1129,
	output wire [127:0] col_1130,
	output wire [127:0] col_1131,
	output wire [127:0] col_1132,
	output wire [127:0] col_1133,
	output wire [127:0] col_1134,
	output wire [127:0] col_1135,
	output wire [127:0] col_1136,
	output wire [127:0] col_1137,
	output wire [127:0] col_1138,
	output wire [127:0] col_1139,
	output wire [127:0] col_1140,
	output wire [127:0] col_1141,
	output wire [127:0] col_1142,
	output wire [127:0] col_1143,
	output wire [127:0] col_1144,
	output wire [127:0] col_1145,
	output wire [127:0] col_1146,
	output wire [127:0] col_1147,
	output wire [127:0] col_1148,
	output wire [127:0] col_1149,
	output wire [127:0] col_1150,
	output wire [127:0] col_1151,
	output wire [127:0] col_1152,
	output wire [127:0] col_1153,
	output wire [127:0] col_1154,
	output wire [127:0] col_1155,
	output wire [127:0] col_1156,
	output wire [127:0] col_1157,
	output wire [127:0] col_1158,
	output wire [127:0] col_1159,
	output wire [127:0] col_1160,
	output wire [127:0] col_1161,
	output wire [127:0] col_1162,
	output wire [127:0] col_1163,
	output wire [127:0] col_1164,
	output wire [127:0] col_1165,
	output wire [127:0] col_1166,
	output wire [127:0] col_1167,
	output wire [127:0] col_1168,
	output wire [127:0] col_1169,
	output wire [127:0] col_1170,
	output wire [127:0] col_1171,
	output wire [127:0] col_1172,
	output wire [127:0] col_1173,
	output wire [127:0] col_1174,
	output wire [127:0] col_1175,
	output wire [127:0] col_1176,
	output wire [127:0] col_1177,
	output wire [127:0] col_1178,
	output wire [127:0] col_1179,
	output wire [127:0] col_1180,
	output wire [127:0] col_1181,
	output wire [127:0] col_1182,
	output wire [127:0] col_1183,
	output wire [127:0] col_1184,
	output wire [127:0] col_1185,
	output wire [127:0] col_1186,
	output wire [127:0] col_1187,
	output wire [127:0] col_1188,
	output wire [127:0] col_1189,
	output wire [127:0] col_1190,
	output wire [127:0] col_1191,
	output wire [127:0] col_1192,
	output wire [127:0] col_1193,
	output wire [127:0] col_1194,
	output wire [127:0] col_1195,
	output wire [127:0] col_1196,
	output wire [127:0] col_1197,
	output wire [127:0] col_1198,
	output wire [127:0] col_1199,
	output wire [127:0] col_1200,
	output wire [127:0] col_1201,
	output wire [127:0] col_1202,
	output wire [127:0] col_1203,
	output wire [127:0] col_1204,
	output wire [127:0] col_1205,
	output wire [127:0] col_1206,
	output wire [127:0] col_1207,
	output wire [127:0] col_1208,
	output wire [127:0] col_1209,
	output wire [127:0] col_1210,
	output wire [127:0] col_1211,
	output wire [127:0] col_1212,
	output wire [127:0] col_1213,
	output wire [127:0] col_1214,
	output wire [127:0] col_1215,
	output wire [127:0] col_1216,
	output wire [127:0] col_1217,
	output wire [127:0] col_1218,
	output wire [127:0] col_1219,
	output wire [127:0] col_1220,
	output wire [127:0] col_1221,
	output wire [127:0] col_1222,
	output wire [127:0] col_1223,
	output wire [127:0] col_1224,
	output wire [127:0] col_1225,
	output wire [127:0] col_1226,
	output wire [127:0] col_1227,
	output wire [127:0] col_1228,
	output wire [127:0] col_1229,
	output wire [127:0] col_1230,
	output wire [127:0] col_1231,
	output wire [127:0] col_1232,
	output wire [127:0] col_1233,
	output wire [127:0] col_1234,
	output wire [127:0] col_1235,
	output wire [127:0] col_1236,
	output wire [127:0] col_1237,
	output wire [127:0] col_1238,
	output wire [127:0] col_1239,
	output wire [127:0] col_1240,
	output wire [127:0] col_1241,
	output wire [127:0] col_1242,
	output wire [127:0] col_1243,
	output wire [127:0] col_1244,
	output wire [127:0] col_1245,
	output wire [127:0] col_1246,
	output wire [127:0] col_1247,
	output wire [127:0] col_1248,
	output wire [127:0] col_1249,
	output wire [127:0] col_1250,
	output wire [127:0] col_1251,
	output wire [127:0] col_1252,
	output wire [127:0] col_1253,
	output wire [127:0] col_1254,
	output wire [127:0] col_1255,
	output wire [127:0] col_1256,
	output wire [127:0] col_1257,
	output wire [127:0] col_1258,
	output wire [127:0] col_1259,
	output wire [127:0] col_1260,
	output wire [127:0] col_1261,
	output wire [127:0] col_1262,
	output wire [127:0] col_1263,
	output wire [127:0] col_1264,
	output wire [127:0] col_1265,
	output wire [127:0] col_1266,
	output wire [127:0] col_1267,
	output wire [127:0] col_1268,
	output wire [127:0] col_1269,
	output wire [127:0] col_1270,
	output wire [127:0] col_1271,
	output wire [127:0] col_1272,
	output wire [127:0] col_1273,
	output wire [127:0] col_1274,
	output wire [127:0] col_1275,
	output wire [127:0] col_1276,
	output wire [127:0] col_1277,
	output wire [127:0] col_1278,
	output wire [127:0] col_1279
);


wire [1021:0] ctrl_1;
wire [1021:0] ctrl_2;
wire [1021:0] ctrl_3;
wire [1021:0] ctrl_4;
wire [1021:0] ctrl_5;
wire [1021:0] ctrl_6;
wire [1021:0] ctrl_7;
wire [1021:0] ctrl_8;
wire [1021:0] ctrl_9;
wire [1021:0] ctrl_10;
wire [1021:0] ctrl_11;
wire [1021:0] ctrl_12;
wire [1021:0] ctrl_13;
wire [1021:0] ctrl_14;
wire [1021:0] ctrl_15;
wire [1021:0] ctrl_16;
wire [1021:0] ctrl_17;
wire [1021:0] ctrl_18;
wire [1021:0] ctrl_19;
wire [1021:0] ctrl_20;
wire [1021:0] ctrl_21;
wire [1021:0] ctrl_22;
wire [1021:0] ctrl_23;
wire [1021:0] ctrl_24;
wire [1021:0] ctrl_25;
wire [1021:0] ctrl_26;
wire [1021:0] ctrl_27;
wire [1021:0] ctrl_28;
wire [1021:0] ctrl_29;
wire [1021:0] ctrl_30;
wire [1021:0] ctrl_31;
wire [1021:0] ctrl_32;
wire [1021:0] ctrl_33;
wire [1021:0] ctrl_34;
wire [1021:0] ctrl_35;
wire [1021:0] ctrl_36;
wire [1021:0] ctrl_37;
wire [1021:0] ctrl_38;
wire [1021:0] ctrl_39;
wire [1021:0] ctrl_40;
wire [1021:0] ctrl_41;
wire [1021:0] ctrl_42;
wire [1021:0] ctrl_43;
wire [1021:0] ctrl_44;
wire [1021:0] ctrl_45;
wire [1021:0] ctrl_46;
wire [1021:0] ctrl_47;
wire [1021:0] ctrl_48;
wire [1021:0] ctrl_49;
wire [1021:0] ctrl_50;
wire [1021:0] ctrl_51;
wire [1021:0] ctrl_52;
wire [1021:0] ctrl_53;
wire [1021:0] ctrl_54;
wire [1021:0] ctrl_55;
wire [1021:0] ctrl_56;
wire [1021:0] ctrl_57;
wire [1021:0] ctrl_58;
wire [1021:0] ctrl_59;
wire [1021:0] ctrl_60;
wire [1021:0] ctrl_61;
wire [1021:0] ctrl_62;
wire [1021:0] ctrl_63;
wire [1021:0] ctrl_64;
wire [1021:0] ctrl_65;
wire [1021:0] ctrl_66;
wire [1021:0] ctrl_67;
wire [1021:0] ctrl_68;
wire [1021:0] ctrl_69;
wire [1021:0] ctrl_70;
wire [1021:0] ctrl_71;
wire [1021:0] ctrl_72;
wire [1021:0] ctrl_73;
wire [1021:0] ctrl_74;
wire [1021:0] ctrl_75;
wire [1021:0] ctrl_76;
wire [1021:0] ctrl_77;
wire [1021:0] ctrl_78;
wire [1021:0] ctrl_79;
wire [1021:0] ctrl_80;
wire [1021:0] ctrl_81;
wire [1021:0] ctrl_82;
wire [1021:0] ctrl_83;
wire [1021:0] ctrl_84;
wire [1021:0] ctrl_85;
wire [1021:0] ctrl_86;
wire [1021:0] ctrl_87;
wire [1021:0] ctrl_88;
wire [1021:0] ctrl_89;
wire [1021:0] ctrl_90;
wire [1021:0] ctrl_91;
wire [1021:0] ctrl_92;
wire [1021:0] ctrl_93;
wire [1021:0] ctrl_94;
wire [1021:0] ctrl_95;
wire [1021:0] ctrl_96;
wire [1021:0] ctrl_97;
wire [1021:0] ctrl_98;
wire [1021:0] ctrl_99;
wire [1021:0] ctrl_100;
wire [1021:0] ctrl_101;
wire [1021:0] ctrl_102;
wire [1021:0] ctrl_103;
wire [1021:0] ctrl_104;
wire [1021:0] ctrl_105;
wire [1021:0] ctrl_106;
wire [1021:0] ctrl_107;
wire [1021:0] ctrl_108;
wire [1021:0] ctrl_109;
wire [1021:0] ctrl_110;
wire [1021:0] ctrl_111;
wire [1021:0] ctrl_112;
wire [1021:0] ctrl_113;
wire [1021:0] ctrl_114;
wire [1021:0] ctrl_115;
wire [1021:0] ctrl_116;
wire [1021:0] ctrl_117;
wire [1021:0] ctrl_118;
wire [1021:0] ctrl_119;
wire [1021:0] ctrl_120;
wire [1021:0] ctrl_121;
wire [1021:0] ctrl_122;
wire [1021:0] ctrl_123;
wire [1021:0] ctrl_124;
wire [1021:0] ctrl_125;
wire [1021:0] ctrl_126;
wire [1021:0] ctrl_127;
wire [1021:0] ctrl_128;

wire [1021:0] a_left_1;
wire [1021:0] a_left_2;
wire [1021:0] a_left_3;
wire [1021:0] a_left_4;
wire [1021:0] a_left_5;
wire [1021:0] a_left_6;
wire [1021:0] a_left_7;
wire [1021:0] a_left_8;
wire [1021:0] a_left_9;
wire [1021:0] a_left_10;
wire [1021:0] a_left_11;
wire [1021:0] a_left_12;
wire [1021:0] a_left_13;
wire [1021:0] a_left_14;
wire [1021:0] a_left_15;
wire [1021:0] a_left_16;
wire [1021:0] a_left_17;
wire [1021:0] a_left_18;
wire [1021:0] a_left_19;
wire [1021:0] a_left_20;
wire [1021:0] a_left_21;
wire [1021:0] a_left_22;
wire [1021:0] a_left_23;
wire [1021:0] a_left_24;
wire [1021:0] a_left_25;
wire [1021:0] a_left_26;
wire [1021:0] a_left_27;
wire [1021:0] a_left_28;
wire [1021:0] a_left_29;
wire [1021:0] a_left_30;
wire [1021:0] a_left_31;
wire [1021:0] a_left_32;
wire [1021:0] a_left_33;
wire [1021:0] a_left_34;
wire [1021:0] a_left_35;
wire [1021:0] a_left_36;
wire [1021:0] a_left_37;
wire [1021:0] a_left_38;
wire [1021:0] a_left_39;
wire [1021:0] a_left_40;
wire [1021:0] a_left_41;
wire [1021:0] a_left_42;
wire [1021:0] a_left_43;
wire [1021:0] a_left_44;
wire [1021:0] a_left_45;
wire [1021:0] a_left_46;
wire [1021:0] a_left_47;
wire [1021:0] a_left_48;
wire [1021:0] a_left_49;
wire [1021:0] a_left_50;
wire [1021:0] a_left_51;
wire [1021:0] a_left_52;
wire [1021:0] a_left_53;
wire [1021:0] a_left_54;
wire [1021:0] a_left_55;
wire [1021:0] a_left_56;
wire [1021:0] a_left_57;
wire [1021:0] a_left_58;
wire [1021:0] a_left_59;
wire [1021:0] a_left_60;
wire [1021:0] a_left_61;
wire [1021:0] a_left_62;
wire [1021:0] a_left_63;
wire [1021:0] a_left_64;
wire [1021:0] a_left_65;
wire [1021:0] a_left_66;
wire [1021:0] a_left_67;
wire [1021:0] a_left_68;
wire [1021:0] a_left_69;
wire [1021:0] a_left_70;
wire [1021:0] a_left_71;
wire [1021:0] a_left_72;
wire [1021:0] a_left_73;
wire [1021:0] a_left_74;
wire [1021:0] a_left_75;
wire [1021:0] a_left_76;
wire [1021:0] a_left_77;
wire [1021:0] a_left_78;
wire [1021:0] a_left_79;
wire [1021:0] a_left_80;
wire [1021:0] a_left_81;
wire [1021:0] a_left_82;
wire [1021:0] a_left_83;
wire [1021:0] a_left_84;
wire [1021:0] a_left_85;
wire [1021:0] a_left_86;
wire [1021:0] a_left_87;
wire [1021:0] a_left_88;
wire [1021:0] a_left_89;
wire [1021:0] a_left_90;
wire [1021:0] a_left_91;
wire [1021:0] a_left_92;
wire [1021:0] a_left_93;
wire [1021:0] a_left_94;
wire [1021:0] a_left_95;
wire [1021:0] a_left_96;
wire [1021:0] a_left_97;
wire [1021:0] a_left_98;
wire [1021:0] a_left_99;
wire [1021:0] a_left_100;
wire [1021:0] a_left_101;
wire [1021:0] a_left_102;
wire [1021:0] a_left_103;
wire [1021:0] a_left_104;
wire [1021:0] a_left_105;
wire [1021:0] a_left_106;
wire [1021:0] a_left_107;
wire [1021:0] a_left_108;
wire [1021:0] a_left_109;
wire [1021:0] a_left_110;
wire [1021:0] a_left_111;
wire [1021:0] a_left_112;
wire [1021:0] a_left_113;
wire [1021:0] a_left_114;
wire [1021:0] a_left_115;
wire [1021:0] a_left_116;
wire [1021:0] a_left_117;
wire [1021:0] a_left_118;
wire [1021:0] a_left_119;
wire [1021:0] a_left_120;
wire [1021:0] a_left_121;
wire [1021:0] a_left_122;
wire [1021:0] a_left_123;
wire [1021:0] a_left_124;
wire [1021:0] a_left_125;
wire [1021:0] a_left_126;
wire [1021:0] a_left_127;
wire [1021:0] a_left_128;

wire [1021:0] a_right_1;
wire [1021:0] a_right_2;
wire [1021:0] a_right_3;
wire [1021:0] a_right_4;
wire [1021:0] a_right_5;
wire [1021:0] a_right_6;
wire [1021:0] a_right_7;
wire [1021:0] a_right_8;
wire [1021:0] a_right_9;
wire [1021:0] a_right_10;
wire [1021:0] a_right_11;
wire [1021:0] a_right_12;
wire [1021:0] a_right_13;
wire [1021:0] a_right_14;
wire [1021:0] a_right_15;
wire [1021:0] a_right_16;
wire [1021:0] a_right_17;
wire [1021:0] a_right_18;
wire [1021:0] a_right_19;
wire [1021:0] a_right_20;
wire [1021:0] a_right_21;
wire [1021:0] a_right_22;
wire [1021:0] a_right_23;
wire [1021:0] a_right_24;
wire [1021:0] a_right_25;
wire [1021:0] a_right_26;
wire [1021:0] a_right_27;
wire [1021:0] a_right_28;
wire [1021:0] a_right_29;
wire [1021:0] a_right_30;
wire [1021:0] a_right_31;
wire [1021:0] a_right_32;
wire [1021:0] a_right_33;
wire [1021:0] a_right_34;
wire [1021:0] a_right_35;
wire [1021:0] a_right_36;
wire [1021:0] a_right_37;
wire [1021:0] a_right_38;
wire [1021:0] a_right_39;
wire [1021:0] a_right_40;
wire [1021:0] a_right_41;
wire [1021:0] a_right_42;
wire [1021:0] a_right_43;
wire [1021:0] a_right_44;
wire [1021:0] a_right_45;
wire [1021:0] a_right_46;
wire [1021:0] a_right_47;
wire [1021:0] a_right_48;
wire [1021:0] a_right_49;
wire [1021:0] a_right_50;
wire [1021:0] a_right_51;
wire [1021:0] a_right_52;
wire [1021:0] a_right_53;
wire [1021:0] a_right_54;
wire [1021:0] a_right_55;
wire [1021:0] a_right_56;
wire [1021:0] a_right_57;
wire [1021:0] a_right_58;
wire [1021:0] a_right_59;
wire [1021:0] a_right_60;
wire [1021:0] a_right_61;
wire [1021:0] a_right_62;
wire [1021:0] a_right_63;
wire [1021:0] a_right_64;
wire [1021:0] a_right_65;
wire [1021:0] a_right_66;
wire [1021:0] a_right_67;
wire [1021:0] a_right_68;
wire [1021:0] a_right_69;
wire [1021:0] a_right_70;
wire [1021:0] a_right_71;
wire [1021:0] a_right_72;
wire [1021:0] a_right_73;
wire [1021:0] a_right_74;
wire [1021:0] a_right_75;
wire [1021:0] a_right_76;
wire [1021:0] a_right_77;
wire [1021:0] a_right_78;
wire [1021:0] a_right_79;
wire [1021:0] a_right_80;
wire [1021:0] a_right_81;
wire [1021:0] a_right_82;
wire [1021:0] a_right_83;
wire [1021:0] a_right_84;
wire [1021:0] a_right_85;
wire [1021:0] a_right_86;
wire [1021:0] a_right_87;
wire [1021:0] a_right_88;
wire [1021:0] a_right_89;
wire [1021:0] a_right_90;
wire [1021:0] a_right_91;
wire [1021:0] a_right_92;
wire [1021:0] a_right_93;
wire [1021:0] a_right_94;
wire [1021:0] a_right_95;
wire [1021:0] a_right_96;
wire [1021:0] a_right_97;
wire [1021:0] a_right_98;
wire [1021:0] a_right_99;
wire [1021:0] a_right_100;
wire [1021:0] a_right_101;
wire [1021:0] a_right_102;
wire [1021:0] a_right_103;
wire [1021:0] a_right_104;
wire [1021:0] a_right_105;
wire [1021:0] a_right_106;
wire [1021:0] a_right_107;
wire [1021:0] a_right_108;
wire [1021:0] a_right_109;
wire [1021:0] a_right_110;
wire [1021:0] a_right_111;
wire [1021:0] a_right_112;
wire [1021:0] a_right_113;
wire [1021:0] a_right_114;
wire [1021:0] a_right_115;
wire [1021:0] a_right_116;
wire [1021:0] a_right_117;
wire [1021:0] a_right_118;
wire [1021:0] a_right_119;
wire [1021:0] a_right_120;
wire [1021:0] a_right_121;
wire [1021:0] a_right_122;
wire [1021:0] a_right_123;
wire [1021:0] a_right_124;
wire [1021:0] a_right_125;
wire [1021:0] a_right_126;
wire [1021:0] a_right_127;
wire [1021:0] a_right_128;

wire [1025:0] line_1;
wire [1025:0] line_2;
wire [1025:0] line_3;
wire [1025:0] line_4;
wire [1025:0] line_5;
wire [1025:0] line_6;
wire [1025:0] line_7;
wire [1025:0] line_8;
wire [1025:0] line_9;
wire [1025:0] line_10;
wire [1025:0] line_11;
wire [1025:0] line_12;
wire [1025:0] line_13;
wire [1025:0] line_14;
wire [1025:0] line_15;
wire [1025:0] line_16;
wire [1025:0] line_17;
wire [1025:0] line_18;
wire [1025:0] line_19;
wire [1025:0] line_20;
wire [1025:0] line_21;
wire [1025:0] line_22;
wire [1025:0] line_23;
wire [1025:0] line_24;
wire [1025:0] line_25;
wire [1025:0] line_26;
wire [1025:0] line_27;
wire [1025:0] line_28;
wire [1025:0] line_29;
wire [1025:0] line_30;
wire [1025:0] line_31;
wire [1025:0] line_32;
wire [1025:0] line_33;
wire [1025:0] line_34;
wire [1025:0] line_35;
wire [1025:0] line_36;
wire [1025:0] line_37;
wire [1025:0] line_38;
wire [1025:0] line_39;
wire [1025:0] line_40;
wire [1025:0] line_41;
wire [1025:0] line_42;
wire [1025:0] line_43;
wire [1025:0] line_44;
wire [1025:0] line_45;
wire [1025:0] line_46;
wire [1025:0] line_47;
wire [1025:0] line_48;
wire [1025:0] line_49;
wire [1025:0] line_50;
wire [1025:0] line_51;
wire [1025:0] line_52;
wire [1025:0] line_53;
wire [1025:0] line_54;
wire [1025:0] line_55;
wire [1025:0] line_56;
wire [1025:0] line_57;
wire [1025:0] line_58;
wire [1025:0] line_59;
wire [1025:0] line_60;
wire [1025:0] line_61;
wire [1025:0] line_62;
wire [1025:0] line_63;
wire [1025:0] line_64;
wire [1025:0] line_65;
wire [1025:0] line_66;
wire [1025:0] line_67;
wire [1025:0] line_68;
wire [1025:0] line_69;
wire [1025:0] line_70;
wire [1025:0] line_71;
wire [1025:0] line_72;
wire [1025:0] line_73;
wire [1025:0] line_74;
wire [1025:0] line_75;
wire [1025:0] line_76;
wire [1025:0] line_77;
wire [1025:0] line_78;
wire [1025:0] line_79;
wire [1025:0] line_80;
wire [1025:0] line_81;
wire [1025:0] line_82;
wire [1025:0] line_83;
wire [1025:0] line_84;
wire [1025:0] line_85;
wire [1025:0] line_86;
wire [1025:0] line_87;
wire [1025:0] line_88;
wire [1025:0] line_89;
wire [1025:0] line_90;
wire [1025:0] line_91;
wire [1025:0] line_92;
wire [1025:0] line_93;
wire [1025:0] line_94;
wire [1025:0] line_95;
wire [1025:0] line_96;
wire [1025:0] line_97;
wire [1025:0] line_98;
wire [1025:0] line_99;
wire [1025:0] line_100;
wire [1025:0] line_101;
wire [1025:0] line_102;
wire [1025:0] line_103;
wire [1025:0] line_104;
wire [1025:0] line_105;
wire [1025:0] line_106;
wire [1025:0] line_107;
wire [1025:0] line_108;
wire [1025:0] line_109;
wire [1025:0] line_110;
wire [1025:0] line_111;
wire [1025:0] line_112;
wire [1025:0] line_113;
wire [1025:0] line_114;
wire [1025:0] line_115;
wire [1025:0] line_116;
wire [1025:0] line_117;
wire [1025:0] line_118;
wire [1025:0] line_119;
wire [1025:0] line_120;
wire [1025:0] line_121;
wire [1025:0] line_122;
wire [1025:0] line_123;
wire [1025:0] line_124;
wire [1025:0] line_125;
wire [1025:0] line_126;
wire [1025:0] line_127;
wire [1025:0] line_128;

ctrl_gene ctrl_gene (
	.sel(sel),
	.ctrl_1(ctrl_1),
	.ctrl_2(ctrl_2),
	.ctrl_3(ctrl_3),
	.ctrl_4(ctrl_4),
	.ctrl_5(ctrl_5),
	.ctrl_6(ctrl_6),
	.ctrl_7(ctrl_7),
	.ctrl_8(ctrl_8),
	.ctrl_9(ctrl_9),
	.ctrl_10(ctrl_10),
	.ctrl_11(ctrl_11),
	.ctrl_12(ctrl_12),
	.ctrl_13(ctrl_13),
	.ctrl_14(ctrl_14),
	.ctrl_15(ctrl_15),
	.ctrl_16(ctrl_16),
	.ctrl_17(ctrl_17),
	.ctrl_18(ctrl_18),
	.ctrl_19(ctrl_19),
	.ctrl_20(ctrl_20),
	.ctrl_21(ctrl_21),
	.ctrl_22(ctrl_22),
	.ctrl_23(ctrl_23),
	.ctrl_24(ctrl_24),
	.ctrl_25(ctrl_25),
	.ctrl_26(ctrl_26),
	.ctrl_27(ctrl_27),
	.ctrl_28(ctrl_28),
	.ctrl_29(ctrl_29),
	.ctrl_30(ctrl_30),
	.ctrl_31(ctrl_31),
	.ctrl_32(ctrl_32),
	.ctrl_33(ctrl_33),
	.ctrl_34(ctrl_34),
	.ctrl_35(ctrl_35),
	.ctrl_36(ctrl_36),
	.ctrl_37(ctrl_37),
	.ctrl_38(ctrl_38),
	.ctrl_39(ctrl_39),
	.ctrl_40(ctrl_40),
	.ctrl_41(ctrl_41),
	.ctrl_42(ctrl_42),
	.ctrl_43(ctrl_43),
	.ctrl_44(ctrl_44),
	.ctrl_45(ctrl_45),
	.ctrl_46(ctrl_46),
	.ctrl_47(ctrl_47),
	.ctrl_48(ctrl_48),
	.ctrl_49(ctrl_49),
	.ctrl_50(ctrl_50),
	.ctrl_51(ctrl_51),
	.ctrl_52(ctrl_52),
	.ctrl_53(ctrl_53),
	.ctrl_54(ctrl_54),
	.ctrl_55(ctrl_55),
	.ctrl_56(ctrl_56),
	.ctrl_57(ctrl_57),
	.ctrl_58(ctrl_58),
	.ctrl_59(ctrl_59),
	.ctrl_60(ctrl_60),
	.ctrl_61(ctrl_61),
	.ctrl_62(ctrl_62),
	.ctrl_63(ctrl_63),
	.ctrl_64(ctrl_64),
	.ctrl_65(ctrl_65),
	.ctrl_66(ctrl_66),
	.ctrl_67(ctrl_67),
	.ctrl_68(ctrl_68),
	.ctrl_69(ctrl_69),
	.ctrl_70(ctrl_70),
	.ctrl_71(ctrl_71),
	.ctrl_72(ctrl_72),
	.ctrl_73(ctrl_73),
	.ctrl_74(ctrl_74),
	.ctrl_75(ctrl_75),
	.ctrl_76(ctrl_76),
	.ctrl_77(ctrl_77),
	.ctrl_78(ctrl_78),
	.ctrl_79(ctrl_79),
	.ctrl_80(ctrl_80),
	.ctrl_81(ctrl_81),
	.ctrl_82(ctrl_82),
	.ctrl_83(ctrl_83),
	.ctrl_84(ctrl_84),
	.ctrl_85(ctrl_85),
	.ctrl_86(ctrl_86),
	.ctrl_87(ctrl_87),
	.ctrl_88(ctrl_88),
	.ctrl_89(ctrl_89),
	.ctrl_90(ctrl_90),
	.ctrl_91(ctrl_91),
	.ctrl_92(ctrl_92),
	.ctrl_93(ctrl_93),
	.ctrl_94(ctrl_94),
	.ctrl_95(ctrl_95),
	.ctrl_96(ctrl_96),
	.ctrl_97(ctrl_97),
	.ctrl_98(ctrl_98),
	.ctrl_99(ctrl_99),
	.ctrl_100(ctrl_100),
	.ctrl_101(ctrl_101),
	.ctrl_102(ctrl_102),
	.ctrl_103(ctrl_103),
	.ctrl_104(ctrl_104),
	.ctrl_105(ctrl_105),
	.ctrl_106(ctrl_106),
	.ctrl_107(ctrl_107),
	.ctrl_108(ctrl_108),
	.ctrl_109(ctrl_109),
	.ctrl_110(ctrl_110),
	.ctrl_111(ctrl_111),
	.ctrl_112(ctrl_112),
	.ctrl_113(ctrl_113),
	.ctrl_114(ctrl_114),
	.ctrl_115(ctrl_115),
	.ctrl_116(ctrl_116),
	.ctrl_117(ctrl_117),
	.ctrl_118(ctrl_118),
	.ctrl_119(ctrl_119),
	.ctrl_120(ctrl_120),
	.ctrl_121(ctrl_121),
	.ctrl_122(ctrl_122),
	.ctrl_123(ctrl_123),
	.ctrl_124(ctrl_124),
	.ctrl_125(ctrl_125),
	.ctrl_126(ctrl_126),
	.ctrl_127(ctrl_127),
	.ctrl_128(ctrl_128)
);

sel_and_array_in sel_and_array_in (
	.al(al),
	.ctrl_1(ctrl_1),
	.ctrl_2(ctrl_2),
	.ctrl_3(ctrl_3),
	.ctrl_4(ctrl_4),
	.ctrl_5(ctrl_5),
	.ctrl_6(ctrl_6),
	.ctrl_7(ctrl_7),
	.ctrl_8(ctrl_8),
	.ctrl_9(ctrl_9),
	.ctrl_10(ctrl_10),
	.ctrl_11(ctrl_11),
	.ctrl_12(ctrl_12),
	.ctrl_13(ctrl_13),
	.ctrl_14(ctrl_14),
	.ctrl_15(ctrl_15),
	.ctrl_16(ctrl_16),
	.ctrl_17(ctrl_17),
	.ctrl_18(ctrl_18),
	.ctrl_19(ctrl_19),
	.ctrl_20(ctrl_20),
	.ctrl_21(ctrl_21),
	.ctrl_22(ctrl_22),
	.ctrl_23(ctrl_23),
	.ctrl_24(ctrl_24),
	.ctrl_25(ctrl_25),
	.ctrl_26(ctrl_26),
	.ctrl_27(ctrl_27),
	.ctrl_28(ctrl_28),
	.ctrl_29(ctrl_29),
	.ctrl_30(ctrl_30),
	.ctrl_31(ctrl_31),
	.ctrl_32(ctrl_32),
	.ctrl_33(ctrl_33),
	.ctrl_34(ctrl_34),
	.ctrl_35(ctrl_35),
	.ctrl_36(ctrl_36),
	.ctrl_37(ctrl_37),
	.ctrl_38(ctrl_38),
	.ctrl_39(ctrl_39),
	.ctrl_40(ctrl_40),
	.ctrl_41(ctrl_41),
	.ctrl_42(ctrl_42),
	.ctrl_43(ctrl_43),
	.ctrl_44(ctrl_44),
	.ctrl_45(ctrl_45),
	.ctrl_46(ctrl_46),
	.ctrl_47(ctrl_47),
	.ctrl_48(ctrl_48),
	.ctrl_49(ctrl_49),
	.ctrl_50(ctrl_50),
	.ctrl_51(ctrl_51),
	.ctrl_52(ctrl_52),
	.ctrl_53(ctrl_53),
	.ctrl_54(ctrl_54),
	.ctrl_55(ctrl_55),
	.ctrl_56(ctrl_56),
	.ctrl_57(ctrl_57),
	.ctrl_58(ctrl_58),
	.ctrl_59(ctrl_59),
	.ctrl_60(ctrl_60),
	.ctrl_61(ctrl_61),
	.ctrl_62(ctrl_62),
	.ctrl_63(ctrl_63),
	.ctrl_64(ctrl_64),
	.ctrl_65(ctrl_65),
	.ctrl_66(ctrl_66),
	.ctrl_67(ctrl_67),
	.ctrl_68(ctrl_68),
	.ctrl_69(ctrl_69),
	.ctrl_70(ctrl_70),
	.ctrl_71(ctrl_71),
	.ctrl_72(ctrl_72),
	.ctrl_73(ctrl_73),
	.ctrl_74(ctrl_74),
	.ctrl_75(ctrl_75),
	.ctrl_76(ctrl_76),
	.ctrl_77(ctrl_77),
	.ctrl_78(ctrl_78),
	.ctrl_79(ctrl_79),
	.ctrl_80(ctrl_80),
	.ctrl_81(ctrl_81),
	.ctrl_82(ctrl_82),
	.ctrl_83(ctrl_83),
	.ctrl_84(ctrl_84),
	.ctrl_85(ctrl_85),
	.ctrl_86(ctrl_86),
	.ctrl_87(ctrl_87),
	.ctrl_88(ctrl_88),
	.ctrl_89(ctrl_89),
	.ctrl_90(ctrl_90),
	.ctrl_91(ctrl_91),
	.ctrl_92(ctrl_92),
	.ctrl_93(ctrl_93),
	.ctrl_94(ctrl_94),
	.ctrl_95(ctrl_95),
	.ctrl_96(ctrl_96),
	.ctrl_97(ctrl_97),
	.ctrl_98(ctrl_98),
	.ctrl_99(ctrl_99),
	.ctrl_100(ctrl_100),
	.ctrl_101(ctrl_101),
	.ctrl_102(ctrl_102),
	.ctrl_103(ctrl_103),
	.ctrl_104(ctrl_104),
	.ctrl_105(ctrl_105),
	.ctrl_106(ctrl_106),
	.ctrl_107(ctrl_107),
	.ctrl_108(ctrl_108),
	.ctrl_109(ctrl_109),
	.ctrl_110(ctrl_110),
	.ctrl_111(ctrl_111),
	.ctrl_112(ctrl_112),
	.ctrl_113(ctrl_113),
	.ctrl_114(ctrl_114),
	.ctrl_115(ctrl_115),
	.ctrl_116(ctrl_116),
	.ctrl_117(ctrl_117),
	.ctrl_118(ctrl_118),
	.ctrl_119(ctrl_119),
	.ctrl_120(ctrl_120),
	.ctrl_121(ctrl_121),
	.ctrl_122(ctrl_122),
	.ctrl_123(ctrl_123),
	.ctrl_124(ctrl_124),
	.ctrl_125(ctrl_125),
	.ctrl_126(ctrl_126),
	.ctrl_127(ctrl_127),
	.ctrl_128(ctrl_128),
	.a_left_1(a_left_1),
	.a_left_2(a_left_2),
	.a_left_3(a_left_3),
	.a_left_4(a_left_4),
	.a_left_5(a_left_5),
	.a_left_6(a_left_6),
	.a_left_7(a_left_7),
	.a_left_8(a_left_8),
	.a_left_9(a_left_9),
	.a_left_10(a_left_10),
	.a_left_11(a_left_11),
	.a_left_12(a_left_12),
	.a_left_13(a_left_13),
	.a_left_14(a_left_14),
	.a_left_15(a_left_15),
	.a_left_16(a_left_16),
	.a_left_17(a_left_17),
	.a_left_18(a_left_18),
	.a_left_19(a_left_19),
	.a_left_20(a_left_20),
	.a_left_21(a_left_21),
	.a_left_22(a_left_22),
	.a_left_23(a_left_23),
	.a_left_24(a_left_24),
	.a_left_25(a_left_25),
	.a_left_26(a_left_26),
	.a_left_27(a_left_27),
	.a_left_28(a_left_28),
	.a_left_29(a_left_29),
	.a_left_30(a_left_30),
	.a_left_31(a_left_31),
	.a_left_32(a_left_32),
	.a_left_33(a_left_33),
	.a_left_34(a_left_34),
	.a_left_35(a_left_35),
	.a_left_36(a_left_36),
	.a_left_37(a_left_37),
	.a_left_38(a_left_38),
	.a_left_39(a_left_39),
	.a_left_40(a_left_40),
	.a_left_41(a_left_41),
	.a_left_42(a_left_42),
	.a_left_43(a_left_43),
	.a_left_44(a_left_44),
	.a_left_45(a_left_45),
	.a_left_46(a_left_46),
	.a_left_47(a_left_47),
	.a_left_48(a_left_48),
	.a_left_49(a_left_49),
	.a_left_50(a_left_50),
	.a_left_51(a_left_51),
	.a_left_52(a_left_52),
	.a_left_53(a_left_53),
	.a_left_54(a_left_54),
	.a_left_55(a_left_55),
	.a_left_56(a_left_56),
	.a_left_57(a_left_57),
	.a_left_58(a_left_58),
	.a_left_59(a_left_59),
	.a_left_60(a_left_60),
	.a_left_61(a_left_61),
	.a_left_62(a_left_62),
	.a_left_63(a_left_63),
	.a_left_64(a_left_64),
	.a_left_65(a_left_65),
	.a_left_66(a_left_66),
	.a_left_67(a_left_67),
	.a_left_68(a_left_68),
	.a_left_69(a_left_69),
	.a_left_70(a_left_70),
	.a_left_71(a_left_71),
	.a_left_72(a_left_72),
	.a_left_73(a_left_73),
	.a_left_74(a_left_74),
	.a_left_75(a_left_75),
	.a_left_76(a_left_76),
	.a_left_77(a_left_77),
	.a_left_78(a_left_78),
	.a_left_79(a_left_79),
	.a_left_80(a_left_80),
	.a_left_81(a_left_81),
	.a_left_82(a_left_82),
	.a_left_83(a_left_83),
	.a_left_84(a_left_84),
	.a_left_85(a_left_85),
	.a_left_86(a_left_86),
	.a_left_87(a_left_87),
	.a_left_88(a_left_88),
	.a_left_89(a_left_89),
	.a_left_90(a_left_90),
	.a_left_91(a_left_91),
	.a_left_92(a_left_92),
	.a_left_93(a_left_93),
	.a_left_94(a_left_94),
	.a_left_95(a_left_95),
	.a_left_96(a_left_96),
	.a_left_97(a_left_97),
	.a_left_98(a_left_98),
	.a_left_99(a_left_99),
	.a_left_100(a_left_100),
	.a_left_101(a_left_101),
	.a_left_102(a_left_102),
	.a_left_103(a_left_103),
	.a_left_104(a_left_104),
	.a_left_105(a_left_105),
	.a_left_106(a_left_106),
	.a_left_107(a_left_107),
	.a_left_108(a_left_108),
	.a_left_109(a_left_109),
	.a_left_110(a_left_110),
	.a_left_111(a_left_111),
	.a_left_112(a_left_112),
	.a_left_113(a_left_113),
	.a_left_114(a_left_114),
	.a_left_115(a_left_115),
	.a_left_116(a_left_116),
	.a_left_117(a_left_117),
	.a_left_118(a_left_118),
	.a_left_119(a_left_119),
	.a_left_120(a_left_120),
	.a_left_121(a_left_121),
	.a_left_122(a_left_122),
	.a_left_123(a_left_123),
	.a_left_124(a_left_124),
	.a_left_125(a_left_125),
	.a_left_126(a_left_126),
	.a_left_127(a_left_127),
	.a_left_128(a_left_128),
	.a_right_1(a_right_1),
	.a_right_2(a_right_2),
	.a_right_3(a_right_3),
	.a_right_4(a_right_4),
	.a_right_5(a_right_5),
	.a_right_6(a_right_6),
	.a_right_7(a_right_7),
	.a_right_8(a_right_8),
	.a_right_9(a_right_9),
	.a_right_10(a_right_10),
	.a_right_11(a_right_11),
	.a_right_12(a_right_12),
	.a_right_13(a_right_13),
	.a_right_14(a_right_14),
	.a_right_15(a_right_15),
	.a_right_16(a_right_16),
	.a_right_17(a_right_17),
	.a_right_18(a_right_18),
	.a_right_19(a_right_19),
	.a_right_20(a_right_20),
	.a_right_21(a_right_21),
	.a_right_22(a_right_22),
	.a_right_23(a_right_23),
	.a_right_24(a_right_24),
	.a_right_25(a_right_25),
	.a_right_26(a_right_26),
	.a_right_27(a_right_27),
	.a_right_28(a_right_28),
	.a_right_29(a_right_29),
	.a_right_30(a_right_30),
	.a_right_31(a_right_31),
	.a_right_32(a_right_32),
	.a_right_33(a_right_33),
	.a_right_34(a_right_34),
	.a_right_35(a_right_35),
	.a_right_36(a_right_36),
	.a_right_37(a_right_37),
	.a_right_38(a_right_38),
	.a_right_39(a_right_39),
	.a_right_40(a_right_40),
	.a_right_41(a_right_41),
	.a_right_42(a_right_42),
	.a_right_43(a_right_43),
	.a_right_44(a_right_44),
	.a_right_45(a_right_45),
	.a_right_46(a_right_46),
	.a_right_47(a_right_47),
	.a_right_48(a_right_48),
	.a_right_49(a_right_49),
	.a_right_50(a_right_50),
	.a_right_51(a_right_51),
	.a_right_52(a_right_52),
	.a_right_53(a_right_53),
	.a_right_54(a_right_54),
	.a_right_55(a_right_55),
	.a_right_56(a_right_56),
	.a_right_57(a_right_57),
	.a_right_58(a_right_58),
	.a_right_59(a_right_59),
	.a_right_60(a_right_60),
	.a_right_61(a_right_61),
	.a_right_62(a_right_62),
	.a_right_63(a_right_63),
	.a_right_64(a_right_64),
	.a_right_65(a_right_65),
	.a_right_66(a_right_66),
	.a_right_67(a_right_67),
	.a_right_68(a_right_68),
	.a_right_69(a_right_69),
	.a_right_70(a_right_70),
	.a_right_71(a_right_71),
	.a_right_72(a_right_72),
	.a_right_73(a_right_73),
	.a_right_74(a_right_74),
	.a_right_75(a_right_75),
	.a_right_76(a_right_76),
	.a_right_77(a_right_77),
	.a_right_78(a_right_78),
	.a_right_79(a_right_79),
	.a_right_80(a_right_80),
	.a_right_81(a_right_81),
	.a_right_82(a_right_82),
	.a_right_83(a_right_83),
	.a_right_84(a_right_84),
	.a_right_85(a_right_85),
	.a_right_86(a_right_86),
	.a_right_87(a_right_87),
	.a_right_88(a_right_88),
	.a_right_89(a_right_89),
	.a_right_90(a_right_90),
	.a_right_91(a_right_91),
	.a_right_92(a_right_92),
	.a_right_93(a_right_93),
	.a_right_94(a_right_94),
	.a_right_95(a_right_95),
	.a_right_96(a_right_96),
	.a_right_97(a_right_97),
	.a_right_98(a_right_98),
	.a_right_99(a_right_99),
	.a_right_100(a_right_100),
	.a_right_101(a_right_101),
	.a_right_102(a_right_102),
	.a_right_103(a_right_103),
	.a_right_104(a_right_104),
	.a_right_105(a_right_105),
	.a_right_106(a_right_106),
	.a_right_107(a_right_107),
	.a_right_108(a_right_108),
	.a_right_109(a_right_109),
	.a_right_110(a_right_110),
	.a_right_111(a_right_111),
	.a_right_112(a_right_112),
	.a_right_113(a_right_113),
	.a_right_114(a_right_114),
	.a_right_115(a_right_115),
	.a_right_116(a_right_116),
	.a_right_117(a_right_117),
	.a_right_118(a_right_118),
	.a_right_119(a_right_119),
	.a_right_120(a_right_120),
	.a_right_121(a_right_121),
	.a_right_122(a_right_122),
	.a_right_123(a_right_123),
	.a_right_124(a_right_124),
	.a_right_125(a_right_125),
	.a_right_126(a_right_126),
	.a_right_127(a_right_127),
	.a_right_128(a_right_128)
);

and_array and_array (
	.al(al),
	.a_left_1(a_left_1),
	.a_left_2(a_left_2),
	.a_left_3(a_left_3),
	.a_left_4(a_left_4),
	.a_left_5(a_left_5),
	.a_left_6(a_left_6),
	.a_left_7(a_left_7),
	.a_left_8(a_left_8),
	.a_left_9(a_left_9),
	.a_left_10(a_left_10),
	.a_left_11(a_left_11),
	.a_left_12(a_left_12),
	.a_left_13(a_left_13),
	.a_left_14(a_left_14),
	.a_left_15(a_left_15),
	.a_left_16(a_left_16),
	.a_left_17(a_left_17),
	.a_left_18(a_left_18),
	.a_left_19(a_left_19),
	.a_left_20(a_left_20),
	.a_left_21(a_left_21),
	.a_left_22(a_left_22),
	.a_left_23(a_left_23),
	.a_left_24(a_left_24),
	.a_left_25(a_left_25),
	.a_left_26(a_left_26),
	.a_left_27(a_left_27),
	.a_left_28(a_left_28),
	.a_left_29(a_left_29),
	.a_left_30(a_left_30),
	.a_left_31(a_left_31),
	.a_left_32(a_left_32),
	.a_left_33(a_left_33),
	.a_left_34(a_left_34),
	.a_left_35(a_left_35),
	.a_left_36(a_left_36),
	.a_left_37(a_left_37),
	.a_left_38(a_left_38),
	.a_left_39(a_left_39),
	.a_left_40(a_left_40),
	.a_left_41(a_left_41),
	.a_left_42(a_left_42),
	.a_left_43(a_left_43),
	.a_left_44(a_left_44),
	.a_left_45(a_left_45),
	.a_left_46(a_left_46),
	.a_left_47(a_left_47),
	.a_left_48(a_left_48),
	.a_left_49(a_left_49),
	.a_left_50(a_left_50),
	.a_left_51(a_left_51),
	.a_left_52(a_left_52),
	.a_left_53(a_left_53),
	.a_left_54(a_left_54),
	.a_left_55(a_left_55),
	.a_left_56(a_left_56),
	.a_left_57(a_left_57),
	.a_left_58(a_left_58),
	.a_left_59(a_left_59),
	.a_left_60(a_left_60),
	.a_left_61(a_left_61),
	.a_left_62(a_left_62),
	.a_left_63(a_left_63),
	.a_left_64(a_left_64),
	.a_left_65(a_left_65),
	.a_left_66(a_left_66),
	.a_left_67(a_left_67),
	.a_left_68(a_left_68),
	.a_left_69(a_left_69),
	.a_left_70(a_left_70),
	.a_left_71(a_left_71),
	.a_left_72(a_left_72),
	.a_left_73(a_left_73),
	.a_left_74(a_left_74),
	.a_left_75(a_left_75),
	.a_left_76(a_left_76),
	.a_left_77(a_left_77),
	.a_left_78(a_left_78),
	.a_left_79(a_left_79),
	.a_left_80(a_left_80),
	.a_left_81(a_left_81),
	.a_left_82(a_left_82),
	.a_left_83(a_left_83),
	.a_left_84(a_left_84),
	.a_left_85(a_left_85),
	.a_left_86(a_left_86),
	.a_left_87(a_left_87),
	.a_left_88(a_left_88),
	.a_left_89(a_left_89),
	.a_left_90(a_left_90),
	.a_left_91(a_left_91),
	.a_left_92(a_left_92),
	.a_left_93(a_left_93),
	.a_left_94(a_left_94),
	.a_left_95(a_left_95),
	.a_left_96(a_left_96),
	.a_left_97(a_left_97),
	.a_left_98(a_left_98),
	.a_left_99(a_left_99),
	.a_left_100(a_left_100),
	.a_left_101(a_left_101),
	.a_left_102(a_left_102),
	.a_left_103(a_left_103),
	.a_left_104(a_left_104),
	.a_left_105(a_left_105),
	.a_left_106(a_left_106),
	.a_left_107(a_left_107),
	.a_left_108(a_left_108),
	.a_left_109(a_left_109),
	.a_left_110(a_left_110),
	.a_left_111(a_left_111),
	.a_left_112(a_left_112),
	.a_left_113(a_left_113),
	.a_left_114(a_left_114),
	.a_left_115(a_left_115),
	.a_left_116(a_left_116),
	.a_left_117(a_left_117),
	.a_left_118(a_left_118),
	.a_left_119(a_left_119),
	.a_left_120(a_left_120),
	.a_left_121(a_left_121),
	.a_left_122(a_left_122),
	.a_left_123(a_left_123),
	.a_left_124(a_left_124),
	.a_left_125(a_left_125),
	.a_left_126(a_left_126),
	.a_left_127(a_left_127),
	.a_left_128(a_left_128),
	.a_right_1(a_right_1),
	.a_right_2(a_right_2),
	.a_right_3(a_right_3),
	.a_right_4(a_right_4),
	.a_right_5(a_right_5),
	.a_right_6(a_right_6),
	.a_right_7(a_right_7),
	.a_right_8(a_right_8),
	.a_right_9(a_right_9),
	.a_right_10(a_right_10),
	.a_right_11(a_right_11),
	.a_right_12(a_right_12),
	.a_right_13(a_right_13),
	.a_right_14(a_right_14),
	.a_right_15(a_right_15),
	.a_right_16(a_right_16),
	.a_right_17(a_right_17),
	.a_right_18(a_right_18),
	.a_right_19(a_right_19),
	.a_right_20(a_right_20),
	.a_right_21(a_right_21),
	.a_right_22(a_right_22),
	.a_right_23(a_right_23),
	.a_right_24(a_right_24),
	.a_right_25(a_right_25),
	.a_right_26(a_right_26),
	.a_right_27(a_right_27),
	.a_right_28(a_right_28),
	.a_right_29(a_right_29),
	.a_right_30(a_right_30),
	.a_right_31(a_right_31),
	.a_right_32(a_right_32),
	.a_right_33(a_right_33),
	.a_right_34(a_right_34),
	.a_right_35(a_right_35),
	.a_right_36(a_right_36),
	.a_right_37(a_right_37),
	.a_right_38(a_right_38),
	.a_right_39(a_right_39),
	.a_right_40(a_right_40),
	.a_right_41(a_right_41),
	.a_right_42(a_right_42),
	.a_right_43(a_right_43),
	.a_right_44(a_right_44),
	.a_right_45(a_right_45),
	.a_right_46(a_right_46),
	.a_right_47(a_right_47),
	.a_right_48(a_right_48),
	.a_right_49(a_right_49),
	.a_right_50(a_right_50),
	.a_right_51(a_right_51),
	.a_right_52(a_right_52),
	.a_right_53(a_right_53),
	.a_right_54(a_right_54),
	.a_right_55(a_right_55),
	.a_right_56(a_right_56),
	.a_right_57(a_right_57),
	.a_right_58(a_right_58),
	.a_right_59(a_right_59),
	.a_right_60(a_right_60),
	.a_right_61(a_right_61),
	.a_right_62(a_right_62),
	.a_right_63(a_right_63),
	.a_right_64(a_right_64),
	.a_right_65(a_right_65),
	.a_right_66(a_right_66),
	.a_right_67(a_right_67),
	.a_right_68(a_right_68),
	.a_right_69(a_right_69),
	.a_right_70(a_right_70),
	.a_right_71(a_right_71),
	.a_right_72(a_right_72),
	.a_right_73(a_right_73),
	.a_right_74(a_right_74),
	.a_right_75(a_right_75),
	.a_right_76(a_right_76),
	.a_right_77(a_right_77),
	.a_right_78(a_right_78),
	.a_right_79(a_right_79),
	.a_right_80(a_right_80),
	.a_right_81(a_right_81),
	.a_right_82(a_right_82),
	.a_right_83(a_right_83),
	.a_right_84(a_right_84),
	.a_right_85(a_right_85),
	.a_right_86(a_right_86),
	.a_right_87(a_right_87),
	.a_right_88(a_right_88),
	.a_right_89(a_right_89),
	.a_right_90(a_right_90),
	.a_right_91(a_right_91),
	.a_right_92(a_right_92),
	.a_right_93(a_right_93),
	.a_right_94(a_right_94),
	.a_right_95(a_right_95),
	.a_right_96(a_right_96),
	.a_right_97(a_right_97),
	.a_right_98(a_right_98),
	.a_right_99(a_right_99),
	.a_right_100(a_right_100),
	.a_right_101(a_right_101),
	.a_right_102(a_right_102),
	.a_right_103(a_right_103),
	.a_right_104(a_right_104),
	.a_right_105(a_right_105),
	.a_right_106(a_right_106),
	.a_right_107(a_right_107),
	.a_right_108(a_right_108),
	.a_right_109(a_right_109),
	.a_right_110(a_right_110),
	.a_right_111(a_right_111),
	.a_right_112(a_right_112),
	.a_right_113(a_right_113),
	.a_right_114(a_right_114),
	.a_right_115(a_right_115),
	.a_right_116(a_right_116),
	.a_right_117(a_right_117),
	.a_right_118(a_right_118),
	.a_right_119(a_right_119),
	.a_right_120(a_right_120),
	.a_right_121(a_right_121),
	.a_right_122(a_right_122),
	.a_right_123(a_right_123),
	.a_right_124(a_right_124),
	.a_right_125(a_right_125),
	.a_right_126(a_right_126),
	.a_right_127(a_right_127),
	.a_right_128(a_right_128),
	.line_1(line_1),
	.line_2(line_2),
	.line_3(line_3),
	.line_4(line_4),
	.line_5(line_5),
	.line_6(line_6),
	.line_7(line_7),
	.line_8(line_8),
	.line_9(line_9),
	.line_10(line_10),
	.line_11(line_11),
	.line_12(line_12),
	.line_13(line_13),
	.line_14(line_14),
	.line_15(line_15),
	.line_16(line_16),
	.line_17(line_17),
	.line_18(line_18),
	.line_19(line_19),
	.line_20(line_20),
	.line_21(line_21),
	.line_22(line_22),
	.line_23(line_23),
	.line_24(line_24),
	.line_25(line_25),
	.line_26(line_26),
	.line_27(line_27),
	.line_28(line_28),
	.line_29(line_29),
	.line_30(line_30),
	.line_31(line_31),
	.line_32(line_32),
	.line_33(line_33),
	.line_34(line_34),
	.line_35(line_35),
	.line_36(line_36),
	.line_37(line_37),
	.line_38(line_38),
	.line_39(line_39),
	.line_40(line_40),
	.line_41(line_41),
	.line_42(line_42),
	.line_43(line_43),
	.line_44(line_44),
	.line_45(line_45),
	.line_46(line_46),
	.line_47(line_47),
	.line_48(line_48),
	.line_49(line_49),
	.line_50(line_50),
	.line_51(line_51),
	.line_52(line_52),
	.line_53(line_53),
	.line_54(line_54),
	.line_55(line_55),
	.line_56(line_56),
	.line_57(line_57),
	.line_58(line_58),
	.line_59(line_59),
	.line_60(line_60),
	.line_61(line_61),
	.line_62(line_62),
	.line_63(line_63),
	.line_64(line_64),
	.line_65(line_65),
	.line_66(line_66),
	.line_67(line_67),
	.line_68(line_68),
	.line_69(line_69),
	.line_70(line_70),
	.line_71(line_71),
	.line_72(line_72),
	.line_73(line_73),
	.line_74(line_74),
	.line_75(line_75),
	.line_76(line_76),
	.line_77(line_77),
	.line_78(line_78),
	.line_79(line_79),
	.line_80(line_80),
	.line_81(line_81),
	.line_82(line_82),
	.line_83(line_83),
	.line_84(line_84),
	.line_85(line_85),
	.line_86(line_86),
	.line_87(line_87),
	.line_88(line_88),
	.line_89(line_89),
	.line_90(line_90),
	.line_91(line_91),
	.line_92(line_92),
	.line_93(line_93),
	.line_94(line_94),
	.line_95(line_95),
	.line_96(line_96),
	.line_97(line_97),
	.line_98(line_98),
	.line_99(line_99),
	.line_100(line_100),
	.line_101(line_101),
	.line_102(line_102),
	.line_103(line_103),
	.line_104(line_104),
	.line_105(line_105),
	.line_106(line_106),
	.line_107(line_107),
	.line_108(line_108),
	.line_109(line_109),
	.line_110(line_110),
	.line_111(line_111),
	.line_112(line_112),
	.line_113(line_113),
	.line_114(line_114),
	.line_115(line_115),
	.line_116(line_116),
	.line_117(line_117),
	.line_118(line_118),
	.line_119(line_119),
	.line_120(line_120),
	.line_121(line_121),
	.line_122(line_122),
	.line_123(line_123),
	.line_124(line_124),
	.line_125(line_125),
	.line_126(line_126),
	.line_127(line_127),
	.line_128(line_128)
);

assign col_0 = {line_128[0], 127'b0};
assign col_1 = {line_128[1], 127'b0};
assign col_2 = {line_128[2], line_127[0], 126'b0};
assign col_3 = {line_128[3], line_127[1], 126'b0};
assign col_4 = {line_128[4], line_127[2], line_126[0], 125'b0};
assign col_5 = {line_128[5], line_127[3], line_126[1], 125'b0};
assign col_6 = {line_128[6], line_127[4], line_126[2], line_125[0], 124'b0};
assign col_7 = {line_128[7], line_127[5], line_126[3], line_125[1], 124'b0};
assign col_8 = {line_128[8], line_127[6], line_126[4], line_125[2], line_124[0], 123'b0};
assign col_9 = {line_128[9], line_127[7], line_126[5], line_125[3], line_124[1], 123'b0};
assign col_10 = {line_128[10], line_127[8], line_126[6], line_125[4], line_124[2], line_123[0], 122'b0};
assign col_11 = {line_128[11], line_127[9], line_126[7], line_125[5], line_124[3], line_123[1], 122'b0};
assign col_12 = {line_128[12], line_127[10], line_126[8], line_125[6], line_124[4], line_123[2], line_122[0], 121'b0};
assign col_13 = {line_128[13], line_127[11], line_126[9], line_125[7], line_124[5], line_123[3], line_122[1], 121'b0};
assign col_14 = {line_128[14], line_127[12], line_126[10], line_125[8], line_124[6], line_123[4], line_122[2], line_121[0], 120'b0};
assign col_15 = {line_128[15], line_127[13], line_126[11], line_125[9], line_124[7], line_123[5], line_122[3], line_121[1], 120'b0};
assign col_16 = {line_128[16], line_127[14], line_126[12], line_125[10], line_124[8], line_123[6], line_122[4], line_121[2], line_120[0], 119'b0};
assign col_17 = {line_128[17], line_127[15], line_126[13], line_125[11], line_124[9], line_123[7], line_122[5], line_121[3], line_120[1], 119'b0};
assign col_18 = {line_128[18], line_127[16], line_126[14], line_125[12], line_124[10], line_123[8], line_122[6], line_121[4], line_120[2], line_119[0], 118'b0};
assign col_19 = {line_128[19], line_127[17], line_126[15], line_125[13], line_124[11], line_123[9], line_122[7], line_121[5], line_120[3], line_119[1], 118'b0};
assign col_20 = {line_128[20], line_127[18], line_126[16], line_125[14], line_124[12], line_123[10], line_122[8], line_121[6], line_120[4], line_119[2], line_118[0], 117'b0};
assign col_21 = {line_128[21], line_127[19], line_126[17], line_125[15], line_124[13], line_123[11], line_122[9], line_121[7], line_120[5], line_119[3], line_118[1], 117'b0};
assign col_22 = {line_128[22], line_127[20], line_126[18], line_125[16], line_124[14], line_123[12], line_122[10], line_121[8], line_120[6], line_119[4], line_118[2], line_117[0], 116'b0};
assign col_23 = {line_128[23], line_127[21], line_126[19], line_125[17], line_124[15], line_123[13], line_122[11], line_121[9], line_120[7], line_119[5], line_118[3], line_117[1], 116'b0};
assign col_24 = {line_128[24], line_127[22], line_126[20], line_125[18], line_124[16], line_123[14], line_122[12], line_121[10], line_120[8], line_119[6], line_118[4], line_117[2], line_116[0], 115'b0};
assign col_25 = {line_128[25], line_127[23], line_126[21], line_125[19], line_124[17], line_123[15], line_122[13], line_121[11], line_120[9], line_119[7], line_118[5], line_117[3], line_116[1], 115'b0};
assign col_26 = {line_128[26], line_127[24], line_126[22], line_125[20], line_124[18], line_123[16], line_122[14], line_121[12], line_120[10], line_119[8], line_118[6], line_117[4], line_116[2], line_115[0], 114'b0};
assign col_27 = {line_128[27], line_127[25], line_126[23], line_125[21], line_124[19], line_123[17], line_122[15], line_121[13], line_120[11], line_119[9], line_118[7], line_117[5], line_116[3], line_115[1], 114'b0};
assign col_28 = {line_128[28], line_127[26], line_126[24], line_125[22], line_124[20], line_123[18], line_122[16], line_121[14], line_120[12], line_119[10], line_118[8], line_117[6], line_116[4], line_115[2], line_114[0], 113'b0};
assign col_29 = {line_128[29], line_127[27], line_126[25], line_125[23], line_124[21], line_123[19], line_122[17], line_121[15], line_120[13], line_119[11], line_118[9], line_117[7], line_116[5], line_115[3], line_114[1], 113'b0};
assign col_30 = {line_128[30], line_127[28], line_126[26], line_125[24], line_124[22], line_123[20], line_122[18], line_121[16], line_120[14], line_119[12], line_118[10], line_117[8], line_116[6], line_115[4], line_114[2], line_113[0], 112'b0};
assign col_31 = {line_128[31], line_127[29], line_126[27], line_125[25], line_124[23], line_123[21], line_122[19], line_121[17], line_120[15], line_119[13], line_118[11], line_117[9], line_116[7], line_115[5], line_114[3], line_113[1], 112'b0};
assign col_32 = {line_128[32], line_127[30], line_126[28], line_125[26], line_124[24], line_123[22], line_122[20], line_121[18], line_120[16], line_119[14], line_118[12], line_117[10], line_116[8], line_115[6], line_114[4], line_113[2], line_112[0], 111'b0};
assign col_33 = {line_128[33], line_127[31], line_126[29], line_125[27], line_124[25], line_123[23], line_122[21], line_121[19], line_120[17], line_119[15], line_118[13], line_117[11], line_116[9], line_115[7], line_114[5], line_113[3], line_112[1], 111'b0};
assign col_34 = {line_128[34], line_127[32], line_126[30], line_125[28], line_124[26], line_123[24], line_122[22], line_121[20], line_120[18], line_119[16], line_118[14], line_117[12], line_116[10], line_115[8], line_114[6], line_113[4], line_112[2], line_111[0], 110'b0};
assign col_35 = {line_128[35], line_127[33], line_126[31], line_125[29], line_124[27], line_123[25], line_122[23], line_121[21], line_120[19], line_119[17], line_118[15], line_117[13], line_116[11], line_115[9], line_114[7], line_113[5], line_112[3], line_111[1], 110'b0};
assign col_36 = {line_128[36], line_127[34], line_126[32], line_125[30], line_124[28], line_123[26], line_122[24], line_121[22], line_120[20], line_119[18], line_118[16], line_117[14], line_116[12], line_115[10], line_114[8], line_113[6], line_112[4], line_111[2], line_110[0], 109'b0};
assign col_37 = {line_128[37], line_127[35], line_126[33], line_125[31], line_124[29], line_123[27], line_122[25], line_121[23], line_120[21], line_119[19], line_118[17], line_117[15], line_116[13], line_115[11], line_114[9], line_113[7], line_112[5], line_111[3], line_110[1], 109'b0};
assign col_38 = {line_128[38], line_127[36], line_126[34], line_125[32], line_124[30], line_123[28], line_122[26], line_121[24], line_120[22], line_119[20], line_118[18], line_117[16], line_116[14], line_115[12], line_114[10], line_113[8], line_112[6], line_111[4], line_110[2], line_109[0], 108'b0};
assign col_39 = {line_128[39], line_127[37], line_126[35], line_125[33], line_124[31], line_123[29], line_122[27], line_121[25], line_120[23], line_119[21], line_118[19], line_117[17], line_116[15], line_115[13], line_114[11], line_113[9], line_112[7], line_111[5], line_110[3], line_109[1], 108'b0};
assign col_40 = {line_128[40], line_127[38], line_126[36], line_125[34], line_124[32], line_123[30], line_122[28], line_121[26], line_120[24], line_119[22], line_118[20], line_117[18], line_116[16], line_115[14], line_114[12], line_113[10], line_112[8], line_111[6], line_110[4], line_109[2], line_108[0], 107'b0};
assign col_41 = {line_128[41], line_127[39], line_126[37], line_125[35], line_124[33], line_123[31], line_122[29], line_121[27], line_120[25], line_119[23], line_118[21], line_117[19], line_116[17], line_115[15], line_114[13], line_113[11], line_112[9], line_111[7], line_110[5], line_109[3], line_108[1], 107'b0};
assign col_42 = {line_128[42], line_127[40], line_126[38], line_125[36], line_124[34], line_123[32], line_122[30], line_121[28], line_120[26], line_119[24], line_118[22], line_117[20], line_116[18], line_115[16], line_114[14], line_113[12], line_112[10], line_111[8], line_110[6], line_109[4], line_108[2], line_107[0], 106'b0};
assign col_43 = {line_128[43], line_127[41], line_126[39], line_125[37], line_124[35], line_123[33], line_122[31], line_121[29], line_120[27], line_119[25], line_118[23], line_117[21], line_116[19], line_115[17], line_114[15], line_113[13], line_112[11], line_111[9], line_110[7], line_109[5], line_108[3], line_107[1], 106'b0};
assign col_44 = {line_128[44], line_127[42], line_126[40], line_125[38], line_124[36], line_123[34], line_122[32], line_121[30], line_120[28], line_119[26], line_118[24], line_117[22], line_116[20], line_115[18], line_114[16], line_113[14], line_112[12], line_111[10], line_110[8], line_109[6], line_108[4], line_107[2], line_106[0], 105'b0};
assign col_45 = {line_128[45], line_127[43], line_126[41], line_125[39], line_124[37], line_123[35], line_122[33], line_121[31], line_120[29], line_119[27], line_118[25], line_117[23], line_116[21], line_115[19], line_114[17], line_113[15], line_112[13], line_111[11], line_110[9], line_109[7], line_108[5], line_107[3], line_106[1], 105'b0};
assign col_46 = {line_128[46], line_127[44], line_126[42], line_125[40], line_124[38], line_123[36], line_122[34], line_121[32], line_120[30], line_119[28], line_118[26], line_117[24], line_116[22], line_115[20], line_114[18], line_113[16], line_112[14], line_111[12], line_110[10], line_109[8], line_108[6], line_107[4], line_106[2], line_105[0], 104'b0};
assign col_47 = {line_128[47], line_127[45], line_126[43], line_125[41], line_124[39], line_123[37], line_122[35], line_121[33], line_120[31], line_119[29], line_118[27], line_117[25], line_116[23], line_115[21], line_114[19], line_113[17], line_112[15], line_111[13], line_110[11], line_109[9], line_108[7], line_107[5], line_106[3], line_105[1], 104'b0};
assign col_48 = {line_128[48], line_127[46], line_126[44], line_125[42], line_124[40], line_123[38], line_122[36], line_121[34], line_120[32], line_119[30], line_118[28], line_117[26], line_116[24], line_115[22], line_114[20], line_113[18], line_112[16], line_111[14], line_110[12], line_109[10], line_108[8], line_107[6], line_106[4], line_105[2], line_104[0], 103'b0};
assign col_49 = {line_128[49], line_127[47], line_126[45], line_125[43], line_124[41], line_123[39], line_122[37], line_121[35], line_120[33], line_119[31], line_118[29], line_117[27], line_116[25], line_115[23], line_114[21], line_113[19], line_112[17], line_111[15], line_110[13], line_109[11], line_108[9], line_107[7], line_106[5], line_105[3], line_104[1], 103'b0};
assign col_50 = {line_128[50], line_127[48], line_126[46], line_125[44], line_124[42], line_123[40], line_122[38], line_121[36], line_120[34], line_119[32], line_118[30], line_117[28], line_116[26], line_115[24], line_114[22], line_113[20], line_112[18], line_111[16], line_110[14], line_109[12], line_108[10], line_107[8], line_106[6], line_105[4], line_104[2], line_103[0], 102'b0};
assign col_51 = {line_128[51], line_127[49], line_126[47], line_125[45], line_124[43], line_123[41], line_122[39], line_121[37], line_120[35], line_119[33], line_118[31], line_117[29], line_116[27], line_115[25], line_114[23], line_113[21], line_112[19], line_111[17], line_110[15], line_109[13], line_108[11], line_107[9], line_106[7], line_105[5], line_104[3], line_103[1], 102'b0};
assign col_52 = {line_128[52], line_127[50], line_126[48], line_125[46], line_124[44], line_123[42], line_122[40], line_121[38], line_120[36], line_119[34], line_118[32], line_117[30], line_116[28], line_115[26], line_114[24], line_113[22], line_112[20], line_111[18], line_110[16], line_109[14], line_108[12], line_107[10], line_106[8], line_105[6], line_104[4], line_103[2], line_102[0], 101'b0};
assign col_53 = {line_128[53], line_127[51], line_126[49], line_125[47], line_124[45], line_123[43], line_122[41], line_121[39], line_120[37], line_119[35], line_118[33], line_117[31], line_116[29], line_115[27], line_114[25], line_113[23], line_112[21], line_111[19], line_110[17], line_109[15], line_108[13], line_107[11], line_106[9], line_105[7], line_104[5], line_103[3], line_102[1], 101'b0};
assign col_54 = {line_128[54], line_127[52], line_126[50], line_125[48], line_124[46], line_123[44], line_122[42], line_121[40], line_120[38], line_119[36], line_118[34], line_117[32], line_116[30], line_115[28], line_114[26], line_113[24], line_112[22], line_111[20], line_110[18], line_109[16], line_108[14], line_107[12], line_106[10], line_105[8], line_104[6], line_103[4], line_102[2], line_101[0], 100'b0};
assign col_55 = {line_128[55], line_127[53], line_126[51], line_125[49], line_124[47], line_123[45], line_122[43], line_121[41], line_120[39], line_119[37], line_118[35], line_117[33], line_116[31], line_115[29], line_114[27], line_113[25], line_112[23], line_111[21], line_110[19], line_109[17], line_108[15], line_107[13], line_106[11], line_105[9], line_104[7], line_103[5], line_102[3], line_101[1], 100'b0};
assign col_56 = {line_128[56], line_127[54], line_126[52], line_125[50], line_124[48], line_123[46], line_122[44], line_121[42], line_120[40], line_119[38], line_118[36], line_117[34], line_116[32], line_115[30], line_114[28], line_113[26], line_112[24], line_111[22], line_110[20], line_109[18], line_108[16], line_107[14], line_106[12], line_105[10], line_104[8], line_103[6], line_102[4], line_101[2], line_100[0], 99'b0};
assign col_57 = {line_128[57], line_127[55], line_126[53], line_125[51], line_124[49], line_123[47], line_122[45], line_121[43], line_120[41], line_119[39], line_118[37], line_117[35], line_116[33], line_115[31], line_114[29], line_113[27], line_112[25], line_111[23], line_110[21], line_109[19], line_108[17], line_107[15], line_106[13], line_105[11], line_104[9], line_103[7], line_102[5], line_101[3], line_100[1], 99'b0};
assign col_58 = {line_128[58], line_127[56], line_126[54], line_125[52], line_124[50], line_123[48], line_122[46], line_121[44], line_120[42], line_119[40], line_118[38], line_117[36], line_116[34], line_115[32], line_114[30], line_113[28], line_112[26], line_111[24], line_110[22], line_109[20], line_108[18], line_107[16], line_106[14], line_105[12], line_104[10], line_103[8], line_102[6], line_101[4], line_100[2], line_99[0], 98'b0};
assign col_59 = {line_128[59], line_127[57], line_126[55], line_125[53], line_124[51], line_123[49], line_122[47], line_121[45], line_120[43], line_119[41], line_118[39], line_117[37], line_116[35], line_115[33], line_114[31], line_113[29], line_112[27], line_111[25], line_110[23], line_109[21], line_108[19], line_107[17], line_106[15], line_105[13], line_104[11], line_103[9], line_102[7], line_101[5], line_100[3], line_99[1], 98'b0};
assign col_60 = {line_128[60], line_127[58], line_126[56], line_125[54], line_124[52], line_123[50], line_122[48], line_121[46], line_120[44], line_119[42], line_118[40], line_117[38], line_116[36], line_115[34], line_114[32], line_113[30], line_112[28], line_111[26], line_110[24], line_109[22], line_108[20], line_107[18], line_106[16], line_105[14], line_104[12], line_103[10], line_102[8], line_101[6], line_100[4], line_99[2], line_98[0], 97'b0};
assign col_61 = {line_128[61], line_127[59], line_126[57], line_125[55], line_124[53], line_123[51], line_122[49], line_121[47], line_120[45], line_119[43], line_118[41], line_117[39], line_116[37], line_115[35], line_114[33], line_113[31], line_112[29], line_111[27], line_110[25], line_109[23], line_108[21], line_107[19], line_106[17], line_105[15], line_104[13], line_103[11], line_102[9], line_101[7], line_100[5], line_99[3], line_98[1], 97'b0};
assign col_62 = {line_128[62], line_127[60], line_126[58], line_125[56], line_124[54], line_123[52], line_122[50], line_121[48], line_120[46], line_119[44], line_118[42], line_117[40], line_116[38], line_115[36], line_114[34], line_113[32], line_112[30], line_111[28], line_110[26], line_109[24], line_108[22], line_107[20], line_106[18], line_105[16], line_104[14], line_103[12], line_102[10], line_101[8], line_100[6], line_99[4], line_98[2], line_97[0], 96'b0};
assign col_63 = {line_128[63], line_127[61], line_126[59], line_125[57], line_124[55], line_123[53], line_122[51], line_121[49], line_120[47], line_119[45], line_118[43], line_117[41], line_116[39], line_115[37], line_114[35], line_113[33], line_112[31], line_111[29], line_110[27], line_109[25], line_108[23], line_107[21], line_106[19], line_105[17], line_104[15], line_103[13], line_102[11], line_101[9], line_100[7], line_99[5], line_98[3], line_97[1], 96'b0};
assign col_64 = {line_128[64], line_127[62], line_126[60], line_125[58], line_124[56], line_123[54], line_122[52], line_121[50], line_120[48], line_119[46], line_118[44], line_117[42], line_116[40], line_115[38], line_114[36], line_113[34], line_112[32], line_111[30], line_110[28], line_109[26], line_108[24], line_107[22], line_106[20], line_105[18], line_104[16], line_103[14], line_102[12], line_101[10], line_100[8], line_99[6], line_98[4], line_97[2], line_96[0], 95'b0};
assign col_65 = {line_128[65], line_127[63], line_126[61], line_125[59], line_124[57], line_123[55], line_122[53], line_121[51], line_120[49], line_119[47], line_118[45], line_117[43], line_116[41], line_115[39], line_114[37], line_113[35], line_112[33], line_111[31], line_110[29], line_109[27], line_108[25], line_107[23], line_106[21], line_105[19], line_104[17], line_103[15], line_102[13], line_101[11], line_100[9], line_99[7], line_98[5], line_97[3], line_96[1], 95'b0};
assign col_66 = {line_128[66], line_127[64], line_126[62], line_125[60], line_124[58], line_123[56], line_122[54], line_121[52], line_120[50], line_119[48], line_118[46], line_117[44], line_116[42], line_115[40], line_114[38], line_113[36], line_112[34], line_111[32], line_110[30], line_109[28], line_108[26], line_107[24], line_106[22], line_105[20], line_104[18], line_103[16], line_102[14], line_101[12], line_100[10], line_99[8], line_98[6], line_97[4], line_96[2], line_95[0], 94'b0};
assign col_67 = {line_128[67], line_127[65], line_126[63], line_125[61], line_124[59], line_123[57], line_122[55], line_121[53], line_120[51], line_119[49], line_118[47], line_117[45], line_116[43], line_115[41], line_114[39], line_113[37], line_112[35], line_111[33], line_110[31], line_109[29], line_108[27], line_107[25], line_106[23], line_105[21], line_104[19], line_103[17], line_102[15], line_101[13], line_100[11], line_99[9], line_98[7], line_97[5], line_96[3], line_95[1], 94'b0};
assign col_68 = {line_128[68], line_127[66], line_126[64], line_125[62], line_124[60], line_123[58], line_122[56], line_121[54], line_120[52], line_119[50], line_118[48], line_117[46], line_116[44], line_115[42], line_114[40], line_113[38], line_112[36], line_111[34], line_110[32], line_109[30], line_108[28], line_107[26], line_106[24], line_105[22], line_104[20], line_103[18], line_102[16], line_101[14], line_100[12], line_99[10], line_98[8], line_97[6], line_96[4], line_95[2], line_94[0], 93'b0};
assign col_69 = {line_128[69], line_127[67], line_126[65], line_125[63], line_124[61], line_123[59], line_122[57], line_121[55], line_120[53], line_119[51], line_118[49], line_117[47], line_116[45], line_115[43], line_114[41], line_113[39], line_112[37], line_111[35], line_110[33], line_109[31], line_108[29], line_107[27], line_106[25], line_105[23], line_104[21], line_103[19], line_102[17], line_101[15], line_100[13], line_99[11], line_98[9], line_97[7], line_96[5], line_95[3], line_94[1], 93'b0};
assign col_70 = {line_128[70], line_127[68], line_126[66], line_125[64], line_124[62], line_123[60], line_122[58], line_121[56], line_120[54], line_119[52], line_118[50], line_117[48], line_116[46], line_115[44], line_114[42], line_113[40], line_112[38], line_111[36], line_110[34], line_109[32], line_108[30], line_107[28], line_106[26], line_105[24], line_104[22], line_103[20], line_102[18], line_101[16], line_100[14], line_99[12], line_98[10], line_97[8], line_96[6], line_95[4], line_94[2], line_93[0], 92'b0};
assign col_71 = {line_128[71], line_127[69], line_126[67], line_125[65], line_124[63], line_123[61], line_122[59], line_121[57], line_120[55], line_119[53], line_118[51], line_117[49], line_116[47], line_115[45], line_114[43], line_113[41], line_112[39], line_111[37], line_110[35], line_109[33], line_108[31], line_107[29], line_106[27], line_105[25], line_104[23], line_103[21], line_102[19], line_101[17], line_100[15], line_99[13], line_98[11], line_97[9], line_96[7], line_95[5], line_94[3], line_93[1], 92'b0};
assign col_72 = {line_128[72], line_127[70], line_126[68], line_125[66], line_124[64], line_123[62], line_122[60], line_121[58], line_120[56], line_119[54], line_118[52], line_117[50], line_116[48], line_115[46], line_114[44], line_113[42], line_112[40], line_111[38], line_110[36], line_109[34], line_108[32], line_107[30], line_106[28], line_105[26], line_104[24], line_103[22], line_102[20], line_101[18], line_100[16], line_99[14], line_98[12], line_97[10], line_96[8], line_95[6], line_94[4], line_93[2], line_92[0], 91'b0};
assign col_73 = {line_128[73], line_127[71], line_126[69], line_125[67], line_124[65], line_123[63], line_122[61], line_121[59], line_120[57], line_119[55], line_118[53], line_117[51], line_116[49], line_115[47], line_114[45], line_113[43], line_112[41], line_111[39], line_110[37], line_109[35], line_108[33], line_107[31], line_106[29], line_105[27], line_104[25], line_103[23], line_102[21], line_101[19], line_100[17], line_99[15], line_98[13], line_97[11], line_96[9], line_95[7], line_94[5], line_93[3], line_92[1], 91'b0};
assign col_74 = {line_128[74], line_127[72], line_126[70], line_125[68], line_124[66], line_123[64], line_122[62], line_121[60], line_120[58], line_119[56], line_118[54], line_117[52], line_116[50], line_115[48], line_114[46], line_113[44], line_112[42], line_111[40], line_110[38], line_109[36], line_108[34], line_107[32], line_106[30], line_105[28], line_104[26], line_103[24], line_102[22], line_101[20], line_100[18], line_99[16], line_98[14], line_97[12], line_96[10], line_95[8], line_94[6], line_93[4], line_92[2], line_91[0], 90'b0};
assign col_75 = {line_128[75], line_127[73], line_126[71], line_125[69], line_124[67], line_123[65], line_122[63], line_121[61], line_120[59], line_119[57], line_118[55], line_117[53], line_116[51], line_115[49], line_114[47], line_113[45], line_112[43], line_111[41], line_110[39], line_109[37], line_108[35], line_107[33], line_106[31], line_105[29], line_104[27], line_103[25], line_102[23], line_101[21], line_100[19], line_99[17], line_98[15], line_97[13], line_96[11], line_95[9], line_94[7], line_93[5], line_92[3], line_91[1], 90'b0};
assign col_76 = {line_128[76], line_127[74], line_126[72], line_125[70], line_124[68], line_123[66], line_122[64], line_121[62], line_120[60], line_119[58], line_118[56], line_117[54], line_116[52], line_115[50], line_114[48], line_113[46], line_112[44], line_111[42], line_110[40], line_109[38], line_108[36], line_107[34], line_106[32], line_105[30], line_104[28], line_103[26], line_102[24], line_101[22], line_100[20], line_99[18], line_98[16], line_97[14], line_96[12], line_95[10], line_94[8], line_93[6], line_92[4], line_91[2], line_90[0], 89'b0};
assign col_77 = {line_128[77], line_127[75], line_126[73], line_125[71], line_124[69], line_123[67], line_122[65], line_121[63], line_120[61], line_119[59], line_118[57], line_117[55], line_116[53], line_115[51], line_114[49], line_113[47], line_112[45], line_111[43], line_110[41], line_109[39], line_108[37], line_107[35], line_106[33], line_105[31], line_104[29], line_103[27], line_102[25], line_101[23], line_100[21], line_99[19], line_98[17], line_97[15], line_96[13], line_95[11], line_94[9], line_93[7], line_92[5], line_91[3], line_90[1], 89'b0};
assign col_78 = {line_128[78], line_127[76], line_126[74], line_125[72], line_124[70], line_123[68], line_122[66], line_121[64], line_120[62], line_119[60], line_118[58], line_117[56], line_116[54], line_115[52], line_114[50], line_113[48], line_112[46], line_111[44], line_110[42], line_109[40], line_108[38], line_107[36], line_106[34], line_105[32], line_104[30], line_103[28], line_102[26], line_101[24], line_100[22], line_99[20], line_98[18], line_97[16], line_96[14], line_95[12], line_94[10], line_93[8], line_92[6], line_91[4], line_90[2], line_89[0], 88'b0};
assign col_79 = {line_128[79], line_127[77], line_126[75], line_125[73], line_124[71], line_123[69], line_122[67], line_121[65], line_120[63], line_119[61], line_118[59], line_117[57], line_116[55], line_115[53], line_114[51], line_113[49], line_112[47], line_111[45], line_110[43], line_109[41], line_108[39], line_107[37], line_106[35], line_105[33], line_104[31], line_103[29], line_102[27], line_101[25], line_100[23], line_99[21], line_98[19], line_97[17], line_96[15], line_95[13], line_94[11], line_93[9], line_92[7], line_91[5], line_90[3], line_89[1], 88'b0};
assign col_80 = {line_128[80], line_127[78], line_126[76], line_125[74], line_124[72], line_123[70], line_122[68], line_121[66], line_120[64], line_119[62], line_118[60], line_117[58], line_116[56], line_115[54], line_114[52], line_113[50], line_112[48], line_111[46], line_110[44], line_109[42], line_108[40], line_107[38], line_106[36], line_105[34], line_104[32], line_103[30], line_102[28], line_101[26], line_100[24], line_99[22], line_98[20], line_97[18], line_96[16], line_95[14], line_94[12], line_93[10], line_92[8], line_91[6], line_90[4], line_89[2], line_88[0], 87'b0};
assign col_81 = {line_128[81], line_127[79], line_126[77], line_125[75], line_124[73], line_123[71], line_122[69], line_121[67], line_120[65], line_119[63], line_118[61], line_117[59], line_116[57], line_115[55], line_114[53], line_113[51], line_112[49], line_111[47], line_110[45], line_109[43], line_108[41], line_107[39], line_106[37], line_105[35], line_104[33], line_103[31], line_102[29], line_101[27], line_100[25], line_99[23], line_98[21], line_97[19], line_96[17], line_95[15], line_94[13], line_93[11], line_92[9], line_91[7], line_90[5], line_89[3], line_88[1], 87'b0};
assign col_82 = {line_128[82], line_127[80], line_126[78], line_125[76], line_124[74], line_123[72], line_122[70], line_121[68], line_120[66], line_119[64], line_118[62], line_117[60], line_116[58], line_115[56], line_114[54], line_113[52], line_112[50], line_111[48], line_110[46], line_109[44], line_108[42], line_107[40], line_106[38], line_105[36], line_104[34], line_103[32], line_102[30], line_101[28], line_100[26], line_99[24], line_98[22], line_97[20], line_96[18], line_95[16], line_94[14], line_93[12], line_92[10], line_91[8], line_90[6], line_89[4], line_88[2], line_87[0], 86'b0};
assign col_83 = {line_128[83], line_127[81], line_126[79], line_125[77], line_124[75], line_123[73], line_122[71], line_121[69], line_120[67], line_119[65], line_118[63], line_117[61], line_116[59], line_115[57], line_114[55], line_113[53], line_112[51], line_111[49], line_110[47], line_109[45], line_108[43], line_107[41], line_106[39], line_105[37], line_104[35], line_103[33], line_102[31], line_101[29], line_100[27], line_99[25], line_98[23], line_97[21], line_96[19], line_95[17], line_94[15], line_93[13], line_92[11], line_91[9], line_90[7], line_89[5], line_88[3], line_87[1], 86'b0};
assign col_84 = {line_128[84], line_127[82], line_126[80], line_125[78], line_124[76], line_123[74], line_122[72], line_121[70], line_120[68], line_119[66], line_118[64], line_117[62], line_116[60], line_115[58], line_114[56], line_113[54], line_112[52], line_111[50], line_110[48], line_109[46], line_108[44], line_107[42], line_106[40], line_105[38], line_104[36], line_103[34], line_102[32], line_101[30], line_100[28], line_99[26], line_98[24], line_97[22], line_96[20], line_95[18], line_94[16], line_93[14], line_92[12], line_91[10], line_90[8], line_89[6], line_88[4], line_87[2], line_86[0], 85'b0};
assign col_85 = {line_128[85], line_127[83], line_126[81], line_125[79], line_124[77], line_123[75], line_122[73], line_121[71], line_120[69], line_119[67], line_118[65], line_117[63], line_116[61], line_115[59], line_114[57], line_113[55], line_112[53], line_111[51], line_110[49], line_109[47], line_108[45], line_107[43], line_106[41], line_105[39], line_104[37], line_103[35], line_102[33], line_101[31], line_100[29], line_99[27], line_98[25], line_97[23], line_96[21], line_95[19], line_94[17], line_93[15], line_92[13], line_91[11], line_90[9], line_89[7], line_88[5], line_87[3], line_86[1], 85'b0};
assign col_86 = {line_128[86], line_127[84], line_126[82], line_125[80], line_124[78], line_123[76], line_122[74], line_121[72], line_120[70], line_119[68], line_118[66], line_117[64], line_116[62], line_115[60], line_114[58], line_113[56], line_112[54], line_111[52], line_110[50], line_109[48], line_108[46], line_107[44], line_106[42], line_105[40], line_104[38], line_103[36], line_102[34], line_101[32], line_100[30], line_99[28], line_98[26], line_97[24], line_96[22], line_95[20], line_94[18], line_93[16], line_92[14], line_91[12], line_90[10], line_89[8], line_88[6], line_87[4], line_86[2], line_85[0], 84'b0};
assign col_87 = {line_128[87], line_127[85], line_126[83], line_125[81], line_124[79], line_123[77], line_122[75], line_121[73], line_120[71], line_119[69], line_118[67], line_117[65], line_116[63], line_115[61], line_114[59], line_113[57], line_112[55], line_111[53], line_110[51], line_109[49], line_108[47], line_107[45], line_106[43], line_105[41], line_104[39], line_103[37], line_102[35], line_101[33], line_100[31], line_99[29], line_98[27], line_97[25], line_96[23], line_95[21], line_94[19], line_93[17], line_92[15], line_91[13], line_90[11], line_89[9], line_88[7], line_87[5], line_86[3], line_85[1], 84'b0};
assign col_88 = {line_128[88], line_127[86], line_126[84], line_125[82], line_124[80], line_123[78], line_122[76], line_121[74], line_120[72], line_119[70], line_118[68], line_117[66], line_116[64], line_115[62], line_114[60], line_113[58], line_112[56], line_111[54], line_110[52], line_109[50], line_108[48], line_107[46], line_106[44], line_105[42], line_104[40], line_103[38], line_102[36], line_101[34], line_100[32], line_99[30], line_98[28], line_97[26], line_96[24], line_95[22], line_94[20], line_93[18], line_92[16], line_91[14], line_90[12], line_89[10], line_88[8], line_87[6], line_86[4], line_85[2], line_84[0], 83'b0};
assign col_89 = {line_128[89], line_127[87], line_126[85], line_125[83], line_124[81], line_123[79], line_122[77], line_121[75], line_120[73], line_119[71], line_118[69], line_117[67], line_116[65], line_115[63], line_114[61], line_113[59], line_112[57], line_111[55], line_110[53], line_109[51], line_108[49], line_107[47], line_106[45], line_105[43], line_104[41], line_103[39], line_102[37], line_101[35], line_100[33], line_99[31], line_98[29], line_97[27], line_96[25], line_95[23], line_94[21], line_93[19], line_92[17], line_91[15], line_90[13], line_89[11], line_88[9], line_87[7], line_86[5], line_85[3], line_84[1], 83'b0};
assign col_90 = {line_128[90], line_127[88], line_126[86], line_125[84], line_124[82], line_123[80], line_122[78], line_121[76], line_120[74], line_119[72], line_118[70], line_117[68], line_116[66], line_115[64], line_114[62], line_113[60], line_112[58], line_111[56], line_110[54], line_109[52], line_108[50], line_107[48], line_106[46], line_105[44], line_104[42], line_103[40], line_102[38], line_101[36], line_100[34], line_99[32], line_98[30], line_97[28], line_96[26], line_95[24], line_94[22], line_93[20], line_92[18], line_91[16], line_90[14], line_89[12], line_88[10], line_87[8], line_86[6], line_85[4], line_84[2], line_83[0], 82'b0};
assign col_91 = {line_128[91], line_127[89], line_126[87], line_125[85], line_124[83], line_123[81], line_122[79], line_121[77], line_120[75], line_119[73], line_118[71], line_117[69], line_116[67], line_115[65], line_114[63], line_113[61], line_112[59], line_111[57], line_110[55], line_109[53], line_108[51], line_107[49], line_106[47], line_105[45], line_104[43], line_103[41], line_102[39], line_101[37], line_100[35], line_99[33], line_98[31], line_97[29], line_96[27], line_95[25], line_94[23], line_93[21], line_92[19], line_91[17], line_90[15], line_89[13], line_88[11], line_87[9], line_86[7], line_85[5], line_84[3], line_83[1], 82'b0};
assign col_92 = {line_128[92], line_127[90], line_126[88], line_125[86], line_124[84], line_123[82], line_122[80], line_121[78], line_120[76], line_119[74], line_118[72], line_117[70], line_116[68], line_115[66], line_114[64], line_113[62], line_112[60], line_111[58], line_110[56], line_109[54], line_108[52], line_107[50], line_106[48], line_105[46], line_104[44], line_103[42], line_102[40], line_101[38], line_100[36], line_99[34], line_98[32], line_97[30], line_96[28], line_95[26], line_94[24], line_93[22], line_92[20], line_91[18], line_90[16], line_89[14], line_88[12], line_87[10], line_86[8], line_85[6], line_84[4], line_83[2], line_82[0], 81'b0};
assign col_93 = {line_128[93], line_127[91], line_126[89], line_125[87], line_124[85], line_123[83], line_122[81], line_121[79], line_120[77], line_119[75], line_118[73], line_117[71], line_116[69], line_115[67], line_114[65], line_113[63], line_112[61], line_111[59], line_110[57], line_109[55], line_108[53], line_107[51], line_106[49], line_105[47], line_104[45], line_103[43], line_102[41], line_101[39], line_100[37], line_99[35], line_98[33], line_97[31], line_96[29], line_95[27], line_94[25], line_93[23], line_92[21], line_91[19], line_90[17], line_89[15], line_88[13], line_87[11], line_86[9], line_85[7], line_84[5], line_83[3], line_82[1], 81'b0};
assign col_94 = {line_128[94], line_127[92], line_126[90], line_125[88], line_124[86], line_123[84], line_122[82], line_121[80], line_120[78], line_119[76], line_118[74], line_117[72], line_116[70], line_115[68], line_114[66], line_113[64], line_112[62], line_111[60], line_110[58], line_109[56], line_108[54], line_107[52], line_106[50], line_105[48], line_104[46], line_103[44], line_102[42], line_101[40], line_100[38], line_99[36], line_98[34], line_97[32], line_96[30], line_95[28], line_94[26], line_93[24], line_92[22], line_91[20], line_90[18], line_89[16], line_88[14], line_87[12], line_86[10], line_85[8], line_84[6], line_83[4], line_82[2], line_81[0], 80'b0};
assign col_95 = {line_128[95], line_127[93], line_126[91], line_125[89], line_124[87], line_123[85], line_122[83], line_121[81], line_120[79], line_119[77], line_118[75], line_117[73], line_116[71], line_115[69], line_114[67], line_113[65], line_112[63], line_111[61], line_110[59], line_109[57], line_108[55], line_107[53], line_106[51], line_105[49], line_104[47], line_103[45], line_102[43], line_101[41], line_100[39], line_99[37], line_98[35], line_97[33], line_96[31], line_95[29], line_94[27], line_93[25], line_92[23], line_91[21], line_90[19], line_89[17], line_88[15], line_87[13], line_86[11], line_85[9], line_84[7], line_83[5], line_82[3], line_81[1], 80'b0};
assign col_96 = {line_128[96], line_127[94], line_126[92], line_125[90], line_124[88], line_123[86], line_122[84], line_121[82], line_120[80], line_119[78], line_118[76], line_117[74], line_116[72], line_115[70], line_114[68], line_113[66], line_112[64], line_111[62], line_110[60], line_109[58], line_108[56], line_107[54], line_106[52], line_105[50], line_104[48], line_103[46], line_102[44], line_101[42], line_100[40], line_99[38], line_98[36], line_97[34], line_96[32], line_95[30], line_94[28], line_93[26], line_92[24], line_91[22], line_90[20], line_89[18], line_88[16], line_87[14], line_86[12], line_85[10], line_84[8], line_83[6], line_82[4], line_81[2], line_80[0], 79'b0};
assign col_97 = {line_128[97], line_127[95], line_126[93], line_125[91], line_124[89], line_123[87], line_122[85], line_121[83], line_120[81], line_119[79], line_118[77], line_117[75], line_116[73], line_115[71], line_114[69], line_113[67], line_112[65], line_111[63], line_110[61], line_109[59], line_108[57], line_107[55], line_106[53], line_105[51], line_104[49], line_103[47], line_102[45], line_101[43], line_100[41], line_99[39], line_98[37], line_97[35], line_96[33], line_95[31], line_94[29], line_93[27], line_92[25], line_91[23], line_90[21], line_89[19], line_88[17], line_87[15], line_86[13], line_85[11], line_84[9], line_83[7], line_82[5], line_81[3], line_80[1], 79'b0};
assign col_98 = {line_128[98], line_127[96], line_126[94], line_125[92], line_124[90], line_123[88], line_122[86], line_121[84], line_120[82], line_119[80], line_118[78], line_117[76], line_116[74], line_115[72], line_114[70], line_113[68], line_112[66], line_111[64], line_110[62], line_109[60], line_108[58], line_107[56], line_106[54], line_105[52], line_104[50], line_103[48], line_102[46], line_101[44], line_100[42], line_99[40], line_98[38], line_97[36], line_96[34], line_95[32], line_94[30], line_93[28], line_92[26], line_91[24], line_90[22], line_89[20], line_88[18], line_87[16], line_86[14], line_85[12], line_84[10], line_83[8], line_82[6], line_81[4], line_80[2], line_79[0], 78'b0};
assign col_99 = {line_128[99], line_127[97], line_126[95], line_125[93], line_124[91], line_123[89], line_122[87], line_121[85], line_120[83], line_119[81], line_118[79], line_117[77], line_116[75], line_115[73], line_114[71], line_113[69], line_112[67], line_111[65], line_110[63], line_109[61], line_108[59], line_107[57], line_106[55], line_105[53], line_104[51], line_103[49], line_102[47], line_101[45], line_100[43], line_99[41], line_98[39], line_97[37], line_96[35], line_95[33], line_94[31], line_93[29], line_92[27], line_91[25], line_90[23], line_89[21], line_88[19], line_87[17], line_86[15], line_85[13], line_84[11], line_83[9], line_82[7], line_81[5], line_80[3], line_79[1], 78'b0};
assign col_100 = {line_128[100], line_127[98], line_126[96], line_125[94], line_124[92], line_123[90], line_122[88], line_121[86], line_120[84], line_119[82], line_118[80], line_117[78], line_116[76], line_115[74], line_114[72], line_113[70], line_112[68], line_111[66], line_110[64], line_109[62], line_108[60], line_107[58], line_106[56], line_105[54], line_104[52], line_103[50], line_102[48], line_101[46], line_100[44], line_99[42], line_98[40], line_97[38], line_96[36], line_95[34], line_94[32], line_93[30], line_92[28], line_91[26], line_90[24], line_89[22], line_88[20], line_87[18], line_86[16], line_85[14], line_84[12], line_83[10], line_82[8], line_81[6], line_80[4], line_79[2], line_78[0], 77'b0};
assign col_101 = {line_128[101], line_127[99], line_126[97], line_125[95], line_124[93], line_123[91], line_122[89], line_121[87], line_120[85], line_119[83], line_118[81], line_117[79], line_116[77], line_115[75], line_114[73], line_113[71], line_112[69], line_111[67], line_110[65], line_109[63], line_108[61], line_107[59], line_106[57], line_105[55], line_104[53], line_103[51], line_102[49], line_101[47], line_100[45], line_99[43], line_98[41], line_97[39], line_96[37], line_95[35], line_94[33], line_93[31], line_92[29], line_91[27], line_90[25], line_89[23], line_88[21], line_87[19], line_86[17], line_85[15], line_84[13], line_83[11], line_82[9], line_81[7], line_80[5], line_79[3], line_78[1], 77'b0};
assign col_102 = {line_128[102], line_127[100], line_126[98], line_125[96], line_124[94], line_123[92], line_122[90], line_121[88], line_120[86], line_119[84], line_118[82], line_117[80], line_116[78], line_115[76], line_114[74], line_113[72], line_112[70], line_111[68], line_110[66], line_109[64], line_108[62], line_107[60], line_106[58], line_105[56], line_104[54], line_103[52], line_102[50], line_101[48], line_100[46], line_99[44], line_98[42], line_97[40], line_96[38], line_95[36], line_94[34], line_93[32], line_92[30], line_91[28], line_90[26], line_89[24], line_88[22], line_87[20], line_86[18], line_85[16], line_84[14], line_83[12], line_82[10], line_81[8], line_80[6], line_79[4], line_78[2], line_77[0], 76'b0};
assign col_103 = {line_128[103], line_127[101], line_126[99], line_125[97], line_124[95], line_123[93], line_122[91], line_121[89], line_120[87], line_119[85], line_118[83], line_117[81], line_116[79], line_115[77], line_114[75], line_113[73], line_112[71], line_111[69], line_110[67], line_109[65], line_108[63], line_107[61], line_106[59], line_105[57], line_104[55], line_103[53], line_102[51], line_101[49], line_100[47], line_99[45], line_98[43], line_97[41], line_96[39], line_95[37], line_94[35], line_93[33], line_92[31], line_91[29], line_90[27], line_89[25], line_88[23], line_87[21], line_86[19], line_85[17], line_84[15], line_83[13], line_82[11], line_81[9], line_80[7], line_79[5], line_78[3], line_77[1], 76'b0};
assign col_104 = {line_128[104], line_127[102], line_126[100], line_125[98], line_124[96], line_123[94], line_122[92], line_121[90], line_120[88], line_119[86], line_118[84], line_117[82], line_116[80], line_115[78], line_114[76], line_113[74], line_112[72], line_111[70], line_110[68], line_109[66], line_108[64], line_107[62], line_106[60], line_105[58], line_104[56], line_103[54], line_102[52], line_101[50], line_100[48], line_99[46], line_98[44], line_97[42], line_96[40], line_95[38], line_94[36], line_93[34], line_92[32], line_91[30], line_90[28], line_89[26], line_88[24], line_87[22], line_86[20], line_85[18], line_84[16], line_83[14], line_82[12], line_81[10], line_80[8], line_79[6], line_78[4], line_77[2], line_76[0], 75'b0};
assign col_105 = {line_128[105], line_127[103], line_126[101], line_125[99], line_124[97], line_123[95], line_122[93], line_121[91], line_120[89], line_119[87], line_118[85], line_117[83], line_116[81], line_115[79], line_114[77], line_113[75], line_112[73], line_111[71], line_110[69], line_109[67], line_108[65], line_107[63], line_106[61], line_105[59], line_104[57], line_103[55], line_102[53], line_101[51], line_100[49], line_99[47], line_98[45], line_97[43], line_96[41], line_95[39], line_94[37], line_93[35], line_92[33], line_91[31], line_90[29], line_89[27], line_88[25], line_87[23], line_86[21], line_85[19], line_84[17], line_83[15], line_82[13], line_81[11], line_80[9], line_79[7], line_78[5], line_77[3], line_76[1], 75'b0};
assign col_106 = {line_128[106], line_127[104], line_126[102], line_125[100], line_124[98], line_123[96], line_122[94], line_121[92], line_120[90], line_119[88], line_118[86], line_117[84], line_116[82], line_115[80], line_114[78], line_113[76], line_112[74], line_111[72], line_110[70], line_109[68], line_108[66], line_107[64], line_106[62], line_105[60], line_104[58], line_103[56], line_102[54], line_101[52], line_100[50], line_99[48], line_98[46], line_97[44], line_96[42], line_95[40], line_94[38], line_93[36], line_92[34], line_91[32], line_90[30], line_89[28], line_88[26], line_87[24], line_86[22], line_85[20], line_84[18], line_83[16], line_82[14], line_81[12], line_80[10], line_79[8], line_78[6], line_77[4], line_76[2], line_75[0], 74'b0};
assign col_107 = {line_128[107], line_127[105], line_126[103], line_125[101], line_124[99], line_123[97], line_122[95], line_121[93], line_120[91], line_119[89], line_118[87], line_117[85], line_116[83], line_115[81], line_114[79], line_113[77], line_112[75], line_111[73], line_110[71], line_109[69], line_108[67], line_107[65], line_106[63], line_105[61], line_104[59], line_103[57], line_102[55], line_101[53], line_100[51], line_99[49], line_98[47], line_97[45], line_96[43], line_95[41], line_94[39], line_93[37], line_92[35], line_91[33], line_90[31], line_89[29], line_88[27], line_87[25], line_86[23], line_85[21], line_84[19], line_83[17], line_82[15], line_81[13], line_80[11], line_79[9], line_78[7], line_77[5], line_76[3], line_75[1], 74'b0};
assign col_108 = {line_128[108], line_127[106], line_126[104], line_125[102], line_124[100], line_123[98], line_122[96], line_121[94], line_120[92], line_119[90], line_118[88], line_117[86], line_116[84], line_115[82], line_114[80], line_113[78], line_112[76], line_111[74], line_110[72], line_109[70], line_108[68], line_107[66], line_106[64], line_105[62], line_104[60], line_103[58], line_102[56], line_101[54], line_100[52], line_99[50], line_98[48], line_97[46], line_96[44], line_95[42], line_94[40], line_93[38], line_92[36], line_91[34], line_90[32], line_89[30], line_88[28], line_87[26], line_86[24], line_85[22], line_84[20], line_83[18], line_82[16], line_81[14], line_80[12], line_79[10], line_78[8], line_77[6], line_76[4], line_75[2], line_74[0], 73'b0};
assign col_109 = {line_128[109], line_127[107], line_126[105], line_125[103], line_124[101], line_123[99], line_122[97], line_121[95], line_120[93], line_119[91], line_118[89], line_117[87], line_116[85], line_115[83], line_114[81], line_113[79], line_112[77], line_111[75], line_110[73], line_109[71], line_108[69], line_107[67], line_106[65], line_105[63], line_104[61], line_103[59], line_102[57], line_101[55], line_100[53], line_99[51], line_98[49], line_97[47], line_96[45], line_95[43], line_94[41], line_93[39], line_92[37], line_91[35], line_90[33], line_89[31], line_88[29], line_87[27], line_86[25], line_85[23], line_84[21], line_83[19], line_82[17], line_81[15], line_80[13], line_79[11], line_78[9], line_77[7], line_76[5], line_75[3], line_74[1], 73'b0};
assign col_110 = {line_128[110], line_127[108], line_126[106], line_125[104], line_124[102], line_123[100], line_122[98], line_121[96], line_120[94], line_119[92], line_118[90], line_117[88], line_116[86], line_115[84], line_114[82], line_113[80], line_112[78], line_111[76], line_110[74], line_109[72], line_108[70], line_107[68], line_106[66], line_105[64], line_104[62], line_103[60], line_102[58], line_101[56], line_100[54], line_99[52], line_98[50], line_97[48], line_96[46], line_95[44], line_94[42], line_93[40], line_92[38], line_91[36], line_90[34], line_89[32], line_88[30], line_87[28], line_86[26], line_85[24], line_84[22], line_83[20], line_82[18], line_81[16], line_80[14], line_79[12], line_78[10], line_77[8], line_76[6], line_75[4], line_74[2], line_73[0], 72'b0};
assign col_111 = {line_128[111], line_127[109], line_126[107], line_125[105], line_124[103], line_123[101], line_122[99], line_121[97], line_120[95], line_119[93], line_118[91], line_117[89], line_116[87], line_115[85], line_114[83], line_113[81], line_112[79], line_111[77], line_110[75], line_109[73], line_108[71], line_107[69], line_106[67], line_105[65], line_104[63], line_103[61], line_102[59], line_101[57], line_100[55], line_99[53], line_98[51], line_97[49], line_96[47], line_95[45], line_94[43], line_93[41], line_92[39], line_91[37], line_90[35], line_89[33], line_88[31], line_87[29], line_86[27], line_85[25], line_84[23], line_83[21], line_82[19], line_81[17], line_80[15], line_79[13], line_78[11], line_77[9], line_76[7], line_75[5], line_74[3], line_73[1], 72'b0};
assign col_112 = {line_128[112], line_127[110], line_126[108], line_125[106], line_124[104], line_123[102], line_122[100], line_121[98], line_120[96], line_119[94], line_118[92], line_117[90], line_116[88], line_115[86], line_114[84], line_113[82], line_112[80], line_111[78], line_110[76], line_109[74], line_108[72], line_107[70], line_106[68], line_105[66], line_104[64], line_103[62], line_102[60], line_101[58], line_100[56], line_99[54], line_98[52], line_97[50], line_96[48], line_95[46], line_94[44], line_93[42], line_92[40], line_91[38], line_90[36], line_89[34], line_88[32], line_87[30], line_86[28], line_85[26], line_84[24], line_83[22], line_82[20], line_81[18], line_80[16], line_79[14], line_78[12], line_77[10], line_76[8], line_75[6], line_74[4], line_73[2], line_72[0], 71'b0};
assign col_113 = {line_128[113], line_127[111], line_126[109], line_125[107], line_124[105], line_123[103], line_122[101], line_121[99], line_120[97], line_119[95], line_118[93], line_117[91], line_116[89], line_115[87], line_114[85], line_113[83], line_112[81], line_111[79], line_110[77], line_109[75], line_108[73], line_107[71], line_106[69], line_105[67], line_104[65], line_103[63], line_102[61], line_101[59], line_100[57], line_99[55], line_98[53], line_97[51], line_96[49], line_95[47], line_94[45], line_93[43], line_92[41], line_91[39], line_90[37], line_89[35], line_88[33], line_87[31], line_86[29], line_85[27], line_84[25], line_83[23], line_82[21], line_81[19], line_80[17], line_79[15], line_78[13], line_77[11], line_76[9], line_75[7], line_74[5], line_73[3], line_72[1], 71'b0};
assign col_114 = {line_128[114], line_127[112], line_126[110], line_125[108], line_124[106], line_123[104], line_122[102], line_121[100], line_120[98], line_119[96], line_118[94], line_117[92], line_116[90], line_115[88], line_114[86], line_113[84], line_112[82], line_111[80], line_110[78], line_109[76], line_108[74], line_107[72], line_106[70], line_105[68], line_104[66], line_103[64], line_102[62], line_101[60], line_100[58], line_99[56], line_98[54], line_97[52], line_96[50], line_95[48], line_94[46], line_93[44], line_92[42], line_91[40], line_90[38], line_89[36], line_88[34], line_87[32], line_86[30], line_85[28], line_84[26], line_83[24], line_82[22], line_81[20], line_80[18], line_79[16], line_78[14], line_77[12], line_76[10], line_75[8], line_74[6], line_73[4], line_72[2], line_71[0], 70'b0};
assign col_115 = {line_128[115], line_127[113], line_126[111], line_125[109], line_124[107], line_123[105], line_122[103], line_121[101], line_120[99], line_119[97], line_118[95], line_117[93], line_116[91], line_115[89], line_114[87], line_113[85], line_112[83], line_111[81], line_110[79], line_109[77], line_108[75], line_107[73], line_106[71], line_105[69], line_104[67], line_103[65], line_102[63], line_101[61], line_100[59], line_99[57], line_98[55], line_97[53], line_96[51], line_95[49], line_94[47], line_93[45], line_92[43], line_91[41], line_90[39], line_89[37], line_88[35], line_87[33], line_86[31], line_85[29], line_84[27], line_83[25], line_82[23], line_81[21], line_80[19], line_79[17], line_78[15], line_77[13], line_76[11], line_75[9], line_74[7], line_73[5], line_72[3], line_71[1], 70'b0};
assign col_116 = {line_128[116], line_127[114], line_126[112], line_125[110], line_124[108], line_123[106], line_122[104], line_121[102], line_120[100], line_119[98], line_118[96], line_117[94], line_116[92], line_115[90], line_114[88], line_113[86], line_112[84], line_111[82], line_110[80], line_109[78], line_108[76], line_107[74], line_106[72], line_105[70], line_104[68], line_103[66], line_102[64], line_101[62], line_100[60], line_99[58], line_98[56], line_97[54], line_96[52], line_95[50], line_94[48], line_93[46], line_92[44], line_91[42], line_90[40], line_89[38], line_88[36], line_87[34], line_86[32], line_85[30], line_84[28], line_83[26], line_82[24], line_81[22], line_80[20], line_79[18], line_78[16], line_77[14], line_76[12], line_75[10], line_74[8], line_73[6], line_72[4], line_71[2], line_70[0], 69'b0};
assign col_117 = {line_128[117], line_127[115], line_126[113], line_125[111], line_124[109], line_123[107], line_122[105], line_121[103], line_120[101], line_119[99], line_118[97], line_117[95], line_116[93], line_115[91], line_114[89], line_113[87], line_112[85], line_111[83], line_110[81], line_109[79], line_108[77], line_107[75], line_106[73], line_105[71], line_104[69], line_103[67], line_102[65], line_101[63], line_100[61], line_99[59], line_98[57], line_97[55], line_96[53], line_95[51], line_94[49], line_93[47], line_92[45], line_91[43], line_90[41], line_89[39], line_88[37], line_87[35], line_86[33], line_85[31], line_84[29], line_83[27], line_82[25], line_81[23], line_80[21], line_79[19], line_78[17], line_77[15], line_76[13], line_75[11], line_74[9], line_73[7], line_72[5], line_71[3], line_70[1], 69'b0};
assign col_118 = {line_128[118], line_127[116], line_126[114], line_125[112], line_124[110], line_123[108], line_122[106], line_121[104], line_120[102], line_119[100], line_118[98], line_117[96], line_116[94], line_115[92], line_114[90], line_113[88], line_112[86], line_111[84], line_110[82], line_109[80], line_108[78], line_107[76], line_106[74], line_105[72], line_104[70], line_103[68], line_102[66], line_101[64], line_100[62], line_99[60], line_98[58], line_97[56], line_96[54], line_95[52], line_94[50], line_93[48], line_92[46], line_91[44], line_90[42], line_89[40], line_88[38], line_87[36], line_86[34], line_85[32], line_84[30], line_83[28], line_82[26], line_81[24], line_80[22], line_79[20], line_78[18], line_77[16], line_76[14], line_75[12], line_74[10], line_73[8], line_72[6], line_71[4], line_70[2], line_69[0], 68'b0};
assign col_119 = {line_128[119], line_127[117], line_126[115], line_125[113], line_124[111], line_123[109], line_122[107], line_121[105], line_120[103], line_119[101], line_118[99], line_117[97], line_116[95], line_115[93], line_114[91], line_113[89], line_112[87], line_111[85], line_110[83], line_109[81], line_108[79], line_107[77], line_106[75], line_105[73], line_104[71], line_103[69], line_102[67], line_101[65], line_100[63], line_99[61], line_98[59], line_97[57], line_96[55], line_95[53], line_94[51], line_93[49], line_92[47], line_91[45], line_90[43], line_89[41], line_88[39], line_87[37], line_86[35], line_85[33], line_84[31], line_83[29], line_82[27], line_81[25], line_80[23], line_79[21], line_78[19], line_77[17], line_76[15], line_75[13], line_74[11], line_73[9], line_72[7], line_71[5], line_70[3], line_69[1], 68'b0};
assign col_120 = {line_128[120], line_127[118], line_126[116], line_125[114], line_124[112], line_123[110], line_122[108], line_121[106], line_120[104], line_119[102], line_118[100], line_117[98], line_116[96], line_115[94], line_114[92], line_113[90], line_112[88], line_111[86], line_110[84], line_109[82], line_108[80], line_107[78], line_106[76], line_105[74], line_104[72], line_103[70], line_102[68], line_101[66], line_100[64], line_99[62], line_98[60], line_97[58], line_96[56], line_95[54], line_94[52], line_93[50], line_92[48], line_91[46], line_90[44], line_89[42], line_88[40], line_87[38], line_86[36], line_85[34], line_84[32], line_83[30], line_82[28], line_81[26], line_80[24], line_79[22], line_78[20], line_77[18], line_76[16], line_75[14], line_74[12], line_73[10], line_72[8], line_71[6], line_70[4], line_69[2], line_68[0], 67'b0};
assign col_121 = {line_128[121], line_127[119], line_126[117], line_125[115], line_124[113], line_123[111], line_122[109], line_121[107], line_120[105], line_119[103], line_118[101], line_117[99], line_116[97], line_115[95], line_114[93], line_113[91], line_112[89], line_111[87], line_110[85], line_109[83], line_108[81], line_107[79], line_106[77], line_105[75], line_104[73], line_103[71], line_102[69], line_101[67], line_100[65], line_99[63], line_98[61], line_97[59], line_96[57], line_95[55], line_94[53], line_93[51], line_92[49], line_91[47], line_90[45], line_89[43], line_88[41], line_87[39], line_86[37], line_85[35], line_84[33], line_83[31], line_82[29], line_81[27], line_80[25], line_79[23], line_78[21], line_77[19], line_76[17], line_75[15], line_74[13], line_73[11], line_72[9], line_71[7], line_70[5], line_69[3], line_68[1], 67'b0};
assign col_122 = {line_128[122], line_127[120], line_126[118], line_125[116], line_124[114], line_123[112], line_122[110], line_121[108], line_120[106], line_119[104], line_118[102], line_117[100], line_116[98], line_115[96], line_114[94], line_113[92], line_112[90], line_111[88], line_110[86], line_109[84], line_108[82], line_107[80], line_106[78], line_105[76], line_104[74], line_103[72], line_102[70], line_101[68], line_100[66], line_99[64], line_98[62], line_97[60], line_96[58], line_95[56], line_94[54], line_93[52], line_92[50], line_91[48], line_90[46], line_89[44], line_88[42], line_87[40], line_86[38], line_85[36], line_84[34], line_83[32], line_82[30], line_81[28], line_80[26], line_79[24], line_78[22], line_77[20], line_76[18], line_75[16], line_74[14], line_73[12], line_72[10], line_71[8], line_70[6], line_69[4], line_68[2], line_67[0], 66'b0};
assign col_123 = {line_128[123], line_127[121], line_126[119], line_125[117], line_124[115], line_123[113], line_122[111], line_121[109], line_120[107], line_119[105], line_118[103], line_117[101], line_116[99], line_115[97], line_114[95], line_113[93], line_112[91], line_111[89], line_110[87], line_109[85], line_108[83], line_107[81], line_106[79], line_105[77], line_104[75], line_103[73], line_102[71], line_101[69], line_100[67], line_99[65], line_98[63], line_97[61], line_96[59], line_95[57], line_94[55], line_93[53], line_92[51], line_91[49], line_90[47], line_89[45], line_88[43], line_87[41], line_86[39], line_85[37], line_84[35], line_83[33], line_82[31], line_81[29], line_80[27], line_79[25], line_78[23], line_77[21], line_76[19], line_75[17], line_74[15], line_73[13], line_72[11], line_71[9], line_70[7], line_69[5], line_68[3], line_67[1], 66'b0};
assign col_124 = {line_128[124], line_127[122], line_126[120], line_125[118], line_124[116], line_123[114], line_122[112], line_121[110], line_120[108], line_119[106], line_118[104], line_117[102], line_116[100], line_115[98], line_114[96], line_113[94], line_112[92], line_111[90], line_110[88], line_109[86], line_108[84], line_107[82], line_106[80], line_105[78], line_104[76], line_103[74], line_102[72], line_101[70], line_100[68], line_99[66], line_98[64], line_97[62], line_96[60], line_95[58], line_94[56], line_93[54], line_92[52], line_91[50], line_90[48], line_89[46], line_88[44], line_87[42], line_86[40], line_85[38], line_84[36], line_83[34], line_82[32], line_81[30], line_80[28], line_79[26], line_78[24], line_77[22], line_76[20], line_75[18], line_74[16], line_73[14], line_72[12], line_71[10], line_70[8], line_69[6], line_68[4], line_67[2], line_66[0], 65'b0};
assign col_125 = {line_128[125], line_127[123], line_126[121], line_125[119], line_124[117], line_123[115], line_122[113], line_121[111], line_120[109], line_119[107], line_118[105], line_117[103], line_116[101], line_115[99], line_114[97], line_113[95], line_112[93], line_111[91], line_110[89], line_109[87], line_108[85], line_107[83], line_106[81], line_105[79], line_104[77], line_103[75], line_102[73], line_101[71], line_100[69], line_99[67], line_98[65], line_97[63], line_96[61], line_95[59], line_94[57], line_93[55], line_92[53], line_91[51], line_90[49], line_89[47], line_88[45], line_87[43], line_86[41], line_85[39], line_84[37], line_83[35], line_82[33], line_81[31], line_80[29], line_79[27], line_78[25], line_77[23], line_76[21], line_75[19], line_74[17], line_73[15], line_72[13], line_71[11], line_70[9], line_69[7], line_68[5], line_67[3], line_66[1], 65'b0};
assign col_126 = {line_128[126], line_127[124], line_126[122], line_125[120], line_124[118], line_123[116], line_122[114], line_121[112], line_120[110], line_119[108], line_118[106], line_117[104], line_116[102], line_115[100], line_114[98], line_113[96], line_112[94], line_111[92], line_110[90], line_109[88], line_108[86], line_107[84], line_106[82], line_105[80], line_104[78], line_103[76], line_102[74], line_101[72], line_100[70], line_99[68], line_98[66], line_97[64], line_96[62], line_95[60], line_94[58], line_93[56], line_92[54], line_91[52], line_90[50], line_89[48], line_88[46], line_87[44], line_86[42], line_85[40], line_84[38], line_83[36], line_82[34], line_81[32], line_80[30], line_79[28], line_78[26], line_77[24], line_76[22], line_75[20], line_74[18], line_73[16], line_72[14], line_71[12], line_70[10], line_69[8], line_68[6], line_67[4], line_66[2], line_65[0], 64'b0};
assign col_127 = {line_128[127], line_127[125], line_126[123], line_125[121], line_124[119], line_123[117], line_122[115], line_121[113], line_120[111], line_119[109], line_118[107], line_117[105], line_116[103], line_115[101], line_114[99], line_113[97], line_112[95], line_111[93], line_110[91], line_109[89], line_108[87], line_107[85], line_106[83], line_105[81], line_104[79], line_103[77], line_102[75], line_101[73], line_100[71], line_99[69], line_98[67], line_97[65], line_96[63], line_95[61], line_94[59], line_93[57], line_92[55], line_91[53], line_90[51], line_89[49], line_88[47], line_87[45], line_86[43], line_85[41], line_84[39], line_83[37], line_82[35], line_81[33], line_80[31], line_79[29], line_78[27], line_77[25], line_76[23], line_75[21], line_74[19], line_73[17], line_72[15], line_71[13], line_70[11], line_69[9], line_68[7], line_67[5], line_66[3], line_65[1], 64'b0};
assign col_128 = {line_128[128], line_127[126], line_126[124], line_125[122], line_124[120], line_123[118], line_122[116], line_121[114], line_120[112], line_119[110], line_118[108], line_117[106], line_116[104], line_115[102], line_114[100], line_113[98], line_112[96], line_111[94], line_110[92], line_109[90], line_108[88], line_107[86], line_106[84], line_105[82], line_104[80], line_103[78], line_102[76], line_101[74], line_100[72], line_99[70], line_98[68], line_97[66], line_96[64], line_95[62], line_94[60], line_93[58], line_92[56], line_91[54], line_90[52], line_89[50], line_88[48], line_87[46], line_86[44], line_85[42], line_84[40], line_83[38], line_82[36], line_81[34], line_80[32], line_79[30], line_78[28], line_77[26], line_76[24], line_75[22], line_74[20], line_73[18], line_72[16], line_71[14], line_70[12], line_69[10], line_68[8], line_67[6], line_66[4], line_65[2], line_64[0], 63'b0};
assign col_129 = {line_128[129], line_127[127], line_126[125], line_125[123], line_124[121], line_123[119], line_122[117], line_121[115], line_120[113], line_119[111], line_118[109], line_117[107], line_116[105], line_115[103], line_114[101], line_113[99], line_112[97], line_111[95], line_110[93], line_109[91], line_108[89], line_107[87], line_106[85], line_105[83], line_104[81], line_103[79], line_102[77], line_101[75], line_100[73], line_99[71], line_98[69], line_97[67], line_96[65], line_95[63], line_94[61], line_93[59], line_92[57], line_91[55], line_90[53], line_89[51], line_88[49], line_87[47], line_86[45], line_85[43], line_84[41], line_83[39], line_82[37], line_81[35], line_80[33], line_79[31], line_78[29], line_77[27], line_76[25], line_75[23], line_74[21], line_73[19], line_72[17], line_71[15], line_70[13], line_69[11], line_68[9], line_67[7], line_66[5], line_65[3], line_64[1], 63'b0};
assign col_130 = {line_128[130], line_127[128], line_126[126], line_125[124], line_124[122], line_123[120], line_122[118], line_121[116], line_120[114], line_119[112], line_118[110], line_117[108], line_116[106], line_115[104], line_114[102], line_113[100], line_112[98], line_111[96], line_110[94], line_109[92], line_108[90], line_107[88], line_106[86], line_105[84], line_104[82], line_103[80], line_102[78], line_101[76], line_100[74], line_99[72], line_98[70], line_97[68], line_96[66], line_95[64], line_94[62], line_93[60], line_92[58], line_91[56], line_90[54], line_89[52], line_88[50], line_87[48], line_86[46], line_85[44], line_84[42], line_83[40], line_82[38], line_81[36], line_80[34], line_79[32], line_78[30], line_77[28], line_76[26], line_75[24], line_74[22], line_73[20], line_72[18], line_71[16], line_70[14], line_69[12], line_68[10], line_67[8], line_66[6], line_65[4], line_64[2], line_63[0], 62'b0};
assign col_131 = {line_128[131], line_127[129], line_126[127], line_125[125], line_124[123], line_123[121], line_122[119], line_121[117], line_120[115], line_119[113], line_118[111], line_117[109], line_116[107], line_115[105], line_114[103], line_113[101], line_112[99], line_111[97], line_110[95], line_109[93], line_108[91], line_107[89], line_106[87], line_105[85], line_104[83], line_103[81], line_102[79], line_101[77], line_100[75], line_99[73], line_98[71], line_97[69], line_96[67], line_95[65], line_94[63], line_93[61], line_92[59], line_91[57], line_90[55], line_89[53], line_88[51], line_87[49], line_86[47], line_85[45], line_84[43], line_83[41], line_82[39], line_81[37], line_80[35], line_79[33], line_78[31], line_77[29], line_76[27], line_75[25], line_74[23], line_73[21], line_72[19], line_71[17], line_70[15], line_69[13], line_68[11], line_67[9], line_66[7], line_65[5], line_64[3], line_63[1], 62'b0};
assign col_132 = {line_128[132], line_127[130], line_126[128], line_125[126], line_124[124], line_123[122], line_122[120], line_121[118], line_120[116], line_119[114], line_118[112], line_117[110], line_116[108], line_115[106], line_114[104], line_113[102], line_112[100], line_111[98], line_110[96], line_109[94], line_108[92], line_107[90], line_106[88], line_105[86], line_104[84], line_103[82], line_102[80], line_101[78], line_100[76], line_99[74], line_98[72], line_97[70], line_96[68], line_95[66], line_94[64], line_93[62], line_92[60], line_91[58], line_90[56], line_89[54], line_88[52], line_87[50], line_86[48], line_85[46], line_84[44], line_83[42], line_82[40], line_81[38], line_80[36], line_79[34], line_78[32], line_77[30], line_76[28], line_75[26], line_74[24], line_73[22], line_72[20], line_71[18], line_70[16], line_69[14], line_68[12], line_67[10], line_66[8], line_65[6], line_64[4], line_63[2], line_62[0], 61'b0};
assign col_133 = {line_128[133], line_127[131], line_126[129], line_125[127], line_124[125], line_123[123], line_122[121], line_121[119], line_120[117], line_119[115], line_118[113], line_117[111], line_116[109], line_115[107], line_114[105], line_113[103], line_112[101], line_111[99], line_110[97], line_109[95], line_108[93], line_107[91], line_106[89], line_105[87], line_104[85], line_103[83], line_102[81], line_101[79], line_100[77], line_99[75], line_98[73], line_97[71], line_96[69], line_95[67], line_94[65], line_93[63], line_92[61], line_91[59], line_90[57], line_89[55], line_88[53], line_87[51], line_86[49], line_85[47], line_84[45], line_83[43], line_82[41], line_81[39], line_80[37], line_79[35], line_78[33], line_77[31], line_76[29], line_75[27], line_74[25], line_73[23], line_72[21], line_71[19], line_70[17], line_69[15], line_68[13], line_67[11], line_66[9], line_65[7], line_64[5], line_63[3], line_62[1], 61'b0};
assign col_134 = {line_128[134], line_127[132], line_126[130], line_125[128], line_124[126], line_123[124], line_122[122], line_121[120], line_120[118], line_119[116], line_118[114], line_117[112], line_116[110], line_115[108], line_114[106], line_113[104], line_112[102], line_111[100], line_110[98], line_109[96], line_108[94], line_107[92], line_106[90], line_105[88], line_104[86], line_103[84], line_102[82], line_101[80], line_100[78], line_99[76], line_98[74], line_97[72], line_96[70], line_95[68], line_94[66], line_93[64], line_92[62], line_91[60], line_90[58], line_89[56], line_88[54], line_87[52], line_86[50], line_85[48], line_84[46], line_83[44], line_82[42], line_81[40], line_80[38], line_79[36], line_78[34], line_77[32], line_76[30], line_75[28], line_74[26], line_73[24], line_72[22], line_71[20], line_70[18], line_69[16], line_68[14], line_67[12], line_66[10], line_65[8], line_64[6], line_63[4], line_62[2], line_61[0], 60'b0};
assign col_135 = {line_128[135], line_127[133], line_126[131], line_125[129], line_124[127], line_123[125], line_122[123], line_121[121], line_120[119], line_119[117], line_118[115], line_117[113], line_116[111], line_115[109], line_114[107], line_113[105], line_112[103], line_111[101], line_110[99], line_109[97], line_108[95], line_107[93], line_106[91], line_105[89], line_104[87], line_103[85], line_102[83], line_101[81], line_100[79], line_99[77], line_98[75], line_97[73], line_96[71], line_95[69], line_94[67], line_93[65], line_92[63], line_91[61], line_90[59], line_89[57], line_88[55], line_87[53], line_86[51], line_85[49], line_84[47], line_83[45], line_82[43], line_81[41], line_80[39], line_79[37], line_78[35], line_77[33], line_76[31], line_75[29], line_74[27], line_73[25], line_72[23], line_71[21], line_70[19], line_69[17], line_68[15], line_67[13], line_66[11], line_65[9], line_64[7], line_63[5], line_62[3], line_61[1], 60'b0};
assign col_136 = {line_128[136], line_127[134], line_126[132], line_125[130], line_124[128], line_123[126], line_122[124], line_121[122], line_120[120], line_119[118], line_118[116], line_117[114], line_116[112], line_115[110], line_114[108], line_113[106], line_112[104], line_111[102], line_110[100], line_109[98], line_108[96], line_107[94], line_106[92], line_105[90], line_104[88], line_103[86], line_102[84], line_101[82], line_100[80], line_99[78], line_98[76], line_97[74], line_96[72], line_95[70], line_94[68], line_93[66], line_92[64], line_91[62], line_90[60], line_89[58], line_88[56], line_87[54], line_86[52], line_85[50], line_84[48], line_83[46], line_82[44], line_81[42], line_80[40], line_79[38], line_78[36], line_77[34], line_76[32], line_75[30], line_74[28], line_73[26], line_72[24], line_71[22], line_70[20], line_69[18], line_68[16], line_67[14], line_66[12], line_65[10], line_64[8], line_63[6], line_62[4], line_61[2], line_60[0], 59'b0};
assign col_137 = {line_128[137], line_127[135], line_126[133], line_125[131], line_124[129], line_123[127], line_122[125], line_121[123], line_120[121], line_119[119], line_118[117], line_117[115], line_116[113], line_115[111], line_114[109], line_113[107], line_112[105], line_111[103], line_110[101], line_109[99], line_108[97], line_107[95], line_106[93], line_105[91], line_104[89], line_103[87], line_102[85], line_101[83], line_100[81], line_99[79], line_98[77], line_97[75], line_96[73], line_95[71], line_94[69], line_93[67], line_92[65], line_91[63], line_90[61], line_89[59], line_88[57], line_87[55], line_86[53], line_85[51], line_84[49], line_83[47], line_82[45], line_81[43], line_80[41], line_79[39], line_78[37], line_77[35], line_76[33], line_75[31], line_74[29], line_73[27], line_72[25], line_71[23], line_70[21], line_69[19], line_68[17], line_67[15], line_66[13], line_65[11], line_64[9], line_63[7], line_62[5], line_61[3], line_60[1], 59'b0};
assign col_138 = {line_128[138], line_127[136], line_126[134], line_125[132], line_124[130], line_123[128], line_122[126], line_121[124], line_120[122], line_119[120], line_118[118], line_117[116], line_116[114], line_115[112], line_114[110], line_113[108], line_112[106], line_111[104], line_110[102], line_109[100], line_108[98], line_107[96], line_106[94], line_105[92], line_104[90], line_103[88], line_102[86], line_101[84], line_100[82], line_99[80], line_98[78], line_97[76], line_96[74], line_95[72], line_94[70], line_93[68], line_92[66], line_91[64], line_90[62], line_89[60], line_88[58], line_87[56], line_86[54], line_85[52], line_84[50], line_83[48], line_82[46], line_81[44], line_80[42], line_79[40], line_78[38], line_77[36], line_76[34], line_75[32], line_74[30], line_73[28], line_72[26], line_71[24], line_70[22], line_69[20], line_68[18], line_67[16], line_66[14], line_65[12], line_64[10], line_63[8], line_62[6], line_61[4], line_60[2], line_59[0], 58'b0};
assign col_139 = {line_128[139], line_127[137], line_126[135], line_125[133], line_124[131], line_123[129], line_122[127], line_121[125], line_120[123], line_119[121], line_118[119], line_117[117], line_116[115], line_115[113], line_114[111], line_113[109], line_112[107], line_111[105], line_110[103], line_109[101], line_108[99], line_107[97], line_106[95], line_105[93], line_104[91], line_103[89], line_102[87], line_101[85], line_100[83], line_99[81], line_98[79], line_97[77], line_96[75], line_95[73], line_94[71], line_93[69], line_92[67], line_91[65], line_90[63], line_89[61], line_88[59], line_87[57], line_86[55], line_85[53], line_84[51], line_83[49], line_82[47], line_81[45], line_80[43], line_79[41], line_78[39], line_77[37], line_76[35], line_75[33], line_74[31], line_73[29], line_72[27], line_71[25], line_70[23], line_69[21], line_68[19], line_67[17], line_66[15], line_65[13], line_64[11], line_63[9], line_62[7], line_61[5], line_60[3], line_59[1], 58'b0};
assign col_140 = {line_128[140], line_127[138], line_126[136], line_125[134], line_124[132], line_123[130], line_122[128], line_121[126], line_120[124], line_119[122], line_118[120], line_117[118], line_116[116], line_115[114], line_114[112], line_113[110], line_112[108], line_111[106], line_110[104], line_109[102], line_108[100], line_107[98], line_106[96], line_105[94], line_104[92], line_103[90], line_102[88], line_101[86], line_100[84], line_99[82], line_98[80], line_97[78], line_96[76], line_95[74], line_94[72], line_93[70], line_92[68], line_91[66], line_90[64], line_89[62], line_88[60], line_87[58], line_86[56], line_85[54], line_84[52], line_83[50], line_82[48], line_81[46], line_80[44], line_79[42], line_78[40], line_77[38], line_76[36], line_75[34], line_74[32], line_73[30], line_72[28], line_71[26], line_70[24], line_69[22], line_68[20], line_67[18], line_66[16], line_65[14], line_64[12], line_63[10], line_62[8], line_61[6], line_60[4], line_59[2], line_58[0], 57'b0};
assign col_141 = {line_128[141], line_127[139], line_126[137], line_125[135], line_124[133], line_123[131], line_122[129], line_121[127], line_120[125], line_119[123], line_118[121], line_117[119], line_116[117], line_115[115], line_114[113], line_113[111], line_112[109], line_111[107], line_110[105], line_109[103], line_108[101], line_107[99], line_106[97], line_105[95], line_104[93], line_103[91], line_102[89], line_101[87], line_100[85], line_99[83], line_98[81], line_97[79], line_96[77], line_95[75], line_94[73], line_93[71], line_92[69], line_91[67], line_90[65], line_89[63], line_88[61], line_87[59], line_86[57], line_85[55], line_84[53], line_83[51], line_82[49], line_81[47], line_80[45], line_79[43], line_78[41], line_77[39], line_76[37], line_75[35], line_74[33], line_73[31], line_72[29], line_71[27], line_70[25], line_69[23], line_68[21], line_67[19], line_66[17], line_65[15], line_64[13], line_63[11], line_62[9], line_61[7], line_60[5], line_59[3], line_58[1], 57'b0};
assign col_142 = {line_128[142], line_127[140], line_126[138], line_125[136], line_124[134], line_123[132], line_122[130], line_121[128], line_120[126], line_119[124], line_118[122], line_117[120], line_116[118], line_115[116], line_114[114], line_113[112], line_112[110], line_111[108], line_110[106], line_109[104], line_108[102], line_107[100], line_106[98], line_105[96], line_104[94], line_103[92], line_102[90], line_101[88], line_100[86], line_99[84], line_98[82], line_97[80], line_96[78], line_95[76], line_94[74], line_93[72], line_92[70], line_91[68], line_90[66], line_89[64], line_88[62], line_87[60], line_86[58], line_85[56], line_84[54], line_83[52], line_82[50], line_81[48], line_80[46], line_79[44], line_78[42], line_77[40], line_76[38], line_75[36], line_74[34], line_73[32], line_72[30], line_71[28], line_70[26], line_69[24], line_68[22], line_67[20], line_66[18], line_65[16], line_64[14], line_63[12], line_62[10], line_61[8], line_60[6], line_59[4], line_58[2], line_57[0], 56'b0};
assign col_143 = {line_128[143], line_127[141], line_126[139], line_125[137], line_124[135], line_123[133], line_122[131], line_121[129], line_120[127], line_119[125], line_118[123], line_117[121], line_116[119], line_115[117], line_114[115], line_113[113], line_112[111], line_111[109], line_110[107], line_109[105], line_108[103], line_107[101], line_106[99], line_105[97], line_104[95], line_103[93], line_102[91], line_101[89], line_100[87], line_99[85], line_98[83], line_97[81], line_96[79], line_95[77], line_94[75], line_93[73], line_92[71], line_91[69], line_90[67], line_89[65], line_88[63], line_87[61], line_86[59], line_85[57], line_84[55], line_83[53], line_82[51], line_81[49], line_80[47], line_79[45], line_78[43], line_77[41], line_76[39], line_75[37], line_74[35], line_73[33], line_72[31], line_71[29], line_70[27], line_69[25], line_68[23], line_67[21], line_66[19], line_65[17], line_64[15], line_63[13], line_62[11], line_61[9], line_60[7], line_59[5], line_58[3], line_57[1], 56'b0};
assign col_144 = {line_128[144], line_127[142], line_126[140], line_125[138], line_124[136], line_123[134], line_122[132], line_121[130], line_120[128], line_119[126], line_118[124], line_117[122], line_116[120], line_115[118], line_114[116], line_113[114], line_112[112], line_111[110], line_110[108], line_109[106], line_108[104], line_107[102], line_106[100], line_105[98], line_104[96], line_103[94], line_102[92], line_101[90], line_100[88], line_99[86], line_98[84], line_97[82], line_96[80], line_95[78], line_94[76], line_93[74], line_92[72], line_91[70], line_90[68], line_89[66], line_88[64], line_87[62], line_86[60], line_85[58], line_84[56], line_83[54], line_82[52], line_81[50], line_80[48], line_79[46], line_78[44], line_77[42], line_76[40], line_75[38], line_74[36], line_73[34], line_72[32], line_71[30], line_70[28], line_69[26], line_68[24], line_67[22], line_66[20], line_65[18], line_64[16], line_63[14], line_62[12], line_61[10], line_60[8], line_59[6], line_58[4], line_57[2], line_56[0], 55'b0};
assign col_145 = {line_128[145], line_127[143], line_126[141], line_125[139], line_124[137], line_123[135], line_122[133], line_121[131], line_120[129], line_119[127], line_118[125], line_117[123], line_116[121], line_115[119], line_114[117], line_113[115], line_112[113], line_111[111], line_110[109], line_109[107], line_108[105], line_107[103], line_106[101], line_105[99], line_104[97], line_103[95], line_102[93], line_101[91], line_100[89], line_99[87], line_98[85], line_97[83], line_96[81], line_95[79], line_94[77], line_93[75], line_92[73], line_91[71], line_90[69], line_89[67], line_88[65], line_87[63], line_86[61], line_85[59], line_84[57], line_83[55], line_82[53], line_81[51], line_80[49], line_79[47], line_78[45], line_77[43], line_76[41], line_75[39], line_74[37], line_73[35], line_72[33], line_71[31], line_70[29], line_69[27], line_68[25], line_67[23], line_66[21], line_65[19], line_64[17], line_63[15], line_62[13], line_61[11], line_60[9], line_59[7], line_58[5], line_57[3], line_56[1], 55'b0};
assign col_146 = {line_128[146], line_127[144], line_126[142], line_125[140], line_124[138], line_123[136], line_122[134], line_121[132], line_120[130], line_119[128], line_118[126], line_117[124], line_116[122], line_115[120], line_114[118], line_113[116], line_112[114], line_111[112], line_110[110], line_109[108], line_108[106], line_107[104], line_106[102], line_105[100], line_104[98], line_103[96], line_102[94], line_101[92], line_100[90], line_99[88], line_98[86], line_97[84], line_96[82], line_95[80], line_94[78], line_93[76], line_92[74], line_91[72], line_90[70], line_89[68], line_88[66], line_87[64], line_86[62], line_85[60], line_84[58], line_83[56], line_82[54], line_81[52], line_80[50], line_79[48], line_78[46], line_77[44], line_76[42], line_75[40], line_74[38], line_73[36], line_72[34], line_71[32], line_70[30], line_69[28], line_68[26], line_67[24], line_66[22], line_65[20], line_64[18], line_63[16], line_62[14], line_61[12], line_60[10], line_59[8], line_58[6], line_57[4], line_56[2], line_55[0], 54'b0};
assign col_147 = {line_128[147], line_127[145], line_126[143], line_125[141], line_124[139], line_123[137], line_122[135], line_121[133], line_120[131], line_119[129], line_118[127], line_117[125], line_116[123], line_115[121], line_114[119], line_113[117], line_112[115], line_111[113], line_110[111], line_109[109], line_108[107], line_107[105], line_106[103], line_105[101], line_104[99], line_103[97], line_102[95], line_101[93], line_100[91], line_99[89], line_98[87], line_97[85], line_96[83], line_95[81], line_94[79], line_93[77], line_92[75], line_91[73], line_90[71], line_89[69], line_88[67], line_87[65], line_86[63], line_85[61], line_84[59], line_83[57], line_82[55], line_81[53], line_80[51], line_79[49], line_78[47], line_77[45], line_76[43], line_75[41], line_74[39], line_73[37], line_72[35], line_71[33], line_70[31], line_69[29], line_68[27], line_67[25], line_66[23], line_65[21], line_64[19], line_63[17], line_62[15], line_61[13], line_60[11], line_59[9], line_58[7], line_57[5], line_56[3], line_55[1], 54'b0};
assign col_148 = {line_128[148], line_127[146], line_126[144], line_125[142], line_124[140], line_123[138], line_122[136], line_121[134], line_120[132], line_119[130], line_118[128], line_117[126], line_116[124], line_115[122], line_114[120], line_113[118], line_112[116], line_111[114], line_110[112], line_109[110], line_108[108], line_107[106], line_106[104], line_105[102], line_104[100], line_103[98], line_102[96], line_101[94], line_100[92], line_99[90], line_98[88], line_97[86], line_96[84], line_95[82], line_94[80], line_93[78], line_92[76], line_91[74], line_90[72], line_89[70], line_88[68], line_87[66], line_86[64], line_85[62], line_84[60], line_83[58], line_82[56], line_81[54], line_80[52], line_79[50], line_78[48], line_77[46], line_76[44], line_75[42], line_74[40], line_73[38], line_72[36], line_71[34], line_70[32], line_69[30], line_68[28], line_67[26], line_66[24], line_65[22], line_64[20], line_63[18], line_62[16], line_61[14], line_60[12], line_59[10], line_58[8], line_57[6], line_56[4], line_55[2], line_54[0], 53'b0};
assign col_149 = {line_128[149], line_127[147], line_126[145], line_125[143], line_124[141], line_123[139], line_122[137], line_121[135], line_120[133], line_119[131], line_118[129], line_117[127], line_116[125], line_115[123], line_114[121], line_113[119], line_112[117], line_111[115], line_110[113], line_109[111], line_108[109], line_107[107], line_106[105], line_105[103], line_104[101], line_103[99], line_102[97], line_101[95], line_100[93], line_99[91], line_98[89], line_97[87], line_96[85], line_95[83], line_94[81], line_93[79], line_92[77], line_91[75], line_90[73], line_89[71], line_88[69], line_87[67], line_86[65], line_85[63], line_84[61], line_83[59], line_82[57], line_81[55], line_80[53], line_79[51], line_78[49], line_77[47], line_76[45], line_75[43], line_74[41], line_73[39], line_72[37], line_71[35], line_70[33], line_69[31], line_68[29], line_67[27], line_66[25], line_65[23], line_64[21], line_63[19], line_62[17], line_61[15], line_60[13], line_59[11], line_58[9], line_57[7], line_56[5], line_55[3], line_54[1], 53'b0};
assign col_150 = {line_128[150], line_127[148], line_126[146], line_125[144], line_124[142], line_123[140], line_122[138], line_121[136], line_120[134], line_119[132], line_118[130], line_117[128], line_116[126], line_115[124], line_114[122], line_113[120], line_112[118], line_111[116], line_110[114], line_109[112], line_108[110], line_107[108], line_106[106], line_105[104], line_104[102], line_103[100], line_102[98], line_101[96], line_100[94], line_99[92], line_98[90], line_97[88], line_96[86], line_95[84], line_94[82], line_93[80], line_92[78], line_91[76], line_90[74], line_89[72], line_88[70], line_87[68], line_86[66], line_85[64], line_84[62], line_83[60], line_82[58], line_81[56], line_80[54], line_79[52], line_78[50], line_77[48], line_76[46], line_75[44], line_74[42], line_73[40], line_72[38], line_71[36], line_70[34], line_69[32], line_68[30], line_67[28], line_66[26], line_65[24], line_64[22], line_63[20], line_62[18], line_61[16], line_60[14], line_59[12], line_58[10], line_57[8], line_56[6], line_55[4], line_54[2], line_53[0], 52'b0};
assign col_151 = {line_128[151], line_127[149], line_126[147], line_125[145], line_124[143], line_123[141], line_122[139], line_121[137], line_120[135], line_119[133], line_118[131], line_117[129], line_116[127], line_115[125], line_114[123], line_113[121], line_112[119], line_111[117], line_110[115], line_109[113], line_108[111], line_107[109], line_106[107], line_105[105], line_104[103], line_103[101], line_102[99], line_101[97], line_100[95], line_99[93], line_98[91], line_97[89], line_96[87], line_95[85], line_94[83], line_93[81], line_92[79], line_91[77], line_90[75], line_89[73], line_88[71], line_87[69], line_86[67], line_85[65], line_84[63], line_83[61], line_82[59], line_81[57], line_80[55], line_79[53], line_78[51], line_77[49], line_76[47], line_75[45], line_74[43], line_73[41], line_72[39], line_71[37], line_70[35], line_69[33], line_68[31], line_67[29], line_66[27], line_65[25], line_64[23], line_63[21], line_62[19], line_61[17], line_60[15], line_59[13], line_58[11], line_57[9], line_56[7], line_55[5], line_54[3], line_53[1], 52'b0};
assign col_152 = {line_128[152], line_127[150], line_126[148], line_125[146], line_124[144], line_123[142], line_122[140], line_121[138], line_120[136], line_119[134], line_118[132], line_117[130], line_116[128], line_115[126], line_114[124], line_113[122], line_112[120], line_111[118], line_110[116], line_109[114], line_108[112], line_107[110], line_106[108], line_105[106], line_104[104], line_103[102], line_102[100], line_101[98], line_100[96], line_99[94], line_98[92], line_97[90], line_96[88], line_95[86], line_94[84], line_93[82], line_92[80], line_91[78], line_90[76], line_89[74], line_88[72], line_87[70], line_86[68], line_85[66], line_84[64], line_83[62], line_82[60], line_81[58], line_80[56], line_79[54], line_78[52], line_77[50], line_76[48], line_75[46], line_74[44], line_73[42], line_72[40], line_71[38], line_70[36], line_69[34], line_68[32], line_67[30], line_66[28], line_65[26], line_64[24], line_63[22], line_62[20], line_61[18], line_60[16], line_59[14], line_58[12], line_57[10], line_56[8], line_55[6], line_54[4], line_53[2], line_52[0], 51'b0};
assign col_153 = {line_128[153], line_127[151], line_126[149], line_125[147], line_124[145], line_123[143], line_122[141], line_121[139], line_120[137], line_119[135], line_118[133], line_117[131], line_116[129], line_115[127], line_114[125], line_113[123], line_112[121], line_111[119], line_110[117], line_109[115], line_108[113], line_107[111], line_106[109], line_105[107], line_104[105], line_103[103], line_102[101], line_101[99], line_100[97], line_99[95], line_98[93], line_97[91], line_96[89], line_95[87], line_94[85], line_93[83], line_92[81], line_91[79], line_90[77], line_89[75], line_88[73], line_87[71], line_86[69], line_85[67], line_84[65], line_83[63], line_82[61], line_81[59], line_80[57], line_79[55], line_78[53], line_77[51], line_76[49], line_75[47], line_74[45], line_73[43], line_72[41], line_71[39], line_70[37], line_69[35], line_68[33], line_67[31], line_66[29], line_65[27], line_64[25], line_63[23], line_62[21], line_61[19], line_60[17], line_59[15], line_58[13], line_57[11], line_56[9], line_55[7], line_54[5], line_53[3], line_52[1], 51'b0};
assign col_154 = {line_128[154], line_127[152], line_126[150], line_125[148], line_124[146], line_123[144], line_122[142], line_121[140], line_120[138], line_119[136], line_118[134], line_117[132], line_116[130], line_115[128], line_114[126], line_113[124], line_112[122], line_111[120], line_110[118], line_109[116], line_108[114], line_107[112], line_106[110], line_105[108], line_104[106], line_103[104], line_102[102], line_101[100], line_100[98], line_99[96], line_98[94], line_97[92], line_96[90], line_95[88], line_94[86], line_93[84], line_92[82], line_91[80], line_90[78], line_89[76], line_88[74], line_87[72], line_86[70], line_85[68], line_84[66], line_83[64], line_82[62], line_81[60], line_80[58], line_79[56], line_78[54], line_77[52], line_76[50], line_75[48], line_74[46], line_73[44], line_72[42], line_71[40], line_70[38], line_69[36], line_68[34], line_67[32], line_66[30], line_65[28], line_64[26], line_63[24], line_62[22], line_61[20], line_60[18], line_59[16], line_58[14], line_57[12], line_56[10], line_55[8], line_54[6], line_53[4], line_52[2], line_51[0], 50'b0};
assign col_155 = {line_128[155], line_127[153], line_126[151], line_125[149], line_124[147], line_123[145], line_122[143], line_121[141], line_120[139], line_119[137], line_118[135], line_117[133], line_116[131], line_115[129], line_114[127], line_113[125], line_112[123], line_111[121], line_110[119], line_109[117], line_108[115], line_107[113], line_106[111], line_105[109], line_104[107], line_103[105], line_102[103], line_101[101], line_100[99], line_99[97], line_98[95], line_97[93], line_96[91], line_95[89], line_94[87], line_93[85], line_92[83], line_91[81], line_90[79], line_89[77], line_88[75], line_87[73], line_86[71], line_85[69], line_84[67], line_83[65], line_82[63], line_81[61], line_80[59], line_79[57], line_78[55], line_77[53], line_76[51], line_75[49], line_74[47], line_73[45], line_72[43], line_71[41], line_70[39], line_69[37], line_68[35], line_67[33], line_66[31], line_65[29], line_64[27], line_63[25], line_62[23], line_61[21], line_60[19], line_59[17], line_58[15], line_57[13], line_56[11], line_55[9], line_54[7], line_53[5], line_52[3], line_51[1], 50'b0};
assign col_156 = {line_128[156], line_127[154], line_126[152], line_125[150], line_124[148], line_123[146], line_122[144], line_121[142], line_120[140], line_119[138], line_118[136], line_117[134], line_116[132], line_115[130], line_114[128], line_113[126], line_112[124], line_111[122], line_110[120], line_109[118], line_108[116], line_107[114], line_106[112], line_105[110], line_104[108], line_103[106], line_102[104], line_101[102], line_100[100], line_99[98], line_98[96], line_97[94], line_96[92], line_95[90], line_94[88], line_93[86], line_92[84], line_91[82], line_90[80], line_89[78], line_88[76], line_87[74], line_86[72], line_85[70], line_84[68], line_83[66], line_82[64], line_81[62], line_80[60], line_79[58], line_78[56], line_77[54], line_76[52], line_75[50], line_74[48], line_73[46], line_72[44], line_71[42], line_70[40], line_69[38], line_68[36], line_67[34], line_66[32], line_65[30], line_64[28], line_63[26], line_62[24], line_61[22], line_60[20], line_59[18], line_58[16], line_57[14], line_56[12], line_55[10], line_54[8], line_53[6], line_52[4], line_51[2], line_50[0], 49'b0};
assign col_157 = {line_128[157], line_127[155], line_126[153], line_125[151], line_124[149], line_123[147], line_122[145], line_121[143], line_120[141], line_119[139], line_118[137], line_117[135], line_116[133], line_115[131], line_114[129], line_113[127], line_112[125], line_111[123], line_110[121], line_109[119], line_108[117], line_107[115], line_106[113], line_105[111], line_104[109], line_103[107], line_102[105], line_101[103], line_100[101], line_99[99], line_98[97], line_97[95], line_96[93], line_95[91], line_94[89], line_93[87], line_92[85], line_91[83], line_90[81], line_89[79], line_88[77], line_87[75], line_86[73], line_85[71], line_84[69], line_83[67], line_82[65], line_81[63], line_80[61], line_79[59], line_78[57], line_77[55], line_76[53], line_75[51], line_74[49], line_73[47], line_72[45], line_71[43], line_70[41], line_69[39], line_68[37], line_67[35], line_66[33], line_65[31], line_64[29], line_63[27], line_62[25], line_61[23], line_60[21], line_59[19], line_58[17], line_57[15], line_56[13], line_55[11], line_54[9], line_53[7], line_52[5], line_51[3], line_50[1], 49'b0};
assign col_158 = {line_128[158], line_127[156], line_126[154], line_125[152], line_124[150], line_123[148], line_122[146], line_121[144], line_120[142], line_119[140], line_118[138], line_117[136], line_116[134], line_115[132], line_114[130], line_113[128], line_112[126], line_111[124], line_110[122], line_109[120], line_108[118], line_107[116], line_106[114], line_105[112], line_104[110], line_103[108], line_102[106], line_101[104], line_100[102], line_99[100], line_98[98], line_97[96], line_96[94], line_95[92], line_94[90], line_93[88], line_92[86], line_91[84], line_90[82], line_89[80], line_88[78], line_87[76], line_86[74], line_85[72], line_84[70], line_83[68], line_82[66], line_81[64], line_80[62], line_79[60], line_78[58], line_77[56], line_76[54], line_75[52], line_74[50], line_73[48], line_72[46], line_71[44], line_70[42], line_69[40], line_68[38], line_67[36], line_66[34], line_65[32], line_64[30], line_63[28], line_62[26], line_61[24], line_60[22], line_59[20], line_58[18], line_57[16], line_56[14], line_55[12], line_54[10], line_53[8], line_52[6], line_51[4], line_50[2], line_49[0], 48'b0};
assign col_159 = {line_128[159], line_127[157], line_126[155], line_125[153], line_124[151], line_123[149], line_122[147], line_121[145], line_120[143], line_119[141], line_118[139], line_117[137], line_116[135], line_115[133], line_114[131], line_113[129], line_112[127], line_111[125], line_110[123], line_109[121], line_108[119], line_107[117], line_106[115], line_105[113], line_104[111], line_103[109], line_102[107], line_101[105], line_100[103], line_99[101], line_98[99], line_97[97], line_96[95], line_95[93], line_94[91], line_93[89], line_92[87], line_91[85], line_90[83], line_89[81], line_88[79], line_87[77], line_86[75], line_85[73], line_84[71], line_83[69], line_82[67], line_81[65], line_80[63], line_79[61], line_78[59], line_77[57], line_76[55], line_75[53], line_74[51], line_73[49], line_72[47], line_71[45], line_70[43], line_69[41], line_68[39], line_67[37], line_66[35], line_65[33], line_64[31], line_63[29], line_62[27], line_61[25], line_60[23], line_59[21], line_58[19], line_57[17], line_56[15], line_55[13], line_54[11], line_53[9], line_52[7], line_51[5], line_50[3], line_49[1], 48'b0};
assign col_160 = {line_128[160], line_127[158], line_126[156], line_125[154], line_124[152], line_123[150], line_122[148], line_121[146], line_120[144], line_119[142], line_118[140], line_117[138], line_116[136], line_115[134], line_114[132], line_113[130], line_112[128], line_111[126], line_110[124], line_109[122], line_108[120], line_107[118], line_106[116], line_105[114], line_104[112], line_103[110], line_102[108], line_101[106], line_100[104], line_99[102], line_98[100], line_97[98], line_96[96], line_95[94], line_94[92], line_93[90], line_92[88], line_91[86], line_90[84], line_89[82], line_88[80], line_87[78], line_86[76], line_85[74], line_84[72], line_83[70], line_82[68], line_81[66], line_80[64], line_79[62], line_78[60], line_77[58], line_76[56], line_75[54], line_74[52], line_73[50], line_72[48], line_71[46], line_70[44], line_69[42], line_68[40], line_67[38], line_66[36], line_65[34], line_64[32], line_63[30], line_62[28], line_61[26], line_60[24], line_59[22], line_58[20], line_57[18], line_56[16], line_55[14], line_54[12], line_53[10], line_52[8], line_51[6], line_50[4], line_49[2], line_48[0], 47'b0};
assign col_161 = {line_128[161], line_127[159], line_126[157], line_125[155], line_124[153], line_123[151], line_122[149], line_121[147], line_120[145], line_119[143], line_118[141], line_117[139], line_116[137], line_115[135], line_114[133], line_113[131], line_112[129], line_111[127], line_110[125], line_109[123], line_108[121], line_107[119], line_106[117], line_105[115], line_104[113], line_103[111], line_102[109], line_101[107], line_100[105], line_99[103], line_98[101], line_97[99], line_96[97], line_95[95], line_94[93], line_93[91], line_92[89], line_91[87], line_90[85], line_89[83], line_88[81], line_87[79], line_86[77], line_85[75], line_84[73], line_83[71], line_82[69], line_81[67], line_80[65], line_79[63], line_78[61], line_77[59], line_76[57], line_75[55], line_74[53], line_73[51], line_72[49], line_71[47], line_70[45], line_69[43], line_68[41], line_67[39], line_66[37], line_65[35], line_64[33], line_63[31], line_62[29], line_61[27], line_60[25], line_59[23], line_58[21], line_57[19], line_56[17], line_55[15], line_54[13], line_53[11], line_52[9], line_51[7], line_50[5], line_49[3], line_48[1], 47'b0};
assign col_162 = {line_128[162], line_127[160], line_126[158], line_125[156], line_124[154], line_123[152], line_122[150], line_121[148], line_120[146], line_119[144], line_118[142], line_117[140], line_116[138], line_115[136], line_114[134], line_113[132], line_112[130], line_111[128], line_110[126], line_109[124], line_108[122], line_107[120], line_106[118], line_105[116], line_104[114], line_103[112], line_102[110], line_101[108], line_100[106], line_99[104], line_98[102], line_97[100], line_96[98], line_95[96], line_94[94], line_93[92], line_92[90], line_91[88], line_90[86], line_89[84], line_88[82], line_87[80], line_86[78], line_85[76], line_84[74], line_83[72], line_82[70], line_81[68], line_80[66], line_79[64], line_78[62], line_77[60], line_76[58], line_75[56], line_74[54], line_73[52], line_72[50], line_71[48], line_70[46], line_69[44], line_68[42], line_67[40], line_66[38], line_65[36], line_64[34], line_63[32], line_62[30], line_61[28], line_60[26], line_59[24], line_58[22], line_57[20], line_56[18], line_55[16], line_54[14], line_53[12], line_52[10], line_51[8], line_50[6], line_49[4], line_48[2], line_47[0], 46'b0};
assign col_163 = {line_128[163], line_127[161], line_126[159], line_125[157], line_124[155], line_123[153], line_122[151], line_121[149], line_120[147], line_119[145], line_118[143], line_117[141], line_116[139], line_115[137], line_114[135], line_113[133], line_112[131], line_111[129], line_110[127], line_109[125], line_108[123], line_107[121], line_106[119], line_105[117], line_104[115], line_103[113], line_102[111], line_101[109], line_100[107], line_99[105], line_98[103], line_97[101], line_96[99], line_95[97], line_94[95], line_93[93], line_92[91], line_91[89], line_90[87], line_89[85], line_88[83], line_87[81], line_86[79], line_85[77], line_84[75], line_83[73], line_82[71], line_81[69], line_80[67], line_79[65], line_78[63], line_77[61], line_76[59], line_75[57], line_74[55], line_73[53], line_72[51], line_71[49], line_70[47], line_69[45], line_68[43], line_67[41], line_66[39], line_65[37], line_64[35], line_63[33], line_62[31], line_61[29], line_60[27], line_59[25], line_58[23], line_57[21], line_56[19], line_55[17], line_54[15], line_53[13], line_52[11], line_51[9], line_50[7], line_49[5], line_48[3], line_47[1], 46'b0};
assign col_164 = {line_128[164], line_127[162], line_126[160], line_125[158], line_124[156], line_123[154], line_122[152], line_121[150], line_120[148], line_119[146], line_118[144], line_117[142], line_116[140], line_115[138], line_114[136], line_113[134], line_112[132], line_111[130], line_110[128], line_109[126], line_108[124], line_107[122], line_106[120], line_105[118], line_104[116], line_103[114], line_102[112], line_101[110], line_100[108], line_99[106], line_98[104], line_97[102], line_96[100], line_95[98], line_94[96], line_93[94], line_92[92], line_91[90], line_90[88], line_89[86], line_88[84], line_87[82], line_86[80], line_85[78], line_84[76], line_83[74], line_82[72], line_81[70], line_80[68], line_79[66], line_78[64], line_77[62], line_76[60], line_75[58], line_74[56], line_73[54], line_72[52], line_71[50], line_70[48], line_69[46], line_68[44], line_67[42], line_66[40], line_65[38], line_64[36], line_63[34], line_62[32], line_61[30], line_60[28], line_59[26], line_58[24], line_57[22], line_56[20], line_55[18], line_54[16], line_53[14], line_52[12], line_51[10], line_50[8], line_49[6], line_48[4], line_47[2], line_46[0], 45'b0};
assign col_165 = {line_128[165], line_127[163], line_126[161], line_125[159], line_124[157], line_123[155], line_122[153], line_121[151], line_120[149], line_119[147], line_118[145], line_117[143], line_116[141], line_115[139], line_114[137], line_113[135], line_112[133], line_111[131], line_110[129], line_109[127], line_108[125], line_107[123], line_106[121], line_105[119], line_104[117], line_103[115], line_102[113], line_101[111], line_100[109], line_99[107], line_98[105], line_97[103], line_96[101], line_95[99], line_94[97], line_93[95], line_92[93], line_91[91], line_90[89], line_89[87], line_88[85], line_87[83], line_86[81], line_85[79], line_84[77], line_83[75], line_82[73], line_81[71], line_80[69], line_79[67], line_78[65], line_77[63], line_76[61], line_75[59], line_74[57], line_73[55], line_72[53], line_71[51], line_70[49], line_69[47], line_68[45], line_67[43], line_66[41], line_65[39], line_64[37], line_63[35], line_62[33], line_61[31], line_60[29], line_59[27], line_58[25], line_57[23], line_56[21], line_55[19], line_54[17], line_53[15], line_52[13], line_51[11], line_50[9], line_49[7], line_48[5], line_47[3], line_46[1], 45'b0};
assign col_166 = {line_128[166], line_127[164], line_126[162], line_125[160], line_124[158], line_123[156], line_122[154], line_121[152], line_120[150], line_119[148], line_118[146], line_117[144], line_116[142], line_115[140], line_114[138], line_113[136], line_112[134], line_111[132], line_110[130], line_109[128], line_108[126], line_107[124], line_106[122], line_105[120], line_104[118], line_103[116], line_102[114], line_101[112], line_100[110], line_99[108], line_98[106], line_97[104], line_96[102], line_95[100], line_94[98], line_93[96], line_92[94], line_91[92], line_90[90], line_89[88], line_88[86], line_87[84], line_86[82], line_85[80], line_84[78], line_83[76], line_82[74], line_81[72], line_80[70], line_79[68], line_78[66], line_77[64], line_76[62], line_75[60], line_74[58], line_73[56], line_72[54], line_71[52], line_70[50], line_69[48], line_68[46], line_67[44], line_66[42], line_65[40], line_64[38], line_63[36], line_62[34], line_61[32], line_60[30], line_59[28], line_58[26], line_57[24], line_56[22], line_55[20], line_54[18], line_53[16], line_52[14], line_51[12], line_50[10], line_49[8], line_48[6], line_47[4], line_46[2], line_45[0], 44'b0};
assign col_167 = {line_128[167], line_127[165], line_126[163], line_125[161], line_124[159], line_123[157], line_122[155], line_121[153], line_120[151], line_119[149], line_118[147], line_117[145], line_116[143], line_115[141], line_114[139], line_113[137], line_112[135], line_111[133], line_110[131], line_109[129], line_108[127], line_107[125], line_106[123], line_105[121], line_104[119], line_103[117], line_102[115], line_101[113], line_100[111], line_99[109], line_98[107], line_97[105], line_96[103], line_95[101], line_94[99], line_93[97], line_92[95], line_91[93], line_90[91], line_89[89], line_88[87], line_87[85], line_86[83], line_85[81], line_84[79], line_83[77], line_82[75], line_81[73], line_80[71], line_79[69], line_78[67], line_77[65], line_76[63], line_75[61], line_74[59], line_73[57], line_72[55], line_71[53], line_70[51], line_69[49], line_68[47], line_67[45], line_66[43], line_65[41], line_64[39], line_63[37], line_62[35], line_61[33], line_60[31], line_59[29], line_58[27], line_57[25], line_56[23], line_55[21], line_54[19], line_53[17], line_52[15], line_51[13], line_50[11], line_49[9], line_48[7], line_47[5], line_46[3], line_45[1], 44'b0};
assign col_168 = {line_128[168], line_127[166], line_126[164], line_125[162], line_124[160], line_123[158], line_122[156], line_121[154], line_120[152], line_119[150], line_118[148], line_117[146], line_116[144], line_115[142], line_114[140], line_113[138], line_112[136], line_111[134], line_110[132], line_109[130], line_108[128], line_107[126], line_106[124], line_105[122], line_104[120], line_103[118], line_102[116], line_101[114], line_100[112], line_99[110], line_98[108], line_97[106], line_96[104], line_95[102], line_94[100], line_93[98], line_92[96], line_91[94], line_90[92], line_89[90], line_88[88], line_87[86], line_86[84], line_85[82], line_84[80], line_83[78], line_82[76], line_81[74], line_80[72], line_79[70], line_78[68], line_77[66], line_76[64], line_75[62], line_74[60], line_73[58], line_72[56], line_71[54], line_70[52], line_69[50], line_68[48], line_67[46], line_66[44], line_65[42], line_64[40], line_63[38], line_62[36], line_61[34], line_60[32], line_59[30], line_58[28], line_57[26], line_56[24], line_55[22], line_54[20], line_53[18], line_52[16], line_51[14], line_50[12], line_49[10], line_48[8], line_47[6], line_46[4], line_45[2], line_44[0], 43'b0};
assign col_169 = {line_128[169], line_127[167], line_126[165], line_125[163], line_124[161], line_123[159], line_122[157], line_121[155], line_120[153], line_119[151], line_118[149], line_117[147], line_116[145], line_115[143], line_114[141], line_113[139], line_112[137], line_111[135], line_110[133], line_109[131], line_108[129], line_107[127], line_106[125], line_105[123], line_104[121], line_103[119], line_102[117], line_101[115], line_100[113], line_99[111], line_98[109], line_97[107], line_96[105], line_95[103], line_94[101], line_93[99], line_92[97], line_91[95], line_90[93], line_89[91], line_88[89], line_87[87], line_86[85], line_85[83], line_84[81], line_83[79], line_82[77], line_81[75], line_80[73], line_79[71], line_78[69], line_77[67], line_76[65], line_75[63], line_74[61], line_73[59], line_72[57], line_71[55], line_70[53], line_69[51], line_68[49], line_67[47], line_66[45], line_65[43], line_64[41], line_63[39], line_62[37], line_61[35], line_60[33], line_59[31], line_58[29], line_57[27], line_56[25], line_55[23], line_54[21], line_53[19], line_52[17], line_51[15], line_50[13], line_49[11], line_48[9], line_47[7], line_46[5], line_45[3], line_44[1], 43'b0};
assign col_170 = {line_128[170], line_127[168], line_126[166], line_125[164], line_124[162], line_123[160], line_122[158], line_121[156], line_120[154], line_119[152], line_118[150], line_117[148], line_116[146], line_115[144], line_114[142], line_113[140], line_112[138], line_111[136], line_110[134], line_109[132], line_108[130], line_107[128], line_106[126], line_105[124], line_104[122], line_103[120], line_102[118], line_101[116], line_100[114], line_99[112], line_98[110], line_97[108], line_96[106], line_95[104], line_94[102], line_93[100], line_92[98], line_91[96], line_90[94], line_89[92], line_88[90], line_87[88], line_86[86], line_85[84], line_84[82], line_83[80], line_82[78], line_81[76], line_80[74], line_79[72], line_78[70], line_77[68], line_76[66], line_75[64], line_74[62], line_73[60], line_72[58], line_71[56], line_70[54], line_69[52], line_68[50], line_67[48], line_66[46], line_65[44], line_64[42], line_63[40], line_62[38], line_61[36], line_60[34], line_59[32], line_58[30], line_57[28], line_56[26], line_55[24], line_54[22], line_53[20], line_52[18], line_51[16], line_50[14], line_49[12], line_48[10], line_47[8], line_46[6], line_45[4], line_44[2], line_43[0], 42'b0};
assign col_171 = {line_128[171], line_127[169], line_126[167], line_125[165], line_124[163], line_123[161], line_122[159], line_121[157], line_120[155], line_119[153], line_118[151], line_117[149], line_116[147], line_115[145], line_114[143], line_113[141], line_112[139], line_111[137], line_110[135], line_109[133], line_108[131], line_107[129], line_106[127], line_105[125], line_104[123], line_103[121], line_102[119], line_101[117], line_100[115], line_99[113], line_98[111], line_97[109], line_96[107], line_95[105], line_94[103], line_93[101], line_92[99], line_91[97], line_90[95], line_89[93], line_88[91], line_87[89], line_86[87], line_85[85], line_84[83], line_83[81], line_82[79], line_81[77], line_80[75], line_79[73], line_78[71], line_77[69], line_76[67], line_75[65], line_74[63], line_73[61], line_72[59], line_71[57], line_70[55], line_69[53], line_68[51], line_67[49], line_66[47], line_65[45], line_64[43], line_63[41], line_62[39], line_61[37], line_60[35], line_59[33], line_58[31], line_57[29], line_56[27], line_55[25], line_54[23], line_53[21], line_52[19], line_51[17], line_50[15], line_49[13], line_48[11], line_47[9], line_46[7], line_45[5], line_44[3], line_43[1], 42'b0};
assign col_172 = {line_128[172], line_127[170], line_126[168], line_125[166], line_124[164], line_123[162], line_122[160], line_121[158], line_120[156], line_119[154], line_118[152], line_117[150], line_116[148], line_115[146], line_114[144], line_113[142], line_112[140], line_111[138], line_110[136], line_109[134], line_108[132], line_107[130], line_106[128], line_105[126], line_104[124], line_103[122], line_102[120], line_101[118], line_100[116], line_99[114], line_98[112], line_97[110], line_96[108], line_95[106], line_94[104], line_93[102], line_92[100], line_91[98], line_90[96], line_89[94], line_88[92], line_87[90], line_86[88], line_85[86], line_84[84], line_83[82], line_82[80], line_81[78], line_80[76], line_79[74], line_78[72], line_77[70], line_76[68], line_75[66], line_74[64], line_73[62], line_72[60], line_71[58], line_70[56], line_69[54], line_68[52], line_67[50], line_66[48], line_65[46], line_64[44], line_63[42], line_62[40], line_61[38], line_60[36], line_59[34], line_58[32], line_57[30], line_56[28], line_55[26], line_54[24], line_53[22], line_52[20], line_51[18], line_50[16], line_49[14], line_48[12], line_47[10], line_46[8], line_45[6], line_44[4], line_43[2], line_42[0], 41'b0};
assign col_173 = {line_128[173], line_127[171], line_126[169], line_125[167], line_124[165], line_123[163], line_122[161], line_121[159], line_120[157], line_119[155], line_118[153], line_117[151], line_116[149], line_115[147], line_114[145], line_113[143], line_112[141], line_111[139], line_110[137], line_109[135], line_108[133], line_107[131], line_106[129], line_105[127], line_104[125], line_103[123], line_102[121], line_101[119], line_100[117], line_99[115], line_98[113], line_97[111], line_96[109], line_95[107], line_94[105], line_93[103], line_92[101], line_91[99], line_90[97], line_89[95], line_88[93], line_87[91], line_86[89], line_85[87], line_84[85], line_83[83], line_82[81], line_81[79], line_80[77], line_79[75], line_78[73], line_77[71], line_76[69], line_75[67], line_74[65], line_73[63], line_72[61], line_71[59], line_70[57], line_69[55], line_68[53], line_67[51], line_66[49], line_65[47], line_64[45], line_63[43], line_62[41], line_61[39], line_60[37], line_59[35], line_58[33], line_57[31], line_56[29], line_55[27], line_54[25], line_53[23], line_52[21], line_51[19], line_50[17], line_49[15], line_48[13], line_47[11], line_46[9], line_45[7], line_44[5], line_43[3], line_42[1], 41'b0};
assign col_174 = {line_128[174], line_127[172], line_126[170], line_125[168], line_124[166], line_123[164], line_122[162], line_121[160], line_120[158], line_119[156], line_118[154], line_117[152], line_116[150], line_115[148], line_114[146], line_113[144], line_112[142], line_111[140], line_110[138], line_109[136], line_108[134], line_107[132], line_106[130], line_105[128], line_104[126], line_103[124], line_102[122], line_101[120], line_100[118], line_99[116], line_98[114], line_97[112], line_96[110], line_95[108], line_94[106], line_93[104], line_92[102], line_91[100], line_90[98], line_89[96], line_88[94], line_87[92], line_86[90], line_85[88], line_84[86], line_83[84], line_82[82], line_81[80], line_80[78], line_79[76], line_78[74], line_77[72], line_76[70], line_75[68], line_74[66], line_73[64], line_72[62], line_71[60], line_70[58], line_69[56], line_68[54], line_67[52], line_66[50], line_65[48], line_64[46], line_63[44], line_62[42], line_61[40], line_60[38], line_59[36], line_58[34], line_57[32], line_56[30], line_55[28], line_54[26], line_53[24], line_52[22], line_51[20], line_50[18], line_49[16], line_48[14], line_47[12], line_46[10], line_45[8], line_44[6], line_43[4], line_42[2], line_41[0], 40'b0};
assign col_175 = {line_128[175], line_127[173], line_126[171], line_125[169], line_124[167], line_123[165], line_122[163], line_121[161], line_120[159], line_119[157], line_118[155], line_117[153], line_116[151], line_115[149], line_114[147], line_113[145], line_112[143], line_111[141], line_110[139], line_109[137], line_108[135], line_107[133], line_106[131], line_105[129], line_104[127], line_103[125], line_102[123], line_101[121], line_100[119], line_99[117], line_98[115], line_97[113], line_96[111], line_95[109], line_94[107], line_93[105], line_92[103], line_91[101], line_90[99], line_89[97], line_88[95], line_87[93], line_86[91], line_85[89], line_84[87], line_83[85], line_82[83], line_81[81], line_80[79], line_79[77], line_78[75], line_77[73], line_76[71], line_75[69], line_74[67], line_73[65], line_72[63], line_71[61], line_70[59], line_69[57], line_68[55], line_67[53], line_66[51], line_65[49], line_64[47], line_63[45], line_62[43], line_61[41], line_60[39], line_59[37], line_58[35], line_57[33], line_56[31], line_55[29], line_54[27], line_53[25], line_52[23], line_51[21], line_50[19], line_49[17], line_48[15], line_47[13], line_46[11], line_45[9], line_44[7], line_43[5], line_42[3], line_41[1], 40'b0};
assign col_176 = {line_128[176], line_127[174], line_126[172], line_125[170], line_124[168], line_123[166], line_122[164], line_121[162], line_120[160], line_119[158], line_118[156], line_117[154], line_116[152], line_115[150], line_114[148], line_113[146], line_112[144], line_111[142], line_110[140], line_109[138], line_108[136], line_107[134], line_106[132], line_105[130], line_104[128], line_103[126], line_102[124], line_101[122], line_100[120], line_99[118], line_98[116], line_97[114], line_96[112], line_95[110], line_94[108], line_93[106], line_92[104], line_91[102], line_90[100], line_89[98], line_88[96], line_87[94], line_86[92], line_85[90], line_84[88], line_83[86], line_82[84], line_81[82], line_80[80], line_79[78], line_78[76], line_77[74], line_76[72], line_75[70], line_74[68], line_73[66], line_72[64], line_71[62], line_70[60], line_69[58], line_68[56], line_67[54], line_66[52], line_65[50], line_64[48], line_63[46], line_62[44], line_61[42], line_60[40], line_59[38], line_58[36], line_57[34], line_56[32], line_55[30], line_54[28], line_53[26], line_52[24], line_51[22], line_50[20], line_49[18], line_48[16], line_47[14], line_46[12], line_45[10], line_44[8], line_43[6], line_42[4], line_41[2], line_40[0], 39'b0};
assign col_177 = {line_128[177], line_127[175], line_126[173], line_125[171], line_124[169], line_123[167], line_122[165], line_121[163], line_120[161], line_119[159], line_118[157], line_117[155], line_116[153], line_115[151], line_114[149], line_113[147], line_112[145], line_111[143], line_110[141], line_109[139], line_108[137], line_107[135], line_106[133], line_105[131], line_104[129], line_103[127], line_102[125], line_101[123], line_100[121], line_99[119], line_98[117], line_97[115], line_96[113], line_95[111], line_94[109], line_93[107], line_92[105], line_91[103], line_90[101], line_89[99], line_88[97], line_87[95], line_86[93], line_85[91], line_84[89], line_83[87], line_82[85], line_81[83], line_80[81], line_79[79], line_78[77], line_77[75], line_76[73], line_75[71], line_74[69], line_73[67], line_72[65], line_71[63], line_70[61], line_69[59], line_68[57], line_67[55], line_66[53], line_65[51], line_64[49], line_63[47], line_62[45], line_61[43], line_60[41], line_59[39], line_58[37], line_57[35], line_56[33], line_55[31], line_54[29], line_53[27], line_52[25], line_51[23], line_50[21], line_49[19], line_48[17], line_47[15], line_46[13], line_45[11], line_44[9], line_43[7], line_42[5], line_41[3], line_40[1], 39'b0};
assign col_178 = {line_128[178], line_127[176], line_126[174], line_125[172], line_124[170], line_123[168], line_122[166], line_121[164], line_120[162], line_119[160], line_118[158], line_117[156], line_116[154], line_115[152], line_114[150], line_113[148], line_112[146], line_111[144], line_110[142], line_109[140], line_108[138], line_107[136], line_106[134], line_105[132], line_104[130], line_103[128], line_102[126], line_101[124], line_100[122], line_99[120], line_98[118], line_97[116], line_96[114], line_95[112], line_94[110], line_93[108], line_92[106], line_91[104], line_90[102], line_89[100], line_88[98], line_87[96], line_86[94], line_85[92], line_84[90], line_83[88], line_82[86], line_81[84], line_80[82], line_79[80], line_78[78], line_77[76], line_76[74], line_75[72], line_74[70], line_73[68], line_72[66], line_71[64], line_70[62], line_69[60], line_68[58], line_67[56], line_66[54], line_65[52], line_64[50], line_63[48], line_62[46], line_61[44], line_60[42], line_59[40], line_58[38], line_57[36], line_56[34], line_55[32], line_54[30], line_53[28], line_52[26], line_51[24], line_50[22], line_49[20], line_48[18], line_47[16], line_46[14], line_45[12], line_44[10], line_43[8], line_42[6], line_41[4], line_40[2], line_39[0], 38'b0};
assign col_179 = {line_128[179], line_127[177], line_126[175], line_125[173], line_124[171], line_123[169], line_122[167], line_121[165], line_120[163], line_119[161], line_118[159], line_117[157], line_116[155], line_115[153], line_114[151], line_113[149], line_112[147], line_111[145], line_110[143], line_109[141], line_108[139], line_107[137], line_106[135], line_105[133], line_104[131], line_103[129], line_102[127], line_101[125], line_100[123], line_99[121], line_98[119], line_97[117], line_96[115], line_95[113], line_94[111], line_93[109], line_92[107], line_91[105], line_90[103], line_89[101], line_88[99], line_87[97], line_86[95], line_85[93], line_84[91], line_83[89], line_82[87], line_81[85], line_80[83], line_79[81], line_78[79], line_77[77], line_76[75], line_75[73], line_74[71], line_73[69], line_72[67], line_71[65], line_70[63], line_69[61], line_68[59], line_67[57], line_66[55], line_65[53], line_64[51], line_63[49], line_62[47], line_61[45], line_60[43], line_59[41], line_58[39], line_57[37], line_56[35], line_55[33], line_54[31], line_53[29], line_52[27], line_51[25], line_50[23], line_49[21], line_48[19], line_47[17], line_46[15], line_45[13], line_44[11], line_43[9], line_42[7], line_41[5], line_40[3], line_39[1], 38'b0};
assign col_180 = {line_128[180], line_127[178], line_126[176], line_125[174], line_124[172], line_123[170], line_122[168], line_121[166], line_120[164], line_119[162], line_118[160], line_117[158], line_116[156], line_115[154], line_114[152], line_113[150], line_112[148], line_111[146], line_110[144], line_109[142], line_108[140], line_107[138], line_106[136], line_105[134], line_104[132], line_103[130], line_102[128], line_101[126], line_100[124], line_99[122], line_98[120], line_97[118], line_96[116], line_95[114], line_94[112], line_93[110], line_92[108], line_91[106], line_90[104], line_89[102], line_88[100], line_87[98], line_86[96], line_85[94], line_84[92], line_83[90], line_82[88], line_81[86], line_80[84], line_79[82], line_78[80], line_77[78], line_76[76], line_75[74], line_74[72], line_73[70], line_72[68], line_71[66], line_70[64], line_69[62], line_68[60], line_67[58], line_66[56], line_65[54], line_64[52], line_63[50], line_62[48], line_61[46], line_60[44], line_59[42], line_58[40], line_57[38], line_56[36], line_55[34], line_54[32], line_53[30], line_52[28], line_51[26], line_50[24], line_49[22], line_48[20], line_47[18], line_46[16], line_45[14], line_44[12], line_43[10], line_42[8], line_41[6], line_40[4], line_39[2], line_38[0], 37'b0};
assign col_181 = {line_128[181], line_127[179], line_126[177], line_125[175], line_124[173], line_123[171], line_122[169], line_121[167], line_120[165], line_119[163], line_118[161], line_117[159], line_116[157], line_115[155], line_114[153], line_113[151], line_112[149], line_111[147], line_110[145], line_109[143], line_108[141], line_107[139], line_106[137], line_105[135], line_104[133], line_103[131], line_102[129], line_101[127], line_100[125], line_99[123], line_98[121], line_97[119], line_96[117], line_95[115], line_94[113], line_93[111], line_92[109], line_91[107], line_90[105], line_89[103], line_88[101], line_87[99], line_86[97], line_85[95], line_84[93], line_83[91], line_82[89], line_81[87], line_80[85], line_79[83], line_78[81], line_77[79], line_76[77], line_75[75], line_74[73], line_73[71], line_72[69], line_71[67], line_70[65], line_69[63], line_68[61], line_67[59], line_66[57], line_65[55], line_64[53], line_63[51], line_62[49], line_61[47], line_60[45], line_59[43], line_58[41], line_57[39], line_56[37], line_55[35], line_54[33], line_53[31], line_52[29], line_51[27], line_50[25], line_49[23], line_48[21], line_47[19], line_46[17], line_45[15], line_44[13], line_43[11], line_42[9], line_41[7], line_40[5], line_39[3], line_38[1], 37'b0};
assign col_182 = {line_128[182], line_127[180], line_126[178], line_125[176], line_124[174], line_123[172], line_122[170], line_121[168], line_120[166], line_119[164], line_118[162], line_117[160], line_116[158], line_115[156], line_114[154], line_113[152], line_112[150], line_111[148], line_110[146], line_109[144], line_108[142], line_107[140], line_106[138], line_105[136], line_104[134], line_103[132], line_102[130], line_101[128], line_100[126], line_99[124], line_98[122], line_97[120], line_96[118], line_95[116], line_94[114], line_93[112], line_92[110], line_91[108], line_90[106], line_89[104], line_88[102], line_87[100], line_86[98], line_85[96], line_84[94], line_83[92], line_82[90], line_81[88], line_80[86], line_79[84], line_78[82], line_77[80], line_76[78], line_75[76], line_74[74], line_73[72], line_72[70], line_71[68], line_70[66], line_69[64], line_68[62], line_67[60], line_66[58], line_65[56], line_64[54], line_63[52], line_62[50], line_61[48], line_60[46], line_59[44], line_58[42], line_57[40], line_56[38], line_55[36], line_54[34], line_53[32], line_52[30], line_51[28], line_50[26], line_49[24], line_48[22], line_47[20], line_46[18], line_45[16], line_44[14], line_43[12], line_42[10], line_41[8], line_40[6], line_39[4], line_38[2], line_37[0], 36'b0};
assign col_183 = {line_128[183], line_127[181], line_126[179], line_125[177], line_124[175], line_123[173], line_122[171], line_121[169], line_120[167], line_119[165], line_118[163], line_117[161], line_116[159], line_115[157], line_114[155], line_113[153], line_112[151], line_111[149], line_110[147], line_109[145], line_108[143], line_107[141], line_106[139], line_105[137], line_104[135], line_103[133], line_102[131], line_101[129], line_100[127], line_99[125], line_98[123], line_97[121], line_96[119], line_95[117], line_94[115], line_93[113], line_92[111], line_91[109], line_90[107], line_89[105], line_88[103], line_87[101], line_86[99], line_85[97], line_84[95], line_83[93], line_82[91], line_81[89], line_80[87], line_79[85], line_78[83], line_77[81], line_76[79], line_75[77], line_74[75], line_73[73], line_72[71], line_71[69], line_70[67], line_69[65], line_68[63], line_67[61], line_66[59], line_65[57], line_64[55], line_63[53], line_62[51], line_61[49], line_60[47], line_59[45], line_58[43], line_57[41], line_56[39], line_55[37], line_54[35], line_53[33], line_52[31], line_51[29], line_50[27], line_49[25], line_48[23], line_47[21], line_46[19], line_45[17], line_44[15], line_43[13], line_42[11], line_41[9], line_40[7], line_39[5], line_38[3], line_37[1], 36'b0};
assign col_184 = {line_128[184], line_127[182], line_126[180], line_125[178], line_124[176], line_123[174], line_122[172], line_121[170], line_120[168], line_119[166], line_118[164], line_117[162], line_116[160], line_115[158], line_114[156], line_113[154], line_112[152], line_111[150], line_110[148], line_109[146], line_108[144], line_107[142], line_106[140], line_105[138], line_104[136], line_103[134], line_102[132], line_101[130], line_100[128], line_99[126], line_98[124], line_97[122], line_96[120], line_95[118], line_94[116], line_93[114], line_92[112], line_91[110], line_90[108], line_89[106], line_88[104], line_87[102], line_86[100], line_85[98], line_84[96], line_83[94], line_82[92], line_81[90], line_80[88], line_79[86], line_78[84], line_77[82], line_76[80], line_75[78], line_74[76], line_73[74], line_72[72], line_71[70], line_70[68], line_69[66], line_68[64], line_67[62], line_66[60], line_65[58], line_64[56], line_63[54], line_62[52], line_61[50], line_60[48], line_59[46], line_58[44], line_57[42], line_56[40], line_55[38], line_54[36], line_53[34], line_52[32], line_51[30], line_50[28], line_49[26], line_48[24], line_47[22], line_46[20], line_45[18], line_44[16], line_43[14], line_42[12], line_41[10], line_40[8], line_39[6], line_38[4], line_37[2], line_36[0], 35'b0};
assign col_185 = {line_128[185], line_127[183], line_126[181], line_125[179], line_124[177], line_123[175], line_122[173], line_121[171], line_120[169], line_119[167], line_118[165], line_117[163], line_116[161], line_115[159], line_114[157], line_113[155], line_112[153], line_111[151], line_110[149], line_109[147], line_108[145], line_107[143], line_106[141], line_105[139], line_104[137], line_103[135], line_102[133], line_101[131], line_100[129], line_99[127], line_98[125], line_97[123], line_96[121], line_95[119], line_94[117], line_93[115], line_92[113], line_91[111], line_90[109], line_89[107], line_88[105], line_87[103], line_86[101], line_85[99], line_84[97], line_83[95], line_82[93], line_81[91], line_80[89], line_79[87], line_78[85], line_77[83], line_76[81], line_75[79], line_74[77], line_73[75], line_72[73], line_71[71], line_70[69], line_69[67], line_68[65], line_67[63], line_66[61], line_65[59], line_64[57], line_63[55], line_62[53], line_61[51], line_60[49], line_59[47], line_58[45], line_57[43], line_56[41], line_55[39], line_54[37], line_53[35], line_52[33], line_51[31], line_50[29], line_49[27], line_48[25], line_47[23], line_46[21], line_45[19], line_44[17], line_43[15], line_42[13], line_41[11], line_40[9], line_39[7], line_38[5], line_37[3], line_36[1], 35'b0};
assign col_186 = {line_128[186], line_127[184], line_126[182], line_125[180], line_124[178], line_123[176], line_122[174], line_121[172], line_120[170], line_119[168], line_118[166], line_117[164], line_116[162], line_115[160], line_114[158], line_113[156], line_112[154], line_111[152], line_110[150], line_109[148], line_108[146], line_107[144], line_106[142], line_105[140], line_104[138], line_103[136], line_102[134], line_101[132], line_100[130], line_99[128], line_98[126], line_97[124], line_96[122], line_95[120], line_94[118], line_93[116], line_92[114], line_91[112], line_90[110], line_89[108], line_88[106], line_87[104], line_86[102], line_85[100], line_84[98], line_83[96], line_82[94], line_81[92], line_80[90], line_79[88], line_78[86], line_77[84], line_76[82], line_75[80], line_74[78], line_73[76], line_72[74], line_71[72], line_70[70], line_69[68], line_68[66], line_67[64], line_66[62], line_65[60], line_64[58], line_63[56], line_62[54], line_61[52], line_60[50], line_59[48], line_58[46], line_57[44], line_56[42], line_55[40], line_54[38], line_53[36], line_52[34], line_51[32], line_50[30], line_49[28], line_48[26], line_47[24], line_46[22], line_45[20], line_44[18], line_43[16], line_42[14], line_41[12], line_40[10], line_39[8], line_38[6], line_37[4], line_36[2], line_35[0], 34'b0};
assign col_187 = {line_128[187], line_127[185], line_126[183], line_125[181], line_124[179], line_123[177], line_122[175], line_121[173], line_120[171], line_119[169], line_118[167], line_117[165], line_116[163], line_115[161], line_114[159], line_113[157], line_112[155], line_111[153], line_110[151], line_109[149], line_108[147], line_107[145], line_106[143], line_105[141], line_104[139], line_103[137], line_102[135], line_101[133], line_100[131], line_99[129], line_98[127], line_97[125], line_96[123], line_95[121], line_94[119], line_93[117], line_92[115], line_91[113], line_90[111], line_89[109], line_88[107], line_87[105], line_86[103], line_85[101], line_84[99], line_83[97], line_82[95], line_81[93], line_80[91], line_79[89], line_78[87], line_77[85], line_76[83], line_75[81], line_74[79], line_73[77], line_72[75], line_71[73], line_70[71], line_69[69], line_68[67], line_67[65], line_66[63], line_65[61], line_64[59], line_63[57], line_62[55], line_61[53], line_60[51], line_59[49], line_58[47], line_57[45], line_56[43], line_55[41], line_54[39], line_53[37], line_52[35], line_51[33], line_50[31], line_49[29], line_48[27], line_47[25], line_46[23], line_45[21], line_44[19], line_43[17], line_42[15], line_41[13], line_40[11], line_39[9], line_38[7], line_37[5], line_36[3], line_35[1], 34'b0};
assign col_188 = {line_128[188], line_127[186], line_126[184], line_125[182], line_124[180], line_123[178], line_122[176], line_121[174], line_120[172], line_119[170], line_118[168], line_117[166], line_116[164], line_115[162], line_114[160], line_113[158], line_112[156], line_111[154], line_110[152], line_109[150], line_108[148], line_107[146], line_106[144], line_105[142], line_104[140], line_103[138], line_102[136], line_101[134], line_100[132], line_99[130], line_98[128], line_97[126], line_96[124], line_95[122], line_94[120], line_93[118], line_92[116], line_91[114], line_90[112], line_89[110], line_88[108], line_87[106], line_86[104], line_85[102], line_84[100], line_83[98], line_82[96], line_81[94], line_80[92], line_79[90], line_78[88], line_77[86], line_76[84], line_75[82], line_74[80], line_73[78], line_72[76], line_71[74], line_70[72], line_69[70], line_68[68], line_67[66], line_66[64], line_65[62], line_64[60], line_63[58], line_62[56], line_61[54], line_60[52], line_59[50], line_58[48], line_57[46], line_56[44], line_55[42], line_54[40], line_53[38], line_52[36], line_51[34], line_50[32], line_49[30], line_48[28], line_47[26], line_46[24], line_45[22], line_44[20], line_43[18], line_42[16], line_41[14], line_40[12], line_39[10], line_38[8], line_37[6], line_36[4], line_35[2], line_34[0], 33'b0};
assign col_189 = {line_128[189], line_127[187], line_126[185], line_125[183], line_124[181], line_123[179], line_122[177], line_121[175], line_120[173], line_119[171], line_118[169], line_117[167], line_116[165], line_115[163], line_114[161], line_113[159], line_112[157], line_111[155], line_110[153], line_109[151], line_108[149], line_107[147], line_106[145], line_105[143], line_104[141], line_103[139], line_102[137], line_101[135], line_100[133], line_99[131], line_98[129], line_97[127], line_96[125], line_95[123], line_94[121], line_93[119], line_92[117], line_91[115], line_90[113], line_89[111], line_88[109], line_87[107], line_86[105], line_85[103], line_84[101], line_83[99], line_82[97], line_81[95], line_80[93], line_79[91], line_78[89], line_77[87], line_76[85], line_75[83], line_74[81], line_73[79], line_72[77], line_71[75], line_70[73], line_69[71], line_68[69], line_67[67], line_66[65], line_65[63], line_64[61], line_63[59], line_62[57], line_61[55], line_60[53], line_59[51], line_58[49], line_57[47], line_56[45], line_55[43], line_54[41], line_53[39], line_52[37], line_51[35], line_50[33], line_49[31], line_48[29], line_47[27], line_46[25], line_45[23], line_44[21], line_43[19], line_42[17], line_41[15], line_40[13], line_39[11], line_38[9], line_37[7], line_36[5], line_35[3], line_34[1], 33'b0};
assign col_190 = {line_128[190], line_127[188], line_126[186], line_125[184], line_124[182], line_123[180], line_122[178], line_121[176], line_120[174], line_119[172], line_118[170], line_117[168], line_116[166], line_115[164], line_114[162], line_113[160], line_112[158], line_111[156], line_110[154], line_109[152], line_108[150], line_107[148], line_106[146], line_105[144], line_104[142], line_103[140], line_102[138], line_101[136], line_100[134], line_99[132], line_98[130], line_97[128], line_96[126], line_95[124], line_94[122], line_93[120], line_92[118], line_91[116], line_90[114], line_89[112], line_88[110], line_87[108], line_86[106], line_85[104], line_84[102], line_83[100], line_82[98], line_81[96], line_80[94], line_79[92], line_78[90], line_77[88], line_76[86], line_75[84], line_74[82], line_73[80], line_72[78], line_71[76], line_70[74], line_69[72], line_68[70], line_67[68], line_66[66], line_65[64], line_64[62], line_63[60], line_62[58], line_61[56], line_60[54], line_59[52], line_58[50], line_57[48], line_56[46], line_55[44], line_54[42], line_53[40], line_52[38], line_51[36], line_50[34], line_49[32], line_48[30], line_47[28], line_46[26], line_45[24], line_44[22], line_43[20], line_42[18], line_41[16], line_40[14], line_39[12], line_38[10], line_37[8], line_36[6], line_35[4], line_34[2], line_33[0], 32'b0};
assign col_191 = {line_128[191], line_127[189], line_126[187], line_125[185], line_124[183], line_123[181], line_122[179], line_121[177], line_120[175], line_119[173], line_118[171], line_117[169], line_116[167], line_115[165], line_114[163], line_113[161], line_112[159], line_111[157], line_110[155], line_109[153], line_108[151], line_107[149], line_106[147], line_105[145], line_104[143], line_103[141], line_102[139], line_101[137], line_100[135], line_99[133], line_98[131], line_97[129], line_96[127], line_95[125], line_94[123], line_93[121], line_92[119], line_91[117], line_90[115], line_89[113], line_88[111], line_87[109], line_86[107], line_85[105], line_84[103], line_83[101], line_82[99], line_81[97], line_80[95], line_79[93], line_78[91], line_77[89], line_76[87], line_75[85], line_74[83], line_73[81], line_72[79], line_71[77], line_70[75], line_69[73], line_68[71], line_67[69], line_66[67], line_65[65], line_64[63], line_63[61], line_62[59], line_61[57], line_60[55], line_59[53], line_58[51], line_57[49], line_56[47], line_55[45], line_54[43], line_53[41], line_52[39], line_51[37], line_50[35], line_49[33], line_48[31], line_47[29], line_46[27], line_45[25], line_44[23], line_43[21], line_42[19], line_41[17], line_40[15], line_39[13], line_38[11], line_37[9], line_36[7], line_35[5], line_34[3], line_33[1], 32'b0};
assign col_192 = {line_128[192], line_127[190], line_126[188], line_125[186], line_124[184], line_123[182], line_122[180], line_121[178], line_120[176], line_119[174], line_118[172], line_117[170], line_116[168], line_115[166], line_114[164], line_113[162], line_112[160], line_111[158], line_110[156], line_109[154], line_108[152], line_107[150], line_106[148], line_105[146], line_104[144], line_103[142], line_102[140], line_101[138], line_100[136], line_99[134], line_98[132], line_97[130], line_96[128], line_95[126], line_94[124], line_93[122], line_92[120], line_91[118], line_90[116], line_89[114], line_88[112], line_87[110], line_86[108], line_85[106], line_84[104], line_83[102], line_82[100], line_81[98], line_80[96], line_79[94], line_78[92], line_77[90], line_76[88], line_75[86], line_74[84], line_73[82], line_72[80], line_71[78], line_70[76], line_69[74], line_68[72], line_67[70], line_66[68], line_65[66], line_64[64], line_63[62], line_62[60], line_61[58], line_60[56], line_59[54], line_58[52], line_57[50], line_56[48], line_55[46], line_54[44], line_53[42], line_52[40], line_51[38], line_50[36], line_49[34], line_48[32], line_47[30], line_46[28], line_45[26], line_44[24], line_43[22], line_42[20], line_41[18], line_40[16], line_39[14], line_38[12], line_37[10], line_36[8], line_35[6], line_34[4], line_33[2], line_32[0], 31'b0};
assign col_193 = {line_128[193], line_127[191], line_126[189], line_125[187], line_124[185], line_123[183], line_122[181], line_121[179], line_120[177], line_119[175], line_118[173], line_117[171], line_116[169], line_115[167], line_114[165], line_113[163], line_112[161], line_111[159], line_110[157], line_109[155], line_108[153], line_107[151], line_106[149], line_105[147], line_104[145], line_103[143], line_102[141], line_101[139], line_100[137], line_99[135], line_98[133], line_97[131], line_96[129], line_95[127], line_94[125], line_93[123], line_92[121], line_91[119], line_90[117], line_89[115], line_88[113], line_87[111], line_86[109], line_85[107], line_84[105], line_83[103], line_82[101], line_81[99], line_80[97], line_79[95], line_78[93], line_77[91], line_76[89], line_75[87], line_74[85], line_73[83], line_72[81], line_71[79], line_70[77], line_69[75], line_68[73], line_67[71], line_66[69], line_65[67], line_64[65], line_63[63], line_62[61], line_61[59], line_60[57], line_59[55], line_58[53], line_57[51], line_56[49], line_55[47], line_54[45], line_53[43], line_52[41], line_51[39], line_50[37], line_49[35], line_48[33], line_47[31], line_46[29], line_45[27], line_44[25], line_43[23], line_42[21], line_41[19], line_40[17], line_39[15], line_38[13], line_37[11], line_36[9], line_35[7], line_34[5], line_33[3], line_32[1], 31'b0};
assign col_194 = {line_128[194], line_127[192], line_126[190], line_125[188], line_124[186], line_123[184], line_122[182], line_121[180], line_120[178], line_119[176], line_118[174], line_117[172], line_116[170], line_115[168], line_114[166], line_113[164], line_112[162], line_111[160], line_110[158], line_109[156], line_108[154], line_107[152], line_106[150], line_105[148], line_104[146], line_103[144], line_102[142], line_101[140], line_100[138], line_99[136], line_98[134], line_97[132], line_96[130], line_95[128], line_94[126], line_93[124], line_92[122], line_91[120], line_90[118], line_89[116], line_88[114], line_87[112], line_86[110], line_85[108], line_84[106], line_83[104], line_82[102], line_81[100], line_80[98], line_79[96], line_78[94], line_77[92], line_76[90], line_75[88], line_74[86], line_73[84], line_72[82], line_71[80], line_70[78], line_69[76], line_68[74], line_67[72], line_66[70], line_65[68], line_64[66], line_63[64], line_62[62], line_61[60], line_60[58], line_59[56], line_58[54], line_57[52], line_56[50], line_55[48], line_54[46], line_53[44], line_52[42], line_51[40], line_50[38], line_49[36], line_48[34], line_47[32], line_46[30], line_45[28], line_44[26], line_43[24], line_42[22], line_41[20], line_40[18], line_39[16], line_38[14], line_37[12], line_36[10], line_35[8], line_34[6], line_33[4], line_32[2], line_31[0], 30'b0};
assign col_195 = {line_128[195], line_127[193], line_126[191], line_125[189], line_124[187], line_123[185], line_122[183], line_121[181], line_120[179], line_119[177], line_118[175], line_117[173], line_116[171], line_115[169], line_114[167], line_113[165], line_112[163], line_111[161], line_110[159], line_109[157], line_108[155], line_107[153], line_106[151], line_105[149], line_104[147], line_103[145], line_102[143], line_101[141], line_100[139], line_99[137], line_98[135], line_97[133], line_96[131], line_95[129], line_94[127], line_93[125], line_92[123], line_91[121], line_90[119], line_89[117], line_88[115], line_87[113], line_86[111], line_85[109], line_84[107], line_83[105], line_82[103], line_81[101], line_80[99], line_79[97], line_78[95], line_77[93], line_76[91], line_75[89], line_74[87], line_73[85], line_72[83], line_71[81], line_70[79], line_69[77], line_68[75], line_67[73], line_66[71], line_65[69], line_64[67], line_63[65], line_62[63], line_61[61], line_60[59], line_59[57], line_58[55], line_57[53], line_56[51], line_55[49], line_54[47], line_53[45], line_52[43], line_51[41], line_50[39], line_49[37], line_48[35], line_47[33], line_46[31], line_45[29], line_44[27], line_43[25], line_42[23], line_41[21], line_40[19], line_39[17], line_38[15], line_37[13], line_36[11], line_35[9], line_34[7], line_33[5], line_32[3], line_31[1], 30'b0};
assign col_196 = {line_128[196], line_127[194], line_126[192], line_125[190], line_124[188], line_123[186], line_122[184], line_121[182], line_120[180], line_119[178], line_118[176], line_117[174], line_116[172], line_115[170], line_114[168], line_113[166], line_112[164], line_111[162], line_110[160], line_109[158], line_108[156], line_107[154], line_106[152], line_105[150], line_104[148], line_103[146], line_102[144], line_101[142], line_100[140], line_99[138], line_98[136], line_97[134], line_96[132], line_95[130], line_94[128], line_93[126], line_92[124], line_91[122], line_90[120], line_89[118], line_88[116], line_87[114], line_86[112], line_85[110], line_84[108], line_83[106], line_82[104], line_81[102], line_80[100], line_79[98], line_78[96], line_77[94], line_76[92], line_75[90], line_74[88], line_73[86], line_72[84], line_71[82], line_70[80], line_69[78], line_68[76], line_67[74], line_66[72], line_65[70], line_64[68], line_63[66], line_62[64], line_61[62], line_60[60], line_59[58], line_58[56], line_57[54], line_56[52], line_55[50], line_54[48], line_53[46], line_52[44], line_51[42], line_50[40], line_49[38], line_48[36], line_47[34], line_46[32], line_45[30], line_44[28], line_43[26], line_42[24], line_41[22], line_40[20], line_39[18], line_38[16], line_37[14], line_36[12], line_35[10], line_34[8], line_33[6], line_32[4], line_31[2], line_30[0], 29'b0};
assign col_197 = {line_128[197], line_127[195], line_126[193], line_125[191], line_124[189], line_123[187], line_122[185], line_121[183], line_120[181], line_119[179], line_118[177], line_117[175], line_116[173], line_115[171], line_114[169], line_113[167], line_112[165], line_111[163], line_110[161], line_109[159], line_108[157], line_107[155], line_106[153], line_105[151], line_104[149], line_103[147], line_102[145], line_101[143], line_100[141], line_99[139], line_98[137], line_97[135], line_96[133], line_95[131], line_94[129], line_93[127], line_92[125], line_91[123], line_90[121], line_89[119], line_88[117], line_87[115], line_86[113], line_85[111], line_84[109], line_83[107], line_82[105], line_81[103], line_80[101], line_79[99], line_78[97], line_77[95], line_76[93], line_75[91], line_74[89], line_73[87], line_72[85], line_71[83], line_70[81], line_69[79], line_68[77], line_67[75], line_66[73], line_65[71], line_64[69], line_63[67], line_62[65], line_61[63], line_60[61], line_59[59], line_58[57], line_57[55], line_56[53], line_55[51], line_54[49], line_53[47], line_52[45], line_51[43], line_50[41], line_49[39], line_48[37], line_47[35], line_46[33], line_45[31], line_44[29], line_43[27], line_42[25], line_41[23], line_40[21], line_39[19], line_38[17], line_37[15], line_36[13], line_35[11], line_34[9], line_33[7], line_32[5], line_31[3], line_30[1], 29'b0};
assign col_198 = {line_128[198], line_127[196], line_126[194], line_125[192], line_124[190], line_123[188], line_122[186], line_121[184], line_120[182], line_119[180], line_118[178], line_117[176], line_116[174], line_115[172], line_114[170], line_113[168], line_112[166], line_111[164], line_110[162], line_109[160], line_108[158], line_107[156], line_106[154], line_105[152], line_104[150], line_103[148], line_102[146], line_101[144], line_100[142], line_99[140], line_98[138], line_97[136], line_96[134], line_95[132], line_94[130], line_93[128], line_92[126], line_91[124], line_90[122], line_89[120], line_88[118], line_87[116], line_86[114], line_85[112], line_84[110], line_83[108], line_82[106], line_81[104], line_80[102], line_79[100], line_78[98], line_77[96], line_76[94], line_75[92], line_74[90], line_73[88], line_72[86], line_71[84], line_70[82], line_69[80], line_68[78], line_67[76], line_66[74], line_65[72], line_64[70], line_63[68], line_62[66], line_61[64], line_60[62], line_59[60], line_58[58], line_57[56], line_56[54], line_55[52], line_54[50], line_53[48], line_52[46], line_51[44], line_50[42], line_49[40], line_48[38], line_47[36], line_46[34], line_45[32], line_44[30], line_43[28], line_42[26], line_41[24], line_40[22], line_39[20], line_38[18], line_37[16], line_36[14], line_35[12], line_34[10], line_33[8], line_32[6], line_31[4], line_30[2], line_29[0], 28'b0};
assign col_199 = {line_128[199], line_127[197], line_126[195], line_125[193], line_124[191], line_123[189], line_122[187], line_121[185], line_120[183], line_119[181], line_118[179], line_117[177], line_116[175], line_115[173], line_114[171], line_113[169], line_112[167], line_111[165], line_110[163], line_109[161], line_108[159], line_107[157], line_106[155], line_105[153], line_104[151], line_103[149], line_102[147], line_101[145], line_100[143], line_99[141], line_98[139], line_97[137], line_96[135], line_95[133], line_94[131], line_93[129], line_92[127], line_91[125], line_90[123], line_89[121], line_88[119], line_87[117], line_86[115], line_85[113], line_84[111], line_83[109], line_82[107], line_81[105], line_80[103], line_79[101], line_78[99], line_77[97], line_76[95], line_75[93], line_74[91], line_73[89], line_72[87], line_71[85], line_70[83], line_69[81], line_68[79], line_67[77], line_66[75], line_65[73], line_64[71], line_63[69], line_62[67], line_61[65], line_60[63], line_59[61], line_58[59], line_57[57], line_56[55], line_55[53], line_54[51], line_53[49], line_52[47], line_51[45], line_50[43], line_49[41], line_48[39], line_47[37], line_46[35], line_45[33], line_44[31], line_43[29], line_42[27], line_41[25], line_40[23], line_39[21], line_38[19], line_37[17], line_36[15], line_35[13], line_34[11], line_33[9], line_32[7], line_31[5], line_30[3], line_29[1], 28'b0};
assign col_200 = {line_128[200], line_127[198], line_126[196], line_125[194], line_124[192], line_123[190], line_122[188], line_121[186], line_120[184], line_119[182], line_118[180], line_117[178], line_116[176], line_115[174], line_114[172], line_113[170], line_112[168], line_111[166], line_110[164], line_109[162], line_108[160], line_107[158], line_106[156], line_105[154], line_104[152], line_103[150], line_102[148], line_101[146], line_100[144], line_99[142], line_98[140], line_97[138], line_96[136], line_95[134], line_94[132], line_93[130], line_92[128], line_91[126], line_90[124], line_89[122], line_88[120], line_87[118], line_86[116], line_85[114], line_84[112], line_83[110], line_82[108], line_81[106], line_80[104], line_79[102], line_78[100], line_77[98], line_76[96], line_75[94], line_74[92], line_73[90], line_72[88], line_71[86], line_70[84], line_69[82], line_68[80], line_67[78], line_66[76], line_65[74], line_64[72], line_63[70], line_62[68], line_61[66], line_60[64], line_59[62], line_58[60], line_57[58], line_56[56], line_55[54], line_54[52], line_53[50], line_52[48], line_51[46], line_50[44], line_49[42], line_48[40], line_47[38], line_46[36], line_45[34], line_44[32], line_43[30], line_42[28], line_41[26], line_40[24], line_39[22], line_38[20], line_37[18], line_36[16], line_35[14], line_34[12], line_33[10], line_32[8], line_31[6], line_30[4], line_29[2], line_28[0], 27'b0};
assign col_201 = {line_128[201], line_127[199], line_126[197], line_125[195], line_124[193], line_123[191], line_122[189], line_121[187], line_120[185], line_119[183], line_118[181], line_117[179], line_116[177], line_115[175], line_114[173], line_113[171], line_112[169], line_111[167], line_110[165], line_109[163], line_108[161], line_107[159], line_106[157], line_105[155], line_104[153], line_103[151], line_102[149], line_101[147], line_100[145], line_99[143], line_98[141], line_97[139], line_96[137], line_95[135], line_94[133], line_93[131], line_92[129], line_91[127], line_90[125], line_89[123], line_88[121], line_87[119], line_86[117], line_85[115], line_84[113], line_83[111], line_82[109], line_81[107], line_80[105], line_79[103], line_78[101], line_77[99], line_76[97], line_75[95], line_74[93], line_73[91], line_72[89], line_71[87], line_70[85], line_69[83], line_68[81], line_67[79], line_66[77], line_65[75], line_64[73], line_63[71], line_62[69], line_61[67], line_60[65], line_59[63], line_58[61], line_57[59], line_56[57], line_55[55], line_54[53], line_53[51], line_52[49], line_51[47], line_50[45], line_49[43], line_48[41], line_47[39], line_46[37], line_45[35], line_44[33], line_43[31], line_42[29], line_41[27], line_40[25], line_39[23], line_38[21], line_37[19], line_36[17], line_35[15], line_34[13], line_33[11], line_32[9], line_31[7], line_30[5], line_29[3], line_28[1], 27'b0};
assign col_202 = {line_128[202], line_127[200], line_126[198], line_125[196], line_124[194], line_123[192], line_122[190], line_121[188], line_120[186], line_119[184], line_118[182], line_117[180], line_116[178], line_115[176], line_114[174], line_113[172], line_112[170], line_111[168], line_110[166], line_109[164], line_108[162], line_107[160], line_106[158], line_105[156], line_104[154], line_103[152], line_102[150], line_101[148], line_100[146], line_99[144], line_98[142], line_97[140], line_96[138], line_95[136], line_94[134], line_93[132], line_92[130], line_91[128], line_90[126], line_89[124], line_88[122], line_87[120], line_86[118], line_85[116], line_84[114], line_83[112], line_82[110], line_81[108], line_80[106], line_79[104], line_78[102], line_77[100], line_76[98], line_75[96], line_74[94], line_73[92], line_72[90], line_71[88], line_70[86], line_69[84], line_68[82], line_67[80], line_66[78], line_65[76], line_64[74], line_63[72], line_62[70], line_61[68], line_60[66], line_59[64], line_58[62], line_57[60], line_56[58], line_55[56], line_54[54], line_53[52], line_52[50], line_51[48], line_50[46], line_49[44], line_48[42], line_47[40], line_46[38], line_45[36], line_44[34], line_43[32], line_42[30], line_41[28], line_40[26], line_39[24], line_38[22], line_37[20], line_36[18], line_35[16], line_34[14], line_33[12], line_32[10], line_31[8], line_30[6], line_29[4], line_28[2], line_27[0], 26'b0};
assign col_203 = {line_128[203], line_127[201], line_126[199], line_125[197], line_124[195], line_123[193], line_122[191], line_121[189], line_120[187], line_119[185], line_118[183], line_117[181], line_116[179], line_115[177], line_114[175], line_113[173], line_112[171], line_111[169], line_110[167], line_109[165], line_108[163], line_107[161], line_106[159], line_105[157], line_104[155], line_103[153], line_102[151], line_101[149], line_100[147], line_99[145], line_98[143], line_97[141], line_96[139], line_95[137], line_94[135], line_93[133], line_92[131], line_91[129], line_90[127], line_89[125], line_88[123], line_87[121], line_86[119], line_85[117], line_84[115], line_83[113], line_82[111], line_81[109], line_80[107], line_79[105], line_78[103], line_77[101], line_76[99], line_75[97], line_74[95], line_73[93], line_72[91], line_71[89], line_70[87], line_69[85], line_68[83], line_67[81], line_66[79], line_65[77], line_64[75], line_63[73], line_62[71], line_61[69], line_60[67], line_59[65], line_58[63], line_57[61], line_56[59], line_55[57], line_54[55], line_53[53], line_52[51], line_51[49], line_50[47], line_49[45], line_48[43], line_47[41], line_46[39], line_45[37], line_44[35], line_43[33], line_42[31], line_41[29], line_40[27], line_39[25], line_38[23], line_37[21], line_36[19], line_35[17], line_34[15], line_33[13], line_32[11], line_31[9], line_30[7], line_29[5], line_28[3], line_27[1], 26'b0};
assign col_204 = {line_128[204], line_127[202], line_126[200], line_125[198], line_124[196], line_123[194], line_122[192], line_121[190], line_120[188], line_119[186], line_118[184], line_117[182], line_116[180], line_115[178], line_114[176], line_113[174], line_112[172], line_111[170], line_110[168], line_109[166], line_108[164], line_107[162], line_106[160], line_105[158], line_104[156], line_103[154], line_102[152], line_101[150], line_100[148], line_99[146], line_98[144], line_97[142], line_96[140], line_95[138], line_94[136], line_93[134], line_92[132], line_91[130], line_90[128], line_89[126], line_88[124], line_87[122], line_86[120], line_85[118], line_84[116], line_83[114], line_82[112], line_81[110], line_80[108], line_79[106], line_78[104], line_77[102], line_76[100], line_75[98], line_74[96], line_73[94], line_72[92], line_71[90], line_70[88], line_69[86], line_68[84], line_67[82], line_66[80], line_65[78], line_64[76], line_63[74], line_62[72], line_61[70], line_60[68], line_59[66], line_58[64], line_57[62], line_56[60], line_55[58], line_54[56], line_53[54], line_52[52], line_51[50], line_50[48], line_49[46], line_48[44], line_47[42], line_46[40], line_45[38], line_44[36], line_43[34], line_42[32], line_41[30], line_40[28], line_39[26], line_38[24], line_37[22], line_36[20], line_35[18], line_34[16], line_33[14], line_32[12], line_31[10], line_30[8], line_29[6], line_28[4], line_27[2], line_26[0], 25'b0};
assign col_205 = {line_128[205], line_127[203], line_126[201], line_125[199], line_124[197], line_123[195], line_122[193], line_121[191], line_120[189], line_119[187], line_118[185], line_117[183], line_116[181], line_115[179], line_114[177], line_113[175], line_112[173], line_111[171], line_110[169], line_109[167], line_108[165], line_107[163], line_106[161], line_105[159], line_104[157], line_103[155], line_102[153], line_101[151], line_100[149], line_99[147], line_98[145], line_97[143], line_96[141], line_95[139], line_94[137], line_93[135], line_92[133], line_91[131], line_90[129], line_89[127], line_88[125], line_87[123], line_86[121], line_85[119], line_84[117], line_83[115], line_82[113], line_81[111], line_80[109], line_79[107], line_78[105], line_77[103], line_76[101], line_75[99], line_74[97], line_73[95], line_72[93], line_71[91], line_70[89], line_69[87], line_68[85], line_67[83], line_66[81], line_65[79], line_64[77], line_63[75], line_62[73], line_61[71], line_60[69], line_59[67], line_58[65], line_57[63], line_56[61], line_55[59], line_54[57], line_53[55], line_52[53], line_51[51], line_50[49], line_49[47], line_48[45], line_47[43], line_46[41], line_45[39], line_44[37], line_43[35], line_42[33], line_41[31], line_40[29], line_39[27], line_38[25], line_37[23], line_36[21], line_35[19], line_34[17], line_33[15], line_32[13], line_31[11], line_30[9], line_29[7], line_28[5], line_27[3], line_26[1], 25'b0};
assign col_206 = {line_128[206], line_127[204], line_126[202], line_125[200], line_124[198], line_123[196], line_122[194], line_121[192], line_120[190], line_119[188], line_118[186], line_117[184], line_116[182], line_115[180], line_114[178], line_113[176], line_112[174], line_111[172], line_110[170], line_109[168], line_108[166], line_107[164], line_106[162], line_105[160], line_104[158], line_103[156], line_102[154], line_101[152], line_100[150], line_99[148], line_98[146], line_97[144], line_96[142], line_95[140], line_94[138], line_93[136], line_92[134], line_91[132], line_90[130], line_89[128], line_88[126], line_87[124], line_86[122], line_85[120], line_84[118], line_83[116], line_82[114], line_81[112], line_80[110], line_79[108], line_78[106], line_77[104], line_76[102], line_75[100], line_74[98], line_73[96], line_72[94], line_71[92], line_70[90], line_69[88], line_68[86], line_67[84], line_66[82], line_65[80], line_64[78], line_63[76], line_62[74], line_61[72], line_60[70], line_59[68], line_58[66], line_57[64], line_56[62], line_55[60], line_54[58], line_53[56], line_52[54], line_51[52], line_50[50], line_49[48], line_48[46], line_47[44], line_46[42], line_45[40], line_44[38], line_43[36], line_42[34], line_41[32], line_40[30], line_39[28], line_38[26], line_37[24], line_36[22], line_35[20], line_34[18], line_33[16], line_32[14], line_31[12], line_30[10], line_29[8], line_28[6], line_27[4], line_26[2], line_25[0], 24'b0};
assign col_207 = {line_128[207], line_127[205], line_126[203], line_125[201], line_124[199], line_123[197], line_122[195], line_121[193], line_120[191], line_119[189], line_118[187], line_117[185], line_116[183], line_115[181], line_114[179], line_113[177], line_112[175], line_111[173], line_110[171], line_109[169], line_108[167], line_107[165], line_106[163], line_105[161], line_104[159], line_103[157], line_102[155], line_101[153], line_100[151], line_99[149], line_98[147], line_97[145], line_96[143], line_95[141], line_94[139], line_93[137], line_92[135], line_91[133], line_90[131], line_89[129], line_88[127], line_87[125], line_86[123], line_85[121], line_84[119], line_83[117], line_82[115], line_81[113], line_80[111], line_79[109], line_78[107], line_77[105], line_76[103], line_75[101], line_74[99], line_73[97], line_72[95], line_71[93], line_70[91], line_69[89], line_68[87], line_67[85], line_66[83], line_65[81], line_64[79], line_63[77], line_62[75], line_61[73], line_60[71], line_59[69], line_58[67], line_57[65], line_56[63], line_55[61], line_54[59], line_53[57], line_52[55], line_51[53], line_50[51], line_49[49], line_48[47], line_47[45], line_46[43], line_45[41], line_44[39], line_43[37], line_42[35], line_41[33], line_40[31], line_39[29], line_38[27], line_37[25], line_36[23], line_35[21], line_34[19], line_33[17], line_32[15], line_31[13], line_30[11], line_29[9], line_28[7], line_27[5], line_26[3], line_25[1], 24'b0};
assign col_208 = {line_128[208], line_127[206], line_126[204], line_125[202], line_124[200], line_123[198], line_122[196], line_121[194], line_120[192], line_119[190], line_118[188], line_117[186], line_116[184], line_115[182], line_114[180], line_113[178], line_112[176], line_111[174], line_110[172], line_109[170], line_108[168], line_107[166], line_106[164], line_105[162], line_104[160], line_103[158], line_102[156], line_101[154], line_100[152], line_99[150], line_98[148], line_97[146], line_96[144], line_95[142], line_94[140], line_93[138], line_92[136], line_91[134], line_90[132], line_89[130], line_88[128], line_87[126], line_86[124], line_85[122], line_84[120], line_83[118], line_82[116], line_81[114], line_80[112], line_79[110], line_78[108], line_77[106], line_76[104], line_75[102], line_74[100], line_73[98], line_72[96], line_71[94], line_70[92], line_69[90], line_68[88], line_67[86], line_66[84], line_65[82], line_64[80], line_63[78], line_62[76], line_61[74], line_60[72], line_59[70], line_58[68], line_57[66], line_56[64], line_55[62], line_54[60], line_53[58], line_52[56], line_51[54], line_50[52], line_49[50], line_48[48], line_47[46], line_46[44], line_45[42], line_44[40], line_43[38], line_42[36], line_41[34], line_40[32], line_39[30], line_38[28], line_37[26], line_36[24], line_35[22], line_34[20], line_33[18], line_32[16], line_31[14], line_30[12], line_29[10], line_28[8], line_27[6], line_26[4], line_25[2], line_24[0], 23'b0};
assign col_209 = {line_128[209], line_127[207], line_126[205], line_125[203], line_124[201], line_123[199], line_122[197], line_121[195], line_120[193], line_119[191], line_118[189], line_117[187], line_116[185], line_115[183], line_114[181], line_113[179], line_112[177], line_111[175], line_110[173], line_109[171], line_108[169], line_107[167], line_106[165], line_105[163], line_104[161], line_103[159], line_102[157], line_101[155], line_100[153], line_99[151], line_98[149], line_97[147], line_96[145], line_95[143], line_94[141], line_93[139], line_92[137], line_91[135], line_90[133], line_89[131], line_88[129], line_87[127], line_86[125], line_85[123], line_84[121], line_83[119], line_82[117], line_81[115], line_80[113], line_79[111], line_78[109], line_77[107], line_76[105], line_75[103], line_74[101], line_73[99], line_72[97], line_71[95], line_70[93], line_69[91], line_68[89], line_67[87], line_66[85], line_65[83], line_64[81], line_63[79], line_62[77], line_61[75], line_60[73], line_59[71], line_58[69], line_57[67], line_56[65], line_55[63], line_54[61], line_53[59], line_52[57], line_51[55], line_50[53], line_49[51], line_48[49], line_47[47], line_46[45], line_45[43], line_44[41], line_43[39], line_42[37], line_41[35], line_40[33], line_39[31], line_38[29], line_37[27], line_36[25], line_35[23], line_34[21], line_33[19], line_32[17], line_31[15], line_30[13], line_29[11], line_28[9], line_27[7], line_26[5], line_25[3], line_24[1], 23'b0};
assign col_210 = {line_128[210], line_127[208], line_126[206], line_125[204], line_124[202], line_123[200], line_122[198], line_121[196], line_120[194], line_119[192], line_118[190], line_117[188], line_116[186], line_115[184], line_114[182], line_113[180], line_112[178], line_111[176], line_110[174], line_109[172], line_108[170], line_107[168], line_106[166], line_105[164], line_104[162], line_103[160], line_102[158], line_101[156], line_100[154], line_99[152], line_98[150], line_97[148], line_96[146], line_95[144], line_94[142], line_93[140], line_92[138], line_91[136], line_90[134], line_89[132], line_88[130], line_87[128], line_86[126], line_85[124], line_84[122], line_83[120], line_82[118], line_81[116], line_80[114], line_79[112], line_78[110], line_77[108], line_76[106], line_75[104], line_74[102], line_73[100], line_72[98], line_71[96], line_70[94], line_69[92], line_68[90], line_67[88], line_66[86], line_65[84], line_64[82], line_63[80], line_62[78], line_61[76], line_60[74], line_59[72], line_58[70], line_57[68], line_56[66], line_55[64], line_54[62], line_53[60], line_52[58], line_51[56], line_50[54], line_49[52], line_48[50], line_47[48], line_46[46], line_45[44], line_44[42], line_43[40], line_42[38], line_41[36], line_40[34], line_39[32], line_38[30], line_37[28], line_36[26], line_35[24], line_34[22], line_33[20], line_32[18], line_31[16], line_30[14], line_29[12], line_28[10], line_27[8], line_26[6], line_25[4], line_24[2], line_23[0], 22'b0};
assign col_211 = {line_128[211], line_127[209], line_126[207], line_125[205], line_124[203], line_123[201], line_122[199], line_121[197], line_120[195], line_119[193], line_118[191], line_117[189], line_116[187], line_115[185], line_114[183], line_113[181], line_112[179], line_111[177], line_110[175], line_109[173], line_108[171], line_107[169], line_106[167], line_105[165], line_104[163], line_103[161], line_102[159], line_101[157], line_100[155], line_99[153], line_98[151], line_97[149], line_96[147], line_95[145], line_94[143], line_93[141], line_92[139], line_91[137], line_90[135], line_89[133], line_88[131], line_87[129], line_86[127], line_85[125], line_84[123], line_83[121], line_82[119], line_81[117], line_80[115], line_79[113], line_78[111], line_77[109], line_76[107], line_75[105], line_74[103], line_73[101], line_72[99], line_71[97], line_70[95], line_69[93], line_68[91], line_67[89], line_66[87], line_65[85], line_64[83], line_63[81], line_62[79], line_61[77], line_60[75], line_59[73], line_58[71], line_57[69], line_56[67], line_55[65], line_54[63], line_53[61], line_52[59], line_51[57], line_50[55], line_49[53], line_48[51], line_47[49], line_46[47], line_45[45], line_44[43], line_43[41], line_42[39], line_41[37], line_40[35], line_39[33], line_38[31], line_37[29], line_36[27], line_35[25], line_34[23], line_33[21], line_32[19], line_31[17], line_30[15], line_29[13], line_28[11], line_27[9], line_26[7], line_25[5], line_24[3], line_23[1], 22'b0};
assign col_212 = {line_128[212], line_127[210], line_126[208], line_125[206], line_124[204], line_123[202], line_122[200], line_121[198], line_120[196], line_119[194], line_118[192], line_117[190], line_116[188], line_115[186], line_114[184], line_113[182], line_112[180], line_111[178], line_110[176], line_109[174], line_108[172], line_107[170], line_106[168], line_105[166], line_104[164], line_103[162], line_102[160], line_101[158], line_100[156], line_99[154], line_98[152], line_97[150], line_96[148], line_95[146], line_94[144], line_93[142], line_92[140], line_91[138], line_90[136], line_89[134], line_88[132], line_87[130], line_86[128], line_85[126], line_84[124], line_83[122], line_82[120], line_81[118], line_80[116], line_79[114], line_78[112], line_77[110], line_76[108], line_75[106], line_74[104], line_73[102], line_72[100], line_71[98], line_70[96], line_69[94], line_68[92], line_67[90], line_66[88], line_65[86], line_64[84], line_63[82], line_62[80], line_61[78], line_60[76], line_59[74], line_58[72], line_57[70], line_56[68], line_55[66], line_54[64], line_53[62], line_52[60], line_51[58], line_50[56], line_49[54], line_48[52], line_47[50], line_46[48], line_45[46], line_44[44], line_43[42], line_42[40], line_41[38], line_40[36], line_39[34], line_38[32], line_37[30], line_36[28], line_35[26], line_34[24], line_33[22], line_32[20], line_31[18], line_30[16], line_29[14], line_28[12], line_27[10], line_26[8], line_25[6], line_24[4], line_23[2], line_22[0], 21'b0};
assign col_213 = {line_128[213], line_127[211], line_126[209], line_125[207], line_124[205], line_123[203], line_122[201], line_121[199], line_120[197], line_119[195], line_118[193], line_117[191], line_116[189], line_115[187], line_114[185], line_113[183], line_112[181], line_111[179], line_110[177], line_109[175], line_108[173], line_107[171], line_106[169], line_105[167], line_104[165], line_103[163], line_102[161], line_101[159], line_100[157], line_99[155], line_98[153], line_97[151], line_96[149], line_95[147], line_94[145], line_93[143], line_92[141], line_91[139], line_90[137], line_89[135], line_88[133], line_87[131], line_86[129], line_85[127], line_84[125], line_83[123], line_82[121], line_81[119], line_80[117], line_79[115], line_78[113], line_77[111], line_76[109], line_75[107], line_74[105], line_73[103], line_72[101], line_71[99], line_70[97], line_69[95], line_68[93], line_67[91], line_66[89], line_65[87], line_64[85], line_63[83], line_62[81], line_61[79], line_60[77], line_59[75], line_58[73], line_57[71], line_56[69], line_55[67], line_54[65], line_53[63], line_52[61], line_51[59], line_50[57], line_49[55], line_48[53], line_47[51], line_46[49], line_45[47], line_44[45], line_43[43], line_42[41], line_41[39], line_40[37], line_39[35], line_38[33], line_37[31], line_36[29], line_35[27], line_34[25], line_33[23], line_32[21], line_31[19], line_30[17], line_29[15], line_28[13], line_27[11], line_26[9], line_25[7], line_24[5], line_23[3], line_22[1], 21'b0};
assign col_214 = {line_128[214], line_127[212], line_126[210], line_125[208], line_124[206], line_123[204], line_122[202], line_121[200], line_120[198], line_119[196], line_118[194], line_117[192], line_116[190], line_115[188], line_114[186], line_113[184], line_112[182], line_111[180], line_110[178], line_109[176], line_108[174], line_107[172], line_106[170], line_105[168], line_104[166], line_103[164], line_102[162], line_101[160], line_100[158], line_99[156], line_98[154], line_97[152], line_96[150], line_95[148], line_94[146], line_93[144], line_92[142], line_91[140], line_90[138], line_89[136], line_88[134], line_87[132], line_86[130], line_85[128], line_84[126], line_83[124], line_82[122], line_81[120], line_80[118], line_79[116], line_78[114], line_77[112], line_76[110], line_75[108], line_74[106], line_73[104], line_72[102], line_71[100], line_70[98], line_69[96], line_68[94], line_67[92], line_66[90], line_65[88], line_64[86], line_63[84], line_62[82], line_61[80], line_60[78], line_59[76], line_58[74], line_57[72], line_56[70], line_55[68], line_54[66], line_53[64], line_52[62], line_51[60], line_50[58], line_49[56], line_48[54], line_47[52], line_46[50], line_45[48], line_44[46], line_43[44], line_42[42], line_41[40], line_40[38], line_39[36], line_38[34], line_37[32], line_36[30], line_35[28], line_34[26], line_33[24], line_32[22], line_31[20], line_30[18], line_29[16], line_28[14], line_27[12], line_26[10], line_25[8], line_24[6], line_23[4], line_22[2], line_21[0], 20'b0};
assign col_215 = {line_128[215], line_127[213], line_126[211], line_125[209], line_124[207], line_123[205], line_122[203], line_121[201], line_120[199], line_119[197], line_118[195], line_117[193], line_116[191], line_115[189], line_114[187], line_113[185], line_112[183], line_111[181], line_110[179], line_109[177], line_108[175], line_107[173], line_106[171], line_105[169], line_104[167], line_103[165], line_102[163], line_101[161], line_100[159], line_99[157], line_98[155], line_97[153], line_96[151], line_95[149], line_94[147], line_93[145], line_92[143], line_91[141], line_90[139], line_89[137], line_88[135], line_87[133], line_86[131], line_85[129], line_84[127], line_83[125], line_82[123], line_81[121], line_80[119], line_79[117], line_78[115], line_77[113], line_76[111], line_75[109], line_74[107], line_73[105], line_72[103], line_71[101], line_70[99], line_69[97], line_68[95], line_67[93], line_66[91], line_65[89], line_64[87], line_63[85], line_62[83], line_61[81], line_60[79], line_59[77], line_58[75], line_57[73], line_56[71], line_55[69], line_54[67], line_53[65], line_52[63], line_51[61], line_50[59], line_49[57], line_48[55], line_47[53], line_46[51], line_45[49], line_44[47], line_43[45], line_42[43], line_41[41], line_40[39], line_39[37], line_38[35], line_37[33], line_36[31], line_35[29], line_34[27], line_33[25], line_32[23], line_31[21], line_30[19], line_29[17], line_28[15], line_27[13], line_26[11], line_25[9], line_24[7], line_23[5], line_22[3], line_21[1], 20'b0};
assign col_216 = {line_128[216], line_127[214], line_126[212], line_125[210], line_124[208], line_123[206], line_122[204], line_121[202], line_120[200], line_119[198], line_118[196], line_117[194], line_116[192], line_115[190], line_114[188], line_113[186], line_112[184], line_111[182], line_110[180], line_109[178], line_108[176], line_107[174], line_106[172], line_105[170], line_104[168], line_103[166], line_102[164], line_101[162], line_100[160], line_99[158], line_98[156], line_97[154], line_96[152], line_95[150], line_94[148], line_93[146], line_92[144], line_91[142], line_90[140], line_89[138], line_88[136], line_87[134], line_86[132], line_85[130], line_84[128], line_83[126], line_82[124], line_81[122], line_80[120], line_79[118], line_78[116], line_77[114], line_76[112], line_75[110], line_74[108], line_73[106], line_72[104], line_71[102], line_70[100], line_69[98], line_68[96], line_67[94], line_66[92], line_65[90], line_64[88], line_63[86], line_62[84], line_61[82], line_60[80], line_59[78], line_58[76], line_57[74], line_56[72], line_55[70], line_54[68], line_53[66], line_52[64], line_51[62], line_50[60], line_49[58], line_48[56], line_47[54], line_46[52], line_45[50], line_44[48], line_43[46], line_42[44], line_41[42], line_40[40], line_39[38], line_38[36], line_37[34], line_36[32], line_35[30], line_34[28], line_33[26], line_32[24], line_31[22], line_30[20], line_29[18], line_28[16], line_27[14], line_26[12], line_25[10], line_24[8], line_23[6], line_22[4], line_21[2], line_20[0], 19'b0};
assign col_217 = {line_128[217], line_127[215], line_126[213], line_125[211], line_124[209], line_123[207], line_122[205], line_121[203], line_120[201], line_119[199], line_118[197], line_117[195], line_116[193], line_115[191], line_114[189], line_113[187], line_112[185], line_111[183], line_110[181], line_109[179], line_108[177], line_107[175], line_106[173], line_105[171], line_104[169], line_103[167], line_102[165], line_101[163], line_100[161], line_99[159], line_98[157], line_97[155], line_96[153], line_95[151], line_94[149], line_93[147], line_92[145], line_91[143], line_90[141], line_89[139], line_88[137], line_87[135], line_86[133], line_85[131], line_84[129], line_83[127], line_82[125], line_81[123], line_80[121], line_79[119], line_78[117], line_77[115], line_76[113], line_75[111], line_74[109], line_73[107], line_72[105], line_71[103], line_70[101], line_69[99], line_68[97], line_67[95], line_66[93], line_65[91], line_64[89], line_63[87], line_62[85], line_61[83], line_60[81], line_59[79], line_58[77], line_57[75], line_56[73], line_55[71], line_54[69], line_53[67], line_52[65], line_51[63], line_50[61], line_49[59], line_48[57], line_47[55], line_46[53], line_45[51], line_44[49], line_43[47], line_42[45], line_41[43], line_40[41], line_39[39], line_38[37], line_37[35], line_36[33], line_35[31], line_34[29], line_33[27], line_32[25], line_31[23], line_30[21], line_29[19], line_28[17], line_27[15], line_26[13], line_25[11], line_24[9], line_23[7], line_22[5], line_21[3], line_20[1], 19'b0};
assign col_218 = {line_128[218], line_127[216], line_126[214], line_125[212], line_124[210], line_123[208], line_122[206], line_121[204], line_120[202], line_119[200], line_118[198], line_117[196], line_116[194], line_115[192], line_114[190], line_113[188], line_112[186], line_111[184], line_110[182], line_109[180], line_108[178], line_107[176], line_106[174], line_105[172], line_104[170], line_103[168], line_102[166], line_101[164], line_100[162], line_99[160], line_98[158], line_97[156], line_96[154], line_95[152], line_94[150], line_93[148], line_92[146], line_91[144], line_90[142], line_89[140], line_88[138], line_87[136], line_86[134], line_85[132], line_84[130], line_83[128], line_82[126], line_81[124], line_80[122], line_79[120], line_78[118], line_77[116], line_76[114], line_75[112], line_74[110], line_73[108], line_72[106], line_71[104], line_70[102], line_69[100], line_68[98], line_67[96], line_66[94], line_65[92], line_64[90], line_63[88], line_62[86], line_61[84], line_60[82], line_59[80], line_58[78], line_57[76], line_56[74], line_55[72], line_54[70], line_53[68], line_52[66], line_51[64], line_50[62], line_49[60], line_48[58], line_47[56], line_46[54], line_45[52], line_44[50], line_43[48], line_42[46], line_41[44], line_40[42], line_39[40], line_38[38], line_37[36], line_36[34], line_35[32], line_34[30], line_33[28], line_32[26], line_31[24], line_30[22], line_29[20], line_28[18], line_27[16], line_26[14], line_25[12], line_24[10], line_23[8], line_22[6], line_21[4], line_20[2], line_19[0], 18'b0};
assign col_219 = {line_128[219], line_127[217], line_126[215], line_125[213], line_124[211], line_123[209], line_122[207], line_121[205], line_120[203], line_119[201], line_118[199], line_117[197], line_116[195], line_115[193], line_114[191], line_113[189], line_112[187], line_111[185], line_110[183], line_109[181], line_108[179], line_107[177], line_106[175], line_105[173], line_104[171], line_103[169], line_102[167], line_101[165], line_100[163], line_99[161], line_98[159], line_97[157], line_96[155], line_95[153], line_94[151], line_93[149], line_92[147], line_91[145], line_90[143], line_89[141], line_88[139], line_87[137], line_86[135], line_85[133], line_84[131], line_83[129], line_82[127], line_81[125], line_80[123], line_79[121], line_78[119], line_77[117], line_76[115], line_75[113], line_74[111], line_73[109], line_72[107], line_71[105], line_70[103], line_69[101], line_68[99], line_67[97], line_66[95], line_65[93], line_64[91], line_63[89], line_62[87], line_61[85], line_60[83], line_59[81], line_58[79], line_57[77], line_56[75], line_55[73], line_54[71], line_53[69], line_52[67], line_51[65], line_50[63], line_49[61], line_48[59], line_47[57], line_46[55], line_45[53], line_44[51], line_43[49], line_42[47], line_41[45], line_40[43], line_39[41], line_38[39], line_37[37], line_36[35], line_35[33], line_34[31], line_33[29], line_32[27], line_31[25], line_30[23], line_29[21], line_28[19], line_27[17], line_26[15], line_25[13], line_24[11], line_23[9], line_22[7], line_21[5], line_20[3], line_19[1], 18'b0};
assign col_220 = {line_128[220], line_127[218], line_126[216], line_125[214], line_124[212], line_123[210], line_122[208], line_121[206], line_120[204], line_119[202], line_118[200], line_117[198], line_116[196], line_115[194], line_114[192], line_113[190], line_112[188], line_111[186], line_110[184], line_109[182], line_108[180], line_107[178], line_106[176], line_105[174], line_104[172], line_103[170], line_102[168], line_101[166], line_100[164], line_99[162], line_98[160], line_97[158], line_96[156], line_95[154], line_94[152], line_93[150], line_92[148], line_91[146], line_90[144], line_89[142], line_88[140], line_87[138], line_86[136], line_85[134], line_84[132], line_83[130], line_82[128], line_81[126], line_80[124], line_79[122], line_78[120], line_77[118], line_76[116], line_75[114], line_74[112], line_73[110], line_72[108], line_71[106], line_70[104], line_69[102], line_68[100], line_67[98], line_66[96], line_65[94], line_64[92], line_63[90], line_62[88], line_61[86], line_60[84], line_59[82], line_58[80], line_57[78], line_56[76], line_55[74], line_54[72], line_53[70], line_52[68], line_51[66], line_50[64], line_49[62], line_48[60], line_47[58], line_46[56], line_45[54], line_44[52], line_43[50], line_42[48], line_41[46], line_40[44], line_39[42], line_38[40], line_37[38], line_36[36], line_35[34], line_34[32], line_33[30], line_32[28], line_31[26], line_30[24], line_29[22], line_28[20], line_27[18], line_26[16], line_25[14], line_24[12], line_23[10], line_22[8], line_21[6], line_20[4], line_19[2], line_18[0], 17'b0};
assign col_221 = {line_128[221], line_127[219], line_126[217], line_125[215], line_124[213], line_123[211], line_122[209], line_121[207], line_120[205], line_119[203], line_118[201], line_117[199], line_116[197], line_115[195], line_114[193], line_113[191], line_112[189], line_111[187], line_110[185], line_109[183], line_108[181], line_107[179], line_106[177], line_105[175], line_104[173], line_103[171], line_102[169], line_101[167], line_100[165], line_99[163], line_98[161], line_97[159], line_96[157], line_95[155], line_94[153], line_93[151], line_92[149], line_91[147], line_90[145], line_89[143], line_88[141], line_87[139], line_86[137], line_85[135], line_84[133], line_83[131], line_82[129], line_81[127], line_80[125], line_79[123], line_78[121], line_77[119], line_76[117], line_75[115], line_74[113], line_73[111], line_72[109], line_71[107], line_70[105], line_69[103], line_68[101], line_67[99], line_66[97], line_65[95], line_64[93], line_63[91], line_62[89], line_61[87], line_60[85], line_59[83], line_58[81], line_57[79], line_56[77], line_55[75], line_54[73], line_53[71], line_52[69], line_51[67], line_50[65], line_49[63], line_48[61], line_47[59], line_46[57], line_45[55], line_44[53], line_43[51], line_42[49], line_41[47], line_40[45], line_39[43], line_38[41], line_37[39], line_36[37], line_35[35], line_34[33], line_33[31], line_32[29], line_31[27], line_30[25], line_29[23], line_28[21], line_27[19], line_26[17], line_25[15], line_24[13], line_23[11], line_22[9], line_21[7], line_20[5], line_19[3], line_18[1], 17'b0};
assign col_222 = {line_128[222], line_127[220], line_126[218], line_125[216], line_124[214], line_123[212], line_122[210], line_121[208], line_120[206], line_119[204], line_118[202], line_117[200], line_116[198], line_115[196], line_114[194], line_113[192], line_112[190], line_111[188], line_110[186], line_109[184], line_108[182], line_107[180], line_106[178], line_105[176], line_104[174], line_103[172], line_102[170], line_101[168], line_100[166], line_99[164], line_98[162], line_97[160], line_96[158], line_95[156], line_94[154], line_93[152], line_92[150], line_91[148], line_90[146], line_89[144], line_88[142], line_87[140], line_86[138], line_85[136], line_84[134], line_83[132], line_82[130], line_81[128], line_80[126], line_79[124], line_78[122], line_77[120], line_76[118], line_75[116], line_74[114], line_73[112], line_72[110], line_71[108], line_70[106], line_69[104], line_68[102], line_67[100], line_66[98], line_65[96], line_64[94], line_63[92], line_62[90], line_61[88], line_60[86], line_59[84], line_58[82], line_57[80], line_56[78], line_55[76], line_54[74], line_53[72], line_52[70], line_51[68], line_50[66], line_49[64], line_48[62], line_47[60], line_46[58], line_45[56], line_44[54], line_43[52], line_42[50], line_41[48], line_40[46], line_39[44], line_38[42], line_37[40], line_36[38], line_35[36], line_34[34], line_33[32], line_32[30], line_31[28], line_30[26], line_29[24], line_28[22], line_27[20], line_26[18], line_25[16], line_24[14], line_23[12], line_22[10], line_21[8], line_20[6], line_19[4], line_18[2], line_17[0], 16'b0};
assign col_223 = {line_128[223], line_127[221], line_126[219], line_125[217], line_124[215], line_123[213], line_122[211], line_121[209], line_120[207], line_119[205], line_118[203], line_117[201], line_116[199], line_115[197], line_114[195], line_113[193], line_112[191], line_111[189], line_110[187], line_109[185], line_108[183], line_107[181], line_106[179], line_105[177], line_104[175], line_103[173], line_102[171], line_101[169], line_100[167], line_99[165], line_98[163], line_97[161], line_96[159], line_95[157], line_94[155], line_93[153], line_92[151], line_91[149], line_90[147], line_89[145], line_88[143], line_87[141], line_86[139], line_85[137], line_84[135], line_83[133], line_82[131], line_81[129], line_80[127], line_79[125], line_78[123], line_77[121], line_76[119], line_75[117], line_74[115], line_73[113], line_72[111], line_71[109], line_70[107], line_69[105], line_68[103], line_67[101], line_66[99], line_65[97], line_64[95], line_63[93], line_62[91], line_61[89], line_60[87], line_59[85], line_58[83], line_57[81], line_56[79], line_55[77], line_54[75], line_53[73], line_52[71], line_51[69], line_50[67], line_49[65], line_48[63], line_47[61], line_46[59], line_45[57], line_44[55], line_43[53], line_42[51], line_41[49], line_40[47], line_39[45], line_38[43], line_37[41], line_36[39], line_35[37], line_34[35], line_33[33], line_32[31], line_31[29], line_30[27], line_29[25], line_28[23], line_27[21], line_26[19], line_25[17], line_24[15], line_23[13], line_22[11], line_21[9], line_20[7], line_19[5], line_18[3], line_17[1], 16'b0};
assign col_224 = {line_128[224], line_127[222], line_126[220], line_125[218], line_124[216], line_123[214], line_122[212], line_121[210], line_120[208], line_119[206], line_118[204], line_117[202], line_116[200], line_115[198], line_114[196], line_113[194], line_112[192], line_111[190], line_110[188], line_109[186], line_108[184], line_107[182], line_106[180], line_105[178], line_104[176], line_103[174], line_102[172], line_101[170], line_100[168], line_99[166], line_98[164], line_97[162], line_96[160], line_95[158], line_94[156], line_93[154], line_92[152], line_91[150], line_90[148], line_89[146], line_88[144], line_87[142], line_86[140], line_85[138], line_84[136], line_83[134], line_82[132], line_81[130], line_80[128], line_79[126], line_78[124], line_77[122], line_76[120], line_75[118], line_74[116], line_73[114], line_72[112], line_71[110], line_70[108], line_69[106], line_68[104], line_67[102], line_66[100], line_65[98], line_64[96], line_63[94], line_62[92], line_61[90], line_60[88], line_59[86], line_58[84], line_57[82], line_56[80], line_55[78], line_54[76], line_53[74], line_52[72], line_51[70], line_50[68], line_49[66], line_48[64], line_47[62], line_46[60], line_45[58], line_44[56], line_43[54], line_42[52], line_41[50], line_40[48], line_39[46], line_38[44], line_37[42], line_36[40], line_35[38], line_34[36], line_33[34], line_32[32], line_31[30], line_30[28], line_29[26], line_28[24], line_27[22], line_26[20], line_25[18], line_24[16], line_23[14], line_22[12], line_21[10], line_20[8], line_19[6], line_18[4], line_17[2], line_16[0], 15'b0};
assign col_225 = {line_128[225], line_127[223], line_126[221], line_125[219], line_124[217], line_123[215], line_122[213], line_121[211], line_120[209], line_119[207], line_118[205], line_117[203], line_116[201], line_115[199], line_114[197], line_113[195], line_112[193], line_111[191], line_110[189], line_109[187], line_108[185], line_107[183], line_106[181], line_105[179], line_104[177], line_103[175], line_102[173], line_101[171], line_100[169], line_99[167], line_98[165], line_97[163], line_96[161], line_95[159], line_94[157], line_93[155], line_92[153], line_91[151], line_90[149], line_89[147], line_88[145], line_87[143], line_86[141], line_85[139], line_84[137], line_83[135], line_82[133], line_81[131], line_80[129], line_79[127], line_78[125], line_77[123], line_76[121], line_75[119], line_74[117], line_73[115], line_72[113], line_71[111], line_70[109], line_69[107], line_68[105], line_67[103], line_66[101], line_65[99], line_64[97], line_63[95], line_62[93], line_61[91], line_60[89], line_59[87], line_58[85], line_57[83], line_56[81], line_55[79], line_54[77], line_53[75], line_52[73], line_51[71], line_50[69], line_49[67], line_48[65], line_47[63], line_46[61], line_45[59], line_44[57], line_43[55], line_42[53], line_41[51], line_40[49], line_39[47], line_38[45], line_37[43], line_36[41], line_35[39], line_34[37], line_33[35], line_32[33], line_31[31], line_30[29], line_29[27], line_28[25], line_27[23], line_26[21], line_25[19], line_24[17], line_23[15], line_22[13], line_21[11], line_20[9], line_19[7], line_18[5], line_17[3], line_16[1], 15'b0};
assign col_226 = {line_128[226], line_127[224], line_126[222], line_125[220], line_124[218], line_123[216], line_122[214], line_121[212], line_120[210], line_119[208], line_118[206], line_117[204], line_116[202], line_115[200], line_114[198], line_113[196], line_112[194], line_111[192], line_110[190], line_109[188], line_108[186], line_107[184], line_106[182], line_105[180], line_104[178], line_103[176], line_102[174], line_101[172], line_100[170], line_99[168], line_98[166], line_97[164], line_96[162], line_95[160], line_94[158], line_93[156], line_92[154], line_91[152], line_90[150], line_89[148], line_88[146], line_87[144], line_86[142], line_85[140], line_84[138], line_83[136], line_82[134], line_81[132], line_80[130], line_79[128], line_78[126], line_77[124], line_76[122], line_75[120], line_74[118], line_73[116], line_72[114], line_71[112], line_70[110], line_69[108], line_68[106], line_67[104], line_66[102], line_65[100], line_64[98], line_63[96], line_62[94], line_61[92], line_60[90], line_59[88], line_58[86], line_57[84], line_56[82], line_55[80], line_54[78], line_53[76], line_52[74], line_51[72], line_50[70], line_49[68], line_48[66], line_47[64], line_46[62], line_45[60], line_44[58], line_43[56], line_42[54], line_41[52], line_40[50], line_39[48], line_38[46], line_37[44], line_36[42], line_35[40], line_34[38], line_33[36], line_32[34], line_31[32], line_30[30], line_29[28], line_28[26], line_27[24], line_26[22], line_25[20], line_24[18], line_23[16], line_22[14], line_21[12], line_20[10], line_19[8], line_18[6], line_17[4], line_16[2], line_15[0], 14'b0};
assign col_227 = {line_128[227], line_127[225], line_126[223], line_125[221], line_124[219], line_123[217], line_122[215], line_121[213], line_120[211], line_119[209], line_118[207], line_117[205], line_116[203], line_115[201], line_114[199], line_113[197], line_112[195], line_111[193], line_110[191], line_109[189], line_108[187], line_107[185], line_106[183], line_105[181], line_104[179], line_103[177], line_102[175], line_101[173], line_100[171], line_99[169], line_98[167], line_97[165], line_96[163], line_95[161], line_94[159], line_93[157], line_92[155], line_91[153], line_90[151], line_89[149], line_88[147], line_87[145], line_86[143], line_85[141], line_84[139], line_83[137], line_82[135], line_81[133], line_80[131], line_79[129], line_78[127], line_77[125], line_76[123], line_75[121], line_74[119], line_73[117], line_72[115], line_71[113], line_70[111], line_69[109], line_68[107], line_67[105], line_66[103], line_65[101], line_64[99], line_63[97], line_62[95], line_61[93], line_60[91], line_59[89], line_58[87], line_57[85], line_56[83], line_55[81], line_54[79], line_53[77], line_52[75], line_51[73], line_50[71], line_49[69], line_48[67], line_47[65], line_46[63], line_45[61], line_44[59], line_43[57], line_42[55], line_41[53], line_40[51], line_39[49], line_38[47], line_37[45], line_36[43], line_35[41], line_34[39], line_33[37], line_32[35], line_31[33], line_30[31], line_29[29], line_28[27], line_27[25], line_26[23], line_25[21], line_24[19], line_23[17], line_22[15], line_21[13], line_20[11], line_19[9], line_18[7], line_17[5], line_16[3], line_15[1], 14'b0};
assign col_228 = {line_128[228], line_127[226], line_126[224], line_125[222], line_124[220], line_123[218], line_122[216], line_121[214], line_120[212], line_119[210], line_118[208], line_117[206], line_116[204], line_115[202], line_114[200], line_113[198], line_112[196], line_111[194], line_110[192], line_109[190], line_108[188], line_107[186], line_106[184], line_105[182], line_104[180], line_103[178], line_102[176], line_101[174], line_100[172], line_99[170], line_98[168], line_97[166], line_96[164], line_95[162], line_94[160], line_93[158], line_92[156], line_91[154], line_90[152], line_89[150], line_88[148], line_87[146], line_86[144], line_85[142], line_84[140], line_83[138], line_82[136], line_81[134], line_80[132], line_79[130], line_78[128], line_77[126], line_76[124], line_75[122], line_74[120], line_73[118], line_72[116], line_71[114], line_70[112], line_69[110], line_68[108], line_67[106], line_66[104], line_65[102], line_64[100], line_63[98], line_62[96], line_61[94], line_60[92], line_59[90], line_58[88], line_57[86], line_56[84], line_55[82], line_54[80], line_53[78], line_52[76], line_51[74], line_50[72], line_49[70], line_48[68], line_47[66], line_46[64], line_45[62], line_44[60], line_43[58], line_42[56], line_41[54], line_40[52], line_39[50], line_38[48], line_37[46], line_36[44], line_35[42], line_34[40], line_33[38], line_32[36], line_31[34], line_30[32], line_29[30], line_28[28], line_27[26], line_26[24], line_25[22], line_24[20], line_23[18], line_22[16], line_21[14], line_20[12], line_19[10], line_18[8], line_17[6], line_16[4], line_15[2], line_14[0], 13'b0};
assign col_229 = {line_128[229], line_127[227], line_126[225], line_125[223], line_124[221], line_123[219], line_122[217], line_121[215], line_120[213], line_119[211], line_118[209], line_117[207], line_116[205], line_115[203], line_114[201], line_113[199], line_112[197], line_111[195], line_110[193], line_109[191], line_108[189], line_107[187], line_106[185], line_105[183], line_104[181], line_103[179], line_102[177], line_101[175], line_100[173], line_99[171], line_98[169], line_97[167], line_96[165], line_95[163], line_94[161], line_93[159], line_92[157], line_91[155], line_90[153], line_89[151], line_88[149], line_87[147], line_86[145], line_85[143], line_84[141], line_83[139], line_82[137], line_81[135], line_80[133], line_79[131], line_78[129], line_77[127], line_76[125], line_75[123], line_74[121], line_73[119], line_72[117], line_71[115], line_70[113], line_69[111], line_68[109], line_67[107], line_66[105], line_65[103], line_64[101], line_63[99], line_62[97], line_61[95], line_60[93], line_59[91], line_58[89], line_57[87], line_56[85], line_55[83], line_54[81], line_53[79], line_52[77], line_51[75], line_50[73], line_49[71], line_48[69], line_47[67], line_46[65], line_45[63], line_44[61], line_43[59], line_42[57], line_41[55], line_40[53], line_39[51], line_38[49], line_37[47], line_36[45], line_35[43], line_34[41], line_33[39], line_32[37], line_31[35], line_30[33], line_29[31], line_28[29], line_27[27], line_26[25], line_25[23], line_24[21], line_23[19], line_22[17], line_21[15], line_20[13], line_19[11], line_18[9], line_17[7], line_16[5], line_15[3], line_14[1], 13'b0};
assign col_230 = {line_128[230], line_127[228], line_126[226], line_125[224], line_124[222], line_123[220], line_122[218], line_121[216], line_120[214], line_119[212], line_118[210], line_117[208], line_116[206], line_115[204], line_114[202], line_113[200], line_112[198], line_111[196], line_110[194], line_109[192], line_108[190], line_107[188], line_106[186], line_105[184], line_104[182], line_103[180], line_102[178], line_101[176], line_100[174], line_99[172], line_98[170], line_97[168], line_96[166], line_95[164], line_94[162], line_93[160], line_92[158], line_91[156], line_90[154], line_89[152], line_88[150], line_87[148], line_86[146], line_85[144], line_84[142], line_83[140], line_82[138], line_81[136], line_80[134], line_79[132], line_78[130], line_77[128], line_76[126], line_75[124], line_74[122], line_73[120], line_72[118], line_71[116], line_70[114], line_69[112], line_68[110], line_67[108], line_66[106], line_65[104], line_64[102], line_63[100], line_62[98], line_61[96], line_60[94], line_59[92], line_58[90], line_57[88], line_56[86], line_55[84], line_54[82], line_53[80], line_52[78], line_51[76], line_50[74], line_49[72], line_48[70], line_47[68], line_46[66], line_45[64], line_44[62], line_43[60], line_42[58], line_41[56], line_40[54], line_39[52], line_38[50], line_37[48], line_36[46], line_35[44], line_34[42], line_33[40], line_32[38], line_31[36], line_30[34], line_29[32], line_28[30], line_27[28], line_26[26], line_25[24], line_24[22], line_23[20], line_22[18], line_21[16], line_20[14], line_19[12], line_18[10], line_17[8], line_16[6], line_15[4], line_14[2], line_13[0], 12'b0};
assign col_231 = {line_128[231], line_127[229], line_126[227], line_125[225], line_124[223], line_123[221], line_122[219], line_121[217], line_120[215], line_119[213], line_118[211], line_117[209], line_116[207], line_115[205], line_114[203], line_113[201], line_112[199], line_111[197], line_110[195], line_109[193], line_108[191], line_107[189], line_106[187], line_105[185], line_104[183], line_103[181], line_102[179], line_101[177], line_100[175], line_99[173], line_98[171], line_97[169], line_96[167], line_95[165], line_94[163], line_93[161], line_92[159], line_91[157], line_90[155], line_89[153], line_88[151], line_87[149], line_86[147], line_85[145], line_84[143], line_83[141], line_82[139], line_81[137], line_80[135], line_79[133], line_78[131], line_77[129], line_76[127], line_75[125], line_74[123], line_73[121], line_72[119], line_71[117], line_70[115], line_69[113], line_68[111], line_67[109], line_66[107], line_65[105], line_64[103], line_63[101], line_62[99], line_61[97], line_60[95], line_59[93], line_58[91], line_57[89], line_56[87], line_55[85], line_54[83], line_53[81], line_52[79], line_51[77], line_50[75], line_49[73], line_48[71], line_47[69], line_46[67], line_45[65], line_44[63], line_43[61], line_42[59], line_41[57], line_40[55], line_39[53], line_38[51], line_37[49], line_36[47], line_35[45], line_34[43], line_33[41], line_32[39], line_31[37], line_30[35], line_29[33], line_28[31], line_27[29], line_26[27], line_25[25], line_24[23], line_23[21], line_22[19], line_21[17], line_20[15], line_19[13], line_18[11], line_17[9], line_16[7], line_15[5], line_14[3], line_13[1], 12'b0};
assign col_232 = {line_128[232], line_127[230], line_126[228], line_125[226], line_124[224], line_123[222], line_122[220], line_121[218], line_120[216], line_119[214], line_118[212], line_117[210], line_116[208], line_115[206], line_114[204], line_113[202], line_112[200], line_111[198], line_110[196], line_109[194], line_108[192], line_107[190], line_106[188], line_105[186], line_104[184], line_103[182], line_102[180], line_101[178], line_100[176], line_99[174], line_98[172], line_97[170], line_96[168], line_95[166], line_94[164], line_93[162], line_92[160], line_91[158], line_90[156], line_89[154], line_88[152], line_87[150], line_86[148], line_85[146], line_84[144], line_83[142], line_82[140], line_81[138], line_80[136], line_79[134], line_78[132], line_77[130], line_76[128], line_75[126], line_74[124], line_73[122], line_72[120], line_71[118], line_70[116], line_69[114], line_68[112], line_67[110], line_66[108], line_65[106], line_64[104], line_63[102], line_62[100], line_61[98], line_60[96], line_59[94], line_58[92], line_57[90], line_56[88], line_55[86], line_54[84], line_53[82], line_52[80], line_51[78], line_50[76], line_49[74], line_48[72], line_47[70], line_46[68], line_45[66], line_44[64], line_43[62], line_42[60], line_41[58], line_40[56], line_39[54], line_38[52], line_37[50], line_36[48], line_35[46], line_34[44], line_33[42], line_32[40], line_31[38], line_30[36], line_29[34], line_28[32], line_27[30], line_26[28], line_25[26], line_24[24], line_23[22], line_22[20], line_21[18], line_20[16], line_19[14], line_18[12], line_17[10], line_16[8], line_15[6], line_14[4], line_13[2], line_12[0], 11'b0};
assign col_233 = {line_128[233], line_127[231], line_126[229], line_125[227], line_124[225], line_123[223], line_122[221], line_121[219], line_120[217], line_119[215], line_118[213], line_117[211], line_116[209], line_115[207], line_114[205], line_113[203], line_112[201], line_111[199], line_110[197], line_109[195], line_108[193], line_107[191], line_106[189], line_105[187], line_104[185], line_103[183], line_102[181], line_101[179], line_100[177], line_99[175], line_98[173], line_97[171], line_96[169], line_95[167], line_94[165], line_93[163], line_92[161], line_91[159], line_90[157], line_89[155], line_88[153], line_87[151], line_86[149], line_85[147], line_84[145], line_83[143], line_82[141], line_81[139], line_80[137], line_79[135], line_78[133], line_77[131], line_76[129], line_75[127], line_74[125], line_73[123], line_72[121], line_71[119], line_70[117], line_69[115], line_68[113], line_67[111], line_66[109], line_65[107], line_64[105], line_63[103], line_62[101], line_61[99], line_60[97], line_59[95], line_58[93], line_57[91], line_56[89], line_55[87], line_54[85], line_53[83], line_52[81], line_51[79], line_50[77], line_49[75], line_48[73], line_47[71], line_46[69], line_45[67], line_44[65], line_43[63], line_42[61], line_41[59], line_40[57], line_39[55], line_38[53], line_37[51], line_36[49], line_35[47], line_34[45], line_33[43], line_32[41], line_31[39], line_30[37], line_29[35], line_28[33], line_27[31], line_26[29], line_25[27], line_24[25], line_23[23], line_22[21], line_21[19], line_20[17], line_19[15], line_18[13], line_17[11], line_16[9], line_15[7], line_14[5], line_13[3], line_12[1], 11'b0};
assign col_234 = {line_128[234], line_127[232], line_126[230], line_125[228], line_124[226], line_123[224], line_122[222], line_121[220], line_120[218], line_119[216], line_118[214], line_117[212], line_116[210], line_115[208], line_114[206], line_113[204], line_112[202], line_111[200], line_110[198], line_109[196], line_108[194], line_107[192], line_106[190], line_105[188], line_104[186], line_103[184], line_102[182], line_101[180], line_100[178], line_99[176], line_98[174], line_97[172], line_96[170], line_95[168], line_94[166], line_93[164], line_92[162], line_91[160], line_90[158], line_89[156], line_88[154], line_87[152], line_86[150], line_85[148], line_84[146], line_83[144], line_82[142], line_81[140], line_80[138], line_79[136], line_78[134], line_77[132], line_76[130], line_75[128], line_74[126], line_73[124], line_72[122], line_71[120], line_70[118], line_69[116], line_68[114], line_67[112], line_66[110], line_65[108], line_64[106], line_63[104], line_62[102], line_61[100], line_60[98], line_59[96], line_58[94], line_57[92], line_56[90], line_55[88], line_54[86], line_53[84], line_52[82], line_51[80], line_50[78], line_49[76], line_48[74], line_47[72], line_46[70], line_45[68], line_44[66], line_43[64], line_42[62], line_41[60], line_40[58], line_39[56], line_38[54], line_37[52], line_36[50], line_35[48], line_34[46], line_33[44], line_32[42], line_31[40], line_30[38], line_29[36], line_28[34], line_27[32], line_26[30], line_25[28], line_24[26], line_23[24], line_22[22], line_21[20], line_20[18], line_19[16], line_18[14], line_17[12], line_16[10], line_15[8], line_14[6], line_13[4], line_12[2], line_11[0], 10'b0};
assign col_235 = {line_128[235], line_127[233], line_126[231], line_125[229], line_124[227], line_123[225], line_122[223], line_121[221], line_120[219], line_119[217], line_118[215], line_117[213], line_116[211], line_115[209], line_114[207], line_113[205], line_112[203], line_111[201], line_110[199], line_109[197], line_108[195], line_107[193], line_106[191], line_105[189], line_104[187], line_103[185], line_102[183], line_101[181], line_100[179], line_99[177], line_98[175], line_97[173], line_96[171], line_95[169], line_94[167], line_93[165], line_92[163], line_91[161], line_90[159], line_89[157], line_88[155], line_87[153], line_86[151], line_85[149], line_84[147], line_83[145], line_82[143], line_81[141], line_80[139], line_79[137], line_78[135], line_77[133], line_76[131], line_75[129], line_74[127], line_73[125], line_72[123], line_71[121], line_70[119], line_69[117], line_68[115], line_67[113], line_66[111], line_65[109], line_64[107], line_63[105], line_62[103], line_61[101], line_60[99], line_59[97], line_58[95], line_57[93], line_56[91], line_55[89], line_54[87], line_53[85], line_52[83], line_51[81], line_50[79], line_49[77], line_48[75], line_47[73], line_46[71], line_45[69], line_44[67], line_43[65], line_42[63], line_41[61], line_40[59], line_39[57], line_38[55], line_37[53], line_36[51], line_35[49], line_34[47], line_33[45], line_32[43], line_31[41], line_30[39], line_29[37], line_28[35], line_27[33], line_26[31], line_25[29], line_24[27], line_23[25], line_22[23], line_21[21], line_20[19], line_19[17], line_18[15], line_17[13], line_16[11], line_15[9], line_14[7], line_13[5], line_12[3], line_11[1], 10'b0};
assign col_236 = {line_128[236], line_127[234], line_126[232], line_125[230], line_124[228], line_123[226], line_122[224], line_121[222], line_120[220], line_119[218], line_118[216], line_117[214], line_116[212], line_115[210], line_114[208], line_113[206], line_112[204], line_111[202], line_110[200], line_109[198], line_108[196], line_107[194], line_106[192], line_105[190], line_104[188], line_103[186], line_102[184], line_101[182], line_100[180], line_99[178], line_98[176], line_97[174], line_96[172], line_95[170], line_94[168], line_93[166], line_92[164], line_91[162], line_90[160], line_89[158], line_88[156], line_87[154], line_86[152], line_85[150], line_84[148], line_83[146], line_82[144], line_81[142], line_80[140], line_79[138], line_78[136], line_77[134], line_76[132], line_75[130], line_74[128], line_73[126], line_72[124], line_71[122], line_70[120], line_69[118], line_68[116], line_67[114], line_66[112], line_65[110], line_64[108], line_63[106], line_62[104], line_61[102], line_60[100], line_59[98], line_58[96], line_57[94], line_56[92], line_55[90], line_54[88], line_53[86], line_52[84], line_51[82], line_50[80], line_49[78], line_48[76], line_47[74], line_46[72], line_45[70], line_44[68], line_43[66], line_42[64], line_41[62], line_40[60], line_39[58], line_38[56], line_37[54], line_36[52], line_35[50], line_34[48], line_33[46], line_32[44], line_31[42], line_30[40], line_29[38], line_28[36], line_27[34], line_26[32], line_25[30], line_24[28], line_23[26], line_22[24], line_21[22], line_20[20], line_19[18], line_18[16], line_17[14], line_16[12], line_15[10], line_14[8], line_13[6], line_12[4], line_11[2], line_10[0], 9'b0};
assign col_237 = {line_128[237], line_127[235], line_126[233], line_125[231], line_124[229], line_123[227], line_122[225], line_121[223], line_120[221], line_119[219], line_118[217], line_117[215], line_116[213], line_115[211], line_114[209], line_113[207], line_112[205], line_111[203], line_110[201], line_109[199], line_108[197], line_107[195], line_106[193], line_105[191], line_104[189], line_103[187], line_102[185], line_101[183], line_100[181], line_99[179], line_98[177], line_97[175], line_96[173], line_95[171], line_94[169], line_93[167], line_92[165], line_91[163], line_90[161], line_89[159], line_88[157], line_87[155], line_86[153], line_85[151], line_84[149], line_83[147], line_82[145], line_81[143], line_80[141], line_79[139], line_78[137], line_77[135], line_76[133], line_75[131], line_74[129], line_73[127], line_72[125], line_71[123], line_70[121], line_69[119], line_68[117], line_67[115], line_66[113], line_65[111], line_64[109], line_63[107], line_62[105], line_61[103], line_60[101], line_59[99], line_58[97], line_57[95], line_56[93], line_55[91], line_54[89], line_53[87], line_52[85], line_51[83], line_50[81], line_49[79], line_48[77], line_47[75], line_46[73], line_45[71], line_44[69], line_43[67], line_42[65], line_41[63], line_40[61], line_39[59], line_38[57], line_37[55], line_36[53], line_35[51], line_34[49], line_33[47], line_32[45], line_31[43], line_30[41], line_29[39], line_28[37], line_27[35], line_26[33], line_25[31], line_24[29], line_23[27], line_22[25], line_21[23], line_20[21], line_19[19], line_18[17], line_17[15], line_16[13], line_15[11], line_14[9], line_13[7], line_12[5], line_11[3], line_10[1], 9'b0};
assign col_238 = {line_128[238], line_127[236], line_126[234], line_125[232], line_124[230], line_123[228], line_122[226], line_121[224], line_120[222], line_119[220], line_118[218], line_117[216], line_116[214], line_115[212], line_114[210], line_113[208], line_112[206], line_111[204], line_110[202], line_109[200], line_108[198], line_107[196], line_106[194], line_105[192], line_104[190], line_103[188], line_102[186], line_101[184], line_100[182], line_99[180], line_98[178], line_97[176], line_96[174], line_95[172], line_94[170], line_93[168], line_92[166], line_91[164], line_90[162], line_89[160], line_88[158], line_87[156], line_86[154], line_85[152], line_84[150], line_83[148], line_82[146], line_81[144], line_80[142], line_79[140], line_78[138], line_77[136], line_76[134], line_75[132], line_74[130], line_73[128], line_72[126], line_71[124], line_70[122], line_69[120], line_68[118], line_67[116], line_66[114], line_65[112], line_64[110], line_63[108], line_62[106], line_61[104], line_60[102], line_59[100], line_58[98], line_57[96], line_56[94], line_55[92], line_54[90], line_53[88], line_52[86], line_51[84], line_50[82], line_49[80], line_48[78], line_47[76], line_46[74], line_45[72], line_44[70], line_43[68], line_42[66], line_41[64], line_40[62], line_39[60], line_38[58], line_37[56], line_36[54], line_35[52], line_34[50], line_33[48], line_32[46], line_31[44], line_30[42], line_29[40], line_28[38], line_27[36], line_26[34], line_25[32], line_24[30], line_23[28], line_22[26], line_21[24], line_20[22], line_19[20], line_18[18], line_17[16], line_16[14], line_15[12], line_14[10], line_13[8], line_12[6], line_11[4], line_10[2], line_9[0], 8'b0};
assign col_239 = {line_128[239], line_127[237], line_126[235], line_125[233], line_124[231], line_123[229], line_122[227], line_121[225], line_120[223], line_119[221], line_118[219], line_117[217], line_116[215], line_115[213], line_114[211], line_113[209], line_112[207], line_111[205], line_110[203], line_109[201], line_108[199], line_107[197], line_106[195], line_105[193], line_104[191], line_103[189], line_102[187], line_101[185], line_100[183], line_99[181], line_98[179], line_97[177], line_96[175], line_95[173], line_94[171], line_93[169], line_92[167], line_91[165], line_90[163], line_89[161], line_88[159], line_87[157], line_86[155], line_85[153], line_84[151], line_83[149], line_82[147], line_81[145], line_80[143], line_79[141], line_78[139], line_77[137], line_76[135], line_75[133], line_74[131], line_73[129], line_72[127], line_71[125], line_70[123], line_69[121], line_68[119], line_67[117], line_66[115], line_65[113], line_64[111], line_63[109], line_62[107], line_61[105], line_60[103], line_59[101], line_58[99], line_57[97], line_56[95], line_55[93], line_54[91], line_53[89], line_52[87], line_51[85], line_50[83], line_49[81], line_48[79], line_47[77], line_46[75], line_45[73], line_44[71], line_43[69], line_42[67], line_41[65], line_40[63], line_39[61], line_38[59], line_37[57], line_36[55], line_35[53], line_34[51], line_33[49], line_32[47], line_31[45], line_30[43], line_29[41], line_28[39], line_27[37], line_26[35], line_25[33], line_24[31], line_23[29], line_22[27], line_21[25], line_20[23], line_19[21], line_18[19], line_17[17], line_16[15], line_15[13], line_14[11], line_13[9], line_12[7], line_11[5], line_10[3], line_9[1], 8'b0};
assign col_240 = {line_128[240], line_127[238], line_126[236], line_125[234], line_124[232], line_123[230], line_122[228], line_121[226], line_120[224], line_119[222], line_118[220], line_117[218], line_116[216], line_115[214], line_114[212], line_113[210], line_112[208], line_111[206], line_110[204], line_109[202], line_108[200], line_107[198], line_106[196], line_105[194], line_104[192], line_103[190], line_102[188], line_101[186], line_100[184], line_99[182], line_98[180], line_97[178], line_96[176], line_95[174], line_94[172], line_93[170], line_92[168], line_91[166], line_90[164], line_89[162], line_88[160], line_87[158], line_86[156], line_85[154], line_84[152], line_83[150], line_82[148], line_81[146], line_80[144], line_79[142], line_78[140], line_77[138], line_76[136], line_75[134], line_74[132], line_73[130], line_72[128], line_71[126], line_70[124], line_69[122], line_68[120], line_67[118], line_66[116], line_65[114], line_64[112], line_63[110], line_62[108], line_61[106], line_60[104], line_59[102], line_58[100], line_57[98], line_56[96], line_55[94], line_54[92], line_53[90], line_52[88], line_51[86], line_50[84], line_49[82], line_48[80], line_47[78], line_46[76], line_45[74], line_44[72], line_43[70], line_42[68], line_41[66], line_40[64], line_39[62], line_38[60], line_37[58], line_36[56], line_35[54], line_34[52], line_33[50], line_32[48], line_31[46], line_30[44], line_29[42], line_28[40], line_27[38], line_26[36], line_25[34], line_24[32], line_23[30], line_22[28], line_21[26], line_20[24], line_19[22], line_18[20], line_17[18], line_16[16], line_15[14], line_14[12], line_13[10], line_12[8], line_11[6], line_10[4], line_9[2], line_8[0], 7'b0};
assign col_241 = {line_128[241], line_127[239], line_126[237], line_125[235], line_124[233], line_123[231], line_122[229], line_121[227], line_120[225], line_119[223], line_118[221], line_117[219], line_116[217], line_115[215], line_114[213], line_113[211], line_112[209], line_111[207], line_110[205], line_109[203], line_108[201], line_107[199], line_106[197], line_105[195], line_104[193], line_103[191], line_102[189], line_101[187], line_100[185], line_99[183], line_98[181], line_97[179], line_96[177], line_95[175], line_94[173], line_93[171], line_92[169], line_91[167], line_90[165], line_89[163], line_88[161], line_87[159], line_86[157], line_85[155], line_84[153], line_83[151], line_82[149], line_81[147], line_80[145], line_79[143], line_78[141], line_77[139], line_76[137], line_75[135], line_74[133], line_73[131], line_72[129], line_71[127], line_70[125], line_69[123], line_68[121], line_67[119], line_66[117], line_65[115], line_64[113], line_63[111], line_62[109], line_61[107], line_60[105], line_59[103], line_58[101], line_57[99], line_56[97], line_55[95], line_54[93], line_53[91], line_52[89], line_51[87], line_50[85], line_49[83], line_48[81], line_47[79], line_46[77], line_45[75], line_44[73], line_43[71], line_42[69], line_41[67], line_40[65], line_39[63], line_38[61], line_37[59], line_36[57], line_35[55], line_34[53], line_33[51], line_32[49], line_31[47], line_30[45], line_29[43], line_28[41], line_27[39], line_26[37], line_25[35], line_24[33], line_23[31], line_22[29], line_21[27], line_20[25], line_19[23], line_18[21], line_17[19], line_16[17], line_15[15], line_14[13], line_13[11], line_12[9], line_11[7], line_10[5], line_9[3], line_8[1], 7'b0};
assign col_242 = {line_128[242], line_127[240], line_126[238], line_125[236], line_124[234], line_123[232], line_122[230], line_121[228], line_120[226], line_119[224], line_118[222], line_117[220], line_116[218], line_115[216], line_114[214], line_113[212], line_112[210], line_111[208], line_110[206], line_109[204], line_108[202], line_107[200], line_106[198], line_105[196], line_104[194], line_103[192], line_102[190], line_101[188], line_100[186], line_99[184], line_98[182], line_97[180], line_96[178], line_95[176], line_94[174], line_93[172], line_92[170], line_91[168], line_90[166], line_89[164], line_88[162], line_87[160], line_86[158], line_85[156], line_84[154], line_83[152], line_82[150], line_81[148], line_80[146], line_79[144], line_78[142], line_77[140], line_76[138], line_75[136], line_74[134], line_73[132], line_72[130], line_71[128], line_70[126], line_69[124], line_68[122], line_67[120], line_66[118], line_65[116], line_64[114], line_63[112], line_62[110], line_61[108], line_60[106], line_59[104], line_58[102], line_57[100], line_56[98], line_55[96], line_54[94], line_53[92], line_52[90], line_51[88], line_50[86], line_49[84], line_48[82], line_47[80], line_46[78], line_45[76], line_44[74], line_43[72], line_42[70], line_41[68], line_40[66], line_39[64], line_38[62], line_37[60], line_36[58], line_35[56], line_34[54], line_33[52], line_32[50], line_31[48], line_30[46], line_29[44], line_28[42], line_27[40], line_26[38], line_25[36], line_24[34], line_23[32], line_22[30], line_21[28], line_20[26], line_19[24], line_18[22], line_17[20], line_16[18], line_15[16], line_14[14], line_13[12], line_12[10], line_11[8], line_10[6], line_9[4], line_8[2], line_7[0], 6'b0};
assign col_243 = {line_128[243], line_127[241], line_126[239], line_125[237], line_124[235], line_123[233], line_122[231], line_121[229], line_120[227], line_119[225], line_118[223], line_117[221], line_116[219], line_115[217], line_114[215], line_113[213], line_112[211], line_111[209], line_110[207], line_109[205], line_108[203], line_107[201], line_106[199], line_105[197], line_104[195], line_103[193], line_102[191], line_101[189], line_100[187], line_99[185], line_98[183], line_97[181], line_96[179], line_95[177], line_94[175], line_93[173], line_92[171], line_91[169], line_90[167], line_89[165], line_88[163], line_87[161], line_86[159], line_85[157], line_84[155], line_83[153], line_82[151], line_81[149], line_80[147], line_79[145], line_78[143], line_77[141], line_76[139], line_75[137], line_74[135], line_73[133], line_72[131], line_71[129], line_70[127], line_69[125], line_68[123], line_67[121], line_66[119], line_65[117], line_64[115], line_63[113], line_62[111], line_61[109], line_60[107], line_59[105], line_58[103], line_57[101], line_56[99], line_55[97], line_54[95], line_53[93], line_52[91], line_51[89], line_50[87], line_49[85], line_48[83], line_47[81], line_46[79], line_45[77], line_44[75], line_43[73], line_42[71], line_41[69], line_40[67], line_39[65], line_38[63], line_37[61], line_36[59], line_35[57], line_34[55], line_33[53], line_32[51], line_31[49], line_30[47], line_29[45], line_28[43], line_27[41], line_26[39], line_25[37], line_24[35], line_23[33], line_22[31], line_21[29], line_20[27], line_19[25], line_18[23], line_17[21], line_16[19], line_15[17], line_14[15], line_13[13], line_12[11], line_11[9], line_10[7], line_9[5], line_8[3], line_7[1], 6'b0};
assign col_244 = {line_128[244], line_127[242], line_126[240], line_125[238], line_124[236], line_123[234], line_122[232], line_121[230], line_120[228], line_119[226], line_118[224], line_117[222], line_116[220], line_115[218], line_114[216], line_113[214], line_112[212], line_111[210], line_110[208], line_109[206], line_108[204], line_107[202], line_106[200], line_105[198], line_104[196], line_103[194], line_102[192], line_101[190], line_100[188], line_99[186], line_98[184], line_97[182], line_96[180], line_95[178], line_94[176], line_93[174], line_92[172], line_91[170], line_90[168], line_89[166], line_88[164], line_87[162], line_86[160], line_85[158], line_84[156], line_83[154], line_82[152], line_81[150], line_80[148], line_79[146], line_78[144], line_77[142], line_76[140], line_75[138], line_74[136], line_73[134], line_72[132], line_71[130], line_70[128], line_69[126], line_68[124], line_67[122], line_66[120], line_65[118], line_64[116], line_63[114], line_62[112], line_61[110], line_60[108], line_59[106], line_58[104], line_57[102], line_56[100], line_55[98], line_54[96], line_53[94], line_52[92], line_51[90], line_50[88], line_49[86], line_48[84], line_47[82], line_46[80], line_45[78], line_44[76], line_43[74], line_42[72], line_41[70], line_40[68], line_39[66], line_38[64], line_37[62], line_36[60], line_35[58], line_34[56], line_33[54], line_32[52], line_31[50], line_30[48], line_29[46], line_28[44], line_27[42], line_26[40], line_25[38], line_24[36], line_23[34], line_22[32], line_21[30], line_20[28], line_19[26], line_18[24], line_17[22], line_16[20], line_15[18], line_14[16], line_13[14], line_12[12], line_11[10], line_10[8], line_9[6], line_8[4], line_7[2], line_6[0], 5'b0};
assign col_245 = {line_128[245], line_127[243], line_126[241], line_125[239], line_124[237], line_123[235], line_122[233], line_121[231], line_120[229], line_119[227], line_118[225], line_117[223], line_116[221], line_115[219], line_114[217], line_113[215], line_112[213], line_111[211], line_110[209], line_109[207], line_108[205], line_107[203], line_106[201], line_105[199], line_104[197], line_103[195], line_102[193], line_101[191], line_100[189], line_99[187], line_98[185], line_97[183], line_96[181], line_95[179], line_94[177], line_93[175], line_92[173], line_91[171], line_90[169], line_89[167], line_88[165], line_87[163], line_86[161], line_85[159], line_84[157], line_83[155], line_82[153], line_81[151], line_80[149], line_79[147], line_78[145], line_77[143], line_76[141], line_75[139], line_74[137], line_73[135], line_72[133], line_71[131], line_70[129], line_69[127], line_68[125], line_67[123], line_66[121], line_65[119], line_64[117], line_63[115], line_62[113], line_61[111], line_60[109], line_59[107], line_58[105], line_57[103], line_56[101], line_55[99], line_54[97], line_53[95], line_52[93], line_51[91], line_50[89], line_49[87], line_48[85], line_47[83], line_46[81], line_45[79], line_44[77], line_43[75], line_42[73], line_41[71], line_40[69], line_39[67], line_38[65], line_37[63], line_36[61], line_35[59], line_34[57], line_33[55], line_32[53], line_31[51], line_30[49], line_29[47], line_28[45], line_27[43], line_26[41], line_25[39], line_24[37], line_23[35], line_22[33], line_21[31], line_20[29], line_19[27], line_18[25], line_17[23], line_16[21], line_15[19], line_14[17], line_13[15], line_12[13], line_11[11], line_10[9], line_9[7], line_8[5], line_7[3], line_6[1], 5'b0};
assign col_246 = {line_128[246], line_127[244], line_126[242], line_125[240], line_124[238], line_123[236], line_122[234], line_121[232], line_120[230], line_119[228], line_118[226], line_117[224], line_116[222], line_115[220], line_114[218], line_113[216], line_112[214], line_111[212], line_110[210], line_109[208], line_108[206], line_107[204], line_106[202], line_105[200], line_104[198], line_103[196], line_102[194], line_101[192], line_100[190], line_99[188], line_98[186], line_97[184], line_96[182], line_95[180], line_94[178], line_93[176], line_92[174], line_91[172], line_90[170], line_89[168], line_88[166], line_87[164], line_86[162], line_85[160], line_84[158], line_83[156], line_82[154], line_81[152], line_80[150], line_79[148], line_78[146], line_77[144], line_76[142], line_75[140], line_74[138], line_73[136], line_72[134], line_71[132], line_70[130], line_69[128], line_68[126], line_67[124], line_66[122], line_65[120], line_64[118], line_63[116], line_62[114], line_61[112], line_60[110], line_59[108], line_58[106], line_57[104], line_56[102], line_55[100], line_54[98], line_53[96], line_52[94], line_51[92], line_50[90], line_49[88], line_48[86], line_47[84], line_46[82], line_45[80], line_44[78], line_43[76], line_42[74], line_41[72], line_40[70], line_39[68], line_38[66], line_37[64], line_36[62], line_35[60], line_34[58], line_33[56], line_32[54], line_31[52], line_30[50], line_29[48], line_28[46], line_27[44], line_26[42], line_25[40], line_24[38], line_23[36], line_22[34], line_21[32], line_20[30], line_19[28], line_18[26], line_17[24], line_16[22], line_15[20], line_14[18], line_13[16], line_12[14], line_11[12], line_10[10], line_9[8], line_8[6], line_7[4], line_6[2], line_5[0], 4'b0};
assign col_247 = {line_128[247], line_127[245], line_126[243], line_125[241], line_124[239], line_123[237], line_122[235], line_121[233], line_120[231], line_119[229], line_118[227], line_117[225], line_116[223], line_115[221], line_114[219], line_113[217], line_112[215], line_111[213], line_110[211], line_109[209], line_108[207], line_107[205], line_106[203], line_105[201], line_104[199], line_103[197], line_102[195], line_101[193], line_100[191], line_99[189], line_98[187], line_97[185], line_96[183], line_95[181], line_94[179], line_93[177], line_92[175], line_91[173], line_90[171], line_89[169], line_88[167], line_87[165], line_86[163], line_85[161], line_84[159], line_83[157], line_82[155], line_81[153], line_80[151], line_79[149], line_78[147], line_77[145], line_76[143], line_75[141], line_74[139], line_73[137], line_72[135], line_71[133], line_70[131], line_69[129], line_68[127], line_67[125], line_66[123], line_65[121], line_64[119], line_63[117], line_62[115], line_61[113], line_60[111], line_59[109], line_58[107], line_57[105], line_56[103], line_55[101], line_54[99], line_53[97], line_52[95], line_51[93], line_50[91], line_49[89], line_48[87], line_47[85], line_46[83], line_45[81], line_44[79], line_43[77], line_42[75], line_41[73], line_40[71], line_39[69], line_38[67], line_37[65], line_36[63], line_35[61], line_34[59], line_33[57], line_32[55], line_31[53], line_30[51], line_29[49], line_28[47], line_27[45], line_26[43], line_25[41], line_24[39], line_23[37], line_22[35], line_21[33], line_20[31], line_19[29], line_18[27], line_17[25], line_16[23], line_15[21], line_14[19], line_13[17], line_12[15], line_11[13], line_10[11], line_9[9], line_8[7], line_7[5], line_6[3], line_5[1], 4'b0};
assign col_248 = {line_128[248], line_127[246], line_126[244], line_125[242], line_124[240], line_123[238], line_122[236], line_121[234], line_120[232], line_119[230], line_118[228], line_117[226], line_116[224], line_115[222], line_114[220], line_113[218], line_112[216], line_111[214], line_110[212], line_109[210], line_108[208], line_107[206], line_106[204], line_105[202], line_104[200], line_103[198], line_102[196], line_101[194], line_100[192], line_99[190], line_98[188], line_97[186], line_96[184], line_95[182], line_94[180], line_93[178], line_92[176], line_91[174], line_90[172], line_89[170], line_88[168], line_87[166], line_86[164], line_85[162], line_84[160], line_83[158], line_82[156], line_81[154], line_80[152], line_79[150], line_78[148], line_77[146], line_76[144], line_75[142], line_74[140], line_73[138], line_72[136], line_71[134], line_70[132], line_69[130], line_68[128], line_67[126], line_66[124], line_65[122], line_64[120], line_63[118], line_62[116], line_61[114], line_60[112], line_59[110], line_58[108], line_57[106], line_56[104], line_55[102], line_54[100], line_53[98], line_52[96], line_51[94], line_50[92], line_49[90], line_48[88], line_47[86], line_46[84], line_45[82], line_44[80], line_43[78], line_42[76], line_41[74], line_40[72], line_39[70], line_38[68], line_37[66], line_36[64], line_35[62], line_34[60], line_33[58], line_32[56], line_31[54], line_30[52], line_29[50], line_28[48], line_27[46], line_26[44], line_25[42], line_24[40], line_23[38], line_22[36], line_21[34], line_20[32], line_19[30], line_18[28], line_17[26], line_16[24], line_15[22], line_14[20], line_13[18], line_12[16], line_11[14], line_10[12], line_9[10], line_8[8], line_7[6], line_6[4], line_5[2], line_4[0], 3'b0};
assign col_249 = {line_128[249], line_127[247], line_126[245], line_125[243], line_124[241], line_123[239], line_122[237], line_121[235], line_120[233], line_119[231], line_118[229], line_117[227], line_116[225], line_115[223], line_114[221], line_113[219], line_112[217], line_111[215], line_110[213], line_109[211], line_108[209], line_107[207], line_106[205], line_105[203], line_104[201], line_103[199], line_102[197], line_101[195], line_100[193], line_99[191], line_98[189], line_97[187], line_96[185], line_95[183], line_94[181], line_93[179], line_92[177], line_91[175], line_90[173], line_89[171], line_88[169], line_87[167], line_86[165], line_85[163], line_84[161], line_83[159], line_82[157], line_81[155], line_80[153], line_79[151], line_78[149], line_77[147], line_76[145], line_75[143], line_74[141], line_73[139], line_72[137], line_71[135], line_70[133], line_69[131], line_68[129], line_67[127], line_66[125], line_65[123], line_64[121], line_63[119], line_62[117], line_61[115], line_60[113], line_59[111], line_58[109], line_57[107], line_56[105], line_55[103], line_54[101], line_53[99], line_52[97], line_51[95], line_50[93], line_49[91], line_48[89], line_47[87], line_46[85], line_45[83], line_44[81], line_43[79], line_42[77], line_41[75], line_40[73], line_39[71], line_38[69], line_37[67], line_36[65], line_35[63], line_34[61], line_33[59], line_32[57], line_31[55], line_30[53], line_29[51], line_28[49], line_27[47], line_26[45], line_25[43], line_24[41], line_23[39], line_22[37], line_21[35], line_20[33], line_19[31], line_18[29], line_17[27], line_16[25], line_15[23], line_14[21], line_13[19], line_12[17], line_11[15], line_10[13], line_9[11], line_8[9], line_7[7], line_6[5], line_5[3], line_4[1], 3'b0};
assign col_250 = {line_128[250], line_127[248], line_126[246], line_125[244], line_124[242], line_123[240], line_122[238], line_121[236], line_120[234], line_119[232], line_118[230], line_117[228], line_116[226], line_115[224], line_114[222], line_113[220], line_112[218], line_111[216], line_110[214], line_109[212], line_108[210], line_107[208], line_106[206], line_105[204], line_104[202], line_103[200], line_102[198], line_101[196], line_100[194], line_99[192], line_98[190], line_97[188], line_96[186], line_95[184], line_94[182], line_93[180], line_92[178], line_91[176], line_90[174], line_89[172], line_88[170], line_87[168], line_86[166], line_85[164], line_84[162], line_83[160], line_82[158], line_81[156], line_80[154], line_79[152], line_78[150], line_77[148], line_76[146], line_75[144], line_74[142], line_73[140], line_72[138], line_71[136], line_70[134], line_69[132], line_68[130], line_67[128], line_66[126], line_65[124], line_64[122], line_63[120], line_62[118], line_61[116], line_60[114], line_59[112], line_58[110], line_57[108], line_56[106], line_55[104], line_54[102], line_53[100], line_52[98], line_51[96], line_50[94], line_49[92], line_48[90], line_47[88], line_46[86], line_45[84], line_44[82], line_43[80], line_42[78], line_41[76], line_40[74], line_39[72], line_38[70], line_37[68], line_36[66], line_35[64], line_34[62], line_33[60], line_32[58], line_31[56], line_30[54], line_29[52], line_28[50], line_27[48], line_26[46], line_25[44], line_24[42], line_23[40], line_22[38], line_21[36], line_20[34], line_19[32], line_18[30], line_17[28], line_16[26], line_15[24], line_14[22], line_13[20], line_12[18], line_11[16], line_10[14], line_9[12], line_8[10], line_7[8], line_6[6], line_5[4], line_4[2], line_3[0], 2'b0};
assign col_251 = {line_128[251], line_127[249], line_126[247], line_125[245], line_124[243], line_123[241], line_122[239], line_121[237], line_120[235], line_119[233], line_118[231], line_117[229], line_116[227], line_115[225], line_114[223], line_113[221], line_112[219], line_111[217], line_110[215], line_109[213], line_108[211], line_107[209], line_106[207], line_105[205], line_104[203], line_103[201], line_102[199], line_101[197], line_100[195], line_99[193], line_98[191], line_97[189], line_96[187], line_95[185], line_94[183], line_93[181], line_92[179], line_91[177], line_90[175], line_89[173], line_88[171], line_87[169], line_86[167], line_85[165], line_84[163], line_83[161], line_82[159], line_81[157], line_80[155], line_79[153], line_78[151], line_77[149], line_76[147], line_75[145], line_74[143], line_73[141], line_72[139], line_71[137], line_70[135], line_69[133], line_68[131], line_67[129], line_66[127], line_65[125], line_64[123], line_63[121], line_62[119], line_61[117], line_60[115], line_59[113], line_58[111], line_57[109], line_56[107], line_55[105], line_54[103], line_53[101], line_52[99], line_51[97], line_50[95], line_49[93], line_48[91], line_47[89], line_46[87], line_45[85], line_44[83], line_43[81], line_42[79], line_41[77], line_40[75], line_39[73], line_38[71], line_37[69], line_36[67], line_35[65], line_34[63], line_33[61], line_32[59], line_31[57], line_30[55], line_29[53], line_28[51], line_27[49], line_26[47], line_25[45], line_24[43], line_23[41], line_22[39], line_21[37], line_20[35], line_19[33], line_18[31], line_17[29], line_16[27], line_15[25], line_14[23], line_13[21], line_12[19], line_11[17], line_10[15], line_9[13], line_8[11], line_7[9], line_6[7], line_5[5], line_4[3], line_3[1], 2'b0};
assign col_252 = {line_128[252], line_127[250], line_126[248], line_125[246], line_124[244], line_123[242], line_122[240], line_121[238], line_120[236], line_119[234], line_118[232], line_117[230], line_116[228], line_115[226], line_114[224], line_113[222], line_112[220], line_111[218], line_110[216], line_109[214], line_108[212], line_107[210], line_106[208], line_105[206], line_104[204], line_103[202], line_102[200], line_101[198], line_100[196], line_99[194], line_98[192], line_97[190], line_96[188], line_95[186], line_94[184], line_93[182], line_92[180], line_91[178], line_90[176], line_89[174], line_88[172], line_87[170], line_86[168], line_85[166], line_84[164], line_83[162], line_82[160], line_81[158], line_80[156], line_79[154], line_78[152], line_77[150], line_76[148], line_75[146], line_74[144], line_73[142], line_72[140], line_71[138], line_70[136], line_69[134], line_68[132], line_67[130], line_66[128], line_65[126], line_64[124], line_63[122], line_62[120], line_61[118], line_60[116], line_59[114], line_58[112], line_57[110], line_56[108], line_55[106], line_54[104], line_53[102], line_52[100], line_51[98], line_50[96], line_49[94], line_48[92], line_47[90], line_46[88], line_45[86], line_44[84], line_43[82], line_42[80], line_41[78], line_40[76], line_39[74], line_38[72], line_37[70], line_36[68], line_35[66], line_34[64], line_33[62], line_32[60], line_31[58], line_30[56], line_29[54], line_28[52], line_27[50], line_26[48], line_25[46], line_24[44], line_23[42], line_22[40], line_21[38], line_20[36], line_19[34], line_18[32], line_17[30], line_16[28], line_15[26], line_14[24], line_13[22], line_12[20], line_11[18], line_10[16], line_9[14], line_8[12], line_7[10], line_6[8], line_5[6], line_4[4], line_3[2], line_2[0], 1'b0};
assign col_253 = {line_128[253], line_127[251], line_126[249], line_125[247], line_124[245], line_123[243], line_122[241], line_121[239], line_120[237], line_119[235], line_118[233], line_117[231], line_116[229], line_115[227], line_114[225], line_113[223], line_112[221], line_111[219], line_110[217], line_109[215], line_108[213], line_107[211], line_106[209], line_105[207], line_104[205], line_103[203], line_102[201], line_101[199], line_100[197], line_99[195], line_98[193], line_97[191], line_96[189], line_95[187], line_94[185], line_93[183], line_92[181], line_91[179], line_90[177], line_89[175], line_88[173], line_87[171], line_86[169], line_85[167], line_84[165], line_83[163], line_82[161], line_81[159], line_80[157], line_79[155], line_78[153], line_77[151], line_76[149], line_75[147], line_74[145], line_73[143], line_72[141], line_71[139], line_70[137], line_69[135], line_68[133], line_67[131], line_66[129], line_65[127], line_64[125], line_63[123], line_62[121], line_61[119], line_60[117], line_59[115], line_58[113], line_57[111], line_56[109], line_55[107], line_54[105], line_53[103], line_52[101], line_51[99], line_50[97], line_49[95], line_48[93], line_47[91], line_46[89], line_45[87], line_44[85], line_43[83], line_42[81], line_41[79], line_40[77], line_39[75], line_38[73], line_37[71], line_36[69], line_35[67], line_34[65], line_33[63], line_32[61], line_31[59], line_30[57], line_29[55], line_28[53], line_27[51], line_26[49], line_25[47], line_24[45], line_23[43], line_22[41], line_21[39], line_20[37], line_19[35], line_18[33], line_17[31], line_16[29], line_15[27], line_14[25], line_13[23], line_12[21], line_11[19], line_10[17], line_9[15], line_8[13], line_7[11], line_6[9], line_5[7], line_4[5], line_3[3], line_2[1], 1'b0};
assign col_254 = {line_128[254], line_127[252], line_126[250], line_125[248], line_124[246], line_123[244], line_122[242], line_121[240], line_120[238], line_119[236], line_118[234], line_117[232], line_116[230], line_115[228], line_114[226], line_113[224], line_112[222], line_111[220], line_110[218], line_109[216], line_108[214], line_107[212], line_106[210], line_105[208], line_104[206], line_103[204], line_102[202], line_101[200], line_100[198], line_99[196], line_98[194], line_97[192], line_96[190], line_95[188], line_94[186], line_93[184], line_92[182], line_91[180], line_90[178], line_89[176], line_88[174], line_87[172], line_86[170], line_85[168], line_84[166], line_83[164], line_82[162], line_81[160], line_80[158], line_79[156], line_78[154], line_77[152], line_76[150], line_75[148], line_74[146], line_73[144], line_72[142], line_71[140], line_70[138], line_69[136], line_68[134], line_67[132], line_66[130], line_65[128], line_64[126], line_63[124], line_62[122], line_61[120], line_60[118], line_59[116], line_58[114], line_57[112], line_56[110], line_55[108], line_54[106], line_53[104], line_52[102], line_51[100], line_50[98], line_49[96], line_48[94], line_47[92], line_46[90], line_45[88], line_44[86], line_43[84], line_42[82], line_41[80], line_40[78], line_39[76], line_38[74], line_37[72], line_36[70], line_35[68], line_34[66], line_33[64], line_32[62], line_31[60], line_30[58], line_29[56], line_28[54], line_27[52], line_26[50], line_25[48], line_24[46], line_23[44], line_22[42], line_21[40], line_20[38], line_19[36], line_18[34], line_17[32], line_16[30], line_15[28], line_14[26], line_13[24], line_12[22], line_11[20], line_10[18], line_9[16], line_8[14], line_7[12], line_6[10], line_5[8], line_4[6], line_3[4], line_2[2], line_1[0]};
assign col_255 = {line_128[255], line_127[253], line_126[251], line_125[249], line_124[247], line_123[245], line_122[243], line_121[241], line_120[239], line_119[237], line_118[235], line_117[233], line_116[231], line_115[229], line_114[227], line_113[225], line_112[223], line_111[221], line_110[219], line_109[217], line_108[215], line_107[213], line_106[211], line_105[209], line_104[207], line_103[205], line_102[203], line_101[201], line_100[199], line_99[197], line_98[195], line_97[193], line_96[191], line_95[189], line_94[187], line_93[185], line_92[183], line_91[181], line_90[179], line_89[177], line_88[175], line_87[173], line_86[171], line_85[169], line_84[167], line_83[165], line_82[163], line_81[161], line_80[159], line_79[157], line_78[155], line_77[153], line_76[151], line_75[149], line_74[147], line_73[145], line_72[143], line_71[141], line_70[139], line_69[137], line_68[135], line_67[133], line_66[131], line_65[129], line_64[127], line_63[125], line_62[123], line_61[121], line_60[119], line_59[117], line_58[115], line_57[113], line_56[111], line_55[109], line_54[107], line_53[105], line_52[103], line_51[101], line_50[99], line_49[97], line_48[95], line_47[93], line_46[91], line_45[89], line_44[87], line_43[85], line_42[83], line_41[81], line_40[79], line_39[77], line_38[75], line_37[73], line_36[71], line_35[69], line_34[67], line_33[65], line_32[63], line_31[61], line_30[59], line_29[57], line_28[55], line_27[53], line_26[51], line_25[49], line_24[47], line_23[45], line_22[43], line_21[41], line_20[39], line_19[37], line_18[35], line_17[33], line_16[31], line_15[29], line_14[27], line_13[25], line_12[23], line_11[21], line_10[19], line_9[17], line_8[15], line_7[13], line_6[11], line_5[9], line_4[7], line_3[5], line_2[3], line_1[1]};

assign col_256 = {line_128[256], line_127[254], line_126[252], line_125[250], line_124[248], line_123[246], line_122[244], line_121[242], line_120[240], line_119[238], line_118[236], line_117[234], line_116[232], line_115[230], line_114[228], line_113[226], line_112[224], line_111[222], line_110[220], line_109[218], line_108[216], line_107[214], line_106[212], line_105[210], line_104[208], line_103[206], line_102[204], line_101[202], line_100[200], line_99[198], line_98[196], line_97[194], line_96[192], line_95[190], line_94[188], line_93[186], line_92[184], line_91[182], line_90[180], line_89[178], line_88[176], line_87[174], line_86[172], line_85[170], line_84[168], line_83[166], line_82[164], line_81[162], line_80[160], line_79[158], line_78[156], line_77[154], line_76[152], line_75[150], line_74[148], line_73[146], line_72[144], line_71[142], line_70[140], line_69[138], line_68[136], line_67[134], line_66[132], line_65[130], line_64[128], line_63[126], line_62[124], line_61[122], line_60[120], line_59[118], line_58[116], line_57[114], line_56[112], line_55[110], line_54[108], line_53[106], line_52[104], line_51[102], line_50[100], line_49[98], line_48[96], line_47[94], line_46[92], line_45[90], line_44[88], line_43[86], line_42[84], line_41[82], line_40[80], line_39[78], line_38[76], line_37[74], line_36[72], line_35[70], line_34[68], line_33[66], line_32[64], line_31[62], line_30[60], line_29[58], line_28[56], line_27[54], line_26[52], line_25[50], line_24[48], line_23[46], line_22[44], line_21[42], line_20[40], line_19[38], line_18[36], line_17[34], line_16[32], line_15[30], line_14[28], line_13[26], line_12[24], line_11[22], line_10[20], line_9[18], line_8[16], line_7[14], line_6[12], line_5[10], line_4[8], line_3[6], line_2[4], line_1[2] };
assign col_257 = {line_128[257], line_127[255], line_126[253], line_125[251], line_124[249], line_123[247], line_122[245], line_121[243], line_120[241], line_119[239], line_118[237], line_117[235], line_116[233], line_115[231], line_114[229], line_113[227], line_112[225], line_111[223], line_110[221], line_109[219], line_108[217], line_107[215], line_106[213], line_105[211], line_104[209], line_103[207], line_102[205], line_101[203], line_100[201], line_99[199], line_98[197], line_97[195], line_96[193], line_95[191], line_94[189], line_93[187], line_92[185], line_91[183], line_90[181], line_89[179], line_88[177], line_87[175], line_86[173], line_85[171], line_84[169], line_83[167], line_82[165], line_81[163], line_80[161], line_79[159], line_78[157], line_77[155], line_76[153], line_75[151], line_74[149], line_73[147], line_72[145], line_71[143], line_70[141], line_69[139], line_68[137], line_67[135], line_66[133], line_65[131], line_64[129], line_63[127], line_62[125], line_61[123], line_60[121], line_59[119], line_58[117], line_57[115], line_56[113], line_55[111], line_54[109], line_53[107], line_52[105], line_51[103], line_50[101], line_49[99], line_48[97], line_47[95], line_46[93], line_45[91], line_44[89], line_43[87], line_42[85], line_41[83], line_40[81], line_39[79], line_38[77], line_37[75], line_36[73], line_35[71], line_34[69], line_33[67], line_32[65], line_31[63], line_30[61], line_29[59], line_28[57], line_27[55], line_26[53], line_25[51], line_24[49], line_23[47], line_22[45], line_21[43], line_20[41], line_19[39], line_18[37], line_17[35], line_16[33], line_15[31], line_14[29], line_13[27], line_12[25], line_11[23], line_10[21], line_9[19], line_8[17], line_7[15], line_6[13], line_5[11], line_4[9], line_3[7], line_2[5], line_1[3] };
assign col_258 = {line_128[258], line_127[256], line_126[254], line_125[252], line_124[250], line_123[248], line_122[246], line_121[244], line_120[242], line_119[240], line_118[238], line_117[236], line_116[234], line_115[232], line_114[230], line_113[228], line_112[226], line_111[224], line_110[222], line_109[220], line_108[218], line_107[216], line_106[214], line_105[212], line_104[210], line_103[208], line_102[206], line_101[204], line_100[202], line_99[200], line_98[198], line_97[196], line_96[194], line_95[192], line_94[190], line_93[188], line_92[186], line_91[184], line_90[182], line_89[180], line_88[178], line_87[176], line_86[174], line_85[172], line_84[170], line_83[168], line_82[166], line_81[164], line_80[162], line_79[160], line_78[158], line_77[156], line_76[154], line_75[152], line_74[150], line_73[148], line_72[146], line_71[144], line_70[142], line_69[140], line_68[138], line_67[136], line_66[134], line_65[132], line_64[130], line_63[128], line_62[126], line_61[124], line_60[122], line_59[120], line_58[118], line_57[116], line_56[114], line_55[112], line_54[110], line_53[108], line_52[106], line_51[104], line_50[102], line_49[100], line_48[98], line_47[96], line_46[94], line_45[92], line_44[90], line_43[88], line_42[86], line_41[84], line_40[82], line_39[80], line_38[78], line_37[76], line_36[74], line_35[72], line_34[70], line_33[68], line_32[66], line_31[64], line_30[62], line_29[60], line_28[58], line_27[56], line_26[54], line_25[52], line_24[50], line_23[48], line_22[46], line_21[44], line_20[42], line_19[40], line_18[38], line_17[36], line_16[34], line_15[32], line_14[30], line_13[28], line_12[26], line_11[24], line_10[22], line_9[20], line_8[18], line_7[16], line_6[14], line_5[12], line_4[10], line_3[8], line_2[6], line_1[4] };
assign col_259 = {line_128[259], line_127[257], line_126[255], line_125[253], line_124[251], line_123[249], line_122[247], line_121[245], line_120[243], line_119[241], line_118[239], line_117[237], line_116[235], line_115[233], line_114[231], line_113[229], line_112[227], line_111[225], line_110[223], line_109[221], line_108[219], line_107[217], line_106[215], line_105[213], line_104[211], line_103[209], line_102[207], line_101[205], line_100[203], line_99[201], line_98[199], line_97[197], line_96[195], line_95[193], line_94[191], line_93[189], line_92[187], line_91[185], line_90[183], line_89[181], line_88[179], line_87[177], line_86[175], line_85[173], line_84[171], line_83[169], line_82[167], line_81[165], line_80[163], line_79[161], line_78[159], line_77[157], line_76[155], line_75[153], line_74[151], line_73[149], line_72[147], line_71[145], line_70[143], line_69[141], line_68[139], line_67[137], line_66[135], line_65[133], line_64[131], line_63[129], line_62[127], line_61[125], line_60[123], line_59[121], line_58[119], line_57[117], line_56[115], line_55[113], line_54[111], line_53[109], line_52[107], line_51[105], line_50[103], line_49[101], line_48[99], line_47[97], line_46[95], line_45[93], line_44[91], line_43[89], line_42[87], line_41[85], line_40[83], line_39[81], line_38[79], line_37[77], line_36[75], line_35[73], line_34[71], line_33[69], line_32[67], line_31[65], line_30[63], line_29[61], line_28[59], line_27[57], line_26[55], line_25[53], line_24[51], line_23[49], line_22[47], line_21[45], line_20[43], line_19[41], line_18[39], line_17[37], line_16[35], line_15[33], line_14[31], line_13[29], line_12[27], line_11[25], line_10[23], line_9[21], line_8[19], line_7[17], line_6[15], line_5[13], line_4[11], line_3[9], line_2[7], line_1[5] };
assign col_260 = {line_128[260], line_127[258], line_126[256], line_125[254], line_124[252], line_123[250], line_122[248], line_121[246], line_120[244], line_119[242], line_118[240], line_117[238], line_116[236], line_115[234], line_114[232], line_113[230], line_112[228], line_111[226], line_110[224], line_109[222], line_108[220], line_107[218], line_106[216], line_105[214], line_104[212], line_103[210], line_102[208], line_101[206], line_100[204], line_99[202], line_98[200], line_97[198], line_96[196], line_95[194], line_94[192], line_93[190], line_92[188], line_91[186], line_90[184], line_89[182], line_88[180], line_87[178], line_86[176], line_85[174], line_84[172], line_83[170], line_82[168], line_81[166], line_80[164], line_79[162], line_78[160], line_77[158], line_76[156], line_75[154], line_74[152], line_73[150], line_72[148], line_71[146], line_70[144], line_69[142], line_68[140], line_67[138], line_66[136], line_65[134], line_64[132], line_63[130], line_62[128], line_61[126], line_60[124], line_59[122], line_58[120], line_57[118], line_56[116], line_55[114], line_54[112], line_53[110], line_52[108], line_51[106], line_50[104], line_49[102], line_48[100], line_47[98], line_46[96], line_45[94], line_44[92], line_43[90], line_42[88], line_41[86], line_40[84], line_39[82], line_38[80], line_37[78], line_36[76], line_35[74], line_34[72], line_33[70], line_32[68], line_31[66], line_30[64], line_29[62], line_28[60], line_27[58], line_26[56], line_25[54], line_24[52], line_23[50], line_22[48], line_21[46], line_20[44], line_19[42], line_18[40], line_17[38], line_16[36], line_15[34], line_14[32], line_13[30], line_12[28], line_11[26], line_10[24], line_9[22], line_8[20], line_7[18], line_6[16], line_5[14], line_4[12], line_3[10], line_2[8], line_1[6] };
assign col_261 = {line_128[261], line_127[259], line_126[257], line_125[255], line_124[253], line_123[251], line_122[249], line_121[247], line_120[245], line_119[243], line_118[241], line_117[239], line_116[237], line_115[235], line_114[233], line_113[231], line_112[229], line_111[227], line_110[225], line_109[223], line_108[221], line_107[219], line_106[217], line_105[215], line_104[213], line_103[211], line_102[209], line_101[207], line_100[205], line_99[203], line_98[201], line_97[199], line_96[197], line_95[195], line_94[193], line_93[191], line_92[189], line_91[187], line_90[185], line_89[183], line_88[181], line_87[179], line_86[177], line_85[175], line_84[173], line_83[171], line_82[169], line_81[167], line_80[165], line_79[163], line_78[161], line_77[159], line_76[157], line_75[155], line_74[153], line_73[151], line_72[149], line_71[147], line_70[145], line_69[143], line_68[141], line_67[139], line_66[137], line_65[135], line_64[133], line_63[131], line_62[129], line_61[127], line_60[125], line_59[123], line_58[121], line_57[119], line_56[117], line_55[115], line_54[113], line_53[111], line_52[109], line_51[107], line_50[105], line_49[103], line_48[101], line_47[99], line_46[97], line_45[95], line_44[93], line_43[91], line_42[89], line_41[87], line_40[85], line_39[83], line_38[81], line_37[79], line_36[77], line_35[75], line_34[73], line_33[71], line_32[69], line_31[67], line_30[65], line_29[63], line_28[61], line_27[59], line_26[57], line_25[55], line_24[53], line_23[51], line_22[49], line_21[47], line_20[45], line_19[43], line_18[41], line_17[39], line_16[37], line_15[35], line_14[33], line_13[31], line_12[29], line_11[27], line_10[25], line_9[23], line_8[21], line_7[19], line_6[17], line_5[15], line_4[13], line_3[11], line_2[9], line_1[7] };
assign col_262 = {line_128[262], line_127[260], line_126[258], line_125[256], line_124[254], line_123[252], line_122[250], line_121[248], line_120[246], line_119[244], line_118[242], line_117[240], line_116[238], line_115[236], line_114[234], line_113[232], line_112[230], line_111[228], line_110[226], line_109[224], line_108[222], line_107[220], line_106[218], line_105[216], line_104[214], line_103[212], line_102[210], line_101[208], line_100[206], line_99[204], line_98[202], line_97[200], line_96[198], line_95[196], line_94[194], line_93[192], line_92[190], line_91[188], line_90[186], line_89[184], line_88[182], line_87[180], line_86[178], line_85[176], line_84[174], line_83[172], line_82[170], line_81[168], line_80[166], line_79[164], line_78[162], line_77[160], line_76[158], line_75[156], line_74[154], line_73[152], line_72[150], line_71[148], line_70[146], line_69[144], line_68[142], line_67[140], line_66[138], line_65[136], line_64[134], line_63[132], line_62[130], line_61[128], line_60[126], line_59[124], line_58[122], line_57[120], line_56[118], line_55[116], line_54[114], line_53[112], line_52[110], line_51[108], line_50[106], line_49[104], line_48[102], line_47[100], line_46[98], line_45[96], line_44[94], line_43[92], line_42[90], line_41[88], line_40[86], line_39[84], line_38[82], line_37[80], line_36[78], line_35[76], line_34[74], line_33[72], line_32[70], line_31[68], line_30[66], line_29[64], line_28[62], line_27[60], line_26[58], line_25[56], line_24[54], line_23[52], line_22[50], line_21[48], line_20[46], line_19[44], line_18[42], line_17[40], line_16[38], line_15[36], line_14[34], line_13[32], line_12[30], line_11[28], line_10[26], line_9[24], line_8[22], line_7[20], line_6[18], line_5[16], line_4[14], line_3[12], line_2[10], line_1[8] };
assign col_263 = {line_128[263], line_127[261], line_126[259], line_125[257], line_124[255], line_123[253], line_122[251], line_121[249], line_120[247], line_119[245], line_118[243], line_117[241], line_116[239], line_115[237], line_114[235], line_113[233], line_112[231], line_111[229], line_110[227], line_109[225], line_108[223], line_107[221], line_106[219], line_105[217], line_104[215], line_103[213], line_102[211], line_101[209], line_100[207], line_99[205], line_98[203], line_97[201], line_96[199], line_95[197], line_94[195], line_93[193], line_92[191], line_91[189], line_90[187], line_89[185], line_88[183], line_87[181], line_86[179], line_85[177], line_84[175], line_83[173], line_82[171], line_81[169], line_80[167], line_79[165], line_78[163], line_77[161], line_76[159], line_75[157], line_74[155], line_73[153], line_72[151], line_71[149], line_70[147], line_69[145], line_68[143], line_67[141], line_66[139], line_65[137], line_64[135], line_63[133], line_62[131], line_61[129], line_60[127], line_59[125], line_58[123], line_57[121], line_56[119], line_55[117], line_54[115], line_53[113], line_52[111], line_51[109], line_50[107], line_49[105], line_48[103], line_47[101], line_46[99], line_45[97], line_44[95], line_43[93], line_42[91], line_41[89], line_40[87], line_39[85], line_38[83], line_37[81], line_36[79], line_35[77], line_34[75], line_33[73], line_32[71], line_31[69], line_30[67], line_29[65], line_28[63], line_27[61], line_26[59], line_25[57], line_24[55], line_23[53], line_22[51], line_21[49], line_20[47], line_19[45], line_18[43], line_17[41], line_16[39], line_15[37], line_14[35], line_13[33], line_12[31], line_11[29], line_10[27], line_9[25], line_8[23], line_7[21], line_6[19], line_5[17], line_4[15], line_3[13], line_2[11], line_1[9] };
assign col_264 = {line_128[264], line_127[262], line_126[260], line_125[258], line_124[256], line_123[254], line_122[252], line_121[250], line_120[248], line_119[246], line_118[244], line_117[242], line_116[240], line_115[238], line_114[236], line_113[234], line_112[232], line_111[230], line_110[228], line_109[226], line_108[224], line_107[222], line_106[220], line_105[218], line_104[216], line_103[214], line_102[212], line_101[210], line_100[208], line_99[206], line_98[204], line_97[202], line_96[200], line_95[198], line_94[196], line_93[194], line_92[192], line_91[190], line_90[188], line_89[186], line_88[184], line_87[182], line_86[180], line_85[178], line_84[176], line_83[174], line_82[172], line_81[170], line_80[168], line_79[166], line_78[164], line_77[162], line_76[160], line_75[158], line_74[156], line_73[154], line_72[152], line_71[150], line_70[148], line_69[146], line_68[144], line_67[142], line_66[140], line_65[138], line_64[136], line_63[134], line_62[132], line_61[130], line_60[128], line_59[126], line_58[124], line_57[122], line_56[120], line_55[118], line_54[116], line_53[114], line_52[112], line_51[110], line_50[108], line_49[106], line_48[104], line_47[102], line_46[100], line_45[98], line_44[96], line_43[94], line_42[92], line_41[90], line_40[88], line_39[86], line_38[84], line_37[82], line_36[80], line_35[78], line_34[76], line_33[74], line_32[72], line_31[70], line_30[68], line_29[66], line_28[64], line_27[62], line_26[60], line_25[58], line_24[56], line_23[54], line_22[52], line_21[50], line_20[48], line_19[46], line_18[44], line_17[42], line_16[40], line_15[38], line_14[36], line_13[34], line_12[32], line_11[30], line_10[28], line_9[26], line_8[24], line_7[22], line_6[20], line_5[18], line_4[16], line_3[14], line_2[12], line_1[10] };
assign col_265 = {line_128[265], line_127[263], line_126[261], line_125[259], line_124[257], line_123[255], line_122[253], line_121[251], line_120[249], line_119[247], line_118[245], line_117[243], line_116[241], line_115[239], line_114[237], line_113[235], line_112[233], line_111[231], line_110[229], line_109[227], line_108[225], line_107[223], line_106[221], line_105[219], line_104[217], line_103[215], line_102[213], line_101[211], line_100[209], line_99[207], line_98[205], line_97[203], line_96[201], line_95[199], line_94[197], line_93[195], line_92[193], line_91[191], line_90[189], line_89[187], line_88[185], line_87[183], line_86[181], line_85[179], line_84[177], line_83[175], line_82[173], line_81[171], line_80[169], line_79[167], line_78[165], line_77[163], line_76[161], line_75[159], line_74[157], line_73[155], line_72[153], line_71[151], line_70[149], line_69[147], line_68[145], line_67[143], line_66[141], line_65[139], line_64[137], line_63[135], line_62[133], line_61[131], line_60[129], line_59[127], line_58[125], line_57[123], line_56[121], line_55[119], line_54[117], line_53[115], line_52[113], line_51[111], line_50[109], line_49[107], line_48[105], line_47[103], line_46[101], line_45[99], line_44[97], line_43[95], line_42[93], line_41[91], line_40[89], line_39[87], line_38[85], line_37[83], line_36[81], line_35[79], line_34[77], line_33[75], line_32[73], line_31[71], line_30[69], line_29[67], line_28[65], line_27[63], line_26[61], line_25[59], line_24[57], line_23[55], line_22[53], line_21[51], line_20[49], line_19[47], line_18[45], line_17[43], line_16[41], line_15[39], line_14[37], line_13[35], line_12[33], line_11[31], line_10[29], line_9[27], line_8[25], line_7[23], line_6[21], line_5[19], line_4[17], line_3[15], line_2[13], line_1[11] };
assign col_266 = {line_128[266], line_127[264], line_126[262], line_125[260], line_124[258], line_123[256], line_122[254], line_121[252], line_120[250], line_119[248], line_118[246], line_117[244], line_116[242], line_115[240], line_114[238], line_113[236], line_112[234], line_111[232], line_110[230], line_109[228], line_108[226], line_107[224], line_106[222], line_105[220], line_104[218], line_103[216], line_102[214], line_101[212], line_100[210], line_99[208], line_98[206], line_97[204], line_96[202], line_95[200], line_94[198], line_93[196], line_92[194], line_91[192], line_90[190], line_89[188], line_88[186], line_87[184], line_86[182], line_85[180], line_84[178], line_83[176], line_82[174], line_81[172], line_80[170], line_79[168], line_78[166], line_77[164], line_76[162], line_75[160], line_74[158], line_73[156], line_72[154], line_71[152], line_70[150], line_69[148], line_68[146], line_67[144], line_66[142], line_65[140], line_64[138], line_63[136], line_62[134], line_61[132], line_60[130], line_59[128], line_58[126], line_57[124], line_56[122], line_55[120], line_54[118], line_53[116], line_52[114], line_51[112], line_50[110], line_49[108], line_48[106], line_47[104], line_46[102], line_45[100], line_44[98], line_43[96], line_42[94], line_41[92], line_40[90], line_39[88], line_38[86], line_37[84], line_36[82], line_35[80], line_34[78], line_33[76], line_32[74], line_31[72], line_30[70], line_29[68], line_28[66], line_27[64], line_26[62], line_25[60], line_24[58], line_23[56], line_22[54], line_21[52], line_20[50], line_19[48], line_18[46], line_17[44], line_16[42], line_15[40], line_14[38], line_13[36], line_12[34], line_11[32], line_10[30], line_9[28], line_8[26], line_7[24], line_6[22], line_5[20], line_4[18], line_3[16], line_2[14], line_1[12] };
assign col_267 = {line_128[267], line_127[265], line_126[263], line_125[261], line_124[259], line_123[257], line_122[255], line_121[253], line_120[251], line_119[249], line_118[247], line_117[245], line_116[243], line_115[241], line_114[239], line_113[237], line_112[235], line_111[233], line_110[231], line_109[229], line_108[227], line_107[225], line_106[223], line_105[221], line_104[219], line_103[217], line_102[215], line_101[213], line_100[211], line_99[209], line_98[207], line_97[205], line_96[203], line_95[201], line_94[199], line_93[197], line_92[195], line_91[193], line_90[191], line_89[189], line_88[187], line_87[185], line_86[183], line_85[181], line_84[179], line_83[177], line_82[175], line_81[173], line_80[171], line_79[169], line_78[167], line_77[165], line_76[163], line_75[161], line_74[159], line_73[157], line_72[155], line_71[153], line_70[151], line_69[149], line_68[147], line_67[145], line_66[143], line_65[141], line_64[139], line_63[137], line_62[135], line_61[133], line_60[131], line_59[129], line_58[127], line_57[125], line_56[123], line_55[121], line_54[119], line_53[117], line_52[115], line_51[113], line_50[111], line_49[109], line_48[107], line_47[105], line_46[103], line_45[101], line_44[99], line_43[97], line_42[95], line_41[93], line_40[91], line_39[89], line_38[87], line_37[85], line_36[83], line_35[81], line_34[79], line_33[77], line_32[75], line_31[73], line_30[71], line_29[69], line_28[67], line_27[65], line_26[63], line_25[61], line_24[59], line_23[57], line_22[55], line_21[53], line_20[51], line_19[49], line_18[47], line_17[45], line_16[43], line_15[41], line_14[39], line_13[37], line_12[35], line_11[33], line_10[31], line_9[29], line_8[27], line_7[25], line_6[23], line_5[21], line_4[19], line_3[17], line_2[15], line_1[13] };
assign col_268 = {line_128[268], line_127[266], line_126[264], line_125[262], line_124[260], line_123[258], line_122[256], line_121[254], line_120[252], line_119[250], line_118[248], line_117[246], line_116[244], line_115[242], line_114[240], line_113[238], line_112[236], line_111[234], line_110[232], line_109[230], line_108[228], line_107[226], line_106[224], line_105[222], line_104[220], line_103[218], line_102[216], line_101[214], line_100[212], line_99[210], line_98[208], line_97[206], line_96[204], line_95[202], line_94[200], line_93[198], line_92[196], line_91[194], line_90[192], line_89[190], line_88[188], line_87[186], line_86[184], line_85[182], line_84[180], line_83[178], line_82[176], line_81[174], line_80[172], line_79[170], line_78[168], line_77[166], line_76[164], line_75[162], line_74[160], line_73[158], line_72[156], line_71[154], line_70[152], line_69[150], line_68[148], line_67[146], line_66[144], line_65[142], line_64[140], line_63[138], line_62[136], line_61[134], line_60[132], line_59[130], line_58[128], line_57[126], line_56[124], line_55[122], line_54[120], line_53[118], line_52[116], line_51[114], line_50[112], line_49[110], line_48[108], line_47[106], line_46[104], line_45[102], line_44[100], line_43[98], line_42[96], line_41[94], line_40[92], line_39[90], line_38[88], line_37[86], line_36[84], line_35[82], line_34[80], line_33[78], line_32[76], line_31[74], line_30[72], line_29[70], line_28[68], line_27[66], line_26[64], line_25[62], line_24[60], line_23[58], line_22[56], line_21[54], line_20[52], line_19[50], line_18[48], line_17[46], line_16[44], line_15[42], line_14[40], line_13[38], line_12[36], line_11[34], line_10[32], line_9[30], line_8[28], line_7[26], line_6[24], line_5[22], line_4[20], line_3[18], line_2[16], line_1[14] };
assign col_269 = {line_128[269], line_127[267], line_126[265], line_125[263], line_124[261], line_123[259], line_122[257], line_121[255], line_120[253], line_119[251], line_118[249], line_117[247], line_116[245], line_115[243], line_114[241], line_113[239], line_112[237], line_111[235], line_110[233], line_109[231], line_108[229], line_107[227], line_106[225], line_105[223], line_104[221], line_103[219], line_102[217], line_101[215], line_100[213], line_99[211], line_98[209], line_97[207], line_96[205], line_95[203], line_94[201], line_93[199], line_92[197], line_91[195], line_90[193], line_89[191], line_88[189], line_87[187], line_86[185], line_85[183], line_84[181], line_83[179], line_82[177], line_81[175], line_80[173], line_79[171], line_78[169], line_77[167], line_76[165], line_75[163], line_74[161], line_73[159], line_72[157], line_71[155], line_70[153], line_69[151], line_68[149], line_67[147], line_66[145], line_65[143], line_64[141], line_63[139], line_62[137], line_61[135], line_60[133], line_59[131], line_58[129], line_57[127], line_56[125], line_55[123], line_54[121], line_53[119], line_52[117], line_51[115], line_50[113], line_49[111], line_48[109], line_47[107], line_46[105], line_45[103], line_44[101], line_43[99], line_42[97], line_41[95], line_40[93], line_39[91], line_38[89], line_37[87], line_36[85], line_35[83], line_34[81], line_33[79], line_32[77], line_31[75], line_30[73], line_29[71], line_28[69], line_27[67], line_26[65], line_25[63], line_24[61], line_23[59], line_22[57], line_21[55], line_20[53], line_19[51], line_18[49], line_17[47], line_16[45], line_15[43], line_14[41], line_13[39], line_12[37], line_11[35], line_10[33], line_9[31], line_8[29], line_7[27], line_6[25], line_5[23], line_4[21], line_3[19], line_2[17], line_1[15] };
assign col_270 = {line_128[270], line_127[268], line_126[266], line_125[264], line_124[262], line_123[260], line_122[258], line_121[256], line_120[254], line_119[252], line_118[250], line_117[248], line_116[246], line_115[244], line_114[242], line_113[240], line_112[238], line_111[236], line_110[234], line_109[232], line_108[230], line_107[228], line_106[226], line_105[224], line_104[222], line_103[220], line_102[218], line_101[216], line_100[214], line_99[212], line_98[210], line_97[208], line_96[206], line_95[204], line_94[202], line_93[200], line_92[198], line_91[196], line_90[194], line_89[192], line_88[190], line_87[188], line_86[186], line_85[184], line_84[182], line_83[180], line_82[178], line_81[176], line_80[174], line_79[172], line_78[170], line_77[168], line_76[166], line_75[164], line_74[162], line_73[160], line_72[158], line_71[156], line_70[154], line_69[152], line_68[150], line_67[148], line_66[146], line_65[144], line_64[142], line_63[140], line_62[138], line_61[136], line_60[134], line_59[132], line_58[130], line_57[128], line_56[126], line_55[124], line_54[122], line_53[120], line_52[118], line_51[116], line_50[114], line_49[112], line_48[110], line_47[108], line_46[106], line_45[104], line_44[102], line_43[100], line_42[98], line_41[96], line_40[94], line_39[92], line_38[90], line_37[88], line_36[86], line_35[84], line_34[82], line_33[80], line_32[78], line_31[76], line_30[74], line_29[72], line_28[70], line_27[68], line_26[66], line_25[64], line_24[62], line_23[60], line_22[58], line_21[56], line_20[54], line_19[52], line_18[50], line_17[48], line_16[46], line_15[44], line_14[42], line_13[40], line_12[38], line_11[36], line_10[34], line_9[32], line_8[30], line_7[28], line_6[26], line_5[24], line_4[22], line_3[20], line_2[18], line_1[16] };
assign col_271 = {line_128[271], line_127[269], line_126[267], line_125[265], line_124[263], line_123[261], line_122[259], line_121[257], line_120[255], line_119[253], line_118[251], line_117[249], line_116[247], line_115[245], line_114[243], line_113[241], line_112[239], line_111[237], line_110[235], line_109[233], line_108[231], line_107[229], line_106[227], line_105[225], line_104[223], line_103[221], line_102[219], line_101[217], line_100[215], line_99[213], line_98[211], line_97[209], line_96[207], line_95[205], line_94[203], line_93[201], line_92[199], line_91[197], line_90[195], line_89[193], line_88[191], line_87[189], line_86[187], line_85[185], line_84[183], line_83[181], line_82[179], line_81[177], line_80[175], line_79[173], line_78[171], line_77[169], line_76[167], line_75[165], line_74[163], line_73[161], line_72[159], line_71[157], line_70[155], line_69[153], line_68[151], line_67[149], line_66[147], line_65[145], line_64[143], line_63[141], line_62[139], line_61[137], line_60[135], line_59[133], line_58[131], line_57[129], line_56[127], line_55[125], line_54[123], line_53[121], line_52[119], line_51[117], line_50[115], line_49[113], line_48[111], line_47[109], line_46[107], line_45[105], line_44[103], line_43[101], line_42[99], line_41[97], line_40[95], line_39[93], line_38[91], line_37[89], line_36[87], line_35[85], line_34[83], line_33[81], line_32[79], line_31[77], line_30[75], line_29[73], line_28[71], line_27[69], line_26[67], line_25[65], line_24[63], line_23[61], line_22[59], line_21[57], line_20[55], line_19[53], line_18[51], line_17[49], line_16[47], line_15[45], line_14[43], line_13[41], line_12[39], line_11[37], line_10[35], line_9[33], line_8[31], line_7[29], line_6[27], line_5[25], line_4[23], line_3[21], line_2[19], line_1[17] };
assign col_272 = {line_128[272], line_127[270], line_126[268], line_125[266], line_124[264], line_123[262], line_122[260], line_121[258], line_120[256], line_119[254], line_118[252], line_117[250], line_116[248], line_115[246], line_114[244], line_113[242], line_112[240], line_111[238], line_110[236], line_109[234], line_108[232], line_107[230], line_106[228], line_105[226], line_104[224], line_103[222], line_102[220], line_101[218], line_100[216], line_99[214], line_98[212], line_97[210], line_96[208], line_95[206], line_94[204], line_93[202], line_92[200], line_91[198], line_90[196], line_89[194], line_88[192], line_87[190], line_86[188], line_85[186], line_84[184], line_83[182], line_82[180], line_81[178], line_80[176], line_79[174], line_78[172], line_77[170], line_76[168], line_75[166], line_74[164], line_73[162], line_72[160], line_71[158], line_70[156], line_69[154], line_68[152], line_67[150], line_66[148], line_65[146], line_64[144], line_63[142], line_62[140], line_61[138], line_60[136], line_59[134], line_58[132], line_57[130], line_56[128], line_55[126], line_54[124], line_53[122], line_52[120], line_51[118], line_50[116], line_49[114], line_48[112], line_47[110], line_46[108], line_45[106], line_44[104], line_43[102], line_42[100], line_41[98], line_40[96], line_39[94], line_38[92], line_37[90], line_36[88], line_35[86], line_34[84], line_33[82], line_32[80], line_31[78], line_30[76], line_29[74], line_28[72], line_27[70], line_26[68], line_25[66], line_24[64], line_23[62], line_22[60], line_21[58], line_20[56], line_19[54], line_18[52], line_17[50], line_16[48], line_15[46], line_14[44], line_13[42], line_12[40], line_11[38], line_10[36], line_9[34], line_8[32], line_7[30], line_6[28], line_5[26], line_4[24], line_3[22], line_2[20], line_1[18] };
assign col_273 = {line_128[273], line_127[271], line_126[269], line_125[267], line_124[265], line_123[263], line_122[261], line_121[259], line_120[257], line_119[255], line_118[253], line_117[251], line_116[249], line_115[247], line_114[245], line_113[243], line_112[241], line_111[239], line_110[237], line_109[235], line_108[233], line_107[231], line_106[229], line_105[227], line_104[225], line_103[223], line_102[221], line_101[219], line_100[217], line_99[215], line_98[213], line_97[211], line_96[209], line_95[207], line_94[205], line_93[203], line_92[201], line_91[199], line_90[197], line_89[195], line_88[193], line_87[191], line_86[189], line_85[187], line_84[185], line_83[183], line_82[181], line_81[179], line_80[177], line_79[175], line_78[173], line_77[171], line_76[169], line_75[167], line_74[165], line_73[163], line_72[161], line_71[159], line_70[157], line_69[155], line_68[153], line_67[151], line_66[149], line_65[147], line_64[145], line_63[143], line_62[141], line_61[139], line_60[137], line_59[135], line_58[133], line_57[131], line_56[129], line_55[127], line_54[125], line_53[123], line_52[121], line_51[119], line_50[117], line_49[115], line_48[113], line_47[111], line_46[109], line_45[107], line_44[105], line_43[103], line_42[101], line_41[99], line_40[97], line_39[95], line_38[93], line_37[91], line_36[89], line_35[87], line_34[85], line_33[83], line_32[81], line_31[79], line_30[77], line_29[75], line_28[73], line_27[71], line_26[69], line_25[67], line_24[65], line_23[63], line_22[61], line_21[59], line_20[57], line_19[55], line_18[53], line_17[51], line_16[49], line_15[47], line_14[45], line_13[43], line_12[41], line_11[39], line_10[37], line_9[35], line_8[33], line_7[31], line_6[29], line_5[27], line_4[25], line_3[23], line_2[21], line_1[19] };
assign col_274 = {line_128[274], line_127[272], line_126[270], line_125[268], line_124[266], line_123[264], line_122[262], line_121[260], line_120[258], line_119[256], line_118[254], line_117[252], line_116[250], line_115[248], line_114[246], line_113[244], line_112[242], line_111[240], line_110[238], line_109[236], line_108[234], line_107[232], line_106[230], line_105[228], line_104[226], line_103[224], line_102[222], line_101[220], line_100[218], line_99[216], line_98[214], line_97[212], line_96[210], line_95[208], line_94[206], line_93[204], line_92[202], line_91[200], line_90[198], line_89[196], line_88[194], line_87[192], line_86[190], line_85[188], line_84[186], line_83[184], line_82[182], line_81[180], line_80[178], line_79[176], line_78[174], line_77[172], line_76[170], line_75[168], line_74[166], line_73[164], line_72[162], line_71[160], line_70[158], line_69[156], line_68[154], line_67[152], line_66[150], line_65[148], line_64[146], line_63[144], line_62[142], line_61[140], line_60[138], line_59[136], line_58[134], line_57[132], line_56[130], line_55[128], line_54[126], line_53[124], line_52[122], line_51[120], line_50[118], line_49[116], line_48[114], line_47[112], line_46[110], line_45[108], line_44[106], line_43[104], line_42[102], line_41[100], line_40[98], line_39[96], line_38[94], line_37[92], line_36[90], line_35[88], line_34[86], line_33[84], line_32[82], line_31[80], line_30[78], line_29[76], line_28[74], line_27[72], line_26[70], line_25[68], line_24[66], line_23[64], line_22[62], line_21[60], line_20[58], line_19[56], line_18[54], line_17[52], line_16[50], line_15[48], line_14[46], line_13[44], line_12[42], line_11[40], line_10[38], line_9[36], line_8[34], line_7[32], line_6[30], line_5[28], line_4[26], line_3[24], line_2[22], line_1[20] };
assign col_275 = {line_128[275], line_127[273], line_126[271], line_125[269], line_124[267], line_123[265], line_122[263], line_121[261], line_120[259], line_119[257], line_118[255], line_117[253], line_116[251], line_115[249], line_114[247], line_113[245], line_112[243], line_111[241], line_110[239], line_109[237], line_108[235], line_107[233], line_106[231], line_105[229], line_104[227], line_103[225], line_102[223], line_101[221], line_100[219], line_99[217], line_98[215], line_97[213], line_96[211], line_95[209], line_94[207], line_93[205], line_92[203], line_91[201], line_90[199], line_89[197], line_88[195], line_87[193], line_86[191], line_85[189], line_84[187], line_83[185], line_82[183], line_81[181], line_80[179], line_79[177], line_78[175], line_77[173], line_76[171], line_75[169], line_74[167], line_73[165], line_72[163], line_71[161], line_70[159], line_69[157], line_68[155], line_67[153], line_66[151], line_65[149], line_64[147], line_63[145], line_62[143], line_61[141], line_60[139], line_59[137], line_58[135], line_57[133], line_56[131], line_55[129], line_54[127], line_53[125], line_52[123], line_51[121], line_50[119], line_49[117], line_48[115], line_47[113], line_46[111], line_45[109], line_44[107], line_43[105], line_42[103], line_41[101], line_40[99], line_39[97], line_38[95], line_37[93], line_36[91], line_35[89], line_34[87], line_33[85], line_32[83], line_31[81], line_30[79], line_29[77], line_28[75], line_27[73], line_26[71], line_25[69], line_24[67], line_23[65], line_22[63], line_21[61], line_20[59], line_19[57], line_18[55], line_17[53], line_16[51], line_15[49], line_14[47], line_13[45], line_12[43], line_11[41], line_10[39], line_9[37], line_8[35], line_7[33], line_6[31], line_5[29], line_4[27], line_3[25], line_2[23], line_1[21] };
assign col_276 = {line_128[276], line_127[274], line_126[272], line_125[270], line_124[268], line_123[266], line_122[264], line_121[262], line_120[260], line_119[258], line_118[256], line_117[254], line_116[252], line_115[250], line_114[248], line_113[246], line_112[244], line_111[242], line_110[240], line_109[238], line_108[236], line_107[234], line_106[232], line_105[230], line_104[228], line_103[226], line_102[224], line_101[222], line_100[220], line_99[218], line_98[216], line_97[214], line_96[212], line_95[210], line_94[208], line_93[206], line_92[204], line_91[202], line_90[200], line_89[198], line_88[196], line_87[194], line_86[192], line_85[190], line_84[188], line_83[186], line_82[184], line_81[182], line_80[180], line_79[178], line_78[176], line_77[174], line_76[172], line_75[170], line_74[168], line_73[166], line_72[164], line_71[162], line_70[160], line_69[158], line_68[156], line_67[154], line_66[152], line_65[150], line_64[148], line_63[146], line_62[144], line_61[142], line_60[140], line_59[138], line_58[136], line_57[134], line_56[132], line_55[130], line_54[128], line_53[126], line_52[124], line_51[122], line_50[120], line_49[118], line_48[116], line_47[114], line_46[112], line_45[110], line_44[108], line_43[106], line_42[104], line_41[102], line_40[100], line_39[98], line_38[96], line_37[94], line_36[92], line_35[90], line_34[88], line_33[86], line_32[84], line_31[82], line_30[80], line_29[78], line_28[76], line_27[74], line_26[72], line_25[70], line_24[68], line_23[66], line_22[64], line_21[62], line_20[60], line_19[58], line_18[56], line_17[54], line_16[52], line_15[50], line_14[48], line_13[46], line_12[44], line_11[42], line_10[40], line_9[38], line_8[36], line_7[34], line_6[32], line_5[30], line_4[28], line_3[26], line_2[24], line_1[22] };
assign col_277 = {line_128[277], line_127[275], line_126[273], line_125[271], line_124[269], line_123[267], line_122[265], line_121[263], line_120[261], line_119[259], line_118[257], line_117[255], line_116[253], line_115[251], line_114[249], line_113[247], line_112[245], line_111[243], line_110[241], line_109[239], line_108[237], line_107[235], line_106[233], line_105[231], line_104[229], line_103[227], line_102[225], line_101[223], line_100[221], line_99[219], line_98[217], line_97[215], line_96[213], line_95[211], line_94[209], line_93[207], line_92[205], line_91[203], line_90[201], line_89[199], line_88[197], line_87[195], line_86[193], line_85[191], line_84[189], line_83[187], line_82[185], line_81[183], line_80[181], line_79[179], line_78[177], line_77[175], line_76[173], line_75[171], line_74[169], line_73[167], line_72[165], line_71[163], line_70[161], line_69[159], line_68[157], line_67[155], line_66[153], line_65[151], line_64[149], line_63[147], line_62[145], line_61[143], line_60[141], line_59[139], line_58[137], line_57[135], line_56[133], line_55[131], line_54[129], line_53[127], line_52[125], line_51[123], line_50[121], line_49[119], line_48[117], line_47[115], line_46[113], line_45[111], line_44[109], line_43[107], line_42[105], line_41[103], line_40[101], line_39[99], line_38[97], line_37[95], line_36[93], line_35[91], line_34[89], line_33[87], line_32[85], line_31[83], line_30[81], line_29[79], line_28[77], line_27[75], line_26[73], line_25[71], line_24[69], line_23[67], line_22[65], line_21[63], line_20[61], line_19[59], line_18[57], line_17[55], line_16[53], line_15[51], line_14[49], line_13[47], line_12[45], line_11[43], line_10[41], line_9[39], line_8[37], line_7[35], line_6[33], line_5[31], line_4[29], line_3[27], line_2[25], line_1[23] };
assign col_278 = {line_128[278], line_127[276], line_126[274], line_125[272], line_124[270], line_123[268], line_122[266], line_121[264], line_120[262], line_119[260], line_118[258], line_117[256], line_116[254], line_115[252], line_114[250], line_113[248], line_112[246], line_111[244], line_110[242], line_109[240], line_108[238], line_107[236], line_106[234], line_105[232], line_104[230], line_103[228], line_102[226], line_101[224], line_100[222], line_99[220], line_98[218], line_97[216], line_96[214], line_95[212], line_94[210], line_93[208], line_92[206], line_91[204], line_90[202], line_89[200], line_88[198], line_87[196], line_86[194], line_85[192], line_84[190], line_83[188], line_82[186], line_81[184], line_80[182], line_79[180], line_78[178], line_77[176], line_76[174], line_75[172], line_74[170], line_73[168], line_72[166], line_71[164], line_70[162], line_69[160], line_68[158], line_67[156], line_66[154], line_65[152], line_64[150], line_63[148], line_62[146], line_61[144], line_60[142], line_59[140], line_58[138], line_57[136], line_56[134], line_55[132], line_54[130], line_53[128], line_52[126], line_51[124], line_50[122], line_49[120], line_48[118], line_47[116], line_46[114], line_45[112], line_44[110], line_43[108], line_42[106], line_41[104], line_40[102], line_39[100], line_38[98], line_37[96], line_36[94], line_35[92], line_34[90], line_33[88], line_32[86], line_31[84], line_30[82], line_29[80], line_28[78], line_27[76], line_26[74], line_25[72], line_24[70], line_23[68], line_22[66], line_21[64], line_20[62], line_19[60], line_18[58], line_17[56], line_16[54], line_15[52], line_14[50], line_13[48], line_12[46], line_11[44], line_10[42], line_9[40], line_8[38], line_7[36], line_6[34], line_5[32], line_4[30], line_3[28], line_2[26], line_1[24] };
assign col_279 = {line_128[279], line_127[277], line_126[275], line_125[273], line_124[271], line_123[269], line_122[267], line_121[265], line_120[263], line_119[261], line_118[259], line_117[257], line_116[255], line_115[253], line_114[251], line_113[249], line_112[247], line_111[245], line_110[243], line_109[241], line_108[239], line_107[237], line_106[235], line_105[233], line_104[231], line_103[229], line_102[227], line_101[225], line_100[223], line_99[221], line_98[219], line_97[217], line_96[215], line_95[213], line_94[211], line_93[209], line_92[207], line_91[205], line_90[203], line_89[201], line_88[199], line_87[197], line_86[195], line_85[193], line_84[191], line_83[189], line_82[187], line_81[185], line_80[183], line_79[181], line_78[179], line_77[177], line_76[175], line_75[173], line_74[171], line_73[169], line_72[167], line_71[165], line_70[163], line_69[161], line_68[159], line_67[157], line_66[155], line_65[153], line_64[151], line_63[149], line_62[147], line_61[145], line_60[143], line_59[141], line_58[139], line_57[137], line_56[135], line_55[133], line_54[131], line_53[129], line_52[127], line_51[125], line_50[123], line_49[121], line_48[119], line_47[117], line_46[115], line_45[113], line_44[111], line_43[109], line_42[107], line_41[105], line_40[103], line_39[101], line_38[99], line_37[97], line_36[95], line_35[93], line_34[91], line_33[89], line_32[87], line_31[85], line_30[83], line_29[81], line_28[79], line_27[77], line_26[75], line_25[73], line_24[71], line_23[69], line_22[67], line_21[65], line_20[63], line_19[61], line_18[59], line_17[57], line_16[55], line_15[53], line_14[51], line_13[49], line_12[47], line_11[45], line_10[43], line_9[41], line_8[39], line_7[37], line_6[35], line_5[33], line_4[31], line_3[29], line_2[27], line_1[25] };
assign col_280 = {line_128[280], line_127[278], line_126[276], line_125[274], line_124[272], line_123[270], line_122[268], line_121[266], line_120[264], line_119[262], line_118[260], line_117[258], line_116[256], line_115[254], line_114[252], line_113[250], line_112[248], line_111[246], line_110[244], line_109[242], line_108[240], line_107[238], line_106[236], line_105[234], line_104[232], line_103[230], line_102[228], line_101[226], line_100[224], line_99[222], line_98[220], line_97[218], line_96[216], line_95[214], line_94[212], line_93[210], line_92[208], line_91[206], line_90[204], line_89[202], line_88[200], line_87[198], line_86[196], line_85[194], line_84[192], line_83[190], line_82[188], line_81[186], line_80[184], line_79[182], line_78[180], line_77[178], line_76[176], line_75[174], line_74[172], line_73[170], line_72[168], line_71[166], line_70[164], line_69[162], line_68[160], line_67[158], line_66[156], line_65[154], line_64[152], line_63[150], line_62[148], line_61[146], line_60[144], line_59[142], line_58[140], line_57[138], line_56[136], line_55[134], line_54[132], line_53[130], line_52[128], line_51[126], line_50[124], line_49[122], line_48[120], line_47[118], line_46[116], line_45[114], line_44[112], line_43[110], line_42[108], line_41[106], line_40[104], line_39[102], line_38[100], line_37[98], line_36[96], line_35[94], line_34[92], line_33[90], line_32[88], line_31[86], line_30[84], line_29[82], line_28[80], line_27[78], line_26[76], line_25[74], line_24[72], line_23[70], line_22[68], line_21[66], line_20[64], line_19[62], line_18[60], line_17[58], line_16[56], line_15[54], line_14[52], line_13[50], line_12[48], line_11[46], line_10[44], line_9[42], line_8[40], line_7[38], line_6[36], line_5[34], line_4[32], line_3[30], line_2[28], line_1[26] };
assign col_281 = {line_128[281], line_127[279], line_126[277], line_125[275], line_124[273], line_123[271], line_122[269], line_121[267], line_120[265], line_119[263], line_118[261], line_117[259], line_116[257], line_115[255], line_114[253], line_113[251], line_112[249], line_111[247], line_110[245], line_109[243], line_108[241], line_107[239], line_106[237], line_105[235], line_104[233], line_103[231], line_102[229], line_101[227], line_100[225], line_99[223], line_98[221], line_97[219], line_96[217], line_95[215], line_94[213], line_93[211], line_92[209], line_91[207], line_90[205], line_89[203], line_88[201], line_87[199], line_86[197], line_85[195], line_84[193], line_83[191], line_82[189], line_81[187], line_80[185], line_79[183], line_78[181], line_77[179], line_76[177], line_75[175], line_74[173], line_73[171], line_72[169], line_71[167], line_70[165], line_69[163], line_68[161], line_67[159], line_66[157], line_65[155], line_64[153], line_63[151], line_62[149], line_61[147], line_60[145], line_59[143], line_58[141], line_57[139], line_56[137], line_55[135], line_54[133], line_53[131], line_52[129], line_51[127], line_50[125], line_49[123], line_48[121], line_47[119], line_46[117], line_45[115], line_44[113], line_43[111], line_42[109], line_41[107], line_40[105], line_39[103], line_38[101], line_37[99], line_36[97], line_35[95], line_34[93], line_33[91], line_32[89], line_31[87], line_30[85], line_29[83], line_28[81], line_27[79], line_26[77], line_25[75], line_24[73], line_23[71], line_22[69], line_21[67], line_20[65], line_19[63], line_18[61], line_17[59], line_16[57], line_15[55], line_14[53], line_13[51], line_12[49], line_11[47], line_10[45], line_9[43], line_8[41], line_7[39], line_6[37], line_5[35], line_4[33], line_3[31], line_2[29], line_1[27] };
assign col_282 = {line_128[282], line_127[280], line_126[278], line_125[276], line_124[274], line_123[272], line_122[270], line_121[268], line_120[266], line_119[264], line_118[262], line_117[260], line_116[258], line_115[256], line_114[254], line_113[252], line_112[250], line_111[248], line_110[246], line_109[244], line_108[242], line_107[240], line_106[238], line_105[236], line_104[234], line_103[232], line_102[230], line_101[228], line_100[226], line_99[224], line_98[222], line_97[220], line_96[218], line_95[216], line_94[214], line_93[212], line_92[210], line_91[208], line_90[206], line_89[204], line_88[202], line_87[200], line_86[198], line_85[196], line_84[194], line_83[192], line_82[190], line_81[188], line_80[186], line_79[184], line_78[182], line_77[180], line_76[178], line_75[176], line_74[174], line_73[172], line_72[170], line_71[168], line_70[166], line_69[164], line_68[162], line_67[160], line_66[158], line_65[156], line_64[154], line_63[152], line_62[150], line_61[148], line_60[146], line_59[144], line_58[142], line_57[140], line_56[138], line_55[136], line_54[134], line_53[132], line_52[130], line_51[128], line_50[126], line_49[124], line_48[122], line_47[120], line_46[118], line_45[116], line_44[114], line_43[112], line_42[110], line_41[108], line_40[106], line_39[104], line_38[102], line_37[100], line_36[98], line_35[96], line_34[94], line_33[92], line_32[90], line_31[88], line_30[86], line_29[84], line_28[82], line_27[80], line_26[78], line_25[76], line_24[74], line_23[72], line_22[70], line_21[68], line_20[66], line_19[64], line_18[62], line_17[60], line_16[58], line_15[56], line_14[54], line_13[52], line_12[50], line_11[48], line_10[46], line_9[44], line_8[42], line_7[40], line_6[38], line_5[36], line_4[34], line_3[32], line_2[30], line_1[28] };
assign col_283 = {line_128[283], line_127[281], line_126[279], line_125[277], line_124[275], line_123[273], line_122[271], line_121[269], line_120[267], line_119[265], line_118[263], line_117[261], line_116[259], line_115[257], line_114[255], line_113[253], line_112[251], line_111[249], line_110[247], line_109[245], line_108[243], line_107[241], line_106[239], line_105[237], line_104[235], line_103[233], line_102[231], line_101[229], line_100[227], line_99[225], line_98[223], line_97[221], line_96[219], line_95[217], line_94[215], line_93[213], line_92[211], line_91[209], line_90[207], line_89[205], line_88[203], line_87[201], line_86[199], line_85[197], line_84[195], line_83[193], line_82[191], line_81[189], line_80[187], line_79[185], line_78[183], line_77[181], line_76[179], line_75[177], line_74[175], line_73[173], line_72[171], line_71[169], line_70[167], line_69[165], line_68[163], line_67[161], line_66[159], line_65[157], line_64[155], line_63[153], line_62[151], line_61[149], line_60[147], line_59[145], line_58[143], line_57[141], line_56[139], line_55[137], line_54[135], line_53[133], line_52[131], line_51[129], line_50[127], line_49[125], line_48[123], line_47[121], line_46[119], line_45[117], line_44[115], line_43[113], line_42[111], line_41[109], line_40[107], line_39[105], line_38[103], line_37[101], line_36[99], line_35[97], line_34[95], line_33[93], line_32[91], line_31[89], line_30[87], line_29[85], line_28[83], line_27[81], line_26[79], line_25[77], line_24[75], line_23[73], line_22[71], line_21[69], line_20[67], line_19[65], line_18[63], line_17[61], line_16[59], line_15[57], line_14[55], line_13[53], line_12[51], line_11[49], line_10[47], line_9[45], line_8[43], line_7[41], line_6[39], line_5[37], line_4[35], line_3[33], line_2[31], line_1[29] };
assign col_284 = {line_128[284], line_127[282], line_126[280], line_125[278], line_124[276], line_123[274], line_122[272], line_121[270], line_120[268], line_119[266], line_118[264], line_117[262], line_116[260], line_115[258], line_114[256], line_113[254], line_112[252], line_111[250], line_110[248], line_109[246], line_108[244], line_107[242], line_106[240], line_105[238], line_104[236], line_103[234], line_102[232], line_101[230], line_100[228], line_99[226], line_98[224], line_97[222], line_96[220], line_95[218], line_94[216], line_93[214], line_92[212], line_91[210], line_90[208], line_89[206], line_88[204], line_87[202], line_86[200], line_85[198], line_84[196], line_83[194], line_82[192], line_81[190], line_80[188], line_79[186], line_78[184], line_77[182], line_76[180], line_75[178], line_74[176], line_73[174], line_72[172], line_71[170], line_70[168], line_69[166], line_68[164], line_67[162], line_66[160], line_65[158], line_64[156], line_63[154], line_62[152], line_61[150], line_60[148], line_59[146], line_58[144], line_57[142], line_56[140], line_55[138], line_54[136], line_53[134], line_52[132], line_51[130], line_50[128], line_49[126], line_48[124], line_47[122], line_46[120], line_45[118], line_44[116], line_43[114], line_42[112], line_41[110], line_40[108], line_39[106], line_38[104], line_37[102], line_36[100], line_35[98], line_34[96], line_33[94], line_32[92], line_31[90], line_30[88], line_29[86], line_28[84], line_27[82], line_26[80], line_25[78], line_24[76], line_23[74], line_22[72], line_21[70], line_20[68], line_19[66], line_18[64], line_17[62], line_16[60], line_15[58], line_14[56], line_13[54], line_12[52], line_11[50], line_10[48], line_9[46], line_8[44], line_7[42], line_6[40], line_5[38], line_4[36], line_3[34], line_2[32], line_1[30] };
assign col_285 = {line_128[285], line_127[283], line_126[281], line_125[279], line_124[277], line_123[275], line_122[273], line_121[271], line_120[269], line_119[267], line_118[265], line_117[263], line_116[261], line_115[259], line_114[257], line_113[255], line_112[253], line_111[251], line_110[249], line_109[247], line_108[245], line_107[243], line_106[241], line_105[239], line_104[237], line_103[235], line_102[233], line_101[231], line_100[229], line_99[227], line_98[225], line_97[223], line_96[221], line_95[219], line_94[217], line_93[215], line_92[213], line_91[211], line_90[209], line_89[207], line_88[205], line_87[203], line_86[201], line_85[199], line_84[197], line_83[195], line_82[193], line_81[191], line_80[189], line_79[187], line_78[185], line_77[183], line_76[181], line_75[179], line_74[177], line_73[175], line_72[173], line_71[171], line_70[169], line_69[167], line_68[165], line_67[163], line_66[161], line_65[159], line_64[157], line_63[155], line_62[153], line_61[151], line_60[149], line_59[147], line_58[145], line_57[143], line_56[141], line_55[139], line_54[137], line_53[135], line_52[133], line_51[131], line_50[129], line_49[127], line_48[125], line_47[123], line_46[121], line_45[119], line_44[117], line_43[115], line_42[113], line_41[111], line_40[109], line_39[107], line_38[105], line_37[103], line_36[101], line_35[99], line_34[97], line_33[95], line_32[93], line_31[91], line_30[89], line_29[87], line_28[85], line_27[83], line_26[81], line_25[79], line_24[77], line_23[75], line_22[73], line_21[71], line_20[69], line_19[67], line_18[65], line_17[63], line_16[61], line_15[59], line_14[57], line_13[55], line_12[53], line_11[51], line_10[49], line_9[47], line_8[45], line_7[43], line_6[41], line_5[39], line_4[37], line_3[35], line_2[33], line_1[31] };
assign col_286 = {line_128[286], line_127[284], line_126[282], line_125[280], line_124[278], line_123[276], line_122[274], line_121[272], line_120[270], line_119[268], line_118[266], line_117[264], line_116[262], line_115[260], line_114[258], line_113[256], line_112[254], line_111[252], line_110[250], line_109[248], line_108[246], line_107[244], line_106[242], line_105[240], line_104[238], line_103[236], line_102[234], line_101[232], line_100[230], line_99[228], line_98[226], line_97[224], line_96[222], line_95[220], line_94[218], line_93[216], line_92[214], line_91[212], line_90[210], line_89[208], line_88[206], line_87[204], line_86[202], line_85[200], line_84[198], line_83[196], line_82[194], line_81[192], line_80[190], line_79[188], line_78[186], line_77[184], line_76[182], line_75[180], line_74[178], line_73[176], line_72[174], line_71[172], line_70[170], line_69[168], line_68[166], line_67[164], line_66[162], line_65[160], line_64[158], line_63[156], line_62[154], line_61[152], line_60[150], line_59[148], line_58[146], line_57[144], line_56[142], line_55[140], line_54[138], line_53[136], line_52[134], line_51[132], line_50[130], line_49[128], line_48[126], line_47[124], line_46[122], line_45[120], line_44[118], line_43[116], line_42[114], line_41[112], line_40[110], line_39[108], line_38[106], line_37[104], line_36[102], line_35[100], line_34[98], line_33[96], line_32[94], line_31[92], line_30[90], line_29[88], line_28[86], line_27[84], line_26[82], line_25[80], line_24[78], line_23[76], line_22[74], line_21[72], line_20[70], line_19[68], line_18[66], line_17[64], line_16[62], line_15[60], line_14[58], line_13[56], line_12[54], line_11[52], line_10[50], line_9[48], line_8[46], line_7[44], line_6[42], line_5[40], line_4[38], line_3[36], line_2[34], line_1[32] };
assign col_287 = {line_128[287], line_127[285], line_126[283], line_125[281], line_124[279], line_123[277], line_122[275], line_121[273], line_120[271], line_119[269], line_118[267], line_117[265], line_116[263], line_115[261], line_114[259], line_113[257], line_112[255], line_111[253], line_110[251], line_109[249], line_108[247], line_107[245], line_106[243], line_105[241], line_104[239], line_103[237], line_102[235], line_101[233], line_100[231], line_99[229], line_98[227], line_97[225], line_96[223], line_95[221], line_94[219], line_93[217], line_92[215], line_91[213], line_90[211], line_89[209], line_88[207], line_87[205], line_86[203], line_85[201], line_84[199], line_83[197], line_82[195], line_81[193], line_80[191], line_79[189], line_78[187], line_77[185], line_76[183], line_75[181], line_74[179], line_73[177], line_72[175], line_71[173], line_70[171], line_69[169], line_68[167], line_67[165], line_66[163], line_65[161], line_64[159], line_63[157], line_62[155], line_61[153], line_60[151], line_59[149], line_58[147], line_57[145], line_56[143], line_55[141], line_54[139], line_53[137], line_52[135], line_51[133], line_50[131], line_49[129], line_48[127], line_47[125], line_46[123], line_45[121], line_44[119], line_43[117], line_42[115], line_41[113], line_40[111], line_39[109], line_38[107], line_37[105], line_36[103], line_35[101], line_34[99], line_33[97], line_32[95], line_31[93], line_30[91], line_29[89], line_28[87], line_27[85], line_26[83], line_25[81], line_24[79], line_23[77], line_22[75], line_21[73], line_20[71], line_19[69], line_18[67], line_17[65], line_16[63], line_15[61], line_14[59], line_13[57], line_12[55], line_11[53], line_10[51], line_9[49], line_8[47], line_7[45], line_6[43], line_5[41], line_4[39], line_3[37], line_2[35], line_1[33] };
assign col_288 = {line_128[288], line_127[286], line_126[284], line_125[282], line_124[280], line_123[278], line_122[276], line_121[274], line_120[272], line_119[270], line_118[268], line_117[266], line_116[264], line_115[262], line_114[260], line_113[258], line_112[256], line_111[254], line_110[252], line_109[250], line_108[248], line_107[246], line_106[244], line_105[242], line_104[240], line_103[238], line_102[236], line_101[234], line_100[232], line_99[230], line_98[228], line_97[226], line_96[224], line_95[222], line_94[220], line_93[218], line_92[216], line_91[214], line_90[212], line_89[210], line_88[208], line_87[206], line_86[204], line_85[202], line_84[200], line_83[198], line_82[196], line_81[194], line_80[192], line_79[190], line_78[188], line_77[186], line_76[184], line_75[182], line_74[180], line_73[178], line_72[176], line_71[174], line_70[172], line_69[170], line_68[168], line_67[166], line_66[164], line_65[162], line_64[160], line_63[158], line_62[156], line_61[154], line_60[152], line_59[150], line_58[148], line_57[146], line_56[144], line_55[142], line_54[140], line_53[138], line_52[136], line_51[134], line_50[132], line_49[130], line_48[128], line_47[126], line_46[124], line_45[122], line_44[120], line_43[118], line_42[116], line_41[114], line_40[112], line_39[110], line_38[108], line_37[106], line_36[104], line_35[102], line_34[100], line_33[98], line_32[96], line_31[94], line_30[92], line_29[90], line_28[88], line_27[86], line_26[84], line_25[82], line_24[80], line_23[78], line_22[76], line_21[74], line_20[72], line_19[70], line_18[68], line_17[66], line_16[64], line_15[62], line_14[60], line_13[58], line_12[56], line_11[54], line_10[52], line_9[50], line_8[48], line_7[46], line_6[44], line_5[42], line_4[40], line_3[38], line_2[36], line_1[34] };
assign col_289 = {line_128[289], line_127[287], line_126[285], line_125[283], line_124[281], line_123[279], line_122[277], line_121[275], line_120[273], line_119[271], line_118[269], line_117[267], line_116[265], line_115[263], line_114[261], line_113[259], line_112[257], line_111[255], line_110[253], line_109[251], line_108[249], line_107[247], line_106[245], line_105[243], line_104[241], line_103[239], line_102[237], line_101[235], line_100[233], line_99[231], line_98[229], line_97[227], line_96[225], line_95[223], line_94[221], line_93[219], line_92[217], line_91[215], line_90[213], line_89[211], line_88[209], line_87[207], line_86[205], line_85[203], line_84[201], line_83[199], line_82[197], line_81[195], line_80[193], line_79[191], line_78[189], line_77[187], line_76[185], line_75[183], line_74[181], line_73[179], line_72[177], line_71[175], line_70[173], line_69[171], line_68[169], line_67[167], line_66[165], line_65[163], line_64[161], line_63[159], line_62[157], line_61[155], line_60[153], line_59[151], line_58[149], line_57[147], line_56[145], line_55[143], line_54[141], line_53[139], line_52[137], line_51[135], line_50[133], line_49[131], line_48[129], line_47[127], line_46[125], line_45[123], line_44[121], line_43[119], line_42[117], line_41[115], line_40[113], line_39[111], line_38[109], line_37[107], line_36[105], line_35[103], line_34[101], line_33[99], line_32[97], line_31[95], line_30[93], line_29[91], line_28[89], line_27[87], line_26[85], line_25[83], line_24[81], line_23[79], line_22[77], line_21[75], line_20[73], line_19[71], line_18[69], line_17[67], line_16[65], line_15[63], line_14[61], line_13[59], line_12[57], line_11[55], line_10[53], line_9[51], line_8[49], line_7[47], line_6[45], line_5[43], line_4[41], line_3[39], line_2[37], line_1[35] };
assign col_290 = {line_128[290], line_127[288], line_126[286], line_125[284], line_124[282], line_123[280], line_122[278], line_121[276], line_120[274], line_119[272], line_118[270], line_117[268], line_116[266], line_115[264], line_114[262], line_113[260], line_112[258], line_111[256], line_110[254], line_109[252], line_108[250], line_107[248], line_106[246], line_105[244], line_104[242], line_103[240], line_102[238], line_101[236], line_100[234], line_99[232], line_98[230], line_97[228], line_96[226], line_95[224], line_94[222], line_93[220], line_92[218], line_91[216], line_90[214], line_89[212], line_88[210], line_87[208], line_86[206], line_85[204], line_84[202], line_83[200], line_82[198], line_81[196], line_80[194], line_79[192], line_78[190], line_77[188], line_76[186], line_75[184], line_74[182], line_73[180], line_72[178], line_71[176], line_70[174], line_69[172], line_68[170], line_67[168], line_66[166], line_65[164], line_64[162], line_63[160], line_62[158], line_61[156], line_60[154], line_59[152], line_58[150], line_57[148], line_56[146], line_55[144], line_54[142], line_53[140], line_52[138], line_51[136], line_50[134], line_49[132], line_48[130], line_47[128], line_46[126], line_45[124], line_44[122], line_43[120], line_42[118], line_41[116], line_40[114], line_39[112], line_38[110], line_37[108], line_36[106], line_35[104], line_34[102], line_33[100], line_32[98], line_31[96], line_30[94], line_29[92], line_28[90], line_27[88], line_26[86], line_25[84], line_24[82], line_23[80], line_22[78], line_21[76], line_20[74], line_19[72], line_18[70], line_17[68], line_16[66], line_15[64], line_14[62], line_13[60], line_12[58], line_11[56], line_10[54], line_9[52], line_8[50], line_7[48], line_6[46], line_5[44], line_4[42], line_3[40], line_2[38], line_1[36] };
assign col_291 = {line_128[291], line_127[289], line_126[287], line_125[285], line_124[283], line_123[281], line_122[279], line_121[277], line_120[275], line_119[273], line_118[271], line_117[269], line_116[267], line_115[265], line_114[263], line_113[261], line_112[259], line_111[257], line_110[255], line_109[253], line_108[251], line_107[249], line_106[247], line_105[245], line_104[243], line_103[241], line_102[239], line_101[237], line_100[235], line_99[233], line_98[231], line_97[229], line_96[227], line_95[225], line_94[223], line_93[221], line_92[219], line_91[217], line_90[215], line_89[213], line_88[211], line_87[209], line_86[207], line_85[205], line_84[203], line_83[201], line_82[199], line_81[197], line_80[195], line_79[193], line_78[191], line_77[189], line_76[187], line_75[185], line_74[183], line_73[181], line_72[179], line_71[177], line_70[175], line_69[173], line_68[171], line_67[169], line_66[167], line_65[165], line_64[163], line_63[161], line_62[159], line_61[157], line_60[155], line_59[153], line_58[151], line_57[149], line_56[147], line_55[145], line_54[143], line_53[141], line_52[139], line_51[137], line_50[135], line_49[133], line_48[131], line_47[129], line_46[127], line_45[125], line_44[123], line_43[121], line_42[119], line_41[117], line_40[115], line_39[113], line_38[111], line_37[109], line_36[107], line_35[105], line_34[103], line_33[101], line_32[99], line_31[97], line_30[95], line_29[93], line_28[91], line_27[89], line_26[87], line_25[85], line_24[83], line_23[81], line_22[79], line_21[77], line_20[75], line_19[73], line_18[71], line_17[69], line_16[67], line_15[65], line_14[63], line_13[61], line_12[59], line_11[57], line_10[55], line_9[53], line_8[51], line_7[49], line_6[47], line_5[45], line_4[43], line_3[41], line_2[39], line_1[37] };
assign col_292 = {line_128[292], line_127[290], line_126[288], line_125[286], line_124[284], line_123[282], line_122[280], line_121[278], line_120[276], line_119[274], line_118[272], line_117[270], line_116[268], line_115[266], line_114[264], line_113[262], line_112[260], line_111[258], line_110[256], line_109[254], line_108[252], line_107[250], line_106[248], line_105[246], line_104[244], line_103[242], line_102[240], line_101[238], line_100[236], line_99[234], line_98[232], line_97[230], line_96[228], line_95[226], line_94[224], line_93[222], line_92[220], line_91[218], line_90[216], line_89[214], line_88[212], line_87[210], line_86[208], line_85[206], line_84[204], line_83[202], line_82[200], line_81[198], line_80[196], line_79[194], line_78[192], line_77[190], line_76[188], line_75[186], line_74[184], line_73[182], line_72[180], line_71[178], line_70[176], line_69[174], line_68[172], line_67[170], line_66[168], line_65[166], line_64[164], line_63[162], line_62[160], line_61[158], line_60[156], line_59[154], line_58[152], line_57[150], line_56[148], line_55[146], line_54[144], line_53[142], line_52[140], line_51[138], line_50[136], line_49[134], line_48[132], line_47[130], line_46[128], line_45[126], line_44[124], line_43[122], line_42[120], line_41[118], line_40[116], line_39[114], line_38[112], line_37[110], line_36[108], line_35[106], line_34[104], line_33[102], line_32[100], line_31[98], line_30[96], line_29[94], line_28[92], line_27[90], line_26[88], line_25[86], line_24[84], line_23[82], line_22[80], line_21[78], line_20[76], line_19[74], line_18[72], line_17[70], line_16[68], line_15[66], line_14[64], line_13[62], line_12[60], line_11[58], line_10[56], line_9[54], line_8[52], line_7[50], line_6[48], line_5[46], line_4[44], line_3[42], line_2[40], line_1[38] };
assign col_293 = {line_128[293], line_127[291], line_126[289], line_125[287], line_124[285], line_123[283], line_122[281], line_121[279], line_120[277], line_119[275], line_118[273], line_117[271], line_116[269], line_115[267], line_114[265], line_113[263], line_112[261], line_111[259], line_110[257], line_109[255], line_108[253], line_107[251], line_106[249], line_105[247], line_104[245], line_103[243], line_102[241], line_101[239], line_100[237], line_99[235], line_98[233], line_97[231], line_96[229], line_95[227], line_94[225], line_93[223], line_92[221], line_91[219], line_90[217], line_89[215], line_88[213], line_87[211], line_86[209], line_85[207], line_84[205], line_83[203], line_82[201], line_81[199], line_80[197], line_79[195], line_78[193], line_77[191], line_76[189], line_75[187], line_74[185], line_73[183], line_72[181], line_71[179], line_70[177], line_69[175], line_68[173], line_67[171], line_66[169], line_65[167], line_64[165], line_63[163], line_62[161], line_61[159], line_60[157], line_59[155], line_58[153], line_57[151], line_56[149], line_55[147], line_54[145], line_53[143], line_52[141], line_51[139], line_50[137], line_49[135], line_48[133], line_47[131], line_46[129], line_45[127], line_44[125], line_43[123], line_42[121], line_41[119], line_40[117], line_39[115], line_38[113], line_37[111], line_36[109], line_35[107], line_34[105], line_33[103], line_32[101], line_31[99], line_30[97], line_29[95], line_28[93], line_27[91], line_26[89], line_25[87], line_24[85], line_23[83], line_22[81], line_21[79], line_20[77], line_19[75], line_18[73], line_17[71], line_16[69], line_15[67], line_14[65], line_13[63], line_12[61], line_11[59], line_10[57], line_9[55], line_8[53], line_7[51], line_6[49], line_5[47], line_4[45], line_3[43], line_2[41], line_1[39] };
assign col_294 = {line_128[294], line_127[292], line_126[290], line_125[288], line_124[286], line_123[284], line_122[282], line_121[280], line_120[278], line_119[276], line_118[274], line_117[272], line_116[270], line_115[268], line_114[266], line_113[264], line_112[262], line_111[260], line_110[258], line_109[256], line_108[254], line_107[252], line_106[250], line_105[248], line_104[246], line_103[244], line_102[242], line_101[240], line_100[238], line_99[236], line_98[234], line_97[232], line_96[230], line_95[228], line_94[226], line_93[224], line_92[222], line_91[220], line_90[218], line_89[216], line_88[214], line_87[212], line_86[210], line_85[208], line_84[206], line_83[204], line_82[202], line_81[200], line_80[198], line_79[196], line_78[194], line_77[192], line_76[190], line_75[188], line_74[186], line_73[184], line_72[182], line_71[180], line_70[178], line_69[176], line_68[174], line_67[172], line_66[170], line_65[168], line_64[166], line_63[164], line_62[162], line_61[160], line_60[158], line_59[156], line_58[154], line_57[152], line_56[150], line_55[148], line_54[146], line_53[144], line_52[142], line_51[140], line_50[138], line_49[136], line_48[134], line_47[132], line_46[130], line_45[128], line_44[126], line_43[124], line_42[122], line_41[120], line_40[118], line_39[116], line_38[114], line_37[112], line_36[110], line_35[108], line_34[106], line_33[104], line_32[102], line_31[100], line_30[98], line_29[96], line_28[94], line_27[92], line_26[90], line_25[88], line_24[86], line_23[84], line_22[82], line_21[80], line_20[78], line_19[76], line_18[74], line_17[72], line_16[70], line_15[68], line_14[66], line_13[64], line_12[62], line_11[60], line_10[58], line_9[56], line_8[54], line_7[52], line_6[50], line_5[48], line_4[46], line_3[44], line_2[42], line_1[40] };
assign col_295 = {line_128[295], line_127[293], line_126[291], line_125[289], line_124[287], line_123[285], line_122[283], line_121[281], line_120[279], line_119[277], line_118[275], line_117[273], line_116[271], line_115[269], line_114[267], line_113[265], line_112[263], line_111[261], line_110[259], line_109[257], line_108[255], line_107[253], line_106[251], line_105[249], line_104[247], line_103[245], line_102[243], line_101[241], line_100[239], line_99[237], line_98[235], line_97[233], line_96[231], line_95[229], line_94[227], line_93[225], line_92[223], line_91[221], line_90[219], line_89[217], line_88[215], line_87[213], line_86[211], line_85[209], line_84[207], line_83[205], line_82[203], line_81[201], line_80[199], line_79[197], line_78[195], line_77[193], line_76[191], line_75[189], line_74[187], line_73[185], line_72[183], line_71[181], line_70[179], line_69[177], line_68[175], line_67[173], line_66[171], line_65[169], line_64[167], line_63[165], line_62[163], line_61[161], line_60[159], line_59[157], line_58[155], line_57[153], line_56[151], line_55[149], line_54[147], line_53[145], line_52[143], line_51[141], line_50[139], line_49[137], line_48[135], line_47[133], line_46[131], line_45[129], line_44[127], line_43[125], line_42[123], line_41[121], line_40[119], line_39[117], line_38[115], line_37[113], line_36[111], line_35[109], line_34[107], line_33[105], line_32[103], line_31[101], line_30[99], line_29[97], line_28[95], line_27[93], line_26[91], line_25[89], line_24[87], line_23[85], line_22[83], line_21[81], line_20[79], line_19[77], line_18[75], line_17[73], line_16[71], line_15[69], line_14[67], line_13[65], line_12[63], line_11[61], line_10[59], line_9[57], line_8[55], line_7[53], line_6[51], line_5[49], line_4[47], line_3[45], line_2[43], line_1[41] };
assign col_296 = {line_128[296], line_127[294], line_126[292], line_125[290], line_124[288], line_123[286], line_122[284], line_121[282], line_120[280], line_119[278], line_118[276], line_117[274], line_116[272], line_115[270], line_114[268], line_113[266], line_112[264], line_111[262], line_110[260], line_109[258], line_108[256], line_107[254], line_106[252], line_105[250], line_104[248], line_103[246], line_102[244], line_101[242], line_100[240], line_99[238], line_98[236], line_97[234], line_96[232], line_95[230], line_94[228], line_93[226], line_92[224], line_91[222], line_90[220], line_89[218], line_88[216], line_87[214], line_86[212], line_85[210], line_84[208], line_83[206], line_82[204], line_81[202], line_80[200], line_79[198], line_78[196], line_77[194], line_76[192], line_75[190], line_74[188], line_73[186], line_72[184], line_71[182], line_70[180], line_69[178], line_68[176], line_67[174], line_66[172], line_65[170], line_64[168], line_63[166], line_62[164], line_61[162], line_60[160], line_59[158], line_58[156], line_57[154], line_56[152], line_55[150], line_54[148], line_53[146], line_52[144], line_51[142], line_50[140], line_49[138], line_48[136], line_47[134], line_46[132], line_45[130], line_44[128], line_43[126], line_42[124], line_41[122], line_40[120], line_39[118], line_38[116], line_37[114], line_36[112], line_35[110], line_34[108], line_33[106], line_32[104], line_31[102], line_30[100], line_29[98], line_28[96], line_27[94], line_26[92], line_25[90], line_24[88], line_23[86], line_22[84], line_21[82], line_20[80], line_19[78], line_18[76], line_17[74], line_16[72], line_15[70], line_14[68], line_13[66], line_12[64], line_11[62], line_10[60], line_9[58], line_8[56], line_7[54], line_6[52], line_5[50], line_4[48], line_3[46], line_2[44], line_1[42] };
assign col_297 = {line_128[297], line_127[295], line_126[293], line_125[291], line_124[289], line_123[287], line_122[285], line_121[283], line_120[281], line_119[279], line_118[277], line_117[275], line_116[273], line_115[271], line_114[269], line_113[267], line_112[265], line_111[263], line_110[261], line_109[259], line_108[257], line_107[255], line_106[253], line_105[251], line_104[249], line_103[247], line_102[245], line_101[243], line_100[241], line_99[239], line_98[237], line_97[235], line_96[233], line_95[231], line_94[229], line_93[227], line_92[225], line_91[223], line_90[221], line_89[219], line_88[217], line_87[215], line_86[213], line_85[211], line_84[209], line_83[207], line_82[205], line_81[203], line_80[201], line_79[199], line_78[197], line_77[195], line_76[193], line_75[191], line_74[189], line_73[187], line_72[185], line_71[183], line_70[181], line_69[179], line_68[177], line_67[175], line_66[173], line_65[171], line_64[169], line_63[167], line_62[165], line_61[163], line_60[161], line_59[159], line_58[157], line_57[155], line_56[153], line_55[151], line_54[149], line_53[147], line_52[145], line_51[143], line_50[141], line_49[139], line_48[137], line_47[135], line_46[133], line_45[131], line_44[129], line_43[127], line_42[125], line_41[123], line_40[121], line_39[119], line_38[117], line_37[115], line_36[113], line_35[111], line_34[109], line_33[107], line_32[105], line_31[103], line_30[101], line_29[99], line_28[97], line_27[95], line_26[93], line_25[91], line_24[89], line_23[87], line_22[85], line_21[83], line_20[81], line_19[79], line_18[77], line_17[75], line_16[73], line_15[71], line_14[69], line_13[67], line_12[65], line_11[63], line_10[61], line_9[59], line_8[57], line_7[55], line_6[53], line_5[51], line_4[49], line_3[47], line_2[45], line_1[43] };
assign col_298 = {line_128[298], line_127[296], line_126[294], line_125[292], line_124[290], line_123[288], line_122[286], line_121[284], line_120[282], line_119[280], line_118[278], line_117[276], line_116[274], line_115[272], line_114[270], line_113[268], line_112[266], line_111[264], line_110[262], line_109[260], line_108[258], line_107[256], line_106[254], line_105[252], line_104[250], line_103[248], line_102[246], line_101[244], line_100[242], line_99[240], line_98[238], line_97[236], line_96[234], line_95[232], line_94[230], line_93[228], line_92[226], line_91[224], line_90[222], line_89[220], line_88[218], line_87[216], line_86[214], line_85[212], line_84[210], line_83[208], line_82[206], line_81[204], line_80[202], line_79[200], line_78[198], line_77[196], line_76[194], line_75[192], line_74[190], line_73[188], line_72[186], line_71[184], line_70[182], line_69[180], line_68[178], line_67[176], line_66[174], line_65[172], line_64[170], line_63[168], line_62[166], line_61[164], line_60[162], line_59[160], line_58[158], line_57[156], line_56[154], line_55[152], line_54[150], line_53[148], line_52[146], line_51[144], line_50[142], line_49[140], line_48[138], line_47[136], line_46[134], line_45[132], line_44[130], line_43[128], line_42[126], line_41[124], line_40[122], line_39[120], line_38[118], line_37[116], line_36[114], line_35[112], line_34[110], line_33[108], line_32[106], line_31[104], line_30[102], line_29[100], line_28[98], line_27[96], line_26[94], line_25[92], line_24[90], line_23[88], line_22[86], line_21[84], line_20[82], line_19[80], line_18[78], line_17[76], line_16[74], line_15[72], line_14[70], line_13[68], line_12[66], line_11[64], line_10[62], line_9[60], line_8[58], line_7[56], line_6[54], line_5[52], line_4[50], line_3[48], line_2[46], line_1[44] };
assign col_299 = {line_128[299], line_127[297], line_126[295], line_125[293], line_124[291], line_123[289], line_122[287], line_121[285], line_120[283], line_119[281], line_118[279], line_117[277], line_116[275], line_115[273], line_114[271], line_113[269], line_112[267], line_111[265], line_110[263], line_109[261], line_108[259], line_107[257], line_106[255], line_105[253], line_104[251], line_103[249], line_102[247], line_101[245], line_100[243], line_99[241], line_98[239], line_97[237], line_96[235], line_95[233], line_94[231], line_93[229], line_92[227], line_91[225], line_90[223], line_89[221], line_88[219], line_87[217], line_86[215], line_85[213], line_84[211], line_83[209], line_82[207], line_81[205], line_80[203], line_79[201], line_78[199], line_77[197], line_76[195], line_75[193], line_74[191], line_73[189], line_72[187], line_71[185], line_70[183], line_69[181], line_68[179], line_67[177], line_66[175], line_65[173], line_64[171], line_63[169], line_62[167], line_61[165], line_60[163], line_59[161], line_58[159], line_57[157], line_56[155], line_55[153], line_54[151], line_53[149], line_52[147], line_51[145], line_50[143], line_49[141], line_48[139], line_47[137], line_46[135], line_45[133], line_44[131], line_43[129], line_42[127], line_41[125], line_40[123], line_39[121], line_38[119], line_37[117], line_36[115], line_35[113], line_34[111], line_33[109], line_32[107], line_31[105], line_30[103], line_29[101], line_28[99], line_27[97], line_26[95], line_25[93], line_24[91], line_23[89], line_22[87], line_21[85], line_20[83], line_19[81], line_18[79], line_17[77], line_16[75], line_15[73], line_14[71], line_13[69], line_12[67], line_11[65], line_10[63], line_9[61], line_8[59], line_7[57], line_6[55], line_5[53], line_4[51], line_3[49], line_2[47], line_1[45] };
assign col_300 = {line_128[300], line_127[298], line_126[296], line_125[294], line_124[292], line_123[290], line_122[288], line_121[286], line_120[284], line_119[282], line_118[280], line_117[278], line_116[276], line_115[274], line_114[272], line_113[270], line_112[268], line_111[266], line_110[264], line_109[262], line_108[260], line_107[258], line_106[256], line_105[254], line_104[252], line_103[250], line_102[248], line_101[246], line_100[244], line_99[242], line_98[240], line_97[238], line_96[236], line_95[234], line_94[232], line_93[230], line_92[228], line_91[226], line_90[224], line_89[222], line_88[220], line_87[218], line_86[216], line_85[214], line_84[212], line_83[210], line_82[208], line_81[206], line_80[204], line_79[202], line_78[200], line_77[198], line_76[196], line_75[194], line_74[192], line_73[190], line_72[188], line_71[186], line_70[184], line_69[182], line_68[180], line_67[178], line_66[176], line_65[174], line_64[172], line_63[170], line_62[168], line_61[166], line_60[164], line_59[162], line_58[160], line_57[158], line_56[156], line_55[154], line_54[152], line_53[150], line_52[148], line_51[146], line_50[144], line_49[142], line_48[140], line_47[138], line_46[136], line_45[134], line_44[132], line_43[130], line_42[128], line_41[126], line_40[124], line_39[122], line_38[120], line_37[118], line_36[116], line_35[114], line_34[112], line_33[110], line_32[108], line_31[106], line_30[104], line_29[102], line_28[100], line_27[98], line_26[96], line_25[94], line_24[92], line_23[90], line_22[88], line_21[86], line_20[84], line_19[82], line_18[80], line_17[78], line_16[76], line_15[74], line_14[72], line_13[70], line_12[68], line_11[66], line_10[64], line_9[62], line_8[60], line_7[58], line_6[56], line_5[54], line_4[52], line_3[50], line_2[48], line_1[46] };
assign col_301 = {line_128[301], line_127[299], line_126[297], line_125[295], line_124[293], line_123[291], line_122[289], line_121[287], line_120[285], line_119[283], line_118[281], line_117[279], line_116[277], line_115[275], line_114[273], line_113[271], line_112[269], line_111[267], line_110[265], line_109[263], line_108[261], line_107[259], line_106[257], line_105[255], line_104[253], line_103[251], line_102[249], line_101[247], line_100[245], line_99[243], line_98[241], line_97[239], line_96[237], line_95[235], line_94[233], line_93[231], line_92[229], line_91[227], line_90[225], line_89[223], line_88[221], line_87[219], line_86[217], line_85[215], line_84[213], line_83[211], line_82[209], line_81[207], line_80[205], line_79[203], line_78[201], line_77[199], line_76[197], line_75[195], line_74[193], line_73[191], line_72[189], line_71[187], line_70[185], line_69[183], line_68[181], line_67[179], line_66[177], line_65[175], line_64[173], line_63[171], line_62[169], line_61[167], line_60[165], line_59[163], line_58[161], line_57[159], line_56[157], line_55[155], line_54[153], line_53[151], line_52[149], line_51[147], line_50[145], line_49[143], line_48[141], line_47[139], line_46[137], line_45[135], line_44[133], line_43[131], line_42[129], line_41[127], line_40[125], line_39[123], line_38[121], line_37[119], line_36[117], line_35[115], line_34[113], line_33[111], line_32[109], line_31[107], line_30[105], line_29[103], line_28[101], line_27[99], line_26[97], line_25[95], line_24[93], line_23[91], line_22[89], line_21[87], line_20[85], line_19[83], line_18[81], line_17[79], line_16[77], line_15[75], line_14[73], line_13[71], line_12[69], line_11[67], line_10[65], line_9[63], line_8[61], line_7[59], line_6[57], line_5[55], line_4[53], line_3[51], line_2[49], line_1[47] };
assign col_302 = {line_128[302], line_127[300], line_126[298], line_125[296], line_124[294], line_123[292], line_122[290], line_121[288], line_120[286], line_119[284], line_118[282], line_117[280], line_116[278], line_115[276], line_114[274], line_113[272], line_112[270], line_111[268], line_110[266], line_109[264], line_108[262], line_107[260], line_106[258], line_105[256], line_104[254], line_103[252], line_102[250], line_101[248], line_100[246], line_99[244], line_98[242], line_97[240], line_96[238], line_95[236], line_94[234], line_93[232], line_92[230], line_91[228], line_90[226], line_89[224], line_88[222], line_87[220], line_86[218], line_85[216], line_84[214], line_83[212], line_82[210], line_81[208], line_80[206], line_79[204], line_78[202], line_77[200], line_76[198], line_75[196], line_74[194], line_73[192], line_72[190], line_71[188], line_70[186], line_69[184], line_68[182], line_67[180], line_66[178], line_65[176], line_64[174], line_63[172], line_62[170], line_61[168], line_60[166], line_59[164], line_58[162], line_57[160], line_56[158], line_55[156], line_54[154], line_53[152], line_52[150], line_51[148], line_50[146], line_49[144], line_48[142], line_47[140], line_46[138], line_45[136], line_44[134], line_43[132], line_42[130], line_41[128], line_40[126], line_39[124], line_38[122], line_37[120], line_36[118], line_35[116], line_34[114], line_33[112], line_32[110], line_31[108], line_30[106], line_29[104], line_28[102], line_27[100], line_26[98], line_25[96], line_24[94], line_23[92], line_22[90], line_21[88], line_20[86], line_19[84], line_18[82], line_17[80], line_16[78], line_15[76], line_14[74], line_13[72], line_12[70], line_11[68], line_10[66], line_9[64], line_8[62], line_7[60], line_6[58], line_5[56], line_4[54], line_3[52], line_2[50], line_1[48] };
assign col_303 = {line_128[303], line_127[301], line_126[299], line_125[297], line_124[295], line_123[293], line_122[291], line_121[289], line_120[287], line_119[285], line_118[283], line_117[281], line_116[279], line_115[277], line_114[275], line_113[273], line_112[271], line_111[269], line_110[267], line_109[265], line_108[263], line_107[261], line_106[259], line_105[257], line_104[255], line_103[253], line_102[251], line_101[249], line_100[247], line_99[245], line_98[243], line_97[241], line_96[239], line_95[237], line_94[235], line_93[233], line_92[231], line_91[229], line_90[227], line_89[225], line_88[223], line_87[221], line_86[219], line_85[217], line_84[215], line_83[213], line_82[211], line_81[209], line_80[207], line_79[205], line_78[203], line_77[201], line_76[199], line_75[197], line_74[195], line_73[193], line_72[191], line_71[189], line_70[187], line_69[185], line_68[183], line_67[181], line_66[179], line_65[177], line_64[175], line_63[173], line_62[171], line_61[169], line_60[167], line_59[165], line_58[163], line_57[161], line_56[159], line_55[157], line_54[155], line_53[153], line_52[151], line_51[149], line_50[147], line_49[145], line_48[143], line_47[141], line_46[139], line_45[137], line_44[135], line_43[133], line_42[131], line_41[129], line_40[127], line_39[125], line_38[123], line_37[121], line_36[119], line_35[117], line_34[115], line_33[113], line_32[111], line_31[109], line_30[107], line_29[105], line_28[103], line_27[101], line_26[99], line_25[97], line_24[95], line_23[93], line_22[91], line_21[89], line_20[87], line_19[85], line_18[83], line_17[81], line_16[79], line_15[77], line_14[75], line_13[73], line_12[71], line_11[69], line_10[67], line_9[65], line_8[63], line_7[61], line_6[59], line_5[57], line_4[55], line_3[53], line_2[51], line_1[49] };
assign col_304 = {line_128[304], line_127[302], line_126[300], line_125[298], line_124[296], line_123[294], line_122[292], line_121[290], line_120[288], line_119[286], line_118[284], line_117[282], line_116[280], line_115[278], line_114[276], line_113[274], line_112[272], line_111[270], line_110[268], line_109[266], line_108[264], line_107[262], line_106[260], line_105[258], line_104[256], line_103[254], line_102[252], line_101[250], line_100[248], line_99[246], line_98[244], line_97[242], line_96[240], line_95[238], line_94[236], line_93[234], line_92[232], line_91[230], line_90[228], line_89[226], line_88[224], line_87[222], line_86[220], line_85[218], line_84[216], line_83[214], line_82[212], line_81[210], line_80[208], line_79[206], line_78[204], line_77[202], line_76[200], line_75[198], line_74[196], line_73[194], line_72[192], line_71[190], line_70[188], line_69[186], line_68[184], line_67[182], line_66[180], line_65[178], line_64[176], line_63[174], line_62[172], line_61[170], line_60[168], line_59[166], line_58[164], line_57[162], line_56[160], line_55[158], line_54[156], line_53[154], line_52[152], line_51[150], line_50[148], line_49[146], line_48[144], line_47[142], line_46[140], line_45[138], line_44[136], line_43[134], line_42[132], line_41[130], line_40[128], line_39[126], line_38[124], line_37[122], line_36[120], line_35[118], line_34[116], line_33[114], line_32[112], line_31[110], line_30[108], line_29[106], line_28[104], line_27[102], line_26[100], line_25[98], line_24[96], line_23[94], line_22[92], line_21[90], line_20[88], line_19[86], line_18[84], line_17[82], line_16[80], line_15[78], line_14[76], line_13[74], line_12[72], line_11[70], line_10[68], line_9[66], line_8[64], line_7[62], line_6[60], line_5[58], line_4[56], line_3[54], line_2[52], line_1[50] };
assign col_305 = {line_128[305], line_127[303], line_126[301], line_125[299], line_124[297], line_123[295], line_122[293], line_121[291], line_120[289], line_119[287], line_118[285], line_117[283], line_116[281], line_115[279], line_114[277], line_113[275], line_112[273], line_111[271], line_110[269], line_109[267], line_108[265], line_107[263], line_106[261], line_105[259], line_104[257], line_103[255], line_102[253], line_101[251], line_100[249], line_99[247], line_98[245], line_97[243], line_96[241], line_95[239], line_94[237], line_93[235], line_92[233], line_91[231], line_90[229], line_89[227], line_88[225], line_87[223], line_86[221], line_85[219], line_84[217], line_83[215], line_82[213], line_81[211], line_80[209], line_79[207], line_78[205], line_77[203], line_76[201], line_75[199], line_74[197], line_73[195], line_72[193], line_71[191], line_70[189], line_69[187], line_68[185], line_67[183], line_66[181], line_65[179], line_64[177], line_63[175], line_62[173], line_61[171], line_60[169], line_59[167], line_58[165], line_57[163], line_56[161], line_55[159], line_54[157], line_53[155], line_52[153], line_51[151], line_50[149], line_49[147], line_48[145], line_47[143], line_46[141], line_45[139], line_44[137], line_43[135], line_42[133], line_41[131], line_40[129], line_39[127], line_38[125], line_37[123], line_36[121], line_35[119], line_34[117], line_33[115], line_32[113], line_31[111], line_30[109], line_29[107], line_28[105], line_27[103], line_26[101], line_25[99], line_24[97], line_23[95], line_22[93], line_21[91], line_20[89], line_19[87], line_18[85], line_17[83], line_16[81], line_15[79], line_14[77], line_13[75], line_12[73], line_11[71], line_10[69], line_9[67], line_8[65], line_7[63], line_6[61], line_5[59], line_4[57], line_3[55], line_2[53], line_1[51] };
assign col_306 = {line_128[306], line_127[304], line_126[302], line_125[300], line_124[298], line_123[296], line_122[294], line_121[292], line_120[290], line_119[288], line_118[286], line_117[284], line_116[282], line_115[280], line_114[278], line_113[276], line_112[274], line_111[272], line_110[270], line_109[268], line_108[266], line_107[264], line_106[262], line_105[260], line_104[258], line_103[256], line_102[254], line_101[252], line_100[250], line_99[248], line_98[246], line_97[244], line_96[242], line_95[240], line_94[238], line_93[236], line_92[234], line_91[232], line_90[230], line_89[228], line_88[226], line_87[224], line_86[222], line_85[220], line_84[218], line_83[216], line_82[214], line_81[212], line_80[210], line_79[208], line_78[206], line_77[204], line_76[202], line_75[200], line_74[198], line_73[196], line_72[194], line_71[192], line_70[190], line_69[188], line_68[186], line_67[184], line_66[182], line_65[180], line_64[178], line_63[176], line_62[174], line_61[172], line_60[170], line_59[168], line_58[166], line_57[164], line_56[162], line_55[160], line_54[158], line_53[156], line_52[154], line_51[152], line_50[150], line_49[148], line_48[146], line_47[144], line_46[142], line_45[140], line_44[138], line_43[136], line_42[134], line_41[132], line_40[130], line_39[128], line_38[126], line_37[124], line_36[122], line_35[120], line_34[118], line_33[116], line_32[114], line_31[112], line_30[110], line_29[108], line_28[106], line_27[104], line_26[102], line_25[100], line_24[98], line_23[96], line_22[94], line_21[92], line_20[90], line_19[88], line_18[86], line_17[84], line_16[82], line_15[80], line_14[78], line_13[76], line_12[74], line_11[72], line_10[70], line_9[68], line_8[66], line_7[64], line_6[62], line_5[60], line_4[58], line_3[56], line_2[54], line_1[52] };
assign col_307 = {line_128[307], line_127[305], line_126[303], line_125[301], line_124[299], line_123[297], line_122[295], line_121[293], line_120[291], line_119[289], line_118[287], line_117[285], line_116[283], line_115[281], line_114[279], line_113[277], line_112[275], line_111[273], line_110[271], line_109[269], line_108[267], line_107[265], line_106[263], line_105[261], line_104[259], line_103[257], line_102[255], line_101[253], line_100[251], line_99[249], line_98[247], line_97[245], line_96[243], line_95[241], line_94[239], line_93[237], line_92[235], line_91[233], line_90[231], line_89[229], line_88[227], line_87[225], line_86[223], line_85[221], line_84[219], line_83[217], line_82[215], line_81[213], line_80[211], line_79[209], line_78[207], line_77[205], line_76[203], line_75[201], line_74[199], line_73[197], line_72[195], line_71[193], line_70[191], line_69[189], line_68[187], line_67[185], line_66[183], line_65[181], line_64[179], line_63[177], line_62[175], line_61[173], line_60[171], line_59[169], line_58[167], line_57[165], line_56[163], line_55[161], line_54[159], line_53[157], line_52[155], line_51[153], line_50[151], line_49[149], line_48[147], line_47[145], line_46[143], line_45[141], line_44[139], line_43[137], line_42[135], line_41[133], line_40[131], line_39[129], line_38[127], line_37[125], line_36[123], line_35[121], line_34[119], line_33[117], line_32[115], line_31[113], line_30[111], line_29[109], line_28[107], line_27[105], line_26[103], line_25[101], line_24[99], line_23[97], line_22[95], line_21[93], line_20[91], line_19[89], line_18[87], line_17[85], line_16[83], line_15[81], line_14[79], line_13[77], line_12[75], line_11[73], line_10[71], line_9[69], line_8[67], line_7[65], line_6[63], line_5[61], line_4[59], line_3[57], line_2[55], line_1[53] };
assign col_308 = {line_128[308], line_127[306], line_126[304], line_125[302], line_124[300], line_123[298], line_122[296], line_121[294], line_120[292], line_119[290], line_118[288], line_117[286], line_116[284], line_115[282], line_114[280], line_113[278], line_112[276], line_111[274], line_110[272], line_109[270], line_108[268], line_107[266], line_106[264], line_105[262], line_104[260], line_103[258], line_102[256], line_101[254], line_100[252], line_99[250], line_98[248], line_97[246], line_96[244], line_95[242], line_94[240], line_93[238], line_92[236], line_91[234], line_90[232], line_89[230], line_88[228], line_87[226], line_86[224], line_85[222], line_84[220], line_83[218], line_82[216], line_81[214], line_80[212], line_79[210], line_78[208], line_77[206], line_76[204], line_75[202], line_74[200], line_73[198], line_72[196], line_71[194], line_70[192], line_69[190], line_68[188], line_67[186], line_66[184], line_65[182], line_64[180], line_63[178], line_62[176], line_61[174], line_60[172], line_59[170], line_58[168], line_57[166], line_56[164], line_55[162], line_54[160], line_53[158], line_52[156], line_51[154], line_50[152], line_49[150], line_48[148], line_47[146], line_46[144], line_45[142], line_44[140], line_43[138], line_42[136], line_41[134], line_40[132], line_39[130], line_38[128], line_37[126], line_36[124], line_35[122], line_34[120], line_33[118], line_32[116], line_31[114], line_30[112], line_29[110], line_28[108], line_27[106], line_26[104], line_25[102], line_24[100], line_23[98], line_22[96], line_21[94], line_20[92], line_19[90], line_18[88], line_17[86], line_16[84], line_15[82], line_14[80], line_13[78], line_12[76], line_11[74], line_10[72], line_9[70], line_8[68], line_7[66], line_6[64], line_5[62], line_4[60], line_3[58], line_2[56], line_1[54] };
assign col_309 = {line_128[309], line_127[307], line_126[305], line_125[303], line_124[301], line_123[299], line_122[297], line_121[295], line_120[293], line_119[291], line_118[289], line_117[287], line_116[285], line_115[283], line_114[281], line_113[279], line_112[277], line_111[275], line_110[273], line_109[271], line_108[269], line_107[267], line_106[265], line_105[263], line_104[261], line_103[259], line_102[257], line_101[255], line_100[253], line_99[251], line_98[249], line_97[247], line_96[245], line_95[243], line_94[241], line_93[239], line_92[237], line_91[235], line_90[233], line_89[231], line_88[229], line_87[227], line_86[225], line_85[223], line_84[221], line_83[219], line_82[217], line_81[215], line_80[213], line_79[211], line_78[209], line_77[207], line_76[205], line_75[203], line_74[201], line_73[199], line_72[197], line_71[195], line_70[193], line_69[191], line_68[189], line_67[187], line_66[185], line_65[183], line_64[181], line_63[179], line_62[177], line_61[175], line_60[173], line_59[171], line_58[169], line_57[167], line_56[165], line_55[163], line_54[161], line_53[159], line_52[157], line_51[155], line_50[153], line_49[151], line_48[149], line_47[147], line_46[145], line_45[143], line_44[141], line_43[139], line_42[137], line_41[135], line_40[133], line_39[131], line_38[129], line_37[127], line_36[125], line_35[123], line_34[121], line_33[119], line_32[117], line_31[115], line_30[113], line_29[111], line_28[109], line_27[107], line_26[105], line_25[103], line_24[101], line_23[99], line_22[97], line_21[95], line_20[93], line_19[91], line_18[89], line_17[87], line_16[85], line_15[83], line_14[81], line_13[79], line_12[77], line_11[75], line_10[73], line_9[71], line_8[69], line_7[67], line_6[65], line_5[63], line_4[61], line_3[59], line_2[57], line_1[55] };
assign col_310 = {line_128[310], line_127[308], line_126[306], line_125[304], line_124[302], line_123[300], line_122[298], line_121[296], line_120[294], line_119[292], line_118[290], line_117[288], line_116[286], line_115[284], line_114[282], line_113[280], line_112[278], line_111[276], line_110[274], line_109[272], line_108[270], line_107[268], line_106[266], line_105[264], line_104[262], line_103[260], line_102[258], line_101[256], line_100[254], line_99[252], line_98[250], line_97[248], line_96[246], line_95[244], line_94[242], line_93[240], line_92[238], line_91[236], line_90[234], line_89[232], line_88[230], line_87[228], line_86[226], line_85[224], line_84[222], line_83[220], line_82[218], line_81[216], line_80[214], line_79[212], line_78[210], line_77[208], line_76[206], line_75[204], line_74[202], line_73[200], line_72[198], line_71[196], line_70[194], line_69[192], line_68[190], line_67[188], line_66[186], line_65[184], line_64[182], line_63[180], line_62[178], line_61[176], line_60[174], line_59[172], line_58[170], line_57[168], line_56[166], line_55[164], line_54[162], line_53[160], line_52[158], line_51[156], line_50[154], line_49[152], line_48[150], line_47[148], line_46[146], line_45[144], line_44[142], line_43[140], line_42[138], line_41[136], line_40[134], line_39[132], line_38[130], line_37[128], line_36[126], line_35[124], line_34[122], line_33[120], line_32[118], line_31[116], line_30[114], line_29[112], line_28[110], line_27[108], line_26[106], line_25[104], line_24[102], line_23[100], line_22[98], line_21[96], line_20[94], line_19[92], line_18[90], line_17[88], line_16[86], line_15[84], line_14[82], line_13[80], line_12[78], line_11[76], line_10[74], line_9[72], line_8[70], line_7[68], line_6[66], line_5[64], line_4[62], line_3[60], line_2[58], line_1[56] };
assign col_311 = {line_128[311], line_127[309], line_126[307], line_125[305], line_124[303], line_123[301], line_122[299], line_121[297], line_120[295], line_119[293], line_118[291], line_117[289], line_116[287], line_115[285], line_114[283], line_113[281], line_112[279], line_111[277], line_110[275], line_109[273], line_108[271], line_107[269], line_106[267], line_105[265], line_104[263], line_103[261], line_102[259], line_101[257], line_100[255], line_99[253], line_98[251], line_97[249], line_96[247], line_95[245], line_94[243], line_93[241], line_92[239], line_91[237], line_90[235], line_89[233], line_88[231], line_87[229], line_86[227], line_85[225], line_84[223], line_83[221], line_82[219], line_81[217], line_80[215], line_79[213], line_78[211], line_77[209], line_76[207], line_75[205], line_74[203], line_73[201], line_72[199], line_71[197], line_70[195], line_69[193], line_68[191], line_67[189], line_66[187], line_65[185], line_64[183], line_63[181], line_62[179], line_61[177], line_60[175], line_59[173], line_58[171], line_57[169], line_56[167], line_55[165], line_54[163], line_53[161], line_52[159], line_51[157], line_50[155], line_49[153], line_48[151], line_47[149], line_46[147], line_45[145], line_44[143], line_43[141], line_42[139], line_41[137], line_40[135], line_39[133], line_38[131], line_37[129], line_36[127], line_35[125], line_34[123], line_33[121], line_32[119], line_31[117], line_30[115], line_29[113], line_28[111], line_27[109], line_26[107], line_25[105], line_24[103], line_23[101], line_22[99], line_21[97], line_20[95], line_19[93], line_18[91], line_17[89], line_16[87], line_15[85], line_14[83], line_13[81], line_12[79], line_11[77], line_10[75], line_9[73], line_8[71], line_7[69], line_6[67], line_5[65], line_4[63], line_3[61], line_2[59], line_1[57] };
assign col_312 = {line_128[312], line_127[310], line_126[308], line_125[306], line_124[304], line_123[302], line_122[300], line_121[298], line_120[296], line_119[294], line_118[292], line_117[290], line_116[288], line_115[286], line_114[284], line_113[282], line_112[280], line_111[278], line_110[276], line_109[274], line_108[272], line_107[270], line_106[268], line_105[266], line_104[264], line_103[262], line_102[260], line_101[258], line_100[256], line_99[254], line_98[252], line_97[250], line_96[248], line_95[246], line_94[244], line_93[242], line_92[240], line_91[238], line_90[236], line_89[234], line_88[232], line_87[230], line_86[228], line_85[226], line_84[224], line_83[222], line_82[220], line_81[218], line_80[216], line_79[214], line_78[212], line_77[210], line_76[208], line_75[206], line_74[204], line_73[202], line_72[200], line_71[198], line_70[196], line_69[194], line_68[192], line_67[190], line_66[188], line_65[186], line_64[184], line_63[182], line_62[180], line_61[178], line_60[176], line_59[174], line_58[172], line_57[170], line_56[168], line_55[166], line_54[164], line_53[162], line_52[160], line_51[158], line_50[156], line_49[154], line_48[152], line_47[150], line_46[148], line_45[146], line_44[144], line_43[142], line_42[140], line_41[138], line_40[136], line_39[134], line_38[132], line_37[130], line_36[128], line_35[126], line_34[124], line_33[122], line_32[120], line_31[118], line_30[116], line_29[114], line_28[112], line_27[110], line_26[108], line_25[106], line_24[104], line_23[102], line_22[100], line_21[98], line_20[96], line_19[94], line_18[92], line_17[90], line_16[88], line_15[86], line_14[84], line_13[82], line_12[80], line_11[78], line_10[76], line_9[74], line_8[72], line_7[70], line_6[68], line_5[66], line_4[64], line_3[62], line_2[60], line_1[58] };
assign col_313 = {line_128[313], line_127[311], line_126[309], line_125[307], line_124[305], line_123[303], line_122[301], line_121[299], line_120[297], line_119[295], line_118[293], line_117[291], line_116[289], line_115[287], line_114[285], line_113[283], line_112[281], line_111[279], line_110[277], line_109[275], line_108[273], line_107[271], line_106[269], line_105[267], line_104[265], line_103[263], line_102[261], line_101[259], line_100[257], line_99[255], line_98[253], line_97[251], line_96[249], line_95[247], line_94[245], line_93[243], line_92[241], line_91[239], line_90[237], line_89[235], line_88[233], line_87[231], line_86[229], line_85[227], line_84[225], line_83[223], line_82[221], line_81[219], line_80[217], line_79[215], line_78[213], line_77[211], line_76[209], line_75[207], line_74[205], line_73[203], line_72[201], line_71[199], line_70[197], line_69[195], line_68[193], line_67[191], line_66[189], line_65[187], line_64[185], line_63[183], line_62[181], line_61[179], line_60[177], line_59[175], line_58[173], line_57[171], line_56[169], line_55[167], line_54[165], line_53[163], line_52[161], line_51[159], line_50[157], line_49[155], line_48[153], line_47[151], line_46[149], line_45[147], line_44[145], line_43[143], line_42[141], line_41[139], line_40[137], line_39[135], line_38[133], line_37[131], line_36[129], line_35[127], line_34[125], line_33[123], line_32[121], line_31[119], line_30[117], line_29[115], line_28[113], line_27[111], line_26[109], line_25[107], line_24[105], line_23[103], line_22[101], line_21[99], line_20[97], line_19[95], line_18[93], line_17[91], line_16[89], line_15[87], line_14[85], line_13[83], line_12[81], line_11[79], line_10[77], line_9[75], line_8[73], line_7[71], line_6[69], line_5[67], line_4[65], line_3[63], line_2[61], line_1[59] };
assign col_314 = {line_128[314], line_127[312], line_126[310], line_125[308], line_124[306], line_123[304], line_122[302], line_121[300], line_120[298], line_119[296], line_118[294], line_117[292], line_116[290], line_115[288], line_114[286], line_113[284], line_112[282], line_111[280], line_110[278], line_109[276], line_108[274], line_107[272], line_106[270], line_105[268], line_104[266], line_103[264], line_102[262], line_101[260], line_100[258], line_99[256], line_98[254], line_97[252], line_96[250], line_95[248], line_94[246], line_93[244], line_92[242], line_91[240], line_90[238], line_89[236], line_88[234], line_87[232], line_86[230], line_85[228], line_84[226], line_83[224], line_82[222], line_81[220], line_80[218], line_79[216], line_78[214], line_77[212], line_76[210], line_75[208], line_74[206], line_73[204], line_72[202], line_71[200], line_70[198], line_69[196], line_68[194], line_67[192], line_66[190], line_65[188], line_64[186], line_63[184], line_62[182], line_61[180], line_60[178], line_59[176], line_58[174], line_57[172], line_56[170], line_55[168], line_54[166], line_53[164], line_52[162], line_51[160], line_50[158], line_49[156], line_48[154], line_47[152], line_46[150], line_45[148], line_44[146], line_43[144], line_42[142], line_41[140], line_40[138], line_39[136], line_38[134], line_37[132], line_36[130], line_35[128], line_34[126], line_33[124], line_32[122], line_31[120], line_30[118], line_29[116], line_28[114], line_27[112], line_26[110], line_25[108], line_24[106], line_23[104], line_22[102], line_21[100], line_20[98], line_19[96], line_18[94], line_17[92], line_16[90], line_15[88], line_14[86], line_13[84], line_12[82], line_11[80], line_10[78], line_9[76], line_8[74], line_7[72], line_6[70], line_5[68], line_4[66], line_3[64], line_2[62], line_1[60] };
assign col_315 = {line_128[315], line_127[313], line_126[311], line_125[309], line_124[307], line_123[305], line_122[303], line_121[301], line_120[299], line_119[297], line_118[295], line_117[293], line_116[291], line_115[289], line_114[287], line_113[285], line_112[283], line_111[281], line_110[279], line_109[277], line_108[275], line_107[273], line_106[271], line_105[269], line_104[267], line_103[265], line_102[263], line_101[261], line_100[259], line_99[257], line_98[255], line_97[253], line_96[251], line_95[249], line_94[247], line_93[245], line_92[243], line_91[241], line_90[239], line_89[237], line_88[235], line_87[233], line_86[231], line_85[229], line_84[227], line_83[225], line_82[223], line_81[221], line_80[219], line_79[217], line_78[215], line_77[213], line_76[211], line_75[209], line_74[207], line_73[205], line_72[203], line_71[201], line_70[199], line_69[197], line_68[195], line_67[193], line_66[191], line_65[189], line_64[187], line_63[185], line_62[183], line_61[181], line_60[179], line_59[177], line_58[175], line_57[173], line_56[171], line_55[169], line_54[167], line_53[165], line_52[163], line_51[161], line_50[159], line_49[157], line_48[155], line_47[153], line_46[151], line_45[149], line_44[147], line_43[145], line_42[143], line_41[141], line_40[139], line_39[137], line_38[135], line_37[133], line_36[131], line_35[129], line_34[127], line_33[125], line_32[123], line_31[121], line_30[119], line_29[117], line_28[115], line_27[113], line_26[111], line_25[109], line_24[107], line_23[105], line_22[103], line_21[101], line_20[99], line_19[97], line_18[95], line_17[93], line_16[91], line_15[89], line_14[87], line_13[85], line_12[83], line_11[81], line_10[79], line_9[77], line_8[75], line_7[73], line_6[71], line_5[69], line_4[67], line_3[65], line_2[63], line_1[61] };
assign col_316 = {line_128[316], line_127[314], line_126[312], line_125[310], line_124[308], line_123[306], line_122[304], line_121[302], line_120[300], line_119[298], line_118[296], line_117[294], line_116[292], line_115[290], line_114[288], line_113[286], line_112[284], line_111[282], line_110[280], line_109[278], line_108[276], line_107[274], line_106[272], line_105[270], line_104[268], line_103[266], line_102[264], line_101[262], line_100[260], line_99[258], line_98[256], line_97[254], line_96[252], line_95[250], line_94[248], line_93[246], line_92[244], line_91[242], line_90[240], line_89[238], line_88[236], line_87[234], line_86[232], line_85[230], line_84[228], line_83[226], line_82[224], line_81[222], line_80[220], line_79[218], line_78[216], line_77[214], line_76[212], line_75[210], line_74[208], line_73[206], line_72[204], line_71[202], line_70[200], line_69[198], line_68[196], line_67[194], line_66[192], line_65[190], line_64[188], line_63[186], line_62[184], line_61[182], line_60[180], line_59[178], line_58[176], line_57[174], line_56[172], line_55[170], line_54[168], line_53[166], line_52[164], line_51[162], line_50[160], line_49[158], line_48[156], line_47[154], line_46[152], line_45[150], line_44[148], line_43[146], line_42[144], line_41[142], line_40[140], line_39[138], line_38[136], line_37[134], line_36[132], line_35[130], line_34[128], line_33[126], line_32[124], line_31[122], line_30[120], line_29[118], line_28[116], line_27[114], line_26[112], line_25[110], line_24[108], line_23[106], line_22[104], line_21[102], line_20[100], line_19[98], line_18[96], line_17[94], line_16[92], line_15[90], line_14[88], line_13[86], line_12[84], line_11[82], line_10[80], line_9[78], line_8[76], line_7[74], line_6[72], line_5[70], line_4[68], line_3[66], line_2[64], line_1[62] };
assign col_317 = {line_128[317], line_127[315], line_126[313], line_125[311], line_124[309], line_123[307], line_122[305], line_121[303], line_120[301], line_119[299], line_118[297], line_117[295], line_116[293], line_115[291], line_114[289], line_113[287], line_112[285], line_111[283], line_110[281], line_109[279], line_108[277], line_107[275], line_106[273], line_105[271], line_104[269], line_103[267], line_102[265], line_101[263], line_100[261], line_99[259], line_98[257], line_97[255], line_96[253], line_95[251], line_94[249], line_93[247], line_92[245], line_91[243], line_90[241], line_89[239], line_88[237], line_87[235], line_86[233], line_85[231], line_84[229], line_83[227], line_82[225], line_81[223], line_80[221], line_79[219], line_78[217], line_77[215], line_76[213], line_75[211], line_74[209], line_73[207], line_72[205], line_71[203], line_70[201], line_69[199], line_68[197], line_67[195], line_66[193], line_65[191], line_64[189], line_63[187], line_62[185], line_61[183], line_60[181], line_59[179], line_58[177], line_57[175], line_56[173], line_55[171], line_54[169], line_53[167], line_52[165], line_51[163], line_50[161], line_49[159], line_48[157], line_47[155], line_46[153], line_45[151], line_44[149], line_43[147], line_42[145], line_41[143], line_40[141], line_39[139], line_38[137], line_37[135], line_36[133], line_35[131], line_34[129], line_33[127], line_32[125], line_31[123], line_30[121], line_29[119], line_28[117], line_27[115], line_26[113], line_25[111], line_24[109], line_23[107], line_22[105], line_21[103], line_20[101], line_19[99], line_18[97], line_17[95], line_16[93], line_15[91], line_14[89], line_13[87], line_12[85], line_11[83], line_10[81], line_9[79], line_8[77], line_7[75], line_6[73], line_5[71], line_4[69], line_3[67], line_2[65], line_1[63] };
assign col_318 = {line_128[318], line_127[316], line_126[314], line_125[312], line_124[310], line_123[308], line_122[306], line_121[304], line_120[302], line_119[300], line_118[298], line_117[296], line_116[294], line_115[292], line_114[290], line_113[288], line_112[286], line_111[284], line_110[282], line_109[280], line_108[278], line_107[276], line_106[274], line_105[272], line_104[270], line_103[268], line_102[266], line_101[264], line_100[262], line_99[260], line_98[258], line_97[256], line_96[254], line_95[252], line_94[250], line_93[248], line_92[246], line_91[244], line_90[242], line_89[240], line_88[238], line_87[236], line_86[234], line_85[232], line_84[230], line_83[228], line_82[226], line_81[224], line_80[222], line_79[220], line_78[218], line_77[216], line_76[214], line_75[212], line_74[210], line_73[208], line_72[206], line_71[204], line_70[202], line_69[200], line_68[198], line_67[196], line_66[194], line_65[192], line_64[190], line_63[188], line_62[186], line_61[184], line_60[182], line_59[180], line_58[178], line_57[176], line_56[174], line_55[172], line_54[170], line_53[168], line_52[166], line_51[164], line_50[162], line_49[160], line_48[158], line_47[156], line_46[154], line_45[152], line_44[150], line_43[148], line_42[146], line_41[144], line_40[142], line_39[140], line_38[138], line_37[136], line_36[134], line_35[132], line_34[130], line_33[128], line_32[126], line_31[124], line_30[122], line_29[120], line_28[118], line_27[116], line_26[114], line_25[112], line_24[110], line_23[108], line_22[106], line_21[104], line_20[102], line_19[100], line_18[98], line_17[96], line_16[94], line_15[92], line_14[90], line_13[88], line_12[86], line_11[84], line_10[82], line_9[80], line_8[78], line_7[76], line_6[74], line_5[72], line_4[70], line_3[68], line_2[66], line_1[64] };
assign col_319 = {line_128[319], line_127[317], line_126[315], line_125[313], line_124[311], line_123[309], line_122[307], line_121[305], line_120[303], line_119[301], line_118[299], line_117[297], line_116[295], line_115[293], line_114[291], line_113[289], line_112[287], line_111[285], line_110[283], line_109[281], line_108[279], line_107[277], line_106[275], line_105[273], line_104[271], line_103[269], line_102[267], line_101[265], line_100[263], line_99[261], line_98[259], line_97[257], line_96[255], line_95[253], line_94[251], line_93[249], line_92[247], line_91[245], line_90[243], line_89[241], line_88[239], line_87[237], line_86[235], line_85[233], line_84[231], line_83[229], line_82[227], line_81[225], line_80[223], line_79[221], line_78[219], line_77[217], line_76[215], line_75[213], line_74[211], line_73[209], line_72[207], line_71[205], line_70[203], line_69[201], line_68[199], line_67[197], line_66[195], line_65[193], line_64[191], line_63[189], line_62[187], line_61[185], line_60[183], line_59[181], line_58[179], line_57[177], line_56[175], line_55[173], line_54[171], line_53[169], line_52[167], line_51[165], line_50[163], line_49[161], line_48[159], line_47[157], line_46[155], line_45[153], line_44[151], line_43[149], line_42[147], line_41[145], line_40[143], line_39[141], line_38[139], line_37[137], line_36[135], line_35[133], line_34[131], line_33[129], line_32[127], line_31[125], line_30[123], line_29[121], line_28[119], line_27[117], line_26[115], line_25[113], line_24[111], line_23[109], line_22[107], line_21[105], line_20[103], line_19[101], line_18[99], line_17[97], line_16[95], line_15[93], line_14[91], line_13[89], line_12[87], line_11[85], line_10[83], line_9[81], line_8[79], line_7[77], line_6[75], line_5[73], line_4[71], line_3[69], line_2[67], line_1[65] };
assign col_320 = {line_128[320], line_127[318], line_126[316], line_125[314], line_124[312], line_123[310], line_122[308], line_121[306], line_120[304], line_119[302], line_118[300], line_117[298], line_116[296], line_115[294], line_114[292], line_113[290], line_112[288], line_111[286], line_110[284], line_109[282], line_108[280], line_107[278], line_106[276], line_105[274], line_104[272], line_103[270], line_102[268], line_101[266], line_100[264], line_99[262], line_98[260], line_97[258], line_96[256], line_95[254], line_94[252], line_93[250], line_92[248], line_91[246], line_90[244], line_89[242], line_88[240], line_87[238], line_86[236], line_85[234], line_84[232], line_83[230], line_82[228], line_81[226], line_80[224], line_79[222], line_78[220], line_77[218], line_76[216], line_75[214], line_74[212], line_73[210], line_72[208], line_71[206], line_70[204], line_69[202], line_68[200], line_67[198], line_66[196], line_65[194], line_64[192], line_63[190], line_62[188], line_61[186], line_60[184], line_59[182], line_58[180], line_57[178], line_56[176], line_55[174], line_54[172], line_53[170], line_52[168], line_51[166], line_50[164], line_49[162], line_48[160], line_47[158], line_46[156], line_45[154], line_44[152], line_43[150], line_42[148], line_41[146], line_40[144], line_39[142], line_38[140], line_37[138], line_36[136], line_35[134], line_34[132], line_33[130], line_32[128], line_31[126], line_30[124], line_29[122], line_28[120], line_27[118], line_26[116], line_25[114], line_24[112], line_23[110], line_22[108], line_21[106], line_20[104], line_19[102], line_18[100], line_17[98], line_16[96], line_15[94], line_14[92], line_13[90], line_12[88], line_11[86], line_10[84], line_9[82], line_8[80], line_7[78], line_6[76], line_5[74], line_4[72], line_3[70], line_2[68], line_1[66] };
assign col_321 = {line_128[321], line_127[319], line_126[317], line_125[315], line_124[313], line_123[311], line_122[309], line_121[307], line_120[305], line_119[303], line_118[301], line_117[299], line_116[297], line_115[295], line_114[293], line_113[291], line_112[289], line_111[287], line_110[285], line_109[283], line_108[281], line_107[279], line_106[277], line_105[275], line_104[273], line_103[271], line_102[269], line_101[267], line_100[265], line_99[263], line_98[261], line_97[259], line_96[257], line_95[255], line_94[253], line_93[251], line_92[249], line_91[247], line_90[245], line_89[243], line_88[241], line_87[239], line_86[237], line_85[235], line_84[233], line_83[231], line_82[229], line_81[227], line_80[225], line_79[223], line_78[221], line_77[219], line_76[217], line_75[215], line_74[213], line_73[211], line_72[209], line_71[207], line_70[205], line_69[203], line_68[201], line_67[199], line_66[197], line_65[195], line_64[193], line_63[191], line_62[189], line_61[187], line_60[185], line_59[183], line_58[181], line_57[179], line_56[177], line_55[175], line_54[173], line_53[171], line_52[169], line_51[167], line_50[165], line_49[163], line_48[161], line_47[159], line_46[157], line_45[155], line_44[153], line_43[151], line_42[149], line_41[147], line_40[145], line_39[143], line_38[141], line_37[139], line_36[137], line_35[135], line_34[133], line_33[131], line_32[129], line_31[127], line_30[125], line_29[123], line_28[121], line_27[119], line_26[117], line_25[115], line_24[113], line_23[111], line_22[109], line_21[107], line_20[105], line_19[103], line_18[101], line_17[99], line_16[97], line_15[95], line_14[93], line_13[91], line_12[89], line_11[87], line_10[85], line_9[83], line_8[81], line_7[79], line_6[77], line_5[75], line_4[73], line_3[71], line_2[69], line_1[67] };
assign col_322 = {line_128[322], line_127[320], line_126[318], line_125[316], line_124[314], line_123[312], line_122[310], line_121[308], line_120[306], line_119[304], line_118[302], line_117[300], line_116[298], line_115[296], line_114[294], line_113[292], line_112[290], line_111[288], line_110[286], line_109[284], line_108[282], line_107[280], line_106[278], line_105[276], line_104[274], line_103[272], line_102[270], line_101[268], line_100[266], line_99[264], line_98[262], line_97[260], line_96[258], line_95[256], line_94[254], line_93[252], line_92[250], line_91[248], line_90[246], line_89[244], line_88[242], line_87[240], line_86[238], line_85[236], line_84[234], line_83[232], line_82[230], line_81[228], line_80[226], line_79[224], line_78[222], line_77[220], line_76[218], line_75[216], line_74[214], line_73[212], line_72[210], line_71[208], line_70[206], line_69[204], line_68[202], line_67[200], line_66[198], line_65[196], line_64[194], line_63[192], line_62[190], line_61[188], line_60[186], line_59[184], line_58[182], line_57[180], line_56[178], line_55[176], line_54[174], line_53[172], line_52[170], line_51[168], line_50[166], line_49[164], line_48[162], line_47[160], line_46[158], line_45[156], line_44[154], line_43[152], line_42[150], line_41[148], line_40[146], line_39[144], line_38[142], line_37[140], line_36[138], line_35[136], line_34[134], line_33[132], line_32[130], line_31[128], line_30[126], line_29[124], line_28[122], line_27[120], line_26[118], line_25[116], line_24[114], line_23[112], line_22[110], line_21[108], line_20[106], line_19[104], line_18[102], line_17[100], line_16[98], line_15[96], line_14[94], line_13[92], line_12[90], line_11[88], line_10[86], line_9[84], line_8[82], line_7[80], line_6[78], line_5[76], line_4[74], line_3[72], line_2[70], line_1[68] };
assign col_323 = {line_128[323], line_127[321], line_126[319], line_125[317], line_124[315], line_123[313], line_122[311], line_121[309], line_120[307], line_119[305], line_118[303], line_117[301], line_116[299], line_115[297], line_114[295], line_113[293], line_112[291], line_111[289], line_110[287], line_109[285], line_108[283], line_107[281], line_106[279], line_105[277], line_104[275], line_103[273], line_102[271], line_101[269], line_100[267], line_99[265], line_98[263], line_97[261], line_96[259], line_95[257], line_94[255], line_93[253], line_92[251], line_91[249], line_90[247], line_89[245], line_88[243], line_87[241], line_86[239], line_85[237], line_84[235], line_83[233], line_82[231], line_81[229], line_80[227], line_79[225], line_78[223], line_77[221], line_76[219], line_75[217], line_74[215], line_73[213], line_72[211], line_71[209], line_70[207], line_69[205], line_68[203], line_67[201], line_66[199], line_65[197], line_64[195], line_63[193], line_62[191], line_61[189], line_60[187], line_59[185], line_58[183], line_57[181], line_56[179], line_55[177], line_54[175], line_53[173], line_52[171], line_51[169], line_50[167], line_49[165], line_48[163], line_47[161], line_46[159], line_45[157], line_44[155], line_43[153], line_42[151], line_41[149], line_40[147], line_39[145], line_38[143], line_37[141], line_36[139], line_35[137], line_34[135], line_33[133], line_32[131], line_31[129], line_30[127], line_29[125], line_28[123], line_27[121], line_26[119], line_25[117], line_24[115], line_23[113], line_22[111], line_21[109], line_20[107], line_19[105], line_18[103], line_17[101], line_16[99], line_15[97], line_14[95], line_13[93], line_12[91], line_11[89], line_10[87], line_9[85], line_8[83], line_7[81], line_6[79], line_5[77], line_4[75], line_3[73], line_2[71], line_1[69] };
assign col_324 = {line_128[324], line_127[322], line_126[320], line_125[318], line_124[316], line_123[314], line_122[312], line_121[310], line_120[308], line_119[306], line_118[304], line_117[302], line_116[300], line_115[298], line_114[296], line_113[294], line_112[292], line_111[290], line_110[288], line_109[286], line_108[284], line_107[282], line_106[280], line_105[278], line_104[276], line_103[274], line_102[272], line_101[270], line_100[268], line_99[266], line_98[264], line_97[262], line_96[260], line_95[258], line_94[256], line_93[254], line_92[252], line_91[250], line_90[248], line_89[246], line_88[244], line_87[242], line_86[240], line_85[238], line_84[236], line_83[234], line_82[232], line_81[230], line_80[228], line_79[226], line_78[224], line_77[222], line_76[220], line_75[218], line_74[216], line_73[214], line_72[212], line_71[210], line_70[208], line_69[206], line_68[204], line_67[202], line_66[200], line_65[198], line_64[196], line_63[194], line_62[192], line_61[190], line_60[188], line_59[186], line_58[184], line_57[182], line_56[180], line_55[178], line_54[176], line_53[174], line_52[172], line_51[170], line_50[168], line_49[166], line_48[164], line_47[162], line_46[160], line_45[158], line_44[156], line_43[154], line_42[152], line_41[150], line_40[148], line_39[146], line_38[144], line_37[142], line_36[140], line_35[138], line_34[136], line_33[134], line_32[132], line_31[130], line_30[128], line_29[126], line_28[124], line_27[122], line_26[120], line_25[118], line_24[116], line_23[114], line_22[112], line_21[110], line_20[108], line_19[106], line_18[104], line_17[102], line_16[100], line_15[98], line_14[96], line_13[94], line_12[92], line_11[90], line_10[88], line_9[86], line_8[84], line_7[82], line_6[80], line_5[78], line_4[76], line_3[74], line_2[72], line_1[70] };
assign col_325 = {line_128[325], line_127[323], line_126[321], line_125[319], line_124[317], line_123[315], line_122[313], line_121[311], line_120[309], line_119[307], line_118[305], line_117[303], line_116[301], line_115[299], line_114[297], line_113[295], line_112[293], line_111[291], line_110[289], line_109[287], line_108[285], line_107[283], line_106[281], line_105[279], line_104[277], line_103[275], line_102[273], line_101[271], line_100[269], line_99[267], line_98[265], line_97[263], line_96[261], line_95[259], line_94[257], line_93[255], line_92[253], line_91[251], line_90[249], line_89[247], line_88[245], line_87[243], line_86[241], line_85[239], line_84[237], line_83[235], line_82[233], line_81[231], line_80[229], line_79[227], line_78[225], line_77[223], line_76[221], line_75[219], line_74[217], line_73[215], line_72[213], line_71[211], line_70[209], line_69[207], line_68[205], line_67[203], line_66[201], line_65[199], line_64[197], line_63[195], line_62[193], line_61[191], line_60[189], line_59[187], line_58[185], line_57[183], line_56[181], line_55[179], line_54[177], line_53[175], line_52[173], line_51[171], line_50[169], line_49[167], line_48[165], line_47[163], line_46[161], line_45[159], line_44[157], line_43[155], line_42[153], line_41[151], line_40[149], line_39[147], line_38[145], line_37[143], line_36[141], line_35[139], line_34[137], line_33[135], line_32[133], line_31[131], line_30[129], line_29[127], line_28[125], line_27[123], line_26[121], line_25[119], line_24[117], line_23[115], line_22[113], line_21[111], line_20[109], line_19[107], line_18[105], line_17[103], line_16[101], line_15[99], line_14[97], line_13[95], line_12[93], line_11[91], line_10[89], line_9[87], line_8[85], line_7[83], line_6[81], line_5[79], line_4[77], line_3[75], line_2[73], line_1[71] };
assign col_326 = {line_128[326], line_127[324], line_126[322], line_125[320], line_124[318], line_123[316], line_122[314], line_121[312], line_120[310], line_119[308], line_118[306], line_117[304], line_116[302], line_115[300], line_114[298], line_113[296], line_112[294], line_111[292], line_110[290], line_109[288], line_108[286], line_107[284], line_106[282], line_105[280], line_104[278], line_103[276], line_102[274], line_101[272], line_100[270], line_99[268], line_98[266], line_97[264], line_96[262], line_95[260], line_94[258], line_93[256], line_92[254], line_91[252], line_90[250], line_89[248], line_88[246], line_87[244], line_86[242], line_85[240], line_84[238], line_83[236], line_82[234], line_81[232], line_80[230], line_79[228], line_78[226], line_77[224], line_76[222], line_75[220], line_74[218], line_73[216], line_72[214], line_71[212], line_70[210], line_69[208], line_68[206], line_67[204], line_66[202], line_65[200], line_64[198], line_63[196], line_62[194], line_61[192], line_60[190], line_59[188], line_58[186], line_57[184], line_56[182], line_55[180], line_54[178], line_53[176], line_52[174], line_51[172], line_50[170], line_49[168], line_48[166], line_47[164], line_46[162], line_45[160], line_44[158], line_43[156], line_42[154], line_41[152], line_40[150], line_39[148], line_38[146], line_37[144], line_36[142], line_35[140], line_34[138], line_33[136], line_32[134], line_31[132], line_30[130], line_29[128], line_28[126], line_27[124], line_26[122], line_25[120], line_24[118], line_23[116], line_22[114], line_21[112], line_20[110], line_19[108], line_18[106], line_17[104], line_16[102], line_15[100], line_14[98], line_13[96], line_12[94], line_11[92], line_10[90], line_9[88], line_8[86], line_7[84], line_6[82], line_5[80], line_4[78], line_3[76], line_2[74], line_1[72] };
assign col_327 = {line_128[327], line_127[325], line_126[323], line_125[321], line_124[319], line_123[317], line_122[315], line_121[313], line_120[311], line_119[309], line_118[307], line_117[305], line_116[303], line_115[301], line_114[299], line_113[297], line_112[295], line_111[293], line_110[291], line_109[289], line_108[287], line_107[285], line_106[283], line_105[281], line_104[279], line_103[277], line_102[275], line_101[273], line_100[271], line_99[269], line_98[267], line_97[265], line_96[263], line_95[261], line_94[259], line_93[257], line_92[255], line_91[253], line_90[251], line_89[249], line_88[247], line_87[245], line_86[243], line_85[241], line_84[239], line_83[237], line_82[235], line_81[233], line_80[231], line_79[229], line_78[227], line_77[225], line_76[223], line_75[221], line_74[219], line_73[217], line_72[215], line_71[213], line_70[211], line_69[209], line_68[207], line_67[205], line_66[203], line_65[201], line_64[199], line_63[197], line_62[195], line_61[193], line_60[191], line_59[189], line_58[187], line_57[185], line_56[183], line_55[181], line_54[179], line_53[177], line_52[175], line_51[173], line_50[171], line_49[169], line_48[167], line_47[165], line_46[163], line_45[161], line_44[159], line_43[157], line_42[155], line_41[153], line_40[151], line_39[149], line_38[147], line_37[145], line_36[143], line_35[141], line_34[139], line_33[137], line_32[135], line_31[133], line_30[131], line_29[129], line_28[127], line_27[125], line_26[123], line_25[121], line_24[119], line_23[117], line_22[115], line_21[113], line_20[111], line_19[109], line_18[107], line_17[105], line_16[103], line_15[101], line_14[99], line_13[97], line_12[95], line_11[93], line_10[91], line_9[89], line_8[87], line_7[85], line_6[83], line_5[81], line_4[79], line_3[77], line_2[75], line_1[73] };
assign col_328 = {line_128[328], line_127[326], line_126[324], line_125[322], line_124[320], line_123[318], line_122[316], line_121[314], line_120[312], line_119[310], line_118[308], line_117[306], line_116[304], line_115[302], line_114[300], line_113[298], line_112[296], line_111[294], line_110[292], line_109[290], line_108[288], line_107[286], line_106[284], line_105[282], line_104[280], line_103[278], line_102[276], line_101[274], line_100[272], line_99[270], line_98[268], line_97[266], line_96[264], line_95[262], line_94[260], line_93[258], line_92[256], line_91[254], line_90[252], line_89[250], line_88[248], line_87[246], line_86[244], line_85[242], line_84[240], line_83[238], line_82[236], line_81[234], line_80[232], line_79[230], line_78[228], line_77[226], line_76[224], line_75[222], line_74[220], line_73[218], line_72[216], line_71[214], line_70[212], line_69[210], line_68[208], line_67[206], line_66[204], line_65[202], line_64[200], line_63[198], line_62[196], line_61[194], line_60[192], line_59[190], line_58[188], line_57[186], line_56[184], line_55[182], line_54[180], line_53[178], line_52[176], line_51[174], line_50[172], line_49[170], line_48[168], line_47[166], line_46[164], line_45[162], line_44[160], line_43[158], line_42[156], line_41[154], line_40[152], line_39[150], line_38[148], line_37[146], line_36[144], line_35[142], line_34[140], line_33[138], line_32[136], line_31[134], line_30[132], line_29[130], line_28[128], line_27[126], line_26[124], line_25[122], line_24[120], line_23[118], line_22[116], line_21[114], line_20[112], line_19[110], line_18[108], line_17[106], line_16[104], line_15[102], line_14[100], line_13[98], line_12[96], line_11[94], line_10[92], line_9[90], line_8[88], line_7[86], line_6[84], line_5[82], line_4[80], line_3[78], line_2[76], line_1[74] };
assign col_329 = {line_128[329], line_127[327], line_126[325], line_125[323], line_124[321], line_123[319], line_122[317], line_121[315], line_120[313], line_119[311], line_118[309], line_117[307], line_116[305], line_115[303], line_114[301], line_113[299], line_112[297], line_111[295], line_110[293], line_109[291], line_108[289], line_107[287], line_106[285], line_105[283], line_104[281], line_103[279], line_102[277], line_101[275], line_100[273], line_99[271], line_98[269], line_97[267], line_96[265], line_95[263], line_94[261], line_93[259], line_92[257], line_91[255], line_90[253], line_89[251], line_88[249], line_87[247], line_86[245], line_85[243], line_84[241], line_83[239], line_82[237], line_81[235], line_80[233], line_79[231], line_78[229], line_77[227], line_76[225], line_75[223], line_74[221], line_73[219], line_72[217], line_71[215], line_70[213], line_69[211], line_68[209], line_67[207], line_66[205], line_65[203], line_64[201], line_63[199], line_62[197], line_61[195], line_60[193], line_59[191], line_58[189], line_57[187], line_56[185], line_55[183], line_54[181], line_53[179], line_52[177], line_51[175], line_50[173], line_49[171], line_48[169], line_47[167], line_46[165], line_45[163], line_44[161], line_43[159], line_42[157], line_41[155], line_40[153], line_39[151], line_38[149], line_37[147], line_36[145], line_35[143], line_34[141], line_33[139], line_32[137], line_31[135], line_30[133], line_29[131], line_28[129], line_27[127], line_26[125], line_25[123], line_24[121], line_23[119], line_22[117], line_21[115], line_20[113], line_19[111], line_18[109], line_17[107], line_16[105], line_15[103], line_14[101], line_13[99], line_12[97], line_11[95], line_10[93], line_9[91], line_8[89], line_7[87], line_6[85], line_5[83], line_4[81], line_3[79], line_2[77], line_1[75] };
assign col_330 = {line_128[330], line_127[328], line_126[326], line_125[324], line_124[322], line_123[320], line_122[318], line_121[316], line_120[314], line_119[312], line_118[310], line_117[308], line_116[306], line_115[304], line_114[302], line_113[300], line_112[298], line_111[296], line_110[294], line_109[292], line_108[290], line_107[288], line_106[286], line_105[284], line_104[282], line_103[280], line_102[278], line_101[276], line_100[274], line_99[272], line_98[270], line_97[268], line_96[266], line_95[264], line_94[262], line_93[260], line_92[258], line_91[256], line_90[254], line_89[252], line_88[250], line_87[248], line_86[246], line_85[244], line_84[242], line_83[240], line_82[238], line_81[236], line_80[234], line_79[232], line_78[230], line_77[228], line_76[226], line_75[224], line_74[222], line_73[220], line_72[218], line_71[216], line_70[214], line_69[212], line_68[210], line_67[208], line_66[206], line_65[204], line_64[202], line_63[200], line_62[198], line_61[196], line_60[194], line_59[192], line_58[190], line_57[188], line_56[186], line_55[184], line_54[182], line_53[180], line_52[178], line_51[176], line_50[174], line_49[172], line_48[170], line_47[168], line_46[166], line_45[164], line_44[162], line_43[160], line_42[158], line_41[156], line_40[154], line_39[152], line_38[150], line_37[148], line_36[146], line_35[144], line_34[142], line_33[140], line_32[138], line_31[136], line_30[134], line_29[132], line_28[130], line_27[128], line_26[126], line_25[124], line_24[122], line_23[120], line_22[118], line_21[116], line_20[114], line_19[112], line_18[110], line_17[108], line_16[106], line_15[104], line_14[102], line_13[100], line_12[98], line_11[96], line_10[94], line_9[92], line_8[90], line_7[88], line_6[86], line_5[84], line_4[82], line_3[80], line_2[78], line_1[76] };
assign col_331 = {line_128[331], line_127[329], line_126[327], line_125[325], line_124[323], line_123[321], line_122[319], line_121[317], line_120[315], line_119[313], line_118[311], line_117[309], line_116[307], line_115[305], line_114[303], line_113[301], line_112[299], line_111[297], line_110[295], line_109[293], line_108[291], line_107[289], line_106[287], line_105[285], line_104[283], line_103[281], line_102[279], line_101[277], line_100[275], line_99[273], line_98[271], line_97[269], line_96[267], line_95[265], line_94[263], line_93[261], line_92[259], line_91[257], line_90[255], line_89[253], line_88[251], line_87[249], line_86[247], line_85[245], line_84[243], line_83[241], line_82[239], line_81[237], line_80[235], line_79[233], line_78[231], line_77[229], line_76[227], line_75[225], line_74[223], line_73[221], line_72[219], line_71[217], line_70[215], line_69[213], line_68[211], line_67[209], line_66[207], line_65[205], line_64[203], line_63[201], line_62[199], line_61[197], line_60[195], line_59[193], line_58[191], line_57[189], line_56[187], line_55[185], line_54[183], line_53[181], line_52[179], line_51[177], line_50[175], line_49[173], line_48[171], line_47[169], line_46[167], line_45[165], line_44[163], line_43[161], line_42[159], line_41[157], line_40[155], line_39[153], line_38[151], line_37[149], line_36[147], line_35[145], line_34[143], line_33[141], line_32[139], line_31[137], line_30[135], line_29[133], line_28[131], line_27[129], line_26[127], line_25[125], line_24[123], line_23[121], line_22[119], line_21[117], line_20[115], line_19[113], line_18[111], line_17[109], line_16[107], line_15[105], line_14[103], line_13[101], line_12[99], line_11[97], line_10[95], line_9[93], line_8[91], line_7[89], line_6[87], line_5[85], line_4[83], line_3[81], line_2[79], line_1[77] };
assign col_332 = {line_128[332], line_127[330], line_126[328], line_125[326], line_124[324], line_123[322], line_122[320], line_121[318], line_120[316], line_119[314], line_118[312], line_117[310], line_116[308], line_115[306], line_114[304], line_113[302], line_112[300], line_111[298], line_110[296], line_109[294], line_108[292], line_107[290], line_106[288], line_105[286], line_104[284], line_103[282], line_102[280], line_101[278], line_100[276], line_99[274], line_98[272], line_97[270], line_96[268], line_95[266], line_94[264], line_93[262], line_92[260], line_91[258], line_90[256], line_89[254], line_88[252], line_87[250], line_86[248], line_85[246], line_84[244], line_83[242], line_82[240], line_81[238], line_80[236], line_79[234], line_78[232], line_77[230], line_76[228], line_75[226], line_74[224], line_73[222], line_72[220], line_71[218], line_70[216], line_69[214], line_68[212], line_67[210], line_66[208], line_65[206], line_64[204], line_63[202], line_62[200], line_61[198], line_60[196], line_59[194], line_58[192], line_57[190], line_56[188], line_55[186], line_54[184], line_53[182], line_52[180], line_51[178], line_50[176], line_49[174], line_48[172], line_47[170], line_46[168], line_45[166], line_44[164], line_43[162], line_42[160], line_41[158], line_40[156], line_39[154], line_38[152], line_37[150], line_36[148], line_35[146], line_34[144], line_33[142], line_32[140], line_31[138], line_30[136], line_29[134], line_28[132], line_27[130], line_26[128], line_25[126], line_24[124], line_23[122], line_22[120], line_21[118], line_20[116], line_19[114], line_18[112], line_17[110], line_16[108], line_15[106], line_14[104], line_13[102], line_12[100], line_11[98], line_10[96], line_9[94], line_8[92], line_7[90], line_6[88], line_5[86], line_4[84], line_3[82], line_2[80], line_1[78] };
assign col_333 = {line_128[333], line_127[331], line_126[329], line_125[327], line_124[325], line_123[323], line_122[321], line_121[319], line_120[317], line_119[315], line_118[313], line_117[311], line_116[309], line_115[307], line_114[305], line_113[303], line_112[301], line_111[299], line_110[297], line_109[295], line_108[293], line_107[291], line_106[289], line_105[287], line_104[285], line_103[283], line_102[281], line_101[279], line_100[277], line_99[275], line_98[273], line_97[271], line_96[269], line_95[267], line_94[265], line_93[263], line_92[261], line_91[259], line_90[257], line_89[255], line_88[253], line_87[251], line_86[249], line_85[247], line_84[245], line_83[243], line_82[241], line_81[239], line_80[237], line_79[235], line_78[233], line_77[231], line_76[229], line_75[227], line_74[225], line_73[223], line_72[221], line_71[219], line_70[217], line_69[215], line_68[213], line_67[211], line_66[209], line_65[207], line_64[205], line_63[203], line_62[201], line_61[199], line_60[197], line_59[195], line_58[193], line_57[191], line_56[189], line_55[187], line_54[185], line_53[183], line_52[181], line_51[179], line_50[177], line_49[175], line_48[173], line_47[171], line_46[169], line_45[167], line_44[165], line_43[163], line_42[161], line_41[159], line_40[157], line_39[155], line_38[153], line_37[151], line_36[149], line_35[147], line_34[145], line_33[143], line_32[141], line_31[139], line_30[137], line_29[135], line_28[133], line_27[131], line_26[129], line_25[127], line_24[125], line_23[123], line_22[121], line_21[119], line_20[117], line_19[115], line_18[113], line_17[111], line_16[109], line_15[107], line_14[105], line_13[103], line_12[101], line_11[99], line_10[97], line_9[95], line_8[93], line_7[91], line_6[89], line_5[87], line_4[85], line_3[83], line_2[81], line_1[79] };
assign col_334 = {line_128[334], line_127[332], line_126[330], line_125[328], line_124[326], line_123[324], line_122[322], line_121[320], line_120[318], line_119[316], line_118[314], line_117[312], line_116[310], line_115[308], line_114[306], line_113[304], line_112[302], line_111[300], line_110[298], line_109[296], line_108[294], line_107[292], line_106[290], line_105[288], line_104[286], line_103[284], line_102[282], line_101[280], line_100[278], line_99[276], line_98[274], line_97[272], line_96[270], line_95[268], line_94[266], line_93[264], line_92[262], line_91[260], line_90[258], line_89[256], line_88[254], line_87[252], line_86[250], line_85[248], line_84[246], line_83[244], line_82[242], line_81[240], line_80[238], line_79[236], line_78[234], line_77[232], line_76[230], line_75[228], line_74[226], line_73[224], line_72[222], line_71[220], line_70[218], line_69[216], line_68[214], line_67[212], line_66[210], line_65[208], line_64[206], line_63[204], line_62[202], line_61[200], line_60[198], line_59[196], line_58[194], line_57[192], line_56[190], line_55[188], line_54[186], line_53[184], line_52[182], line_51[180], line_50[178], line_49[176], line_48[174], line_47[172], line_46[170], line_45[168], line_44[166], line_43[164], line_42[162], line_41[160], line_40[158], line_39[156], line_38[154], line_37[152], line_36[150], line_35[148], line_34[146], line_33[144], line_32[142], line_31[140], line_30[138], line_29[136], line_28[134], line_27[132], line_26[130], line_25[128], line_24[126], line_23[124], line_22[122], line_21[120], line_20[118], line_19[116], line_18[114], line_17[112], line_16[110], line_15[108], line_14[106], line_13[104], line_12[102], line_11[100], line_10[98], line_9[96], line_8[94], line_7[92], line_6[90], line_5[88], line_4[86], line_3[84], line_2[82], line_1[80] };
assign col_335 = {line_128[335], line_127[333], line_126[331], line_125[329], line_124[327], line_123[325], line_122[323], line_121[321], line_120[319], line_119[317], line_118[315], line_117[313], line_116[311], line_115[309], line_114[307], line_113[305], line_112[303], line_111[301], line_110[299], line_109[297], line_108[295], line_107[293], line_106[291], line_105[289], line_104[287], line_103[285], line_102[283], line_101[281], line_100[279], line_99[277], line_98[275], line_97[273], line_96[271], line_95[269], line_94[267], line_93[265], line_92[263], line_91[261], line_90[259], line_89[257], line_88[255], line_87[253], line_86[251], line_85[249], line_84[247], line_83[245], line_82[243], line_81[241], line_80[239], line_79[237], line_78[235], line_77[233], line_76[231], line_75[229], line_74[227], line_73[225], line_72[223], line_71[221], line_70[219], line_69[217], line_68[215], line_67[213], line_66[211], line_65[209], line_64[207], line_63[205], line_62[203], line_61[201], line_60[199], line_59[197], line_58[195], line_57[193], line_56[191], line_55[189], line_54[187], line_53[185], line_52[183], line_51[181], line_50[179], line_49[177], line_48[175], line_47[173], line_46[171], line_45[169], line_44[167], line_43[165], line_42[163], line_41[161], line_40[159], line_39[157], line_38[155], line_37[153], line_36[151], line_35[149], line_34[147], line_33[145], line_32[143], line_31[141], line_30[139], line_29[137], line_28[135], line_27[133], line_26[131], line_25[129], line_24[127], line_23[125], line_22[123], line_21[121], line_20[119], line_19[117], line_18[115], line_17[113], line_16[111], line_15[109], line_14[107], line_13[105], line_12[103], line_11[101], line_10[99], line_9[97], line_8[95], line_7[93], line_6[91], line_5[89], line_4[87], line_3[85], line_2[83], line_1[81] };
assign col_336 = {line_128[336], line_127[334], line_126[332], line_125[330], line_124[328], line_123[326], line_122[324], line_121[322], line_120[320], line_119[318], line_118[316], line_117[314], line_116[312], line_115[310], line_114[308], line_113[306], line_112[304], line_111[302], line_110[300], line_109[298], line_108[296], line_107[294], line_106[292], line_105[290], line_104[288], line_103[286], line_102[284], line_101[282], line_100[280], line_99[278], line_98[276], line_97[274], line_96[272], line_95[270], line_94[268], line_93[266], line_92[264], line_91[262], line_90[260], line_89[258], line_88[256], line_87[254], line_86[252], line_85[250], line_84[248], line_83[246], line_82[244], line_81[242], line_80[240], line_79[238], line_78[236], line_77[234], line_76[232], line_75[230], line_74[228], line_73[226], line_72[224], line_71[222], line_70[220], line_69[218], line_68[216], line_67[214], line_66[212], line_65[210], line_64[208], line_63[206], line_62[204], line_61[202], line_60[200], line_59[198], line_58[196], line_57[194], line_56[192], line_55[190], line_54[188], line_53[186], line_52[184], line_51[182], line_50[180], line_49[178], line_48[176], line_47[174], line_46[172], line_45[170], line_44[168], line_43[166], line_42[164], line_41[162], line_40[160], line_39[158], line_38[156], line_37[154], line_36[152], line_35[150], line_34[148], line_33[146], line_32[144], line_31[142], line_30[140], line_29[138], line_28[136], line_27[134], line_26[132], line_25[130], line_24[128], line_23[126], line_22[124], line_21[122], line_20[120], line_19[118], line_18[116], line_17[114], line_16[112], line_15[110], line_14[108], line_13[106], line_12[104], line_11[102], line_10[100], line_9[98], line_8[96], line_7[94], line_6[92], line_5[90], line_4[88], line_3[86], line_2[84], line_1[82] };
assign col_337 = {line_128[337], line_127[335], line_126[333], line_125[331], line_124[329], line_123[327], line_122[325], line_121[323], line_120[321], line_119[319], line_118[317], line_117[315], line_116[313], line_115[311], line_114[309], line_113[307], line_112[305], line_111[303], line_110[301], line_109[299], line_108[297], line_107[295], line_106[293], line_105[291], line_104[289], line_103[287], line_102[285], line_101[283], line_100[281], line_99[279], line_98[277], line_97[275], line_96[273], line_95[271], line_94[269], line_93[267], line_92[265], line_91[263], line_90[261], line_89[259], line_88[257], line_87[255], line_86[253], line_85[251], line_84[249], line_83[247], line_82[245], line_81[243], line_80[241], line_79[239], line_78[237], line_77[235], line_76[233], line_75[231], line_74[229], line_73[227], line_72[225], line_71[223], line_70[221], line_69[219], line_68[217], line_67[215], line_66[213], line_65[211], line_64[209], line_63[207], line_62[205], line_61[203], line_60[201], line_59[199], line_58[197], line_57[195], line_56[193], line_55[191], line_54[189], line_53[187], line_52[185], line_51[183], line_50[181], line_49[179], line_48[177], line_47[175], line_46[173], line_45[171], line_44[169], line_43[167], line_42[165], line_41[163], line_40[161], line_39[159], line_38[157], line_37[155], line_36[153], line_35[151], line_34[149], line_33[147], line_32[145], line_31[143], line_30[141], line_29[139], line_28[137], line_27[135], line_26[133], line_25[131], line_24[129], line_23[127], line_22[125], line_21[123], line_20[121], line_19[119], line_18[117], line_17[115], line_16[113], line_15[111], line_14[109], line_13[107], line_12[105], line_11[103], line_10[101], line_9[99], line_8[97], line_7[95], line_6[93], line_5[91], line_4[89], line_3[87], line_2[85], line_1[83] };
assign col_338 = {line_128[338], line_127[336], line_126[334], line_125[332], line_124[330], line_123[328], line_122[326], line_121[324], line_120[322], line_119[320], line_118[318], line_117[316], line_116[314], line_115[312], line_114[310], line_113[308], line_112[306], line_111[304], line_110[302], line_109[300], line_108[298], line_107[296], line_106[294], line_105[292], line_104[290], line_103[288], line_102[286], line_101[284], line_100[282], line_99[280], line_98[278], line_97[276], line_96[274], line_95[272], line_94[270], line_93[268], line_92[266], line_91[264], line_90[262], line_89[260], line_88[258], line_87[256], line_86[254], line_85[252], line_84[250], line_83[248], line_82[246], line_81[244], line_80[242], line_79[240], line_78[238], line_77[236], line_76[234], line_75[232], line_74[230], line_73[228], line_72[226], line_71[224], line_70[222], line_69[220], line_68[218], line_67[216], line_66[214], line_65[212], line_64[210], line_63[208], line_62[206], line_61[204], line_60[202], line_59[200], line_58[198], line_57[196], line_56[194], line_55[192], line_54[190], line_53[188], line_52[186], line_51[184], line_50[182], line_49[180], line_48[178], line_47[176], line_46[174], line_45[172], line_44[170], line_43[168], line_42[166], line_41[164], line_40[162], line_39[160], line_38[158], line_37[156], line_36[154], line_35[152], line_34[150], line_33[148], line_32[146], line_31[144], line_30[142], line_29[140], line_28[138], line_27[136], line_26[134], line_25[132], line_24[130], line_23[128], line_22[126], line_21[124], line_20[122], line_19[120], line_18[118], line_17[116], line_16[114], line_15[112], line_14[110], line_13[108], line_12[106], line_11[104], line_10[102], line_9[100], line_8[98], line_7[96], line_6[94], line_5[92], line_4[90], line_3[88], line_2[86], line_1[84] };
assign col_339 = {line_128[339], line_127[337], line_126[335], line_125[333], line_124[331], line_123[329], line_122[327], line_121[325], line_120[323], line_119[321], line_118[319], line_117[317], line_116[315], line_115[313], line_114[311], line_113[309], line_112[307], line_111[305], line_110[303], line_109[301], line_108[299], line_107[297], line_106[295], line_105[293], line_104[291], line_103[289], line_102[287], line_101[285], line_100[283], line_99[281], line_98[279], line_97[277], line_96[275], line_95[273], line_94[271], line_93[269], line_92[267], line_91[265], line_90[263], line_89[261], line_88[259], line_87[257], line_86[255], line_85[253], line_84[251], line_83[249], line_82[247], line_81[245], line_80[243], line_79[241], line_78[239], line_77[237], line_76[235], line_75[233], line_74[231], line_73[229], line_72[227], line_71[225], line_70[223], line_69[221], line_68[219], line_67[217], line_66[215], line_65[213], line_64[211], line_63[209], line_62[207], line_61[205], line_60[203], line_59[201], line_58[199], line_57[197], line_56[195], line_55[193], line_54[191], line_53[189], line_52[187], line_51[185], line_50[183], line_49[181], line_48[179], line_47[177], line_46[175], line_45[173], line_44[171], line_43[169], line_42[167], line_41[165], line_40[163], line_39[161], line_38[159], line_37[157], line_36[155], line_35[153], line_34[151], line_33[149], line_32[147], line_31[145], line_30[143], line_29[141], line_28[139], line_27[137], line_26[135], line_25[133], line_24[131], line_23[129], line_22[127], line_21[125], line_20[123], line_19[121], line_18[119], line_17[117], line_16[115], line_15[113], line_14[111], line_13[109], line_12[107], line_11[105], line_10[103], line_9[101], line_8[99], line_7[97], line_6[95], line_5[93], line_4[91], line_3[89], line_2[87], line_1[85] };
assign col_340 = {line_128[340], line_127[338], line_126[336], line_125[334], line_124[332], line_123[330], line_122[328], line_121[326], line_120[324], line_119[322], line_118[320], line_117[318], line_116[316], line_115[314], line_114[312], line_113[310], line_112[308], line_111[306], line_110[304], line_109[302], line_108[300], line_107[298], line_106[296], line_105[294], line_104[292], line_103[290], line_102[288], line_101[286], line_100[284], line_99[282], line_98[280], line_97[278], line_96[276], line_95[274], line_94[272], line_93[270], line_92[268], line_91[266], line_90[264], line_89[262], line_88[260], line_87[258], line_86[256], line_85[254], line_84[252], line_83[250], line_82[248], line_81[246], line_80[244], line_79[242], line_78[240], line_77[238], line_76[236], line_75[234], line_74[232], line_73[230], line_72[228], line_71[226], line_70[224], line_69[222], line_68[220], line_67[218], line_66[216], line_65[214], line_64[212], line_63[210], line_62[208], line_61[206], line_60[204], line_59[202], line_58[200], line_57[198], line_56[196], line_55[194], line_54[192], line_53[190], line_52[188], line_51[186], line_50[184], line_49[182], line_48[180], line_47[178], line_46[176], line_45[174], line_44[172], line_43[170], line_42[168], line_41[166], line_40[164], line_39[162], line_38[160], line_37[158], line_36[156], line_35[154], line_34[152], line_33[150], line_32[148], line_31[146], line_30[144], line_29[142], line_28[140], line_27[138], line_26[136], line_25[134], line_24[132], line_23[130], line_22[128], line_21[126], line_20[124], line_19[122], line_18[120], line_17[118], line_16[116], line_15[114], line_14[112], line_13[110], line_12[108], line_11[106], line_10[104], line_9[102], line_8[100], line_7[98], line_6[96], line_5[94], line_4[92], line_3[90], line_2[88], line_1[86] };
assign col_341 = {line_128[341], line_127[339], line_126[337], line_125[335], line_124[333], line_123[331], line_122[329], line_121[327], line_120[325], line_119[323], line_118[321], line_117[319], line_116[317], line_115[315], line_114[313], line_113[311], line_112[309], line_111[307], line_110[305], line_109[303], line_108[301], line_107[299], line_106[297], line_105[295], line_104[293], line_103[291], line_102[289], line_101[287], line_100[285], line_99[283], line_98[281], line_97[279], line_96[277], line_95[275], line_94[273], line_93[271], line_92[269], line_91[267], line_90[265], line_89[263], line_88[261], line_87[259], line_86[257], line_85[255], line_84[253], line_83[251], line_82[249], line_81[247], line_80[245], line_79[243], line_78[241], line_77[239], line_76[237], line_75[235], line_74[233], line_73[231], line_72[229], line_71[227], line_70[225], line_69[223], line_68[221], line_67[219], line_66[217], line_65[215], line_64[213], line_63[211], line_62[209], line_61[207], line_60[205], line_59[203], line_58[201], line_57[199], line_56[197], line_55[195], line_54[193], line_53[191], line_52[189], line_51[187], line_50[185], line_49[183], line_48[181], line_47[179], line_46[177], line_45[175], line_44[173], line_43[171], line_42[169], line_41[167], line_40[165], line_39[163], line_38[161], line_37[159], line_36[157], line_35[155], line_34[153], line_33[151], line_32[149], line_31[147], line_30[145], line_29[143], line_28[141], line_27[139], line_26[137], line_25[135], line_24[133], line_23[131], line_22[129], line_21[127], line_20[125], line_19[123], line_18[121], line_17[119], line_16[117], line_15[115], line_14[113], line_13[111], line_12[109], line_11[107], line_10[105], line_9[103], line_8[101], line_7[99], line_6[97], line_5[95], line_4[93], line_3[91], line_2[89], line_1[87] };
assign col_342 = {line_128[342], line_127[340], line_126[338], line_125[336], line_124[334], line_123[332], line_122[330], line_121[328], line_120[326], line_119[324], line_118[322], line_117[320], line_116[318], line_115[316], line_114[314], line_113[312], line_112[310], line_111[308], line_110[306], line_109[304], line_108[302], line_107[300], line_106[298], line_105[296], line_104[294], line_103[292], line_102[290], line_101[288], line_100[286], line_99[284], line_98[282], line_97[280], line_96[278], line_95[276], line_94[274], line_93[272], line_92[270], line_91[268], line_90[266], line_89[264], line_88[262], line_87[260], line_86[258], line_85[256], line_84[254], line_83[252], line_82[250], line_81[248], line_80[246], line_79[244], line_78[242], line_77[240], line_76[238], line_75[236], line_74[234], line_73[232], line_72[230], line_71[228], line_70[226], line_69[224], line_68[222], line_67[220], line_66[218], line_65[216], line_64[214], line_63[212], line_62[210], line_61[208], line_60[206], line_59[204], line_58[202], line_57[200], line_56[198], line_55[196], line_54[194], line_53[192], line_52[190], line_51[188], line_50[186], line_49[184], line_48[182], line_47[180], line_46[178], line_45[176], line_44[174], line_43[172], line_42[170], line_41[168], line_40[166], line_39[164], line_38[162], line_37[160], line_36[158], line_35[156], line_34[154], line_33[152], line_32[150], line_31[148], line_30[146], line_29[144], line_28[142], line_27[140], line_26[138], line_25[136], line_24[134], line_23[132], line_22[130], line_21[128], line_20[126], line_19[124], line_18[122], line_17[120], line_16[118], line_15[116], line_14[114], line_13[112], line_12[110], line_11[108], line_10[106], line_9[104], line_8[102], line_7[100], line_6[98], line_5[96], line_4[94], line_3[92], line_2[90], line_1[88] };
assign col_343 = {line_128[343], line_127[341], line_126[339], line_125[337], line_124[335], line_123[333], line_122[331], line_121[329], line_120[327], line_119[325], line_118[323], line_117[321], line_116[319], line_115[317], line_114[315], line_113[313], line_112[311], line_111[309], line_110[307], line_109[305], line_108[303], line_107[301], line_106[299], line_105[297], line_104[295], line_103[293], line_102[291], line_101[289], line_100[287], line_99[285], line_98[283], line_97[281], line_96[279], line_95[277], line_94[275], line_93[273], line_92[271], line_91[269], line_90[267], line_89[265], line_88[263], line_87[261], line_86[259], line_85[257], line_84[255], line_83[253], line_82[251], line_81[249], line_80[247], line_79[245], line_78[243], line_77[241], line_76[239], line_75[237], line_74[235], line_73[233], line_72[231], line_71[229], line_70[227], line_69[225], line_68[223], line_67[221], line_66[219], line_65[217], line_64[215], line_63[213], line_62[211], line_61[209], line_60[207], line_59[205], line_58[203], line_57[201], line_56[199], line_55[197], line_54[195], line_53[193], line_52[191], line_51[189], line_50[187], line_49[185], line_48[183], line_47[181], line_46[179], line_45[177], line_44[175], line_43[173], line_42[171], line_41[169], line_40[167], line_39[165], line_38[163], line_37[161], line_36[159], line_35[157], line_34[155], line_33[153], line_32[151], line_31[149], line_30[147], line_29[145], line_28[143], line_27[141], line_26[139], line_25[137], line_24[135], line_23[133], line_22[131], line_21[129], line_20[127], line_19[125], line_18[123], line_17[121], line_16[119], line_15[117], line_14[115], line_13[113], line_12[111], line_11[109], line_10[107], line_9[105], line_8[103], line_7[101], line_6[99], line_5[97], line_4[95], line_3[93], line_2[91], line_1[89] };
assign col_344 = {line_128[344], line_127[342], line_126[340], line_125[338], line_124[336], line_123[334], line_122[332], line_121[330], line_120[328], line_119[326], line_118[324], line_117[322], line_116[320], line_115[318], line_114[316], line_113[314], line_112[312], line_111[310], line_110[308], line_109[306], line_108[304], line_107[302], line_106[300], line_105[298], line_104[296], line_103[294], line_102[292], line_101[290], line_100[288], line_99[286], line_98[284], line_97[282], line_96[280], line_95[278], line_94[276], line_93[274], line_92[272], line_91[270], line_90[268], line_89[266], line_88[264], line_87[262], line_86[260], line_85[258], line_84[256], line_83[254], line_82[252], line_81[250], line_80[248], line_79[246], line_78[244], line_77[242], line_76[240], line_75[238], line_74[236], line_73[234], line_72[232], line_71[230], line_70[228], line_69[226], line_68[224], line_67[222], line_66[220], line_65[218], line_64[216], line_63[214], line_62[212], line_61[210], line_60[208], line_59[206], line_58[204], line_57[202], line_56[200], line_55[198], line_54[196], line_53[194], line_52[192], line_51[190], line_50[188], line_49[186], line_48[184], line_47[182], line_46[180], line_45[178], line_44[176], line_43[174], line_42[172], line_41[170], line_40[168], line_39[166], line_38[164], line_37[162], line_36[160], line_35[158], line_34[156], line_33[154], line_32[152], line_31[150], line_30[148], line_29[146], line_28[144], line_27[142], line_26[140], line_25[138], line_24[136], line_23[134], line_22[132], line_21[130], line_20[128], line_19[126], line_18[124], line_17[122], line_16[120], line_15[118], line_14[116], line_13[114], line_12[112], line_11[110], line_10[108], line_9[106], line_8[104], line_7[102], line_6[100], line_5[98], line_4[96], line_3[94], line_2[92], line_1[90] };
assign col_345 = {line_128[345], line_127[343], line_126[341], line_125[339], line_124[337], line_123[335], line_122[333], line_121[331], line_120[329], line_119[327], line_118[325], line_117[323], line_116[321], line_115[319], line_114[317], line_113[315], line_112[313], line_111[311], line_110[309], line_109[307], line_108[305], line_107[303], line_106[301], line_105[299], line_104[297], line_103[295], line_102[293], line_101[291], line_100[289], line_99[287], line_98[285], line_97[283], line_96[281], line_95[279], line_94[277], line_93[275], line_92[273], line_91[271], line_90[269], line_89[267], line_88[265], line_87[263], line_86[261], line_85[259], line_84[257], line_83[255], line_82[253], line_81[251], line_80[249], line_79[247], line_78[245], line_77[243], line_76[241], line_75[239], line_74[237], line_73[235], line_72[233], line_71[231], line_70[229], line_69[227], line_68[225], line_67[223], line_66[221], line_65[219], line_64[217], line_63[215], line_62[213], line_61[211], line_60[209], line_59[207], line_58[205], line_57[203], line_56[201], line_55[199], line_54[197], line_53[195], line_52[193], line_51[191], line_50[189], line_49[187], line_48[185], line_47[183], line_46[181], line_45[179], line_44[177], line_43[175], line_42[173], line_41[171], line_40[169], line_39[167], line_38[165], line_37[163], line_36[161], line_35[159], line_34[157], line_33[155], line_32[153], line_31[151], line_30[149], line_29[147], line_28[145], line_27[143], line_26[141], line_25[139], line_24[137], line_23[135], line_22[133], line_21[131], line_20[129], line_19[127], line_18[125], line_17[123], line_16[121], line_15[119], line_14[117], line_13[115], line_12[113], line_11[111], line_10[109], line_9[107], line_8[105], line_7[103], line_6[101], line_5[99], line_4[97], line_3[95], line_2[93], line_1[91] };
assign col_346 = {line_128[346], line_127[344], line_126[342], line_125[340], line_124[338], line_123[336], line_122[334], line_121[332], line_120[330], line_119[328], line_118[326], line_117[324], line_116[322], line_115[320], line_114[318], line_113[316], line_112[314], line_111[312], line_110[310], line_109[308], line_108[306], line_107[304], line_106[302], line_105[300], line_104[298], line_103[296], line_102[294], line_101[292], line_100[290], line_99[288], line_98[286], line_97[284], line_96[282], line_95[280], line_94[278], line_93[276], line_92[274], line_91[272], line_90[270], line_89[268], line_88[266], line_87[264], line_86[262], line_85[260], line_84[258], line_83[256], line_82[254], line_81[252], line_80[250], line_79[248], line_78[246], line_77[244], line_76[242], line_75[240], line_74[238], line_73[236], line_72[234], line_71[232], line_70[230], line_69[228], line_68[226], line_67[224], line_66[222], line_65[220], line_64[218], line_63[216], line_62[214], line_61[212], line_60[210], line_59[208], line_58[206], line_57[204], line_56[202], line_55[200], line_54[198], line_53[196], line_52[194], line_51[192], line_50[190], line_49[188], line_48[186], line_47[184], line_46[182], line_45[180], line_44[178], line_43[176], line_42[174], line_41[172], line_40[170], line_39[168], line_38[166], line_37[164], line_36[162], line_35[160], line_34[158], line_33[156], line_32[154], line_31[152], line_30[150], line_29[148], line_28[146], line_27[144], line_26[142], line_25[140], line_24[138], line_23[136], line_22[134], line_21[132], line_20[130], line_19[128], line_18[126], line_17[124], line_16[122], line_15[120], line_14[118], line_13[116], line_12[114], line_11[112], line_10[110], line_9[108], line_8[106], line_7[104], line_6[102], line_5[100], line_4[98], line_3[96], line_2[94], line_1[92] };
assign col_347 = {line_128[347], line_127[345], line_126[343], line_125[341], line_124[339], line_123[337], line_122[335], line_121[333], line_120[331], line_119[329], line_118[327], line_117[325], line_116[323], line_115[321], line_114[319], line_113[317], line_112[315], line_111[313], line_110[311], line_109[309], line_108[307], line_107[305], line_106[303], line_105[301], line_104[299], line_103[297], line_102[295], line_101[293], line_100[291], line_99[289], line_98[287], line_97[285], line_96[283], line_95[281], line_94[279], line_93[277], line_92[275], line_91[273], line_90[271], line_89[269], line_88[267], line_87[265], line_86[263], line_85[261], line_84[259], line_83[257], line_82[255], line_81[253], line_80[251], line_79[249], line_78[247], line_77[245], line_76[243], line_75[241], line_74[239], line_73[237], line_72[235], line_71[233], line_70[231], line_69[229], line_68[227], line_67[225], line_66[223], line_65[221], line_64[219], line_63[217], line_62[215], line_61[213], line_60[211], line_59[209], line_58[207], line_57[205], line_56[203], line_55[201], line_54[199], line_53[197], line_52[195], line_51[193], line_50[191], line_49[189], line_48[187], line_47[185], line_46[183], line_45[181], line_44[179], line_43[177], line_42[175], line_41[173], line_40[171], line_39[169], line_38[167], line_37[165], line_36[163], line_35[161], line_34[159], line_33[157], line_32[155], line_31[153], line_30[151], line_29[149], line_28[147], line_27[145], line_26[143], line_25[141], line_24[139], line_23[137], line_22[135], line_21[133], line_20[131], line_19[129], line_18[127], line_17[125], line_16[123], line_15[121], line_14[119], line_13[117], line_12[115], line_11[113], line_10[111], line_9[109], line_8[107], line_7[105], line_6[103], line_5[101], line_4[99], line_3[97], line_2[95], line_1[93] };
assign col_348 = {line_128[348], line_127[346], line_126[344], line_125[342], line_124[340], line_123[338], line_122[336], line_121[334], line_120[332], line_119[330], line_118[328], line_117[326], line_116[324], line_115[322], line_114[320], line_113[318], line_112[316], line_111[314], line_110[312], line_109[310], line_108[308], line_107[306], line_106[304], line_105[302], line_104[300], line_103[298], line_102[296], line_101[294], line_100[292], line_99[290], line_98[288], line_97[286], line_96[284], line_95[282], line_94[280], line_93[278], line_92[276], line_91[274], line_90[272], line_89[270], line_88[268], line_87[266], line_86[264], line_85[262], line_84[260], line_83[258], line_82[256], line_81[254], line_80[252], line_79[250], line_78[248], line_77[246], line_76[244], line_75[242], line_74[240], line_73[238], line_72[236], line_71[234], line_70[232], line_69[230], line_68[228], line_67[226], line_66[224], line_65[222], line_64[220], line_63[218], line_62[216], line_61[214], line_60[212], line_59[210], line_58[208], line_57[206], line_56[204], line_55[202], line_54[200], line_53[198], line_52[196], line_51[194], line_50[192], line_49[190], line_48[188], line_47[186], line_46[184], line_45[182], line_44[180], line_43[178], line_42[176], line_41[174], line_40[172], line_39[170], line_38[168], line_37[166], line_36[164], line_35[162], line_34[160], line_33[158], line_32[156], line_31[154], line_30[152], line_29[150], line_28[148], line_27[146], line_26[144], line_25[142], line_24[140], line_23[138], line_22[136], line_21[134], line_20[132], line_19[130], line_18[128], line_17[126], line_16[124], line_15[122], line_14[120], line_13[118], line_12[116], line_11[114], line_10[112], line_9[110], line_8[108], line_7[106], line_6[104], line_5[102], line_4[100], line_3[98], line_2[96], line_1[94] };
assign col_349 = {line_128[349], line_127[347], line_126[345], line_125[343], line_124[341], line_123[339], line_122[337], line_121[335], line_120[333], line_119[331], line_118[329], line_117[327], line_116[325], line_115[323], line_114[321], line_113[319], line_112[317], line_111[315], line_110[313], line_109[311], line_108[309], line_107[307], line_106[305], line_105[303], line_104[301], line_103[299], line_102[297], line_101[295], line_100[293], line_99[291], line_98[289], line_97[287], line_96[285], line_95[283], line_94[281], line_93[279], line_92[277], line_91[275], line_90[273], line_89[271], line_88[269], line_87[267], line_86[265], line_85[263], line_84[261], line_83[259], line_82[257], line_81[255], line_80[253], line_79[251], line_78[249], line_77[247], line_76[245], line_75[243], line_74[241], line_73[239], line_72[237], line_71[235], line_70[233], line_69[231], line_68[229], line_67[227], line_66[225], line_65[223], line_64[221], line_63[219], line_62[217], line_61[215], line_60[213], line_59[211], line_58[209], line_57[207], line_56[205], line_55[203], line_54[201], line_53[199], line_52[197], line_51[195], line_50[193], line_49[191], line_48[189], line_47[187], line_46[185], line_45[183], line_44[181], line_43[179], line_42[177], line_41[175], line_40[173], line_39[171], line_38[169], line_37[167], line_36[165], line_35[163], line_34[161], line_33[159], line_32[157], line_31[155], line_30[153], line_29[151], line_28[149], line_27[147], line_26[145], line_25[143], line_24[141], line_23[139], line_22[137], line_21[135], line_20[133], line_19[131], line_18[129], line_17[127], line_16[125], line_15[123], line_14[121], line_13[119], line_12[117], line_11[115], line_10[113], line_9[111], line_8[109], line_7[107], line_6[105], line_5[103], line_4[101], line_3[99], line_2[97], line_1[95] };
assign col_350 = {line_128[350], line_127[348], line_126[346], line_125[344], line_124[342], line_123[340], line_122[338], line_121[336], line_120[334], line_119[332], line_118[330], line_117[328], line_116[326], line_115[324], line_114[322], line_113[320], line_112[318], line_111[316], line_110[314], line_109[312], line_108[310], line_107[308], line_106[306], line_105[304], line_104[302], line_103[300], line_102[298], line_101[296], line_100[294], line_99[292], line_98[290], line_97[288], line_96[286], line_95[284], line_94[282], line_93[280], line_92[278], line_91[276], line_90[274], line_89[272], line_88[270], line_87[268], line_86[266], line_85[264], line_84[262], line_83[260], line_82[258], line_81[256], line_80[254], line_79[252], line_78[250], line_77[248], line_76[246], line_75[244], line_74[242], line_73[240], line_72[238], line_71[236], line_70[234], line_69[232], line_68[230], line_67[228], line_66[226], line_65[224], line_64[222], line_63[220], line_62[218], line_61[216], line_60[214], line_59[212], line_58[210], line_57[208], line_56[206], line_55[204], line_54[202], line_53[200], line_52[198], line_51[196], line_50[194], line_49[192], line_48[190], line_47[188], line_46[186], line_45[184], line_44[182], line_43[180], line_42[178], line_41[176], line_40[174], line_39[172], line_38[170], line_37[168], line_36[166], line_35[164], line_34[162], line_33[160], line_32[158], line_31[156], line_30[154], line_29[152], line_28[150], line_27[148], line_26[146], line_25[144], line_24[142], line_23[140], line_22[138], line_21[136], line_20[134], line_19[132], line_18[130], line_17[128], line_16[126], line_15[124], line_14[122], line_13[120], line_12[118], line_11[116], line_10[114], line_9[112], line_8[110], line_7[108], line_6[106], line_5[104], line_4[102], line_3[100], line_2[98], line_1[96] };
assign col_351 = {line_128[351], line_127[349], line_126[347], line_125[345], line_124[343], line_123[341], line_122[339], line_121[337], line_120[335], line_119[333], line_118[331], line_117[329], line_116[327], line_115[325], line_114[323], line_113[321], line_112[319], line_111[317], line_110[315], line_109[313], line_108[311], line_107[309], line_106[307], line_105[305], line_104[303], line_103[301], line_102[299], line_101[297], line_100[295], line_99[293], line_98[291], line_97[289], line_96[287], line_95[285], line_94[283], line_93[281], line_92[279], line_91[277], line_90[275], line_89[273], line_88[271], line_87[269], line_86[267], line_85[265], line_84[263], line_83[261], line_82[259], line_81[257], line_80[255], line_79[253], line_78[251], line_77[249], line_76[247], line_75[245], line_74[243], line_73[241], line_72[239], line_71[237], line_70[235], line_69[233], line_68[231], line_67[229], line_66[227], line_65[225], line_64[223], line_63[221], line_62[219], line_61[217], line_60[215], line_59[213], line_58[211], line_57[209], line_56[207], line_55[205], line_54[203], line_53[201], line_52[199], line_51[197], line_50[195], line_49[193], line_48[191], line_47[189], line_46[187], line_45[185], line_44[183], line_43[181], line_42[179], line_41[177], line_40[175], line_39[173], line_38[171], line_37[169], line_36[167], line_35[165], line_34[163], line_33[161], line_32[159], line_31[157], line_30[155], line_29[153], line_28[151], line_27[149], line_26[147], line_25[145], line_24[143], line_23[141], line_22[139], line_21[137], line_20[135], line_19[133], line_18[131], line_17[129], line_16[127], line_15[125], line_14[123], line_13[121], line_12[119], line_11[117], line_10[115], line_9[113], line_8[111], line_7[109], line_6[107], line_5[105], line_4[103], line_3[101], line_2[99], line_1[97] };
assign col_352 = {line_128[352], line_127[350], line_126[348], line_125[346], line_124[344], line_123[342], line_122[340], line_121[338], line_120[336], line_119[334], line_118[332], line_117[330], line_116[328], line_115[326], line_114[324], line_113[322], line_112[320], line_111[318], line_110[316], line_109[314], line_108[312], line_107[310], line_106[308], line_105[306], line_104[304], line_103[302], line_102[300], line_101[298], line_100[296], line_99[294], line_98[292], line_97[290], line_96[288], line_95[286], line_94[284], line_93[282], line_92[280], line_91[278], line_90[276], line_89[274], line_88[272], line_87[270], line_86[268], line_85[266], line_84[264], line_83[262], line_82[260], line_81[258], line_80[256], line_79[254], line_78[252], line_77[250], line_76[248], line_75[246], line_74[244], line_73[242], line_72[240], line_71[238], line_70[236], line_69[234], line_68[232], line_67[230], line_66[228], line_65[226], line_64[224], line_63[222], line_62[220], line_61[218], line_60[216], line_59[214], line_58[212], line_57[210], line_56[208], line_55[206], line_54[204], line_53[202], line_52[200], line_51[198], line_50[196], line_49[194], line_48[192], line_47[190], line_46[188], line_45[186], line_44[184], line_43[182], line_42[180], line_41[178], line_40[176], line_39[174], line_38[172], line_37[170], line_36[168], line_35[166], line_34[164], line_33[162], line_32[160], line_31[158], line_30[156], line_29[154], line_28[152], line_27[150], line_26[148], line_25[146], line_24[144], line_23[142], line_22[140], line_21[138], line_20[136], line_19[134], line_18[132], line_17[130], line_16[128], line_15[126], line_14[124], line_13[122], line_12[120], line_11[118], line_10[116], line_9[114], line_8[112], line_7[110], line_6[108], line_5[106], line_4[104], line_3[102], line_2[100], line_1[98] };
assign col_353 = {line_128[353], line_127[351], line_126[349], line_125[347], line_124[345], line_123[343], line_122[341], line_121[339], line_120[337], line_119[335], line_118[333], line_117[331], line_116[329], line_115[327], line_114[325], line_113[323], line_112[321], line_111[319], line_110[317], line_109[315], line_108[313], line_107[311], line_106[309], line_105[307], line_104[305], line_103[303], line_102[301], line_101[299], line_100[297], line_99[295], line_98[293], line_97[291], line_96[289], line_95[287], line_94[285], line_93[283], line_92[281], line_91[279], line_90[277], line_89[275], line_88[273], line_87[271], line_86[269], line_85[267], line_84[265], line_83[263], line_82[261], line_81[259], line_80[257], line_79[255], line_78[253], line_77[251], line_76[249], line_75[247], line_74[245], line_73[243], line_72[241], line_71[239], line_70[237], line_69[235], line_68[233], line_67[231], line_66[229], line_65[227], line_64[225], line_63[223], line_62[221], line_61[219], line_60[217], line_59[215], line_58[213], line_57[211], line_56[209], line_55[207], line_54[205], line_53[203], line_52[201], line_51[199], line_50[197], line_49[195], line_48[193], line_47[191], line_46[189], line_45[187], line_44[185], line_43[183], line_42[181], line_41[179], line_40[177], line_39[175], line_38[173], line_37[171], line_36[169], line_35[167], line_34[165], line_33[163], line_32[161], line_31[159], line_30[157], line_29[155], line_28[153], line_27[151], line_26[149], line_25[147], line_24[145], line_23[143], line_22[141], line_21[139], line_20[137], line_19[135], line_18[133], line_17[131], line_16[129], line_15[127], line_14[125], line_13[123], line_12[121], line_11[119], line_10[117], line_9[115], line_8[113], line_7[111], line_6[109], line_5[107], line_4[105], line_3[103], line_2[101], line_1[99] };
assign col_354 = {line_128[354], line_127[352], line_126[350], line_125[348], line_124[346], line_123[344], line_122[342], line_121[340], line_120[338], line_119[336], line_118[334], line_117[332], line_116[330], line_115[328], line_114[326], line_113[324], line_112[322], line_111[320], line_110[318], line_109[316], line_108[314], line_107[312], line_106[310], line_105[308], line_104[306], line_103[304], line_102[302], line_101[300], line_100[298], line_99[296], line_98[294], line_97[292], line_96[290], line_95[288], line_94[286], line_93[284], line_92[282], line_91[280], line_90[278], line_89[276], line_88[274], line_87[272], line_86[270], line_85[268], line_84[266], line_83[264], line_82[262], line_81[260], line_80[258], line_79[256], line_78[254], line_77[252], line_76[250], line_75[248], line_74[246], line_73[244], line_72[242], line_71[240], line_70[238], line_69[236], line_68[234], line_67[232], line_66[230], line_65[228], line_64[226], line_63[224], line_62[222], line_61[220], line_60[218], line_59[216], line_58[214], line_57[212], line_56[210], line_55[208], line_54[206], line_53[204], line_52[202], line_51[200], line_50[198], line_49[196], line_48[194], line_47[192], line_46[190], line_45[188], line_44[186], line_43[184], line_42[182], line_41[180], line_40[178], line_39[176], line_38[174], line_37[172], line_36[170], line_35[168], line_34[166], line_33[164], line_32[162], line_31[160], line_30[158], line_29[156], line_28[154], line_27[152], line_26[150], line_25[148], line_24[146], line_23[144], line_22[142], line_21[140], line_20[138], line_19[136], line_18[134], line_17[132], line_16[130], line_15[128], line_14[126], line_13[124], line_12[122], line_11[120], line_10[118], line_9[116], line_8[114], line_7[112], line_6[110], line_5[108], line_4[106], line_3[104], line_2[102], line_1[100] };
assign col_355 = {line_128[355], line_127[353], line_126[351], line_125[349], line_124[347], line_123[345], line_122[343], line_121[341], line_120[339], line_119[337], line_118[335], line_117[333], line_116[331], line_115[329], line_114[327], line_113[325], line_112[323], line_111[321], line_110[319], line_109[317], line_108[315], line_107[313], line_106[311], line_105[309], line_104[307], line_103[305], line_102[303], line_101[301], line_100[299], line_99[297], line_98[295], line_97[293], line_96[291], line_95[289], line_94[287], line_93[285], line_92[283], line_91[281], line_90[279], line_89[277], line_88[275], line_87[273], line_86[271], line_85[269], line_84[267], line_83[265], line_82[263], line_81[261], line_80[259], line_79[257], line_78[255], line_77[253], line_76[251], line_75[249], line_74[247], line_73[245], line_72[243], line_71[241], line_70[239], line_69[237], line_68[235], line_67[233], line_66[231], line_65[229], line_64[227], line_63[225], line_62[223], line_61[221], line_60[219], line_59[217], line_58[215], line_57[213], line_56[211], line_55[209], line_54[207], line_53[205], line_52[203], line_51[201], line_50[199], line_49[197], line_48[195], line_47[193], line_46[191], line_45[189], line_44[187], line_43[185], line_42[183], line_41[181], line_40[179], line_39[177], line_38[175], line_37[173], line_36[171], line_35[169], line_34[167], line_33[165], line_32[163], line_31[161], line_30[159], line_29[157], line_28[155], line_27[153], line_26[151], line_25[149], line_24[147], line_23[145], line_22[143], line_21[141], line_20[139], line_19[137], line_18[135], line_17[133], line_16[131], line_15[129], line_14[127], line_13[125], line_12[123], line_11[121], line_10[119], line_9[117], line_8[115], line_7[113], line_6[111], line_5[109], line_4[107], line_3[105], line_2[103], line_1[101] };
assign col_356 = {line_128[356], line_127[354], line_126[352], line_125[350], line_124[348], line_123[346], line_122[344], line_121[342], line_120[340], line_119[338], line_118[336], line_117[334], line_116[332], line_115[330], line_114[328], line_113[326], line_112[324], line_111[322], line_110[320], line_109[318], line_108[316], line_107[314], line_106[312], line_105[310], line_104[308], line_103[306], line_102[304], line_101[302], line_100[300], line_99[298], line_98[296], line_97[294], line_96[292], line_95[290], line_94[288], line_93[286], line_92[284], line_91[282], line_90[280], line_89[278], line_88[276], line_87[274], line_86[272], line_85[270], line_84[268], line_83[266], line_82[264], line_81[262], line_80[260], line_79[258], line_78[256], line_77[254], line_76[252], line_75[250], line_74[248], line_73[246], line_72[244], line_71[242], line_70[240], line_69[238], line_68[236], line_67[234], line_66[232], line_65[230], line_64[228], line_63[226], line_62[224], line_61[222], line_60[220], line_59[218], line_58[216], line_57[214], line_56[212], line_55[210], line_54[208], line_53[206], line_52[204], line_51[202], line_50[200], line_49[198], line_48[196], line_47[194], line_46[192], line_45[190], line_44[188], line_43[186], line_42[184], line_41[182], line_40[180], line_39[178], line_38[176], line_37[174], line_36[172], line_35[170], line_34[168], line_33[166], line_32[164], line_31[162], line_30[160], line_29[158], line_28[156], line_27[154], line_26[152], line_25[150], line_24[148], line_23[146], line_22[144], line_21[142], line_20[140], line_19[138], line_18[136], line_17[134], line_16[132], line_15[130], line_14[128], line_13[126], line_12[124], line_11[122], line_10[120], line_9[118], line_8[116], line_7[114], line_6[112], line_5[110], line_4[108], line_3[106], line_2[104], line_1[102] };
assign col_357 = {line_128[357], line_127[355], line_126[353], line_125[351], line_124[349], line_123[347], line_122[345], line_121[343], line_120[341], line_119[339], line_118[337], line_117[335], line_116[333], line_115[331], line_114[329], line_113[327], line_112[325], line_111[323], line_110[321], line_109[319], line_108[317], line_107[315], line_106[313], line_105[311], line_104[309], line_103[307], line_102[305], line_101[303], line_100[301], line_99[299], line_98[297], line_97[295], line_96[293], line_95[291], line_94[289], line_93[287], line_92[285], line_91[283], line_90[281], line_89[279], line_88[277], line_87[275], line_86[273], line_85[271], line_84[269], line_83[267], line_82[265], line_81[263], line_80[261], line_79[259], line_78[257], line_77[255], line_76[253], line_75[251], line_74[249], line_73[247], line_72[245], line_71[243], line_70[241], line_69[239], line_68[237], line_67[235], line_66[233], line_65[231], line_64[229], line_63[227], line_62[225], line_61[223], line_60[221], line_59[219], line_58[217], line_57[215], line_56[213], line_55[211], line_54[209], line_53[207], line_52[205], line_51[203], line_50[201], line_49[199], line_48[197], line_47[195], line_46[193], line_45[191], line_44[189], line_43[187], line_42[185], line_41[183], line_40[181], line_39[179], line_38[177], line_37[175], line_36[173], line_35[171], line_34[169], line_33[167], line_32[165], line_31[163], line_30[161], line_29[159], line_28[157], line_27[155], line_26[153], line_25[151], line_24[149], line_23[147], line_22[145], line_21[143], line_20[141], line_19[139], line_18[137], line_17[135], line_16[133], line_15[131], line_14[129], line_13[127], line_12[125], line_11[123], line_10[121], line_9[119], line_8[117], line_7[115], line_6[113], line_5[111], line_4[109], line_3[107], line_2[105], line_1[103] };
assign col_358 = {line_128[358], line_127[356], line_126[354], line_125[352], line_124[350], line_123[348], line_122[346], line_121[344], line_120[342], line_119[340], line_118[338], line_117[336], line_116[334], line_115[332], line_114[330], line_113[328], line_112[326], line_111[324], line_110[322], line_109[320], line_108[318], line_107[316], line_106[314], line_105[312], line_104[310], line_103[308], line_102[306], line_101[304], line_100[302], line_99[300], line_98[298], line_97[296], line_96[294], line_95[292], line_94[290], line_93[288], line_92[286], line_91[284], line_90[282], line_89[280], line_88[278], line_87[276], line_86[274], line_85[272], line_84[270], line_83[268], line_82[266], line_81[264], line_80[262], line_79[260], line_78[258], line_77[256], line_76[254], line_75[252], line_74[250], line_73[248], line_72[246], line_71[244], line_70[242], line_69[240], line_68[238], line_67[236], line_66[234], line_65[232], line_64[230], line_63[228], line_62[226], line_61[224], line_60[222], line_59[220], line_58[218], line_57[216], line_56[214], line_55[212], line_54[210], line_53[208], line_52[206], line_51[204], line_50[202], line_49[200], line_48[198], line_47[196], line_46[194], line_45[192], line_44[190], line_43[188], line_42[186], line_41[184], line_40[182], line_39[180], line_38[178], line_37[176], line_36[174], line_35[172], line_34[170], line_33[168], line_32[166], line_31[164], line_30[162], line_29[160], line_28[158], line_27[156], line_26[154], line_25[152], line_24[150], line_23[148], line_22[146], line_21[144], line_20[142], line_19[140], line_18[138], line_17[136], line_16[134], line_15[132], line_14[130], line_13[128], line_12[126], line_11[124], line_10[122], line_9[120], line_8[118], line_7[116], line_6[114], line_5[112], line_4[110], line_3[108], line_2[106], line_1[104] };
assign col_359 = {line_128[359], line_127[357], line_126[355], line_125[353], line_124[351], line_123[349], line_122[347], line_121[345], line_120[343], line_119[341], line_118[339], line_117[337], line_116[335], line_115[333], line_114[331], line_113[329], line_112[327], line_111[325], line_110[323], line_109[321], line_108[319], line_107[317], line_106[315], line_105[313], line_104[311], line_103[309], line_102[307], line_101[305], line_100[303], line_99[301], line_98[299], line_97[297], line_96[295], line_95[293], line_94[291], line_93[289], line_92[287], line_91[285], line_90[283], line_89[281], line_88[279], line_87[277], line_86[275], line_85[273], line_84[271], line_83[269], line_82[267], line_81[265], line_80[263], line_79[261], line_78[259], line_77[257], line_76[255], line_75[253], line_74[251], line_73[249], line_72[247], line_71[245], line_70[243], line_69[241], line_68[239], line_67[237], line_66[235], line_65[233], line_64[231], line_63[229], line_62[227], line_61[225], line_60[223], line_59[221], line_58[219], line_57[217], line_56[215], line_55[213], line_54[211], line_53[209], line_52[207], line_51[205], line_50[203], line_49[201], line_48[199], line_47[197], line_46[195], line_45[193], line_44[191], line_43[189], line_42[187], line_41[185], line_40[183], line_39[181], line_38[179], line_37[177], line_36[175], line_35[173], line_34[171], line_33[169], line_32[167], line_31[165], line_30[163], line_29[161], line_28[159], line_27[157], line_26[155], line_25[153], line_24[151], line_23[149], line_22[147], line_21[145], line_20[143], line_19[141], line_18[139], line_17[137], line_16[135], line_15[133], line_14[131], line_13[129], line_12[127], line_11[125], line_10[123], line_9[121], line_8[119], line_7[117], line_6[115], line_5[113], line_4[111], line_3[109], line_2[107], line_1[105] };
assign col_360 = {line_128[360], line_127[358], line_126[356], line_125[354], line_124[352], line_123[350], line_122[348], line_121[346], line_120[344], line_119[342], line_118[340], line_117[338], line_116[336], line_115[334], line_114[332], line_113[330], line_112[328], line_111[326], line_110[324], line_109[322], line_108[320], line_107[318], line_106[316], line_105[314], line_104[312], line_103[310], line_102[308], line_101[306], line_100[304], line_99[302], line_98[300], line_97[298], line_96[296], line_95[294], line_94[292], line_93[290], line_92[288], line_91[286], line_90[284], line_89[282], line_88[280], line_87[278], line_86[276], line_85[274], line_84[272], line_83[270], line_82[268], line_81[266], line_80[264], line_79[262], line_78[260], line_77[258], line_76[256], line_75[254], line_74[252], line_73[250], line_72[248], line_71[246], line_70[244], line_69[242], line_68[240], line_67[238], line_66[236], line_65[234], line_64[232], line_63[230], line_62[228], line_61[226], line_60[224], line_59[222], line_58[220], line_57[218], line_56[216], line_55[214], line_54[212], line_53[210], line_52[208], line_51[206], line_50[204], line_49[202], line_48[200], line_47[198], line_46[196], line_45[194], line_44[192], line_43[190], line_42[188], line_41[186], line_40[184], line_39[182], line_38[180], line_37[178], line_36[176], line_35[174], line_34[172], line_33[170], line_32[168], line_31[166], line_30[164], line_29[162], line_28[160], line_27[158], line_26[156], line_25[154], line_24[152], line_23[150], line_22[148], line_21[146], line_20[144], line_19[142], line_18[140], line_17[138], line_16[136], line_15[134], line_14[132], line_13[130], line_12[128], line_11[126], line_10[124], line_9[122], line_8[120], line_7[118], line_6[116], line_5[114], line_4[112], line_3[110], line_2[108], line_1[106] };
assign col_361 = {line_128[361], line_127[359], line_126[357], line_125[355], line_124[353], line_123[351], line_122[349], line_121[347], line_120[345], line_119[343], line_118[341], line_117[339], line_116[337], line_115[335], line_114[333], line_113[331], line_112[329], line_111[327], line_110[325], line_109[323], line_108[321], line_107[319], line_106[317], line_105[315], line_104[313], line_103[311], line_102[309], line_101[307], line_100[305], line_99[303], line_98[301], line_97[299], line_96[297], line_95[295], line_94[293], line_93[291], line_92[289], line_91[287], line_90[285], line_89[283], line_88[281], line_87[279], line_86[277], line_85[275], line_84[273], line_83[271], line_82[269], line_81[267], line_80[265], line_79[263], line_78[261], line_77[259], line_76[257], line_75[255], line_74[253], line_73[251], line_72[249], line_71[247], line_70[245], line_69[243], line_68[241], line_67[239], line_66[237], line_65[235], line_64[233], line_63[231], line_62[229], line_61[227], line_60[225], line_59[223], line_58[221], line_57[219], line_56[217], line_55[215], line_54[213], line_53[211], line_52[209], line_51[207], line_50[205], line_49[203], line_48[201], line_47[199], line_46[197], line_45[195], line_44[193], line_43[191], line_42[189], line_41[187], line_40[185], line_39[183], line_38[181], line_37[179], line_36[177], line_35[175], line_34[173], line_33[171], line_32[169], line_31[167], line_30[165], line_29[163], line_28[161], line_27[159], line_26[157], line_25[155], line_24[153], line_23[151], line_22[149], line_21[147], line_20[145], line_19[143], line_18[141], line_17[139], line_16[137], line_15[135], line_14[133], line_13[131], line_12[129], line_11[127], line_10[125], line_9[123], line_8[121], line_7[119], line_6[117], line_5[115], line_4[113], line_3[111], line_2[109], line_1[107] };
assign col_362 = {line_128[362], line_127[360], line_126[358], line_125[356], line_124[354], line_123[352], line_122[350], line_121[348], line_120[346], line_119[344], line_118[342], line_117[340], line_116[338], line_115[336], line_114[334], line_113[332], line_112[330], line_111[328], line_110[326], line_109[324], line_108[322], line_107[320], line_106[318], line_105[316], line_104[314], line_103[312], line_102[310], line_101[308], line_100[306], line_99[304], line_98[302], line_97[300], line_96[298], line_95[296], line_94[294], line_93[292], line_92[290], line_91[288], line_90[286], line_89[284], line_88[282], line_87[280], line_86[278], line_85[276], line_84[274], line_83[272], line_82[270], line_81[268], line_80[266], line_79[264], line_78[262], line_77[260], line_76[258], line_75[256], line_74[254], line_73[252], line_72[250], line_71[248], line_70[246], line_69[244], line_68[242], line_67[240], line_66[238], line_65[236], line_64[234], line_63[232], line_62[230], line_61[228], line_60[226], line_59[224], line_58[222], line_57[220], line_56[218], line_55[216], line_54[214], line_53[212], line_52[210], line_51[208], line_50[206], line_49[204], line_48[202], line_47[200], line_46[198], line_45[196], line_44[194], line_43[192], line_42[190], line_41[188], line_40[186], line_39[184], line_38[182], line_37[180], line_36[178], line_35[176], line_34[174], line_33[172], line_32[170], line_31[168], line_30[166], line_29[164], line_28[162], line_27[160], line_26[158], line_25[156], line_24[154], line_23[152], line_22[150], line_21[148], line_20[146], line_19[144], line_18[142], line_17[140], line_16[138], line_15[136], line_14[134], line_13[132], line_12[130], line_11[128], line_10[126], line_9[124], line_8[122], line_7[120], line_6[118], line_5[116], line_4[114], line_3[112], line_2[110], line_1[108] };
assign col_363 = {line_128[363], line_127[361], line_126[359], line_125[357], line_124[355], line_123[353], line_122[351], line_121[349], line_120[347], line_119[345], line_118[343], line_117[341], line_116[339], line_115[337], line_114[335], line_113[333], line_112[331], line_111[329], line_110[327], line_109[325], line_108[323], line_107[321], line_106[319], line_105[317], line_104[315], line_103[313], line_102[311], line_101[309], line_100[307], line_99[305], line_98[303], line_97[301], line_96[299], line_95[297], line_94[295], line_93[293], line_92[291], line_91[289], line_90[287], line_89[285], line_88[283], line_87[281], line_86[279], line_85[277], line_84[275], line_83[273], line_82[271], line_81[269], line_80[267], line_79[265], line_78[263], line_77[261], line_76[259], line_75[257], line_74[255], line_73[253], line_72[251], line_71[249], line_70[247], line_69[245], line_68[243], line_67[241], line_66[239], line_65[237], line_64[235], line_63[233], line_62[231], line_61[229], line_60[227], line_59[225], line_58[223], line_57[221], line_56[219], line_55[217], line_54[215], line_53[213], line_52[211], line_51[209], line_50[207], line_49[205], line_48[203], line_47[201], line_46[199], line_45[197], line_44[195], line_43[193], line_42[191], line_41[189], line_40[187], line_39[185], line_38[183], line_37[181], line_36[179], line_35[177], line_34[175], line_33[173], line_32[171], line_31[169], line_30[167], line_29[165], line_28[163], line_27[161], line_26[159], line_25[157], line_24[155], line_23[153], line_22[151], line_21[149], line_20[147], line_19[145], line_18[143], line_17[141], line_16[139], line_15[137], line_14[135], line_13[133], line_12[131], line_11[129], line_10[127], line_9[125], line_8[123], line_7[121], line_6[119], line_5[117], line_4[115], line_3[113], line_2[111], line_1[109] };
assign col_364 = {line_128[364], line_127[362], line_126[360], line_125[358], line_124[356], line_123[354], line_122[352], line_121[350], line_120[348], line_119[346], line_118[344], line_117[342], line_116[340], line_115[338], line_114[336], line_113[334], line_112[332], line_111[330], line_110[328], line_109[326], line_108[324], line_107[322], line_106[320], line_105[318], line_104[316], line_103[314], line_102[312], line_101[310], line_100[308], line_99[306], line_98[304], line_97[302], line_96[300], line_95[298], line_94[296], line_93[294], line_92[292], line_91[290], line_90[288], line_89[286], line_88[284], line_87[282], line_86[280], line_85[278], line_84[276], line_83[274], line_82[272], line_81[270], line_80[268], line_79[266], line_78[264], line_77[262], line_76[260], line_75[258], line_74[256], line_73[254], line_72[252], line_71[250], line_70[248], line_69[246], line_68[244], line_67[242], line_66[240], line_65[238], line_64[236], line_63[234], line_62[232], line_61[230], line_60[228], line_59[226], line_58[224], line_57[222], line_56[220], line_55[218], line_54[216], line_53[214], line_52[212], line_51[210], line_50[208], line_49[206], line_48[204], line_47[202], line_46[200], line_45[198], line_44[196], line_43[194], line_42[192], line_41[190], line_40[188], line_39[186], line_38[184], line_37[182], line_36[180], line_35[178], line_34[176], line_33[174], line_32[172], line_31[170], line_30[168], line_29[166], line_28[164], line_27[162], line_26[160], line_25[158], line_24[156], line_23[154], line_22[152], line_21[150], line_20[148], line_19[146], line_18[144], line_17[142], line_16[140], line_15[138], line_14[136], line_13[134], line_12[132], line_11[130], line_10[128], line_9[126], line_8[124], line_7[122], line_6[120], line_5[118], line_4[116], line_3[114], line_2[112], line_1[110] };
assign col_365 = {line_128[365], line_127[363], line_126[361], line_125[359], line_124[357], line_123[355], line_122[353], line_121[351], line_120[349], line_119[347], line_118[345], line_117[343], line_116[341], line_115[339], line_114[337], line_113[335], line_112[333], line_111[331], line_110[329], line_109[327], line_108[325], line_107[323], line_106[321], line_105[319], line_104[317], line_103[315], line_102[313], line_101[311], line_100[309], line_99[307], line_98[305], line_97[303], line_96[301], line_95[299], line_94[297], line_93[295], line_92[293], line_91[291], line_90[289], line_89[287], line_88[285], line_87[283], line_86[281], line_85[279], line_84[277], line_83[275], line_82[273], line_81[271], line_80[269], line_79[267], line_78[265], line_77[263], line_76[261], line_75[259], line_74[257], line_73[255], line_72[253], line_71[251], line_70[249], line_69[247], line_68[245], line_67[243], line_66[241], line_65[239], line_64[237], line_63[235], line_62[233], line_61[231], line_60[229], line_59[227], line_58[225], line_57[223], line_56[221], line_55[219], line_54[217], line_53[215], line_52[213], line_51[211], line_50[209], line_49[207], line_48[205], line_47[203], line_46[201], line_45[199], line_44[197], line_43[195], line_42[193], line_41[191], line_40[189], line_39[187], line_38[185], line_37[183], line_36[181], line_35[179], line_34[177], line_33[175], line_32[173], line_31[171], line_30[169], line_29[167], line_28[165], line_27[163], line_26[161], line_25[159], line_24[157], line_23[155], line_22[153], line_21[151], line_20[149], line_19[147], line_18[145], line_17[143], line_16[141], line_15[139], line_14[137], line_13[135], line_12[133], line_11[131], line_10[129], line_9[127], line_8[125], line_7[123], line_6[121], line_5[119], line_4[117], line_3[115], line_2[113], line_1[111] };
assign col_366 = {line_128[366], line_127[364], line_126[362], line_125[360], line_124[358], line_123[356], line_122[354], line_121[352], line_120[350], line_119[348], line_118[346], line_117[344], line_116[342], line_115[340], line_114[338], line_113[336], line_112[334], line_111[332], line_110[330], line_109[328], line_108[326], line_107[324], line_106[322], line_105[320], line_104[318], line_103[316], line_102[314], line_101[312], line_100[310], line_99[308], line_98[306], line_97[304], line_96[302], line_95[300], line_94[298], line_93[296], line_92[294], line_91[292], line_90[290], line_89[288], line_88[286], line_87[284], line_86[282], line_85[280], line_84[278], line_83[276], line_82[274], line_81[272], line_80[270], line_79[268], line_78[266], line_77[264], line_76[262], line_75[260], line_74[258], line_73[256], line_72[254], line_71[252], line_70[250], line_69[248], line_68[246], line_67[244], line_66[242], line_65[240], line_64[238], line_63[236], line_62[234], line_61[232], line_60[230], line_59[228], line_58[226], line_57[224], line_56[222], line_55[220], line_54[218], line_53[216], line_52[214], line_51[212], line_50[210], line_49[208], line_48[206], line_47[204], line_46[202], line_45[200], line_44[198], line_43[196], line_42[194], line_41[192], line_40[190], line_39[188], line_38[186], line_37[184], line_36[182], line_35[180], line_34[178], line_33[176], line_32[174], line_31[172], line_30[170], line_29[168], line_28[166], line_27[164], line_26[162], line_25[160], line_24[158], line_23[156], line_22[154], line_21[152], line_20[150], line_19[148], line_18[146], line_17[144], line_16[142], line_15[140], line_14[138], line_13[136], line_12[134], line_11[132], line_10[130], line_9[128], line_8[126], line_7[124], line_6[122], line_5[120], line_4[118], line_3[116], line_2[114], line_1[112] };
assign col_367 = {line_128[367], line_127[365], line_126[363], line_125[361], line_124[359], line_123[357], line_122[355], line_121[353], line_120[351], line_119[349], line_118[347], line_117[345], line_116[343], line_115[341], line_114[339], line_113[337], line_112[335], line_111[333], line_110[331], line_109[329], line_108[327], line_107[325], line_106[323], line_105[321], line_104[319], line_103[317], line_102[315], line_101[313], line_100[311], line_99[309], line_98[307], line_97[305], line_96[303], line_95[301], line_94[299], line_93[297], line_92[295], line_91[293], line_90[291], line_89[289], line_88[287], line_87[285], line_86[283], line_85[281], line_84[279], line_83[277], line_82[275], line_81[273], line_80[271], line_79[269], line_78[267], line_77[265], line_76[263], line_75[261], line_74[259], line_73[257], line_72[255], line_71[253], line_70[251], line_69[249], line_68[247], line_67[245], line_66[243], line_65[241], line_64[239], line_63[237], line_62[235], line_61[233], line_60[231], line_59[229], line_58[227], line_57[225], line_56[223], line_55[221], line_54[219], line_53[217], line_52[215], line_51[213], line_50[211], line_49[209], line_48[207], line_47[205], line_46[203], line_45[201], line_44[199], line_43[197], line_42[195], line_41[193], line_40[191], line_39[189], line_38[187], line_37[185], line_36[183], line_35[181], line_34[179], line_33[177], line_32[175], line_31[173], line_30[171], line_29[169], line_28[167], line_27[165], line_26[163], line_25[161], line_24[159], line_23[157], line_22[155], line_21[153], line_20[151], line_19[149], line_18[147], line_17[145], line_16[143], line_15[141], line_14[139], line_13[137], line_12[135], line_11[133], line_10[131], line_9[129], line_8[127], line_7[125], line_6[123], line_5[121], line_4[119], line_3[117], line_2[115], line_1[113] };
assign col_368 = {line_128[368], line_127[366], line_126[364], line_125[362], line_124[360], line_123[358], line_122[356], line_121[354], line_120[352], line_119[350], line_118[348], line_117[346], line_116[344], line_115[342], line_114[340], line_113[338], line_112[336], line_111[334], line_110[332], line_109[330], line_108[328], line_107[326], line_106[324], line_105[322], line_104[320], line_103[318], line_102[316], line_101[314], line_100[312], line_99[310], line_98[308], line_97[306], line_96[304], line_95[302], line_94[300], line_93[298], line_92[296], line_91[294], line_90[292], line_89[290], line_88[288], line_87[286], line_86[284], line_85[282], line_84[280], line_83[278], line_82[276], line_81[274], line_80[272], line_79[270], line_78[268], line_77[266], line_76[264], line_75[262], line_74[260], line_73[258], line_72[256], line_71[254], line_70[252], line_69[250], line_68[248], line_67[246], line_66[244], line_65[242], line_64[240], line_63[238], line_62[236], line_61[234], line_60[232], line_59[230], line_58[228], line_57[226], line_56[224], line_55[222], line_54[220], line_53[218], line_52[216], line_51[214], line_50[212], line_49[210], line_48[208], line_47[206], line_46[204], line_45[202], line_44[200], line_43[198], line_42[196], line_41[194], line_40[192], line_39[190], line_38[188], line_37[186], line_36[184], line_35[182], line_34[180], line_33[178], line_32[176], line_31[174], line_30[172], line_29[170], line_28[168], line_27[166], line_26[164], line_25[162], line_24[160], line_23[158], line_22[156], line_21[154], line_20[152], line_19[150], line_18[148], line_17[146], line_16[144], line_15[142], line_14[140], line_13[138], line_12[136], line_11[134], line_10[132], line_9[130], line_8[128], line_7[126], line_6[124], line_5[122], line_4[120], line_3[118], line_2[116], line_1[114] };
assign col_369 = {line_128[369], line_127[367], line_126[365], line_125[363], line_124[361], line_123[359], line_122[357], line_121[355], line_120[353], line_119[351], line_118[349], line_117[347], line_116[345], line_115[343], line_114[341], line_113[339], line_112[337], line_111[335], line_110[333], line_109[331], line_108[329], line_107[327], line_106[325], line_105[323], line_104[321], line_103[319], line_102[317], line_101[315], line_100[313], line_99[311], line_98[309], line_97[307], line_96[305], line_95[303], line_94[301], line_93[299], line_92[297], line_91[295], line_90[293], line_89[291], line_88[289], line_87[287], line_86[285], line_85[283], line_84[281], line_83[279], line_82[277], line_81[275], line_80[273], line_79[271], line_78[269], line_77[267], line_76[265], line_75[263], line_74[261], line_73[259], line_72[257], line_71[255], line_70[253], line_69[251], line_68[249], line_67[247], line_66[245], line_65[243], line_64[241], line_63[239], line_62[237], line_61[235], line_60[233], line_59[231], line_58[229], line_57[227], line_56[225], line_55[223], line_54[221], line_53[219], line_52[217], line_51[215], line_50[213], line_49[211], line_48[209], line_47[207], line_46[205], line_45[203], line_44[201], line_43[199], line_42[197], line_41[195], line_40[193], line_39[191], line_38[189], line_37[187], line_36[185], line_35[183], line_34[181], line_33[179], line_32[177], line_31[175], line_30[173], line_29[171], line_28[169], line_27[167], line_26[165], line_25[163], line_24[161], line_23[159], line_22[157], line_21[155], line_20[153], line_19[151], line_18[149], line_17[147], line_16[145], line_15[143], line_14[141], line_13[139], line_12[137], line_11[135], line_10[133], line_9[131], line_8[129], line_7[127], line_6[125], line_5[123], line_4[121], line_3[119], line_2[117], line_1[115] };
assign col_370 = {line_128[370], line_127[368], line_126[366], line_125[364], line_124[362], line_123[360], line_122[358], line_121[356], line_120[354], line_119[352], line_118[350], line_117[348], line_116[346], line_115[344], line_114[342], line_113[340], line_112[338], line_111[336], line_110[334], line_109[332], line_108[330], line_107[328], line_106[326], line_105[324], line_104[322], line_103[320], line_102[318], line_101[316], line_100[314], line_99[312], line_98[310], line_97[308], line_96[306], line_95[304], line_94[302], line_93[300], line_92[298], line_91[296], line_90[294], line_89[292], line_88[290], line_87[288], line_86[286], line_85[284], line_84[282], line_83[280], line_82[278], line_81[276], line_80[274], line_79[272], line_78[270], line_77[268], line_76[266], line_75[264], line_74[262], line_73[260], line_72[258], line_71[256], line_70[254], line_69[252], line_68[250], line_67[248], line_66[246], line_65[244], line_64[242], line_63[240], line_62[238], line_61[236], line_60[234], line_59[232], line_58[230], line_57[228], line_56[226], line_55[224], line_54[222], line_53[220], line_52[218], line_51[216], line_50[214], line_49[212], line_48[210], line_47[208], line_46[206], line_45[204], line_44[202], line_43[200], line_42[198], line_41[196], line_40[194], line_39[192], line_38[190], line_37[188], line_36[186], line_35[184], line_34[182], line_33[180], line_32[178], line_31[176], line_30[174], line_29[172], line_28[170], line_27[168], line_26[166], line_25[164], line_24[162], line_23[160], line_22[158], line_21[156], line_20[154], line_19[152], line_18[150], line_17[148], line_16[146], line_15[144], line_14[142], line_13[140], line_12[138], line_11[136], line_10[134], line_9[132], line_8[130], line_7[128], line_6[126], line_5[124], line_4[122], line_3[120], line_2[118], line_1[116] };
assign col_371 = {line_128[371], line_127[369], line_126[367], line_125[365], line_124[363], line_123[361], line_122[359], line_121[357], line_120[355], line_119[353], line_118[351], line_117[349], line_116[347], line_115[345], line_114[343], line_113[341], line_112[339], line_111[337], line_110[335], line_109[333], line_108[331], line_107[329], line_106[327], line_105[325], line_104[323], line_103[321], line_102[319], line_101[317], line_100[315], line_99[313], line_98[311], line_97[309], line_96[307], line_95[305], line_94[303], line_93[301], line_92[299], line_91[297], line_90[295], line_89[293], line_88[291], line_87[289], line_86[287], line_85[285], line_84[283], line_83[281], line_82[279], line_81[277], line_80[275], line_79[273], line_78[271], line_77[269], line_76[267], line_75[265], line_74[263], line_73[261], line_72[259], line_71[257], line_70[255], line_69[253], line_68[251], line_67[249], line_66[247], line_65[245], line_64[243], line_63[241], line_62[239], line_61[237], line_60[235], line_59[233], line_58[231], line_57[229], line_56[227], line_55[225], line_54[223], line_53[221], line_52[219], line_51[217], line_50[215], line_49[213], line_48[211], line_47[209], line_46[207], line_45[205], line_44[203], line_43[201], line_42[199], line_41[197], line_40[195], line_39[193], line_38[191], line_37[189], line_36[187], line_35[185], line_34[183], line_33[181], line_32[179], line_31[177], line_30[175], line_29[173], line_28[171], line_27[169], line_26[167], line_25[165], line_24[163], line_23[161], line_22[159], line_21[157], line_20[155], line_19[153], line_18[151], line_17[149], line_16[147], line_15[145], line_14[143], line_13[141], line_12[139], line_11[137], line_10[135], line_9[133], line_8[131], line_7[129], line_6[127], line_5[125], line_4[123], line_3[121], line_2[119], line_1[117] };
assign col_372 = {line_128[372], line_127[370], line_126[368], line_125[366], line_124[364], line_123[362], line_122[360], line_121[358], line_120[356], line_119[354], line_118[352], line_117[350], line_116[348], line_115[346], line_114[344], line_113[342], line_112[340], line_111[338], line_110[336], line_109[334], line_108[332], line_107[330], line_106[328], line_105[326], line_104[324], line_103[322], line_102[320], line_101[318], line_100[316], line_99[314], line_98[312], line_97[310], line_96[308], line_95[306], line_94[304], line_93[302], line_92[300], line_91[298], line_90[296], line_89[294], line_88[292], line_87[290], line_86[288], line_85[286], line_84[284], line_83[282], line_82[280], line_81[278], line_80[276], line_79[274], line_78[272], line_77[270], line_76[268], line_75[266], line_74[264], line_73[262], line_72[260], line_71[258], line_70[256], line_69[254], line_68[252], line_67[250], line_66[248], line_65[246], line_64[244], line_63[242], line_62[240], line_61[238], line_60[236], line_59[234], line_58[232], line_57[230], line_56[228], line_55[226], line_54[224], line_53[222], line_52[220], line_51[218], line_50[216], line_49[214], line_48[212], line_47[210], line_46[208], line_45[206], line_44[204], line_43[202], line_42[200], line_41[198], line_40[196], line_39[194], line_38[192], line_37[190], line_36[188], line_35[186], line_34[184], line_33[182], line_32[180], line_31[178], line_30[176], line_29[174], line_28[172], line_27[170], line_26[168], line_25[166], line_24[164], line_23[162], line_22[160], line_21[158], line_20[156], line_19[154], line_18[152], line_17[150], line_16[148], line_15[146], line_14[144], line_13[142], line_12[140], line_11[138], line_10[136], line_9[134], line_8[132], line_7[130], line_6[128], line_5[126], line_4[124], line_3[122], line_2[120], line_1[118] };
assign col_373 = {line_128[373], line_127[371], line_126[369], line_125[367], line_124[365], line_123[363], line_122[361], line_121[359], line_120[357], line_119[355], line_118[353], line_117[351], line_116[349], line_115[347], line_114[345], line_113[343], line_112[341], line_111[339], line_110[337], line_109[335], line_108[333], line_107[331], line_106[329], line_105[327], line_104[325], line_103[323], line_102[321], line_101[319], line_100[317], line_99[315], line_98[313], line_97[311], line_96[309], line_95[307], line_94[305], line_93[303], line_92[301], line_91[299], line_90[297], line_89[295], line_88[293], line_87[291], line_86[289], line_85[287], line_84[285], line_83[283], line_82[281], line_81[279], line_80[277], line_79[275], line_78[273], line_77[271], line_76[269], line_75[267], line_74[265], line_73[263], line_72[261], line_71[259], line_70[257], line_69[255], line_68[253], line_67[251], line_66[249], line_65[247], line_64[245], line_63[243], line_62[241], line_61[239], line_60[237], line_59[235], line_58[233], line_57[231], line_56[229], line_55[227], line_54[225], line_53[223], line_52[221], line_51[219], line_50[217], line_49[215], line_48[213], line_47[211], line_46[209], line_45[207], line_44[205], line_43[203], line_42[201], line_41[199], line_40[197], line_39[195], line_38[193], line_37[191], line_36[189], line_35[187], line_34[185], line_33[183], line_32[181], line_31[179], line_30[177], line_29[175], line_28[173], line_27[171], line_26[169], line_25[167], line_24[165], line_23[163], line_22[161], line_21[159], line_20[157], line_19[155], line_18[153], line_17[151], line_16[149], line_15[147], line_14[145], line_13[143], line_12[141], line_11[139], line_10[137], line_9[135], line_8[133], line_7[131], line_6[129], line_5[127], line_4[125], line_3[123], line_2[121], line_1[119] };
assign col_374 = {line_128[374], line_127[372], line_126[370], line_125[368], line_124[366], line_123[364], line_122[362], line_121[360], line_120[358], line_119[356], line_118[354], line_117[352], line_116[350], line_115[348], line_114[346], line_113[344], line_112[342], line_111[340], line_110[338], line_109[336], line_108[334], line_107[332], line_106[330], line_105[328], line_104[326], line_103[324], line_102[322], line_101[320], line_100[318], line_99[316], line_98[314], line_97[312], line_96[310], line_95[308], line_94[306], line_93[304], line_92[302], line_91[300], line_90[298], line_89[296], line_88[294], line_87[292], line_86[290], line_85[288], line_84[286], line_83[284], line_82[282], line_81[280], line_80[278], line_79[276], line_78[274], line_77[272], line_76[270], line_75[268], line_74[266], line_73[264], line_72[262], line_71[260], line_70[258], line_69[256], line_68[254], line_67[252], line_66[250], line_65[248], line_64[246], line_63[244], line_62[242], line_61[240], line_60[238], line_59[236], line_58[234], line_57[232], line_56[230], line_55[228], line_54[226], line_53[224], line_52[222], line_51[220], line_50[218], line_49[216], line_48[214], line_47[212], line_46[210], line_45[208], line_44[206], line_43[204], line_42[202], line_41[200], line_40[198], line_39[196], line_38[194], line_37[192], line_36[190], line_35[188], line_34[186], line_33[184], line_32[182], line_31[180], line_30[178], line_29[176], line_28[174], line_27[172], line_26[170], line_25[168], line_24[166], line_23[164], line_22[162], line_21[160], line_20[158], line_19[156], line_18[154], line_17[152], line_16[150], line_15[148], line_14[146], line_13[144], line_12[142], line_11[140], line_10[138], line_9[136], line_8[134], line_7[132], line_6[130], line_5[128], line_4[126], line_3[124], line_2[122], line_1[120] };
assign col_375 = {line_128[375], line_127[373], line_126[371], line_125[369], line_124[367], line_123[365], line_122[363], line_121[361], line_120[359], line_119[357], line_118[355], line_117[353], line_116[351], line_115[349], line_114[347], line_113[345], line_112[343], line_111[341], line_110[339], line_109[337], line_108[335], line_107[333], line_106[331], line_105[329], line_104[327], line_103[325], line_102[323], line_101[321], line_100[319], line_99[317], line_98[315], line_97[313], line_96[311], line_95[309], line_94[307], line_93[305], line_92[303], line_91[301], line_90[299], line_89[297], line_88[295], line_87[293], line_86[291], line_85[289], line_84[287], line_83[285], line_82[283], line_81[281], line_80[279], line_79[277], line_78[275], line_77[273], line_76[271], line_75[269], line_74[267], line_73[265], line_72[263], line_71[261], line_70[259], line_69[257], line_68[255], line_67[253], line_66[251], line_65[249], line_64[247], line_63[245], line_62[243], line_61[241], line_60[239], line_59[237], line_58[235], line_57[233], line_56[231], line_55[229], line_54[227], line_53[225], line_52[223], line_51[221], line_50[219], line_49[217], line_48[215], line_47[213], line_46[211], line_45[209], line_44[207], line_43[205], line_42[203], line_41[201], line_40[199], line_39[197], line_38[195], line_37[193], line_36[191], line_35[189], line_34[187], line_33[185], line_32[183], line_31[181], line_30[179], line_29[177], line_28[175], line_27[173], line_26[171], line_25[169], line_24[167], line_23[165], line_22[163], line_21[161], line_20[159], line_19[157], line_18[155], line_17[153], line_16[151], line_15[149], line_14[147], line_13[145], line_12[143], line_11[141], line_10[139], line_9[137], line_8[135], line_7[133], line_6[131], line_5[129], line_4[127], line_3[125], line_2[123], line_1[121] };
assign col_376 = {line_128[376], line_127[374], line_126[372], line_125[370], line_124[368], line_123[366], line_122[364], line_121[362], line_120[360], line_119[358], line_118[356], line_117[354], line_116[352], line_115[350], line_114[348], line_113[346], line_112[344], line_111[342], line_110[340], line_109[338], line_108[336], line_107[334], line_106[332], line_105[330], line_104[328], line_103[326], line_102[324], line_101[322], line_100[320], line_99[318], line_98[316], line_97[314], line_96[312], line_95[310], line_94[308], line_93[306], line_92[304], line_91[302], line_90[300], line_89[298], line_88[296], line_87[294], line_86[292], line_85[290], line_84[288], line_83[286], line_82[284], line_81[282], line_80[280], line_79[278], line_78[276], line_77[274], line_76[272], line_75[270], line_74[268], line_73[266], line_72[264], line_71[262], line_70[260], line_69[258], line_68[256], line_67[254], line_66[252], line_65[250], line_64[248], line_63[246], line_62[244], line_61[242], line_60[240], line_59[238], line_58[236], line_57[234], line_56[232], line_55[230], line_54[228], line_53[226], line_52[224], line_51[222], line_50[220], line_49[218], line_48[216], line_47[214], line_46[212], line_45[210], line_44[208], line_43[206], line_42[204], line_41[202], line_40[200], line_39[198], line_38[196], line_37[194], line_36[192], line_35[190], line_34[188], line_33[186], line_32[184], line_31[182], line_30[180], line_29[178], line_28[176], line_27[174], line_26[172], line_25[170], line_24[168], line_23[166], line_22[164], line_21[162], line_20[160], line_19[158], line_18[156], line_17[154], line_16[152], line_15[150], line_14[148], line_13[146], line_12[144], line_11[142], line_10[140], line_9[138], line_8[136], line_7[134], line_6[132], line_5[130], line_4[128], line_3[126], line_2[124], line_1[122] };
assign col_377 = {line_128[377], line_127[375], line_126[373], line_125[371], line_124[369], line_123[367], line_122[365], line_121[363], line_120[361], line_119[359], line_118[357], line_117[355], line_116[353], line_115[351], line_114[349], line_113[347], line_112[345], line_111[343], line_110[341], line_109[339], line_108[337], line_107[335], line_106[333], line_105[331], line_104[329], line_103[327], line_102[325], line_101[323], line_100[321], line_99[319], line_98[317], line_97[315], line_96[313], line_95[311], line_94[309], line_93[307], line_92[305], line_91[303], line_90[301], line_89[299], line_88[297], line_87[295], line_86[293], line_85[291], line_84[289], line_83[287], line_82[285], line_81[283], line_80[281], line_79[279], line_78[277], line_77[275], line_76[273], line_75[271], line_74[269], line_73[267], line_72[265], line_71[263], line_70[261], line_69[259], line_68[257], line_67[255], line_66[253], line_65[251], line_64[249], line_63[247], line_62[245], line_61[243], line_60[241], line_59[239], line_58[237], line_57[235], line_56[233], line_55[231], line_54[229], line_53[227], line_52[225], line_51[223], line_50[221], line_49[219], line_48[217], line_47[215], line_46[213], line_45[211], line_44[209], line_43[207], line_42[205], line_41[203], line_40[201], line_39[199], line_38[197], line_37[195], line_36[193], line_35[191], line_34[189], line_33[187], line_32[185], line_31[183], line_30[181], line_29[179], line_28[177], line_27[175], line_26[173], line_25[171], line_24[169], line_23[167], line_22[165], line_21[163], line_20[161], line_19[159], line_18[157], line_17[155], line_16[153], line_15[151], line_14[149], line_13[147], line_12[145], line_11[143], line_10[141], line_9[139], line_8[137], line_7[135], line_6[133], line_5[131], line_4[129], line_3[127], line_2[125], line_1[123] };
assign col_378 = {line_128[378], line_127[376], line_126[374], line_125[372], line_124[370], line_123[368], line_122[366], line_121[364], line_120[362], line_119[360], line_118[358], line_117[356], line_116[354], line_115[352], line_114[350], line_113[348], line_112[346], line_111[344], line_110[342], line_109[340], line_108[338], line_107[336], line_106[334], line_105[332], line_104[330], line_103[328], line_102[326], line_101[324], line_100[322], line_99[320], line_98[318], line_97[316], line_96[314], line_95[312], line_94[310], line_93[308], line_92[306], line_91[304], line_90[302], line_89[300], line_88[298], line_87[296], line_86[294], line_85[292], line_84[290], line_83[288], line_82[286], line_81[284], line_80[282], line_79[280], line_78[278], line_77[276], line_76[274], line_75[272], line_74[270], line_73[268], line_72[266], line_71[264], line_70[262], line_69[260], line_68[258], line_67[256], line_66[254], line_65[252], line_64[250], line_63[248], line_62[246], line_61[244], line_60[242], line_59[240], line_58[238], line_57[236], line_56[234], line_55[232], line_54[230], line_53[228], line_52[226], line_51[224], line_50[222], line_49[220], line_48[218], line_47[216], line_46[214], line_45[212], line_44[210], line_43[208], line_42[206], line_41[204], line_40[202], line_39[200], line_38[198], line_37[196], line_36[194], line_35[192], line_34[190], line_33[188], line_32[186], line_31[184], line_30[182], line_29[180], line_28[178], line_27[176], line_26[174], line_25[172], line_24[170], line_23[168], line_22[166], line_21[164], line_20[162], line_19[160], line_18[158], line_17[156], line_16[154], line_15[152], line_14[150], line_13[148], line_12[146], line_11[144], line_10[142], line_9[140], line_8[138], line_7[136], line_6[134], line_5[132], line_4[130], line_3[128], line_2[126], line_1[124] };
assign col_379 = {line_128[379], line_127[377], line_126[375], line_125[373], line_124[371], line_123[369], line_122[367], line_121[365], line_120[363], line_119[361], line_118[359], line_117[357], line_116[355], line_115[353], line_114[351], line_113[349], line_112[347], line_111[345], line_110[343], line_109[341], line_108[339], line_107[337], line_106[335], line_105[333], line_104[331], line_103[329], line_102[327], line_101[325], line_100[323], line_99[321], line_98[319], line_97[317], line_96[315], line_95[313], line_94[311], line_93[309], line_92[307], line_91[305], line_90[303], line_89[301], line_88[299], line_87[297], line_86[295], line_85[293], line_84[291], line_83[289], line_82[287], line_81[285], line_80[283], line_79[281], line_78[279], line_77[277], line_76[275], line_75[273], line_74[271], line_73[269], line_72[267], line_71[265], line_70[263], line_69[261], line_68[259], line_67[257], line_66[255], line_65[253], line_64[251], line_63[249], line_62[247], line_61[245], line_60[243], line_59[241], line_58[239], line_57[237], line_56[235], line_55[233], line_54[231], line_53[229], line_52[227], line_51[225], line_50[223], line_49[221], line_48[219], line_47[217], line_46[215], line_45[213], line_44[211], line_43[209], line_42[207], line_41[205], line_40[203], line_39[201], line_38[199], line_37[197], line_36[195], line_35[193], line_34[191], line_33[189], line_32[187], line_31[185], line_30[183], line_29[181], line_28[179], line_27[177], line_26[175], line_25[173], line_24[171], line_23[169], line_22[167], line_21[165], line_20[163], line_19[161], line_18[159], line_17[157], line_16[155], line_15[153], line_14[151], line_13[149], line_12[147], line_11[145], line_10[143], line_9[141], line_8[139], line_7[137], line_6[135], line_5[133], line_4[131], line_3[129], line_2[127], line_1[125] };
assign col_380 = {line_128[380], line_127[378], line_126[376], line_125[374], line_124[372], line_123[370], line_122[368], line_121[366], line_120[364], line_119[362], line_118[360], line_117[358], line_116[356], line_115[354], line_114[352], line_113[350], line_112[348], line_111[346], line_110[344], line_109[342], line_108[340], line_107[338], line_106[336], line_105[334], line_104[332], line_103[330], line_102[328], line_101[326], line_100[324], line_99[322], line_98[320], line_97[318], line_96[316], line_95[314], line_94[312], line_93[310], line_92[308], line_91[306], line_90[304], line_89[302], line_88[300], line_87[298], line_86[296], line_85[294], line_84[292], line_83[290], line_82[288], line_81[286], line_80[284], line_79[282], line_78[280], line_77[278], line_76[276], line_75[274], line_74[272], line_73[270], line_72[268], line_71[266], line_70[264], line_69[262], line_68[260], line_67[258], line_66[256], line_65[254], line_64[252], line_63[250], line_62[248], line_61[246], line_60[244], line_59[242], line_58[240], line_57[238], line_56[236], line_55[234], line_54[232], line_53[230], line_52[228], line_51[226], line_50[224], line_49[222], line_48[220], line_47[218], line_46[216], line_45[214], line_44[212], line_43[210], line_42[208], line_41[206], line_40[204], line_39[202], line_38[200], line_37[198], line_36[196], line_35[194], line_34[192], line_33[190], line_32[188], line_31[186], line_30[184], line_29[182], line_28[180], line_27[178], line_26[176], line_25[174], line_24[172], line_23[170], line_22[168], line_21[166], line_20[164], line_19[162], line_18[160], line_17[158], line_16[156], line_15[154], line_14[152], line_13[150], line_12[148], line_11[146], line_10[144], line_9[142], line_8[140], line_7[138], line_6[136], line_5[134], line_4[132], line_3[130], line_2[128], line_1[126] };
assign col_381 = {line_128[381], line_127[379], line_126[377], line_125[375], line_124[373], line_123[371], line_122[369], line_121[367], line_120[365], line_119[363], line_118[361], line_117[359], line_116[357], line_115[355], line_114[353], line_113[351], line_112[349], line_111[347], line_110[345], line_109[343], line_108[341], line_107[339], line_106[337], line_105[335], line_104[333], line_103[331], line_102[329], line_101[327], line_100[325], line_99[323], line_98[321], line_97[319], line_96[317], line_95[315], line_94[313], line_93[311], line_92[309], line_91[307], line_90[305], line_89[303], line_88[301], line_87[299], line_86[297], line_85[295], line_84[293], line_83[291], line_82[289], line_81[287], line_80[285], line_79[283], line_78[281], line_77[279], line_76[277], line_75[275], line_74[273], line_73[271], line_72[269], line_71[267], line_70[265], line_69[263], line_68[261], line_67[259], line_66[257], line_65[255], line_64[253], line_63[251], line_62[249], line_61[247], line_60[245], line_59[243], line_58[241], line_57[239], line_56[237], line_55[235], line_54[233], line_53[231], line_52[229], line_51[227], line_50[225], line_49[223], line_48[221], line_47[219], line_46[217], line_45[215], line_44[213], line_43[211], line_42[209], line_41[207], line_40[205], line_39[203], line_38[201], line_37[199], line_36[197], line_35[195], line_34[193], line_33[191], line_32[189], line_31[187], line_30[185], line_29[183], line_28[181], line_27[179], line_26[177], line_25[175], line_24[173], line_23[171], line_22[169], line_21[167], line_20[165], line_19[163], line_18[161], line_17[159], line_16[157], line_15[155], line_14[153], line_13[151], line_12[149], line_11[147], line_10[145], line_9[143], line_8[141], line_7[139], line_6[137], line_5[135], line_4[133], line_3[131], line_2[129], line_1[127] };
assign col_382 = {line_128[382], line_127[380], line_126[378], line_125[376], line_124[374], line_123[372], line_122[370], line_121[368], line_120[366], line_119[364], line_118[362], line_117[360], line_116[358], line_115[356], line_114[354], line_113[352], line_112[350], line_111[348], line_110[346], line_109[344], line_108[342], line_107[340], line_106[338], line_105[336], line_104[334], line_103[332], line_102[330], line_101[328], line_100[326], line_99[324], line_98[322], line_97[320], line_96[318], line_95[316], line_94[314], line_93[312], line_92[310], line_91[308], line_90[306], line_89[304], line_88[302], line_87[300], line_86[298], line_85[296], line_84[294], line_83[292], line_82[290], line_81[288], line_80[286], line_79[284], line_78[282], line_77[280], line_76[278], line_75[276], line_74[274], line_73[272], line_72[270], line_71[268], line_70[266], line_69[264], line_68[262], line_67[260], line_66[258], line_65[256], line_64[254], line_63[252], line_62[250], line_61[248], line_60[246], line_59[244], line_58[242], line_57[240], line_56[238], line_55[236], line_54[234], line_53[232], line_52[230], line_51[228], line_50[226], line_49[224], line_48[222], line_47[220], line_46[218], line_45[216], line_44[214], line_43[212], line_42[210], line_41[208], line_40[206], line_39[204], line_38[202], line_37[200], line_36[198], line_35[196], line_34[194], line_33[192], line_32[190], line_31[188], line_30[186], line_29[184], line_28[182], line_27[180], line_26[178], line_25[176], line_24[174], line_23[172], line_22[170], line_21[168], line_20[166], line_19[164], line_18[162], line_17[160], line_16[158], line_15[156], line_14[154], line_13[152], line_12[150], line_11[148], line_10[146], line_9[144], line_8[142], line_7[140], line_6[138], line_5[136], line_4[134], line_3[132], line_2[130], line_1[128] };
assign col_383 = {line_128[383], line_127[381], line_126[379], line_125[377], line_124[375], line_123[373], line_122[371], line_121[369], line_120[367], line_119[365], line_118[363], line_117[361], line_116[359], line_115[357], line_114[355], line_113[353], line_112[351], line_111[349], line_110[347], line_109[345], line_108[343], line_107[341], line_106[339], line_105[337], line_104[335], line_103[333], line_102[331], line_101[329], line_100[327], line_99[325], line_98[323], line_97[321], line_96[319], line_95[317], line_94[315], line_93[313], line_92[311], line_91[309], line_90[307], line_89[305], line_88[303], line_87[301], line_86[299], line_85[297], line_84[295], line_83[293], line_82[291], line_81[289], line_80[287], line_79[285], line_78[283], line_77[281], line_76[279], line_75[277], line_74[275], line_73[273], line_72[271], line_71[269], line_70[267], line_69[265], line_68[263], line_67[261], line_66[259], line_65[257], line_64[255], line_63[253], line_62[251], line_61[249], line_60[247], line_59[245], line_58[243], line_57[241], line_56[239], line_55[237], line_54[235], line_53[233], line_52[231], line_51[229], line_50[227], line_49[225], line_48[223], line_47[221], line_46[219], line_45[217], line_44[215], line_43[213], line_42[211], line_41[209], line_40[207], line_39[205], line_38[203], line_37[201], line_36[199], line_35[197], line_34[195], line_33[193], line_32[191], line_31[189], line_30[187], line_29[185], line_28[183], line_27[181], line_26[179], line_25[177], line_24[175], line_23[173], line_22[171], line_21[169], line_20[167], line_19[165], line_18[163], line_17[161], line_16[159], line_15[157], line_14[155], line_13[153], line_12[151], line_11[149], line_10[147], line_9[145], line_8[143], line_7[141], line_6[139], line_5[137], line_4[135], line_3[133], line_2[131], line_1[129] };
assign col_384 = {line_128[384], line_127[382], line_126[380], line_125[378], line_124[376], line_123[374], line_122[372], line_121[370], line_120[368], line_119[366], line_118[364], line_117[362], line_116[360], line_115[358], line_114[356], line_113[354], line_112[352], line_111[350], line_110[348], line_109[346], line_108[344], line_107[342], line_106[340], line_105[338], line_104[336], line_103[334], line_102[332], line_101[330], line_100[328], line_99[326], line_98[324], line_97[322], line_96[320], line_95[318], line_94[316], line_93[314], line_92[312], line_91[310], line_90[308], line_89[306], line_88[304], line_87[302], line_86[300], line_85[298], line_84[296], line_83[294], line_82[292], line_81[290], line_80[288], line_79[286], line_78[284], line_77[282], line_76[280], line_75[278], line_74[276], line_73[274], line_72[272], line_71[270], line_70[268], line_69[266], line_68[264], line_67[262], line_66[260], line_65[258], line_64[256], line_63[254], line_62[252], line_61[250], line_60[248], line_59[246], line_58[244], line_57[242], line_56[240], line_55[238], line_54[236], line_53[234], line_52[232], line_51[230], line_50[228], line_49[226], line_48[224], line_47[222], line_46[220], line_45[218], line_44[216], line_43[214], line_42[212], line_41[210], line_40[208], line_39[206], line_38[204], line_37[202], line_36[200], line_35[198], line_34[196], line_33[194], line_32[192], line_31[190], line_30[188], line_29[186], line_28[184], line_27[182], line_26[180], line_25[178], line_24[176], line_23[174], line_22[172], line_21[170], line_20[168], line_19[166], line_18[164], line_17[162], line_16[160], line_15[158], line_14[156], line_13[154], line_12[152], line_11[150], line_10[148], line_9[146], line_8[144], line_7[142], line_6[140], line_5[138], line_4[136], line_3[134], line_2[132], line_1[130] };
assign col_385 = {line_128[385], line_127[383], line_126[381], line_125[379], line_124[377], line_123[375], line_122[373], line_121[371], line_120[369], line_119[367], line_118[365], line_117[363], line_116[361], line_115[359], line_114[357], line_113[355], line_112[353], line_111[351], line_110[349], line_109[347], line_108[345], line_107[343], line_106[341], line_105[339], line_104[337], line_103[335], line_102[333], line_101[331], line_100[329], line_99[327], line_98[325], line_97[323], line_96[321], line_95[319], line_94[317], line_93[315], line_92[313], line_91[311], line_90[309], line_89[307], line_88[305], line_87[303], line_86[301], line_85[299], line_84[297], line_83[295], line_82[293], line_81[291], line_80[289], line_79[287], line_78[285], line_77[283], line_76[281], line_75[279], line_74[277], line_73[275], line_72[273], line_71[271], line_70[269], line_69[267], line_68[265], line_67[263], line_66[261], line_65[259], line_64[257], line_63[255], line_62[253], line_61[251], line_60[249], line_59[247], line_58[245], line_57[243], line_56[241], line_55[239], line_54[237], line_53[235], line_52[233], line_51[231], line_50[229], line_49[227], line_48[225], line_47[223], line_46[221], line_45[219], line_44[217], line_43[215], line_42[213], line_41[211], line_40[209], line_39[207], line_38[205], line_37[203], line_36[201], line_35[199], line_34[197], line_33[195], line_32[193], line_31[191], line_30[189], line_29[187], line_28[185], line_27[183], line_26[181], line_25[179], line_24[177], line_23[175], line_22[173], line_21[171], line_20[169], line_19[167], line_18[165], line_17[163], line_16[161], line_15[159], line_14[157], line_13[155], line_12[153], line_11[151], line_10[149], line_9[147], line_8[145], line_7[143], line_6[141], line_5[139], line_4[137], line_3[135], line_2[133], line_1[131] };
assign col_386 = {line_128[386], line_127[384], line_126[382], line_125[380], line_124[378], line_123[376], line_122[374], line_121[372], line_120[370], line_119[368], line_118[366], line_117[364], line_116[362], line_115[360], line_114[358], line_113[356], line_112[354], line_111[352], line_110[350], line_109[348], line_108[346], line_107[344], line_106[342], line_105[340], line_104[338], line_103[336], line_102[334], line_101[332], line_100[330], line_99[328], line_98[326], line_97[324], line_96[322], line_95[320], line_94[318], line_93[316], line_92[314], line_91[312], line_90[310], line_89[308], line_88[306], line_87[304], line_86[302], line_85[300], line_84[298], line_83[296], line_82[294], line_81[292], line_80[290], line_79[288], line_78[286], line_77[284], line_76[282], line_75[280], line_74[278], line_73[276], line_72[274], line_71[272], line_70[270], line_69[268], line_68[266], line_67[264], line_66[262], line_65[260], line_64[258], line_63[256], line_62[254], line_61[252], line_60[250], line_59[248], line_58[246], line_57[244], line_56[242], line_55[240], line_54[238], line_53[236], line_52[234], line_51[232], line_50[230], line_49[228], line_48[226], line_47[224], line_46[222], line_45[220], line_44[218], line_43[216], line_42[214], line_41[212], line_40[210], line_39[208], line_38[206], line_37[204], line_36[202], line_35[200], line_34[198], line_33[196], line_32[194], line_31[192], line_30[190], line_29[188], line_28[186], line_27[184], line_26[182], line_25[180], line_24[178], line_23[176], line_22[174], line_21[172], line_20[170], line_19[168], line_18[166], line_17[164], line_16[162], line_15[160], line_14[158], line_13[156], line_12[154], line_11[152], line_10[150], line_9[148], line_8[146], line_7[144], line_6[142], line_5[140], line_4[138], line_3[136], line_2[134], line_1[132] };
assign col_387 = {line_128[387], line_127[385], line_126[383], line_125[381], line_124[379], line_123[377], line_122[375], line_121[373], line_120[371], line_119[369], line_118[367], line_117[365], line_116[363], line_115[361], line_114[359], line_113[357], line_112[355], line_111[353], line_110[351], line_109[349], line_108[347], line_107[345], line_106[343], line_105[341], line_104[339], line_103[337], line_102[335], line_101[333], line_100[331], line_99[329], line_98[327], line_97[325], line_96[323], line_95[321], line_94[319], line_93[317], line_92[315], line_91[313], line_90[311], line_89[309], line_88[307], line_87[305], line_86[303], line_85[301], line_84[299], line_83[297], line_82[295], line_81[293], line_80[291], line_79[289], line_78[287], line_77[285], line_76[283], line_75[281], line_74[279], line_73[277], line_72[275], line_71[273], line_70[271], line_69[269], line_68[267], line_67[265], line_66[263], line_65[261], line_64[259], line_63[257], line_62[255], line_61[253], line_60[251], line_59[249], line_58[247], line_57[245], line_56[243], line_55[241], line_54[239], line_53[237], line_52[235], line_51[233], line_50[231], line_49[229], line_48[227], line_47[225], line_46[223], line_45[221], line_44[219], line_43[217], line_42[215], line_41[213], line_40[211], line_39[209], line_38[207], line_37[205], line_36[203], line_35[201], line_34[199], line_33[197], line_32[195], line_31[193], line_30[191], line_29[189], line_28[187], line_27[185], line_26[183], line_25[181], line_24[179], line_23[177], line_22[175], line_21[173], line_20[171], line_19[169], line_18[167], line_17[165], line_16[163], line_15[161], line_14[159], line_13[157], line_12[155], line_11[153], line_10[151], line_9[149], line_8[147], line_7[145], line_6[143], line_5[141], line_4[139], line_3[137], line_2[135], line_1[133] };
assign col_388 = {line_128[388], line_127[386], line_126[384], line_125[382], line_124[380], line_123[378], line_122[376], line_121[374], line_120[372], line_119[370], line_118[368], line_117[366], line_116[364], line_115[362], line_114[360], line_113[358], line_112[356], line_111[354], line_110[352], line_109[350], line_108[348], line_107[346], line_106[344], line_105[342], line_104[340], line_103[338], line_102[336], line_101[334], line_100[332], line_99[330], line_98[328], line_97[326], line_96[324], line_95[322], line_94[320], line_93[318], line_92[316], line_91[314], line_90[312], line_89[310], line_88[308], line_87[306], line_86[304], line_85[302], line_84[300], line_83[298], line_82[296], line_81[294], line_80[292], line_79[290], line_78[288], line_77[286], line_76[284], line_75[282], line_74[280], line_73[278], line_72[276], line_71[274], line_70[272], line_69[270], line_68[268], line_67[266], line_66[264], line_65[262], line_64[260], line_63[258], line_62[256], line_61[254], line_60[252], line_59[250], line_58[248], line_57[246], line_56[244], line_55[242], line_54[240], line_53[238], line_52[236], line_51[234], line_50[232], line_49[230], line_48[228], line_47[226], line_46[224], line_45[222], line_44[220], line_43[218], line_42[216], line_41[214], line_40[212], line_39[210], line_38[208], line_37[206], line_36[204], line_35[202], line_34[200], line_33[198], line_32[196], line_31[194], line_30[192], line_29[190], line_28[188], line_27[186], line_26[184], line_25[182], line_24[180], line_23[178], line_22[176], line_21[174], line_20[172], line_19[170], line_18[168], line_17[166], line_16[164], line_15[162], line_14[160], line_13[158], line_12[156], line_11[154], line_10[152], line_9[150], line_8[148], line_7[146], line_6[144], line_5[142], line_4[140], line_3[138], line_2[136], line_1[134] };
assign col_389 = {line_128[389], line_127[387], line_126[385], line_125[383], line_124[381], line_123[379], line_122[377], line_121[375], line_120[373], line_119[371], line_118[369], line_117[367], line_116[365], line_115[363], line_114[361], line_113[359], line_112[357], line_111[355], line_110[353], line_109[351], line_108[349], line_107[347], line_106[345], line_105[343], line_104[341], line_103[339], line_102[337], line_101[335], line_100[333], line_99[331], line_98[329], line_97[327], line_96[325], line_95[323], line_94[321], line_93[319], line_92[317], line_91[315], line_90[313], line_89[311], line_88[309], line_87[307], line_86[305], line_85[303], line_84[301], line_83[299], line_82[297], line_81[295], line_80[293], line_79[291], line_78[289], line_77[287], line_76[285], line_75[283], line_74[281], line_73[279], line_72[277], line_71[275], line_70[273], line_69[271], line_68[269], line_67[267], line_66[265], line_65[263], line_64[261], line_63[259], line_62[257], line_61[255], line_60[253], line_59[251], line_58[249], line_57[247], line_56[245], line_55[243], line_54[241], line_53[239], line_52[237], line_51[235], line_50[233], line_49[231], line_48[229], line_47[227], line_46[225], line_45[223], line_44[221], line_43[219], line_42[217], line_41[215], line_40[213], line_39[211], line_38[209], line_37[207], line_36[205], line_35[203], line_34[201], line_33[199], line_32[197], line_31[195], line_30[193], line_29[191], line_28[189], line_27[187], line_26[185], line_25[183], line_24[181], line_23[179], line_22[177], line_21[175], line_20[173], line_19[171], line_18[169], line_17[167], line_16[165], line_15[163], line_14[161], line_13[159], line_12[157], line_11[155], line_10[153], line_9[151], line_8[149], line_7[147], line_6[145], line_5[143], line_4[141], line_3[139], line_2[137], line_1[135] };
assign col_390 = {line_128[390], line_127[388], line_126[386], line_125[384], line_124[382], line_123[380], line_122[378], line_121[376], line_120[374], line_119[372], line_118[370], line_117[368], line_116[366], line_115[364], line_114[362], line_113[360], line_112[358], line_111[356], line_110[354], line_109[352], line_108[350], line_107[348], line_106[346], line_105[344], line_104[342], line_103[340], line_102[338], line_101[336], line_100[334], line_99[332], line_98[330], line_97[328], line_96[326], line_95[324], line_94[322], line_93[320], line_92[318], line_91[316], line_90[314], line_89[312], line_88[310], line_87[308], line_86[306], line_85[304], line_84[302], line_83[300], line_82[298], line_81[296], line_80[294], line_79[292], line_78[290], line_77[288], line_76[286], line_75[284], line_74[282], line_73[280], line_72[278], line_71[276], line_70[274], line_69[272], line_68[270], line_67[268], line_66[266], line_65[264], line_64[262], line_63[260], line_62[258], line_61[256], line_60[254], line_59[252], line_58[250], line_57[248], line_56[246], line_55[244], line_54[242], line_53[240], line_52[238], line_51[236], line_50[234], line_49[232], line_48[230], line_47[228], line_46[226], line_45[224], line_44[222], line_43[220], line_42[218], line_41[216], line_40[214], line_39[212], line_38[210], line_37[208], line_36[206], line_35[204], line_34[202], line_33[200], line_32[198], line_31[196], line_30[194], line_29[192], line_28[190], line_27[188], line_26[186], line_25[184], line_24[182], line_23[180], line_22[178], line_21[176], line_20[174], line_19[172], line_18[170], line_17[168], line_16[166], line_15[164], line_14[162], line_13[160], line_12[158], line_11[156], line_10[154], line_9[152], line_8[150], line_7[148], line_6[146], line_5[144], line_4[142], line_3[140], line_2[138], line_1[136] };
assign col_391 = {line_128[391], line_127[389], line_126[387], line_125[385], line_124[383], line_123[381], line_122[379], line_121[377], line_120[375], line_119[373], line_118[371], line_117[369], line_116[367], line_115[365], line_114[363], line_113[361], line_112[359], line_111[357], line_110[355], line_109[353], line_108[351], line_107[349], line_106[347], line_105[345], line_104[343], line_103[341], line_102[339], line_101[337], line_100[335], line_99[333], line_98[331], line_97[329], line_96[327], line_95[325], line_94[323], line_93[321], line_92[319], line_91[317], line_90[315], line_89[313], line_88[311], line_87[309], line_86[307], line_85[305], line_84[303], line_83[301], line_82[299], line_81[297], line_80[295], line_79[293], line_78[291], line_77[289], line_76[287], line_75[285], line_74[283], line_73[281], line_72[279], line_71[277], line_70[275], line_69[273], line_68[271], line_67[269], line_66[267], line_65[265], line_64[263], line_63[261], line_62[259], line_61[257], line_60[255], line_59[253], line_58[251], line_57[249], line_56[247], line_55[245], line_54[243], line_53[241], line_52[239], line_51[237], line_50[235], line_49[233], line_48[231], line_47[229], line_46[227], line_45[225], line_44[223], line_43[221], line_42[219], line_41[217], line_40[215], line_39[213], line_38[211], line_37[209], line_36[207], line_35[205], line_34[203], line_33[201], line_32[199], line_31[197], line_30[195], line_29[193], line_28[191], line_27[189], line_26[187], line_25[185], line_24[183], line_23[181], line_22[179], line_21[177], line_20[175], line_19[173], line_18[171], line_17[169], line_16[167], line_15[165], line_14[163], line_13[161], line_12[159], line_11[157], line_10[155], line_9[153], line_8[151], line_7[149], line_6[147], line_5[145], line_4[143], line_3[141], line_2[139], line_1[137] };
assign col_392 = {line_128[392], line_127[390], line_126[388], line_125[386], line_124[384], line_123[382], line_122[380], line_121[378], line_120[376], line_119[374], line_118[372], line_117[370], line_116[368], line_115[366], line_114[364], line_113[362], line_112[360], line_111[358], line_110[356], line_109[354], line_108[352], line_107[350], line_106[348], line_105[346], line_104[344], line_103[342], line_102[340], line_101[338], line_100[336], line_99[334], line_98[332], line_97[330], line_96[328], line_95[326], line_94[324], line_93[322], line_92[320], line_91[318], line_90[316], line_89[314], line_88[312], line_87[310], line_86[308], line_85[306], line_84[304], line_83[302], line_82[300], line_81[298], line_80[296], line_79[294], line_78[292], line_77[290], line_76[288], line_75[286], line_74[284], line_73[282], line_72[280], line_71[278], line_70[276], line_69[274], line_68[272], line_67[270], line_66[268], line_65[266], line_64[264], line_63[262], line_62[260], line_61[258], line_60[256], line_59[254], line_58[252], line_57[250], line_56[248], line_55[246], line_54[244], line_53[242], line_52[240], line_51[238], line_50[236], line_49[234], line_48[232], line_47[230], line_46[228], line_45[226], line_44[224], line_43[222], line_42[220], line_41[218], line_40[216], line_39[214], line_38[212], line_37[210], line_36[208], line_35[206], line_34[204], line_33[202], line_32[200], line_31[198], line_30[196], line_29[194], line_28[192], line_27[190], line_26[188], line_25[186], line_24[184], line_23[182], line_22[180], line_21[178], line_20[176], line_19[174], line_18[172], line_17[170], line_16[168], line_15[166], line_14[164], line_13[162], line_12[160], line_11[158], line_10[156], line_9[154], line_8[152], line_7[150], line_6[148], line_5[146], line_4[144], line_3[142], line_2[140], line_1[138] };
assign col_393 = {line_128[393], line_127[391], line_126[389], line_125[387], line_124[385], line_123[383], line_122[381], line_121[379], line_120[377], line_119[375], line_118[373], line_117[371], line_116[369], line_115[367], line_114[365], line_113[363], line_112[361], line_111[359], line_110[357], line_109[355], line_108[353], line_107[351], line_106[349], line_105[347], line_104[345], line_103[343], line_102[341], line_101[339], line_100[337], line_99[335], line_98[333], line_97[331], line_96[329], line_95[327], line_94[325], line_93[323], line_92[321], line_91[319], line_90[317], line_89[315], line_88[313], line_87[311], line_86[309], line_85[307], line_84[305], line_83[303], line_82[301], line_81[299], line_80[297], line_79[295], line_78[293], line_77[291], line_76[289], line_75[287], line_74[285], line_73[283], line_72[281], line_71[279], line_70[277], line_69[275], line_68[273], line_67[271], line_66[269], line_65[267], line_64[265], line_63[263], line_62[261], line_61[259], line_60[257], line_59[255], line_58[253], line_57[251], line_56[249], line_55[247], line_54[245], line_53[243], line_52[241], line_51[239], line_50[237], line_49[235], line_48[233], line_47[231], line_46[229], line_45[227], line_44[225], line_43[223], line_42[221], line_41[219], line_40[217], line_39[215], line_38[213], line_37[211], line_36[209], line_35[207], line_34[205], line_33[203], line_32[201], line_31[199], line_30[197], line_29[195], line_28[193], line_27[191], line_26[189], line_25[187], line_24[185], line_23[183], line_22[181], line_21[179], line_20[177], line_19[175], line_18[173], line_17[171], line_16[169], line_15[167], line_14[165], line_13[163], line_12[161], line_11[159], line_10[157], line_9[155], line_8[153], line_7[151], line_6[149], line_5[147], line_4[145], line_3[143], line_2[141], line_1[139] };
assign col_394 = {line_128[394], line_127[392], line_126[390], line_125[388], line_124[386], line_123[384], line_122[382], line_121[380], line_120[378], line_119[376], line_118[374], line_117[372], line_116[370], line_115[368], line_114[366], line_113[364], line_112[362], line_111[360], line_110[358], line_109[356], line_108[354], line_107[352], line_106[350], line_105[348], line_104[346], line_103[344], line_102[342], line_101[340], line_100[338], line_99[336], line_98[334], line_97[332], line_96[330], line_95[328], line_94[326], line_93[324], line_92[322], line_91[320], line_90[318], line_89[316], line_88[314], line_87[312], line_86[310], line_85[308], line_84[306], line_83[304], line_82[302], line_81[300], line_80[298], line_79[296], line_78[294], line_77[292], line_76[290], line_75[288], line_74[286], line_73[284], line_72[282], line_71[280], line_70[278], line_69[276], line_68[274], line_67[272], line_66[270], line_65[268], line_64[266], line_63[264], line_62[262], line_61[260], line_60[258], line_59[256], line_58[254], line_57[252], line_56[250], line_55[248], line_54[246], line_53[244], line_52[242], line_51[240], line_50[238], line_49[236], line_48[234], line_47[232], line_46[230], line_45[228], line_44[226], line_43[224], line_42[222], line_41[220], line_40[218], line_39[216], line_38[214], line_37[212], line_36[210], line_35[208], line_34[206], line_33[204], line_32[202], line_31[200], line_30[198], line_29[196], line_28[194], line_27[192], line_26[190], line_25[188], line_24[186], line_23[184], line_22[182], line_21[180], line_20[178], line_19[176], line_18[174], line_17[172], line_16[170], line_15[168], line_14[166], line_13[164], line_12[162], line_11[160], line_10[158], line_9[156], line_8[154], line_7[152], line_6[150], line_5[148], line_4[146], line_3[144], line_2[142], line_1[140] };
assign col_395 = {line_128[395], line_127[393], line_126[391], line_125[389], line_124[387], line_123[385], line_122[383], line_121[381], line_120[379], line_119[377], line_118[375], line_117[373], line_116[371], line_115[369], line_114[367], line_113[365], line_112[363], line_111[361], line_110[359], line_109[357], line_108[355], line_107[353], line_106[351], line_105[349], line_104[347], line_103[345], line_102[343], line_101[341], line_100[339], line_99[337], line_98[335], line_97[333], line_96[331], line_95[329], line_94[327], line_93[325], line_92[323], line_91[321], line_90[319], line_89[317], line_88[315], line_87[313], line_86[311], line_85[309], line_84[307], line_83[305], line_82[303], line_81[301], line_80[299], line_79[297], line_78[295], line_77[293], line_76[291], line_75[289], line_74[287], line_73[285], line_72[283], line_71[281], line_70[279], line_69[277], line_68[275], line_67[273], line_66[271], line_65[269], line_64[267], line_63[265], line_62[263], line_61[261], line_60[259], line_59[257], line_58[255], line_57[253], line_56[251], line_55[249], line_54[247], line_53[245], line_52[243], line_51[241], line_50[239], line_49[237], line_48[235], line_47[233], line_46[231], line_45[229], line_44[227], line_43[225], line_42[223], line_41[221], line_40[219], line_39[217], line_38[215], line_37[213], line_36[211], line_35[209], line_34[207], line_33[205], line_32[203], line_31[201], line_30[199], line_29[197], line_28[195], line_27[193], line_26[191], line_25[189], line_24[187], line_23[185], line_22[183], line_21[181], line_20[179], line_19[177], line_18[175], line_17[173], line_16[171], line_15[169], line_14[167], line_13[165], line_12[163], line_11[161], line_10[159], line_9[157], line_8[155], line_7[153], line_6[151], line_5[149], line_4[147], line_3[145], line_2[143], line_1[141] };
assign col_396 = {line_128[396], line_127[394], line_126[392], line_125[390], line_124[388], line_123[386], line_122[384], line_121[382], line_120[380], line_119[378], line_118[376], line_117[374], line_116[372], line_115[370], line_114[368], line_113[366], line_112[364], line_111[362], line_110[360], line_109[358], line_108[356], line_107[354], line_106[352], line_105[350], line_104[348], line_103[346], line_102[344], line_101[342], line_100[340], line_99[338], line_98[336], line_97[334], line_96[332], line_95[330], line_94[328], line_93[326], line_92[324], line_91[322], line_90[320], line_89[318], line_88[316], line_87[314], line_86[312], line_85[310], line_84[308], line_83[306], line_82[304], line_81[302], line_80[300], line_79[298], line_78[296], line_77[294], line_76[292], line_75[290], line_74[288], line_73[286], line_72[284], line_71[282], line_70[280], line_69[278], line_68[276], line_67[274], line_66[272], line_65[270], line_64[268], line_63[266], line_62[264], line_61[262], line_60[260], line_59[258], line_58[256], line_57[254], line_56[252], line_55[250], line_54[248], line_53[246], line_52[244], line_51[242], line_50[240], line_49[238], line_48[236], line_47[234], line_46[232], line_45[230], line_44[228], line_43[226], line_42[224], line_41[222], line_40[220], line_39[218], line_38[216], line_37[214], line_36[212], line_35[210], line_34[208], line_33[206], line_32[204], line_31[202], line_30[200], line_29[198], line_28[196], line_27[194], line_26[192], line_25[190], line_24[188], line_23[186], line_22[184], line_21[182], line_20[180], line_19[178], line_18[176], line_17[174], line_16[172], line_15[170], line_14[168], line_13[166], line_12[164], line_11[162], line_10[160], line_9[158], line_8[156], line_7[154], line_6[152], line_5[150], line_4[148], line_3[146], line_2[144], line_1[142] };
assign col_397 = {line_128[397], line_127[395], line_126[393], line_125[391], line_124[389], line_123[387], line_122[385], line_121[383], line_120[381], line_119[379], line_118[377], line_117[375], line_116[373], line_115[371], line_114[369], line_113[367], line_112[365], line_111[363], line_110[361], line_109[359], line_108[357], line_107[355], line_106[353], line_105[351], line_104[349], line_103[347], line_102[345], line_101[343], line_100[341], line_99[339], line_98[337], line_97[335], line_96[333], line_95[331], line_94[329], line_93[327], line_92[325], line_91[323], line_90[321], line_89[319], line_88[317], line_87[315], line_86[313], line_85[311], line_84[309], line_83[307], line_82[305], line_81[303], line_80[301], line_79[299], line_78[297], line_77[295], line_76[293], line_75[291], line_74[289], line_73[287], line_72[285], line_71[283], line_70[281], line_69[279], line_68[277], line_67[275], line_66[273], line_65[271], line_64[269], line_63[267], line_62[265], line_61[263], line_60[261], line_59[259], line_58[257], line_57[255], line_56[253], line_55[251], line_54[249], line_53[247], line_52[245], line_51[243], line_50[241], line_49[239], line_48[237], line_47[235], line_46[233], line_45[231], line_44[229], line_43[227], line_42[225], line_41[223], line_40[221], line_39[219], line_38[217], line_37[215], line_36[213], line_35[211], line_34[209], line_33[207], line_32[205], line_31[203], line_30[201], line_29[199], line_28[197], line_27[195], line_26[193], line_25[191], line_24[189], line_23[187], line_22[185], line_21[183], line_20[181], line_19[179], line_18[177], line_17[175], line_16[173], line_15[171], line_14[169], line_13[167], line_12[165], line_11[163], line_10[161], line_9[159], line_8[157], line_7[155], line_6[153], line_5[151], line_4[149], line_3[147], line_2[145], line_1[143] };
assign col_398 = {line_128[398], line_127[396], line_126[394], line_125[392], line_124[390], line_123[388], line_122[386], line_121[384], line_120[382], line_119[380], line_118[378], line_117[376], line_116[374], line_115[372], line_114[370], line_113[368], line_112[366], line_111[364], line_110[362], line_109[360], line_108[358], line_107[356], line_106[354], line_105[352], line_104[350], line_103[348], line_102[346], line_101[344], line_100[342], line_99[340], line_98[338], line_97[336], line_96[334], line_95[332], line_94[330], line_93[328], line_92[326], line_91[324], line_90[322], line_89[320], line_88[318], line_87[316], line_86[314], line_85[312], line_84[310], line_83[308], line_82[306], line_81[304], line_80[302], line_79[300], line_78[298], line_77[296], line_76[294], line_75[292], line_74[290], line_73[288], line_72[286], line_71[284], line_70[282], line_69[280], line_68[278], line_67[276], line_66[274], line_65[272], line_64[270], line_63[268], line_62[266], line_61[264], line_60[262], line_59[260], line_58[258], line_57[256], line_56[254], line_55[252], line_54[250], line_53[248], line_52[246], line_51[244], line_50[242], line_49[240], line_48[238], line_47[236], line_46[234], line_45[232], line_44[230], line_43[228], line_42[226], line_41[224], line_40[222], line_39[220], line_38[218], line_37[216], line_36[214], line_35[212], line_34[210], line_33[208], line_32[206], line_31[204], line_30[202], line_29[200], line_28[198], line_27[196], line_26[194], line_25[192], line_24[190], line_23[188], line_22[186], line_21[184], line_20[182], line_19[180], line_18[178], line_17[176], line_16[174], line_15[172], line_14[170], line_13[168], line_12[166], line_11[164], line_10[162], line_9[160], line_8[158], line_7[156], line_6[154], line_5[152], line_4[150], line_3[148], line_2[146], line_1[144] };
assign col_399 = {line_128[399], line_127[397], line_126[395], line_125[393], line_124[391], line_123[389], line_122[387], line_121[385], line_120[383], line_119[381], line_118[379], line_117[377], line_116[375], line_115[373], line_114[371], line_113[369], line_112[367], line_111[365], line_110[363], line_109[361], line_108[359], line_107[357], line_106[355], line_105[353], line_104[351], line_103[349], line_102[347], line_101[345], line_100[343], line_99[341], line_98[339], line_97[337], line_96[335], line_95[333], line_94[331], line_93[329], line_92[327], line_91[325], line_90[323], line_89[321], line_88[319], line_87[317], line_86[315], line_85[313], line_84[311], line_83[309], line_82[307], line_81[305], line_80[303], line_79[301], line_78[299], line_77[297], line_76[295], line_75[293], line_74[291], line_73[289], line_72[287], line_71[285], line_70[283], line_69[281], line_68[279], line_67[277], line_66[275], line_65[273], line_64[271], line_63[269], line_62[267], line_61[265], line_60[263], line_59[261], line_58[259], line_57[257], line_56[255], line_55[253], line_54[251], line_53[249], line_52[247], line_51[245], line_50[243], line_49[241], line_48[239], line_47[237], line_46[235], line_45[233], line_44[231], line_43[229], line_42[227], line_41[225], line_40[223], line_39[221], line_38[219], line_37[217], line_36[215], line_35[213], line_34[211], line_33[209], line_32[207], line_31[205], line_30[203], line_29[201], line_28[199], line_27[197], line_26[195], line_25[193], line_24[191], line_23[189], line_22[187], line_21[185], line_20[183], line_19[181], line_18[179], line_17[177], line_16[175], line_15[173], line_14[171], line_13[169], line_12[167], line_11[165], line_10[163], line_9[161], line_8[159], line_7[157], line_6[155], line_5[153], line_4[151], line_3[149], line_2[147], line_1[145] };
assign col_400 = {line_128[400], line_127[398], line_126[396], line_125[394], line_124[392], line_123[390], line_122[388], line_121[386], line_120[384], line_119[382], line_118[380], line_117[378], line_116[376], line_115[374], line_114[372], line_113[370], line_112[368], line_111[366], line_110[364], line_109[362], line_108[360], line_107[358], line_106[356], line_105[354], line_104[352], line_103[350], line_102[348], line_101[346], line_100[344], line_99[342], line_98[340], line_97[338], line_96[336], line_95[334], line_94[332], line_93[330], line_92[328], line_91[326], line_90[324], line_89[322], line_88[320], line_87[318], line_86[316], line_85[314], line_84[312], line_83[310], line_82[308], line_81[306], line_80[304], line_79[302], line_78[300], line_77[298], line_76[296], line_75[294], line_74[292], line_73[290], line_72[288], line_71[286], line_70[284], line_69[282], line_68[280], line_67[278], line_66[276], line_65[274], line_64[272], line_63[270], line_62[268], line_61[266], line_60[264], line_59[262], line_58[260], line_57[258], line_56[256], line_55[254], line_54[252], line_53[250], line_52[248], line_51[246], line_50[244], line_49[242], line_48[240], line_47[238], line_46[236], line_45[234], line_44[232], line_43[230], line_42[228], line_41[226], line_40[224], line_39[222], line_38[220], line_37[218], line_36[216], line_35[214], line_34[212], line_33[210], line_32[208], line_31[206], line_30[204], line_29[202], line_28[200], line_27[198], line_26[196], line_25[194], line_24[192], line_23[190], line_22[188], line_21[186], line_20[184], line_19[182], line_18[180], line_17[178], line_16[176], line_15[174], line_14[172], line_13[170], line_12[168], line_11[166], line_10[164], line_9[162], line_8[160], line_7[158], line_6[156], line_5[154], line_4[152], line_3[150], line_2[148], line_1[146] };
assign col_401 = {line_128[401], line_127[399], line_126[397], line_125[395], line_124[393], line_123[391], line_122[389], line_121[387], line_120[385], line_119[383], line_118[381], line_117[379], line_116[377], line_115[375], line_114[373], line_113[371], line_112[369], line_111[367], line_110[365], line_109[363], line_108[361], line_107[359], line_106[357], line_105[355], line_104[353], line_103[351], line_102[349], line_101[347], line_100[345], line_99[343], line_98[341], line_97[339], line_96[337], line_95[335], line_94[333], line_93[331], line_92[329], line_91[327], line_90[325], line_89[323], line_88[321], line_87[319], line_86[317], line_85[315], line_84[313], line_83[311], line_82[309], line_81[307], line_80[305], line_79[303], line_78[301], line_77[299], line_76[297], line_75[295], line_74[293], line_73[291], line_72[289], line_71[287], line_70[285], line_69[283], line_68[281], line_67[279], line_66[277], line_65[275], line_64[273], line_63[271], line_62[269], line_61[267], line_60[265], line_59[263], line_58[261], line_57[259], line_56[257], line_55[255], line_54[253], line_53[251], line_52[249], line_51[247], line_50[245], line_49[243], line_48[241], line_47[239], line_46[237], line_45[235], line_44[233], line_43[231], line_42[229], line_41[227], line_40[225], line_39[223], line_38[221], line_37[219], line_36[217], line_35[215], line_34[213], line_33[211], line_32[209], line_31[207], line_30[205], line_29[203], line_28[201], line_27[199], line_26[197], line_25[195], line_24[193], line_23[191], line_22[189], line_21[187], line_20[185], line_19[183], line_18[181], line_17[179], line_16[177], line_15[175], line_14[173], line_13[171], line_12[169], line_11[167], line_10[165], line_9[163], line_8[161], line_7[159], line_6[157], line_5[155], line_4[153], line_3[151], line_2[149], line_1[147] };
assign col_402 = {line_128[402], line_127[400], line_126[398], line_125[396], line_124[394], line_123[392], line_122[390], line_121[388], line_120[386], line_119[384], line_118[382], line_117[380], line_116[378], line_115[376], line_114[374], line_113[372], line_112[370], line_111[368], line_110[366], line_109[364], line_108[362], line_107[360], line_106[358], line_105[356], line_104[354], line_103[352], line_102[350], line_101[348], line_100[346], line_99[344], line_98[342], line_97[340], line_96[338], line_95[336], line_94[334], line_93[332], line_92[330], line_91[328], line_90[326], line_89[324], line_88[322], line_87[320], line_86[318], line_85[316], line_84[314], line_83[312], line_82[310], line_81[308], line_80[306], line_79[304], line_78[302], line_77[300], line_76[298], line_75[296], line_74[294], line_73[292], line_72[290], line_71[288], line_70[286], line_69[284], line_68[282], line_67[280], line_66[278], line_65[276], line_64[274], line_63[272], line_62[270], line_61[268], line_60[266], line_59[264], line_58[262], line_57[260], line_56[258], line_55[256], line_54[254], line_53[252], line_52[250], line_51[248], line_50[246], line_49[244], line_48[242], line_47[240], line_46[238], line_45[236], line_44[234], line_43[232], line_42[230], line_41[228], line_40[226], line_39[224], line_38[222], line_37[220], line_36[218], line_35[216], line_34[214], line_33[212], line_32[210], line_31[208], line_30[206], line_29[204], line_28[202], line_27[200], line_26[198], line_25[196], line_24[194], line_23[192], line_22[190], line_21[188], line_20[186], line_19[184], line_18[182], line_17[180], line_16[178], line_15[176], line_14[174], line_13[172], line_12[170], line_11[168], line_10[166], line_9[164], line_8[162], line_7[160], line_6[158], line_5[156], line_4[154], line_3[152], line_2[150], line_1[148] };
assign col_403 = {line_128[403], line_127[401], line_126[399], line_125[397], line_124[395], line_123[393], line_122[391], line_121[389], line_120[387], line_119[385], line_118[383], line_117[381], line_116[379], line_115[377], line_114[375], line_113[373], line_112[371], line_111[369], line_110[367], line_109[365], line_108[363], line_107[361], line_106[359], line_105[357], line_104[355], line_103[353], line_102[351], line_101[349], line_100[347], line_99[345], line_98[343], line_97[341], line_96[339], line_95[337], line_94[335], line_93[333], line_92[331], line_91[329], line_90[327], line_89[325], line_88[323], line_87[321], line_86[319], line_85[317], line_84[315], line_83[313], line_82[311], line_81[309], line_80[307], line_79[305], line_78[303], line_77[301], line_76[299], line_75[297], line_74[295], line_73[293], line_72[291], line_71[289], line_70[287], line_69[285], line_68[283], line_67[281], line_66[279], line_65[277], line_64[275], line_63[273], line_62[271], line_61[269], line_60[267], line_59[265], line_58[263], line_57[261], line_56[259], line_55[257], line_54[255], line_53[253], line_52[251], line_51[249], line_50[247], line_49[245], line_48[243], line_47[241], line_46[239], line_45[237], line_44[235], line_43[233], line_42[231], line_41[229], line_40[227], line_39[225], line_38[223], line_37[221], line_36[219], line_35[217], line_34[215], line_33[213], line_32[211], line_31[209], line_30[207], line_29[205], line_28[203], line_27[201], line_26[199], line_25[197], line_24[195], line_23[193], line_22[191], line_21[189], line_20[187], line_19[185], line_18[183], line_17[181], line_16[179], line_15[177], line_14[175], line_13[173], line_12[171], line_11[169], line_10[167], line_9[165], line_8[163], line_7[161], line_6[159], line_5[157], line_4[155], line_3[153], line_2[151], line_1[149] };
assign col_404 = {line_128[404], line_127[402], line_126[400], line_125[398], line_124[396], line_123[394], line_122[392], line_121[390], line_120[388], line_119[386], line_118[384], line_117[382], line_116[380], line_115[378], line_114[376], line_113[374], line_112[372], line_111[370], line_110[368], line_109[366], line_108[364], line_107[362], line_106[360], line_105[358], line_104[356], line_103[354], line_102[352], line_101[350], line_100[348], line_99[346], line_98[344], line_97[342], line_96[340], line_95[338], line_94[336], line_93[334], line_92[332], line_91[330], line_90[328], line_89[326], line_88[324], line_87[322], line_86[320], line_85[318], line_84[316], line_83[314], line_82[312], line_81[310], line_80[308], line_79[306], line_78[304], line_77[302], line_76[300], line_75[298], line_74[296], line_73[294], line_72[292], line_71[290], line_70[288], line_69[286], line_68[284], line_67[282], line_66[280], line_65[278], line_64[276], line_63[274], line_62[272], line_61[270], line_60[268], line_59[266], line_58[264], line_57[262], line_56[260], line_55[258], line_54[256], line_53[254], line_52[252], line_51[250], line_50[248], line_49[246], line_48[244], line_47[242], line_46[240], line_45[238], line_44[236], line_43[234], line_42[232], line_41[230], line_40[228], line_39[226], line_38[224], line_37[222], line_36[220], line_35[218], line_34[216], line_33[214], line_32[212], line_31[210], line_30[208], line_29[206], line_28[204], line_27[202], line_26[200], line_25[198], line_24[196], line_23[194], line_22[192], line_21[190], line_20[188], line_19[186], line_18[184], line_17[182], line_16[180], line_15[178], line_14[176], line_13[174], line_12[172], line_11[170], line_10[168], line_9[166], line_8[164], line_7[162], line_6[160], line_5[158], line_4[156], line_3[154], line_2[152], line_1[150] };
assign col_405 = {line_128[405], line_127[403], line_126[401], line_125[399], line_124[397], line_123[395], line_122[393], line_121[391], line_120[389], line_119[387], line_118[385], line_117[383], line_116[381], line_115[379], line_114[377], line_113[375], line_112[373], line_111[371], line_110[369], line_109[367], line_108[365], line_107[363], line_106[361], line_105[359], line_104[357], line_103[355], line_102[353], line_101[351], line_100[349], line_99[347], line_98[345], line_97[343], line_96[341], line_95[339], line_94[337], line_93[335], line_92[333], line_91[331], line_90[329], line_89[327], line_88[325], line_87[323], line_86[321], line_85[319], line_84[317], line_83[315], line_82[313], line_81[311], line_80[309], line_79[307], line_78[305], line_77[303], line_76[301], line_75[299], line_74[297], line_73[295], line_72[293], line_71[291], line_70[289], line_69[287], line_68[285], line_67[283], line_66[281], line_65[279], line_64[277], line_63[275], line_62[273], line_61[271], line_60[269], line_59[267], line_58[265], line_57[263], line_56[261], line_55[259], line_54[257], line_53[255], line_52[253], line_51[251], line_50[249], line_49[247], line_48[245], line_47[243], line_46[241], line_45[239], line_44[237], line_43[235], line_42[233], line_41[231], line_40[229], line_39[227], line_38[225], line_37[223], line_36[221], line_35[219], line_34[217], line_33[215], line_32[213], line_31[211], line_30[209], line_29[207], line_28[205], line_27[203], line_26[201], line_25[199], line_24[197], line_23[195], line_22[193], line_21[191], line_20[189], line_19[187], line_18[185], line_17[183], line_16[181], line_15[179], line_14[177], line_13[175], line_12[173], line_11[171], line_10[169], line_9[167], line_8[165], line_7[163], line_6[161], line_5[159], line_4[157], line_3[155], line_2[153], line_1[151] };
assign col_406 = {line_128[406], line_127[404], line_126[402], line_125[400], line_124[398], line_123[396], line_122[394], line_121[392], line_120[390], line_119[388], line_118[386], line_117[384], line_116[382], line_115[380], line_114[378], line_113[376], line_112[374], line_111[372], line_110[370], line_109[368], line_108[366], line_107[364], line_106[362], line_105[360], line_104[358], line_103[356], line_102[354], line_101[352], line_100[350], line_99[348], line_98[346], line_97[344], line_96[342], line_95[340], line_94[338], line_93[336], line_92[334], line_91[332], line_90[330], line_89[328], line_88[326], line_87[324], line_86[322], line_85[320], line_84[318], line_83[316], line_82[314], line_81[312], line_80[310], line_79[308], line_78[306], line_77[304], line_76[302], line_75[300], line_74[298], line_73[296], line_72[294], line_71[292], line_70[290], line_69[288], line_68[286], line_67[284], line_66[282], line_65[280], line_64[278], line_63[276], line_62[274], line_61[272], line_60[270], line_59[268], line_58[266], line_57[264], line_56[262], line_55[260], line_54[258], line_53[256], line_52[254], line_51[252], line_50[250], line_49[248], line_48[246], line_47[244], line_46[242], line_45[240], line_44[238], line_43[236], line_42[234], line_41[232], line_40[230], line_39[228], line_38[226], line_37[224], line_36[222], line_35[220], line_34[218], line_33[216], line_32[214], line_31[212], line_30[210], line_29[208], line_28[206], line_27[204], line_26[202], line_25[200], line_24[198], line_23[196], line_22[194], line_21[192], line_20[190], line_19[188], line_18[186], line_17[184], line_16[182], line_15[180], line_14[178], line_13[176], line_12[174], line_11[172], line_10[170], line_9[168], line_8[166], line_7[164], line_6[162], line_5[160], line_4[158], line_3[156], line_2[154], line_1[152] };
assign col_407 = {line_128[407], line_127[405], line_126[403], line_125[401], line_124[399], line_123[397], line_122[395], line_121[393], line_120[391], line_119[389], line_118[387], line_117[385], line_116[383], line_115[381], line_114[379], line_113[377], line_112[375], line_111[373], line_110[371], line_109[369], line_108[367], line_107[365], line_106[363], line_105[361], line_104[359], line_103[357], line_102[355], line_101[353], line_100[351], line_99[349], line_98[347], line_97[345], line_96[343], line_95[341], line_94[339], line_93[337], line_92[335], line_91[333], line_90[331], line_89[329], line_88[327], line_87[325], line_86[323], line_85[321], line_84[319], line_83[317], line_82[315], line_81[313], line_80[311], line_79[309], line_78[307], line_77[305], line_76[303], line_75[301], line_74[299], line_73[297], line_72[295], line_71[293], line_70[291], line_69[289], line_68[287], line_67[285], line_66[283], line_65[281], line_64[279], line_63[277], line_62[275], line_61[273], line_60[271], line_59[269], line_58[267], line_57[265], line_56[263], line_55[261], line_54[259], line_53[257], line_52[255], line_51[253], line_50[251], line_49[249], line_48[247], line_47[245], line_46[243], line_45[241], line_44[239], line_43[237], line_42[235], line_41[233], line_40[231], line_39[229], line_38[227], line_37[225], line_36[223], line_35[221], line_34[219], line_33[217], line_32[215], line_31[213], line_30[211], line_29[209], line_28[207], line_27[205], line_26[203], line_25[201], line_24[199], line_23[197], line_22[195], line_21[193], line_20[191], line_19[189], line_18[187], line_17[185], line_16[183], line_15[181], line_14[179], line_13[177], line_12[175], line_11[173], line_10[171], line_9[169], line_8[167], line_7[165], line_6[163], line_5[161], line_4[159], line_3[157], line_2[155], line_1[153] };
assign col_408 = {line_128[408], line_127[406], line_126[404], line_125[402], line_124[400], line_123[398], line_122[396], line_121[394], line_120[392], line_119[390], line_118[388], line_117[386], line_116[384], line_115[382], line_114[380], line_113[378], line_112[376], line_111[374], line_110[372], line_109[370], line_108[368], line_107[366], line_106[364], line_105[362], line_104[360], line_103[358], line_102[356], line_101[354], line_100[352], line_99[350], line_98[348], line_97[346], line_96[344], line_95[342], line_94[340], line_93[338], line_92[336], line_91[334], line_90[332], line_89[330], line_88[328], line_87[326], line_86[324], line_85[322], line_84[320], line_83[318], line_82[316], line_81[314], line_80[312], line_79[310], line_78[308], line_77[306], line_76[304], line_75[302], line_74[300], line_73[298], line_72[296], line_71[294], line_70[292], line_69[290], line_68[288], line_67[286], line_66[284], line_65[282], line_64[280], line_63[278], line_62[276], line_61[274], line_60[272], line_59[270], line_58[268], line_57[266], line_56[264], line_55[262], line_54[260], line_53[258], line_52[256], line_51[254], line_50[252], line_49[250], line_48[248], line_47[246], line_46[244], line_45[242], line_44[240], line_43[238], line_42[236], line_41[234], line_40[232], line_39[230], line_38[228], line_37[226], line_36[224], line_35[222], line_34[220], line_33[218], line_32[216], line_31[214], line_30[212], line_29[210], line_28[208], line_27[206], line_26[204], line_25[202], line_24[200], line_23[198], line_22[196], line_21[194], line_20[192], line_19[190], line_18[188], line_17[186], line_16[184], line_15[182], line_14[180], line_13[178], line_12[176], line_11[174], line_10[172], line_9[170], line_8[168], line_7[166], line_6[164], line_5[162], line_4[160], line_3[158], line_2[156], line_1[154] };
assign col_409 = {line_128[409], line_127[407], line_126[405], line_125[403], line_124[401], line_123[399], line_122[397], line_121[395], line_120[393], line_119[391], line_118[389], line_117[387], line_116[385], line_115[383], line_114[381], line_113[379], line_112[377], line_111[375], line_110[373], line_109[371], line_108[369], line_107[367], line_106[365], line_105[363], line_104[361], line_103[359], line_102[357], line_101[355], line_100[353], line_99[351], line_98[349], line_97[347], line_96[345], line_95[343], line_94[341], line_93[339], line_92[337], line_91[335], line_90[333], line_89[331], line_88[329], line_87[327], line_86[325], line_85[323], line_84[321], line_83[319], line_82[317], line_81[315], line_80[313], line_79[311], line_78[309], line_77[307], line_76[305], line_75[303], line_74[301], line_73[299], line_72[297], line_71[295], line_70[293], line_69[291], line_68[289], line_67[287], line_66[285], line_65[283], line_64[281], line_63[279], line_62[277], line_61[275], line_60[273], line_59[271], line_58[269], line_57[267], line_56[265], line_55[263], line_54[261], line_53[259], line_52[257], line_51[255], line_50[253], line_49[251], line_48[249], line_47[247], line_46[245], line_45[243], line_44[241], line_43[239], line_42[237], line_41[235], line_40[233], line_39[231], line_38[229], line_37[227], line_36[225], line_35[223], line_34[221], line_33[219], line_32[217], line_31[215], line_30[213], line_29[211], line_28[209], line_27[207], line_26[205], line_25[203], line_24[201], line_23[199], line_22[197], line_21[195], line_20[193], line_19[191], line_18[189], line_17[187], line_16[185], line_15[183], line_14[181], line_13[179], line_12[177], line_11[175], line_10[173], line_9[171], line_8[169], line_7[167], line_6[165], line_5[163], line_4[161], line_3[159], line_2[157], line_1[155] };
assign col_410 = {line_128[410], line_127[408], line_126[406], line_125[404], line_124[402], line_123[400], line_122[398], line_121[396], line_120[394], line_119[392], line_118[390], line_117[388], line_116[386], line_115[384], line_114[382], line_113[380], line_112[378], line_111[376], line_110[374], line_109[372], line_108[370], line_107[368], line_106[366], line_105[364], line_104[362], line_103[360], line_102[358], line_101[356], line_100[354], line_99[352], line_98[350], line_97[348], line_96[346], line_95[344], line_94[342], line_93[340], line_92[338], line_91[336], line_90[334], line_89[332], line_88[330], line_87[328], line_86[326], line_85[324], line_84[322], line_83[320], line_82[318], line_81[316], line_80[314], line_79[312], line_78[310], line_77[308], line_76[306], line_75[304], line_74[302], line_73[300], line_72[298], line_71[296], line_70[294], line_69[292], line_68[290], line_67[288], line_66[286], line_65[284], line_64[282], line_63[280], line_62[278], line_61[276], line_60[274], line_59[272], line_58[270], line_57[268], line_56[266], line_55[264], line_54[262], line_53[260], line_52[258], line_51[256], line_50[254], line_49[252], line_48[250], line_47[248], line_46[246], line_45[244], line_44[242], line_43[240], line_42[238], line_41[236], line_40[234], line_39[232], line_38[230], line_37[228], line_36[226], line_35[224], line_34[222], line_33[220], line_32[218], line_31[216], line_30[214], line_29[212], line_28[210], line_27[208], line_26[206], line_25[204], line_24[202], line_23[200], line_22[198], line_21[196], line_20[194], line_19[192], line_18[190], line_17[188], line_16[186], line_15[184], line_14[182], line_13[180], line_12[178], line_11[176], line_10[174], line_9[172], line_8[170], line_7[168], line_6[166], line_5[164], line_4[162], line_3[160], line_2[158], line_1[156] };
assign col_411 = {line_128[411], line_127[409], line_126[407], line_125[405], line_124[403], line_123[401], line_122[399], line_121[397], line_120[395], line_119[393], line_118[391], line_117[389], line_116[387], line_115[385], line_114[383], line_113[381], line_112[379], line_111[377], line_110[375], line_109[373], line_108[371], line_107[369], line_106[367], line_105[365], line_104[363], line_103[361], line_102[359], line_101[357], line_100[355], line_99[353], line_98[351], line_97[349], line_96[347], line_95[345], line_94[343], line_93[341], line_92[339], line_91[337], line_90[335], line_89[333], line_88[331], line_87[329], line_86[327], line_85[325], line_84[323], line_83[321], line_82[319], line_81[317], line_80[315], line_79[313], line_78[311], line_77[309], line_76[307], line_75[305], line_74[303], line_73[301], line_72[299], line_71[297], line_70[295], line_69[293], line_68[291], line_67[289], line_66[287], line_65[285], line_64[283], line_63[281], line_62[279], line_61[277], line_60[275], line_59[273], line_58[271], line_57[269], line_56[267], line_55[265], line_54[263], line_53[261], line_52[259], line_51[257], line_50[255], line_49[253], line_48[251], line_47[249], line_46[247], line_45[245], line_44[243], line_43[241], line_42[239], line_41[237], line_40[235], line_39[233], line_38[231], line_37[229], line_36[227], line_35[225], line_34[223], line_33[221], line_32[219], line_31[217], line_30[215], line_29[213], line_28[211], line_27[209], line_26[207], line_25[205], line_24[203], line_23[201], line_22[199], line_21[197], line_20[195], line_19[193], line_18[191], line_17[189], line_16[187], line_15[185], line_14[183], line_13[181], line_12[179], line_11[177], line_10[175], line_9[173], line_8[171], line_7[169], line_6[167], line_5[165], line_4[163], line_3[161], line_2[159], line_1[157] };
assign col_412 = {line_128[412], line_127[410], line_126[408], line_125[406], line_124[404], line_123[402], line_122[400], line_121[398], line_120[396], line_119[394], line_118[392], line_117[390], line_116[388], line_115[386], line_114[384], line_113[382], line_112[380], line_111[378], line_110[376], line_109[374], line_108[372], line_107[370], line_106[368], line_105[366], line_104[364], line_103[362], line_102[360], line_101[358], line_100[356], line_99[354], line_98[352], line_97[350], line_96[348], line_95[346], line_94[344], line_93[342], line_92[340], line_91[338], line_90[336], line_89[334], line_88[332], line_87[330], line_86[328], line_85[326], line_84[324], line_83[322], line_82[320], line_81[318], line_80[316], line_79[314], line_78[312], line_77[310], line_76[308], line_75[306], line_74[304], line_73[302], line_72[300], line_71[298], line_70[296], line_69[294], line_68[292], line_67[290], line_66[288], line_65[286], line_64[284], line_63[282], line_62[280], line_61[278], line_60[276], line_59[274], line_58[272], line_57[270], line_56[268], line_55[266], line_54[264], line_53[262], line_52[260], line_51[258], line_50[256], line_49[254], line_48[252], line_47[250], line_46[248], line_45[246], line_44[244], line_43[242], line_42[240], line_41[238], line_40[236], line_39[234], line_38[232], line_37[230], line_36[228], line_35[226], line_34[224], line_33[222], line_32[220], line_31[218], line_30[216], line_29[214], line_28[212], line_27[210], line_26[208], line_25[206], line_24[204], line_23[202], line_22[200], line_21[198], line_20[196], line_19[194], line_18[192], line_17[190], line_16[188], line_15[186], line_14[184], line_13[182], line_12[180], line_11[178], line_10[176], line_9[174], line_8[172], line_7[170], line_6[168], line_5[166], line_4[164], line_3[162], line_2[160], line_1[158] };
assign col_413 = {line_128[413], line_127[411], line_126[409], line_125[407], line_124[405], line_123[403], line_122[401], line_121[399], line_120[397], line_119[395], line_118[393], line_117[391], line_116[389], line_115[387], line_114[385], line_113[383], line_112[381], line_111[379], line_110[377], line_109[375], line_108[373], line_107[371], line_106[369], line_105[367], line_104[365], line_103[363], line_102[361], line_101[359], line_100[357], line_99[355], line_98[353], line_97[351], line_96[349], line_95[347], line_94[345], line_93[343], line_92[341], line_91[339], line_90[337], line_89[335], line_88[333], line_87[331], line_86[329], line_85[327], line_84[325], line_83[323], line_82[321], line_81[319], line_80[317], line_79[315], line_78[313], line_77[311], line_76[309], line_75[307], line_74[305], line_73[303], line_72[301], line_71[299], line_70[297], line_69[295], line_68[293], line_67[291], line_66[289], line_65[287], line_64[285], line_63[283], line_62[281], line_61[279], line_60[277], line_59[275], line_58[273], line_57[271], line_56[269], line_55[267], line_54[265], line_53[263], line_52[261], line_51[259], line_50[257], line_49[255], line_48[253], line_47[251], line_46[249], line_45[247], line_44[245], line_43[243], line_42[241], line_41[239], line_40[237], line_39[235], line_38[233], line_37[231], line_36[229], line_35[227], line_34[225], line_33[223], line_32[221], line_31[219], line_30[217], line_29[215], line_28[213], line_27[211], line_26[209], line_25[207], line_24[205], line_23[203], line_22[201], line_21[199], line_20[197], line_19[195], line_18[193], line_17[191], line_16[189], line_15[187], line_14[185], line_13[183], line_12[181], line_11[179], line_10[177], line_9[175], line_8[173], line_7[171], line_6[169], line_5[167], line_4[165], line_3[163], line_2[161], line_1[159] };
assign col_414 = {line_128[414], line_127[412], line_126[410], line_125[408], line_124[406], line_123[404], line_122[402], line_121[400], line_120[398], line_119[396], line_118[394], line_117[392], line_116[390], line_115[388], line_114[386], line_113[384], line_112[382], line_111[380], line_110[378], line_109[376], line_108[374], line_107[372], line_106[370], line_105[368], line_104[366], line_103[364], line_102[362], line_101[360], line_100[358], line_99[356], line_98[354], line_97[352], line_96[350], line_95[348], line_94[346], line_93[344], line_92[342], line_91[340], line_90[338], line_89[336], line_88[334], line_87[332], line_86[330], line_85[328], line_84[326], line_83[324], line_82[322], line_81[320], line_80[318], line_79[316], line_78[314], line_77[312], line_76[310], line_75[308], line_74[306], line_73[304], line_72[302], line_71[300], line_70[298], line_69[296], line_68[294], line_67[292], line_66[290], line_65[288], line_64[286], line_63[284], line_62[282], line_61[280], line_60[278], line_59[276], line_58[274], line_57[272], line_56[270], line_55[268], line_54[266], line_53[264], line_52[262], line_51[260], line_50[258], line_49[256], line_48[254], line_47[252], line_46[250], line_45[248], line_44[246], line_43[244], line_42[242], line_41[240], line_40[238], line_39[236], line_38[234], line_37[232], line_36[230], line_35[228], line_34[226], line_33[224], line_32[222], line_31[220], line_30[218], line_29[216], line_28[214], line_27[212], line_26[210], line_25[208], line_24[206], line_23[204], line_22[202], line_21[200], line_20[198], line_19[196], line_18[194], line_17[192], line_16[190], line_15[188], line_14[186], line_13[184], line_12[182], line_11[180], line_10[178], line_9[176], line_8[174], line_7[172], line_6[170], line_5[168], line_4[166], line_3[164], line_2[162], line_1[160] };
assign col_415 = {line_128[415], line_127[413], line_126[411], line_125[409], line_124[407], line_123[405], line_122[403], line_121[401], line_120[399], line_119[397], line_118[395], line_117[393], line_116[391], line_115[389], line_114[387], line_113[385], line_112[383], line_111[381], line_110[379], line_109[377], line_108[375], line_107[373], line_106[371], line_105[369], line_104[367], line_103[365], line_102[363], line_101[361], line_100[359], line_99[357], line_98[355], line_97[353], line_96[351], line_95[349], line_94[347], line_93[345], line_92[343], line_91[341], line_90[339], line_89[337], line_88[335], line_87[333], line_86[331], line_85[329], line_84[327], line_83[325], line_82[323], line_81[321], line_80[319], line_79[317], line_78[315], line_77[313], line_76[311], line_75[309], line_74[307], line_73[305], line_72[303], line_71[301], line_70[299], line_69[297], line_68[295], line_67[293], line_66[291], line_65[289], line_64[287], line_63[285], line_62[283], line_61[281], line_60[279], line_59[277], line_58[275], line_57[273], line_56[271], line_55[269], line_54[267], line_53[265], line_52[263], line_51[261], line_50[259], line_49[257], line_48[255], line_47[253], line_46[251], line_45[249], line_44[247], line_43[245], line_42[243], line_41[241], line_40[239], line_39[237], line_38[235], line_37[233], line_36[231], line_35[229], line_34[227], line_33[225], line_32[223], line_31[221], line_30[219], line_29[217], line_28[215], line_27[213], line_26[211], line_25[209], line_24[207], line_23[205], line_22[203], line_21[201], line_20[199], line_19[197], line_18[195], line_17[193], line_16[191], line_15[189], line_14[187], line_13[185], line_12[183], line_11[181], line_10[179], line_9[177], line_8[175], line_7[173], line_6[171], line_5[169], line_4[167], line_3[165], line_2[163], line_1[161] };
assign col_416 = {line_128[416], line_127[414], line_126[412], line_125[410], line_124[408], line_123[406], line_122[404], line_121[402], line_120[400], line_119[398], line_118[396], line_117[394], line_116[392], line_115[390], line_114[388], line_113[386], line_112[384], line_111[382], line_110[380], line_109[378], line_108[376], line_107[374], line_106[372], line_105[370], line_104[368], line_103[366], line_102[364], line_101[362], line_100[360], line_99[358], line_98[356], line_97[354], line_96[352], line_95[350], line_94[348], line_93[346], line_92[344], line_91[342], line_90[340], line_89[338], line_88[336], line_87[334], line_86[332], line_85[330], line_84[328], line_83[326], line_82[324], line_81[322], line_80[320], line_79[318], line_78[316], line_77[314], line_76[312], line_75[310], line_74[308], line_73[306], line_72[304], line_71[302], line_70[300], line_69[298], line_68[296], line_67[294], line_66[292], line_65[290], line_64[288], line_63[286], line_62[284], line_61[282], line_60[280], line_59[278], line_58[276], line_57[274], line_56[272], line_55[270], line_54[268], line_53[266], line_52[264], line_51[262], line_50[260], line_49[258], line_48[256], line_47[254], line_46[252], line_45[250], line_44[248], line_43[246], line_42[244], line_41[242], line_40[240], line_39[238], line_38[236], line_37[234], line_36[232], line_35[230], line_34[228], line_33[226], line_32[224], line_31[222], line_30[220], line_29[218], line_28[216], line_27[214], line_26[212], line_25[210], line_24[208], line_23[206], line_22[204], line_21[202], line_20[200], line_19[198], line_18[196], line_17[194], line_16[192], line_15[190], line_14[188], line_13[186], line_12[184], line_11[182], line_10[180], line_9[178], line_8[176], line_7[174], line_6[172], line_5[170], line_4[168], line_3[166], line_2[164], line_1[162] };
assign col_417 = {line_128[417], line_127[415], line_126[413], line_125[411], line_124[409], line_123[407], line_122[405], line_121[403], line_120[401], line_119[399], line_118[397], line_117[395], line_116[393], line_115[391], line_114[389], line_113[387], line_112[385], line_111[383], line_110[381], line_109[379], line_108[377], line_107[375], line_106[373], line_105[371], line_104[369], line_103[367], line_102[365], line_101[363], line_100[361], line_99[359], line_98[357], line_97[355], line_96[353], line_95[351], line_94[349], line_93[347], line_92[345], line_91[343], line_90[341], line_89[339], line_88[337], line_87[335], line_86[333], line_85[331], line_84[329], line_83[327], line_82[325], line_81[323], line_80[321], line_79[319], line_78[317], line_77[315], line_76[313], line_75[311], line_74[309], line_73[307], line_72[305], line_71[303], line_70[301], line_69[299], line_68[297], line_67[295], line_66[293], line_65[291], line_64[289], line_63[287], line_62[285], line_61[283], line_60[281], line_59[279], line_58[277], line_57[275], line_56[273], line_55[271], line_54[269], line_53[267], line_52[265], line_51[263], line_50[261], line_49[259], line_48[257], line_47[255], line_46[253], line_45[251], line_44[249], line_43[247], line_42[245], line_41[243], line_40[241], line_39[239], line_38[237], line_37[235], line_36[233], line_35[231], line_34[229], line_33[227], line_32[225], line_31[223], line_30[221], line_29[219], line_28[217], line_27[215], line_26[213], line_25[211], line_24[209], line_23[207], line_22[205], line_21[203], line_20[201], line_19[199], line_18[197], line_17[195], line_16[193], line_15[191], line_14[189], line_13[187], line_12[185], line_11[183], line_10[181], line_9[179], line_8[177], line_7[175], line_6[173], line_5[171], line_4[169], line_3[167], line_2[165], line_1[163] };
assign col_418 = {line_128[418], line_127[416], line_126[414], line_125[412], line_124[410], line_123[408], line_122[406], line_121[404], line_120[402], line_119[400], line_118[398], line_117[396], line_116[394], line_115[392], line_114[390], line_113[388], line_112[386], line_111[384], line_110[382], line_109[380], line_108[378], line_107[376], line_106[374], line_105[372], line_104[370], line_103[368], line_102[366], line_101[364], line_100[362], line_99[360], line_98[358], line_97[356], line_96[354], line_95[352], line_94[350], line_93[348], line_92[346], line_91[344], line_90[342], line_89[340], line_88[338], line_87[336], line_86[334], line_85[332], line_84[330], line_83[328], line_82[326], line_81[324], line_80[322], line_79[320], line_78[318], line_77[316], line_76[314], line_75[312], line_74[310], line_73[308], line_72[306], line_71[304], line_70[302], line_69[300], line_68[298], line_67[296], line_66[294], line_65[292], line_64[290], line_63[288], line_62[286], line_61[284], line_60[282], line_59[280], line_58[278], line_57[276], line_56[274], line_55[272], line_54[270], line_53[268], line_52[266], line_51[264], line_50[262], line_49[260], line_48[258], line_47[256], line_46[254], line_45[252], line_44[250], line_43[248], line_42[246], line_41[244], line_40[242], line_39[240], line_38[238], line_37[236], line_36[234], line_35[232], line_34[230], line_33[228], line_32[226], line_31[224], line_30[222], line_29[220], line_28[218], line_27[216], line_26[214], line_25[212], line_24[210], line_23[208], line_22[206], line_21[204], line_20[202], line_19[200], line_18[198], line_17[196], line_16[194], line_15[192], line_14[190], line_13[188], line_12[186], line_11[184], line_10[182], line_9[180], line_8[178], line_7[176], line_6[174], line_5[172], line_4[170], line_3[168], line_2[166], line_1[164] };
assign col_419 = {line_128[419], line_127[417], line_126[415], line_125[413], line_124[411], line_123[409], line_122[407], line_121[405], line_120[403], line_119[401], line_118[399], line_117[397], line_116[395], line_115[393], line_114[391], line_113[389], line_112[387], line_111[385], line_110[383], line_109[381], line_108[379], line_107[377], line_106[375], line_105[373], line_104[371], line_103[369], line_102[367], line_101[365], line_100[363], line_99[361], line_98[359], line_97[357], line_96[355], line_95[353], line_94[351], line_93[349], line_92[347], line_91[345], line_90[343], line_89[341], line_88[339], line_87[337], line_86[335], line_85[333], line_84[331], line_83[329], line_82[327], line_81[325], line_80[323], line_79[321], line_78[319], line_77[317], line_76[315], line_75[313], line_74[311], line_73[309], line_72[307], line_71[305], line_70[303], line_69[301], line_68[299], line_67[297], line_66[295], line_65[293], line_64[291], line_63[289], line_62[287], line_61[285], line_60[283], line_59[281], line_58[279], line_57[277], line_56[275], line_55[273], line_54[271], line_53[269], line_52[267], line_51[265], line_50[263], line_49[261], line_48[259], line_47[257], line_46[255], line_45[253], line_44[251], line_43[249], line_42[247], line_41[245], line_40[243], line_39[241], line_38[239], line_37[237], line_36[235], line_35[233], line_34[231], line_33[229], line_32[227], line_31[225], line_30[223], line_29[221], line_28[219], line_27[217], line_26[215], line_25[213], line_24[211], line_23[209], line_22[207], line_21[205], line_20[203], line_19[201], line_18[199], line_17[197], line_16[195], line_15[193], line_14[191], line_13[189], line_12[187], line_11[185], line_10[183], line_9[181], line_8[179], line_7[177], line_6[175], line_5[173], line_4[171], line_3[169], line_2[167], line_1[165] };
assign col_420 = {line_128[420], line_127[418], line_126[416], line_125[414], line_124[412], line_123[410], line_122[408], line_121[406], line_120[404], line_119[402], line_118[400], line_117[398], line_116[396], line_115[394], line_114[392], line_113[390], line_112[388], line_111[386], line_110[384], line_109[382], line_108[380], line_107[378], line_106[376], line_105[374], line_104[372], line_103[370], line_102[368], line_101[366], line_100[364], line_99[362], line_98[360], line_97[358], line_96[356], line_95[354], line_94[352], line_93[350], line_92[348], line_91[346], line_90[344], line_89[342], line_88[340], line_87[338], line_86[336], line_85[334], line_84[332], line_83[330], line_82[328], line_81[326], line_80[324], line_79[322], line_78[320], line_77[318], line_76[316], line_75[314], line_74[312], line_73[310], line_72[308], line_71[306], line_70[304], line_69[302], line_68[300], line_67[298], line_66[296], line_65[294], line_64[292], line_63[290], line_62[288], line_61[286], line_60[284], line_59[282], line_58[280], line_57[278], line_56[276], line_55[274], line_54[272], line_53[270], line_52[268], line_51[266], line_50[264], line_49[262], line_48[260], line_47[258], line_46[256], line_45[254], line_44[252], line_43[250], line_42[248], line_41[246], line_40[244], line_39[242], line_38[240], line_37[238], line_36[236], line_35[234], line_34[232], line_33[230], line_32[228], line_31[226], line_30[224], line_29[222], line_28[220], line_27[218], line_26[216], line_25[214], line_24[212], line_23[210], line_22[208], line_21[206], line_20[204], line_19[202], line_18[200], line_17[198], line_16[196], line_15[194], line_14[192], line_13[190], line_12[188], line_11[186], line_10[184], line_9[182], line_8[180], line_7[178], line_6[176], line_5[174], line_4[172], line_3[170], line_2[168], line_1[166] };
assign col_421 = {line_128[421], line_127[419], line_126[417], line_125[415], line_124[413], line_123[411], line_122[409], line_121[407], line_120[405], line_119[403], line_118[401], line_117[399], line_116[397], line_115[395], line_114[393], line_113[391], line_112[389], line_111[387], line_110[385], line_109[383], line_108[381], line_107[379], line_106[377], line_105[375], line_104[373], line_103[371], line_102[369], line_101[367], line_100[365], line_99[363], line_98[361], line_97[359], line_96[357], line_95[355], line_94[353], line_93[351], line_92[349], line_91[347], line_90[345], line_89[343], line_88[341], line_87[339], line_86[337], line_85[335], line_84[333], line_83[331], line_82[329], line_81[327], line_80[325], line_79[323], line_78[321], line_77[319], line_76[317], line_75[315], line_74[313], line_73[311], line_72[309], line_71[307], line_70[305], line_69[303], line_68[301], line_67[299], line_66[297], line_65[295], line_64[293], line_63[291], line_62[289], line_61[287], line_60[285], line_59[283], line_58[281], line_57[279], line_56[277], line_55[275], line_54[273], line_53[271], line_52[269], line_51[267], line_50[265], line_49[263], line_48[261], line_47[259], line_46[257], line_45[255], line_44[253], line_43[251], line_42[249], line_41[247], line_40[245], line_39[243], line_38[241], line_37[239], line_36[237], line_35[235], line_34[233], line_33[231], line_32[229], line_31[227], line_30[225], line_29[223], line_28[221], line_27[219], line_26[217], line_25[215], line_24[213], line_23[211], line_22[209], line_21[207], line_20[205], line_19[203], line_18[201], line_17[199], line_16[197], line_15[195], line_14[193], line_13[191], line_12[189], line_11[187], line_10[185], line_9[183], line_8[181], line_7[179], line_6[177], line_5[175], line_4[173], line_3[171], line_2[169], line_1[167] };
assign col_422 = {line_128[422], line_127[420], line_126[418], line_125[416], line_124[414], line_123[412], line_122[410], line_121[408], line_120[406], line_119[404], line_118[402], line_117[400], line_116[398], line_115[396], line_114[394], line_113[392], line_112[390], line_111[388], line_110[386], line_109[384], line_108[382], line_107[380], line_106[378], line_105[376], line_104[374], line_103[372], line_102[370], line_101[368], line_100[366], line_99[364], line_98[362], line_97[360], line_96[358], line_95[356], line_94[354], line_93[352], line_92[350], line_91[348], line_90[346], line_89[344], line_88[342], line_87[340], line_86[338], line_85[336], line_84[334], line_83[332], line_82[330], line_81[328], line_80[326], line_79[324], line_78[322], line_77[320], line_76[318], line_75[316], line_74[314], line_73[312], line_72[310], line_71[308], line_70[306], line_69[304], line_68[302], line_67[300], line_66[298], line_65[296], line_64[294], line_63[292], line_62[290], line_61[288], line_60[286], line_59[284], line_58[282], line_57[280], line_56[278], line_55[276], line_54[274], line_53[272], line_52[270], line_51[268], line_50[266], line_49[264], line_48[262], line_47[260], line_46[258], line_45[256], line_44[254], line_43[252], line_42[250], line_41[248], line_40[246], line_39[244], line_38[242], line_37[240], line_36[238], line_35[236], line_34[234], line_33[232], line_32[230], line_31[228], line_30[226], line_29[224], line_28[222], line_27[220], line_26[218], line_25[216], line_24[214], line_23[212], line_22[210], line_21[208], line_20[206], line_19[204], line_18[202], line_17[200], line_16[198], line_15[196], line_14[194], line_13[192], line_12[190], line_11[188], line_10[186], line_9[184], line_8[182], line_7[180], line_6[178], line_5[176], line_4[174], line_3[172], line_2[170], line_1[168] };
assign col_423 = {line_128[423], line_127[421], line_126[419], line_125[417], line_124[415], line_123[413], line_122[411], line_121[409], line_120[407], line_119[405], line_118[403], line_117[401], line_116[399], line_115[397], line_114[395], line_113[393], line_112[391], line_111[389], line_110[387], line_109[385], line_108[383], line_107[381], line_106[379], line_105[377], line_104[375], line_103[373], line_102[371], line_101[369], line_100[367], line_99[365], line_98[363], line_97[361], line_96[359], line_95[357], line_94[355], line_93[353], line_92[351], line_91[349], line_90[347], line_89[345], line_88[343], line_87[341], line_86[339], line_85[337], line_84[335], line_83[333], line_82[331], line_81[329], line_80[327], line_79[325], line_78[323], line_77[321], line_76[319], line_75[317], line_74[315], line_73[313], line_72[311], line_71[309], line_70[307], line_69[305], line_68[303], line_67[301], line_66[299], line_65[297], line_64[295], line_63[293], line_62[291], line_61[289], line_60[287], line_59[285], line_58[283], line_57[281], line_56[279], line_55[277], line_54[275], line_53[273], line_52[271], line_51[269], line_50[267], line_49[265], line_48[263], line_47[261], line_46[259], line_45[257], line_44[255], line_43[253], line_42[251], line_41[249], line_40[247], line_39[245], line_38[243], line_37[241], line_36[239], line_35[237], line_34[235], line_33[233], line_32[231], line_31[229], line_30[227], line_29[225], line_28[223], line_27[221], line_26[219], line_25[217], line_24[215], line_23[213], line_22[211], line_21[209], line_20[207], line_19[205], line_18[203], line_17[201], line_16[199], line_15[197], line_14[195], line_13[193], line_12[191], line_11[189], line_10[187], line_9[185], line_8[183], line_7[181], line_6[179], line_5[177], line_4[175], line_3[173], line_2[171], line_1[169] };
assign col_424 = {line_128[424], line_127[422], line_126[420], line_125[418], line_124[416], line_123[414], line_122[412], line_121[410], line_120[408], line_119[406], line_118[404], line_117[402], line_116[400], line_115[398], line_114[396], line_113[394], line_112[392], line_111[390], line_110[388], line_109[386], line_108[384], line_107[382], line_106[380], line_105[378], line_104[376], line_103[374], line_102[372], line_101[370], line_100[368], line_99[366], line_98[364], line_97[362], line_96[360], line_95[358], line_94[356], line_93[354], line_92[352], line_91[350], line_90[348], line_89[346], line_88[344], line_87[342], line_86[340], line_85[338], line_84[336], line_83[334], line_82[332], line_81[330], line_80[328], line_79[326], line_78[324], line_77[322], line_76[320], line_75[318], line_74[316], line_73[314], line_72[312], line_71[310], line_70[308], line_69[306], line_68[304], line_67[302], line_66[300], line_65[298], line_64[296], line_63[294], line_62[292], line_61[290], line_60[288], line_59[286], line_58[284], line_57[282], line_56[280], line_55[278], line_54[276], line_53[274], line_52[272], line_51[270], line_50[268], line_49[266], line_48[264], line_47[262], line_46[260], line_45[258], line_44[256], line_43[254], line_42[252], line_41[250], line_40[248], line_39[246], line_38[244], line_37[242], line_36[240], line_35[238], line_34[236], line_33[234], line_32[232], line_31[230], line_30[228], line_29[226], line_28[224], line_27[222], line_26[220], line_25[218], line_24[216], line_23[214], line_22[212], line_21[210], line_20[208], line_19[206], line_18[204], line_17[202], line_16[200], line_15[198], line_14[196], line_13[194], line_12[192], line_11[190], line_10[188], line_9[186], line_8[184], line_7[182], line_6[180], line_5[178], line_4[176], line_3[174], line_2[172], line_1[170] };
assign col_425 = {line_128[425], line_127[423], line_126[421], line_125[419], line_124[417], line_123[415], line_122[413], line_121[411], line_120[409], line_119[407], line_118[405], line_117[403], line_116[401], line_115[399], line_114[397], line_113[395], line_112[393], line_111[391], line_110[389], line_109[387], line_108[385], line_107[383], line_106[381], line_105[379], line_104[377], line_103[375], line_102[373], line_101[371], line_100[369], line_99[367], line_98[365], line_97[363], line_96[361], line_95[359], line_94[357], line_93[355], line_92[353], line_91[351], line_90[349], line_89[347], line_88[345], line_87[343], line_86[341], line_85[339], line_84[337], line_83[335], line_82[333], line_81[331], line_80[329], line_79[327], line_78[325], line_77[323], line_76[321], line_75[319], line_74[317], line_73[315], line_72[313], line_71[311], line_70[309], line_69[307], line_68[305], line_67[303], line_66[301], line_65[299], line_64[297], line_63[295], line_62[293], line_61[291], line_60[289], line_59[287], line_58[285], line_57[283], line_56[281], line_55[279], line_54[277], line_53[275], line_52[273], line_51[271], line_50[269], line_49[267], line_48[265], line_47[263], line_46[261], line_45[259], line_44[257], line_43[255], line_42[253], line_41[251], line_40[249], line_39[247], line_38[245], line_37[243], line_36[241], line_35[239], line_34[237], line_33[235], line_32[233], line_31[231], line_30[229], line_29[227], line_28[225], line_27[223], line_26[221], line_25[219], line_24[217], line_23[215], line_22[213], line_21[211], line_20[209], line_19[207], line_18[205], line_17[203], line_16[201], line_15[199], line_14[197], line_13[195], line_12[193], line_11[191], line_10[189], line_9[187], line_8[185], line_7[183], line_6[181], line_5[179], line_4[177], line_3[175], line_2[173], line_1[171] };
assign col_426 = {line_128[426], line_127[424], line_126[422], line_125[420], line_124[418], line_123[416], line_122[414], line_121[412], line_120[410], line_119[408], line_118[406], line_117[404], line_116[402], line_115[400], line_114[398], line_113[396], line_112[394], line_111[392], line_110[390], line_109[388], line_108[386], line_107[384], line_106[382], line_105[380], line_104[378], line_103[376], line_102[374], line_101[372], line_100[370], line_99[368], line_98[366], line_97[364], line_96[362], line_95[360], line_94[358], line_93[356], line_92[354], line_91[352], line_90[350], line_89[348], line_88[346], line_87[344], line_86[342], line_85[340], line_84[338], line_83[336], line_82[334], line_81[332], line_80[330], line_79[328], line_78[326], line_77[324], line_76[322], line_75[320], line_74[318], line_73[316], line_72[314], line_71[312], line_70[310], line_69[308], line_68[306], line_67[304], line_66[302], line_65[300], line_64[298], line_63[296], line_62[294], line_61[292], line_60[290], line_59[288], line_58[286], line_57[284], line_56[282], line_55[280], line_54[278], line_53[276], line_52[274], line_51[272], line_50[270], line_49[268], line_48[266], line_47[264], line_46[262], line_45[260], line_44[258], line_43[256], line_42[254], line_41[252], line_40[250], line_39[248], line_38[246], line_37[244], line_36[242], line_35[240], line_34[238], line_33[236], line_32[234], line_31[232], line_30[230], line_29[228], line_28[226], line_27[224], line_26[222], line_25[220], line_24[218], line_23[216], line_22[214], line_21[212], line_20[210], line_19[208], line_18[206], line_17[204], line_16[202], line_15[200], line_14[198], line_13[196], line_12[194], line_11[192], line_10[190], line_9[188], line_8[186], line_7[184], line_6[182], line_5[180], line_4[178], line_3[176], line_2[174], line_1[172] };
assign col_427 = {line_128[427], line_127[425], line_126[423], line_125[421], line_124[419], line_123[417], line_122[415], line_121[413], line_120[411], line_119[409], line_118[407], line_117[405], line_116[403], line_115[401], line_114[399], line_113[397], line_112[395], line_111[393], line_110[391], line_109[389], line_108[387], line_107[385], line_106[383], line_105[381], line_104[379], line_103[377], line_102[375], line_101[373], line_100[371], line_99[369], line_98[367], line_97[365], line_96[363], line_95[361], line_94[359], line_93[357], line_92[355], line_91[353], line_90[351], line_89[349], line_88[347], line_87[345], line_86[343], line_85[341], line_84[339], line_83[337], line_82[335], line_81[333], line_80[331], line_79[329], line_78[327], line_77[325], line_76[323], line_75[321], line_74[319], line_73[317], line_72[315], line_71[313], line_70[311], line_69[309], line_68[307], line_67[305], line_66[303], line_65[301], line_64[299], line_63[297], line_62[295], line_61[293], line_60[291], line_59[289], line_58[287], line_57[285], line_56[283], line_55[281], line_54[279], line_53[277], line_52[275], line_51[273], line_50[271], line_49[269], line_48[267], line_47[265], line_46[263], line_45[261], line_44[259], line_43[257], line_42[255], line_41[253], line_40[251], line_39[249], line_38[247], line_37[245], line_36[243], line_35[241], line_34[239], line_33[237], line_32[235], line_31[233], line_30[231], line_29[229], line_28[227], line_27[225], line_26[223], line_25[221], line_24[219], line_23[217], line_22[215], line_21[213], line_20[211], line_19[209], line_18[207], line_17[205], line_16[203], line_15[201], line_14[199], line_13[197], line_12[195], line_11[193], line_10[191], line_9[189], line_8[187], line_7[185], line_6[183], line_5[181], line_4[179], line_3[177], line_2[175], line_1[173] };
assign col_428 = {line_128[428], line_127[426], line_126[424], line_125[422], line_124[420], line_123[418], line_122[416], line_121[414], line_120[412], line_119[410], line_118[408], line_117[406], line_116[404], line_115[402], line_114[400], line_113[398], line_112[396], line_111[394], line_110[392], line_109[390], line_108[388], line_107[386], line_106[384], line_105[382], line_104[380], line_103[378], line_102[376], line_101[374], line_100[372], line_99[370], line_98[368], line_97[366], line_96[364], line_95[362], line_94[360], line_93[358], line_92[356], line_91[354], line_90[352], line_89[350], line_88[348], line_87[346], line_86[344], line_85[342], line_84[340], line_83[338], line_82[336], line_81[334], line_80[332], line_79[330], line_78[328], line_77[326], line_76[324], line_75[322], line_74[320], line_73[318], line_72[316], line_71[314], line_70[312], line_69[310], line_68[308], line_67[306], line_66[304], line_65[302], line_64[300], line_63[298], line_62[296], line_61[294], line_60[292], line_59[290], line_58[288], line_57[286], line_56[284], line_55[282], line_54[280], line_53[278], line_52[276], line_51[274], line_50[272], line_49[270], line_48[268], line_47[266], line_46[264], line_45[262], line_44[260], line_43[258], line_42[256], line_41[254], line_40[252], line_39[250], line_38[248], line_37[246], line_36[244], line_35[242], line_34[240], line_33[238], line_32[236], line_31[234], line_30[232], line_29[230], line_28[228], line_27[226], line_26[224], line_25[222], line_24[220], line_23[218], line_22[216], line_21[214], line_20[212], line_19[210], line_18[208], line_17[206], line_16[204], line_15[202], line_14[200], line_13[198], line_12[196], line_11[194], line_10[192], line_9[190], line_8[188], line_7[186], line_6[184], line_5[182], line_4[180], line_3[178], line_2[176], line_1[174] };
assign col_429 = {line_128[429], line_127[427], line_126[425], line_125[423], line_124[421], line_123[419], line_122[417], line_121[415], line_120[413], line_119[411], line_118[409], line_117[407], line_116[405], line_115[403], line_114[401], line_113[399], line_112[397], line_111[395], line_110[393], line_109[391], line_108[389], line_107[387], line_106[385], line_105[383], line_104[381], line_103[379], line_102[377], line_101[375], line_100[373], line_99[371], line_98[369], line_97[367], line_96[365], line_95[363], line_94[361], line_93[359], line_92[357], line_91[355], line_90[353], line_89[351], line_88[349], line_87[347], line_86[345], line_85[343], line_84[341], line_83[339], line_82[337], line_81[335], line_80[333], line_79[331], line_78[329], line_77[327], line_76[325], line_75[323], line_74[321], line_73[319], line_72[317], line_71[315], line_70[313], line_69[311], line_68[309], line_67[307], line_66[305], line_65[303], line_64[301], line_63[299], line_62[297], line_61[295], line_60[293], line_59[291], line_58[289], line_57[287], line_56[285], line_55[283], line_54[281], line_53[279], line_52[277], line_51[275], line_50[273], line_49[271], line_48[269], line_47[267], line_46[265], line_45[263], line_44[261], line_43[259], line_42[257], line_41[255], line_40[253], line_39[251], line_38[249], line_37[247], line_36[245], line_35[243], line_34[241], line_33[239], line_32[237], line_31[235], line_30[233], line_29[231], line_28[229], line_27[227], line_26[225], line_25[223], line_24[221], line_23[219], line_22[217], line_21[215], line_20[213], line_19[211], line_18[209], line_17[207], line_16[205], line_15[203], line_14[201], line_13[199], line_12[197], line_11[195], line_10[193], line_9[191], line_8[189], line_7[187], line_6[185], line_5[183], line_4[181], line_3[179], line_2[177], line_1[175] };
assign col_430 = {line_128[430], line_127[428], line_126[426], line_125[424], line_124[422], line_123[420], line_122[418], line_121[416], line_120[414], line_119[412], line_118[410], line_117[408], line_116[406], line_115[404], line_114[402], line_113[400], line_112[398], line_111[396], line_110[394], line_109[392], line_108[390], line_107[388], line_106[386], line_105[384], line_104[382], line_103[380], line_102[378], line_101[376], line_100[374], line_99[372], line_98[370], line_97[368], line_96[366], line_95[364], line_94[362], line_93[360], line_92[358], line_91[356], line_90[354], line_89[352], line_88[350], line_87[348], line_86[346], line_85[344], line_84[342], line_83[340], line_82[338], line_81[336], line_80[334], line_79[332], line_78[330], line_77[328], line_76[326], line_75[324], line_74[322], line_73[320], line_72[318], line_71[316], line_70[314], line_69[312], line_68[310], line_67[308], line_66[306], line_65[304], line_64[302], line_63[300], line_62[298], line_61[296], line_60[294], line_59[292], line_58[290], line_57[288], line_56[286], line_55[284], line_54[282], line_53[280], line_52[278], line_51[276], line_50[274], line_49[272], line_48[270], line_47[268], line_46[266], line_45[264], line_44[262], line_43[260], line_42[258], line_41[256], line_40[254], line_39[252], line_38[250], line_37[248], line_36[246], line_35[244], line_34[242], line_33[240], line_32[238], line_31[236], line_30[234], line_29[232], line_28[230], line_27[228], line_26[226], line_25[224], line_24[222], line_23[220], line_22[218], line_21[216], line_20[214], line_19[212], line_18[210], line_17[208], line_16[206], line_15[204], line_14[202], line_13[200], line_12[198], line_11[196], line_10[194], line_9[192], line_8[190], line_7[188], line_6[186], line_5[184], line_4[182], line_3[180], line_2[178], line_1[176] };
assign col_431 = {line_128[431], line_127[429], line_126[427], line_125[425], line_124[423], line_123[421], line_122[419], line_121[417], line_120[415], line_119[413], line_118[411], line_117[409], line_116[407], line_115[405], line_114[403], line_113[401], line_112[399], line_111[397], line_110[395], line_109[393], line_108[391], line_107[389], line_106[387], line_105[385], line_104[383], line_103[381], line_102[379], line_101[377], line_100[375], line_99[373], line_98[371], line_97[369], line_96[367], line_95[365], line_94[363], line_93[361], line_92[359], line_91[357], line_90[355], line_89[353], line_88[351], line_87[349], line_86[347], line_85[345], line_84[343], line_83[341], line_82[339], line_81[337], line_80[335], line_79[333], line_78[331], line_77[329], line_76[327], line_75[325], line_74[323], line_73[321], line_72[319], line_71[317], line_70[315], line_69[313], line_68[311], line_67[309], line_66[307], line_65[305], line_64[303], line_63[301], line_62[299], line_61[297], line_60[295], line_59[293], line_58[291], line_57[289], line_56[287], line_55[285], line_54[283], line_53[281], line_52[279], line_51[277], line_50[275], line_49[273], line_48[271], line_47[269], line_46[267], line_45[265], line_44[263], line_43[261], line_42[259], line_41[257], line_40[255], line_39[253], line_38[251], line_37[249], line_36[247], line_35[245], line_34[243], line_33[241], line_32[239], line_31[237], line_30[235], line_29[233], line_28[231], line_27[229], line_26[227], line_25[225], line_24[223], line_23[221], line_22[219], line_21[217], line_20[215], line_19[213], line_18[211], line_17[209], line_16[207], line_15[205], line_14[203], line_13[201], line_12[199], line_11[197], line_10[195], line_9[193], line_8[191], line_7[189], line_6[187], line_5[185], line_4[183], line_3[181], line_2[179], line_1[177] };
assign col_432 = {line_128[432], line_127[430], line_126[428], line_125[426], line_124[424], line_123[422], line_122[420], line_121[418], line_120[416], line_119[414], line_118[412], line_117[410], line_116[408], line_115[406], line_114[404], line_113[402], line_112[400], line_111[398], line_110[396], line_109[394], line_108[392], line_107[390], line_106[388], line_105[386], line_104[384], line_103[382], line_102[380], line_101[378], line_100[376], line_99[374], line_98[372], line_97[370], line_96[368], line_95[366], line_94[364], line_93[362], line_92[360], line_91[358], line_90[356], line_89[354], line_88[352], line_87[350], line_86[348], line_85[346], line_84[344], line_83[342], line_82[340], line_81[338], line_80[336], line_79[334], line_78[332], line_77[330], line_76[328], line_75[326], line_74[324], line_73[322], line_72[320], line_71[318], line_70[316], line_69[314], line_68[312], line_67[310], line_66[308], line_65[306], line_64[304], line_63[302], line_62[300], line_61[298], line_60[296], line_59[294], line_58[292], line_57[290], line_56[288], line_55[286], line_54[284], line_53[282], line_52[280], line_51[278], line_50[276], line_49[274], line_48[272], line_47[270], line_46[268], line_45[266], line_44[264], line_43[262], line_42[260], line_41[258], line_40[256], line_39[254], line_38[252], line_37[250], line_36[248], line_35[246], line_34[244], line_33[242], line_32[240], line_31[238], line_30[236], line_29[234], line_28[232], line_27[230], line_26[228], line_25[226], line_24[224], line_23[222], line_22[220], line_21[218], line_20[216], line_19[214], line_18[212], line_17[210], line_16[208], line_15[206], line_14[204], line_13[202], line_12[200], line_11[198], line_10[196], line_9[194], line_8[192], line_7[190], line_6[188], line_5[186], line_4[184], line_3[182], line_2[180], line_1[178] };
assign col_433 = {line_128[433], line_127[431], line_126[429], line_125[427], line_124[425], line_123[423], line_122[421], line_121[419], line_120[417], line_119[415], line_118[413], line_117[411], line_116[409], line_115[407], line_114[405], line_113[403], line_112[401], line_111[399], line_110[397], line_109[395], line_108[393], line_107[391], line_106[389], line_105[387], line_104[385], line_103[383], line_102[381], line_101[379], line_100[377], line_99[375], line_98[373], line_97[371], line_96[369], line_95[367], line_94[365], line_93[363], line_92[361], line_91[359], line_90[357], line_89[355], line_88[353], line_87[351], line_86[349], line_85[347], line_84[345], line_83[343], line_82[341], line_81[339], line_80[337], line_79[335], line_78[333], line_77[331], line_76[329], line_75[327], line_74[325], line_73[323], line_72[321], line_71[319], line_70[317], line_69[315], line_68[313], line_67[311], line_66[309], line_65[307], line_64[305], line_63[303], line_62[301], line_61[299], line_60[297], line_59[295], line_58[293], line_57[291], line_56[289], line_55[287], line_54[285], line_53[283], line_52[281], line_51[279], line_50[277], line_49[275], line_48[273], line_47[271], line_46[269], line_45[267], line_44[265], line_43[263], line_42[261], line_41[259], line_40[257], line_39[255], line_38[253], line_37[251], line_36[249], line_35[247], line_34[245], line_33[243], line_32[241], line_31[239], line_30[237], line_29[235], line_28[233], line_27[231], line_26[229], line_25[227], line_24[225], line_23[223], line_22[221], line_21[219], line_20[217], line_19[215], line_18[213], line_17[211], line_16[209], line_15[207], line_14[205], line_13[203], line_12[201], line_11[199], line_10[197], line_9[195], line_8[193], line_7[191], line_6[189], line_5[187], line_4[185], line_3[183], line_2[181], line_1[179] };
assign col_434 = {line_128[434], line_127[432], line_126[430], line_125[428], line_124[426], line_123[424], line_122[422], line_121[420], line_120[418], line_119[416], line_118[414], line_117[412], line_116[410], line_115[408], line_114[406], line_113[404], line_112[402], line_111[400], line_110[398], line_109[396], line_108[394], line_107[392], line_106[390], line_105[388], line_104[386], line_103[384], line_102[382], line_101[380], line_100[378], line_99[376], line_98[374], line_97[372], line_96[370], line_95[368], line_94[366], line_93[364], line_92[362], line_91[360], line_90[358], line_89[356], line_88[354], line_87[352], line_86[350], line_85[348], line_84[346], line_83[344], line_82[342], line_81[340], line_80[338], line_79[336], line_78[334], line_77[332], line_76[330], line_75[328], line_74[326], line_73[324], line_72[322], line_71[320], line_70[318], line_69[316], line_68[314], line_67[312], line_66[310], line_65[308], line_64[306], line_63[304], line_62[302], line_61[300], line_60[298], line_59[296], line_58[294], line_57[292], line_56[290], line_55[288], line_54[286], line_53[284], line_52[282], line_51[280], line_50[278], line_49[276], line_48[274], line_47[272], line_46[270], line_45[268], line_44[266], line_43[264], line_42[262], line_41[260], line_40[258], line_39[256], line_38[254], line_37[252], line_36[250], line_35[248], line_34[246], line_33[244], line_32[242], line_31[240], line_30[238], line_29[236], line_28[234], line_27[232], line_26[230], line_25[228], line_24[226], line_23[224], line_22[222], line_21[220], line_20[218], line_19[216], line_18[214], line_17[212], line_16[210], line_15[208], line_14[206], line_13[204], line_12[202], line_11[200], line_10[198], line_9[196], line_8[194], line_7[192], line_6[190], line_5[188], line_4[186], line_3[184], line_2[182], line_1[180] };
assign col_435 = {line_128[435], line_127[433], line_126[431], line_125[429], line_124[427], line_123[425], line_122[423], line_121[421], line_120[419], line_119[417], line_118[415], line_117[413], line_116[411], line_115[409], line_114[407], line_113[405], line_112[403], line_111[401], line_110[399], line_109[397], line_108[395], line_107[393], line_106[391], line_105[389], line_104[387], line_103[385], line_102[383], line_101[381], line_100[379], line_99[377], line_98[375], line_97[373], line_96[371], line_95[369], line_94[367], line_93[365], line_92[363], line_91[361], line_90[359], line_89[357], line_88[355], line_87[353], line_86[351], line_85[349], line_84[347], line_83[345], line_82[343], line_81[341], line_80[339], line_79[337], line_78[335], line_77[333], line_76[331], line_75[329], line_74[327], line_73[325], line_72[323], line_71[321], line_70[319], line_69[317], line_68[315], line_67[313], line_66[311], line_65[309], line_64[307], line_63[305], line_62[303], line_61[301], line_60[299], line_59[297], line_58[295], line_57[293], line_56[291], line_55[289], line_54[287], line_53[285], line_52[283], line_51[281], line_50[279], line_49[277], line_48[275], line_47[273], line_46[271], line_45[269], line_44[267], line_43[265], line_42[263], line_41[261], line_40[259], line_39[257], line_38[255], line_37[253], line_36[251], line_35[249], line_34[247], line_33[245], line_32[243], line_31[241], line_30[239], line_29[237], line_28[235], line_27[233], line_26[231], line_25[229], line_24[227], line_23[225], line_22[223], line_21[221], line_20[219], line_19[217], line_18[215], line_17[213], line_16[211], line_15[209], line_14[207], line_13[205], line_12[203], line_11[201], line_10[199], line_9[197], line_8[195], line_7[193], line_6[191], line_5[189], line_4[187], line_3[185], line_2[183], line_1[181] };
assign col_436 = {line_128[436], line_127[434], line_126[432], line_125[430], line_124[428], line_123[426], line_122[424], line_121[422], line_120[420], line_119[418], line_118[416], line_117[414], line_116[412], line_115[410], line_114[408], line_113[406], line_112[404], line_111[402], line_110[400], line_109[398], line_108[396], line_107[394], line_106[392], line_105[390], line_104[388], line_103[386], line_102[384], line_101[382], line_100[380], line_99[378], line_98[376], line_97[374], line_96[372], line_95[370], line_94[368], line_93[366], line_92[364], line_91[362], line_90[360], line_89[358], line_88[356], line_87[354], line_86[352], line_85[350], line_84[348], line_83[346], line_82[344], line_81[342], line_80[340], line_79[338], line_78[336], line_77[334], line_76[332], line_75[330], line_74[328], line_73[326], line_72[324], line_71[322], line_70[320], line_69[318], line_68[316], line_67[314], line_66[312], line_65[310], line_64[308], line_63[306], line_62[304], line_61[302], line_60[300], line_59[298], line_58[296], line_57[294], line_56[292], line_55[290], line_54[288], line_53[286], line_52[284], line_51[282], line_50[280], line_49[278], line_48[276], line_47[274], line_46[272], line_45[270], line_44[268], line_43[266], line_42[264], line_41[262], line_40[260], line_39[258], line_38[256], line_37[254], line_36[252], line_35[250], line_34[248], line_33[246], line_32[244], line_31[242], line_30[240], line_29[238], line_28[236], line_27[234], line_26[232], line_25[230], line_24[228], line_23[226], line_22[224], line_21[222], line_20[220], line_19[218], line_18[216], line_17[214], line_16[212], line_15[210], line_14[208], line_13[206], line_12[204], line_11[202], line_10[200], line_9[198], line_8[196], line_7[194], line_6[192], line_5[190], line_4[188], line_3[186], line_2[184], line_1[182] };
assign col_437 = {line_128[437], line_127[435], line_126[433], line_125[431], line_124[429], line_123[427], line_122[425], line_121[423], line_120[421], line_119[419], line_118[417], line_117[415], line_116[413], line_115[411], line_114[409], line_113[407], line_112[405], line_111[403], line_110[401], line_109[399], line_108[397], line_107[395], line_106[393], line_105[391], line_104[389], line_103[387], line_102[385], line_101[383], line_100[381], line_99[379], line_98[377], line_97[375], line_96[373], line_95[371], line_94[369], line_93[367], line_92[365], line_91[363], line_90[361], line_89[359], line_88[357], line_87[355], line_86[353], line_85[351], line_84[349], line_83[347], line_82[345], line_81[343], line_80[341], line_79[339], line_78[337], line_77[335], line_76[333], line_75[331], line_74[329], line_73[327], line_72[325], line_71[323], line_70[321], line_69[319], line_68[317], line_67[315], line_66[313], line_65[311], line_64[309], line_63[307], line_62[305], line_61[303], line_60[301], line_59[299], line_58[297], line_57[295], line_56[293], line_55[291], line_54[289], line_53[287], line_52[285], line_51[283], line_50[281], line_49[279], line_48[277], line_47[275], line_46[273], line_45[271], line_44[269], line_43[267], line_42[265], line_41[263], line_40[261], line_39[259], line_38[257], line_37[255], line_36[253], line_35[251], line_34[249], line_33[247], line_32[245], line_31[243], line_30[241], line_29[239], line_28[237], line_27[235], line_26[233], line_25[231], line_24[229], line_23[227], line_22[225], line_21[223], line_20[221], line_19[219], line_18[217], line_17[215], line_16[213], line_15[211], line_14[209], line_13[207], line_12[205], line_11[203], line_10[201], line_9[199], line_8[197], line_7[195], line_6[193], line_5[191], line_4[189], line_3[187], line_2[185], line_1[183] };
assign col_438 = {line_128[438], line_127[436], line_126[434], line_125[432], line_124[430], line_123[428], line_122[426], line_121[424], line_120[422], line_119[420], line_118[418], line_117[416], line_116[414], line_115[412], line_114[410], line_113[408], line_112[406], line_111[404], line_110[402], line_109[400], line_108[398], line_107[396], line_106[394], line_105[392], line_104[390], line_103[388], line_102[386], line_101[384], line_100[382], line_99[380], line_98[378], line_97[376], line_96[374], line_95[372], line_94[370], line_93[368], line_92[366], line_91[364], line_90[362], line_89[360], line_88[358], line_87[356], line_86[354], line_85[352], line_84[350], line_83[348], line_82[346], line_81[344], line_80[342], line_79[340], line_78[338], line_77[336], line_76[334], line_75[332], line_74[330], line_73[328], line_72[326], line_71[324], line_70[322], line_69[320], line_68[318], line_67[316], line_66[314], line_65[312], line_64[310], line_63[308], line_62[306], line_61[304], line_60[302], line_59[300], line_58[298], line_57[296], line_56[294], line_55[292], line_54[290], line_53[288], line_52[286], line_51[284], line_50[282], line_49[280], line_48[278], line_47[276], line_46[274], line_45[272], line_44[270], line_43[268], line_42[266], line_41[264], line_40[262], line_39[260], line_38[258], line_37[256], line_36[254], line_35[252], line_34[250], line_33[248], line_32[246], line_31[244], line_30[242], line_29[240], line_28[238], line_27[236], line_26[234], line_25[232], line_24[230], line_23[228], line_22[226], line_21[224], line_20[222], line_19[220], line_18[218], line_17[216], line_16[214], line_15[212], line_14[210], line_13[208], line_12[206], line_11[204], line_10[202], line_9[200], line_8[198], line_7[196], line_6[194], line_5[192], line_4[190], line_3[188], line_2[186], line_1[184] };
assign col_439 = {line_128[439], line_127[437], line_126[435], line_125[433], line_124[431], line_123[429], line_122[427], line_121[425], line_120[423], line_119[421], line_118[419], line_117[417], line_116[415], line_115[413], line_114[411], line_113[409], line_112[407], line_111[405], line_110[403], line_109[401], line_108[399], line_107[397], line_106[395], line_105[393], line_104[391], line_103[389], line_102[387], line_101[385], line_100[383], line_99[381], line_98[379], line_97[377], line_96[375], line_95[373], line_94[371], line_93[369], line_92[367], line_91[365], line_90[363], line_89[361], line_88[359], line_87[357], line_86[355], line_85[353], line_84[351], line_83[349], line_82[347], line_81[345], line_80[343], line_79[341], line_78[339], line_77[337], line_76[335], line_75[333], line_74[331], line_73[329], line_72[327], line_71[325], line_70[323], line_69[321], line_68[319], line_67[317], line_66[315], line_65[313], line_64[311], line_63[309], line_62[307], line_61[305], line_60[303], line_59[301], line_58[299], line_57[297], line_56[295], line_55[293], line_54[291], line_53[289], line_52[287], line_51[285], line_50[283], line_49[281], line_48[279], line_47[277], line_46[275], line_45[273], line_44[271], line_43[269], line_42[267], line_41[265], line_40[263], line_39[261], line_38[259], line_37[257], line_36[255], line_35[253], line_34[251], line_33[249], line_32[247], line_31[245], line_30[243], line_29[241], line_28[239], line_27[237], line_26[235], line_25[233], line_24[231], line_23[229], line_22[227], line_21[225], line_20[223], line_19[221], line_18[219], line_17[217], line_16[215], line_15[213], line_14[211], line_13[209], line_12[207], line_11[205], line_10[203], line_9[201], line_8[199], line_7[197], line_6[195], line_5[193], line_4[191], line_3[189], line_2[187], line_1[185] };
assign col_440 = {line_128[440], line_127[438], line_126[436], line_125[434], line_124[432], line_123[430], line_122[428], line_121[426], line_120[424], line_119[422], line_118[420], line_117[418], line_116[416], line_115[414], line_114[412], line_113[410], line_112[408], line_111[406], line_110[404], line_109[402], line_108[400], line_107[398], line_106[396], line_105[394], line_104[392], line_103[390], line_102[388], line_101[386], line_100[384], line_99[382], line_98[380], line_97[378], line_96[376], line_95[374], line_94[372], line_93[370], line_92[368], line_91[366], line_90[364], line_89[362], line_88[360], line_87[358], line_86[356], line_85[354], line_84[352], line_83[350], line_82[348], line_81[346], line_80[344], line_79[342], line_78[340], line_77[338], line_76[336], line_75[334], line_74[332], line_73[330], line_72[328], line_71[326], line_70[324], line_69[322], line_68[320], line_67[318], line_66[316], line_65[314], line_64[312], line_63[310], line_62[308], line_61[306], line_60[304], line_59[302], line_58[300], line_57[298], line_56[296], line_55[294], line_54[292], line_53[290], line_52[288], line_51[286], line_50[284], line_49[282], line_48[280], line_47[278], line_46[276], line_45[274], line_44[272], line_43[270], line_42[268], line_41[266], line_40[264], line_39[262], line_38[260], line_37[258], line_36[256], line_35[254], line_34[252], line_33[250], line_32[248], line_31[246], line_30[244], line_29[242], line_28[240], line_27[238], line_26[236], line_25[234], line_24[232], line_23[230], line_22[228], line_21[226], line_20[224], line_19[222], line_18[220], line_17[218], line_16[216], line_15[214], line_14[212], line_13[210], line_12[208], line_11[206], line_10[204], line_9[202], line_8[200], line_7[198], line_6[196], line_5[194], line_4[192], line_3[190], line_2[188], line_1[186] };
assign col_441 = {line_128[441], line_127[439], line_126[437], line_125[435], line_124[433], line_123[431], line_122[429], line_121[427], line_120[425], line_119[423], line_118[421], line_117[419], line_116[417], line_115[415], line_114[413], line_113[411], line_112[409], line_111[407], line_110[405], line_109[403], line_108[401], line_107[399], line_106[397], line_105[395], line_104[393], line_103[391], line_102[389], line_101[387], line_100[385], line_99[383], line_98[381], line_97[379], line_96[377], line_95[375], line_94[373], line_93[371], line_92[369], line_91[367], line_90[365], line_89[363], line_88[361], line_87[359], line_86[357], line_85[355], line_84[353], line_83[351], line_82[349], line_81[347], line_80[345], line_79[343], line_78[341], line_77[339], line_76[337], line_75[335], line_74[333], line_73[331], line_72[329], line_71[327], line_70[325], line_69[323], line_68[321], line_67[319], line_66[317], line_65[315], line_64[313], line_63[311], line_62[309], line_61[307], line_60[305], line_59[303], line_58[301], line_57[299], line_56[297], line_55[295], line_54[293], line_53[291], line_52[289], line_51[287], line_50[285], line_49[283], line_48[281], line_47[279], line_46[277], line_45[275], line_44[273], line_43[271], line_42[269], line_41[267], line_40[265], line_39[263], line_38[261], line_37[259], line_36[257], line_35[255], line_34[253], line_33[251], line_32[249], line_31[247], line_30[245], line_29[243], line_28[241], line_27[239], line_26[237], line_25[235], line_24[233], line_23[231], line_22[229], line_21[227], line_20[225], line_19[223], line_18[221], line_17[219], line_16[217], line_15[215], line_14[213], line_13[211], line_12[209], line_11[207], line_10[205], line_9[203], line_8[201], line_7[199], line_6[197], line_5[195], line_4[193], line_3[191], line_2[189], line_1[187] };
assign col_442 = {line_128[442], line_127[440], line_126[438], line_125[436], line_124[434], line_123[432], line_122[430], line_121[428], line_120[426], line_119[424], line_118[422], line_117[420], line_116[418], line_115[416], line_114[414], line_113[412], line_112[410], line_111[408], line_110[406], line_109[404], line_108[402], line_107[400], line_106[398], line_105[396], line_104[394], line_103[392], line_102[390], line_101[388], line_100[386], line_99[384], line_98[382], line_97[380], line_96[378], line_95[376], line_94[374], line_93[372], line_92[370], line_91[368], line_90[366], line_89[364], line_88[362], line_87[360], line_86[358], line_85[356], line_84[354], line_83[352], line_82[350], line_81[348], line_80[346], line_79[344], line_78[342], line_77[340], line_76[338], line_75[336], line_74[334], line_73[332], line_72[330], line_71[328], line_70[326], line_69[324], line_68[322], line_67[320], line_66[318], line_65[316], line_64[314], line_63[312], line_62[310], line_61[308], line_60[306], line_59[304], line_58[302], line_57[300], line_56[298], line_55[296], line_54[294], line_53[292], line_52[290], line_51[288], line_50[286], line_49[284], line_48[282], line_47[280], line_46[278], line_45[276], line_44[274], line_43[272], line_42[270], line_41[268], line_40[266], line_39[264], line_38[262], line_37[260], line_36[258], line_35[256], line_34[254], line_33[252], line_32[250], line_31[248], line_30[246], line_29[244], line_28[242], line_27[240], line_26[238], line_25[236], line_24[234], line_23[232], line_22[230], line_21[228], line_20[226], line_19[224], line_18[222], line_17[220], line_16[218], line_15[216], line_14[214], line_13[212], line_12[210], line_11[208], line_10[206], line_9[204], line_8[202], line_7[200], line_6[198], line_5[196], line_4[194], line_3[192], line_2[190], line_1[188] };
assign col_443 = {line_128[443], line_127[441], line_126[439], line_125[437], line_124[435], line_123[433], line_122[431], line_121[429], line_120[427], line_119[425], line_118[423], line_117[421], line_116[419], line_115[417], line_114[415], line_113[413], line_112[411], line_111[409], line_110[407], line_109[405], line_108[403], line_107[401], line_106[399], line_105[397], line_104[395], line_103[393], line_102[391], line_101[389], line_100[387], line_99[385], line_98[383], line_97[381], line_96[379], line_95[377], line_94[375], line_93[373], line_92[371], line_91[369], line_90[367], line_89[365], line_88[363], line_87[361], line_86[359], line_85[357], line_84[355], line_83[353], line_82[351], line_81[349], line_80[347], line_79[345], line_78[343], line_77[341], line_76[339], line_75[337], line_74[335], line_73[333], line_72[331], line_71[329], line_70[327], line_69[325], line_68[323], line_67[321], line_66[319], line_65[317], line_64[315], line_63[313], line_62[311], line_61[309], line_60[307], line_59[305], line_58[303], line_57[301], line_56[299], line_55[297], line_54[295], line_53[293], line_52[291], line_51[289], line_50[287], line_49[285], line_48[283], line_47[281], line_46[279], line_45[277], line_44[275], line_43[273], line_42[271], line_41[269], line_40[267], line_39[265], line_38[263], line_37[261], line_36[259], line_35[257], line_34[255], line_33[253], line_32[251], line_31[249], line_30[247], line_29[245], line_28[243], line_27[241], line_26[239], line_25[237], line_24[235], line_23[233], line_22[231], line_21[229], line_20[227], line_19[225], line_18[223], line_17[221], line_16[219], line_15[217], line_14[215], line_13[213], line_12[211], line_11[209], line_10[207], line_9[205], line_8[203], line_7[201], line_6[199], line_5[197], line_4[195], line_3[193], line_2[191], line_1[189] };
assign col_444 = {line_128[444], line_127[442], line_126[440], line_125[438], line_124[436], line_123[434], line_122[432], line_121[430], line_120[428], line_119[426], line_118[424], line_117[422], line_116[420], line_115[418], line_114[416], line_113[414], line_112[412], line_111[410], line_110[408], line_109[406], line_108[404], line_107[402], line_106[400], line_105[398], line_104[396], line_103[394], line_102[392], line_101[390], line_100[388], line_99[386], line_98[384], line_97[382], line_96[380], line_95[378], line_94[376], line_93[374], line_92[372], line_91[370], line_90[368], line_89[366], line_88[364], line_87[362], line_86[360], line_85[358], line_84[356], line_83[354], line_82[352], line_81[350], line_80[348], line_79[346], line_78[344], line_77[342], line_76[340], line_75[338], line_74[336], line_73[334], line_72[332], line_71[330], line_70[328], line_69[326], line_68[324], line_67[322], line_66[320], line_65[318], line_64[316], line_63[314], line_62[312], line_61[310], line_60[308], line_59[306], line_58[304], line_57[302], line_56[300], line_55[298], line_54[296], line_53[294], line_52[292], line_51[290], line_50[288], line_49[286], line_48[284], line_47[282], line_46[280], line_45[278], line_44[276], line_43[274], line_42[272], line_41[270], line_40[268], line_39[266], line_38[264], line_37[262], line_36[260], line_35[258], line_34[256], line_33[254], line_32[252], line_31[250], line_30[248], line_29[246], line_28[244], line_27[242], line_26[240], line_25[238], line_24[236], line_23[234], line_22[232], line_21[230], line_20[228], line_19[226], line_18[224], line_17[222], line_16[220], line_15[218], line_14[216], line_13[214], line_12[212], line_11[210], line_10[208], line_9[206], line_8[204], line_7[202], line_6[200], line_5[198], line_4[196], line_3[194], line_2[192], line_1[190] };
assign col_445 = {line_128[445], line_127[443], line_126[441], line_125[439], line_124[437], line_123[435], line_122[433], line_121[431], line_120[429], line_119[427], line_118[425], line_117[423], line_116[421], line_115[419], line_114[417], line_113[415], line_112[413], line_111[411], line_110[409], line_109[407], line_108[405], line_107[403], line_106[401], line_105[399], line_104[397], line_103[395], line_102[393], line_101[391], line_100[389], line_99[387], line_98[385], line_97[383], line_96[381], line_95[379], line_94[377], line_93[375], line_92[373], line_91[371], line_90[369], line_89[367], line_88[365], line_87[363], line_86[361], line_85[359], line_84[357], line_83[355], line_82[353], line_81[351], line_80[349], line_79[347], line_78[345], line_77[343], line_76[341], line_75[339], line_74[337], line_73[335], line_72[333], line_71[331], line_70[329], line_69[327], line_68[325], line_67[323], line_66[321], line_65[319], line_64[317], line_63[315], line_62[313], line_61[311], line_60[309], line_59[307], line_58[305], line_57[303], line_56[301], line_55[299], line_54[297], line_53[295], line_52[293], line_51[291], line_50[289], line_49[287], line_48[285], line_47[283], line_46[281], line_45[279], line_44[277], line_43[275], line_42[273], line_41[271], line_40[269], line_39[267], line_38[265], line_37[263], line_36[261], line_35[259], line_34[257], line_33[255], line_32[253], line_31[251], line_30[249], line_29[247], line_28[245], line_27[243], line_26[241], line_25[239], line_24[237], line_23[235], line_22[233], line_21[231], line_20[229], line_19[227], line_18[225], line_17[223], line_16[221], line_15[219], line_14[217], line_13[215], line_12[213], line_11[211], line_10[209], line_9[207], line_8[205], line_7[203], line_6[201], line_5[199], line_4[197], line_3[195], line_2[193], line_1[191] };
assign col_446 = {line_128[446], line_127[444], line_126[442], line_125[440], line_124[438], line_123[436], line_122[434], line_121[432], line_120[430], line_119[428], line_118[426], line_117[424], line_116[422], line_115[420], line_114[418], line_113[416], line_112[414], line_111[412], line_110[410], line_109[408], line_108[406], line_107[404], line_106[402], line_105[400], line_104[398], line_103[396], line_102[394], line_101[392], line_100[390], line_99[388], line_98[386], line_97[384], line_96[382], line_95[380], line_94[378], line_93[376], line_92[374], line_91[372], line_90[370], line_89[368], line_88[366], line_87[364], line_86[362], line_85[360], line_84[358], line_83[356], line_82[354], line_81[352], line_80[350], line_79[348], line_78[346], line_77[344], line_76[342], line_75[340], line_74[338], line_73[336], line_72[334], line_71[332], line_70[330], line_69[328], line_68[326], line_67[324], line_66[322], line_65[320], line_64[318], line_63[316], line_62[314], line_61[312], line_60[310], line_59[308], line_58[306], line_57[304], line_56[302], line_55[300], line_54[298], line_53[296], line_52[294], line_51[292], line_50[290], line_49[288], line_48[286], line_47[284], line_46[282], line_45[280], line_44[278], line_43[276], line_42[274], line_41[272], line_40[270], line_39[268], line_38[266], line_37[264], line_36[262], line_35[260], line_34[258], line_33[256], line_32[254], line_31[252], line_30[250], line_29[248], line_28[246], line_27[244], line_26[242], line_25[240], line_24[238], line_23[236], line_22[234], line_21[232], line_20[230], line_19[228], line_18[226], line_17[224], line_16[222], line_15[220], line_14[218], line_13[216], line_12[214], line_11[212], line_10[210], line_9[208], line_8[206], line_7[204], line_6[202], line_5[200], line_4[198], line_3[196], line_2[194], line_1[192] };
assign col_447 = {line_128[447], line_127[445], line_126[443], line_125[441], line_124[439], line_123[437], line_122[435], line_121[433], line_120[431], line_119[429], line_118[427], line_117[425], line_116[423], line_115[421], line_114[419], line_113[417], line_112[415], line_111[413], line_110[411], line_109[409], line_108[407], line_107[405], line_106[403], line_105[401], line_104[399], line_103[397], line_102[395], line_101[393], line_100[391], line_99[389], line_98[387], line_97[385], line_96[383], line_95[381], line_94[379], line_93[377], line_92[375], line_91[373], line_90[371], line_89[369], line_88[367], line_87[365], line_86[363], line_85[361], line_84[359], line_83[357], line_82[355], line_81[353], line_80[351], line_79[349], line_78[347], line_77[345], line_76[343], line_75[341], line_74[339], line_73[337], line_72[335], line_71[333], line_70[331], line_69[329], line_68[327], line_67[325], line_66[323], line_65[321], line_64[319], line_63[317], line_62[315], line_61[313], line_60[311], line_59[309], line_58[307], line_57[305], line_56[303], line_55[301], line_54[299], line_53[297], line_52[295], line_51[293], line_50[291], line_49[289], line_48[287], line_47[285], line_46[283], line_45[281], line_44[279], line_43[277], line_42[275], line_41[273], line_40[271], line_39[269], line_38[267], line_37[265], line_36[263], line_35[261], line_34[259], line_33[257], line_32[255], line_31[253], line_30[251], line_29[249], line_28[247], line_27[245], line_26[243], line_25[241], line_24[239], line_23[237], line_22[235], line_21[233], line_20[231], line_19[229], line_18[227], line_17[225], line_16[223], line_15[221], line_14[219], line_13[217], line_12[215], line_11[213], line_10[211], line_9[209], line_8[207], line_7[205], line_6[203], line_5[201], line_4[199], line_3[197], line_2[195], line_1[193] };
assign col_448 = {line_128[448], line_127[446], line_126[444], line_125[442], line_124[440], line_123[438], line_122[436], line_121[434], line_120[432], line_119[430], line_118[428], line_117[426], line_116[424], line_115[422], line_114[420], line_113[418], line_112[416], line_111[414], line_110[412], line_109[410], line_108[408], line_107[406], line_106[404], line_105[402], line_104[400], line_103[398], line_102[396], line_101[394], line_100[392], line_99[390], line_98[388], line_97[386], line_96[384], line_95[382], line_94[380], line_93[378], line_92[376], line_91[374], line_90[372], line_89[370], line_88[368], line_87[366], line_86[364], line_85[362], line_84[360], line_83[358], line_82[356], line_81[354], line_80[352], line_79[350], line_78[348], line_77[346], line_76[344], line_75[342], line_74[340], line_73[338], line_72[336], line_71[334], line_70[332], line_69[330], line_68[328], line_67[326], line_66[324], line_65[322], line_64[320], line_63[318], line_62[316], line_61[314], line_60[312], line_59[310], line_58[308], line_57[306], line_56[304], line_55[302], line_54[300], line_53[298], line_52[296], line_51[294], line_50[292], line_49[290], line_48[288], line_47[286], line_46[284], line_45[282], line_44[280], line_43[278], line_42[276], line_41[274], line_40[272], line_39[270], line_38[268], line_37[266], line_36[264], line_35[262], line_34[260], line_33[258], line_32[256], line_31[254], line_30[252], line_29[250], line_28[248], line_27[246], line_26[244], line_25[242], line_24[240], line_23[238], line_22[236], line_21[234], line_20[232], line_19[230], line_18[228], line_17[226], line_16[224], line_15[222], line_14[220], line_13[218], line_12[216], line_11[214], line_10[212], line_9[210], line_8[208], line_7[206], line_6[204], line_5[202], line_4[200], line_3[198], line_2[196], line_1[194] };
assign col_449 = {line_128[449], line_127[447], line_126[445], line_125[443], line_124[441], line_123[439], line_122[437], line_121[435], line_120[433], line_119[431], line_118[429], line_117[427], line_116[425], line_115[423], line_114[421], line_113[419], line_112[417], line_111[415], line_110[413], line_109[411], line_108[409], line_107[407], line_106[405], line_105[403], line_104[401], line_103[399], line_102[397], line_101[395], line_100[393], line_99[391], line_98[389], line_97[387], line_96[385], line_95[383], line_94[381], line_93[379], line_92[377], line_91[375], line_90[373], line_89[371], line_88[369], line_87[367], line_86[365], line_85[363], line_84[361], line_83[359], line_82[357], line_81[355], line_80[353], line_79[351], line_78[349], line_77[347], line_76[345], line_75[343], line_74[341], line_73[339], line_72[337], line_71[335], line_70[333], line_69[331], line_68[329], line_67[327], line_66[325], line_65[323], line_64[321], line_63[319], line_62[317], line_61[315], line_60[313], line_59[311], line_58[309], line_57[307], line_56[305], line_55[303], line_54[301], line_53[299], line_52[297], line_51[295], line_50[293], line_49[291], line_48[289], line_47[287], line_46[285], line_45[283], line_44[281], line_43[279], line_42[277], line_41[275], line_40[273], line_39[271], line_38[269], line_37[267], line_36[265], line_35[263], line_34[261], line_33[259], line_32[257], line_31[255], line_30[253], line_29[251], line_28[249], line_27[247], line_26[245], line_25[243], line_24[241], line_23[239], line_22[237], line_21[235], line_20[233], line_19[231], line_18[229], line_17[227], line_16[225], line_15[223], line_14[221], line_13[219], line_12[217], line_11[215], line_10[213], line_9[211], line_8[209], line_7[207], line_6[205], line_5[203], line_4[201], line_3[199], line_2[197], line_1[195] };
assign col_450 = {line_128[450], line_127[448], line_126[446], line_125[444], line_124[442], line_123[440], line_122[438], line_121[436], line_120[434], line_119[432], line_118[430], line_117[428], line_116[426], line_115[424], line_114[422], line_113[420], line_112[418], line_111[416], line_110[414], line_109[412], line_108[410], line_107[408], line_106[406], line_105[404], line_104[402], line_103[400], line_102[398], line_101[396], line_100[394], line_99[392], line_98[390], line_97[388], line_96[386], line_95[384], line_94[382], line_93[380], line_92[378], line_91[376], line_90[374], line_89[372], line_88[370], line_87[368], line_86[366], line_85[364], line_84[362], line_83[360], line_82[358], line_81[356], line_80[354], line_79[352], line_78[350], line_77[348], line_76[346], line_75[344], line_74[342], line_73[340], line_72[338], line_71[336], line_70[334], line_69[332], line_68[330], line_67[328], line_66[326], line_65[324], line_64[322], line_63[320], line_62[318], line_61[316], line_60[314], line_59[312], line_58[310], line_57[308], line_56[306], line_55[304], line_54[302], line_53[300], line_52[298], line_51[296], line_50[294], line_49[292], line_48[290], line_47[288], line_46[286], line_45[284], line_44[282], line_43[280], line_42[278], line_41[276], line_40[274], line_39[272], line_38[270], line_37[268], line_36[266], line_35[264], line_34[262], line_33[260], line_32[258], line_31[256], line_30[254], line_29[252], line_28[250], line_27[248], line_26[246], line_25[244], line_24[242], line_23[240], line_22[238], line_21[236], line_20[234], line_19[232], line_18[230], line_17[228], line_16[226], line_15[224], line_14[222], line_13[220], line_12[218], line_11[216], line_10[214], line_9[212], line_8[210], line_7[208], line_6[206], line_5[204], line_4[202], line_3[200], line_2[198], line_1[196] };
assign col_451 = {line_128[451], line_127[449], line_126[447], line_125[445], line_124[443], line_123[441], line_122[439], line_121[437], line_120[435], line_119[433], line_118[431], line_117[429], line_116[427], line_115[425], line_114[423], line_113[421], line_112[419], line_111[417], line_110[415], line_109[413], line_108[411], line_107[409], line_106[407], line_105[405], line_104[403], line_103[401], line_102[399], line_101[397], line_100[395], line_99[393], line_98[391], line_97[389], line_96[387], line_95[385], line_94[383], line_93[381], line_92[379], line_91[377], line_90[375], line_89[373], line_88[371], line_87[369], line_86[367], line_85[365], line_84[363], line_83[361], line_82[359], line_81[357], line_80[355], line_79[353], line_78[351], line_77[349], line_76[347], line_75[345], line_74[343], line_73[341], line_72[339], line_71[337], line_70[335], line_69[333], line_68[331], line_67[329], line_66[327], line_65[325], line_64[323], line_63[321], line_62[319], line_61[317], line_60[315], line_59[313], line_58[311], line_57[309], line_56[307], line_55[305], line_54[303], line_53[301], line_52[299], line_51[297], line_50[295], line_49[293], line_48[291], line_47[289], line_46[287], line_45[285], line_44[283], line_43[281], line_42[279], line_41[277], line_40[275], line_39[273], line_38[271], line_37[269], line_36[267], line_35[265], line_34[263], line_33[261], line_32[259], line_31[257], line_30[255], line_29[253], line_28[251], line_27[249], line_26[247], line_25[245], line_24[243], line_23[241], line_22[239], line_21[237], line_20[235], line_19[233], line_18[231], line_17[229], line_16[227], line_15[225], line_14[223], line_13[221], line_12[219], line_11[217], line_10[215], line_9[213], line_8[211], line_7[209], line_6[207], line_5[205], line_4[203], line_3[201], line_2[199], line_1[197] };
assign col_452 = {line_128[452], line_127[450], line_126[448], line_125[446], line_124[444], line_123[442], line_122[440], line_121[438], line_120[436], line_119[434], line_118[432], line_117[430], line_116[428], line_115[426], line_114[424], line_113[422], line_112[420], line_111[418], line_110[416], line_109[414], line_108[412], line_107[410], line_106[408], line_105[406], line_104[404], line_103[402], line_102[400], line_101[398], line_100[396], line_99[394], line_98[392], line_97[390], line_96[388], line_95[386], line_94[384], line_93[382], line_92[380], line_91[378], line_90[376], line_89[374], line_88[372], line_87[370], line_86[368], line_85[366], line_84[364], line_83[362], line_82[360], line_81[358], line_80[356], line_79[354], line_78[352], line_77[350], line_76[348], line_75[346], line_74[344], line_73[342], line_72[340], line_71[338], line_70[336], line_69[334], line_68[332], line_67[330], line_66[328], line_65[326], line_64[324], line_63[322], line_62[320], line_61[318], line_60[316], line_59[314], line_58[312], line_57[310], line_56[308], line_55[306], line_54[304], line_53[302], line_52[300], line_51[298], line_50[296], line_49[294], line_48[292], line_47[290], line_46[288], line_45[286], line_44[284], line_43[282], line_42[280], line_41[278], line_40[276], line_39[274], line_38[272], line_37[270], line_36[268], line_35[266], line_34[264], line_33[262], line_32[260], line_31[258], line_30[256], line_29[254], line_28[252], line_27[250], line_26[248], line_25[246], line_24[244], line_23[242], line_22[240], line_21[238], line_20[236], line_19[234], line_18[232], line_17[230], line_16[228], line_15[226], line_14[224], line_13[222], line_12[220], line_11[218], line_10[216], line_9[214], line_8[212], line_7[210], line_6[208], line_5[206], line_4[204], line_3[202], line_2[200], line_1[198] };
assign col_453 = {line_128[453], line_127[451], line_126[449], line_125[447], line_124[445], line_123[443], line_122[441], line_121[439], line_120[437], line_119[435], line_118[433], line_117[431], line_116[429], line_115[427], line_114[425], line_113[423], line_112[421], line_111[419], line_110[417], line_109[415], line_108[413], line_107[411], line_106[409], line_105[407], line_104[405], line_103[403], line_102[401], line_101[399], line_100[397], line_99[395], line_98[393], line_97[391], line_96[389], line_95[387], line_94[385], line_93[383], line_92[381], line_91[379], line_90[377], line_89[375], line_88[373], line_87[371], line_86[369], line_85[367], line_84[365], line_83[363], line_82[361], line_81[359], line_80[357], line_79[355], line_78[353], line_77[351], line_76[349], line_75[347], line_74[345], line_73[343], line_72[341], line_71[339], line_70[337], line_69[335], line_68[333], line_67[331], line_66[329], line_65[327], line_64[325], line_63[323], line_62[321], line_61[319], line_60[317], line_59[315], line_58[313], line_57[311], line_56[309], line_55[307], line_54[305], line_53[303], line_52[301], line_51[299], line_50[297], line_49[295], line_48[293], line_47[291], line_46[289], line_45[287], line_44[285], line_43[283], line_42[281], line_41[279], line_40[277], line_39[275], line_38[273], line_37[271], line_36[269], line_35[267], line_34[265], line_33[263], line_32[261], line_31[259], line_30[257], line_29[255], line_28[253], line_27[251], line_26[249], line_25[247], line_24[245], line_23[243], line_22[241], line_21[239], line_20[237], line_19[235], line_18[233], line_17[231], line_16[229], line_15[227], line_14[225], line_13[223], line_12[221], line_11[219], line_10[217], line_9[215], line_8[213], line_7[211], line_6[209], line_5[207], line_4[205], line_3[203], line_2[201], line_1[199] };
assign col_454 = {line_128[454], line_127[452], line_126[450], line_125[448], line_124[446], line_123[444], line_122[442], line_121[440], line_120[438], line_119[436], line_118[434], line_117[432], line_116[430], line_115[428], line_114[426], line_113[424], line_112[422], line_111[420], line_110[418], line_109[416], line_108[414], line_107[412], line_106[410], line_105[408], line_104[406], line_103[404], line_102[402], line_101[400], line_100[398], line_99[396], line_98[394], line_97[392], line_96[390], line_95[388], line_94[386], line_93[384], line_92[382], line_91[380], line_90[378], line_89[376], line_88[374], line_87[372], line_86[370], line_85[368], line_84[366], line_83[364], line_82[362], line_81[360], line_80[358], line_79[356], line_78[354], line_77[352], line_76[350], line_75[348], line_74[346], line_73[344], line_72[342], line_71[340], line_70[338], line_69[336], line_68[334], line_67[332], line_66[330], line_65[328], line_64[326], line_63[324], line_62[322], line_61[320], line_60[318], line_59[316], line_58[314], line_57[312], line_56[310], line_55[308], line_54[306], line_53[304], line_52[302], line_51[300], line_50[298], line_49[296], line_48[294], line_47[292], line_46[290], line_45[288], line_44[286], line_43[284], line_42[282], line_41[280], line_40[278], line_39[276], line_38[274], line_37[272], line_36[270], line_35[268], line_34[266], line_33[264], line_32[262], line_31[260], line_30[258], line_29[256], line_28[254], line_27[252], line_26[250], line_25[248], line_24[246], line_23[244], line_22[242], line_21[240], line_20[238], line_19[236], line_18[234], line_17[232], line_16[230], line_15[228], line_14[226], line_13[224], line_12[222], line_11[220], line_10[218], line_9[216], line_8[214], line_7[212], line_6[210], line_5[208], line_4[206], line_3[204], line_2[202], line_1[200] };
assign col_455 = {line_128[455], line_127[453], line_126[451], line_125[449], line_124[447], line_123[445], line_122[443], line_121[441], line_120[439], line_119[437], line_118[435], line_117[433], line_116[431], line_115[429], line_114[427], line_113[425], line_112[423], line_111[421], line_110[419], line_109[417], line_108[415], line_107[413], line_106[411], line_105[409], line_104[407], line_103[405], line_102[403], line_101[401], line_100[399], line_99[397], line_98[395], line_97[393], line_96[391], line_95[389], line_94[387], line_93[385], line_92[383], line_91[381], line_90[379], line_89[377], line_88[375], line_87[373], line_86[371], line_85[369], line_84[367], line_83[365], line_82[363], line_81[361], line_80[359], line_79[357], line_78[355], line_77[353], line_76[351], line_75[349], line_74[347], line_73[345], line_72[343], line_71[341], line_70[339], line_69[337], line_68[335], line_67[333], line_66[331], line_65[329], line_64[327], line_63[325], line_62[323], line_61[321], line_60[319], line_59[317], line_58[315], line_57[313], line_56[311], line_55[309], line_54[307], line_53[305], line_52[303], line_51[301], line_50[299], line_49[297], line_48[295], line_47[293], line_46[291], line_45[289], line_44[287], line_43[285], line_42[283], line_41[281], line_40[279], line_39[277], line_38[275], line_37[273], line_36[271], line_35[269], line_34[267], line_33[265], line_32[263], line_31[261], line_30[259], line_29[257], line_28[255], line_27[253], line_26[251], line_25[249], line_24[247], line_23[245], line_22[243], line_21[241], line_20[239], line_19[237], line_18[235], line_17[233], line_16[231], line_15[229], line_14[227], line_13[225], line_12[223], line_11[221], line_10[219], line_9[217], line_8[215], line_7[213], line_6[211], line_5[209], line_4[207], line_3[205], line_2[203], line_1[201] };
assign col_456 = {line_128[456], line_127[454], line_126[452], line_125[450], line_124[448], line_123[446], line_122[444], line_121[442], line_120[440], line_119[438], line_118[436], line_117[434], line_116[432], line_115[430], line_114[428], line_113[426], line_112[424], line_111[422], line_110[420], line_109[418], line_108[416], line_107[414], line_106[412], line_105[410], line_104[408], line_103[406], line_102[404], line_101[402], line_100[400], line_99[398], line_98[396], line_97[394], line_96[392], line_95[390], line_94[388], line_93[386], line_92[384], line_91[382], line_90[380], line_89[378], line_88[376], line_87[374], line_86[372], line_85[370], line_84[368], line_83[366], line_82[364], line_81[362], line_80[360], line_79[358], line_78[356], line_77[354], line_76[352], line_75[350], line_74[348], line_73[346], line_72[344], line_71[342], line_70[340], line_69[338], line_68[336], line_67[334], line_66[332], line_65[330], line_64[328], line_63[326], line_62[324], line_61[322], line_60[320], line_59[318], line_58[316], line_57[314], line_56[312], line_55[310], line_54[308], line_53[306], line_52[304], line_51[302], line_50[300], line_49[298], line_48[296], line_47[294], line_46[292], line_45[290], line_44[288], line_43[286], line_42[284], line_41[282], line_40[280], line_39[278], line_38[276], line_37[274], line_36[272], line_35[270], line_34[268], line_33[266], line_32[264], line_31[262], line_30[260], line_29[258], line_28[256], line_27[254], line_26[252], line_25[250], line_24[248], line_23[246], line_22[244], line_21[242], line_20[240], line_19[238], line_18[236], line_17[234], line_16[232], line_15[230], line_14[228], line_13[226], line_12[224], line_11[222], line_10[220], line_9[218], line_8[216], line_7[214], line_6[212], line_5[210], line_4[208], line_3[206], line_2[204], line_1[202] };
assign col_457 = {line_128[457], line_127[455], line_126[453], line_125[451], line_124[449], line_123[447], line_122[445], line_121[443], line_120[441], line_119[439], line_118[437], line_117[435], line_116[433], line_115[431], line_114[429], line_113[427], line_112[425], line_111[423], line_110[421], line_109[419], line_108[417], line_107[415], line_106[413], line_105[411], line_104[409], line_103[407], line_102[405], line_101[403], line_100[401], line_99[399], line_98[397], line_97[395], line_96[393], line_95[391], line_94[389], line_93[387], line_92[385], line_91[383], line_90[381], line_89[379], line_88[377], line_87[375], line_86[373], line_85[371], line_84[369], line_83[367], line_82[365], line_81[363], line_80[361], line_79[359], line_78[357], line_77[355], line_76[353], line_75[351], line_74[349], line_73[347], line_72[345], line_71[343], line_70[341], line_69[339], line_68[337], line_67[335], line_66[333], line_65[331], line_64[329], line_63[327], line_62[325], line_61[323], line_60[321], line_59[319], line_58[317], line_57[315], line_56[313], line_55[311], line_54[309], line_53[307], line_52[305], line_51[303], line_50[301], line_49[299], line_48[297], line_47[295], line_46[293], line_45[291], line_44[289], line_43[287], line_42[285], line_41[283], line_40[281], line_39[279], line_38[277], line_37[275], line_36[273], line_35[271], line_34[269], line_33[267], line_32[265], line_31[263], line_30[261], line_29[259], line_28[257], line_27[255], line_26[253], line_25[251], line_24[249], line_23[247], line_22[245], line_21[243], line_20[241], line_19[239], line_18[237], line_17[235], line_16[233], line_15[231], line_14[229], line_13[227], line_12[225], line_11[223], line_10[221], line_9[219], line_8[217], line_7[215], line_6[213], line_5[211], line_4[209], line_3[207], line_2[205], line_1[203] };
assign col_458 = {line_128[458], line_127[456], line_126[454], line_125[452], line_124[450], line_123[448], line_122[446], line_121[444], line_120[442], line_119[440], line_118[438], line_117[436], line_116[434], line_115[432], line_114[430], line_113[428], line_112[426], line_111[424], line_110[422], line_109[420], line_108[418], line_107[416], line_106[414], line_105[412], line_104[410], line_103[408], line_102[406], line_101[404], line_100[402], line_99[400], line_98[398], line_97[396], line_96[394], line_95[392], line_94[390], line_93[388], line_92[386], line_91[384], line_90[382], line_89[380], line_88[378], line_87[376], line_86[374], line_85[372], line_84[370], line_83[368], line_82[366], line_81[364], line_80[362], line_79[360], line_78[358], line_77[356], line_76[354], line_75[352], line_74[350], line_73[348], line_72[346], line_71[344], line_70[342], line_69[340], line_68[338], line_67[336], line_66[334], line_65[332], line_64[330], line_63[328], line_62[326], line_61[324], line_60[322], line_59[320], line_58[318], line_57[316], line_56[314], line_55[312], line_54[310], line_53[308], line_52[306], line_51[304], line_50[302], line_49[300], line_48[298], line_47[296], line_46[294], line_45[292], line_44[290], line_43[288], line_42[286], line_41[284], line_40[282], line_39[280], line_38[278], line_37[276], line_36[274], line_35[272], line_34[270], line_33[268], line_32[266], line_31[264], line_30[262], line_29[260], line_28[258], line_27[256], line_26[254], line_25[252], line_24[250], line_23[248], line_22[246], line_21[244], line_20[242], line_19[240], line_18[238], line_17[236], line_16[234], line_15[232], line_14[230], line_13[228], line_12[226], line_11[224], line_10[222], line_9[220], line_8[218], line_7[216], line_6[214], line_5[212], line_4[210], line_3[208], line_2[206], line_1[204] };
assign col_459 = {line_128[459], line_127[457], line_126[455], line_125[453], line_124[451], line_123[449], line_122[447], line_121[445], line_120[443], line_119[441], line_118[439], line_117[437], line_116[435], line_115[433], line_114[431], line_113[429], line_112[427], line_111[425], line_110[423], line_109[421], line_108[419], line_107[417], line_106[415], line_105[413], line_104[411], line_103[409], line_102[407], line_101[405], line_100[403], line_99[401], line_98[399], line_97[397], line_96[395], line_95[393], line_94[391], line_93[389], line_92[387], line_91[385], line_90[383], line_89[381], line_88[379], line_87[377], line_86[375], line_85[373], line_84[371], line_83[369], line_82[367], line_81[365], line_80[363], line_79[361], line_78[359], line_77[357], line_76[355], line_75[353], line_74[351], line_73[349], line_72[347], line_71[345], line_70[343], line_69[341], line_68[339], line_67[337], line_66[335], line_65[333], line_64[331], line_63[329], line_62[327], line_61[325], line_60[323], line_59[321], line_58[319], line_57[317], line_56[315], line_55[313], line_54[311], line_53[309], line_52[307], line_51[305], line_50[303], line_49[301], line_48[299], line_47[297], line_46[295], line_45[293], line_44[291], line_43[289], line_42[287], line_41[285], line_40[283], line_39[281], line_38[279], line_37[277], line_36[275], line_35[273], line_34[271], line_33[269], line_32[267], line_31[265], line_30[263], line_29[261], line_28[259], line_27[257], line_26[255], line_25[253], line_24[251], line_23[249], line_22[247], line_21[245], line_20[243], line_19[241], line_18[239], line_17[237], line_16[235], line_15[233], line_14[231], line_13[229], line_12[227], line_11[225], line_10[223], line_9[221], line_8[219], line_7[217], line_6[215], line_5[213], line_4[211], line_3[209], line_2[207], line_1[205] };
assign col_460 = {line_128[460], line_127[458], line_126[456], line_125[454], line_124[452], line_123[450], line_122[448], line_121[446], line_120[444], line_119[442], line_118[440], line_117[438], line_116[436], line_115[434], line_114[432], line_113[430], line_112[428], line_111[426], line_110[424], line_109[422], line_108[420], line_107[418], line_106[416], line_105[414], line_104[412], line_103[410], line_102[408], line_101[406], line_100[404], line_99[402], line_98[400], line_97[398], line_96[396], line_95[394], line_94[392], line_93[390], line_92[388], line_91[386], line_90[384], line_89[382], line_88[380], line_87[378], line_86[376], line_85[374], line_84[372], line_83[370], line_82[368], line_81[366], line_80[364], line_79[362], line_78[360], line_77[358], line_76[356], line_75[354], line_74[352], line_73[350], line_72[348], line_71[346], line_70[344], line_69[342], line_68[340], line_67[338], line_66[336], line_65[334], line_64[332], line_63[330], line_62[328], line_61[326], line_60[324], line_59[322], line_58[320], line_57[318], line_56[316], line_55[314], line_54[312], line_53[310], line_52[308], line_51[306], line_50[304], line_49[302], line_48[300], line_47[298], line_46[296], line_45[294], line_44[292], line_43[290], line_42[288], line_41[286], line_40[284], line_39[282], line_38[280], line_37[278], line_36[276], line_35[274], line_34[272], line_33[270], line_32[268], line_31[266], line_30[264], line_29[262], line_28[260], line_27[258], line_26[256], line_25[254], line_24[252], line_23[250], line_22[248], line_21[246], line_20[244], line_19[242], line_18[240], line_17[238], line_16[236], line_15[234], line_14[232], line_13[230], line_12[228], line_11[226], line_10[224], line_9[222], line_8[220], line_7[218], line_6[216], line_5[214], line_4[212], line_3[210], line_2[208], line_1[206] };
assign col_461 = {line_128[461], line_127[459], line_126[457], line_125[455], line_124[453], line_123[451], line_122[449], line_121[447], line_120[445], line_119[443], line_118[441], line_117[439], line_116[437], line_115[435], line_114[433], line_113[431], line_112[429], line_111[427], line_110[425], line_109[423], line_108[421], line_107[419], line_106[417], line_105[415], line_104[413], line_103[411], line_102[409], line_101[407], line_100[405], line_99[403], line_98[401], line_97[399], line_96[397], line_95[395], line_94[393], line_93[391], line_92[389], line_91[387], line_90[385], line_89[383], line_88[381], line_87[379], line_86[377], line_85[375], line_84[373], line_83[371], line_82[369], line_81[367], line_80[365], line_79[363], line_78[361], line_77[359], line_76[357], line_75[355], line_74[353], line_73[351], line_72[349], line_71[347], line_70[345], line_69[343], line_68[341], line_67[339], line_66[337], line_65[335], line_64[333], line_63[331], line_62[329], line_61[327], line_60[325], line_59[323], line_58[321], line_57[319], line_56[317], line_55[315], line_54[313], line_53[311], line_52[309], line_51[307], line_50[305], line_49[303], line_48[301], line_47[299], line_46[297], line_45[295], line_44[293], line_43[291], line_42[289], line_41[287], line_40[285], line_39[283], line_38[281], line_37[279], line_36[277], line_35[275], line_34[273], line_33[271], line_32[269], line_31[267], line_30[265], line_29[263], line_28[261], line_27[259], line_26[257], line_25[255], line_24[253], line_23[251], line_22[249], line_21[247], line_20[245], line_19[243], line_18[241], line_17[239], line_16[237], line_15[235], line_14[233], line_13[231], line_12[229], line_11[227], line_10[225], line_9[223], line_8[221], line_7[219], line_6[217], line_5[215], line_4[213], line_3[211], line_2[209], line_1[207] };
assign col_462 = {line_128[462], line_127[460], line_126[458], line_125[456], line_124[454], line_123[452], line_122[450], line_121[448], line_120[446], line_119[444], line_118[442], line_117[440], line_116[438], line_115[436], line_114[434], line_113[432], line_112[430], line_111[428], line_110[426], line_109[424], line_108[422], line_107[420], line_106[418], line_105[416], line_104[414], line_103[412], line_102[410], line_101[408], line_100[406], line_99[404], line_98[402], line_97[400], line_96[398], line_95[396], line_94[394], line_93[392], line_92[390], line_91[388], line_90[386], line_89[384], line_88[382], line_87[380], line_86[378], line_85[376], line_84[374], line_83[372], line_82[370], line_81[368], line_80[366], line_79[364], line_78[362], line_77[360], line_76[358], line_75[356], line_74[354], line_73[352], line_72[350], line_71[348], line_70[346], line_69[344], line_68[342], line_67[340], line_66[338], line_65[336], line_64[334], line_63[332], line_62[330], line_61[328], line_60[326], line_59[324], line_58[322], line_57[320], line_56[318], line_55[316], line_54[314], line_53[312], line_52[310], line_51[308], line_50[306], line_49[304], line_48[302], line_47[300], line_46[298], line_45[296], line_44[294], line_43[292], line_42[290], line_41[288], line_40[286], line_39[284], line_38[282], line_37[280], line_36[278], line_35[276], line_34[274], line_33[272], line_32[270], line_31[268], line_30[266], line_29[264], line_28[262], line_27[260], line_26[258], line_25[256], line_24[254], line_23[252], line_22[250], line_21[248], line_20[246], line_19[244], line_18[242], line_17[240], line_16[238], line_15[236], line_14[234], line_13[232], line_12[230], line_11[228], line_10[226], line_9[224], line_8[222], line_7[220], line_6[218], line_5[216], line_4[214], line_3[212], line_2[210], line_1[208] };
assign col_463 = {line_128[463], line_127[461], line_126[459], line_125[457], line_124[455], line_123[453], line_122[451], line_121[449], line_120[447], line_119[445], line_118[443], line_117[441], line_116[439], line_115[437], line_114[435], line_113[433], line_112[431], line_111[429], line_110[427], line_109[425], line_108[423], line_107[421], line_106[419], line_105[417], line_104[415], line_103[413], line_102[411], line_101[409], line_100[407], line_99[405], line_98[403], line_97[401], line_96[399], line_95[397], line_94[395], line_93[393], line_92[391], line_91[389], line_90[387], line_89[385], line_88[383], line_87[381], line_86[379], line_85[377], line_84[375], line_83[373], line_82[371], line_81[369], line_80[367], line_79[365], line_78[363], line_77[361], line_76[359], line_75[357], line_74[355], line_73[353], line_72[351], line_71[349], line_70[347], line_69[345], line_68[343], line_67[341], line_66[339], line_65[337], line_64[335], line_63[333], line_62[331], line_61[329], line_60[327], line_59[325], line_58[323], line_57[321], line_56[319], line_55[317], line_54[315], line_53[313], line_52[311], line_51[309], line_50[307], line_49[305], line_48[303], line_47[301], line_46[299], line_45[297], line_44[295], line_43[293], line_42[291], line_41[289], line_40[287], line_39[285], line_38[283], line_37[281], line_36[279], line_35[277], line_34[275], line_33[273], line_32[271], line_31[269], line_30[267], line_29[265], line_28[263], line_27[261], line_26[259], line_25[257], line_24[255], line_23[253], line_22[251], line_21[249], line_20[247], line_19[245], line_18[243], line_17[241], line_16[239], line_15[237], line_14[235], line_13[233], line_12[231], line_11[229], line_10[227], line_9[225], line_8[223], line_7[221], line_6[219], line_5[217], line_4[215], line_3[213], line_2[211], line_1[209] };
assign col_464 = {line_128[464], line_127[462], line_126[460], line_125[458], line_124[456], line_123[454], line_122[452], line_121[450], line_120[448], line_119[446], line_118[444], line_117[442], line_116[440], line_115[438], line_114[436], line_113[434], line_112[432], line_111[430], line_110[428], line_109[426], line_108[424], line_107[422], line_106[420], line_105[418], line_104[416], line_103[414], line_102[412], line_101[410], line_100[408], line_99[406], line_98[404], line_97[402], line_96[400], line_95[398], line_94[396], line_93[394], line_92[392], line_91[390], line_90[388], line_89[386], line_88[384], line_87[382], line_86[380], line_85[378], line_84[376], line_83[374], line_82[372], line_81[370], line_80[368], line_79[366], line_78[364], line_77[362], line_76[360], line_75[358], line_74[356], line_73[354], line_72[352], line_71[350], line_70[348], line_69[346], line_68[344], line_67[342], line_66[340], line_65[338], line_64[336], line_63[334], line_62[332], line_61[330], line_60[328], line_59[326], line_58[324], line_57[322], line_56[320], line_55[318], line_54[316], line_53[314], line_52[312], line_51[310], line_50[308], line_49[306], line_48[304], line_47[302], line_46[300], line_45[298], line_44[296], line_43[294], line_42[292], line_41[290], line_40[288], line_39[286], line_38[284], line_37[282], line_36[280], line_35[278], line_34[276], line_33[274], line_32[272], line_31[270], line_30[268], line_29[266], line_28[264], line_27[262], line_26[260], line_25[258], line_24[256], line_23[254], line_22[252], line_21[250], line_20[248], line_19[246], line_18[244], line_17[242], line_16[240], line_15[238], line_14[236], line_13[234], line_12[232], line_11[230], line_10[228], line_9[226], line_8[224], line_7[222], line_6[220], line_5[218], line_4[216], line_3[214], line_2[212], line_1[210] };
assign col_465 = {line_128[465], line_127[463], line_126[461], line_125[459], line_124[457], line_123[455], line_122[453], line_121[451], line_120[449], line_119[447], line_118[445], line_117[443], line_116[441], line_115[439], line_114[437], line_113[435], line_112[433], line_111[431], line_110[429], line_109[427], line_108[425], line_107[423], line_106[421], line_105[419], line_104[417], line_103[415], line_102[413], line_101[411], line_100[409], line_99[407], line_98[405], line_97[403], line_96[401], line_95[399], line_94[397], line_93[395], line_92[393], line_91[391], line_90[389], line_89[387], line_88[385], line_87[383], line_86[381], line_85[379], line_84[377], line_83[375], line_82[373], line_81[371], line_80[369], line_79[367], line_78[365], line_77[363], line_76[361], line_75[359], line_74[357], line_73[355], line_72[353], line_71[351], line_70[349], line_69[347], line_68[345], line_67[343], line_66[341], line_65[339], line_64[337], line_63[335], line_62[333], line_61[331], line_60[329], line_59[327], line_58[325], line_57[323], line_56[321], line_55[319], line_54[317], line_53[315], line_52[313], line_51[311], line_50[309], line_49[307], line_48[305], line_47[303], line_46[301], line_45[299], line_44[297], line_43[295], line_42[293], line_41[291], line_40[289], line_39[287], line_38[285], line_37[283], line_36[281], line_35[279], line_34[277], line_33[275], line_32[273], line_31[271], line_30[269], line_29[267], line_28[265], line_27[263], line_26[261], line_25[259], line_24[257], line_23[255], line_22[253], line_21[251], line_20[249], line_19[247], line_18[245], line_17[243], line_16[241], line_15[239], line_14[237], line_13[235], line_12[233], line_11[231], line_10[229], line_9[227], line_8[225], line_7[223], line_6[221], line_5[219], line_4[217], line_3[215], line_2[213], line_1[211] };
assign col_466 = {line_128[466], line_127[464], line_126[462], line_125[460], line_124[458], line_123[456], line_122[454], line_121[452], line_120[450], line_119[448], line_118[446], line_117[444], line_116[442], line_115[440], line_114[438], line_113[436], line_112[434], line_111[432], line_110[430], line_109[428], line_108[426], line_107[424], line_106[422], line_105[420], line_104[418], line_103[416], line_102[414], line_101[412], line_100[410], line_99[408], line_98[406], line_97[404], line_96[402], line_95[400], line_94[398], line_93[396], line_92[394], line_91[392], line_90[390], line_89[388], line_88[386], line_87[384], line_86[382], line_85[380], line_84[378], line_83[376], line_82[374], line_81[372], line_80[370], line_79[368], line_78[366], line_77[364], line_76[362], line_75[360], line_74[358], line_73[356], line_72[354], line_71[352], line_70[350], line_69[348], line_68[346], line_67[344], line_66[342], line_65[340], line_64[338], line_63[336], line_62[334], line_61[332], line_60[330], line_59[328], line_58[326], line_57[324], line_56[322], line_55[320], line_54[318], line_53[316], line_52[314], line_51[312], line_50[310], line_49[308], line_48[306], line_47[304], line_46[302], line_45[300], line_44[298], line_43[296], line_42[294], line_41[292], line_40[290], line_39[288], line_38[286], line_37[284], line_36[282], line_35[280], line_34[278], line_33[276], line_32[274], line_31[272], line_30[270], line_29[268], line_28[266], line_27[264], line_26[262], line_25[260], line_24[258], line_23[256], line_22[254], line_21[252], line_20[250], line_19[248], line_18[246], line_17[244], line_16[242], line_15[240], line_14[238], line_13[236], line_12[234], line_11[232], line_10[230], line_9[228], line_8[226], line_7[224], line_6[222], line_5[220], line_4[218], line_3[216], line_2[214], line_1[212] };
assign col_467 = {line_128[467], line_127[465], line_126[463], line_125[461], line_124[459], line_123[457], line_122[455], line_121[453], line_120[451], line_119[449], line_118[447], line_117[445], line_116[443], line_115[441], line_114[439], line_113[437], line_112[435], line_111[433], line_110[431], line_109[429], line_108[427], line_107[425], line_106[423], line_105[421], line_104[419], line_103[417], line_102[415], line_101[413], line_100[411], line_99[409], line_98[407], line_97[405], line_96[403], line_95[401], line_94[399], line_93[397], line_92[395], line_91[393], line_90[391], line_89[389], line_88[387], line_87[385], line_86[383], line_85[381], line_84[379], line_83[377], line_82[375], line_81[373], line_80[371], line_79[369], line_78[367], line_77[365], line_76[363], line_75[361], line_74[359], line_73[357], line_72[355], line_71[353], line_70[351], line_69[349], line_68[347], line_67[345], line_66[343], line_65[341], line_64[339], line_63[337], line_62[335], line_61[333], line_60[331], line_59[329], line_58[327], line_57[325], line_56[323], line_55[321], line_54[319], line_53[317], line_52[315], line_51[313], line_50[311], line_49[309], line_48[307], line_47[305], line_46[303], line_45[301], line_44[299], line_43[297], line_42[295], line_41[293], line_40[291], line_39[289], line_38[287], line_37[285], line_36[283], line_35[281], line_34[279], line_33[277], line_32[275], line_31[273], line_30[271], line_29[269], line_28[267], line_27[265], line_26[263], line_25[261], line_24[259], line_23[257], line_22[255], line_21[253], line_20[251], line_19[249], line_18[247], line_17[245], line_16[243], line_15[241], line_14[239], line_13[237], line_12[235], line_11[233], line_10[231], line_9[229], line_8[227], line_7[225], line_6[223], line_5[221], line_4[219], line_3[217], line_2[215], line_1[213] };
assign col_468 = {line_128[468], line_127[466], line_126[464], line_125[462], line_124[460], line_123[458], line_122[456], line_121[454], line_120[452], line_119[450], line_118[448], line_117[446], line_116[444], line_115[442], line_114[440], line_113[438], line_112[436], line_111[434], line_110[432], line_109[430], line_108[428], line_107[426], line_106[424], line_105[422], line_104[420], line_103[418], line_102[416], line_101[414], line_100[412], line_99[410], line_98[408], line_97[406], line_96[404], line_95[402], line_94[400], line_93[398], line_92[396], line_91[394], line_90[392], line_89[390], line_88[388], line_87[386], line_86[384], line_85[382], line_84[380], line_83[378], line_82[376], line_81[374], line_80[372], line_79[370], line_78[368], line_77[366], line_76[364], line_75[362], line_74[360], line_73[358], line_72[356], line_71[354], line_70[352], line_69[350], line_68[348], line_67[346], line_66[344], line_65[342], line_64[340], line_63[338], line_62[336], line_61[334], line_60[332], line_59[330], line_58[328], line_57[326], line_56[324], line_55[322], line_54[320], line_53[318], line_52[316], line_51[314], line_50[312], line_49[310], line_48[308], line_47[306], line_46[304], line_45[302], line_44[300], line_43[298], line_42[296], line_41[294], line_40[292], line_39[290], line_38[288], line_37[286], line_36[284], line_35[282], line_34[280], line_33[278], line_32[276], line_31[274], line_30[272], line_29[270], line_28[268], line_27[266], line_26[264], line_25[262], line_24[260], line_23[258], line_22[256], line_21[254], line_20[252], line_19[250], line_18[248], line_17[246], line_16[244], line_15[242], line_14[240], line_13[238], line_12[236], line_11[234], line_10[232], line_9[230], line_8[228], line_7[226], line_6[224], line_5[222], line_4[220], line_3[218], line_2[216], line_1[214] };
assign col_469 = {line_128[469], line_127[467], line_126[465], line_125[463], line_124[461], line_123[459], line_122[457], line_121[455], line_120[453], line_119[451], line_118[449], line_117[447], line_116[445], line_115[443], line_114[441], line_113[439], line_112[437], line_111[435], line_110[433], line_109[431], line_108[429], line_107[427], line_106[425], line_105[423], line_104[421], line_103[419], line_102[417], line_101[415], line_100[413], line_99[411], line_98[409], line_97[407], line_96[405], line_95[403], line_94[401], line_93[399], line_92[397], line_91[395], line_90[393], line_89[391], line_88[389], line_87[387], line_86[385], line_85[383], line_84[381], line_83[379], line_82[377], line_81[375], line_80[373], line_79[371], line_78[369], line_77[367], line_76[365], line_75[363], line_74[361], line_73[359], line_72[357], line_71[355], line_70[353], line_69[351], line_68[349], line_67[347], line_66[345], line_65[343], line_64[341], line_63[339], line_62[337], line_61[335], line_60[333], line_59[331], line_58[329], line_57[327], line_56[325], line_55[323], line_54[321], line_53[319], line_52[317], line_51[315], line_50[313], line_49[311], line_48[309], line_47[307], line_46[305], line_45[303], line_44[301], line_43[299], line_42[297], line_41[295], line_40[293], line_39[291], line_38[289], line_37[287], line_36[285], line_35[283], line_34[281], line_33[279], line_32[277], line_31[275], line_30[273], line_29[271], line_28[269], line_27[267], line_26[265], line_25[263], line_24[261], line_23[259], line_22[257], line_21[255], line_20[253], line_19[251], line_18[249], line_17[247], line_16[245], line_15[243], line_14[241], line_13[239], line_12[237], line_11[235], line_10[233], line_9[231], line_8[229], line_7[227], line_6[225], line_5[223], line_4[221], line_3[219], line_2[217], line_1[215] };
assign col_470 = {line_128[470], line_127[468], line_126[466], line_125[464], line_124[462], line_123[460], line_122[458], line_121[456], line_120[454], line_119[452], line_118[450], line_117[448], line_116[446], line_115[444], line_114[442], line_113[440], line_112[438], line_111[436], line_110[434], line_109[432], line_108[430], line_107[428], line_106[426], line_105[424], line_104[422], line_103[420], line_102[418], line_101[416], line_100[414], line_99[412], line_98[410], line_97[408], line_96[406], line_95[404], line_94[402], line_93[400], line_92[398], line_91[396], line_90[394], line_89[392], line_88[390], line_87[388], line_86[386], line_85[384], line_84[382], line_83[380], line_82[378], line_81[376], line_80[374], line_79[372], line_78[370], line_77[368], line_76[366], line_75[364], line_74[362], line_73[360], line_72[358], line_71[356], line_70[354], line_69[352], line_68[350], line_67[348], line_66[346], line_65[344], line_64[342], line_63[340], line_62[338], line_61[336], line_60[334], line_59[332], line_58[330], line_57[328], line_56[326], line_55[324], line_54[322], line_53[320], line_52[318], line_51[316], line_50[314], line_49[312], line_48[310], line_47[308], line_46[306], line_45[304], line_44[302], line_43[300], line_42[298], line_41[296], line_40[294], line_39[292], line_38[290], line_37[288], line_36[286], line_35[284], line_34[282], line_33[280], line_32[278], line_31[276], line_30[274], line_29[272], line_28[270], line_27[268], line_26[266], line_25[264], line_24[262], line_23[260], line_22[258], line_21[256], line_20[254], line_19[252], line_18[250], line_17[248], line_16[246], line_15[244], line_14[242], line_13[240], line_12[238], line_11[236], line_10[234], line_9[232], line_8[230], line_7[228], line_6[226], line_5[224], line_4[222], line_3[220], line_2[218], line_1[216] };
assign col_471 = {line_128[471], line_127[469], line_126[467], line_125[465], line_124[463], line_123[461], line_122[459], line_121[457], line_120[455], line_119[453], line_118[451], line_117[449], line_116[447], line_115[445], line_114[443], line_113[441], line_112[439], line_111[437], line_110[435], line_109[433], line_108[431], line_107[429], line_106[427], line_105[425], line_104[423], line_103[421], line_102[419], line_101[417], line_100[415], line_99[413], line_98[411], line_97[409], line_96[407], line_95[405], line_94[403], line_93[401], line_92[399], line_91[397], line_90[395], line_89[393], line_88[391], line_87[389], line_86[387], line_85[385], line_84[383], line_83[381], line_82[379], line_81[377], line_80[375], line_79[373], line_78[371], line_77[369], line_76[367], line_75[365], line_74[363], line_73[361], line_72[359], line_71[357], line_70[355], line_69[353], line_68[351], line_67[349], line_66[347], line_65[345], line_64[343], line_63[341], line_62[339], line_61[337], line_60[335], line_59[333], line_58[331], line_57[329], line_56[327], line_55[325], line_54[323], line_53[321], line_52[319], line_51[317], line_50[315], line_49[313], line_48[311], line_47[309], line_46[307], line_45[305], line_44[303], line_43[301], line_42[299], line_41[297], line_40[295], line_39[293], line_38[291], line_37[289], line_36[287], line_35[285], line_34[283], line_33[281], line_32[279], line_31[277], line_30[275], line_29[273], line_28[271], line_27[269], line_26[267], line_25[265], line_24[263], line_23[261], line_22[259], line_21[257], line_20[255], line_19[253], line_18[251], line_17[249], line_16[247], line_15[245], line_14[243], line_13[241], line_12[239], line_11[237], line_10[235], line_9[233], line_8[231], line_7[229], line_6[227], line_5[225], line_4[223], line_3[221], line_2[219], line_1[217] };
assign col_472 = {line_128[472], line_127[470], line_126[468], line_125[466], line_124[464], line_123[462], line_122[460], line_121[458], line_120[456], line_119[454], line_118[452], line_117[450], line_116[448], line_115[446], line_114[444], line_113[442], line_112[440], line_111[438], line_110[436], line_109[434], line_108[432], line_107[430], line_106[428], line_105[426], line_104[424], line_103[422], line_102[420], line_101[418], line_100[416], line_99[414], line_98[412], line_97[410], line_96[408], line_95[406], line_94[404], line_93[402], line_92[400], line_91[398], line_90[396], line_89[394], line_88[392], line_87[390], line_86[388], line_85[386], line_84[384], line_83[382], line_82[380], line_81[378], line_80[376], line_79[374], line_78[372], line_77[370], line_76[368], line_75[366], line_74[364], line_73[362], line_72[360], line_71[358], line_70[356], line_69[354], line_68[352], line_67[350], line_66[348], line_65[346], line_64[344], line_63[342], line_62[340], line_61[338], line_60[336], line_59[334], line_58[332], line_57[330], line_56[328], line_55[326], line_54[324], line_53[322], line_52[320], line_51[318], line_50[316], line_49[314], line_48[312], line_47[310], line_46[308], line_45[306], line_44[304], line_43[302], line_42[300], line_41[298], line_40[296], line_39[294], line_38[292], line_37[290], line_36[288], line_35[286], line_34[284], line_33[282], line_32[280], line_31[278], line_30[276], line_29[274], line_28[272], line_27[270], line_26[268], line_25[266], line_24[264], line_23[262], line_22[260], line_21[258], line_20[256], line_19[254], line_18[252], line_17[250], line_16[248], line_15[246], line_14[244], line_13[242], line_12[240], line_11[238], line_10[236], line_9[234], line_8[232], line_7[230], line_6[228], line_5[226], line_4[224], line_3[222], line_2[220], line_1[218] };
assign col_473 = {line_128[473], line_127[471], line_126[469], line_125[467], line_124[465], line_123[463], line_122[461], line_121[459], line_120[457], line_119[455], line_118[453], line_117[451], line_116[449], line_115[447], line_114[445], line_113[443], line_112[441], line_111[439], line_110[437], line_109[435], line_108[433], line_107[431], line_106[429], line_105[427], line_104[425], line_103[423], line_102[421], line_101[419], line_100[417], line_99[415], line_98[413], line_97[411], line_96[409], line_95[407], line_94[405], line_93[403], line_92[401], line_91[399], line_90[397], line_89[395], line_88[393], line_87[391], line_86[389], line_85[387], line_84[385], line_83[383], line_82[381], line_81[379], line_80[377], line_79[375], line_78[373], line_77[371], line_76[369], line_75[367], line_74[365], line_73[363], line_72[361], line_71[359], line_70[357], line_69[355], line_68[353], line_67[351], line_66[349], line_65[347], line_64[345], line_63[343], line_62[341], line_61[339], line_60[337], line_59[335], line_58[333], line_57[331], line_56[329], line_55[327], line_54[325], line_53[323], line_52[321], line_51[319], line_50[317], line_49[315], line_48[313], line_47[311], line_46[309], line_45[307], line_44[305], line_43[303], line_42[301], line_41[299], line_40[297], line_39[295], line_38[293], line_37[291], line_36[289], line_35[287], line_34[285], line_33[283], line_32[281], line_31[279], line_30[277], line_29[275], line_28[273], line_27[271], line_26[269], line_25[267], line_24[265], line_23[263], line_22[261], line_21[259], line_20[257], line_19[255], line_18[253], line_17[251], line_16[249], line_15[247], line_14[245], line_13[243], line_12[241], line_11[239], line_10[237], line_9[235], line_8[233], line_7[231], line_6[229], line_5[227], line_4[225], line_3[223], line_2[221], line_1[219] };
assign col_474 = {line_128[474], line_127[472], line_126[470], line_125[468], line_124[466], line_123[464], line_122[462], line_121[460], line_120[458], line_119[456], line_118[454], line_117[452], line_116[450], line_115[448], line_114[446], line_113[444], line_112[442], line_111[440], line_110[438], line_109[436], line_108[434], line_107[432], line_106[430], line_105[428], line_104[426], line_103[424], line_102[422], line_101[420], line_100[418], line_99[416], line_98[414], line_97[412], line_96[410], line_95[408], line_94[406], line_93[404], line_92[402], line_91[400], line_90[398], line_89[396], line_88[394], line_87[392], line_86[390], line_85[388], line_84[386], line_83[384], line_82[382], line_81[380], line_80[378], line_79[376], line_78[374], line_77[372], line_76[370], line_75[368], line_74[366], line_73[364], line_72[362], line_71[360], line_70[358], line_69[356], line_68[354], line_67[352], line_66[350], line_65[348], line_64[346], line_63[344], line_62[342], line_61[340], line_60[338], line_59[336], line_58[334], line_57[332], line_56[330], line_55[328], line_54[326], line_53[324], line_52[322], line_51[320], line_50[318], line_49[316], line_48[314], line_47[312], line_46[310], line_45[308], line_44[306], line_43[304], line_42[302], line_41[300], line_40[298], line_39[296], line_38[294], line_37[292], line_36[290], line_35[288], line_34[286], line_33[284], line_32[282], line_31[280], line_30[278], line_29[276], line_28[274], line_27[272], line_26[270], line_25[268], line_24[266], line_23[264], line_22[262], line_21[260], line_20[258], line_19[256], line_18[254], line_17[252], line_16[250], line_15[248], line_14[246], line_13[244], line_12[242], line_11[240], line_10[238], line_9[236], line_8[234], line_7[232], line_6[230], line_5[228], line_4[226], line_3[224], line_2[222], line_1[220] };
assign col_475 = {line_128[475], line_127[473], line_126[471], line_125[469], line_124[467], line_123[465], line_122[463], line_121[461], line_120[459], line_119[457], line_118[455], line_117[453], line_116[451], line_115[449], line_114[447], line_113[445], line_112[443], line_111[441], line_110[439], line_109[437], line_108[435], line_107[433], line_106[431], line_105[429], line_104[427], line_103[425], line_102[423], line_101[421], line_100[419], line_99[417], line_98[415], line_97[413], line_96[411], line_95[409], line_94[407], line_93[405], line_92[403], line_91[401], line_90[399], line_89[397], line_88[395], line_87[393], line_86[391], line_85[389], line_84[387], line_83[385], line_82[383], line_81[381], line_80[379], line_79[377], line_78[375], line_77[373], line_76[371], line_75[369], line_74[367], line_73[365], line_72[363], line_71[361], line_70[359], line_69[357], line_68[355], line_67[353], line_66[351], line_65[349], line_64[347], line_63[345], line_62[343], line_61[341], line_60[339], line_59[337], line_58[335], line_57[333], line_56[331], line_55[329], line_54[327], line_53[325], line_52[323], line_51[321], line_50[319], line_49[317], line_48[315], line_47[313], line_46[311], line_45[309], line_44[307], line_43[305], line_42[303], line_41[301], line_40[299], line_39[297], line_38[295], line_37[293], line_36[291], line_35[289], line_34[287], line_33[285], line_32[283], line_31[281], line_30[279], line_29[277], line_28[275], line_27[273], line_26[271], line_25[269], line_24[267], line_23[265], line_22[263], line_21[261], line_20[259], line_19[257], line_18[255], line_17[253], line_16[251], line_15[249], line_14[247], line_13[245], line_12[243], line_11[241], line_10[239], line_9[237], line_8[235], line_7[233], line_6[231], line_5[229], line_4[227], line_3[225], line_2[223], line_1[221] };
assign col_476 = {line_128[476], line_127[474], line_126[472], line_125[470], line_124[468], line_123[466], line_122[464], line_121[462], line_120[460], line_119[458], line_118[456], line_117[454], line_116[452], line_115[450], line_114[448], line_113[446], line_112[444], line_111[442], line_110[440], line_109[438], line_108[436], line_107[434], line_106[432], line_105[430], line_104[428], line_103[426], line_102[424], line_101[422], line_100[420], line_99[418], line_98[416], line_97[414], line_96[412], line_95[410], line_94[408], line_93[406], line_92[404], line_91[402], line_90[400], line_89[398], line_88[396], line_87[394], line_86[392], line_85[390], line_84[388], line_83[386], line_82[384], line_81[382], line_80[380], line_79[378], line_78[376], line_77[374], line_76[372], line_75[370], line_74[368], line_73[366], line_72[364], line_71[362], line_70[360], line_69[358], line_68[356], line_67[354], line_66[352], line_65[350], line_64[348], line_63[346], line_62[344], line_61[342], line_60[340], line_59[338], line_58[336], line_57[334], line_56[332], line_55[330], line_54[328], line_53[326], line_52[324], line_51[322], line_50[320], line_49[318], line_48[316], line_47[314], line_46[312], line_45[310], line_44[308], line_43[306], line_42[304], line_41[302], line_40[300], line_39[298], line_38[296], line_37[294], line_36[292], line_35[290], line_34[288], line_33[286], line_32[284], line_31[282], line_30[280], line_29[278], line_28[276], line_27[274], line_26[272], line_25[270], line_24[268], line_23[266], line_22[264], line_21[262], line_20[260], line_19[258], line_18[256], line_17[254], line_16[252], line_15[250], line_14[248], line_13[246], line_12[244], line_11[242], line_10[240], line_9[238], line_8[236], line_7[234], line_6[232], line_5[230], line_4[228], line_3[226], line_2[224], line_1[222] };
assign col_477 = {line_128[477], line_127[475], line_126[473], line_125[471], line_124[469], line_123[467], line_122[465], line_121[463], line_120[461], line_119[459], line_118[457], line_117[455], line_116[453], line_115[451], line_114[449], line_113[447], line_112[445], line_111[443], line_110[441], line_109[439], line_108[437], line_107[435], line_106[433], line_105[431], line_104[429], line_103[427], line_102[425], line_101[423], line_100[421], line_99[419], line_98[417], line_97[415], line_96[413], line_95[411], line_94[409], line_93[407], line_92[405], line_91[403], line_90[401], line_89[399], line_88[397], line_87[395], line_86[393], line_85[391], line_84[389], line_83[387], line_82[385], line_81[383], line_80[381], line_79[379], line_78[377], line_77[375], line_76[373], line_75[371], line_74[369], line_73[367], line_72[365], line_71[363], line_70[361], line_69[359], line_68[357], line_67[355], line_66[353], line_65[351], line_64[349], line_63[347], line_62[345], line_61[343], line_60[341], line_59[339], line_58[337], line_57[335], line_56[333], line_55[331], line_54[329], line_53[327], line_52[325], line_51[323], line_50[321], line_49[319], line_48[317], line_47[315], line_46[313], line_45[311], line_44[309], line_43[307], line_42[305], line_41[303], line_40[301], line_39[299], line_38[297], line_37[295], line_36[293], line_35[291], line_34[289], line_33[287], line_32[285], line_31[283], line_30[281], line_29[279], line_28[277], line_27[275], line_26[273], line_25[271], line_24[269], line_23[267], line_22[265], line_21[263], line_20[261], line_19[259], line_18[257], line_17[255], line_16[253], line_15[251], line_14[249], line_13[247], line_12[245], line_11[243], line_10[241], line_9[239], line_8[237], line_7[235], line_6[233], line_5[231], line_4[229], line_3[227], line_2[225], line_1[223] };
assign col_478 = {line_128[478], line_127[476], line_126[474], line_125[472], line_124[470], line_123[468], line_122[466], line_121[464], line_120[462], line_119[460], line_118[458], line_117[456], line_116[454], line_115[452], line_114[450], line_113[448], line_112[446], line_111[444], line_110[442], line_109[440], line_108[438], line_107[436], line_106[434], line_105[432], line_104[430], line_103[428], line_102[426], line_101[424], line_100[422], line_99[420], line_98[418], line_97[416], line_96[414], line_95[412], line_94[410], line_93[408], line_92[406], line_91[404], line_90[402], line_89[400], line_88[398], line_87[396], line_86[394], line_85[392], line_84[390], line_83[388], line_82[386], line_81[384], line_80[382], line_79[380], line_78[378], line_77[376], line_76[374], line_75[372], line_74[370], line_73[368], line_72[366], line_71[364], line_70[362], line_69[360], line_68[358], line_67[356], line_66[354], line_65[352], line_64[350], line_63[348], line_62[346], line_61[344], line_60[342], line_59[340], line_58[338], line_57[336], line_56[334], line_55[332], line_54[330], line_53[328], line_52[326], line_51[324], line_50[322], line_49[320], line_48[318], line_47[316], line_46[314], line_45[312], line_44[310], line_43[308], line_42[306], line_41[304], line_40[302], line_39[300], line_38[298], line_37[296], line_36[294], line_35[292], line_34[290], line_33[288], line_32[286], line_31[284], line_30[282], line_29[280], line_28[278], line_27[276], line_26[274], line_25[272], line_24[270], line_23[268], line_22[266], line_21[264], line_20[262], line_19[260], line_18[258], line_17[256], line_16[254], line_15[252], line_14[250], line_13[248], line_12[246], line_11[244], line_10[242], line_9[240], line_8[238], line_7[236], line_6[234], line_5[232], line_4[230], line_3[228], line_2[226], line_1[224] };
assign col_479 = {line_128[479], line_127[477], line_126[475], line_125[473], line_124[471], line_123[469], line_122[467], line_121[465], line_120[463], line_119[461], line_118[459], line_117[457], line_116[455], line_115[453], line_114[451], line_113[449], line_112[447], line_111[445], line_110[443], line_109[441], line_108[439], line_107[437], line_106[435], line_105[433], line_104[431], line_103[429], line_102[427], line_101[425], line_100[423], line_99[421], line_98[419], line_97[417], line_96[415], line_95[413], line_94[411], line_93[409], line_92[407], line_91[405], line_90[403], line_89[401], line_88[399], line_87[397], line_86[395], line_85[393], line_84[391], line_83[389], line_82[387], line_81[385], line_80[383], line_79[381], line_78[379], line_77[377], line_76[375], line_75[373], line_74[371], line_73[369], line_72[367], line_71[365], line_70[363], line_69[361], line_68[359], line_67[357], line_66[355], line_65[353], line_64[351], line_63[349], line_62[347], line_61[345], line_60[343], line_59[341], line_58[339], line_57[337], line_56[335], line_55[333], line_54[331], line_53[329], line_52[327], line_51[325], line_50[323], line_49[321], line_48[319], line_47[317], line_46[315], line_45[313], line_44[311], line_43[309], line_42[307], line_41[305], line_40[303], line_39[301], line_38[299], line_37[297], line_36[295], line_35[293], line_34[291], line_33[289], line_32[287], line_31[285], line_30[283], line_29[281], line_28[279], line_27[277], line_26[275], line_25[273], line_24[271], line_23[269], line_22[267], line_21[265], line_20[263], line_19[261], line_18[259], line_17[257], line_16[255], line_15[253], line_14[251], line_13[249], line_12[247], line_11[245], line_10[243], line_9[241], line_8[239], line_7[237], line_6[235], line_5[233], line_4[231], line_3[229], line_2[227], line_1[225] };
assign col_480 = {line_128[480], line_127[478], line_126[476], line_125[474], line_124[472], line_123[470], line_122[468], line_121[466], line_120[464], line_119[462], line_118[460], line_117[458], line_116[456], line_115[454], line_114[452], line_113[450], line_112[448], line_111[446], line_110[444], line_109[442], line_108[440], line_107[438], line_106[436], line_105[434], line_104[432], line_103[430], line_102[428], line_101[426], line_100[424], line_99[422], line_98[420], line_97[418], line_96[416], line_95[414], line_94[412], line_93[410], line_92[408], line_91[406], line_90[404], line_89[402], line_88[400], line_87[398], line_86[396], line_85[394], line_84[392], line_83[390], line_82[388], line_81[386], line_80[384], line_79[382], line_78[380], line_77[378], line_76[376], line_75[374], line_74[372], line_73[370], line_72[368], line_71[366], line_70[364], line_69[362], line_68[360], line_67[358], line_66[356], line_65[354], line_64[352], line_63[350], line_62[348], line_61[346], line_60[344], line_59[342], line_58[340], line_57[338], line_56[336], line_55[334], line_54[332], line_53[330], line_52[328], line_51[326], line_50[324], line_49[322], line_48[320], line_47[318], line_46[316], line_45[314], line_44[312], line_43[310], line_42[308], line_41[306], line_40[304], line_39[302], line_38[300], line_37[298], line_36[296], line_35[294], line_34[292], line_33[290], line_32[288], line_31[286], line_30[284], line_29[282], line_28[280], line_27[278], line_26[276], line_25[274], line_24[272], line_23[270], line_22[268], line_21[266], line_20[264], line_19[262], line_18[260], line_17[258], line_16[256], line_15[254], line_14[252], line_13[250], line_12[248], line_11[246], line_10[244], line_9[242], line_8[240], line_7[238], line_6[236], line_5[234], line_4[232], line_3[230], line_2[228], line_1[226] };
assign col_481 = {line_128[481], line_127[479], line_126[477], line_125[475], line_124[473], line_123[471], line_122[469], line_121[467], line_120[465], line_119[463], line_118[461], line_117[459], line_116[457], line_115[455], line_114[453], line_113[451], line_112[449], line_111[447], line_110[445], line_109[443], line_108[441], line_107[439], line_106[437], line_105[435], line_104[433], line_103[431], line_102[429], line_101[427], line_100[425], line_99[423], line_98[421], line_97[419], line_96[417], line_95[415], line_94[413], line_93[411], line_92[409], line_91[407], line_90[405], line_89[403], line_88[401], line_87[399], line_86[397], line_85[395], line_84[393], line_83[391], line_82[389], line_81[387], line_80[385], line_79[383], line_78[381], line_77[379], line_76[377], line_75[375], line_74[373], line_73[371], line_72[369], line_71[367], line_70[365], line_69[363], line_68[361], line_67[359], line_66[357], line_65[355], line_64[353], line_63[351], line_62[349], line_61[347], line_60[345], line_59[343], line_58[341], line_57[339], line_56[337], line_55[335], line_54[333], line_53[331], line_52[329], line_51[327], line_50[325], line_49[323], line_48[321], line_47[319], line_46[317], line_45[315], line_44[313], line_43[311], line_42[309], line_41[307], line_40[305], line_39[303], line_38[301], line_37[299], line_36[297], line_35[295], line_34[293], line_33[291], line_32[289], line_31[287], line_30[285], line_29[283], line_28[281], line_27[279], line_26[277], line_25[275], line_24[273], line_23[271], line_22[269], line_21[267], line_20[265], line_19[263], line_18[261], line_17[259], line_16[257], line_15[255], line_14[253], line_13[251], line_12[249], line_11[247], line_10[245], line_9[243], line_8[241], line_7[239], line_6[237], line_5[235], line_4[233], line_3[231], line_2[229], line_1[227] };
assign col_482 = {line_128[482], line_127[480], line_126[478], line_125[476], line_124[474], line_123[472], line_122[470], line_121[468], line_120[466], line_119[464], line_118[462], line_117[460], line_116[458], line_115[456], line_114[454], line_113[452], line_112[450], line_111[448], line_110[446], line_109[444], line_108[442], line_107[440], line_106[438], line_105[436], line_104[434], line_103[432], line_102[430], line_101[428], line_100[426], line_99[424], line_98[422], line_97[420], line_96[418], line_95[416], line_94[414], line_93[412], line_92[410], line_91[408], line_90[406], line_89[404], line_88[402], line_87[400], line_86[398], line_85[396], line_84[394], line_83[392], line_82[390], line_81[388], line_80[386], line_79[384], line_78[382], line_77[380], line_76[378], line_75[376], line_74[374], line_73[372], line_72[370], line_71[368], line_70[366], line_69[364], line_68[362], line_67[360], line_66[358], line_65[356], line_64[354], line_63[352], line_62[350], line_61[348], line_60[346], line_59[344], line_58[342], line_57[340], line_56[338], line_55[336], line_54[334], line_53[332], line_52[330], line_51[328], line_50[326], line_49[324], line_48[322], line_47[320], line_46[318], line_45[316], line_44[314], line_43[312], line_42[310], line_41[308], line_40[306], line_39[304], line_38[302], line_37[300], line_36[298], line_35[296], line_34[294], line_33[292], line_32[290], line_31[288], line_30[286], line_29[284], line_28[282], line_27[280], line_26[278], line_25[276], line_24[274], line_23[272], line_22[270], line_21[268], line_20[266], line_19[264], line_18[262], line_17[260], line_16[258], line_15[256], line_14[254], line_13[252], line_12[250], line_11[248], line_10[246], line_9[244], line_8[242], line_7[240], line_6[238], line_5[236], line_4[234], line_3[232], line_2[230], line_1[228] };
assign col_483 = {line_128[483], line_127[481], line_126[479], line_125[477], line_124[475], line_123[473], line_122[471], line_121[469], line_120[467], line_119[465], line_118[463], line_117[461], line_116[459], line_115[457], line_114[455], line_113[453], line_112[451], line_111[449], line_110[447], line_109[445], line_108[443], line_107[441], line_106[439], line_105[437], line_104[435], line_103[433], line_102[431], line_101[429], line_100[427], line_99[425], line_98[423], line_97[421], line_96[419], line_95[417], line_94[415], line_93[413], line_92[411], line_91[409], line_90[407], line_89[405], line_88[403], line_87[401], line_86[399], line_85[397], line_84[395], line_83[393], line_82[391], line_81[389], line_80[387], line_79[385], line_78[383], line_77[381], line_76[379], line_75[377], line_74[375], line_73[373], line_72[371], line_71[369], line_70[367], line_69[365], line_68[363], line_67[361], line_66[359], line_65[357], line_64[355], line_63[353], line_62[351], line_61[349], line_60[347], line_59[345], line_58[343], line_57[341], line_56[339], line_55[337], line_54[335], line_53[333], line_52[331], line_51[329], line_50[327], line_49[325], line_48[323], line_47[321], line_46[319], line_45[317], line_44[315], line_43[313], line_42[311], line_41[309], line_40[307], line_39[305], line_38[303], line_37[301], line_36[299], line_35[297], line_34[295], line_33[293], line_32[291], line_31[289], line_30[287], line_29[285], line_28[283], line_27[281], line_26[279], line_25[277], line_24[275], line_23[273], line_22[271], line_21[269], line_20[267], line_19[265], line_18[263], line_17[261], line_16[259], line_15[257], line_14[255], line_13[253], line_12[251], line_11[249], line_10[247], line_9[245], line_8[243], line_7[241], line_6[239], line_5[237], line_4[235], line_3[233], line_2[231], line_1[229] };
assign col_484 = {line_128[484], line_127[482], line_126[480], line_125[478], line_124[476], line_123[474], line_122[472], line_121[470], line_120[468], line_119[466], line_118[464], line_117[462], line_116[460], line_115[458], line_114[456], line_113[454], line_112[452], line_111[450], line_110[448], line_109[446], line_108[444], line_107[442], line_106[440], line_105[438], line_104[436], line_103[434], line_102[432], line_101[430], line_100[428], line_99[426], line_98[424], line_97[422], line_96[420], line_95[418], line_94[416], line_93[414], line_92[412], line_91[410], line_90[408], line_89[406], line_88[404], line_87[402], line_86[400], line_85[398], line_84[396], line_83[394], line_82[392], line_81[390], line_80[388], line_79[386], line_78[384], line_77[382], line_76[380], line_75[378], line_74[376], line_73[374], line_72[372], line_71[370], line_70[368], line_69[366], line_68[364], line_67[362], line_66[360], line_65[358], line_64[356], line_63[354], line_62[352], line_61[350], line_60[348], line_59[346], line_58[344], line_57[342], line_56[340], line_55[338], line_54[336], line_53[334], line_52[332], line_51[330], line_50[328], line_49[326], line_48[324], line_47[322], line_46[320], line_45[318], line_44[316], line_43[314], line_42[312], line_41[310], line_40[308], line_39[306], line_38[304], line_37[302], line_36[300], line_35[298], line_34[296], line_33[294], line_32[292], line_31[290], line_30[288], line_29[286], line_28[284], line_27[282], line_26[280], line_25[278], line_24[276], line_23[274], line_22[272], line_21[270], line_20[268], line_19[266], line_18[264], line_17[262], line_16[260], line_15[258], line_14[256], line_13[254], line_12[252], line_11[250], line_10[248], line_9[246], line_8[244], line_7[242], line_6[240], line_5[238], line_4[236], line_3[234], line_2[232], line_1[230] };
assign col_485 = {line_128[485], line_127[483], line_126[481], line_125[479], line_124[477], line_123[475], line_122[473], line_121[471], line_120[469], line_119[467], line_118[465], line_117[463], line_116[461], line_115[459], line_114[457], line_113[455], line_112[453], line_111[451], line_110[449], line_109[447], line_108[445], line_107[443], line_106[441], line_105[439], line_104[437], line_103[435], line_102[433], line_101[431], line_100[429], line_99[427], line_98[425], line_97[423], line_96[421], line_95[419], line_94[417], line_93[415], line_92[413], line_91[411], line_90[409], line_89[407], line_88[405], line_87[403], line_86[401], line_85[399], line_84[397], line_83[395], line_82[393], line_81[391], line_80[389], line_79[387], line_78[385], line_77[383], line_76[381], line_75[379], line_74[377], line_73[375], line_72[373], line_71[371], line_70[369], line_69[367], line_68[365], line_67[363], line_66[361], line_65[359], line_64[357], line_63[355], line_62[353], line_61[351], line_60[349], line_59[347], line_58[345], line_57[343], line_56[341], line_55[339], line_54[337], line_53[335], line_52[333], line_51[331], line_50[329], line_49[327], line_48[325], line_47[323], line_46[321], line_45[319], line_44[317], line_43[315], line_42[313], line_41[311], line_40[309], line_39[307], line_38[305], line_37[303], line_36[301], line_35[299], line_34[297], line_33[295], line_32[293], line_31[291], line_30[289], line_29[287], line_28[285], line_27[283], line_26[281], line_25[279], line_24[277], line_23[275], line_22[273], line_21[271], line_20[269], line_19[267], line_18[265], line_17[263], line_16[261], line_15[259], line_14[257], line_13[255], line_12[253], line_11[251], line_10[249], line_9[247], line_8[245], line_7[243], line_6[241], line_5[239], line_4[237], line_3[235], line_2[233], line_1[231] };
assign col_486 = {line_128[486], line_127[484], line_126[482], line_125[480], line_124[478], line_123[476], line_122[474], line_121[472], line_120[470], line_119[468], line_118[466], line_117[464], line_116[462], line_115[460], line_114[458], line_113[456], line_112[454], line_111[452], line_110[450], line_109[448], line_108[446], line_107[444], line_106[442], line_105[440], line_104[438], line_103[436], line_102[434], line_101[432], line_100[430], line_99[428], line_98[426], line_97[424], line_96[422], line_95[420], line_94[418], line_93[416], line_92[414], line_91[412], line_90[410], line_89[408], line_88[406], line_87[404], line_86[402], line_85[400], line_84[398], line_83[396], line_82[394], line_81[392], line_80[390], line_79[388], line_78[386], line_77[384], line_76[382], line_75[380], line_74[378], line_73[376], line_72[374], line_71[372], line_70[370], line_69[368], line_68[366], line_67[364], line_66[362], line_65[360], line_64[358], line_63[356], line_62[354], line_61[352], line_60[350], line_59[348], line_58[346], line_57[344], line_56[342], line_55[340], line_54[338], line_53[336], line_52[334], line_51[332], line_50[330], line_49[328], line_48[326], line_47[324], line_46[322], line_45[320], line_44[318], line_43[316], line_42[314], line_41[312], line_40[310], line_39[308], line_38[306], line_37[304], line_36[302], line_35[300], line_34[298], line_33[296], line_32[294], line_31[292], line_30[290], line_29[288], line_28[286], line_27[284], line_26[282], line_25[280], line_24[278], line_23[276], line_22[274], line_21[272], line_20[270], line_19[268], line_18[266], line_17[264], line_16[262], line_15[260], line_14[258], line_13[256], line_12[254], line_11[252], line_10[250], line_9[248], line_8[246], line_7[244], line_6[242], line_5[240], line_4[238], line_3[236], line_2[234], line_1[232] };
assign col_487 = {line_128[487], line_127[485], line_126[483], line_125[481], line_124[479], line_123[477], line_122[475], line_121[473], line_120[471], line_119[469], line_118[467], line_117[465], line_116[463], line_115[461], line_114[459], line_113[457], line_112[455], line_111[453], line_110[451], line_109[449], line_108[447], line_107[445], line_106[443], line_105[441], line_104[439], line_103[437], line_102[435], line_101[433], line_100[431], line_99[429], line_98[427], line_97[425], line_96[423], line_95[421], line_94[419], line_93[417], line_92[415], line_91[413], line_90[411], line_89[409], line_88[407], line_87[405], line_86[403], line_85[401], line_84[399], line_83[397], line_82[395], line_81[393], line_80[391], line_79[389], line_78[387], line_77[385], line_76[383], line_75[381], line_74[379], line_73[377], line_72[375], line_71[373], line_70[371], line_69[369], line_68[367], line_67[365], line_66[363], line_65[361], line_64[359], line_63[357], line_62[355], line_61[353], line_60[351], line_59[349], line_58[347], line_57[345], line_56[343], line_55[341], line_54[339], line_53[337], line_52[335], line_51[333], line_50[331], line_49[329], line_48[327], line_47[325], line_46[323], line_45[321], line_44[319], line_43[317], line_42[315], line_41[313], line_40[311], line_39[309], line_38[307], line_37[305], line_36[303], line_35[301], line_34[299], line_33[297], line_32[295], line_31[293], line_30[291], line_29[289], line_28[287], line_27[285], line_26[283], line_25[281], line_24[279], line_23[277], line_22[275], line_21[273], line_20[271], line_19[269], line_18[267], line_17[265], line_16[263], line_15[261], line_14[259], line_13[257], line_12[255], line_11[253], line_10[251], line_9[249], line_8[247], line_7[245], line_6[243], line_5[241], line_4[239], line_3[237], line_2[235], line_1[233] };
assign col_488 = {line_128[488], line_127[486], line_126[484], line_125[482], line_124[480], line_123[478], line_122[476], line_121[474], line_120[472], line_119[470], line_118[468], line_117[466], line_116[464], line_115[462], line_114[460], line_113[458], line_112[456], line_111[454], line_110[452], line_109[450], line_108[448], line_107[446], line_106[444], line_105[442], line_104[440], line_103[438], line_102[436], line_101[434], line_100[432], line_99[430], line_98[428], line_97[426], line_96[424], line_95[422], line_94[420], line_93[418], line_92[416], line_91[414], line_90[412], line_89[410], line_88[408], line_87[406], line_86[404], line_85[402], line_84[400], line_83[398], line_82[396], line_81[394], line_80[392], line_79[390], line_78[388], line_77[386], line_76[384], line_75[382], line_74[380], line_73[378], line_72[376], line_71[374], line_70[372], line_69[370], line_68[368], line_67[366], line_66[364], line_65[362], line_64[360], line_63[358], line_62[356], line_61[354], line_60[352], line_59[350], line_58[348], line_57[346], line_56[344], line_55[342], line_54[340], line_53[338], line_52[336], line_51[334], line_50[332], line_49[330], line_48[328], line_47[326], line_46[324], line_45[322], line_44[320], line_43[318], line_42[316], line_41[314], line_40[312], line_39[310], line_38[308], line_37[306], line_36[304], line_35[302], line_34[300], line_33[298], line_32[296], line_31[294], line_30[292], line_29[290], line_28[288], line_27[286], line_26[284], line_25[282], line_24[280], line_23[278], line_22[276], line_21[274], line_20[272], line_19[270], line_18[268], line_17[266], line_16[264], line_15[262], line_14[260], line_13[258], line_12[256], line_11[254], line_10[252], line_9[250], line_8[248], line_7[246], line_6[244], line_5[242], line_4[240], line_3[238], line_2[236], line_1[234] };
assign col_489 = {line_128[489], line_127[487], line_126[485], line_125[483], line_124[481], line_123[479], line_122[477], line_121[475], line_120[473], line_119[471], line_118[469], line_117[467], line_116[465], line_115[463], line_114[461], line_113[459], line_112[457], line_111[455], line_110[453], line_109[451], line_108[449], line_107[447], line_106[445], line_105[443], line_104[441], line_103[439], line_102[437], line_101[435], line_100[433], line_99[431], line_98[429], line_97[427], line_96[425], line_95[423], line_94[421], line_93[419], line_92[417], line_91[415], line_90[413], line_89[411], line_88[409], line_87[407], line_86[405], line_85[403], line_84[401], line_83[399], line_82[397], line_81[395], line_80[393], line_79[391], line_78[389], line_77[387], line_76[385], line_75[383], line_74[381], line_73[379], line_72[377], line_71[375], line_70[373], line_69[371], line_68[369], line_67[367], line_66[365], line_65[363], line_64[361], line_63[359], line_62[357], line_61[355], line_60[353], line_59[351], line_58[349], line_57[347], line_56[345], line_55[343], line_54[341], line_53[339], line_52[337], line_51[335], line_50[333], line_49[331], line_48[329], line_47[327], line_46[325], line_45[323], line_44[321], line_43[319], line_42[317], line_41[315], line_40[313], line_39[311], line_38[309], line_37[307], line_36[305], line_35[303], line_34[301], line_33[299], line_32[297], line_31[295], line_30[293], line_29[291], line_28[289], line_27[287], line_26[285], line_25[283], line_24[281], line_23[279], line_22[277], line_21[275], line_20[273], line_19[271], line_18[269], line_17[267], line_16[265], line_15[263], line_14[261], line_13[259], line_12[257], line_11[255], line_10[253], line_9[251], line_8[249], line_7[247], line_6[245], line_5[243], line_4[241], line_3[239], line_2[237], line_1[235] };
assign col_490 = {line_128[490], line_127[488], line_126[486], line_125[484], line_124[482], line_123[480], line_122[478], line_121[476], line_120[474], line_119[472], line_118[470], line_117[468], line_116[466], line_115[464], line_114[462], line_113[460], line_112[458], line_111[456], line_110[454], line_109[452], line_108[450], line_107[448], line_106[446], line_105[444], line_104[442], line_103[440], line_102[438], line_101[436], line_100[434], line_99[432], line_98[430], line_97[428], line_96[426], line_95[424], line_94[422], line_93[420], line_92[418], line_91[416], line_90[414], line_89[412], line_88[410], line_87[408], line_86[406], line_85[404], line_84[402], line_83[400], line_82[398], line_81[396], line_80[394], line_79[392], line_78[390], line_77[388], line_76[386], line_75[384], line_74[382], line_73[380], line_72[378], line_71[376], line_70[374], line_69[372], line_68[370], line_67[368], line_66[366], line_65[364], line_64[362], line_63[360], line_62[358], line_61[356], line_60[354], line_59[352], line_58[350], line_57[348], line_56[346], line_55[344], line_54[342], line_53[340], line_52[338], line_51[336], line_50[334], line_49[332], line_48[330], line_47[328], line_46[326], line_45[324], line_44[322], line_43[320], line_42[318], line_41[316], line_40[314], line_39[312], line_38[310], line_37[308], line_36[306], line_35[304], line_34[302], line_33[300], line_32[298], line_31[296], line_30[294], line_29[292], line_28[290], line_27[288], line_26[286], line_25[284], line_24[282], line_23[280], line_22[278], line_21[276], line_20[274], line_19[272], line_18[270], line_17[268], line_16[266], line_15[264], line_14[262], line_13[260], line_12[258], line_11[256], line_10[254], line_9[252], line_8[250], line_7[248], line_6[246], line_5[244], line_4[242], line_3[240], line_2[238], line_1[236] };
assign col_491 = {line_128[491], line_127[489], line_126[487], line_125[485], line_124[483], line_123[481], line_122[479], line_121[477], line_120[475], line_119[473], line_118[471], line_117[469], line_116[467], line_115[465], line_114[463], line_113[461], line_112[459], line_111[457], line_110[455], line_109[453], line_108[451], line_107[449], line_106[447], line_105[445], line_104[443], line_103[441], line_102[439], line_101[437], line_100[435], line_99[433], line_98[431], line_97[429], line_96[427], line_95[425], line_94[423], line_93[421], line_92[419], line_91[417], line_90[415], line_89[413], line_88[411], line_87[409], line_86[407], line_85[405], line_84[403], line_83[401], line_82[399], line_81[397], line_80[395], line_79[393], line_78[391], line_77[389], line_76[387], line_75[385], line_74[383], line_73[381], line_72[379], line_71[377], line_70[375], line_69[373], line_68[371], line_67[369], line_66[367], line_65[365], line_64[363], line_63[361], line_62[359], line_61[357], line_60[355], line_59[353], line_58[351], line_57[349], line_56[347], line_55[345], line_54[343], line_53[341], line_52[339], line_51[337], line_50[335], line_49[333], line_48[331], line_47[329], line_46[327], line_45[325], line_44[323], line_43[321], line_42[319], line_41[317], line_40[315], line_39[313], line_38[311], line_37[309], line_36[307], line_35[305], line_34[303], line_33[301], line_32[299], line_31[297], line_30[295], line_29[293], line_28[291], line_27[289], line_26[287], line_25[285], line_24[283], line_23[281], line_22[279], line_21[277], line_20[275], line_19[273], line_18[271], line_17[269], line_16[267], line_15[265], line_14[263], line_13[261], line_12[259], line_11[257], line_10[255], line_9[253], line_8[251], line_7[249], line_6[247], line_5[245], line_4[243], line_3[241], line_2[239], line_1[237] };
assign col_492 = {line_128[492], line_127[490], line_126[488], line_125[486], line_124[484], line_123[482], line_122[480], line_121[478], line_120[476], line_119[474], line_118[472], line_117[470], line_116[468], line_115[466], line_114[464], line_113[462], line_112[460], line_111[458], line_110[456], line_109[454], line_108[452], line_107[450], line_106[448], line_105[446], line_104[444], line_103[442], line_102[440], line_101[438], line_100[436], line_99[434], line_98[432], line_97[430], line_96[428], line_95[426], line_94[424], line_93[422], line_92[420], line_91[418], line_90[416], line_89[414], line_88[412], line_87[410], line_86[408], line_85[406], line_84[404], line_83[402], line_82[400], line_81[398], line_80[396], line_79[394], line_78[392], line_77[390], line_76[388], line_75[386], line_74[384], line_73[382], line_72[380], line_71[378], line_70[376], line_69[374], line_68[372], line_67[370], line_66[368], line_65[366], line_64[364], line_63[362], line_62[360], line_61[358], line_60[356], line_59[354], line_58[352], line_57[350], line_56[348], line_55[346], line_54[344], line_53[342], line_52[340], line_51[338], line_50[336], line_49[334], line_48[332], line_47[330], line_46[328], line_45[326], line_44[324], line_43[322], line_42[320], line_41[318], line_40[316], line_39[314], line_38[312], line_37[310], line_36[308], line_35[306], line_34[304], line_33[302], line_32[300], line_31[298], line_30[296], line_29[294], line_28[292], line_27[290], line_26[288], line_25[286], line_24[284], line_23[282], line_22[280], line_21[278], line_20[276], line_19[274], line_18[272], line_17[270], line_16[268], line_15[266], line_14[264], line_13[262], line_12[260], line_11[258], line_10[256], line_9[254], line_8[252], line_7[250], line_6[248], line_5[246], line_4[244], line_3[242], line_2[240], line_1[238] };
assign col_493 = {line_128[493], line_127[491], line_126[489], line_125[487], line_124[485], line_123[483], line_122[481], line_121[479], line_120[477], line_119[475], line_118[473], line_117[471], line_116[469], line_115[467], line_114[465], line_113[463], line_112[461], line_111[459], line_110[457], line_109[455], line_108[453], line_107[451], line_106[449], line_105[447], line_104[445], line_103[443], line_102[441], line_101[439], line_100[437], line_99[435], line_98[433], line_97[431], line_96[429], line_95[427], line_94[425], line_93[423], line_92[421], line_91[419], line_90[417], line_89[415], line_88[413], line_87[411], line_86[409], line_85[407], line_84[405], line_83[403], line_82[401], line_81[399], line_80[397], line_79[395], line_78[393], line_77[391], line_76[389], line_75[387], line_74[385], line_73[383], line_72[381], line_71[379], line_70[377], line_69[375], line_68[373], line_67[371], line_66[369], line_65[367], line_64[365], line_63[363], line_62[361], line_61[359], line_60[357], line_59[355], line_58[353], line_57[351], line_56[349], line_55[347], line_54[345], line_53[343], line_52[341], line_51[339], line_50[337], line_49[335], line_48[333], line_47[331], line_46[329], line_45[327], line_44[325], line_43[323], line_42[321], line_41[319], line_40[317], line_39[315], line_38[313], line_37[311], line_36[309], line_35[307], line_34[305], line_33[303], line_32[301], line_31[299], line_30[297], line_29[295], line_28[293], line_27[291], line_26[289], line_25[287], line_24[285], line_23[283], line_22[281], line_21[279], line_20[277], line_19[275], line_18[273], line_17[271], line_16[269], line_15[267], line_14[265], line_13[263], line_12[261], line_11[259], line_10[257], line_9[255], line_8[253], line_7[251], line_6[249], line_5[247], line_4[245], line_3[243], line_2[241], line_1[239] };
assign col_494 = {line_128[494], line_127[492], line_126[490], line_125[488], line_124[486], line_123[484], line_122[482], line_121[480], line_120[478], line_119[476], line_118[474], line_117[472], line_116[470], line_115[468], line_114[466], line_113[464], line_112[462], line_111[460], line_110[458], line_109[456], line_108[454], line_107[452], line_106[450], line_105[448], line_104[446], line_103[444], line_102[442], line_101[440], line_100[438], line_99[436], line_98[434], line_97[432], line_96[430], line_95[428], line_94[426], line_93[424], line_92[422], line_91[420], line_90[418], line_89[416], line_88[414], line_87[412], line_86[410], line_85[408], line_84[406], line_83[404], line_82[402], line_81[400], line_80[398], line_79[396], line_78[394], line_77[392], line_76[390], line_75[388], line_74[386], line_73[384], line_72[382], line_71[380], line_70[378], line_69[376], line_68[374], line_67[372], line_66[370], line_65[368], line_64[366], line_63[364], line_62[362], line_61[360], line_60[358], line_59[356], line_58[354], line_57[352], line_56[350], line_55[348], line_54[346], line_53[344], line_52[342], line_51[340], line_50[338], line_49[336], line_48[334], line_47[332], line_46[330], line_45[328], line_44[326], line_43[324], line_42[322], line_41[320], line_40[318], line_39[316], line_38[314], line_37[312], line_36[310], line_35[308], line_34[306], line_33[304], line_32[302], line_31[300], line_30[298], line_29[296], line_28[294], line_27[292], line_26[290], line_25[288], line_24[286], line_23[284], line_22[282], line_21[280], line_20[278], line_19[276], line_18[274], line_17[272], line_16[270], line_15[268], line_14[266], line_13[264], line_12[262], line_11[260], line_10[258], line_9[256], line_8[254], line_7[252], line_6[250], line_5[248], line_4[246], line_3[244], line_2[242], line_1[240] };
assign col_495 = {line_128[495], line_127[493], line_126[491], line_125[489], line_124[487], line_123[485], line_122[483], line_121[481], line_120[479], line_119[477], line_118[475], line_117[473], line_116[471], line_115[469], line_114[467], line_113[465], line_112[463], line_111[461], line_110[459], line_109[457], line_108[455], line_107[453], line_106[451], line_105[449], line_104[447], line_103[445], line_102[443], line_101[441], line_100[439], line_99[437], line_98[435], line_97[433], line_96[431], line_95[429], line_94[427], line_93[425], line_92[423], line_91[421], line_90[419], line_89[417], line_88[415], line_87[413], line_86[411], line_85[409], line_84[407], line_83[405], line_82[403], line_81[401], line_80[399], line_79[397], line_78[395], line_77[393], line_76[391], line_75[389], line_74[387], line_73[385], line_72[383], line_71[381], line_70[379], line_69[377], line_68[375], line_67[373], line_66[371], line_65[369], line_64[367], line_63[365], line_62[363], line_61[361], line_60[359], line_59[357], line_58[355], line_57[353], line_56[351], line_55[349], line_54[347], line_53[345], line_52[343], line_51[341], line_50[339], line_49[337], line_48[335], line_47[333], line_46[331], line_45[329], line_44[327], line_43[325], line_42[323], line_41[321], line_40[319], line_39[317], line_38[315], line_37[313], line_36[311], line_35[309], line_34[307], line_33[305], line_32[303], line_31[301], line_30[299], line_29[297], line_28[295], line_27[293], line_26[291], line_25[289], line_24[287], line_23[285], line_22[283], line_21[281], line_20[279], line_19[277], line_18[275], line_17[273], line_16[271], line_15[269], line_14[267], line_13[265], line_12[263], line_11[261], line_10[259], line_9[257], line_8[255], line_7[253], line_6[251], line_5[249], line_4[247], line_3[245], line_2[243], line_1[241] };
assign col_496 = {line_128[496], line_127[494], line_126[492], line_125[490], line_124[488], line_123[486], line_122[484], line_121[482], line_120[480], line_119[478], line_118[476], line_117[474], line_116[472], line_115[470], line_114[468], line_113[466], line_112[464], line_111[462], line_110[460], line_109[458], line_108[456], line_107[454], line_106[452], line_105[450], line_104[448], line_103[446], line_102[444], line_101[442], line_100[440], line_99[438], line_98[436], line_97[434], line_96[432], line_95[430], line_94[428], line_93[426], line_92[424], line_91[422], line_90[420], line_89[418], line_88[416], line_87[414], line_86[412], line_85[410], line_84[408], line_83[406], line_82[404], line_81[402], line_80[400], line_79[398], line_78[396], line_77[394], line_76[392], line_75[390], line_74[388], line_73[386], line_72[384], line_71[382], line_70[380], line_69[378], line_68[376], line_67[374], line_66[372], line_65[370], line_64[368], line_63[366], line_62[364], line_61[362], line_60[360], line_59[358], line_58[356], line_57[354], line_56[352], line_55[350], line_54[348], line_53[346], line_52[344], line_51[342], line_50[340], line_49[338], line_48[336], line_47[334], line_46[332], line_45[330], line_44[328], line_43[326], line_42[324], line_41[322], line_40[320], line_39[318], line_38[316], line_37[314], line_36[312], line_35[310], line_34[308], line_33[306], line_32[304], line_31[302], line_30[300], line_29[298], line_28[296], line_27[294], line_26[292], line_25[290], line_24[288], line_23[286], line_22[284], line_21[282], line_20[280], line_19[278], line_18[276], line_17[274], line_16[272], line_15[270], line_14[268], line_13[266], line_12[264], line_11[262], line_10[260], line_9[258], line_8[256], line_7[254], line_6[252], line_5[250], line_4[248], line_3[246], line_2[244], line_1[242] };
assign col_497 = {line_128[497], line_127[495], line_126[493], line_125[491], line_124[489], line_123[487], line_122[485], line_121[483], line_120[481], line_119[479], line_118[477], line_117[475], line_116[473], line_115[471], line_114[469], line_113[467], line_112[465], line_111[463], line_110[461], line_109[459], line_108[457], line_107[455], line_106[453], line_105[451], line_104[449], line_103[447], line_102[445], line_101[443], line_100[441], line_99[439], line_98[437], line_97[435], line_96[433], line_95[431], line_94[429], line_93[427], line_92[425], line_91[423], line_90[421], line_89[419], line_88[417], line_87[415], line_86[413], line_85[411], line_84[409], line_83[407], line_82[405], line_81[403], line_80[401], line_79[399], line_78[397], line_77[395], line_76[393], line_75[391], line_74[389], line_73[387], line_72[385], line_71[383], line_70[381], line_69[379], line_68[377], line_67[375], line_66[373], line_65[371], line_64[369], line_63[367], line_62[365], line_61[363], line_60[361], line_59[359], line_58[357], line_57[355], line_56[353], line_55[351], line_54[349], line_53[347], line_52[345], line_51[343], line_50[341], line_49[339], line_48[337], line_47[335], line_46[333], line_45[331], line_44[329], line_43[327], line_42[325], line_41[323], line_40[321], line_39[319], line_38[317], line_37[315], line_36[313], line_35[311], line_34[309], line_33[307], line_32[305], line_31[303], line_30[301], line_29[299], line_28[297], line_27[295], line_26[293], line_25[291], line_24[289], line_23[287], line_22[285], line_21[283], line_20[281], line_19[279], line_18[277], line_17[275], line_16[273], line_15[271], line_14[269], line_13[267], line_12[265], line_11[263], line_10[261], line_9[259], line_8[257], line_7[255], line_6[253], line_5[251], line_4[249], line_3[247], line_2[245], line_1[243] };
assign col_498 = {line_128[498], line_127[496], line_126[494], line_125[492], line_124[490], line_123[488], line_122[486], line_121[484], line_120[482], line_119[480], line_118[478], line_117[476], line_116[474], line_115[472], line_114[470], line_113[468], line_112[466], line_111[464], line_110[462], line_109[460], line_108[458], line_107[456], line_106[454], line_105[452], line_104[450], line_103[448], line_102[446], line_101[444], line_100[442], line_99[440], line_98[438], line_97[436], line_96[434], line_95[432], line_94[430], line_93[428], line_92[426], line_91[424], line_90[422], line_89[420], line_88[418], line_87[416], line_86[414], line_85[412], line_84[410], line_83[408], line_82[406], line_81[404], line_80[402], line_79[400], line_78[398], line_77[396], line_76[394], line_75[392], line_74[390], line_73[388], line_72[386], line_71[384], line_70[382], line_69[380], line_68[378], line_67[376], line_66[374], line_65[372], line_64[370], line_63[368], line_62[366], line_61[364], line_60[362], line_59[360], line_58[358], line_57[356], line_56[354], line_55[352], line_54[350], line_53[348], line_52[346], line_51[344], line_50[342], line_49[340], line_48[338], line_47[336], line_46[334], line_45[332], line_44[330], line_43[328], line_42[326], line_41[324], line_40[322], line_39[320], line_38[318], line_37[316], line_36[314], line_35[312], line_34[310], line_33[308], line_32[306], line_31[304], line_30[302], line_29[300], line_28[298], line_27[296], line_26[294], line_25[292], line_24[290], line_23[288], line_22[286], line_21[284], line_20[282], line_19[280], line_18[278], line_17[276], line_16[274], line_15[272], line_14[270], line_13[268], line_12[266], line_11[264], line_10[262], line_9[260], line_8[258], line_7[256], line_6[254], line_5[252], line_4[250], line_3[248], line_2[246], line_1[244] };
assign col_499 = {line_128[499], line_127[497], line_126[495], line_125[493], line_124[491], line_123[489], line_122[487], line_121[485], line_120[483], line_119[481], line_118[479], line_117[477], line_116[475], line_115[473], line_114[471], line_113[469], line_112[467], line_111[465], line_110[463], line_109[461], line_108[459], line_107[457], line_106[455], line_105[453], line_104[451], line_103[449], line_102[447], line_101[445], line_100[443], line_99[441], line_98[439], line_97[437], line_96[435], line_95[433], line_94[431], line_93[429], line_92[427], line_91[425], line_90[423], line_89[421], line_88[419], line_87[417], line_86[415], line_85[413], line_84[411], line_83[409], line_82[407], line_81[405], line_80[403], line_79[401], line_78[399], line_77[397], line_76[395], line_75[393], line_74[391], line_73[389], line_72[387], line_71[385], line_70[383], line_69[381], line_68[379], line_67[377], line_66[375], line_65[373], line_64[371], line_63[369], line_62[367], line_61[365], line_60[363], line_59[361], line_58[359], line_57[357], line_56[355], line_55[353], line_54[351], line_53[349], line_52[347], line_51[345], line_50[343], line_49[341], line_48[339], line_47[337], line_46[335], line_45[333], line_44[331], line_43[329], line_42[327], line_41[325], line_40[323], line_39[321], line_38[319], line_37[317], line_36[315], line_35[313], line_34[311], line_33[309], line_32[307], line_31[305], line_30[303], line_29[301], line_28[299], line_27[297], line_26[295], line_25[293], line_24[291], line_23[289], line_22[287], line_21[285], line_20[283], line_19[281], line_18[279], line_17[277], line_16[275], line_15[273], line_14[271], line_13[269], line_12[267], line_11[265], line_10[263], line_9[261], line_8[259], line_7[257], line_6[255], line_5[253], line_4[251], line_3[249], line_2[247], line_1[245] };
assign col_500 = {line_128[500], line_127[498], line_126[496], line_125[494], line_124[492], line_123[490], line_122[488], line_121[486], line_120[484], line_119[482], line_118[480], line_117[478], line_116[476], line_115[474], line_114[472], line_113[470], line_112[468], line_111[466], line_110[464], line_109[462], line_108[460], line_107[458], line_106[456], line_105[454], line_104[452], line_103[450], line_102[448], line_101[446], line_100[444], line_99[442], line_98[440], line_97[438], line_96[436], line_95[434], line_94[432], line_93[430], line_92[428], line_91[426], line_90[424], line_89[422], line_88[420], line_87[418], line_86[416], line_85[414], line_84[412], line_83[410], line_82[408], line_81[406], line_80[404], line_79[402], line_78[400], line_77[398], line_76[396], line_75[394], line_74[392], line_73[390], line_72[388], line_71[386], line_70[384], line_69[382], line_68[380], line_67[378], line_66[376], line_65[374], line_64[372], line_63[370], line_62[368], line_61[366], line_60[364], line_59[362], line_58[360], line_57[358], line_56[356], line_55[354], line_54[352], line_53[350], line_52[348], line_51[346], line_50[344], line_49[342], line_48[340], line_47[338], line_46[336], line_45[334], line_44[332], line_43[330], line_42[328], line_41[326], line_40[324], line_39[322], line_38[320], line_37[318], line_36[316], line_35[314], line_34[312], line_33[310], line_32[308], line_31[306], line_30[304], line_29[302], line_28[300], line_27[298], line_26[296], line_25[294], line_24[292], line_23[290], line_22[288], line_21[286], line_20[284], line_19[282], line_18[280], line_17[278], line_16[276], line_15[274], line_14[272], line_13[270], line_12[268], line_11[266], line_10[264], line_9[262], line_8[260], line_7[258], line_6[256], line_5[254], line_4[252], line_3[250], line_2[248], line_1[246] };
assign col_501 = {line_128[501], line_127[499], line_126[497], line_125[495], line_124[493], line_123[491], line_122[489], line_121[487], line_120[485], line_119[483], line_118[481], line_117[479], line_116[477], line_115[475], line_114[473], line_113[471], line_112[469], line_111[467], line_110[465], line_109[463], line_108[461], line_107[459], line_106[457], line_105[455], line_104[453], line_103[451], line_102[449], line_101[447], line_100[445], line_99[443], line_98[441], line_97[439], line_96[437], line_95[435], line_94[433], line_93[431], line_92[429], line_91[427], line_90[425], line_89[423], line_88[421], line_87[419], line_86[417], line_85[415], line_84[413], line_83[411], line_82[409], line_81[407], line_80[405], line_79[403], line_78[401], line_77[399], line_76[397], line_75[395], line_74[393], line_73[391], line_72[389], line_71[387], line_70[385], line_69[383], line_68[381], line_67[379], line_66[377], line_65[375], line_64[373], line_63[371], line_62[369], line_61[367], line_60[365], line_59[363], line_58[361], line_57[359], line_56[357], line_55[355], line_54[353], line_53[351], line_52[349], line_51[347], line_50[345], line_49[343], line_48[341], line_47[339], line_46[337], line_45[335], line_44[333], line_43[331], line_42[329], line_41[327], line_40[325], line_39[323], line_38[321], line_37[319], line_36[317], line_35[315], line_34[313], line_33[311], line_32[309], line_31[307], line_30[305], line_29[303], line_28[301], line_27[299], line_26[297], line_25[295], line_24[293], line_23[291], line_22[289], line_21[287], line_20[285], line_19[283], line_18[281], line_17[279], line_16[277], line_15[275], line_14[273], line_13[271], line_12[269], line_11[267], line_10[265], line_9[263], line_8[261], line_7[259], line_6[257], line_5[255], line_4[253], line_3[251], line_2[249], line_1[247] };
assign col_502 = {line_128[502], line_127[500], line_126[498], line_125[496], line_124[494], line_123[492], line_122[490], line_121[488], line_120[486], line_119[484], line_118[482], line_117[480], line_116[478], line_115[476], line_114[474], line_113[472], line_112[470], line_111[468], line_110[466], line_109[464], line_108[462], line_107[460], line_106[458], line_105[456], line_104[454], line_103[452], line_102[450], line_101[448], line_100[446], line_99[444], line_98[442], line_97[440], line_96[438], line_95[436], line_94[434], line_93[432], line_92[430], line_91[428], line_90[426], line_89[424], line_88[422], line_87[420], line_86[418], line_85[416], line_84[414], line_83[412], line_82[410], line_81[408], line_80[406], line_79[404], line_78[402], line_77[400], line_76[398], line_75[396], line_74[394], line_73[392], line_72[390], line_71[388], line_70[386], line_69[384], line_68[382], line_67[380], line_66[378], line_65[376], line_64[374], line_63[372], line_62[370], line_61[368], line_60[366], line_59[364], line_58[362], line_57[360], line_56[358], line_55[356], line_54[354], line_53[352], line_52[350], line_51[348], line_50[346], line_49[344], line_48[342], line_47[340], line_46[338], line_45[336], line_44[334], line_43[332], line_42[330], line_41[328], line_40[326], line_39[324], line_38[322], line_37[320], line_36[318], line_35[316], line_34[314], line_33[312], line_32[310], line_31[308], line_30[306], line_29[304], line_28[302], line_27[300], line_26[298], line_25[296], line_24[294], line_23[292], line_22[290], line_21[288], line_20[286], line_19[284], line_18[282], line_17[280], line_16[278], line_15[276], line_14[274], line_13[272], line_12[270], line_11[268], line_10[266], line_9[264], line_8[262], line_7[260], line_6[258], line_5[256], line_4[254], line_3[252], line_2[250], line_1[248] };
assign col_503 = {line_128[503], line_127[501], line_126[499], line_125[497], line_124[495], line_123[493], line_122[491], line_121[489], line_120[487], line_119[485], line_118[483], line_117[481], line_116[479], line_115[477], line_114[475], line_113[473], line_112[471], line_111[469], line_110[467], line_109[465], line_108[463], line_107[461], line_106[459], line_105[457], line_104[455], line_103[453], line_102[451], line_101[449], line_100[447], line_99[445], line_98[443], line_97[441], line_96[439], line_95[437], line_94[435], line_93[433], line_92[431], line_91[429], line_90[427], line_89[425], line_88[423], line_87[421], line_86[419], line_85[417], line_84[415], line_83[413], line_82[411], line_81[409], line_80[407], line_79[405], line_78[403], line_77[401], line_76[399], line_75[397], line_74[395], line_73[393], line_72[391], line_71[389], line_70[387], line_69[385], line_68[383], line_67[381], line_66[379], line_65[377], line_64[375], line_63[373], line_62[371], line_61[369], line_60[367], line_59[365], line_58[363], line_57[361], line_56[359], line_55[357], line_54[355], line_53[353], line_52[351], line_51[349], line_50[347], line_49[345], line_48[343], line_47[341], line_46[339], line_45[337], line_44[335], line_43[333], line_42[331], line_41[329], line_40[327], line_39[325], line_38[323], line_37[321], line_36[319], line_35[317], line_34[315], line_33[313], line_32[311], line_31[309], line_30[307], line_29[305], line_28[303], line_27[301], line_26[299], line_25[297], line_24[295], line_23[293], line_22[291], line_21[289], line_20[287], line_19[285], line_18[283], line_17[281], line_16[279], line_15[277], line_14[275], line_13[273], line_12[271], line_11[269], line_10[267], line_9[265], line_8[263], line_7[261], line_6[259], line_5[257], line_4[255], line_3[253], line_2[251], line_1[249] };
assign col_504 = {line_128[504], line_127[502], line_126[500], line_125[498], line_124[496], line_123[494], line_122[492], line_121[490], line_120[488], line_119[486], line_118[484], line_117[482], line_116[480], line_115[478], line_114[476], line_113[474], line_112[472], line_111[470], line_110[468], line_109[466], line_108[464], line_107[462], line_106[460], line_105[458], line_104[456], line_103[454], line_102[452], line_101[450], line_100[448], line_99[446], line_98[444], line_97[442], line_96[440], line_95[438], line_94[436], line_93[434], line_92[432], line_91[430], line_90[428], line_89[426], line_88[424], line_87[422], line_86[420], line_85[418], line_84[416], line_83[414], line_82[412], line_81[410], line_80[408], line_79[406], line_78[404], line_77[402], line_76[400], line_75[398], line_74[396], line_73[394], line_72[392], line_71[390], line_70[388], line_69[386], line_68[384], line_67[382], line_66[380], line_65[378], line_64[376], line_63[374], line_62[372], line_61[370], line_60[368], line_59[366], line_58[364], line_57[362], line_56[360], line_55[358], line_54[356], line_53[354], line_52[352], line_51[350], line_50[348], line_49[346], line_48[344], line_47[342], line_46[340], line_45[338], line_44[336], line_43[334], line_42[332], line_41[330], line_40[328], line_39[326], line_38[324], line_37[322], line_36[320], line_35[318], line_34[316], line_33[314], line_32[312], line_31[310], line_30[308], line_29[306], line_28[304], line_27[302], line_26[300], line_25[298], line_24[296], line_23[294], line_22[292], line_21[290], line_20[288], line_19[286], line_18[284], line_17[282], line_16[280], line_15[278], line_14[276], line_13[274], line_12[272], line_11[270], line_10[268], line_9[266], line_8[264], line_7[262], line_6[260], line_5[258], line_4[256], line_3[254], line_2[252], line_1[250] };
assign col_505 = {line_128[505], line_127[503], line_126[501], line_125[499], line_124[497], line_123[495], line_122[493], line_121[491], line_120[489], line_119[487], line_118[485], line_117[483], line_116[481], line_115[479], line_114[477], line_113[475], line_112[473], line_111[471], line_110[469], line_109[467], line_108[465], line_107[463], line_106[461], line_105[459], line_104[457], line_103[455], line_102[453], line_101[451], line_100[449], line_99[447], line_98[445], line_97[443], line_96[441], line_95[439], line_94[437], line_93[435], line_92[433], line_91[431], line_90[429], line_89[427], line_88[425], line_87[423], line_86[421], line_85[419], line_84[417], line_83[415], line_82[413], line_81[411], line_80[409], line_79[407], line_78[405], line_77[403], line_76[401], line_75[399], line_74[397], line_73[395], line_72[393], line_71[391], line_70[389], line_69[387], line_68[385], line_67[383], line_66[381], line_65[379], line_64[377], line_63[375], line_62[373], line_61[371], line_60[369], line_59[367], line_58[365], line_57[363], line_56[361], line_55[359], line_54[357], line_53[355], line_52[353], line_51[351], line_50[349], line_49[347], line_48[345], line_47[343], line_46[341], line_45[339], line_44[337], line_43[335], line_42[333], line_41[331], line_40[329], line_39[327], line_38[325], line_37[323], line_36[321], line_35[319], line_34[317], line_33[315], line_32[313], line_31[311], line_30[309], line_29[307], line_28[305], line_27[303], line_26[301], line_25[299], line_24[297], line_23[295], line_22[293], line_21[291], line_20[289], line_19[287], line_18[285], line_17[283], line_16[281], line_15[279], line_14[277], line_13[275], line_12[273], line_11[271], line_10[269], line_9[267], line_8[265], line_7[263], line_6[261], line_5[259], line_4[257], line_3[255], line_2[253], line_1[251] };
assign col_506 = {line_128[506], line_127[504], line_126[502], line_125[500], line_124[498], line_123[496], line_122[494], line_121[492], line_120[490], line_119[488], line_118[486], line_117[484], line_116[482], line_115[480], line_114[478], line_113[476], line_112[474], line_111[472], line_110[470], line_109[468], line_108[466], line_107[464], line_106[462], line_105[460], line_104[458], line_103[456], line_102[454], line_101[452], line_100[450], line_99[448], line_98[446], line_97[444], line_96[442], line_95[440], line_94[438], line_93[436], line_92[434], line_91[432], line_90[430], line_89[428], line_88[426], line_87[424], line_86[422], line_85[420], line_84[418], line_83[416], line_82[414], line_81[412], line_80[410], line_79[408], line_78[406], line_77[404], line_76[402], line_75[400], line_74[398], line_73[396], line_72[394], line_71[392], line_70[390], line_69[388], line_68[386], line_67[384], line_66[382], line_65[380], line_64[378], line_63[376], line_62[374], line_61[372], line_60[370], line_59[368], line_58[366], line_57[364], line_56[362], line_55[360], line_54[358], line_53[356], line_52[354], line_51[352], line_50[350], line_49[348], line_48[346], line_47[344], line_46[342], line_45[340], line_44[338], line_43[336], line_42[334], line_41[332], line_40[330], line_39[328], line_38[326], line_37[324], line_36[322], line_35[320], line_34[318], line_33[316], line_32[314], line_31[312], line_30[310], line_29[308], line_28[306], line_27[304], line_26[302], line_25[300], line_24[298], line_23[296], line_22[294], line_21[292], line_20[290], line_19[288], line_18[286], line_17[284], line_16[282], line_15[280], line_14[278], line_13[276], line_12[274], line_11[272], line_10[270], line_9[268], line_8[266], line_7[264], line_6[262], line_5[260], line_4[258], line_3[256], line_2[254], line_1[252] };
assign col_507 = {line_128[507], line_127[505], line_126[503], line_125[501], line_124[499], line_123[497], line_122[495], line_121[493], line_120[491], line_119[489], line_118[487], line_117[485], line_116[483], line_115[481], line_114[479], line_113[477], line_112[475], line_111[473], line_110[471], line_109[469], line_108[467], line_107[465], line_106[463], line_105[461], line_104[459], line_103[457], line_102[455], line_101[453], line_100[451], line_99[449], line_98[447], line_97[445], line_96[443], line_95[441], line_94[439], line_93[437], line_92[435], line_91[433], line_90[431], line_89[429], line_88[427], line_87[425], line_86[423], line_85[421], line_84[419], line_83[417], line_82[415], line_81[413], line_80[411], line_79[409], line_78[407], line_77[405], line_76[403], line_75[401], line_74[399], line_73[397], line_72[395], line_71[393], line_70[391], line_69[389], line_68[387], line_67[385], line_66[383], line_65[381], line_64[379], line_63[377], line_62[375], line_61[373], line_60[371], line_59[369], line_58[367], line_57[365], line_56[363], line_55[361], line_54[359], line_53[357], line_52[355], line_51[353], line_50[351], line_49[349], line_48[347], line_47[345], line_46[343], line_45[341], line_44[339], line_43[337], line_42[335], line_41[333], line_40[331], line_39[329], line_38[327], line_37[325], line_36[323], line_35[321], line_34[319], line_33[317], line_32[315], line_31[313], line_30[311], line_29[309], line_28[307], line_27[305], line_26[303], line_25[301], line_24[299], line_23[297], line_22[295], line_21[293], line_20[291], line_19[289], line_18[287], line_17[285], line_16[283], line_15[281], line_14[279], line_13[277], line_12[275], line_11[273], line_10[271], line_9[269], line_8[267], line_7[265], line_6[263], line_5[261], line_4[259], line_3[257], line_2[255], line_1[253] };
assign col_508 = {line_128[508], line_127[506], line_126[504], line_125[502], line_124[500], line_123[498], line_122[496], line_121[494], line_120[492], line_119[490], line_118[488], line_117[486], line_116[484], line_115[482], line_114[480], line_113[478], line_112[476], line_111[474], line_110[472], line_109[470], line_108[468], line_107[466], line_106[464], line_105[462], line_104[460], line_103[458], line_102[456], line_101[454], line_100[452], line_99[450], line_98[448], line_97[446], line_96[444], line_95[442], line_94[440], line_93[438], line_92[436], line_91[434], line_90[432], line_89[430], line_88[428], line_87[426], line_86[424], line_85[422], line_84[420], line_83[418], line_82[416], line_81[414], line_80[412], line_79[410], line_78[408], line_77[406], line_76[404], line_75[402], line_74[400], line_73[398], line_72[396], line_71[394], line_70[392], line_69[390], line_68[388], line_67[386], line_66[384], line_65[382], line_64[380], line_63[378], line_62[376], line_61[374], line_60[372], line_59[370], line_58[368], line_57[366], line_56[364], line_55[362], line_54[360], line_53[358], line_52[356], line_51[354], line_50[352], line_49[350], line_48[348], line_47[346], line_46[344], line_45[342], line_44[340], line_43[338], line_42[336], line_41[334], line_40[332], line_39[330], line_38[328], line_37[326], line_36[324], line_35[322], line_34[320], line_33[318], line_32[316], line_31[314], line_30[312], line_29[310], line_28[308], line_27[306], line_26[304], line_25[302], line_24[300], line_23[298], line_22[296], line_21[294], line_20[292], line_19[290], line_18[288], line_17[286], line_16[284], line_15[282], line_14[280], line_13[278], line_12[276], line_11[274], line_10[272], line_9[270], line_8[268], line_7[266], line_6[264], line_5[262], line_4[260], line_3[258], line_2[256], line_1[254] };
assign col_509 = {line_128[509], line_127[507], line_126[505], line_125[503], line_124[501], line_123[499], line_122[497], line_121[495], line_120[493], line_119[491], line_118[489], line_117[487], line_116[485], line_115[483], line_114[481], line_113[479], line_112[477], line_111[475], line_110[473], line_109[471], line_108[469], line_107[467], line_106[465], line_105[463], line_104[461], line_103[459], line_102[457], line_101[455], line_100[453], line_99[451], line_98[449], line_97[447], line_96[445], line_95[443], line_94[441], line_93[439], line_92[437], line_91[435], line_90[433], line_89[431], line_88[429], line_87[427], line_86[425], line_85[423], line_84[421], line_83[419], line_82[417], line_81[415], line_80[413], line_79[411], line_78[409], line_77[407], line_76[405], line_75[403], line_74[401], line_73[399], line_72[397], line_71[395], line_70[393], line_69[391], line_68[389], line_67[387], line_66[385], line_65[383], line_64[381], line_63[379], line_62[377], line_61[375], line_60[373], line_59[371], line_58[369], line_57[367], line_56[365], line_55[363], line_54[361], line_53[359], line_52[357], line_51[355], line_50[353], line_49[351], line_48[349], line_47[347], line_46[345], line_45[343], line_44[341], line_43[339], line_42[337], line_41[335], line_40[333], line_39[331], line_38[329], line_37[327], line_36[325], line_35[323], line_34[321], line_33[319], line_32[317], line_31[315], line_30[313], line_29[311], line_28[309], line_27[307], line_26[305], line_25[303], line_24[301], line_23[299], line_22[297], line_21[295], line_20[293], line_19[291], line_18[289], line_17[287], line_16[285], line_15[283], line_14[281], line_13[279], line_12[277], line_11[275], line_10[273], line_9[271], line_8[269], line_7[267], line_6[265], line_5[263], line_4[261], line_3[259], line_2[257], line_1[255] };
assign col_510 = {line_128[510], line_127[508], line_126[506], line_125[504], line_124[502], line_123[500], line_122[498], line_121[496], line_120[494], line_119[492], line_118[490], line_117[488], line_116[486], line_115[484], line_114[482], line_113[480], line_112[478], line_111[476], line_110[474], line_109[472], line_108[470], line_107[468], line_106[466], line_105[464], line_104[462], line_103[460], line_102[458], line_101[456], line_100[454], line_99[452], line_98[450], line_97[448], line_96[446], line_95[444], line_94[442], line_93[440], line_92[438], line_91[436], line_90[434], line_89[432], line_88[430], line_87[428], line_86[426], line_85[424], line_84[422], line_83[420], line_82[418], line_81[416], line_80[414], line_79[412], line_78[410], line_77[408], line_76[406], line_75[404], line_74[402], line_73[400], line_72[398], line_71[396], line_70[394], line_69[392], line_68[390], line_67[388], line_66[386], line_65[384], line_64[382], line_63[380], line_62[378], line_61[376], line_60[374], line_59[372], line_58[370], line_57[368], line_56[366], line_55[364], line_54[362], line_53[360], line_52[358], line_51[356], line_50[354], line_49[352], line_48[350], line_47[348], line_46[346], line_45[344], line_44[342], line_43[340], line_42[338], line_41[336], line_40[334], line_39[332], line_38[330], line_37[328], line_36[326], line_35[324], line_34[322], line_33[320], line_32[318], line_31[316], line_30[314], line_29[312], line_28[310], line_27[308], line_26[306], line_25[304], line_24[302], line_23[300], line_22[298], line_21[296], line_20[294], line_19[292], line_18[290], line_17[288], line_16[286], line_15[284], line_14[282], line_13[280], line_12[278], line_11[276], line_10[274], line_9[272], line_8[270], line_7[268], line_6[266], line_5[264], line_4[262], line_3[260], line_2[258], line_1[256] };
assign col_511 = {line_128[511], line_127[509], line_126[507], line_125[505], line_124[503], line_123[501], line_122[499], line_121[497], line_120[495], line_119[493], line_118[491], line_117[489], line_116[487], line_115[485], line_114[483], line_113[481], line_112[479], line_111[477], line_110[475], line_109[473], line_108[471], line_107[469], line_106[467], line_105[465], line_104[463], line_103[461], line_102[459], line_101[457], line_100[455], line_99[453], line_98[451], line_97[449], line_96[447], line_95[445], line_94[443], line_93[441], line_92[439], line_91[437], line_90[435], line_89[433], line_88[431], line_87[429], line_86[427], line_85[425], line_84[423], line_83[421], line_82[419], line_81[417], line_80[415], line_79[413], line_78[411], line_77[409], line_76[407], line_75[405], line_74[403], line_73[401], line_72[399], line_71[397], line_70[395], line_69[393], line_68[391], line_67[389], line_66[387], line_65[385], line_64[383], line_63[381], line_62[379], line_61[377], line_60[375], line_59[373], line_58[371], line_57[369], line_56[367], line_55[365], line_54[363], line_53[361], line_52[359], line_51[357], line_50[355], line_49[353], line_48[351], line_47[349], line_46[347], line_45[345], line_44[343], line_43[341], line_42[339], line_41[337], line_40[335], line_39[333], line_38[331], line_37[329], line_36[327], line_35[325], line_34[323], line_33[321], line_32[319], line_31[317], line_30[315], line_29[313], line_28[311], line_27[309], line_26[307], line_25[305], line_24[303], line_23[301], line_22[299], line_21[297], line_20[295], line_19[293], line_18[291], line_17[289], line_16[287], line_15[285], line_14[283], line_13[281], line_12[279], line_11[277], line_10[275], line_9[273], line_8[271], line_7[269], line_6[267], line_5[265], line_4[263], line_3[261], line_2[259], line_1[257] };
assign col_512 = {line_128[512], line_127[510], line_126[508], line_125[506], line_124[504], line_123[502], line_122[500], line_121[498], line_120[496], line_119[494], line_118[492], line_117[490], line_116[488], line_115[486], line_114[484], line_113[482], line_112[480], line_111[478], line_110[476], line_109[474], line_108[472], line_107[470], line_106[468], line_105[466], line_104[464], line_103[462], line_102[460], line_101[458], line_100[456], line_99[454], line_98[452], line_97[450], line_96[448], line_95[446], line_94[444], line_93[442], line_92[440], line_91[438], line_90[436], line_89[434], line_88[432], line_87[430], line_86[428], line_85[426], line_84[424], line_83[422], line_82[420], line_81[418], line_80[416], line_79[414], line_78[412], line_77[410], line_76[408], line_75[406], line_74[404], line_73[402], line_72[400], line_71[398], line_70[396], line_69[394], line_68[392], line_67[390], line_66[388], line_65[386], line_64[384], line_63[382], line_62[380], line_61[378], line_60[376], line_59[374], line_58[372], line_57[370], line_56[368], line_55[366], line_54[364], line_53[362], line_52[360], line_51[358], line_50[356], line_49[354], line_48[352], line_47[350], line_46[348], line_45[346], line_44[344], line_43[342], line_42[340], line_41[338], line_40[336], line_39[334], line_38[332], line_37[330], line_36[328], line_35[326], line_34[324], line_33[322], line_32[320], line_31[318], line_30[316], line_29[314], line_28[312], line_27[310], line_26[308], line_25[306], line_24[304], line_23[302], line_22[300], line_21[298], line_20[296], line_19[294], line_18[292], line_17[290], line_16[288], line_15[286], line_14[284], line_13[282], line_12[280], line_11[278], line_10[276], line_9[274], line_8[272], line_7[270], line_6[268], line_5[266], line_4[264], line_3[262], line_2[260], line_1[258] };
assign col_513 = {line_128[513], line_127[511], line_126[509], line_125[507], line_124[505], line_123[503], line_122[501], line_121[499], line_120[497], line_119[495], line_118[493], line_117[491], line_116[489], line_115[487], line_114[485], line_113[483], line_112[481], line_111[479], line_110[477], line_109[475], line_108[473], line_107[471], line_106[469], line_105[467], line_104[465], line_103[463], line_102[461], line_101[459], line_100[457], line_99[455], line_98[453], line_97[451], line_96[449], line_95[447], line_94[445], line_93[443], line_92[441], line_91[439], line_90[437], line_89[435], line_88[433], line_87[431], line_86[429], line_85[427], line_84[425], line_83[423], line_82[421], line_81[419], line_80[417], line_79[415], line_78[413], line_77[411], line_76[409], line_75[407], line_74[405], line_73[403], line_72[401], line_71[399], line_70[397], line_69[395], line_68[393], line_67[391], line_66[389], line_65[387], line_64[385], line_63[383], line_62[381], line_61[379], line_60[377], line_59[375], line_58[373], line_57[371], line_56[369], line_55[367], line_54[365], line_53[363], line_52[361], line_51[359], line_50[357], line_49[355], line_48[353], line_47[351], line_46[349], line_45[347], line_44[345], line_43[343], line_42[341], line_41[339], line_40[337], line_39[335], line_38[333], line_37[331], line_36[329], line_35[327], line_34[325], line_33[323], line_32[321], line_31[319], line_30[317], line_29[315], line_28[313], line_27[311], line_26[309], line_25[307], line_24[305], line_23[303], line_22[301], line_21[299], line_20[297], line_19[295], line_18[293], line_17[291], line_16[289], line_15[287], line_14[285], line_13[283], line_12[281], line_11[279], line_10[277], line_9[275], line_8[273], line_7[271], line_6[269], line_5[267], line_4[265], line_3[263], line_2[261], line_1[259] };
assign col_514 = {line_128[514], line_127[512], line_126[510], line_125[508], line_124[506], line_123[504], line_122[502], line_121[500], line_120[498], line_119[496], line_118[494], line_117[492], line_116[490], line_115[488], line_114[486], line_113[484], line_112[482], line_111[480], line_110[478], line_109[476], line_108[474], line_107[472], line_106[470], line_105[468], line_104[466], line_103[464], line_102[462], line_101[460], line_100[458], line_99[456], line_98[454], line_97[452], line_96[450], line_95[448], line_94[446], line_93[444], line_92[442], line_91[440], line_90[438], line_89[436], line_88[434], line_87[432], line_86[430], line_85[428], line_84[426], line_83[424], line_82[422], line_81[420], line_80[418], line_79[416], line_78[414], line_77[412], line_76[410], line_75[408], line_74[406], line_73[404], line_72[402], line_71[400], line_70[398], line_69[396], line_68[394], line_67[392], line_66[390], line_65[388], line_64[386], line_63[384], line_62[382], line_61[380], line_60[378], line_59[376], line_58[374], line_57[372], line_56[370], line_55[368], line_54[366], line_53[364], line_52[362], line_51[360], line_50[358], line_49[356], line_48[354], line_47[352], line_46[350], line_45[348], line_44[346], line_43[344], line_42[342], line_41[340], line_40[338], line_39[336], line_38[334], line_37[332], line_36[330], line_35[328], line_34[326], line_33[324], line_32[322], line_31[320], line_30[318], line_29[316], line_28[314], line_27[312], line_26[310], line_25[308], line_24[306], line_23[304], line_22[302], line_21[300], line_20[298], line_19[296], line_18[294], line_17[292], line_16[290], line_15[288], line_14[286], line_13[284], line_12[282], line_11[280], line_10[278], line_9[276], line_8[274], line_7[272], line_6[270], line_5[268], line_4[266], line_3[264], line_2[262], line_1[260] };
assign col_515 = {line_128[515], line_127[513], line_126[511], line_125[509], line_124[507], line_123[505], line_122[503], line_121[501], line_120[499], line_119[497], line_118[495], line_117[493], line_116[491], line_115[489], line_114[487], line_113[485], line_112[483], line_111[481], line_110[479], line_109[477], line_108[475], line_107[473], line_106[471], line_105[469], line_104[467], line_103[465], line_102[463], line_101[461], line_100[459], line_99[457], line_98[455], line_97[453], line_96[451], line_95[449], line_94[447], line_93[445], line_92[443], line_91[441], line_90[439], line_89[437], line_88[435], line_87[433], line_86[431], line_85[429], line_84[427], line_83[425], line_82[423], line_81[421], line_80[419], line_79[417], line_78[415], line_77[413], line_76[411], line_75[409], line_74[407], line_73[405], line_72[403], line_71[401], line_70[399], line_69[397], line_68[395], line_67[393], line_66[391], line_65[389], line_64[387], line_63[385], line_62[383], line_61[381], line_60[379], line_59[377], line_58[375], line_57[373], line_56[371], line_55[369], line_54[367], line_53[365], line_52[363], line_51[361], line_50[359], line_49[357], line_48[355], line_47[353], line_46[351], line_45[349], line_44[347], line_43[345], line_42[343], line_41[341], line_40[339], line_39[337], line_38[335], line_37[333], line_36[331], line_35[329], line_34[327], line_33[325], line_32[323], line_31[321], line_30[319], line_29[317], line_28[315], line_27[313], line_26[311], line_25[309], line_24[307], line_23[305], line_22[303], line_21[301], line_20[299], line_19[297], line_18[295], line_17[293], line_16[291], line_15[289], line_14[287], line_13[285], line_12[283], line_11[281], line_10[279], line_9[277], line_8[275], line_7[273], line_6[271], line_5[269], line_4[267], line_3[265], line_2[263], line_1[261] };
assign col_516 = {line_128[516], line_127[514], line_126[512], line_125[510], line_124[508], line_123[506], line_122[504], line_121[502], line_120[500], line_119[498], line_118[496], line_117[494], line_116[492], line_115[490], line_114[488], line_113[486], line_112[484], line_111[482], line_110[480], line_109[478], line_108[476], line_107[474], line_106[472], line_105[470], line_104[468], line_103[466], line_102[464], line_101[462], line_100[460], line_99[458], line_98[456], line_97[454], line_96[452], line_95[450], line_94[448], line_93[446], line_92[444], line_91[442], line_90[440], line_89[438], line_88[436], line_87[434], line_86[432], line_85[430], line_84[428], line_83[426], line_82[424], line_81[422], line_80[420], line_79[418], line_78[416], line_77[414], line_76[412], line_75[410], line_74[408], line_73[406], line_72[404], line_71[402], line_70[400], line_69[398], line_68[396], line_67[394], line_66[392], line_65[390], line_64[388], line_63[386], line_62[384], line_61[382], line_60[380], line_59[378], line_58[376], line_57[374], line_56[372], line_55[370], line_54[368], line_53[366], line_52[364], line_51[362], line_50[360], line_49[358], line_48[356], line_47[354], line_46[352], line_45[350], line_44[348], line_43[346], line_42[344], line_41[342], line_40[340], line_39[338], line_38[336], line_37[334], line_36[332], line_35[330], line_34[328], line_33[326], line_32[324], line_31[322], line_30[320], line_29[318], line_28[316], line_27[314], line_26[312], line_25[310], line_24[308], line_23[306], line_22[304], line_21[302], line_20[300], line_19[298], line_18[296], line_17[294], line_16[292], line_15[290], line_14[288], line_13[286], line_12[284], line_11[282], line_10[280], line_9[278], line_8[276], line_7[274], line_6[272], line_5[270], line_4[268], line_3[266], line_2[264], line_1[262] };
assign col_517 = {line_128[517], line_127[515], line_126[513], line_125[511], line_124[509], line_123[507], line_122[505], line_121[503], line_120[501], line_119[499], line_118[497], line_117[495], line_116[493], line_115[491], line_114[489], line_113[487], line_112[485], line_111[483], line_110[481], line_109[479], line_108[477], line_107[475], line_106[473], line_105[471], line_104[469], line_103[467], line_102[465], line_101[463], line_100[461], line_99[459], line_98[457], line_97[455], line_96[453], line_95[451], line_94[449], line_93[447], line_92[445], line_91[443], line_90[441], line_89[439], line_88[437], line_87[435], line_86[433], line_85[431], line_84[429], line_83[427], line_82[425], line_81[423], line_80[421], line_79[419], line_78[417], line_77[415], line_76[413], line_75[411], line_74[409], line_73[407], line_72[405], line_71[403], line_70[401], line_69[399], line_68[397], line_67[395], line_66[393], line_65[391], line_64[389], line_63[387], line_62[385], line_61[383], line_60[381], line_59[379], line_58[377], line_57[375], line_56[373], line_55[371], line_54[369], line_53[367], line_52[365], line_51[363], line_50[361], line_49[359], line_48[357], line_47[355], line_46[353], line_45[351], line_44[349], line_43[347], line_42[345], line_41[343], line_40[341], line_39[339], line_38[337], line_37[335], line_36[333], line_35[331], line_34[329], line_33[327], line_32[325], line_31[323], line_30[321], line_29[319], line_28[317], line_27[315], line_26[313], line_25[311], line_24[309], line_23[307], line_22[305], line_21[303], line_20[301], line_19[299], line_18[297], line_17[295], line_16[293], line_15[291], line_14[289], line_13[287], line_12[285], line_11[283], line_10[281], line_9[279], line_8[277], line_7[275], line_6[273], line_5[271], line_4[269], line_3[267], line_2[265], line_1[263] };
assign col_518 = {line_128[518], line_127[516], line_126[514], line_125[512], line_124[510], line_123[508], line_122[506], line_121[504], line_120[502], line_119[500], line_118[498], line_117[496], line_116[494], line_115[492], line_114[490], line_113[488], line_112[486], line_111[484], line_110[482], line_109[480], line_108[478], line_107[476], line_106[474], line_105[472], line_104[470], line_103[468], line_102[466], line_101[464], line_100[462], line_99[460], line_98[458], line_97[456], line_96[454], line_95[452], line_94[450], line_93[448], line_92[446], line_91[444], line_90[442], line_89[440], line_88[438], line_87[436], line_86[434], line_85[432], line_84[430], line_83[428], line_82[426], line_81[424], line_80[422], line_79[420], line_78[418], line_77[416], line_76[414], line_75[412], line_74[410], line_73[408], line_72[406], line_71[404], line_70[402], line_69[400], line_68[398], line_67[396], line_66[394], line_65[392], line_64[390], line_63[388], line_62[386], line_61[384], line_60[382], line_59[380], line_58[378], line_57[376], line_56[374], line_55[372], line_54[370], line_53[368], line_52[366], line_51[364], line_50[362], line_49[360], line_48[358], line_47[356], line_46[354], line_45[352], line_44[350], line_43[348], line_42[346], line_41[344], line_40[342], line_39[340], line_38[338], line_37[336], line_36[334], line_35[332], line_34[330], line_33[328], line_32[326], line_31[324], line_30[322], line_29[320], line_28[318], line_27[316], line_26[314], line_25[312], line_24[310], line_23[308], line_22[306], line_21[304], line_20[302], line_19[300], line_18[298], line_17[296], line_16[294], line_15[292], line_14[290], line_13[288], line_12[286], line_11[284], line_10[282], line_9[280], line_8[278], line_7[276], line_6[274], line_5[272], line_4[270], line_3[268], line_2[266], line_1[264] };
assign col_519 = {line_128[519], line_127[517], line_126[515], line_125[513], line_124[511], line_123[509], line_122[507], line_121[505], line_120[503], line_119[501], line_118[499], line_117[497], line_116[495], line_115[493], line_114[491], line_113[489], line_112[487], line_111[485], line_110[483], line_109[481], line_108[479], line_107[477], line_106[475], line_105[473], line_104[471], line_103[469], line_102[467], line_101[465], line_100[463], line_99[461], line_98[459], line_97[457], line_96[455], line_95[453], line_94[451], line_93[449], line_92[447], line_91[445], line_90[443], line_89[441], line_88[439], line_87[437], line_86[435], line_85[433], line_84[431], line_83[429], line_82[427], line_81[425], line_80[423], line_79[421], line_78[419], line_77[417], line_76[415], line_75[413], line_74[411], line_73[409], line_72[407], line_71[405], line_70[403], line_69[401], line_68[399], line_67[397], line_66[395], line_65[393], line_64[391], line_63[389], line_62[387], line_61[385], line_60[383], line_59[381], line_58[379], line_57[377], line_56[375], line_55[373], line_54[371], line_53[369], line_52[367], line_51[365], line_50[363], line_49[361], line_48[359], line_47[357], line_46[355], line_45[353], line_44[351], line_43[349], line_42[347], line_41[345], line_40[343], line_39[341], line_38[339], line_37[337], line_36[335], line_35[333], line_34[331], line_33[329], line_32[327], line_31[325], line_30[323], line_29[321], line_28[319], line_27[317], line_26[315], line_25[313], line_24[311], line_23[309], line_22[307], line_21[305], line_20[303], line_19[301], line_18[299], line_17[297], line_16[295], line_15[293], line_14[291], line_13[289], line_12[287], line_11[285], line_10[283], line_9[281], line_8[279], line_7[277], line_6[275], line_5[273], line_4[271], line_3[269], line_2[267], line_1[265] };
assign col_520 = {line_128[520], line_127[518], line_126[516], line_125[514], line_124[512], line_123[510], line_122[508], line_121[506], line_120[504], line_119[502], line_118[500], line_117[498], line_116[496], line_115[494], line_114[492], line_113[490], line_112[488], line_111[486], line_110[484], line_109[482], line_108[480], line_107[478], line_106[476], line_105[474], line_104[472], line_103[470], line_102[468], line_101[466], line_100[464], line_99[462], line_98[460], line_97[458], line_96[456], line_95[454], line_94[452], line_93[450], line_92[448], line_91[446], line_90[444], line_89[442], line_88[440], line_87[438], line_86[436], line_85[434], line_84[432], line_83[430], line_82[428], line_81[426], line_80[424], line_79[422], line_78[420], line_77[418], line_76[416], line_75[414], line_74[412], line_73[410], line_72[408], line_71[406], line_70[404], line_69[402], line_68[400], line_67[398], line_66[396], line_65[394], line_64[392], line_63[390], line_62[388], line_61[386], line_60[384], line_59[382], line_58[380], line_57[378], line_56[376], line_55[374], line_54[372], line_53[370], line_52[368], line_51[366], line_50[364], line_49[362], line_48[360], line_47[358], line_46[356], line_45[354], line_44[352], line_43[350], line_42[348], line_41[346], line_40[344], line_39[342], line_38[340], line_37[338], line_36[336], line_35[334], line_34[332], line_33[330], line_32[328], line_31[326], line_30[324], line_29[322], line_28[320], line_27[318], line_26[316], line_25[314], line_24[312], line_23[310], line_22[308], line_21[306], line_20[304], line_19[302], line_18[300], line_17[298], line_16[296], line_15[294], line_14[292], line_13[290], line_12[288], line_11[286], line_10[284], line_9[282], line_8[280], line_7[278], line_6[276], line_5[274], line_4[272], line_3[270], line_2[268], line_1[266] };
assign col_521 = {line_128[521], line_127[519], line_126[517], line_125[515], line_124[513], line_123[511], line_122[509], line_121[507], line_120[505], line_119[503], line_118[501], line_117[499], line_116[497], line_115[495], line_114[493], line_113[491], line_112[489], line_111[487], line_110[485], line_109[483], line_108[481], line_107[479], line_106[477], line_105[475], line_104[473], line_103[471], line_102[469], line_101[467], line_100[465], line_99[463], line_98[461], line_97[459], line_96[457], line_95[455], line_94[453], line_93[451], line_92[449], line_91[447], line_90[445], line_89[443], line_88[441], line_87[439], line_86[437], line_85[435], line_84[433], line_83[431], line_82[429], line_81[427], line_80[425], line_79[423], line_78[421], line_77[419], line_76[417], line_75[415], line_74[413], line_73[411], line_72[409], line_71[407], line_70[405], line_69[403], line_68[401], line_67[399], line_66[397], line_65[395], line_64[393], line_63[391], line_62[389], line_61[387], line_60[385], line_59[383], line_58[381], line_57[379], line_56[377], line_55[375], line_54[373], line_53[371], line_52[369], line_51[367], line_50[365], line_49[363], line_48[361], line_47[359], line_46[357], line_45[355], line_44[353], line_43[351], line_42[349], line_41[347], line_40[345], line_39[343], line_38[341], line_37[339], line_36[337], line_35[335], line_34[333], line_33[331], line_32[329], line_31[327], line_30[325], line_29[323], line_28[321], line_27[319], line_26[317], line_25[315], line_24[313], line_23[311], line_22[309], line_21[307], line_20[305], line_19[303], line_18[301], line_17[299], line_16[297], line_15[295], line_14[293], line_13[291], line_12[289], line_11[287], line_10[285], line_9[283], line_8[281], line_7[279], line_6[277], line_5[275], line_4[273], line_3[271], line_2[269], line_1[267] };
assign col_522 = {line_128[522], line_127[520], line_126[518], line_125[516], line_124[514], line_123[512], line_122[510], line_121[508], line_120[506], line_119[504], line_118[502], line_117[500], line_116[498], line_115[496], line_114[494], line_113[492], line_112[490], line_111[488], line_110[486], line_109[484], line_108[482], line_107[480], line_106[478], line_105[476], line_104[474], line_103[472], line_102[470], line_101[468], line_100[466], line_99[464], line_98[462], line_97[460], line_96[458], line_95[456], line_94[454], line_93[452], line_92[450], line_91[448], line_90[446], line_89[444], line_88[442], line_87[440], line_86[438], line_85[436], line_84[434], line_83[432], line_82[430], line_81[428], line_80[426], line_79[424], line_78[422], line_77[420], line_76[418], line_75[416], line_74[414], line_73[412], line_72[410], line_71[408], line_70[406], line_69[404], line_68[402], line_67[400], line_66[398], line_65[396], line_64[394], line_63[392], line_62[390], line_61[388], line_60[386], line_59[384], line_58[382], line_57[380], line_56[378], line_55[376], line_54[374], line_53[372], line_52[370], line_51[368], line_50[366], line_49[364], line_48[362], line_47[360], line_46[358], line_45[356], line_44[354], line_43[352], line_42[350], line_41[348], line_40[346], line_39[344], line_38[342], line_37[340], line_36[338], line_35[336], line_34[334], line_33[332], line_32[330], line_31[328], line_30[326], line_29[324], line_28[322], line_27[320], line_26[318], line_25[316], line_24[314], line_23[312], line_22[310], line_21[308], line_20[306], line_19[304], line_18[302], line_17[300], line_16[298], line_15[296], line_14[294], line_13[292], line_12[290], line_11[288], line_10[286], line_9[284], line_8[282], line_7[280], line_6[278], line_5[276], line_4[274], line_3[272], line_2[270], line_1[268] };
assign col_523 = {line_128[523], line_127[521], line_126[519], line_125[517], line_124[515], line_123[513], line_122[511], line_121[509], line_120[507], line_119[505], line_118[503], line_117[501], line_116[499], line_115[497], line_114[495], line_113[493], line_112[491], line_111[489], line_110[487], line_109[485], line_108[483], line_107[481], line_106[479], line_105[477], line_104[475], line_103[473], line_102[471], line_101[469], line_100[467], line_99[465], line_98[463], line_97[461], line_96[459], line_95[457], line_94[455], line_93[453], line_92[451], line_91[449], line_90[447], line_89[445], line_88[443], line_87[441], line_86[439], line_85[437], line_84[435], line_83[433], line_82[431], line_81[429], line_80[427], line_79[425], line_78[423], line_77[421], line_76[419], line_75[417], line_74[415], line_73[413], line_72[411], line_71[409], line_70[407], line_69[405], line_68[403], line_67[401], line_66[399], line_65[397], line_64[395], line_63[393], line_62[391], line_61[389], line_60[387], line_59[385], line_58[383], line_57[381], line_56[379], line_55[377], line_54[375], line_53[373], line_52[371], line_51[369], line_50[367], line_49[365], line_48[363], line_47[361], line_46[359], line_45[357], line_44[355], line_43[353], line_42[351], line_41[349], line_40[347], line_39[345], line_38[343], line_37[341], line_36[339], line_35[337], line_34[335], line_33[333], line_32[331], line_31[329], line_30[327], line_29[325], line_28[323], line_27[321], line_26[319], line_25[317], line_24[315], line_23[313], line_22[311], line_21[309], line_20[307], line_19[305], line_18[303], line_17[301], line_16[299], line_15[297], line_14[295], line_13[293], line_12[291], line_11[289], line_10[287], line_9[285], line_8[283], line_7[281], line_6[279], line_5[277], line_4[275], line_3[273], line_2[271], line_1[269] };
assign col_524 = {line_128[524], line_127[522], line_126[520], line_125[518], line_124[516], line_123[514], line_122[512], line_121[510], line_120[508], line_119[506], line_118[504], line_117[502], line_116[500], line_115[498], line_114[496], line_113[494], line_112[492], line_111[490], line_110[488], line_109[486], line_108[484], line_107[482], line_106[480], line_105[478], line_104[476], line_103[474], line_102[472], line_101[470], line_100[468], line_99[466], line_98[464], line_97[462], line_96[460], line_95[458], line_94[456], line_93[454], line_92[452], line_91[450], line_90[448], line_89[446], line_88[444], line_87[442], line_86[440], line_85[438], line_84[436], line_83[434], line_82[432], line_81[430], line_80[428], line_79[426], line_78[424], line_77[422], line_76[420], line_75[418], line_74[416], line_73[414], line_72[412], line_71[410], line_70[408], line_69[406], line_68[404], line_67[402], line_66[400], line_65[398], line_64[396], line_63[394], line_62[392], line_61[390], line_60[388], line_59[386], line_58[384], line_57[382], line_56[380], line_55[378], line_54[376], line_53[374], line_52[372], line_51[370], line_50[368], line_49[366], line_48[364], line_47[362], line_46[360], line_45[358], line_44[356], line_43[354], line_42[352], line_41[350], line_40[348], line_39[346], line_38[344], line_37[342], line_36[340], line_35[338], line_34[336], line_33[334], line_32[332], line_31[330], line_30[328], line_29[326], line_28[324], line_27[322], line_26[320], line_25[318], line_24[316], line_23[314], line_22[312], line_21[310], line_20[308], line_19[306], line_18[304], line_17[302], line_16[300], line_15[298], line_14[296], line_13[294], line_12[292], line_11[290], line_10[288], line_9[286], line_8[284], line_7[282], line_6[280], line_5[278], line_4[276], line_3[274], line_2[272], line_1[270] };
assign col_525 = {line_128[525], line_127[523], line_126[521], line_125[519], line_124[517], line_123[515], line_122[513], line_121[511], line_120[509], line_119[507], line_118[505], line_117[503], line_116[501], line_115[499], line_114[497], line_113[495], line_112[493], line_111[491], line_110[489], line_109[487], line_108[485], line_107[483], line_106[481], line_105[479], line_104[477], line_103[475], line_102[473], line_101[471], line_100[469], line_99[467], line_98[465], line_97[463], line_96[461], line_95[459], line_94[457], line_93[455], line_92[453], line_91[451], line_90[449], line_89[447], line_88[445], line_87[443], line_86[441], line_85[439], line_84[437], line_83[435], line_82[433], line_81[431], line_80[429], line_79[427], line_78[425], line_77[423], line_76[421], line_75[419], line_74[417], line_73[415], line_72[413], line_71[411], line_70[409], line_69[407], line_68[405], line_67[403], line_66[401], line_65[399], line_64[397], line_63[395], line_62[393], line_61[391], line_60[389], line_59[387], line_58[385], line_57[383], line_56[381], line_55[379], line_54[377], line_53[375], line_52[373], line_51[371], line_50[369], line_49[367], line_48[365], line_47[363], line_46[361], line_45[359], line_44[357], line_43[355], line_42[353], line_41[351], line_40[349], line_39[347], line_38[345], line_37[343], line_36[341], line_35[339], line_34[337], line_33[335], line_32[333], line_31[331], line_30[329], line_29[327], line_28[325], line_27[323], line_26[321], line_25[319], line_24[317], line_23[315], line_22[313], line_21[311], line_20[309], line_19[307], line_18[305], line_17[303], line_16[301], line_15[299], line_14[297], line_13[295], line_12[293], line_11[291], line_10[289], line_9[287], line_8[285], line_7[283], line_6[281], line_5[279], line_4[277], line_3[275], line_2[273], line_1[271] };
assign col_526 = {line_128[526], line_127[524], line_126[522], line_125[520], line_124[518], line_123[516], line_122[514], line_121[512], line_120[510], line_119[508], line_118[506], line_117[504], line_116[502], line_115[500], line_114[498], line_113[496], line_112[494], line_111[492], line_110[490], line_109[488], line_108[486], line_107[484], line_106[482], line_105[480], line_104[478], line_103[476], line_102[474], line_101[472], line_100[470], line_99[468], line_98[466], line_97[464], line_96[462], line_95[460], line_94[458], line_93[456], line_92[454], line_91[452], line_90[450], line_89[448], line_88[446], line_87[444], line_86[442], line_85[440], line_84[438], line_83[436], line_82[434], line_81[432], line_80[430], line_79[428], line_78[426], line_77[424], line_76[422], line_75[420], line_74[418], line_73[416], line_72[414], line_71[412], line_70[410], line_69[408], line_68[406], line_67[404], line_66[402], line_65[400], line_64[398], line_63[396], line_62[394], line_61[392], line_60[390], line_59[388], line_58[386], line_57[384], line_56[382], line_55[380], line_54[378], line_53[376], line_52[374], line_51[372], line_50[370], line_49[368], line_48[366], line_47[364], line_46[362], line_45[360], line_44[358], line_43[356], line_42[354], line_41[352], line_40[350], line_39[348], line_38[346], line_37[344], line_36[342], line_35[340], line_34[338], line_33[336], line_32[334], line_31[332], line_30[330], line_29[328], line_28[326], line_27[324], line_26[322], line_25[320], line_24[318], line_23[316], line_22[314], line_21[312], line_20[310], line_19[308], line_18[306], line_17[304], line_16[302], line_15[300], line_14[298], line_13[296], line_12[294], line_11[292], line_10[290], line_9[288], line_8[286], line_7[284], line_6[282], line_5[280], line_4[278], line_3[276], line_2[274], line_1[272] };
assign col_527 = {line_128[527], line_127[525], line_126[523], line_125[521], line_124[519], line_123[517], line_122[515], line_121[513], line_120[511], line_119[509], line_118[507], line_117[505], line_116[503], line_115[501], line_114[499], line_113[497], line_112[495], line_111[493], line_110[491], line_109[489], line_108[487], line_107[485], line_106[483], line_105[481], line_104[479], line_103[477], line_102[475], line_101[473], line_100[471], line_99[469], line_98[467], line_97[465], line_96[463], line_95[461], line_94[459], line_93[457], line_92[455], line_91[453], line_90[451], line_89[449], line_88[447], line_87[445], line_86[443], line_85[441], line_84[439], line_83[437], line_82[435], line_81[433], line_80[431], line_79[429], line_78[427], line_77[425], line_76[423], line_75[421], line_74[419], line_73[417], line_72[415], line_71[413], line_70[411], line_69[409], line_68[407], line_67[405], line_66[403], line_65[401], line_64[399], line_63[397], line_62[395], line_61[393], line_60[391], line_59[389], line_58[387], line_57[385], line_56[383], line_55[381], line_54[379], line_53[377], line_52[375], line_51[373], line_50[371], line_49[369], line_48[367], line_47[365], line_46[363], line_45[361], line_44[359], line_43[357], line_42[355], line_41[353], line_40[351], line_39[349], line_38[347], line_37[345], line_36[343], line_35[341], line_34[339], line_33[337], line_32[335], line_31[333], line_30[331], line_29[329], line_28[327], line_27[325], line_26[323], line_25[321], line_24[319], line_23[317], line_22[315], line_21[313], line_20[311], line_19[309], line_18[307], line_17[305], line_16[303], line_15[301], line_14[299], line_13[297], line_12[295], line_11[293], line_10[291], line_9[289], line_8[287], line_7[285], line_6[283], line_5[281], line_4[279], line_3[277], line_2[275], line_1[273] };
assign col_528 = {line_128[528], line_127[526], line_126[524], line_125[522], line_124[520], line_123[518], line_122[516], line_121[514], line_120[512], line_119[510], line_118[508], line_117[506], line_116[504], line_115[502], line_114[500], line_113[498], line_112[496], line_111[494], line_110[492], line_109[490], line_108[488], line_107[486], line_106[484], line_105[482], line_104[480], line_103[478], line_102[476], line_101[474], line_100[472], line_99[470], line_98[468], line_97[466], line_96[464], line_95[462], line_94[460], line_93[458], line_92[456], line_91[454], line_90[452], line_89[450], line_88[448], line_87[446], line_86[444], line_85[442], line_84[440], line_83[438], line_82[436], line_81[434], line_80[432], line_79[430], line_78[428], line_77[426], line_76[424], line_75[422], line_74[420], line_73[418], line_72[416], line_71[414], line_70[412], line_69[410], line_68[408], line_67[406], line_66[404], line_65[402], line_64[400], line_63[398], line_62[396], line_61[394], line_60[392], line_59[390], line_58[388], line_57[386], line_56[384], line_55[382], line_54[380], line_53[378], line_52[376], line_51[374], line_50[372], line_49[370], line_48[368], line_47[366], line_46[364], line_45[362], line_44[360], line_43[358], line_42[356], line_41[354], line_40[352], line_39[350], line_38[348], line_37[346], line_36[344], line_35[342], line_34[340], line_33[338], line_32[336], line_31[334], line_30[332], line_29[330], line_28[328], line_27[326], line_26[324], line_25[322], line_24[320], line_23[318], line_22[316], line_21[314], line_20[312], line_19[310], line_18[308], line_17[306], line_16[304], line_15[302], line_14[300], line_13[298], line_12[296], line_11[294], line_10[292], line_9[290], line_8[288], line_7[286], line_6[284], line_5[282], line_4[280], line_3[278], line_2[276], line_1[274] };
assign col_529 = {line_128[529], line_127[527], line_126[525], line_125[523], line_124[521], line_123[519], line_122[517], line_121[515], line_120[513], line_119[511], line_118[509], line_117[507], line_116[505], line_115[503], line_114[501], line_113[499], line_112[497], line_111[495], line_110[493], line_109[491], line_108[489], line_107[487], line_106[485], line_105[483], line_104[481], line_103[479], line_102[477], line_101[475], line_100[473], line_99[471], line_98[469], line_97[467], line_96[465], line_95[463], line_94[461], line_93[459], line_92[457], line_91[455], line_90[453], line_89[451], line_88[449], line_87[447], line_86[445], line_85[443], line_84[441], line_83[439], line_82[437], line_81[435], line_80[433], line_79[431], line_78[429], line_77[427], line_76[425], line_75[423], line_74[421], line_73[419], line_72[417], line_71[415], line_70[413], line_69[411], line_68[409], line_67[407], line_66[405], line_65[403], line_64[401], line_63[399], line_62[397], line_61[395], line_60[393], line_59[391], line_58[389], line_57[387], line_56[385], line_55[383], line_54[381], line_53[379], line_52[377], line_51[375], line_50[373], line_49[371], line_48[369], line_47[367], line_46[365], line_45[363], line_44[361], line_43[359], line_42[357], line_41[355], line_40[353], line_39[351], line_38[349], line_37[347], line_36[345], line_35[343], line_34[341], line_33[339], line_32[337], line_31[335], line_30[333], line_29[331], line_28[329], line_27[327], line_26[325], line_25[323], line_24[321], line_23[319], line_22[317], line_21[315], line_20[313], line_19[311], line_18[309], line_17[307], line_16[305], line_15[303], line_14[301], line_13[299], line_12[297], line_11[295], line_10[293], line_9[291], line_8[289], line_7[287], line_6[285], line_5[283], line_4[281], line_3[279], line_2[277], line_1[275] };
assign col_530 = {line_128[530], line_127[528], line_126[526], line_125[524], line_124[522], line_123[520], line_122[518], line_121[516], line_120[514], line_119[512], line_118[510], line_117[508], line_116[506], line_115[504], line_114[502], line_113[500], line_112[498], line_111[496], line_110[494], line_109[492], line_108[490], line_107[488], line_106[486], line_105[484], line_104[482], line_103[480], line_102[478], line_101[476], line_100[474], line_99[472], line_98[470], line_97[468], line_96[466], line_95[464], line_94[462], line_93[460], line_92[458], line_91[456], line_90[454], line_89[452], line_88[450], line_87[448], line_86[446], line_85[444], line_84[442], line_83[440], line_82[438], line_81[436], line_80[434], line_79[432], line_78[430], line_77[428], line_76[426], line_75[424], line_74[422], line_73[420], line_72[418], line_71[416], line_70[414], line_69[412], line_68[410], line_67[408], line_66[406], line_65[404], line_64[402], line_63[400], line_62[398], line_61[396], line_60[394], line_59[392], line_58[390], line_57[388], line_56[386], line_55[384], line_54[382], line_53[380], line_52[378], line_51[376], line_50[374], line_49[372], line_48[370], line_47[368], line_46[366], line_45[364], line_44[362], line_43[360], line_42[358], line_41[356], line_40[354], line_39[352], line_38[350], line_37[348], line_36[346], line_35[344], line_34[342], line_33[340], line_32[338], line_31[336], line_30[334], line_29[332], line_28[330], line_27[328], line_26[326], line_25[324], line_24[322], line_23[320], line_22[318], line_21[316], line_20[314], line_19[312], line_18[310], line_17[308], line_16[306], line_15[304], line_14[302], line_13[300], line_12[298], line_11[296], line_10[294], line_9[292], line_8[290], line_7[288], line_6[286], line_5[284], line_4[282], line_3[280], line_2[278], line_1[276] };
assign col_531 = {line_128[531], line_127[529], line_126[527], line_125[525], line_124[523], line_123[521], line_122[519], line_121[517], line_120[515], line_119[513], line_118[511], line_117[509], line_116[507], line_115[505], line_114[503], line_113[501], line_112[499], line_111[497], line_110[495], line_109[493], line_108[491], line_107[489], line_106[487], line_105[485], line_104[483], line_103[481], line_102[479], line_101[477], line_100[475], line_99[473], line_98[471], line_97[469], line_96[467], line_95[465], line_94[463], line_93[461], line_92[459], line_91[457], line_90[455], line_89[453], line_88[451], line_87[449], line_86[447], line_85[445], line_84[443], line_83[441], line_82[439], line_81[437], line_80[435], line_79[433], line_78[431], line_77[429], line_76[427], line_75[425], line_74[423], line_73[421], line_72[419], line_71[417], line_70[415], line_69[413], line_68[411], line_67[409], line_66[407], line_65[405], line_64[403], line_63[401], line_62[399], line_61[397], line_60[395], line_59[393], line_58[391], line_57[389], line_56[387], line_55[385], line_54[383], line_53[381], line_52[379], line_51[377], line_50[375], line_49[373], line_48[371], line_47[369], line_46[367], line_45[365], line_44[363], line_43[361], line_42[359], line_41[357], line_40[355], line_39[353], line_38[351], line_37[349], line_36[347], line_35[345], line_34[343], line_33[341], line_32[339], line_31[337], line_30[335], line_29[333], line_28[331], line_27[329], line_26[327], line_25[325], line_24[323], line_23[321], line_22[319], line_21[317], line_20[315], line_19[313], line_18[311], line_17[309], line_16[307], line_15[305], line_14[303], line_13[301], line_12[299], line_11[297], line_10[295], line_9[293], line_8[291], line_7[289], line_6[287], line_5[285], line_4[283], line_3[281], line_2[279], line_1[277] };
assign col_532 = {line_128[532], line_127[530], line_126[528], line_125[526], line_124[524], line_123[522], line_122[520], line_121[518], line_120[516], line_119[514], line_118[512], line_117[510], line_116[508], line_115[506], line_114[504], line_113[502], line_112[500], line_111[498], line_110[496], line_109[494], line_108[492], line_107[490], line_106[488], line_105[486], line_104[484], line_103[482], line_102[480], line_101[478], line_100[476], line_99[474], line_98[472], line_97[470], line_96[468], line_95[466], line_94[464], line_93[462], line_92[460], line_91[458], line_90[456], line_89[454], line_88[452], line_87[450], line_86[448], line_85[446], line_84[444], line_83[442], line_82[440], line_81[438], line_80[436], line_79[434], line_78[432], line_77[430], line_76[428], line_75[426], line_74[424], line_73[422], line_72[420], line_71[418], line_70[416], line_69[414], line_68[412], line_67[410], line_66[408], line_65[406], line_64[404], line_63[402], line_62[400], line_61[398], line_60[396], line_59[394], line_58[392], line_57[390], line_56[388], line_55[386], line_54[384], line_53[382], line_52[380], line_51[378], line_50[376], line_49[374], line_48[372], line_47[370], line_46[368], line_45[366], line_44[364], line_43[362], line_42[360], line_41[358], line_40[356], line_39[354], line_38[352], line_37[350], line_36[348], line_35[346], line_34[344], line_33[342], line_32[340], line_31[338], line_30[336], line_29[334], line_28[332], line_27[330], line_26[328], line_25[326], line_24[324], line_23[322], line_22[320], line_21[318], line_20[316], line_19[314], line_18[312], line_17[310], line_16[308], line_15[306], line_14[304], line_13[302], line_12[300], line_11[298], line_10[296], line_9[294], line_8[292], line_7[290], line_6[288], line_5[286], line_4[284], line_3[282], line_2[280], line_1[278] };
assign col_533 = {line_128[533], line_127[531], line_126[529], line_125[527], line_124[525], line_123[523], line_122[521], line_121[519], line_120[517], line_119[515], line_118[513], line_117[511], line_116[509], line_115[507], line_114[505], line_113[503], line_112[501], line_111[499], line_110[497], line_109[495], line_108[493], line_107[491], line_106[489], line_105[487], line_104[485], line_103[483], line_102[481], line_101[479], line_100[477], line_99[475], line_98[473], line_97[471], line_96[469], line_95[467], line_94[465], line_93[463], line_92[461], line_91[459], line_90[457], line_89[455], line_88[453], line_87[451], line_86[449], line_85[447], line_84[445], line_83[443], line_82[441], line_81[439], line_80[437], line_79[435], line_78[433], line_77[431], line_76[429], line_75[427], line_74[425], line_73[423], line_72[421], line_71[419], line_70[417], line_69[415], line_68[413], line_67[411], line_66[409], line_65[407], line_64[405], line_63[403], line_62[401], line_61[399], line_60[397], line_59[395], line_58[393], line_57[391], line_56[389], line_55[387], line_54[385], line_53[383], line_52[381], line_51[379], line_50[377], line_49[375], line_48[373], line_47[371], line_46[369], line_45[367], line_44[365], line_43[363], line_42[361], line_41[359], line_40[357], line_39[355], line_38[353], line_37[351], line_36[349], line_35[347], line_34[345], line_33[343], line_32[341], line_31[339], line_30[337], line_29[335], line_28[333], line_27[331], line_26[329], line_25[327], line_24[325], line_23[323], line_22[321], line_21[319], line_20[317], line_19[315], line_18[313], line_17[311], line_16[309], line_15[307], line_14[305], line_13[303], line_12[301], line_11[299], line_10[297], line_9[295], line_8[293], line_7[291], line_6[289], line_5[287], line_4[285], line_3[283], line_2[281], line_1[279] };
assign col_534 = {line_128[534], line_127[532], line_126[530], line_125[528], line_124[526], line_123[524], line_122[522], line_121[520], line_120[518], line_119[516], line_118[514], line_117[512], line_116[510], line_115[508], line_114[506], line_113[504], line_112[502], line_111[500], line_110[498], line_109[496], line_108[494], line_107[492], line_106[490], line_105[488], line_104[486], line_103[484], line_102[482], line_101[480], line_100[478], line_99[476], line_98[474], line_97[472], line_96[470], line_95[468], line_94[466], line_93[464], line_92[462], line_91[460], line_90[458], line_89[456], line_88[454], line_87[452], line_86[450], line_85[448], line_84[446], line_83[444], line_82[442], line_81[440], line_80[438], line_79[436], line_78[434], line_77[432], line_76[430], line_75[428], line_74[426], line_73[424], line_72[422], line_71[420], line_70[418], line_69[416], line_68[414], line_67[412], line_66[410], line_65[408], line_64[406], line_63[404], line_62[402], line_61[400], line_60[398], line_59[396], line_58[394], line_57[392], line_56[390], line_55[388], line_54[386], line_53[384], line_52[382], line_51[380], line_50[378], line_49[376], line_48[374], line_47[372], line_46[370], line_45[368], line_44[366], line_43[364], line_42[362], line_41[360], line_40[358], line_39[356], line_38[354], line_37[352], line_36[350], line_35[348], line_34[346], line_33[344], line_32[342], line_31[340], line_30[338], line_29[336], line_28[334], line_27[332], line_26[330], line_25[328], line_24[326], line_23[324], line_22[322], line_21[320], line_20[318], line_19[316], line_18[314], line_17[312], line_16[310], line_15[308], line_14[306], line_13[304], line_12[302], line_11[300], line_10[298], line_9[296], line_8[294], line_7[292], line_6[290], line_5[288], line_4[286], line_3[284], line_2[282], line_1[280] };
assign col_535 = {line_128[535], line_127[533], line_126[531], line_125[529], line_124[527], line_123[525], line_122[523], line_121[521], line_120[519], line_119[517], line_118[515], line_117[513], line_116[511], line_115[509], line_114[507], line_113[505], line_112[503], line_111[501], line_110[499], line_109[497], line_108[495], line_107[493], line_106[491], line_105[489], line_104[487], line_103[485], line_102[483], line_101[481], line_100[479], line_99[477], line_98[475], line_97[473], line_96[471], line_95[469], line_94[467], line_93[465], line_92[463], line_91[461], line_90[459], line_89[457], line_88[455], line_87[453], line_86[451], line_85[449], line_84[447], line_83[445], line_82[443], line_81[441], line_80[439], line_79[437], line_78[435], line_77[433], line_76[431], line_75[429], line_74[427], line_73[425], line_72[423], line_71[421], line_70[419], line_69[417], line_68[415], line_67[413], line_66[411], line_65[409], line_64[407], line_63[405], line_62[403], line_61[401], line_60[399], line_59[397], line_58[395], line_57[393], line_56[391], line_55[389], line_54[387], line_53[385], line_52[383], line_51[381], line_50[379], line_49[377], line_48[375], line_47[373], line_46[371], line_45[369], line_44[367], line_43[365], line_42[363], line_41[361], line_40[359], line_39[357], line_38[355], line_37[353], line_36[351], line_35[349], line_34[347], line_33[345], line_32[343], line_31[341], line_30[339], line_29[337], line_28[335], line_27[333], line_26[331], line_25[329], line_24[327], line_23[325], line_22[323], line_21[321], line_20[319], line_19[317], line_18[315], line_17[313], line_16[311], line_15[309], line_14[307], line_13[305], line_12[303], line_11[301], line_10[299], line_9[297], line_8[295], line_7[293], line_6[291], line_5[289], line_4[287], line_3[285], line_2[283], line_1[281] };
assign col_536 = {line_128[536], line_127[534], line_126[532], line_125[530], line_124[528], line_123[526], line_122[524], line_121[522], line_120[520], line_119[518], line_118[516], line_117[514], line_116[512], line_115[510], line_114[508], line_113[506], line_112[504], line_111[502], line_110[500], line_109[498], line_108[496], line_107[494], line_106[492], line_105[490], line_104[488], line_103[486], line_102[484], line_101[482], line_100[480], line_99[478], line_98[476], line_97[474], line_96[472], line_95[470], line_94[468], line_93[466], line_92[464], line_91[462], line_90[460], line_89[458], line_88[456], line_87[454], line_86[452], line_85[450], line_84[448], line_83[446], line_82[444], line_81[442], line_80[440], line_79[438], line_78[436], line_77[434], line_76[432], line_75[430], line_74[428], line_73[426], line_72[424], line_71[422], line_70[420], line_69[418], line_68[416], line_67[414], line_66[412], line_65[410], line_64[408], line_63[406], line_62[404], line_61[402], line_60[400], line_59[398], line_58[396], line_57[394], line_56[392], line_55[390], line_54[388], line_53[386], line_52[384], line_51[382], line_50[380], line_49[378], line_48[376], line_47[374], line_46[372], line_45[370], line_44[368], line_43[366], line_42[364], line_41[362], line_40[360], line_39[358], line_38[356], line_37[354], line_36[352], line_35[350], line_34[348], line_33[346], line_32[344], line_31[342], line_30[340], line_29[338], line_28[336], line_27[334], line_26[332], line_25[330], line_24[328], line_23[326], line_22[324], line_21[322], line_20[320], line_19[318], line_18[316], line_17[314], line_16[312], line_15[310], line_14[308], line_13[306], line_12[304], line_11[302], line_10[300], line_9[298], line_8[296], line_7[294], line_6[292], line_5[290], line_4[288], line_3[286], line_2[284], line_1[282] };
assign col_537 = {line_128[537], line_127[535], line_126[533], line_125[531], line_124[529], line_123[527], line_122[525], line_121[523], line_120[521], line_119[519], line_118[517], line_117[515], line_116[513], line_115[511], line_114[509], line_113[507], line_112[505], line_111[503], line_110[501], line_109[499], line_108[497], line_107[495], line_106[493], line_105[491], line_104[489], line_103[487], line_102[485], line_101[483], line_100[481], line_99[479], line_98[477], line_97[475], line_96[473], line_95[471], line_94[469], line_93[467], line_92[465], line_91[463], line_90[461], line_89[459], line_88[457], line_87[455], line_86[453], line_85[451], line_84[449], line_83[447], line_82[445], line_81[443], line_80[441], line_79[439], line_78[437], line_77[435], line_76[433], line_75[431], line_74[429], line_73[427], line_72[425], line_71[423], line_70[421], line_69[419], line_68[417], line_67[415], line_66[413], line_65[411], line_64[409], line_63[407], line_62[405], line_61[403], line_60[401], line_59[399], line_58[397], line_57[395], line_56[393], line_55[391], line_54[389], line_53[387], line_52[385], line_51[383], line_50[381], line_49[379], line_48[377], line_47[375], line_46[373], line_45[371], line_44[369], line_43[367], line_42[365], line_41[363], line_40[361], line_39[359], line_38[357], line_37[355], line_36[353], line_35[351], line_34[349], line_33[347], line_32[345], line_31[343], line_30[341], line_29[339], line_28[337], line_27[335], line_26[333], line_25[331], line_24[329], line_23[327], line_22[325], line_21[323], line_20[321], line_19[319], line_18[317], line_17[315], line_16[313], line_15[311], line_14[309], line_13[307], line_12[305], line_11[303], line_10[301], line_9[299], line_8[297], line_7[295], line_6[293], line_5[291], line_4[289], line_3[287], line_2[285], line_1[283] };
assign col_538 = {line_128[538], line_127[536], line_126[534], line_125[532], line_124[530], line_123[528], line_122[526], line_121[524], line_120[522], line_119[520], line_118[518], line_117[516], line_116[514], line_115[512], line_114[510], line_113[508], line_112[506], line_111[504], line_110[502], line_109[500], line_108[498], line_107[496], line_106[494], line_105[492], line_104[490], line_103[488], line_102[486], line_101[484], line_100[482], line_99[480], line_98[478], line_97[476], line_96[474], line_95[472], line_94[470], line_93[468], line_92[466], line_91[464], line_90[462], line_89[460], line_88[458], line_87[456], line_86[454], line_85[452], line_84[450], line_83[448], line_82[446], line_81[444], line_80[442], line_79[440], line_78[438], line_77[436], line_76[434], line_75[432], line_74[430], line_73[428], line_72[426], line_71[424], line_70[422], line_69[420], line_68[418], line_67[416], line_66[414], line_65[412], line_64[410], line_63[408], line_62[406], line_61[404], line_60[402], line_59[400], line_58[398], line_57[396], line_56[394], line_55[392], line_54[390], line_53[388], line_52[386], line_51[384], line_50[382], line_49[380], line_48[378], line_47[376], line_46[374], line_45[372], line_44[370], line_43[368], line_42[366], line_41[364], line_40[362], line_39[360], line_38[358], line_37[356], line_36[354], line_35[352], line_34[350], line_33[348], line_32[346], line_31[344], line_30[342], line_29[340], line_28[338], line_27[336], line_26[334], line_25[332], line_24[330], line_23[328], line_22[326], line_21[324], line_20[322], line_19[320], line_18[318], line_17[316], line_16[314], line_15[312], line_14[310], line_13[308], line_12[306], line_11[304], line_10[302], line_9[300], line_8[298], line_7[296], line_6[294], line_5[292], line_4[290], line_3[288], line_2[286], line_1[284] };
assign col_539 = {line_128[539], line_127[537], line_126[535], line_125[533], line_124[531], line_123[529], line_122[527], line_121[525], line_120[523], line_119[521], line_118[519], line_117[517], line_116[515], line_115[513], line_114[511], line_113[509], line_112[507], line_111[505], line_110[503], line_109[501], line_108[499], line_107[497], line_106[495], line_105[493], line_104[491], line_103[489], line_102[487], line_101[485], line_100[483], line_99[481], line_98[479], line_97[477], line_96[475], line_95[473], line_94[471], line_93[469], line_92[467], line_91[465], line_90[463], line_89[461], line_88[459], line_87[457], line_86[455], line_85[453], line_84[451], line_83[449], line_82[447], line_81[445], line_80[443], line_79[441], line_78[439], line_77[437], line_76[435], line_75[433], line_74[431], line_73[429], line_72[427], line_71[425], line_70[423], line_69[421], line_68[419], line_67[417], line_66[415], line_65[413], line_64[411], line_63[409], line_62[407], line_61[405], line_60[403], line_59[401], line_58[399], line_57[397], line_56[395], line_55[393], line_54[391], line_53[389], line_52[387], line_51[385], line_50[383], line_49[381], line_48[379], line_47[377], line_46[375], line_45[373], line_44[371], line_43[369], line_42[367], line_41[365], line_40[363], line_39[361], line_38[359], line_37[357], line_36[355], line_35[353], line_34[351], line_33[349], line_32[347], line_31[345], line_30[343], line_29[341], line_28[339], line_27[337], line_26[335], line_25[333], line_24[331], line_23[329], line_22[327], line_21[325], line_20[323], line_19[321], line_18[319], line_17[317], line_16[315], line_15[313], line_14[311], line_13[309], line_12[307], line_11[305], line_10[303], line_9[301], line_8[299], line_7[297], line_6[295], line_5[293], line_4[291], line_3[289], line_2[287], line_1[285] };
assign col_540 = {line_128[540], line_127[538], line_126[536], line_125[534], line_124[532], line_123[530], line_122[528], line_121[526], line_120[524], line_119[522], line_118[520], line_117[518], line_116[516], line_115[514], line_114[512], line_113[510], line_112[508], line_111[506], line_110[504], line_109[502], line_108[500], line_107[498], line_106[496], line_105[494], line_104[492], line_103[490], line_102[488], line_101[486], line_100[484], line_99[482], line_98[480], line_97[478], line_96[476], line_95[474], line_94[472], line_93[470], line_92[468], line_91[466], line_90[464], line_89[462], line_88[460], line_87[458], line_86[456], line_85[454], line_84[452], line_83[450], line_82[448], line_81[446], line_80[444], line_79[442], line_78[440], line_77[438], line_76[436], line_75[434], line_74[432], line_73[430], line_72[428], line_71[426], line_70[424], line_69[422], line_68[420], line_67[418], line_66[416], line_65[414], line_64[412], line_63[410], line_62[408], line_61[406], line_60[404], line_59[402], line_58[400], line_57[398], line_56[396], line_55[394], line_54[392], line_53[390], line_52[388], line_51[386], line_50[384], line_49[382], line_48[380], line_47[378], line_46[376], line_45[374], line_44[372], line_43[370], line_42[368], line_41[366], line_40[364], line_39[362], line_38[360], line_37[358], line_36[356], line_35[354], line_34[352], line_33[350], line_32[348], line_31[346], line_30[344], line_29[342], line_28[340], line_27[338], line_26[336], line_25[334], line_24[332], line_23[330], line_22[328], line_21[326], line_20[324], line_19[322], line_18[320], line_17[318], line_16[316], line_15[314], line_14[312], line_13[310], line_12[308], line_11[306], line_10[304], line_9[302], line_8[300], line_7[298], line_6[296], line_5[294], line_4[292], line_3[290], line_2[288], line_1[286] };
assign col_541 = {line_128[541], line_127[539], line_126[537], line_125[535], line_124[533], line_123[531], line_122[529], line_121[527], line_120[525], line_119[523], line_118[521], line_117[519], line_116[517], line_115[515], line_114[513], line_113[511], line_112[509], line_111[507], line_110[505], line_109[503], line_108[501], line_107[499], line_106[497], line_105[495], line_104[493], line_103[491], line_102[489], line_101[487], line_100[485], line_99[483], line_98[481], line_97[479], line_96[477], line_95[475], line_94[473], line_93[471], line_92[469], line_91[467], line_90[465], line_89[463], line_88[461], line_87[459], line_86[457], line_85[455], line_84[453], line_83[451], line_82[449], line_81[447], line_80[445], line_79[443], line_78[441], line_77[439], line_76[437], line_75[435], line_74[433], line_73[431], line_72[429], line_71[427], line_70[425], line_69[423], line_68[421], line_67[419], line_66[417], line_65[415], line_64[413], line_63[411], line_62[409], line_61[407], line_60[405], line_59[403], line_58[401], line_57[399], line_56[397], line_55[395], line_54[393], line_53[391], line_52[389], line_51[387], line_50[385], line_49[383], line_48[381], line_47[379], line_46[377], line_45[375], line_44[373], line_43[371], line_42[369], line_41[367], line_40[365], line_39[363], line_38[361], line_37[359], line_36[357], line_35[355], line_34[353], line_33[351], line_32[349], line_31[347], line_30[345], line_29[343], line_28[341], line_27[339], line_26[337], line_25[335], line_24[333], line_23[331], line_22[329], line_21[327], line_20[325], line_19[323], line_18[321], line_17[319], line_16[317], line_15[315], line_14[313], line_13[311], line_12[309], line_11[307], line_10[305], line_9[303], line_8[301], line_7[299], line_6[297], line_5[295], line_4[293], line_3[291], line_2[289], line_1[287] };
assign col_542 = {line_128[542], line_127[540], line_126[538], line_125[536], line_124[534], line_123[532], line_122[530], line_121[528], line_120[526], line_119[524], line_118[522], line_117[520], line_116[518], line_115[516], line_114[514], line_113[512], line_112[510], line_111[508], line_110[506], line_109[504], line_108[502], line_107[500], line_106[498], line_105[496], line_104[494], line_103[492], line_102[490], line_101[488], line_100[486], line_99[484], line_98[482], line_97[480], line_96[478], line_95[476], line_94[474], line_93[472], line_92[470], line_91[468], line_90[466], line_89[464], line_88[462], line_87[460], line_86[458], line_85[456], line_84[454], line_83[452], line_82[450], line_81[448], line_80[446], line_79[444], line_78[442], line_77[440], line_76[438], line_75[436], line_74[434], line_73[432], line_72[430], line_71[428], line_70[426], line_69[424], line_68[422], line_67[420], line_66[418], line_65[416], line_64[414], line_63[412], line_62[410], line_61[408], line_60[406], line_59[404], line_58[402], line_57[400], line_56[398], line_55[396], line_54[394], line_53[392], line_52[390], line_51[388], line_50[386], line_49[384], line_48[382], line_47[380], line_46[378], line_45[376], line_44[374], line_43[372], line_42[370], line_41[368], line_40[366], line_39[364], line_38[362], line_37[360], line_36[358], line_35[356], line_34[354], line_33[352], line_32[350], line_31[348], line_30[346], line_29[344], line_28[342], line_27[340], line_26[338], line_25[336], line_24[334], line_23[332], line_22[330], line_21[328], line_20[326], line_19[324], line_18[322], line_17[320], line_16[318], line_15[316], line_14[314], line_13[312], line_12[310], line_11[308], line_10[306], line_9[304], line_8[302], line_7[300], line_6[298], line_5[296], line_4[294], line_3[292], line_2[290], line_1[288] };
assign col_543 = {line_128[543], line_127[541], line_126[539], line_125[537], line_124[535], line_123[533], line_122[531], line_121[529], line_120[527], line_119[525], line_118[523], line_117[521], line_116[519], line_115[517], line_114[515], line_113[513], line_112[511], line_111[509], line_110[507], line_109[505], line_108[503], line_107[501], line_106[499], line_105[497], line_104[495], line_103[493], line_102[491], line_101[489], line_100[487], line_99[485], line_98[483], line_97[481], line_96[479], line_95[477], line_94[475], line_93[473], line_92[471], line_91[469], line_90[467], line_89[465], line_88[463], line_87[461], line_86[459], line_85[457], line_84[455], line_83[453], line_82[451], line_81[449], line_80[447], line_79[445], line_78[443], line_77[441], line_76[439], line_75[437], line_74[435], line_73[433], line_72[431], line_71[429], line_70[427], line_69[425], line_68[423], line_67[421], line_66[419], line_65[417], line_64[415], line_63[413], line_62[411], line_61[409], line_60[407], line_59[405], line_58[403], line_57[401], line_56[399], line_55[397], line_54[395], line_53[393], line_52[391], line_51[389], line_50[387], line_49[385], line_48[383], line_47[381], line_46[379], line_45[377], line_44[375], line_43[373], line_42[371], line_41[369], line_40[367], line_39[365], line_38[363], line_37[361], line_36[359], line_35[357], line_34[355], line_33[353], line_32[351], line_31[349], line_30[347], line_29[345], line_28[343], line_27[341], line_26[339], line_25[337], line_24[335], line_23[333], line_22[331], line_21[329], line_20[327], line_19[325], line_18[323], line_17[321], line_16[319], line_15[317], line_14[315], line_13[313], line_12[311], line_11[309], line_10[307], line_9[305], line_8[303], line_7[301], line_6[299], line_5[297], line_4[295], line_3[293], line_2[291], line_1[289] };
assign col_544 = {line_128[544], line_127[542], line_126[540], line_125[538], line_124[536], line_123[534], line_122[532], line_121[530], line_120[528], line_119[526], line_118[524], line_117[522], line_116[520], line_115[518], line_114[516], line_113[514], line_112[512], line_111[510], line_110[508], line_109[506], line_108[504], line_107[502], line_106[500], line_105[498], line_104[496], line_103[494], line_102[492], line_101[490], line_100[488], line_99[486], line_98[484], line_97[482], line_96[480], line_95[478], line_94[476], line_93[474], line_92[472], line_91[470], line_90[468], line_89[466], line_88[464], line_87[462], line_86[460], line_85[458], line_84[456], line_83[454], line_82[452], line_81[450], line_80[448], line_79[446], line_78[444], line_77[442], line_76[440], line_75[438], line_74[436], line_73[434], line_72[432], line_71[430], line_70[428], line_69[426], line_68[424], line_67[422], line_66[420], line_65[418], line_64[416], line_63[414], line_62[412], line_61[410], line_60[408], line_59[406], line_58[404], line_57[402], line_56[400], line_55[398], line_54[396], line_53[394], line_52[392], line_51[390], line_50[388], line_49[386], line_48[384], line_47[382], line_46[380], line_45[378], line_44[376], line_43[374], line_42[372], line_41[370], line_40[368], line_39[366], line_38[364], line_37[362], line_36[360], line_35[358], line_34[356], line_33[354], line_32[352], line_31[350], line_30[348], line_29[346], line_28[344], line_27[342], line_26[340], line_25[338], line_24[336], line_23[334], line_22[332], line_21[330], line_20[328], line_19[326], line_18[324], line_17[322], line_16[320], line_15[318], line_14[316], line_13[314], line_12[312], line_11[310], line_10[308], line_9[306], line_8[304], line_7[302], line_6[300], line_5[298], line_4[296], line_3[294], line_2[292], line_1[290] };
assign col_545 = {line_128[545], line_127[543], line_126[541], line_125[539], line_124[537], line_123[535], line_122[533], line_121[531], line_120[529], line_119[527], line_118[525], line_117[523], line_116[521], line_115[519], line_114[517], line_113[515], line_112[513], line_111[511], line_110[509], line_109[507], line_108[505], line_107[503], line_106[501], line_105[499], line_104[497], line_103[495], line_102[493], line_101[491], line_100[489], line_99[487], line_98[485], line_97[483], line_96[481], line_95[479], line_94[477], line_93[475], line_92[473], line_91[471], line_90[469], line_89[467], line_88[465], line_87[463], line_86[461], line_85[459], line_84[457], line_83[455], line_82[453], line_81[451], line_80[449], line_79[447], line_78[445], line_77[443], line_76[441], line_75[439], line_74[437], line_73[435], line_72[433], line_71[431], line_70[429], line_69[427], line_68[425], line_67[423], line_66[421], line_65[419], line_64[417], line_63[415], line_62[413], line_61[411], line_60[409], line_59[407], line_58[405], line_57[403], line_56[401], line_55[399], line_54[397], line_53[395], line_52[393], line_51[391], line_50[389], line_49[387], line_48[385], line_47[383], line_46[381], line_45[379], line_44[377], line_43[375], line_42[373], line_41[371], line_40[369], line_39[367], line_38[365], line_37[363], line_36[361], line_35[359], line_34[357], line_33[355], line_32[353], line_31[351], line_30[349], line_29[347], line_28[345], line_27[343], line_26[341], line_25[339], line_24[337], line_23[335], line_22[333], line_21[331], line_20[329], line_19[327], line_18[325], line_17[323], line_16[321], line_15[319], line_14[317], line_13[315], line_12[313], line_11[311], line_10[309], line_9[307], line_8[305], line_7[303], line_6[301], line_5[299], line_4[297], line_3[295], line_2[293], line_1[291] };
assign col_546 = {line_128[546], line_127[544], line_126[542], line_125[540], line_124[538], line_123[536], line_122[534], line_121[532], line_120[530], line_119[528], line_118[526], line_117[524], line_116[522], line_115[520], line_114[518], line_113[516], line_112[514], line_111[512], line_110[510], line_109[508], line_108[506], line_107[504], line_106[502], line_105[500], line_104[498], line_103[496], line_102[494], line_101[492], line_100[490], line_99[488], line_98[486], line_97[484], line_96[482], line_95[480], line_94[478], line_93[476], line_92[474], line_91[472], line_90[470], line_89[468], line_88[466], line_87[464], line_86[462], line_85[460], line_84[458], line_83[456], line_82[454], line_81[452], line_80[450], line_79[448], line_78[446], line_77[444], line_76[442], line_75[440], line_74[438], line_73[436], line_72[434], line_71[432], line_70[430], line_69[428], line_68[426], line_67[424], line_66[422], line_65[420], line_64[418], line_63[416], line_62[414], line_61[412], line_60[410], line_59[408], line_58[406], line_57[404], line_56[402], line_55[400], line_54[398], line_53[396], line_52[394], line_51[392], line_50[390], line_49[388], line_48[386], line_47[384], line_46[382], line_45[380], line_44[378], line_43[376], line_42[374], line_41[372], line_40[370], line_39[368], line_38[366], line_37[364], line_36[362], line_35[360], line_34[358], line_33[356], line_32[354], line_31[352], line_30[350], line_29[348], line_28[346], line_27[344], line_26[342], line_25[340], line_24[338], line_23[336], line_22[334], line_21[332], line_20[330], line_19[328], line_18[326], line_17[324], line_16[322], line_15[320], line_14[318], line_13[316], line_12[314], line_11[312], line_10[310], line_9[308], line_8[306], line_7[304], line_6[302], line_5[300], line_4[298], line_3[296], line_2[294], line_1[292] };
assign col_547 = {line_128[547], line_127[545], line_126[543], line_125[541], line_124[539], line_123[537], line_122[535], line_121[533], line_120[531], line_119[529], line_118[527], line_117[525], line_116[523], line_115[521], line_114[519], line_113[517], line_112[515], line_111[513], line_110[511], line_109[509], line_108[507], line_107[505], line_106[503], line_105[501], line_104[499], line_103[497], line_102[495], line_101[493], line_100[491], line_99[489], line_98[487], line_97[485], line_96[483], line_95[481], line_94[479], line_93[477], line_92[475], line_91[473], line_90[471], line_89[469], line_88[467], line_87[465], line_86[463], line_85[461], line_84[459], line_83[457], line_82[455], line_81[453], line_80[451], line_79[449], line_78[447], line_77[445], line_76[443], line_75[441], line_74[439], line_73[437], line_72[435], line_71[433], line_70[431], line_69[429], line_68[427], line_67[425], line_66[423], line_65[421], line_64[419], line_63[417], line_62[415], line_61[413], line_60[411], line_59[409], line_58[407], line_57[405], line_56[403], line_55[401], line_54[399], line_53[397], line_52[395], line_51[393], line_50[391], line_49[389], line_48[387], line_47[385], line_46[383], line_45[381], line_44[379], line_43[377], line_42[375], line_41[373], line_40[371], line_39[369], line_38[367], line_37[365], line_36[363], line_35[361], line_34[359], line_33[357], line_32[355], line_31[353], line_30[351], line_29[349], line_28[347], line_27[345], line_26[343], line_25[341], line_24[339], line_23[337], line_22[335], line_21[333], line_20[331], line_19[329], line_18[327], line_17[325], line_16[323], line_15[321], line_14[319], line_13[317], line_12[315], line_11[313], line_10[311], line_9[309], line_8[307], line_7[305], line_6[303], line_5[301], line_4[299], line_3[297], line_2[295], line_1[293] };
assign col_548 = {line_128[548], line_127[546], line_126[544], line_125[542], line_124[540], line_123[538], line_122[536], line_121[534], line_120[532], line_119[530], line_118[528], line_117[526], line_116[524], line_115[522], line_114[520], line_113[518], line_112[516], line_111[514], line_110[512], line_109[510], line_108[508], line_107[506], line_106[504], line_105[502], line_104[500], line_103[498], line_102[496], line_101[494], line_100[492], line_99[490], line_98[488], line_97[486], line_96[484], line_95[482], line_94[480], line_93[478], line_92[476], line_91[474], line_90[472], line_89[470], line_88[468], line_87[466], line_86[464], line_85[462], line_84[460], line_83[458], line_82[456], line_81[454], line_80[452], line_79[450], line_78[448], line_77[446], line_76[444], line_75[442], line_74[440], line_73[438], line_72[436], line_71[434], line_70[432], line_69[430], line_68[428], line_67[426], line_66[424], line_65[422], line_64[420], line_63[418], line_62[416], line_61[414], line_60[412], line_59[410], line_58[408], line_57[406], line_56[404], line_55[402], line_54[400], line_53[398], line_52[396], line_51[394], line_50[392], line_49[390], line_48[388], line_47[386], line_46[384], line_45[382], line_44[380], line_43[378], line_42[376], line_41[374], line_40[372], line_39[370], line_38[368], line_37[366], line_36[364], line_35[362], line_34[360], line_33[358], line_32[356], line_31[354], line_30[352], line_29[350], line_28[348], line_27[346], line_26[344], line_25[342], line_24[340], line_23[338], line_22[336], line_21[334], line_20[332], line_19[330], line_18[328], line_17[326], line_16[324], line_15[322], line_14[320], line_13[318], line_12[316], line_11[314], line_10[312], line_9[310], line_8[308], line_7[306], line_6[304], line_5[302], line_4[300], line_3[298], line_2[296], line_1[294] };
assign col_549 = {line_128[549], line_127[547], line_126[545], line_125[543], line_124[541], line_123[539], line_122[537], line_121[535], line_120[533], line_119[531], line_118[529], line_117[527], line_116[525], line_115[523], line_114[521], line_113[519], line_112[517], line_111[515], line_110[513], line_109[511], line_108[509], line_107[507], line_106[505], line_105[503], line_104[501], line_103[499], line_102[497], line_101[495], line_100[493], line_99[491], line_98[489], line_97[487], line_96[485], line_95[483], line_94[481], line_93[479], line_92[477], line_91[475], line_90[473], line_89[471], line_88[469], line_87[467], line_86[465], line_85[463], line_84[461], line_83[459], line_82[457], line_81[455], line_80[453], line_79[451], line_78[449], line_77[447], line_76[445], line_75[443], line_74[441], line_73[439], line_72[437], line_71[435], line_70[433], line_69[431], line_68[429], line_67[427], line_66[425], line_65[423], line_64[421], line_63[419], line_62[417], line_61[415], line_60[413], line_59[411], line_58[409], line_57[407], line_56[405], line_55[403], line_54[401], line_53[399], line_52[397], line_51[395], line_50[393], line_49[391], line_48[389], line_47[387], line_46[385], line_45[383], line_44[381], line_43[379], line_42[377], line_41[375], line_40[373], line_39[371], line_38[369], line_37[367], line_36[365], line_35[363], line_34[361], line_33[359], line_32[357], line_31[355], line_30[353], line_29[351], line_28[349], line_27[347], line_26[345], line_25[343], line_24[341], line_23[339], line_22[337], line_21[335], line_20[333], line_19[331], line_18[329], line_17[327], line_16[325], line_15[323], line_14[321], line_13[319], line_12[317], line_11[315], line_10[313], line_9[311], line_8[309], line_7[307], line_6[305], line_5[303], line_4[301], line_3[299], line_2[297], line_1[295] };
assign col_550 = {line_128[550], line_127[548], line_126[546], line_125[544], line_124[542], line_123[540], line_122[538], line_121[536], line_120[534], line_119[532], line_118[530], line_117[528], line_116[526], line_115[524], line_114[522], line_113[520], line_112[518], line_111[516], line_110[514], line_109[512], line_108[510], line_107[508], line_106[506], line_105[504], line_104[502], line_103[500], line_102[498], line_101[496], line_100[494], line_99[492], line_98[490], line_97[488], line_96[486], line_95[484], line_94[482], line_93[480], line_92[478], line_91[476], line_90[474], line_89[472], line_88[470], line_87[468], line_86[466], line_85[464], line_84[462], line_83[460], line_82[458], line_81[456], line_80[454], line_79[452], line_78[450], line_77[448], line_76[446], line_75[444], line_74[442], line_73[440], line_72[438], line_71[436], line_70[434], line_69[432], line_68[430], line_67[428], line_66[426], line_65[424], line_64[422], line_63[420], line_62[418], line_61[416], line_60[414], line_59[412], line_58[410], line_57[408], line_56[406], line_55[404], line_54[402], line_53[400], line_52[398], line_51[396], line_50[394], line_49[392], line_48[390], line_47[388], line_46[386], line_45[384], line_44[382], line_43[380], line_42[378], line_41[376], line_40[374], line_39[372], line_38[370], line_37[368], line_36[366], line_35[364], line_34[362], line_33[360], line_32[358], line_31[356], line_30[354], line_29[352], line_28[350], line_27[348], line_26[346], line_25[344], line_24[342], line_23[340], line_22[338], line_21[336], line_20[334], line_19[332], line_18[330], line_17[328], line_16[326], line_15[324], line_14[322], line_13[320], line_12[318], line_11[316], line_10[314], line_9[312], line_8[310], line_7[308], line_6[306], line_5[304], line_4[302], line_3[300], line_2[298], line_1[296] };
assign col_551 = {line_128[551], line_127[549], line_126[547], line_125[545], line_124[543], line_123[541], line_122[539], line_121[537], line_120[535], line_119[533], line_118[531], line_117[529], line_116[527], line_115[525], line_114[523], line_113[521], line_112[519], line_111[517], line_110[515], line_109[513], line_108[511], line_107[509], line_106[507], line_105[505], line_104[503], line_103[501], line_102[499], line_101[497], line_100[495], line_99[493], line_98[491], line_97[489], line_96[487], line_95[485], line_94[483], line_93[481], line_92[479], line_91[477], line_90[475], line_89[473], line_88[471], line_87[469], line_86[467], line_85[465], line_84[463], line_83[461], line_82[459], line_81[457], line_80[455], line_79[453], line_78[451], line_77[449], line_76[447], line_75[445], line_74[443], line_73[441], line_72[439], line_71[437], line_70[435], line_69[433], line_68[431], line_67[429], line_66[427], line_65[425], line_64[423], line_63[421], line_62[419], line_61[417], line_60[415], line_59[413], line_58[411], line_57[409], line_56[407], line_55[405], line_54[403], line_53[401], line_52[399], line_51[397], line_50[395], line_49[393], line_48[391], line_47[389], line_46[387], line_45[385], line_44[383], line_43[381], line_42[379], line_41[377], line_40[375], line_39[373], line_38[371], line_37[369], line_36[367], line_35[365], line_34[363], line_33[361], line_32[359], line_31[357], line_30[355], line_29[353], line_28[351], line_27[349], line_26[347], line_25[345], line_24[343], line_23[341], line_22[339], line_21[337], line_20[335], line_19[333], line_18[331], line_17[329], line_16[327], line_15[325], line_14[323], line_13[321], line_12[319], line_11[317], line_10[315], line_9[313], line_8[311], line_7[309], line_6[307], line_5[305], line_4[303], line_3[301], line_2[299], line_1[297] };
assign col_552 = {line_128[552], line_127[550], line_126[548], line_125[546], line_124[544], line_123[542], line_122[540], line_121[538], line_120[536], line_119[534], line_118[532], line_117[530], line_116[528], line_115[526], line_114[524], line_113[522], line_112[520], line_111[518], line_110[516], line_109[514], line_108[512], line_107[510], line_106[508], line_105[506], line_104[504], line_103[502], line_102[500], line_101[498], line_100[496], line_99[494], line_98[492], line_97[490], line_96[488], line_95[486], line_94[484], line_93[482], line_92[480], line_91[478], line_90[476], line_89[474], line_88[472], line_87[470], line_86[468], line_85[466], line_84[464], line_83[462], line_82[460], line_81[458], line_80[456], line_79[454], line_78[452], line_77[450], line_76[448], line_75[446], line_74[444], line_73[442], line_72[440], line_71[438], line_70[436], line_69[434], line_68[432], line_67[430], line_66[428], line_65[426], line_64[424], line_63[422], line_62[420], line_61[418], line_60[416], line_59[414], line_58[412], line_57[410], line_56[408], line_55[406], line_54[404], line_53[402], line_52[400], line_51[398], line_50[396], line_49[394], line_48[392], line_47[390], line_46[388], line_45[386], line_44[384], line_43[382], line_42[380], line_41[378], line_40[376], line_39[374], line_38[372], line_37[370], line_36[368], line_35[366], line_34[364], line_33[362], line_32[360], line_31[358], line_30[356], line_29[354], line_28[352], line_27[350], line_26[348], line_25[346], line_24[344], line_23[342], line_22[340], line_21[338], line_20[336], line_19[334], line_18[332], line_17[330], line_16[328], line_15[326], line_14[324], line_13[322], line_12[320], line_11[318], line_10[316], line_9[314], line_8[312], line_7[310], line_6[308], line_5[306], line_4[304], line_3[302], line_2[300], line_1[298] };
assign col_553 = {line_128[553], line_127[551], line_126[549], line_125[547], line_124[545], line_123[543], line_122[541], line_121[539], line_120[537], line_119[535], line_118[533], line_117[531], line_116[529], line_115[527], line_114[525], line_113[523], line_112[521], line_111[519], line_110[517], line_109[515], line_108[513], line_107[511], line_106[509], line_105[507], line_104[505], line_103[503], line_102[501], line_101[499], line_100[497], line_99[495], line_98[493], line_97[491], line_96[489], line_95[487], line_94[485], line_93[483], line_92[481], line_91[479], line_90[477], line_89[475], line_88[473], line_87[471], line_86[469], line_85[467], line_84[465], line_83[463], line_82[461], line_81[459], line_80[457], line_79[455], line_78[453], line_77[451], line_76[449], line_75[447], line_74[445], line_73[443], line_72[441], line_71[439], line_70[437], line_69[435], line_68[433], line_67[431], line_66[429], line_65[427], line_64[425], line_63[423], line_62[421], line_61[419], line_60[417], line_59[415], line_58[413], line_57[411], line_56[409], line_55[407], line_54[405], line_53[403], line_52[401], line_51[399], line_50[397], line_49[395], line_48[393], line_47[391], line_46[389], line_45[387], line_44[385], line_43[383], line_42[381], line_41[379], line_40[377], line_39[375], line_38[373], line_37[371], line_36[369], line_35[367], line_34[365], line_33[363], line_32[361], line_31[359], line_30[357], line_29[355], line_28[353], line_27[351], line_26[349], line_25[347], line_24[345], line_23[343], line_22[341], line_21[339], line_20[337], line_19[335], line_18[333], line_17[331], line_16[329], line_15[327], line_14[325], line_13[323], line_12[321], line_11[319], line_10[317], line_9[315], line_8[313], line_7[311], line_6[309], line_5[307], line_4[305], line_3[303], line_2[301], line_1[299] };
assign col_554 = {line_128[554], line_127[552], line_126[550], line_125[548], line_124[546], line_123[544], line_122[542], line_121[540], line_120[538], line_119[536], line_118[534], line_117[532], line_116[530], line_115[528], line_114[526], line_113[524], line_112[522], line_111[520], line_110[518], line_109[516], line_108[514], line_107[512], line_106[510], line_105[508], line_104[506], line_103[504], line_102[502], line_101[500], line_100[498], line_99[496], line_98[494], line_97[492], line_96[490], line_95[488], line_94[486], line_93[484], line_92[482], line_91[480], line_90[478], line_89[476], line_88[474], line_87[472], line_86[470], line_85[468], line_84[466], line_83[464], line_82[462], line_81[460], line_80[458], line_79[456], line_78[454], line_77[452], line_76[450], line_75[448], line_74[446], line_73[444], line_72[442], line_71[440], line_70[438], line_69[436], line_68[434], line_67[432], line_66[430], line_65[428], line_64[426], line_63[424], line_62[422], line_61[420], line_60[418], line_59[416], line_58[414], line_57[412], line_56[410], line_55[408], line_54[406], line_53[404], line_52[402], line_51[400], line_50[398], line_49[396], line_48[394], line_47[392], line_46[390], line_45[388], line_44[386], line_43[384], line_42[382], line_41[380], line_40[378], line_39[376], line_38[374], line_37[372], line_36[370], line_35[368], line_34[366], line_33[364], line_32[362], line_31[360], line_30[358], line_29[356], line_28[354], line_27[352], line_26[350], line_25[348], line_24[346], line_23[344], line_22[342], line_21[340], line_20[338], line_19[336], line_18[334], line_17[332], line_16[330], line_15[328], line_14[326], line_13[324], line_12[322], line_11[320], line_10[318], line_9[316], line_8[314], line_7[312], line_6[310], line_5[308], line_4[306], line_3[304], line_2[302], line_1[300] };
assign col_555 = {line_128[555], line_127[553], line_126[551], line_125[549], line_124[547], line_123[545], line_122[543], line_121[541], line_120[539], line_119[537], line_118[535], line_117[533], line_116[531], line_115[529], line_114[527], line_113[525], line_112[523], line_111[521], line_110[519], line_109[517], line_108[515], line_107[513], line_106[511], line_105[509], line_104[507], line_103[505], line_102[503], line_101[501], line_100[499], line_99[497], line_98[495], line_97[493], line_96[491], line_95[489], line_94[487], line_93[485], line_92[483], line_91[481], line_90[479], line_89[477], line_88[475], line_87[473], line_86[471], line_85[469], line_84[467], line_83[465], line_82[463], line_81[461], line_80[459], line_79[457], line_78[455], line_77[453], line_76[451], line_75[449], line_74[447], line_73[445], line_72[443], line_71[441], line_70[439], line_69[437], line_68[435], line_67[433], line_66[431], line_65[429], line_64[427], line_63[425], line_62[423], line_61[421], line_60[419], line_59[417], line_58[415], line_57[413], line_56[411], line_55[409], line_54[407], line_53[405], line_52[403], line_51[401], line_50[399], line_49[397], line_48[395], line_47[393], line_46[391], line_45[389], line_44[387], line_43[385], line_42[383], line_41[381], line_40[379], line_39[377], line_38[375], line_37[373], line_36[371], line_35[369], line_34[367], line_33[365], line_32[363], line_31[361], line_30[359], line_29[357], line_28[355], line_27[353], line_26[351], line_25[349], line_24[347], line_23[345], line_22[343], line_21[341], line_20[339], line_19[337], line_18[335], line_17[333], line_16[331], line_15[329], line_14[327], line_13[325], line_12[323], line_11[321], line_10[319], line_9[317], line_8[315], line_7[313], line_6[311], line_5[309], line_4[307], line_3[305], line_2[303], line_1[301] };
assign col_556 = {line_128[556], line_127[554], line_126[552], line_125[550], line_124[548], line_123[546], line_122[544], line_121[542], line_120[540], line_119[538], line_118[536], line_117[534], line_116[532], line_115[530], line_114[528], line_113[526], line_112[524], line_111[522], line_110[520], line_109[518], line_108[516], line_107[514], line_106[512], line_105[510], line_104[508], line_103[506], line_102[504], line_101[502], line_100[500], line_99[498], line_98[496], line_97[494], line_96[492], line_95[490], line_94[488], line_93[486], line_92[484], line_91[482], line_90[480], line_89[478], line_88[476], line_87[474], line_86[472], line_85[470], line_84[468], line_83[466], line_82[464], line_81[462], line_80[460], line_79[458], line_78[456], line_77[454], line_76[452], line_75[450], line_74[448], line_73[446], line_72[444], line_71[442], line_70[440], line_69[438], line_68[436], line_67[434], line_66[432], line_65[430], line_64[428], line_63[426], line_62[424], line_61[422], line_60[420], line_59[418], line_58[416], line_57[414], line_56[412], line_55[410], line_54[408], line_53[406], line_52[404], line_51[402], line_50[400], line_49[398], line_48[396], line_47[394], line_46[392], line_45[390], line_44[388], line_43[386], line_42[384], line_41[382], line_40[380], line_39[378], line_38[376], line_37[374], line_36[372], line_35[370], line_34[368], line_33[366], line_32[364], line_31[362], line_30[360], line_29[358], line_28[356], line_27[354], line_26[352], line_25[350], line_24[348], line_23[346], line_22[344], line_21[342], line_20[340], line_19[338], line_18[336], line_17[334], line_16[332], line_15[330], line_14[328], line_13[326], line_12[324], line_11[322], line_10[320], line_9[318], line_8[316], line_7[314], line_6[312], line_5[310], line_4[308], line_3[306], line_2[304], line_1[302] };
assign col_557 = {line_128[557], line_127[555], line_126[553], line_125[551], line_124[549], line_123[547], line_122[545], line_121[543], line_120[541], line_119[539], line_118[537], line_117[535], line_116[533], line_115[531], line_114[529], line_113[527], line_112[525], line_111[523], line_110[521], line_109[519], line_108[517], line_107[515], line_106[513], line_105[511], line_104[509], line_103[507], line_102[505], line_101[503], line_100[501], line_99[499], line_98[497], line_97[495], line_96[493], line_95[491], line_94[489], line_93[487], line_92[485], line_91[483], line_90[481], line_89[479], line_88[477], line_87[475], line_86[473], line_85[471], line_84[469], line_83[467], line_82[465], line_81[463], line_80[461], line_79[459], line_78[457], line_77[455], line_76[453], line_75[451], line_74[449], line_73[447], line_72[445], line_71[443], line_70[441], line_69[439], line_68[437], line_67[435], line_66[433], line_65[431], line_64[429], line_63[427], line_62[425], line_61[423], line_60[421], line_59[419], line_58[417], line_57[415], line_56[413], line_55[411], line_54[409], line_53[407], line_52[405], line_51[403], line_50[401], line_49[399], line_48[397], line_47[395], line_46[393], line_45[391], line_44[389], line_43[387], line_42[385], line_41[383], line_40[381], line_39[379], line_38[377], line_37[375], line_36[373], line_35[371], line_34[369], line_33[367], line_32[365], line_31[363], line_30[361], line_29[359], line_28[357], line_27[355], line_26[353], line_25[351], line_24[349], line_23[347], line_22[345], line_21[343], line_20[341], line_19[339], line_18[337], line_17[335], line_16[333], line_15[331], line_14[329], line_13[327], line_12[325], line_11[323], line_10[321], line_9[319], line_8[317], line_7[315], line_6[313], line_5[311], line_4[309], line_3[307], line_2[305], line_1[303] };
assign col_558 = {line_128[558], line_127[556], line_126[554], line_125[552], line_124[550], line_123[548], line_122[546], line_121[544], line_120[542], line_119[540], line_118[538], line_117[536], line_116[534], line_115[532], line_114[530], line_113[528], line_112[526], line_111[524], line_110[522], line_109[520], line_108[518], line_107[516], line_106[514], line_105[512], line_104[510], line_103[508], line_102[506], line_101[504], line_100[502], line_99[500], line_98[498], line_97[496], line_96[494], line_95[492], line_94[490], line_93[488], line_92[486], line_91[484], line_90[482], line_89[480], line_88[478], line_87[476], line_86[474], line_85[472], line_84[470], line_83[468], line_82[466], line_81[464], line_80[462], line_79[460], line_78[458], line_77[456], line_76[454], line_75[452], line_74[450], line_73[448], line_72[446], line_71[444], line_70[442], line_69[440], line_68[438], line_67[436], line_66[434], line_65[432], line_64[430], line_63[428], line_62[426], line_61[424], line_60[422], line_59[420], line_58[418], line_57[416], line_56[414], line_55[412], line_54[410], line_53[408], line_52[406], line_51[404], line_50[402], line_49[400], line_48[398], line_47[396], line_46[394], line_45[392], line_44[390], line_43[388], line_42[386], line_41[384], line_40[382], line_39[380], line_38[378], line_37[376], line_36[374], line_35[372], line_34[370], line_33[368], line_32[366], line_31[364], line_30[362], line_29[360], line_28[358], line_27[356], line_26[354], line_25[352], line_24[350], line_23[348], line_22[346], line_21[344], line_20[342], line_19[340], line_18[338], line_17[336], line_16[334], line_15[332], line_14[330], line_13[328], line_12[326], line_11[324], line_10[322], line_9[320], line_8[318], line_7[316], line_6[314], line_5[312], line_4[310], line_3[308], line_2[306], line_1[304] };
assign col_559 = {line_128[559], line_127[557], line_126[555], line_125[553], line_124[551], line_123[549], line_122[547], line_121[545], line_120[543], line_119[541], line_118[539], line_117[537], line_116[535], line_115[533], line_114[531], line_113[529], line_112[527], line_111[525], line_110[523], line_109[521], line_108[519], line_107[517], line_106[515], line_105[513], line_104[511], line_103[509], line_102[507], line_101[505], line_100[503], line_99[501], line_98[499], line_97[497], line_96[495], line_95[493], line_94[491], line_93[489], line_92[487], line_91[485], line_90[483], line_89[481], line_88[479], line_87[477], line_86[475], line_85[473], line_84[471], line_83[469], line_82[467], line_81[465], line_80[463], line_79[461], line_78[459], line_77[457], line_76[455], line_75[453], line_74[451], line_73[449], line_72[447], line_71[445], line_70[443], line_69[441], line_68[439], line_67[437], line_66[435], line_65[433], line_64[431], line_63[429], line_62[427], line_61[425], line_60[423], line_59[421], line_58[419], line_57[417], line_56[415], line_55[413], line_54[411], line_53[409], line_52[407], line_51[405], line_50[403], line_49[401], line_48[399], line_47[397], line_46[395], line_45[393], line_44[391], line_43[389], line_42[387], line_41[385], line_40[383], line_39[381], line_38[379], line_37[377], line_36[375], line_35[373], line_34[371], line_33[369], line_32[367], line_31[365], line_30[363], line_29[361], line_28[359], line_27[357], line_26[355], line_25[353], line_24[351], line_23[349], line_22[347], line_21[345], line_20[343], line_19[341], line_18[339], line_17[337], line_16[335], line_15[333], line_14[331], line_13[329], line_12[327], line_11[325], line_10[323], line_9[321], line_8[319], line_7[317], line_6[315], line_5[313], line_4[311], line_3[309], line_2[307], line_1[305] };
assign col_560 = {line_128[560], line_127[558], line_126[556], line_125[554], line_124[552], line_123[550], line_122[548], line_121[546], line_120[544], line_119[542], line_118[540], line_117[538], line_116[536], line_115[534], line_114[532], line_113[530], line_112[528], line_111[526], line_110[524], line_109[522], line_108[520], line_107[518], line_106[516], line_105[514], line_104[512], line_103[510], line_102[508], line_101[506], line_100[504], line_99[502], line_98[500], line_97[498], line_96[496], line_95[494], line_94[492], line_93[490], line_92[488], line_91[486], line_90[484], line_89[482], line_88[480], line_87[478], line_86[476], line_85[474], line_84[472], line_83[470], line_82[468], line_81[466], line_80[464], line_79[462], line_78[460], line_77[458], line_76[456], line_75[454], line_74[452], line_73[450], line_72[448], line_71[446], line_70[444], line_69[442], line_68[440], line_67[438], line_66[436], line_65[434], line_64[432], line_63[430], line_62[428], line_61[426], line_60[424], line_59[422], line_58[420], line_57[418], line_56[416], line_55[414], line_54[412], line_53[410], line_52[408], line_51[406], line_50[404], line_49[402], line_48[400], line_47[398], line_46[396], line_45[394], line_44[392], line_43[390], line_42[388], line_41[386], line_40[384], line_39[382], line_38[380], line_37[378], line_36[376], line_35[374], line_34[372], line_33[370], line_32[368], line_31[366], line_30[364], line_29[362], line_28[360], line_27[358], line_26[356], line_25[354], line_24[352], line_23[350], line_22[348], line_21[346], line_20[344], line_19[342], line_18[340], line_17[338], line_16[336], line_15[334], line_14[332], line_13[330], line_12[328], line_11[326], line_10[324], line_9[322], line_8[320], line_7[318], line_6[316], line_5[314], line_4[312], line_3[310], line_2[308], line_1[306] };
assign col_561 = {line_128[561], line_127[559], line_126[557], line_125[555], line_124[553], line_123[551], line_122[549], line_121[547], line_120[545], line_119[543], line_118[541], line_117[539], line_116[537], line_115[535], line_114[533], line_113[531], line_112[529], line_111[527], line_110[525], line_109[523], line_108[521], line_107[519], line_106[517], line_105[515], line_104[513], line_103[511], line_102[509], line_101[507], line_100[505], line_99[503], line_98[501], line_97[499], line_96[497], line_95[495], line_94[493], line_93[491], line_92[489], line_91[487], line_90[485], line_89[483], line_88[481], line_87[479], line_86[477], line_85[475], line_84[473], line_83[471], line_82[469], line_81[467], line_80[465], line_79[463], line_78[461], line_77[459], line_76[457], line_75[455], line_74[453], line_73[451], line_72[449], line_71[447], line_70[445], line_69[443], line_68[441], line_67[439], line_66[437], line_65[435], line_64[433], line_63[431], line_62[429], line_61[427], line_60[425], line_59[423], line_58[421], line_57[419], line_56[417], line_55[415], line_54[413], line_53[411], line_52[409], line_51[407], line_50[405], line_49[403], line_48[401], line_47[399], line_46[397], line_45[395], line_44[393], line_43[391], line_42[389], line_41[387], line_40[385], line_39[383], line_38[381], line_37[379], line_36[377], line_35[375], line_34[373], line_33[371], line_32[369], line_31[367], line_30[365], line_29[363], line_28[361], line_27[359], line_26[357], line_25[355], line_24[353], line_23[351], line_22[349], line_21[347], line_20[345], line_19[343], line_18[341], line_17[339], line_16[337], line_15[335], line_14[333], line_13[331], line_12[329], line_11[327], line_10[325], line_9[323], line_8[321], line_7[319], line_6[317], line_5[315], line_4[313], line_3[311], line_2[309], line_1[307] };
assign col_562 = {line_128[562], line_127[560], line_126[558], line_125[556], line_124[554], line_123[552], line_122[550], line_121[548], line_120[546], line_119[544], line_118[542], line_117[540], line_116[538], line_115[536], line_114[534], line_113[532], line_112[530], line_111[528], line_110[526], line_109[524], line_108[522], line_107[520], line_106[518], line_105[516], line_104[514], line_103[512], line_102[510], line_101[508], line_100[506], line_99[504], line_98[502], line_97[500], line_96[498], line_95[496], line_94[494], line_93[492], line_92[490], line_91[488], line_90[486], line_89[484], line_88[482], line_87[480], line_86[478], line_85[476], line_84[474], line_83[472], line_82[470], line_81[468], line_80[466], line_79[464], line_78[462], line_77[460], line_76[458], line_75[456], line_74[454], line_73[452], line_72[450], line_71[448], line_70[446], line_69[444], line_68[442], line_67[440], line_66[438], line_65[436], line_64[434], line_63[432], line_62[430], line_61[428], line_60[426], line_59[424], line_58[422], line_57[420], line_56[418], line_55[416], line_54[414], line_53[412], line_52[410], line_51[408], line_50[406], line_49[404], line_48[402], line_47[400], line_46[398], line_45[396], line_44[394], line_43[392], line_42[390], line_41[388], line_40[386], line_39[384], line_38[382], line_37[380], line_36[378], line_35[376], line_34[374], line_33[372], line_32[370], line_31[368], line_30[366], line_29[364], line_28[362], line_27[360], line_26[358], line_25[356], line_24[354], line_23[352], line_22[350], line_21[348], line_20[346], line_19[344], line_18[342], line_17[340], line_16[338], line_15[336], line_14[334], line_13[332], line_12[330], line_11[328], line_10[326], line_9[324], line_8[322], line_7[320], line_6[318], line_5[316], line_4[314], line_3[312], line_2[310], line_1[308] };
assign col_563 = {line_128[563], line_127[561], line_126[559], line_125[557], line_124[555], line_123[553], line_122[551], line_121[549], line_120[547], line_119[545], line_118[543], line_117[541], line_116[539], line_115[537], line_114[535], line_113[533], line_112[531], line_111[529], line_110[527], line_109[525], line_108[523], line_107[521], line_106[519], line_105[517], line_104[515], line_103[513], line_102[511], line_101[509], line_100[507], line_99[505], line_98[503], line_97[501], line_96[499], line_95[497], line_94[495], line_93[493], line_92[491], line_91[489], line_90[487], line_89[485], line_88[483], line_87[481], line_86[479], line_85[477], line_84[475], line_83[473], line_82[471], line_81[469], line_80[467], line_79[465], line_78[463], line_77[461], line_76[459], line_75[457], line_74[455], line_73[453], line_72[451], line_71[449], line_70[447], line_69[445], line_68[443], line_67[441], line_66[439], line_65[437], line_64[435], line_63[433], line_62[431], line_61[429], line_60[427], line_59[425], line_58[423], line_57[421], line_56[419], line_55[417], line_54[415], line_53[413], line_52[411], line_51[409], line_50[407], line_49[405], line_48[403], line_47[401], line_46[399], line_45[397], line_44[395], line_43[393], line_42[391], line_41[389], line_40[387], line_39[385], line_38[383], line_37[381], line_36[379], line_35[377], line_34[375], line_33[373], line_32[371], line_31[369], line_30[367], line_29[365], line_28[363], line_27[361], line_26[359], line_25[357], line_24[355], line_23[353], line_22[351], line_21[349], line_20[347], line_19[345], line_18[343], line_17[341], line_16[339], line_15[337], line_14[335], line_13[333], line_12[331], line_11[329], line_10[327], line_9[325], line_8[323], line_7[321], line_6[319], line_5[317], line_4[315], line_3[313], line_2[311], line_1[309] };
assign col_564 = {line_128[564], line_127[562], line_126[560], line_125[558], line_124[556], line_123[554], line_122[552], line_121[550], line_120[548], line_119[546], line_118[544], line_117[542], line_116[540], line_115[538], line_114[536], line_113[534], line_112[532], line_111[530], line_110[528], line_109[526], line_108[524], line_107[522], line_106[520], line_105[518], line_104[516], line_103[514], line_102[512], line_101[510], line_100[508], line_99[506], line_98[504], line_97[502], line_96[500], line_95[498], line_94[496], line_93[494], line_92[492], line_91[490], line_90[488], line_89[486], line_88[484], line_87[482], line_86[480], line_85[478], line_84[476], line_83[474], line_82[472], line_81[470], line_80[468], line_79[466], line_78[464], line_77[462], line_76[460], line_75[458], line_74[456], line_73[454], line_72[452], line_71[450], line_70[448], line_69[446], line_68[444], line_67[442], line_66[440], line_65[438], line_64[436], line_63[434], line_62[432], line_61[430], line_60[428], line_59[426], line_58[424], line_57[422], line_56[420], line_55[418], line_54[416], line_53[414], line_52[412], line_51[410], line_50[408], line_49[406], line_48[404], line_47[402], line_46[400], line_45[398], line_44[396], line_43[394], line_42[392], line_41[390], line_40[388], line_39[386], line_38[384], line_37[382], line_36[380], line_35[378], line_34[376], line_33[374], line_32[372], line_31[370], line_30[368], line_29[366], line_28[364], line_27[362], line_26[360], line_25[358], line_24[356], line_23[354], line_22[352], line_21[350], line_20[348], line_19[346], line_18[344], line_17[342], line_16[340], line_15[338], line_14[336], line_13[334], line_12[332], line_11[330], line_10[328], line_9[326], line_8[324], line_7[322], line_6[320], line_5[318], line_4[316], line_3[314], line_2[312], line_1[310] };
assign col_565 = {line_128[565], line_127[563], line_126[561], line_125[559], line_124[557], line_123[555], line_122[553], line_121[551], line_120[549], line_119[547], line_118[545], line_117[543], line_116[541], line_115[539], line_114[537], line_113[535], line_112[533], line_111[531], line_110[529], line_109[527], line_108[525], line_107[523], line_106[521], line_105[519], line_104[517], line_103[515], line_102[513], line_101[511], line_100[509], line_99[507], line_98[505], line_97[503], line_96[501], line_95[499], line_94[497], line_93[495], line_92[493], line_91[491], line_90[489], line_89[487], line_88[485], line_87[483], line_86[481], line_85[479], line_84[477], line_83[475], line_82[473], line_81[471], line_80[469], line_79[467], line_78[465], line_77[463], line_76[461], line_75[459], line_74[457], line_73[455], line_72[453], line_71[451], line_70[449], line_69[447], line_68[445], line_67[443], line_66[441], line_65[439], line_64[437], line_63[435], line_62[433], line_61[431], line_60[429], line_59[427], line_58[425], line_57[423], line_56[421], line_55[419], line_54[417], line_53[415], line_52[413], line_51[411], line_50[409], line_49[407], line_48[405], line_47[403], line_46[401], line_45[399], line_44[397], line_43[395], line_42[393], line_41[391], line_40[389], line_39[387], line_38[385], line_37[383], line_36[381], line_35[379], line_34[377], line_33[375], line_32[373], line_31[371], line_30[369], line_29[367], line_28[365], line_27[363], line_26[361], line_25[359], line_24[357], line_23[355], line_22[353], line_21[351], line_20[349], line_19[347], line_18[345], line_17[343], line_16[341], line_15[339], line_14[337], line_13[335], line_12[333], line_11[331], line_10[329], line_9[327], line_8[325], line_7[323], line_6[321], line_5[319], line_4[317], line_3[315], line_2[313], line_1[311] };
assign col_566 = {line_128[566], line_127[564], line_126[562], line_125[560], line_124[558], line_123[556], line_122[554], line_121[552], line_120[550], line_119[548], line_118[546], line_117[544], line_116[542], line_115[540], line_114[538], line_113[536], line_112[534], line_111[532], line_110[530], line_109[528], line_108[526], line_107[524], line_106[522], line_105[520], line_104[518], line_103[516], line_102[514], line_101[512], line_100[510], line_99[508], line_98[506], line_97[504], line_96[502], line_95[500], line_94[498], line_93[496], line_92[494], line_91[492], line_90[490], line_89[488], line_88[486], line_87[484], line_86[482], line_85[480], line_84[478], line_83[476], line_82[474], line_81[472], line_80[470], line_79[468], line_78[466], line_77[464], line_76[462], line_75[460], line_74[458], line_73[456], line_72[454], line_71[452], line_70[450], line_69[448], line_68[446], line_67[444], line_66[442], line_65[440], line_64[438], line_63[436], line_62[434], line_61[432], line_60[430], line_59[428], line_58[426], line_57[424], line_56[422], line_55[420], line_54[418], line_53[416], line_52[414], line_51[412], line_50[410], line_49[408], line_48[406], line_47[404], line_46[402], line_45[400], line_44[398], line_43[396], line_42[394], line_41[392], line_40[390], line_39[388], line_38[386], line_37[384], line_36[382], line_35[380], line_34[378], line_33[376], line_32[374], line_31[372], line_30[370], line_29[368], line_28[366], line_27[364], line_26[362], line_25[360], line_24[358], line_23[356], line_22[354], line_21[352], line_20[350], line_19[348], line_18[346], line_17[344], line_16[342], line_15[340], line_14[338], line_13[336], line_12[334], line_11[332], line_10[330], line_9[328], line_8[326], line_7[324], line_6[322], line_5[320], line_4[318], line_3[316], line_2[314], line_1[312] };
assign col_567 = {line_128[567], line_127[565], line_126[563], line_125[561], line_124[559], line_123[557], line_122[555], line_121[553], line_120[551], line_119[549], line_118[547], line_117[545], line_116[543], line_115[541], line_114[539], line_113[537], line_112[535], line_111[533], line_110[531], line_109[529], line_108[527], line_107[525], line_106[523], line_105[521], line_104[519], line_103[517], line_102[515], line_101[513], line_100[511], line_99[509], line_98[507], line_97[505], line_96[503], line_95[501], line_94[499], line_93[497], line_92[495], line_91[493], line_90[491], line_89[489], line_88[487], line_87[485], line_86[483], line_85[481], line_84[479], line_83[477], line_82[475], line_81[473], line_80[471], line_79[469], line_78[467], line_77[465], line_76[463], line_75[461], line_74[459], line_73[457], line_72[455], line_71[453], line_70[451], line_69[449], line_68[447], line_67[445], line_66[443], line_65[441], line_64[439], line_63[437], line_62[435], line_61[433], line_60[431], line_59[429], line_58[427], line_57[425], line_56[423], line_55[421], line_54[419], line_53[417], line_52[415], line_51[413], line_50[411], line_49[409], line_48[407], line_47[405], line_46[403], line_45[401], line_44[399], line_43[397], line_42[395], line_41[393], line_40[391], line_39[389], line_38[387], line_37[385], line_36[383], line_35[381], line_34[379], line_33[377], line_32[375], line_31[373], line_30[371], line_29[369], line_28[367], line_27[365], line_26[363], line_25[361], line_24[359], line_23[357], line_22[355], line_21[353], line_20[351], line_19[349], line_18[347], line_17[345], line_16[343], line_15[341], line_14[339], line_13[337], line_12[335], line_11[333], line_10[331], line_9[329], line_8[327], line_7[325], line_6[323], line_5[321], line_4[319], line_3[317], line_2[315], line_1[313] };
assign col_568 = {line_128[568], line_127[566], line_126[564], line_125[562], line_124[560], line_123[558], line_122[556], line_121[554], line_120[552], line_119[550], line_118[548], line_117[546], line_116[544], line_115[542], line_114[540], line_113[538], line_112[536], line_111[534], line_110[532], line_109[530], line_108[528], line_107[526], line_106[524], line_105[522], line_104[520], line_103[518], line_102[516], line_101[514], line_100[512], line_99[510], line_98[508], line_97[506], line_96[504], line_95[502], line_94[500], line_93[498], line_92[496], line_91[494], line_90[492], line_89[490], line_88[488], line_87[486], line_86[484], line_85[482], line_84[480], line_83[478], line_82[476], line_81[474], line_80[472], line_79[470], line_78[468], line_77[466], line_76[464], line_75[462], line_74[460], line_73[458], line_72[456], line_71[454], line_70[452], line_69[450], line_68[448], line_67[446], line_66[444], line_65[442], line_64[440], line_63[438], line_62[436], line_61[434], line_60[432], line_59[430], line_58[428], line_57[426], line_56[424], line_55[422], line_54[420], line_53[418], line_52[416], line_51[414], line_50[412], line_49[410], line_48[408], line_47[406], line_46[404], line_45[402], line_44[400], line_43[398], line_42[396], line_41[394], line_40[392], line_39[390], line_38[388], line_37[386], line_36[384], line_35[382], line_34[380], line_33[378], line_32[376], line_31[374], line_30[372], line_29[370], line_28[368], line_27[366], line_26[364], line_25[362], line_24[360], line_23[358], line_22[356], line_21[354], line_20[352], line_19[350], line_18[348], line_17[346], line_16[344], line_15[342], line_14[340], line_13[338], line_12[336], line_11[334], line_10[332], line_9[330], line_8[328], line_7[326], line_6[324], line_5[322], line_4[320], line_3[318], line_2[316], line_1[314] };
assign col_569 = {line_128[569], line_127[567], line_126[565], line_125[563], line_124[561], line_123[559], line_122[557], line_121[555], line_120[553], line_119[551], line_118[549], line_117[547], line_116[545], line_115[543], line_114[541], line_113[539], line_112[537], line_111[535], line_110[533], line_109[531], line_108[529], line_107[527], line_106[525], line_105[523], line_104[521], line_103[519], line_102[517], line_101[515], line_100[513], line_99[511], line_98[509], line_97[507], line_96[505], line_95[503], line_94[501], line_93[499], line_92[497], line_91[495], line_90[493], line_89[491], line_88[489], line_87[487], line_86[485], line_85[483], line_84[481], line_83[479], line_82[477], line_81[475], line_80[473], line_79[471], line_78[469], line_77[467], line_76[465], line_75[463], line_74[461], line_73[459], line_72[457], line_71[455], line_70[453], line_69[451], line_68[449], line_67[447], line_66[445], line_65[443], line_64[441], line_63[439], line_62[437], line_61[435], line_60[433], line_59[431], line_58[429], line_57[427], line_56[425], line_55[423], line_54[421], line_53[419], line_52[417], line_51[415], line_50[413], line_49[411], line_48[409], line_47[407], line_46[405], line_45[403], line_44[401], line_43[399], line_42[397], line_41[395], line_40[393], line_39[391], line_38[389], line_37[387], line_36[385], line_35[383], line_34[381], line_33[379], line_32[377], line_31[375], line_30[373], line_29[371], line_28[369], line_27[367], line_26[365], line_25[363], line_24[361], line_23[359], line_22[357], line_21[355], line_20[353], line_19[351], line_18[349], line_17[347], line_16[345], line_15[343], line_14[341], line_13[339], line_12[337], line_11[335], line_10[333], line_9[331], line_8[329], line_7[327], line_6[325], line_5[323], line_4[321], line_3[319], line_2[317], line_1[315] };
assign col_570 = {line_128[570], line_127[568], line_126[566], line_125[564], line_124[562], line_123[560], line_122[558], line_121[556], line_120[554], line_119[552], line_118[550], line_117[548], line_116[546], line_115[544], line_114[542], line_113[540], line_112[538], line_111[536], line_110[534], line_109[532], line_108[530], line_107[528], line_106[526], line_105[524], line_104[522], line_103[520], line_102[518], line_101[516], line_100[514], line_99[512], line_98[510], line_97[508], line_96[506], line_95[504], line_94[502], line_93[500], line_92[498], line_91[496], line_90[494], line_89[492], line_88[490], line_87[488], line_86[486], line_85[484], line_84[482], line_83[480], line_82[478], line_81[476], line_80[474], line_79[472], line_78[470], line_77[468], line_76[466], line_75[464], line_74[462], line_73[460], line_72[458], line_71[456], line_70[454], line_69[452], line_68[450], line_67[448], line_66[446], line_65[444], line_64[442], line_63[440], line_62[438], line_61[436], line_60[434], line_59[432], line_58[430], line_57[428], line_56[426], line_55[424], line_54[422], line_53[420], line_52[418], line_51[416], line_50[414], line_49[412], line_48[410], line_47[408], line_46[406], line_45[404], line_44[402], line_43[400], line_42[398], line_41[396], line_40[394], line_39[392], line_38[390], line_37[388], line_36[386], line_35[384], line_34[382], line_33[380], line_32[378], line_31[376], line_30[374], line_29[372], line_28[370], line_27[368], line_26[366], line_25[364], line_24[362], line_23[360], line_22[358], line_21[356], line_20[354], line_19[352], line_18[350], line_17[348], line_16[346], line_15[344], line_14[342], line_13[340], line_12[338], line_11[336], line_10[334], line_9[332], line_8[330], line_7[328], line_6[326], line_5[324], line_4[322], line_3[320], line_2[318], line_1[316] };
assign col_571 = {line_128[571], line_127[569], line_126[567], line_125[565], line_124[563], line_123[561], line_122[559], line_121[557], line_120[555], line_119[553], line_118[551], line_117[549], line_116[547], line_115[545], line_114[543], line_113[541], line_112[539], line_111[537], line_110[535], line_109[533], line_108[531], line_107[529], line_106[527], line_105[525], line_104[523], line_103[521], line_102[519], line_101[517], line_100[515], line_99[513], line_98[511], line_97[509], line_96[507], line_95[505], line_94[503], line_93[501], line_92[499], line_91[497], line_90[495], line_89[493], line_88[491], line_87[489], line_86[487], line_85[485], line_84[483], line_83[481], line_82[479], line_81[477], line_80[475], line_79[473], line_78[471], line_77[469], line_76[467], line_75[465], line_74[463], line_73[461], line_72[459], line_71[457], line_70[455], line_69[453], line_68[451], line_67[449], line_66[447], line_65[445], line_64[443], line_63[441], line_62[439], line_61[437], line_60[435], line_59[433], line_58[431], line_57[429], line_56[427], line_55[425], line_54[423], line_53[421], line_52[419], line_51[417], line_50[415], line_49[413], line_48[411], line_47[409], line_46[407], line_45[405], line_44[403], line_43[401], line_42[399], line_41[397], line_40[395], line_39[393], line_38[391], line_37[389], line_36[387], line_35[385], line_34[383], line_33[381], line_32[379], line_31[377], line_30[375], line_29[373], line_28[371], line_27[369], line_26[367], line_25[365], line_24[363], line_23[361], line_22[359], line_21[357], line_20[355], line_19[353], line_18[351], line_17[349], line_16[347], line_15[345], line_14[343], line_13[341], line_12[339], line_11[337], line_10[335], line_9[333], line_8[331], line_7[329], line_6[327], line_5[325], line_4[323], line_3[321], line_2[319], line_1[317] };
assign col_572 = {line_128[572], line_127[570], line_126[568], line_125[566], line_124[564], line_123[562], line_122[560], line_121[558], line_120[556], line_119[554], line_118[552], line_117[550], line_116[548], line_115[546], line_114[544], line_113[542], line_112[540], line_111[538], line_110[536], line_109[534], line_108[532], line_107[530], line_106[528], line_105[526], line_104[524], line_103[522], line_102[520], line_101[518], line_100[516], line_99[514], line_98[512], line_97[510], line_96[508], line_95[506], line_94[504], line_93[502], line_92[500], line_91[498], line_90[496], line_89[494], line_88[492], line_87[490], line_86[488], line_85[486], line_84[484], line_83[482], line_82[480], line_81[478], line_80[476], line_79[474], line_78[472], line_77[470], line_76[468], line_75[466], line_74[464], line_73[462], line_72[460], line_71[458], line_70[456], line_69[454], line_68[452], line_67[450], line_66[448], line_65[446], line_64[444], line_63[442], line_62[440], line_61[438], line_60[436], line_59[434], line_58[432], line_57[430], line_56[428], line_55[426], line_54[424], line_53[422], line_52[420], line_51[418], line_50[416], line_49[414], line_48[412], line_47[410], line_46[408], line_45[406], line_44[404], line_43[402], line_42[400], line_41[398], line_40[396], line_39[394], line_38[392], line_37[390], line_36[388], line_35[386], line_34[384], line_33[382], line_32[380], line_31[378], line_30[376], line_29[374], line_28[372], line_27[370], line_26[368], line_25[366], line_24[364], line_23[362], line_22[360], line_21[358], line_20[356], line_19[354], line_18[352], line_17[350], line_16[348], line_15[346], line_14[344], line_13[342], line_12[340], line_11[338], line_10[336], line_9[334], line_8[332], line_7[330], line_6[328], line_5[326], line_4[324], line_3[322], line_2[320], line_1[318] };
assign col_573 = {line_128[573], line_127[571], line_126[569], line_125[567], line_124[565], line_123[563], line_122[561], line_121[559], line_120[557], line_119[555], line_118[553], line_117[551], line_116[549], line_115[547], line_114[545], line_113[543], line_112[541], line_111[539], line_110[537], line_109[535], line_108[533], line_107[531], line_106[529], line_105[527], line_104[525], line_103[523], line_102[521], line_101[519], line_100[517], line_99[515], line_98[513], line_97[511], line_96[509], line_95[507], line_94[505], line_93[503], line_92[501], line_91[499], line_90[497], line_89[495], line_88[493], line_87[491], line_86[489], line_85[487], line_84[485], line_83[483], line_82[481], line_81[479], line_80[477], line_79[475], line_78[473], line_77[471], line_76[469], line_75[467], line_74[465], line_73[463], line_72[461], line_71[459], line_70[457], line_69[455], line_68[453], line_67[451], line_66[449], line_65[447], line_64[445], line_63[443], line_62[441], line_61[439], line_60[437], line_59[435], line_58[433], line_57[431], line_56[429], line_55[427], line_54[425], line_53[423], line_52[421], line_51[419], line_50[417], line_49[415], line_48[413], line_47[411], line_46[409], line_45[407], line_44[405], line_43[403], line_42[401], line_41[399], line_40[397], line_39[395], line_38[393], line_37[391], line_36[389], line_35[387], line_34[385], line_33[383], line_32[381], line_31[379], line_30[377], line_29[375], line_28[373], line_27[371], line_26[369], line_25[367], line_24[365], line_23[363], line_22[361], line_21[359], line_20[357], line_19[355], line_18[353], line_17[351], line_16[349], line_15[347], line_14[345], line_13[343], line_12[341], line_11[339], line_10[337], line_9[335], line_8[333], line_7[331], line_6[329], line_5[327], line_4[325], line_3[323], line_2[321], line_1[319] };
assign col_574 = {line_128[574], line_127[572], line_126[570], line_125[568], line_124[566], line_123[564], line_122[562], line_121[560], line_120[558], line_119[556], line_118[554], line_117[552], line_116[550], line_115[548], line_114[546], line_113[544], line_112[542], line_111[540], line_110[538], line_109[536], line_108[534], line_107[532], line_106[530], line_105[528], line_104[526], line_103[524], line_102[522], line_101[520], line_100[518], line_99[516], line_98[514], line_97[512], line_96[510], line_95[508], line_94[506], line_93[504], line_92[502], line_91[500], line_90[498], line_89[496], line_88[494], line_87[492], line_86[490], line_85[488], line_84[486], line_83[484], line_82[482], line_81[480], line_80[478], line_79[476], line_78[474], line_77[472], line_76[470], line_75[468], line_74[466], line_73[464], line_72[462], line_71[460], line_70[458], line_69[456], line_68[454], line_67[452], line_66[450], line_65[448], line_64[446], line_63[444], line_62[442], line_61[440], line_60[438], line_59[436], line_58[434], line_57[432], line_56[430], line_55[428], line_54[426], line_53[424], line_52[422], line_51[420], line_50[418], line_49[416], line_48[414], line_47[412], line_46[410], line_45[408], line_44[406], line_43[404], line_42[402], line_41[400], line_40[398], line_39[396], line_38[394], line_37[392], line_36[390], line_35[388], line_34[386], line_33[384], line_32[382], line_31[380], line_30[378], line_29[376], line_28[374], line_27[372], line_26[370], line_25[368], line_24[366], line_23[364], line_22[362], line_21[360], line_20[358], line_19[356], line_18[354], line_17[352], line_16[350], line_15[348], line_14[346], line_13[344], line_12[342], line_11[340], line_10[338], line_9[336], line_8[334], line_7[332], line_6[330], line_5[328], line_4[326], line_3[324], line_2[322], line_1[320] };
assign col_575 = {line_128[575], line_127[573], line_126[571], line_125[569], line_124[567], line_123[565], line_122[563], line_121[561], line_120[559], line_119[557], line_118[555], line_117[553], line_116[551], line_115[549], line_114[547], line_113[545], line_112[543], line_111[541], line_110[539], line_109[537], line_108[535], line_107[533], line_106[531], line_105[529], line_104[527], line_103[525], line_102[523], line_101[521], line_100[519], line_99[517], line_98[515], line_97[513], line_96[511], line_95[509], line_94[507], line_93[505], line_92[503], line_91[501], line_90[499], line_89[497], line_88[495], line_87[493], line_86[491], line_85[489], line_84[487], line_83[485], line_82[483], line_81[481], line_80[479], line_79[477], line_78[475], line_77[473], line_76[471], line_75[469], line_74[467], line_73[465], line_72[463], line_71[461], line_70[459], line_69[457], line_68[455], line_67[453], line_66[451], line_65[449], line_64[447], line_63[445], line_62[443], line_61[441], line_60[439], line_59[437], line_58[435], line_57[433], line_56[431], line_55[429], line_54[427], line_53[425], line_52[423], line_51[421], line_50[419], line_49[417], line_48[415], line_47[413], line_46[411], line_45[409], line_44[407], line_43[405], line_42[403], line_41[401], line_40[399], line_39[397], line_38[395], line_37[393], line_36[391], line_35[389], line_34[387], line_33[385], line_32[383], line_31[381], line_30[379], line_29[377], line_28[375], line_27[373], line_26[371], line_25[369], line_24[367], line_23[365], line_22[363], line_21[361], line_20[359], line_19[357], line_18[355], line_17[353], line_16[351], line_15[349], line_14[347], line_13[345], line_12[343], line_11[341], line_10[339], line_9[337], line_8[335], line_7[333], line_6[331], line_5[329], line_4[327], line_3[325], line_2[323], line_1[321] };
assign col_576 = {line_128[576], line_127[574], line_126[572], line_125[570], line_124[568], line_123[566], line_122[564], line_121[562], line_120[560], line_119[558], line_118[556], line_117[554], line_116[552], line_115[550], line_114[548], line_113[546], line_112[544], line_111[542], line_110[540], line_109[538], line_108[536], line_107[534], line_106[532], line_105[530], line_104[528], line_103[526], line_102[524], line_101[522], line_100[520], line_99[518], line_98[516], line_97[514], line_96[512], line_95[510], line_94[508], line_93[506], line_92[504], line_91[502], line_90[500], line_89[498], line_88[496], line_87[494], line_86[492], line_85[490], line_84[488], line_83[486], line_82[484], line_81[482], line_80[480], line_79[478], line_78[476], line_77[474], line_76[472], line_75[470], line_74[468], line_73[466], line_72[464], line_71[462], line_70[460], line_69[458], line_68[456], line_67[454], line_66[452], line_65[450], line_64[448], line_63[446], line_62[444], line_61[442], line_60[440], line_59[438], line_58[436], line_57[434], line_56[432], line_55[430], line_54[428], line_53[426], line_52[424], line_51[422], line_50[420], line_49[418], line_48[416], line_47[414], line_46[412], line_45[410], line_44[408], line_43[406], line_42[404], line_41[402], line_40[400], line_39[398], line_38[396], line_37[394], line_36[392], line_35[390], line_34[388], line_33[386], line_32[384], line_31[382], line_30[380], line_29[378], line_28[376], line_27[374], line_26[372], line_25[370], line_24[368], line_23[366], line_22[364], line_21[362], line_20[360], line_19[358], line_18[356], line_17[354], line_16[352], line_15[350], line_14[348], line_13[346], line_12[344], line_11[342], line_10[340], line_9[338], line_8[336], line_7[334], line_6[332], line_5[330], line_4[328], line_3[326], line_2[324], line_1[322] };
assign col_577 = {line_128[577], line_127[575], line_126[573], line_125[571], line_124[569], line_123[567], line_122[565], line_121[563], line_120[561], line_119[559], line_118[557], line_117[555], line_116[553], line_115[551], line_114[549], line_113[547], line_112[545], line_111[543], line_110[541], line_109[539], line_108[537], line_107[535], line_106[533], line_105[531], line_104[529], line_103[527], line_102[525], line_101[523], line_100[521], line_99[519], line_98[517], line_97[515], line_96[513], line_95[511], line_94[509], line_93[507], line_92[505], line_91[503], line_90[501], line_89[499], line_88[497], line_87[495], line_86[493], line_85[491], line_84[489], line_83[487], line_82[485], line_81[483], line_80[481], line_79[479], line_78[477], line_77[475], line_76[473], line_75[471], line_74[469], line_73[467], line_72[465], line_71[463], line_70[461], line_69[459], line_68[457], line_67[455], line_66[453], line_65[451], line_64[449], line_63[447], line_62[445], line_61[443], line_60[441], line_59[439], line_58[437], line_57[435], line_56[433], line_55[431], line_54[429], line_53[427], line_52[425], line_51[423], line_50[421], line_49[419], line_48[417], line_47[415], line_46[413], line_45[411], line_44[409], line_43[407], line_42[405], line_41[403], line_40[401], line_39[399], line_38[397], line_37[395], line_36[393], line_35[391], line_34[389], line_33[387], line_32[385], line_31[383], line_30[381], line_29[379], line_28[377], line_27[375], line_26[373], line_25[371], line_24[369], line_23[367], line_22[365], line_21[363], line_20[361], line_19[359], line_18[357], line_17[355], line_16[353], line_15[351], line_14[349], line_13[347], line_12[345], line_11[343], line_10[341], line_9[339], line_8[337], line_7[335], line_6[333], line_5[331], line_4[329], line_3[327], line_2[325], line_1[323] };
assign col_578 = {line_128[578], line_127[576], line_126[574], line_125[572], line_124[570], line_123[568], line_122[566], line_121[564], line_120[562], line_119[560], line_118[558], line_117[556], line_116[554], line_115[552], line_114[550], line_113[548], line_112[546], line_111[544], line_110[542], line_109[540], line_108[538], line_107[536], line_106[534], line_105[532], line_104[530], line_103[528], line_102[526], line_101[524], line_100[522], line_99[520], line_98[518], line_97[516], line_96[514], line_95[512], line_94[510], line_93[508], line_92[506], line_91[504], line_90[502], line_89[500], line_88[498], line_87[496], line_86[494], line_85[492], line_84[490], line_83[488], line_82[486], line_81[484], line_80[482], line_79[480], line_78[478], line_77[476], line_76[474], line_75[472], line_74[470], line_73[468], line_72[466], line_71[464], line_70[462], line_69[460], line_68[458], line_67[456], line_66[454], line_65[452], line_64[450], line_63[448], line_62[446], line_61[444], line_60[442], line_59[440], line_58[438], line_57[436], line_56[434], line_55[432], line_54[430], line_53[428], line_52[426], line_51[424], line_50[422], line_49[420], line_48[418], line_47[416], line_46[414], line_45[412], line_44[410], line_43[408], line_42[406], line_41[404], line_40[402], line_39[400], line_38[398], line_37[396], line_36[394], line_35[392], line_34[390], line_33[388], line_32[386], line_31[384], line_30[382], line_29[380], line_28[378], line_27[376], line_26[374], line_25[372], line_24[370], line_23[368], line_22[366], line_21[364], line_20[362], line_19[360], line_18[358], line_17[356], line_16[354], line_15[352], line_14[350], line_13[348], line_12[346], line_11[344], line_10[342], line_9[340], line_8[338], line_7[336], line_6[334], line_5[332], line_4[330], line_3[328], line_2[326], line_1[324] };
assign col_579 = {line_128[579], line_127[577], line_126[575], line_125[573], line_124[571], line_123[569], line_122[567], line_121[565], line_120[563], line_119[561], line_118[559], line_117[557], line_116[555], line_115[553], line_114[551], line_113[549], line_112[547], line_111[545], line_110[543], line_109[541], line_108[539], line_107[537], line_106[535], line_105[533], line_104[531], line_103[529], line_102[527], line_101[525], line_100[523], line_99[521], line_98[519], line_97[517], line_96[515], line_95[513], line_94[511], line_93[509], line_92[507], line_91[505], line_90[503], line_89[501], line_88[499], line_87[497], line_86[495], line_85[493], line_84[491], line_83[489], line_82[487], line_81[485], line_80[483], line_79[481], line_78[479], line_77[477], line_76[475], line_75[473], line_74[471], line_73[469], line_72[467], line_71[465], line_70[463], line_69[461], line_68[459], line_67[457], line_66[455], line_65[453], line_64[451], line_63[449], line_62[447], line_61[445], line_60[443], line_59[441], line_58[439], line_57[437], line_56[435], line_55[433], line_54[431], line_53[429], line_52[427], line_51[425], line_50[423], line_49[421], line_48[419], line_47[417], line_46[415], line_45[413], line_44[411], line_43[409], line_42[407], line_41[405], line_40[403], line_39[401], line_38[399], line_37[397], line_36[395], line_35[393], line_34[391], line_33[389], line_32[387], line_31[385], line_30[383], line_29[381], line_28[379], line_27[377], line_26[375], line_25[373], line_24[371], line_23[369], line_22[367], line_21[365], line_20[363], line_19[361], line_18[359], line_17[357], line_16[355], line_15[353], line_14[351], line_13[349], line_12[347], line_11[345], line_10[343], line_9[341], line_8[339], line_7[337], line_6[335], line_5[333], line_4[331], line_3[329], line_2[327], line_1[325] };
assign col_580 = {line_128[580], line_127[578], line_126[576], line_125[574], line_124[572], line_123[570], line_122[568], line_121[566], line_120[564], line_119[562], line_118[560], line_117[558], line_116[556], line_115[554], line_114[552], line_113[550], line_112[548], line_111[546], line_110[544], line_109[542], line_108[540], line_107[538], line_106[536], line_105[534], line_104[532], line_103[530], line_102[528], line_101[526], line_100[524], line_99[522], line_98[520], line_97[518], line_96[516], line_95[514], line_94[512], line_93[510], line_92[508], line_91[506], line_90[504], line_89[502], line_88[500], line_87[498], line_86[496], line_85[494], line_84[492], line_83[490], line_82[488], line_81[486], line_80[484], line_79[482], line_78[480], line_77[478], line_76[476], line_75[474], line_74[472], line_73[470], line_72[468], line_71[466], line_70[464], line_69[462], line_68[460], line_67[458], line_66[456], line_65[454], line_64[452], line_63[450], line_62[448], line_61[446], line_60[444], line_59[442], line_58[440], line_57[438], line_56[436], line_55[434], line_54[432], line_53[430], line_52[428], line_51[426], line_50[424], line_49[422], line_48[420], line_47[418], line_46[416], line_45[414], line_44[412], line_43[410], line_42[408], line_41[406], line_40[404], line_39[402], line_38[400], line_37[398], line_36[396], line_35[394], line_34[392], line_33[390], line_32[388], line_31[386], line_30[384], line_29[382], line_28[380], line_27[378], line_26[376], line_25[374], line_24[372], line_23[370], line_22[368], line_21[366], line_20[364], line_19[362], line_18[360], line_17[358], line_16[356], line_15[354], line_14[352], line_13[350], line_12[348], line_11[346], line_10[344], line_9[342], line_8[340], line_7[338], line_6[336], line_5[334], line_4[332], line_3[330], line_2[328], line_1[326] };
assign col_581 = {line_128[581], line_127[579], line_126[577], line_125[575], line_124[573], line_123[571], line_122[569], line_121[567], line_120[565], line_119[563], line_118[561], line_117[559], line_116[557], line_115[555], line_114[553], line_113[551], line_112[549], line_111[547], line_110[545], line_109[543], line_108[541], line_107[539], line_106[537], line_105[535], line_104[533], line_103[531], line_102[529], line_101[527], line_100[525], line_99[523], line_98[521], line_97[519], line_96[517], line_95[515], line_94[513], line_93[511], line_92[509], line_91[507], line_90[505], line_89[503], line_88[501], line_87[499], line_86[497], line_85[495], line_84[493], line_83[491], line_82[489], line_81[487], line_80[485], line_79[483], line_78[481], line_77[479], line_76[477], line_75[475], line_74[473], line_73[471], line_72[469], line_71[467], line_70[465], line_69[463], line_68[461], line_67[459], line_66[457], line_65[455], line_64[453], line_63[451], line_62[449], line_61[447], line_60[445], line_59[443], line_58[441], line_57[439], line_56[437], line_55[435], line_54[433], line_53[431], line_52[429], line_51[427], line_50[425], line_49[423], line_48[421], line_47[419], line_46[417], line_45[415], line_44[413], line_43[411], line_42[409], line_41[407], line_40[405], line_39[403], line_38[401], line_37[399], line_36[397], line_35[395], line_34[393], line_33[391], line_32[389], line_31[387], line_30[385], line_29[383], line_28[381], line_27[379], line_26[377], line_25[375], line_24[373], line_23[371], line_22[369], line_21[367], line_20[365], line_19[363], line_18[361], line_17[359], line_16[357], line_15[355], line_14[353], line_13[351], line_12[349], line_11[347], line_10[345], line_9[343], line_8[341], line_7[339], line_6[337], line_5[335], line_4[333], line_3[331], line_2[329], line_1[327] };
assign col_582 = {line_128[582], line_127[580], line_126[578], line_125[576], line_124[574], line_123[572], line_122[570], line_121[568], line_120[566], line_119[564], line_118[562], line_117[560], line_116[558], line_115[556], line_114[554], line_113[552], line_112[550], line_111[548], line_110[546], line_109[544], line_108[542], line_107[540], line_106[538], line_105[536], line_104[534], line_103[532], line_102[530], line_101[528], line_100[526], line_99[524], line_98[522], line_97[520], line_96[518], line_95[516], line_94[514], line_93[512], line_92[510], line_91[508], line_90[506], line_89[504], line_88[502], line_87[500], line_86[498], line_85[496], line_84[494], line_83[492], line_82[490], line_81[488], line_80[486], line_79[484], line_78[482], line_77[480], line_76[478], line_75[476], line_74[474], line_73[472], line_72[470], line_71[468], line_70[466], line_69[464], line_68[462], line_67[460], line_66[458], line_65[456], line_64[454], line_63[452], line_62[450], line_61[448], line_60[446], line_59[444], line_58[442], line_57[440], line_56[438], line_55[436], line_54[434], line_53[432], line_52[430], line_51[428], line_50[426], line_49[424], line_48[422], line_47[420], line_46[418], line_45[416], line_44[414], line_43[412], line_42[410], line_41[408], line_40[406], line_39[404], line_38[402], line_37[400], line_36[398], line_35[396], line_34[394], line_33[392], line_32[390], line_31[388], line_30[386], line_29[384], line_28[382], line_27[380], line_26[378], line_25[376], line_24[374], line_23[372], line_22[370], line_21[368], line_20[366], line_19[364], line_18[362], line_17[360], line_16[358], line_15[356], line_14[354], line_13[352], line_12[350], line_11[348], line_10[346], line_9[344], line_8[342], line_7[340], line_6[338], line_5[336], line_4[334], line_3[332], line_2[330], line_1[328] };
assign col_583 = {line_128[583], line_127[581], line_126[579], line_125[577], line_124[575], line_123[573], line_122[571], line_121[569], line_120[567], line_119[565], line_118[563], line_117[561], line_116[559], line_115[557], line_114[555], line_113[553], line_112[551], line_111[549], line_110[547], line_109[545], line_108[543], line_107[541], line_106[539], line_105[537], line_104[535], line_103[533], line_102[531], line_101[529], line_100[527], line_99[525], line_98[523], line_97[521], line_96[519], line_95[517], line_94[515], line_93[513], line_92[511], line_91[509], line_90[507], line_89[505], line_88[503], line_87[501], line_86[499], line_85[497], line_84[495], line_83[493], line_82[491], line_81[489], line_80[487], line_79[485], line_78[483], line_77[481], line_76[479], line_75[477], line_74[475], line_73[473], line_72[471], line_71[469], line_70[467], line_69[465], line_68[463], line_67[461], line_66[459], line_65[457], line_64[455], line_63[453], line_62[451], line_61[449], line_60[447], line_59[445], line_58[443], line_57[441], line_56[439], line_55[437], line_54[435], line_53[433], line_52[431], line_51[429], line_50[427], line_49[425], line_48[423], line_47[421], line_46[419], line_45[417], line_44[415], line_43[413], line_42[411], line_41[409], line_40[407], line_39[405], line_38[403], line_37[401], line_36[399], line_35[397], line_34[395], line_33[393], line_32[391], line_31[389], line_30[387], line_29[385], line_28[383], line_27[381], line_26[379], line_25[377], line_24[375], line_23[373], line_22[371], line_21[369], line_20[367], line_19[365], line_18[363], line_17[361], line_16[359], line_15[357], line_14[355], line_13[353], line_12[351], line_11[349], line_10[347], line_9[345], line_8[343], line_7[341], line_6[339], line_5[337], line_4[335], line_3[333], line_2[331], line_1[329] };
assign col_584 = {line_128[584], line_127[582], line_126[580], line_125[578], line_124[576], line_123[574], line_122[572], line_121[570], line_120[568], line_119[566], line_118[564], line_117[562], line_116[560], line_115[558], line_114[556], line_113[554], line_112[552], line_111[550], line_110[548], line_109[546], line_108[544], line_107[542], line_106[540], line_105[538], line_104[536], line_103[534], line_102[532], line_101[530], line_100[528], line_99[526], line_98[524], line_97[522], line_96[520], line_95[518], line_94[516], line_93[514], line_92[512], line_91[510], line_90[508], line_89[506], line_88[504], line_87[502], line_86[500], line_85[498], line_84[496], line_83[494], line_82[492], line_81[490], line_80[488], line_79[486], line_78[484], line_77[482], line_76[480], line_75[478], line_74[476], line_73[474], line_72[472], line_71[470], line_70[468], line_69[466], line_68[464], line_67[462], line_66[460], line_65[458], line_64[456], line_63[454], line_62[452], line_61[450], line_60[448], line_59[446], line_58[444], line_57[442], line_56[440], line_55[438], line_54[436], line_53[434], line_52[432], line_51[430], line_50[428], line_49[426], line_48[424], line_47[422], line_46[420], line_45[418], line_44[416], line_43[414], line_42[412], line_41[410], line_40[408], line_39[406], line_38[404], line_37[402], line_36[400], line_35[398], line_34[396], line_33[394], line_32[392], line_31[390], line_30[388], line_29[386], line_28[384], line_27[382], line_26[380], line_25[378], line_24[376], line_23[374], line_22[372], line_21[370], line_20[368], line_19[366], line_18[364], line_17[362], line_16[360], line_15[358], line_14[356], line_13[354], line_12[352], line_11[350], line_10[348], line_9[346], line_8[344], line_7[342], line_6[340], line_5[338], line_4[336], line_3[334], line_2[332], line_1[330] };
assign col_585 = {line_128[585], line_127[583], line_126[581], line_125[579], line_124[577], line_123[575], line_122[573], line_121[571], line_120[569], line_119[567], line_118[565], line_117[563], line_116[561], line_115[559], line_114[557], line_113[555], line_112[553], line_111[551], line_110[549], line_109[547], line_108[545], line_107[543], line_106[541], line_105[539], line_104[537], line_103[535], line_102[533], line_101[531], line_100[529], line_99[527], line_98[525], line_97[523], line_96[521], line_95[519], line_94[517], line_93[515], line_92[513], line_91[511], line_90[509], line_89[507], line_88[505], line_87[503], line_86[501], line_85[499], line_84[497], line_83[495], line_82[493], line_81[491], line_80[489], line_79[487], line_78[485], line_77[483], line_76[481], line_75[479], line_74[477], line_73[475], line_72[473], line_71[471], line_70[469], line_69[467], line_68[465], line_67[463], line_66[461], line_65[459], line_64[457], line_63[455], line_62[453], line_61[451], line_60[449], line_59[447], line_58[445], line_57[443], line_56[441], line_55[439], line_54[437], line_53[435], line_52[433], line_51[431], line_50[429], line_49[427], line_48[425], line_47[423], line_46[421], line_45[419], line_44[417], line_43[415], line_42[413], line_41[411], line_40[409], line_39[407], line_38[405], line_37[403], line_36[401], line_35[399], line_34[397], line_33[395], line_32[393], line_31[391], line_30[389], line_29[387], line_28[385], line_27[383], line_26[381], line_25[379], line_24[377], line_23[375], line_22[373], line_21[371], line_20[369], line_19[367], line_18[365], line_17[363], line_16[361], line_15[359], line_14[357], line_13[355], line_12[353], line_11[351], line_10[349], line_9[347], line_8[345], line_7[343], line_6[341], line_5[339], line_4[337], line_3[335], line_2[333], line_1[331] };
assign col_586 = {line_128[586], line_127[584], line_126[582], line_125[580], line_124[578], line_123[576], line_122[574], line_121[572], line_120[570], line_119[568], line_118[566], line_117[564], line_116[562], line_115[560], line_114[558], line_113[556], line_112[554], line_111[552], line_110[550], line_109[548], line_108[546], line_107[544], line_106[542], line_105[540], line_104[538], line_103[536], line_102[534], line_101[532], line_100[530], line_99[528], line_98[526], line_97[524], line_96[522], line_95[520], line_94[518], line_93[516], line_92[514], line_91[512], line_90[510], line_89[508], line_88[506], line_87[504], line_86[502], line_85[500], line_84[498], line_83[496], line_82[494], line_81[492], line_80[490], line_79[488], line_78[486], line_77[484], line_76[482], line_75[480], line_74[478], line_73[476], line_72[474], line_71[472], line_70[470], line_69[468], line_68[466], line_67[464], line_66[462], line_65[460], line_64[458], line_63[456], line_62[454], line_61[452], line_60[450], line_59[448], line_58[446], line_57[444], line_56[442], line_55[440], line_54[438], line_53[436], line_52[434], line_51[432], line_50[430], line_49[428], line_48[426], line_47[424], line_46[422], line_45[420], line_44[418], line_43[416], line_42[414], line_41[412], line_40[410], line_39[408], line_38[406], line_37[404], line_36[402], line_35[400], line_34[398], line_33[396], line_32[394], line_31[392], line_30[390], line_29[388], line_28[386], line_27[384], line_26[382], line_25[380], line_24[378], line_23[376], line_22[374], line_21[372], line_20[370], line_19[368], line_18[366], line_17[364], line_16[362], line_15[360], line_14[358], line_13[356], line_12[354], line_11[352], line_10[350], line_9[348], line_8[346], line_7[344], line_6[342], line_5[340], line_4[338], line_3[336], line_2[334], line_1[332] };
assign col_587 = {line_128[587], line_127[585], line_126[583], line_125[581], line_124[579], line_123[577], line_122[575], line_121[573], line_120[571], line_119[569], line_118[567], line_117[565], line_116[563], line_115[561], line_114[559], line_113[557], line_112[555], line_111[553], line_110[551], line_109[549], line_108[547], line_107[545], line_106[543], line_105[541], line_104[539], line_103[537], line_102[535], line_101[533], line_100[531], line_99[529], line_98[527], line_97[525], line_96[523], line_95[521], line_94[519], line_93[517], line_92[515], line_91[513], line_90[511], line_89[509], line_88[507], line_87[505], line_86[503], line_85[501], line_84[499], line_83[497], line_82[495], line_81[493], line_80[491], line_79[489], line_78[487], line_77[485], line_76[483], line_75[481], line_74[479], line_73[477], line_72[475], line_71[473], line_70[471], line_69[469], line_68[467], line_67[465], line_66[463], line_65[461], line_64[459], line_63[457], line_62[455], line_61[453], line_60[451], line_59[449], line_58[447], line_57[445], line_56[443], line_55[441], line_54[439], line_53[437], line_52[435], line_51[433], line_50[431], line_49[429], line_48[427], line_47[425], line_46[423], line_45[421], line_44[419], line_43[417], line_42[415], line_41[413], line_40[411], line_39[409], line_38[407], line_37[405], line_36[403], line_35[401], line_34[399], line_33[397], line_32[395], line_31[393], line_30[391], line_29[389], line_28[387], line_27[385], line_26[383], line_25[381], line_24[379], line_23[377], line_22[375], line_21[373], line_20[371], line_19[369], line_18[367], line_17[365], line_16[363], line_15[361], line_14[359], line_13[357], line_12[355], line_11[353], line_10[351], line_9[349], line_8[347], line_7[345], line_6[343], line_5[341], line_4[339], line_3[337], line_2[335], line_1[333] };
assign col_588 = {line_128[588], line_127[586], line_126[584], line_125[582], line_124[580], line_123[578], line_122[576], line_121[574], line_120[572], line_119[570], line_118[568], line_117[566], line_116[564], line_115[562], line_114[560], line_113[558], line_112[556], line_111[554], line_110[552], line_109[550], line_108[548], line_107[546], line_106[544], line_105[542], line_104[540], line_103[538], line_102[536], line_101[534], line_100[532], line_99[530], line_98[528], line_97[526], line_96[524], line_95[522], line_94[520], line_93[518], line_92[516], line_91[514], line_90[512], line_89[510], line_88[508], line_87[506], line_86[504], line_85[502], line_84[500], line_83[498], line_82[496], line_81[494], line_80[492], line_79[490], line_78[488], line_77[486], line_76[484], line_75[482], line_74[480], line_73[478], line_72[476], line_71[474], line_70[472], line_69[470], line_68[468], line_67[466], line_66[464], line_65[462], line_64[460], line_63[458], line_62[456], line_61[454], line_60[452], line_59[450], line_58[448], line_57[446], line_56[444], line_55[442], line_54[440], line_53[438], line_52[436], line_51[434], line_50[432], line_49[430], line_48[428], line_47[426], line_46[424], line_45[422], line_44[420], line_43[418], line_42[416], line_41[414], line_40[412], line_39[410], line_38[408], line_37[406], line_36[404], line_35[402], line_34[400], line_33[398], line_32[396], line_31[394], line_30[392], line_29[390], line_28[388], line_27[386], line_26[384], line_25[382], line_24[380], line_23[378], line_22[376], line_21[374], line_20[372], line_19[370], line_18[368], line_17[366], line_16[364], line_15[362], line_14[360], line_13[358], line_12[356], line_11[354], line_10[352], line_9[350], line_8[348], line_7[346], line_6[344], line_5[342], line_4[340], line_3[338], line_2[336], line_1[334] };
assign col_589 = {line_128[589], line_127[587], line_126[585], line_125[583], line_124[581], line_123[579], line_122[577], line_121[575], line_120[573], line_119[571], line_118[569], line_117[567], line_116[565], line_115[563], line_114[561], line_113[559], line_112[557], line_111[555], line_110[553], line_109[551], line_108[549], line_107[547], line_106[545], line_105[543], line_104[541], line_103[539], line_102[537], line_101[535], line_100[533], line_99[531], line_98[529], line_97[527], line_96[525], line_95[523], line_94[521], line_93[519], line_92[517], line_91[515], line_90[513], line_89[511], line_88[509], line_87[507], line_86[505], line_85[503], line_84[501], line_83[499], line_82[497], line_81[495], line_80[493], line_79[491], line_78[489], line_77[487], line_76[485], line_75[483], line_74[481], line_73[479], line_72[477], line_71[475], line_70[473], line_69[471], line_68[469], line_67[467], line_66[465], line_65[463], line_64[461], line_63[459], line_62[457], line_61[455], line_60[453], line_59[451], line_58[449], line_57[447], line_56[445], line_55[443], line_54[441], line_53[439], line_52[437], line_51[435], line_50[433], line_49[431], line_48[429], line_47[427], line_46[425], line_45[423], line_44[421], line_43[419], line_42[417], line_41[415], line_40[413], line_39[411], line_38[409], line_37[407], line_36[405], line_35[403], line_34[401], line_33[399], line_32[397], line_31[395], line_30[393], line_29[391], line_28[389], line_27[387], line_26[385], line_25[383], line_24[381], line_23[379], line_22[377], line_21[375], line_20[373], line_19[371], line_18[369], line_17[367], line_16[365], line_15[363], line_14[361], line_13[359], line_12[357], line_11[355], line_10[353], line_9[351], line_8[349], line_7[347], line_6[345], line_5[343], line_4[341], line_3[339], line_2[337], line_1[335] };
assign col_590 = {line_128[590], line_127[588], line_126[586], line_125[584], line_124[582], line_123[580], line_122[578], line_121[576], line_120[574], line_119[572], line_118[570], line_117[568], line_116[566], line_115[564], line_114[562], line_113[560], line_112[558], line_111[556], line_110[554], line_109[552], line_108[550], line_107[548], line_106[546], line_105[544], line_104[542], line_103[540], line_102[538], line_101[536], line_100[534], line_99[532], line_98[530], line_97[528], line_96[526], line_95[524], line_94[522], line_93[520], line_92[518], line_91[516], line_90[514], line_89[512], line_88[510], line_87[508], line_86[506], line_85[504], line_84[502], line_83[500], line_82[498], line_81[496], line_80[494], line_79[492], line_78[490], line_77[488], line_76[486], line_75[484], line_74[482], line_73[480], line_72[478], line_71[476], line_70[474], line_69[472], line_68[470], line_67[468], line_66[466], line_65[464], line_64[462], line_63[460], line_62[458], line_61[456], line_60[454], line_59[452], line_58[450], line_57[448], line_56[446], line_55[444], line_54[442], line_53[440], line_52[438], line_51[436], line_50[434], line_49[432], line_48[430], line_47[428], line_46[426], line_45[424], line_44[422], line_43[420], line_42[418], line_41[416], line_40[414], line_39[412], line_38[410], line_37[408], line_36[406], line_35[404], line_34[402], line_33[400], line_32[398], line_31[396], line_30[394], line_29[392], line_28[390], line_27[388], line_26[386], line_25[384], line_24[382], line_23[380], line_22[378], line_21[376], line_20[374], line_19[372], line_18[370], line_17[368], line_16[366], line_15[364], line_14[362], line_13[360], line_12[358], line_11[356], line_10[354], line_9[352], line_8[350], line_7[348], line_6[346], line_5[344], line_4[342], line_3[340], line_2[338], line_1[336] };
assign col_591 = {line_128[591], line_127[589], line_126[587], line_125[585], line_124[583], line_123[581], line_122[579], line_121[577], line_120[575], line_119[573], line_118[571], line_117[569], line_116[567], line_115[565], line_114[563], line_113[561], line_112[559], line_111[557], line_110[555], line_109[553], line_108[551], line_107[549], line_106[547], line_105[545], line_104[543], line_103[541], line_102[539], line_101[537], line_100[535], line_99[533], line_98[531], line_97[529], line_96[527], line_95[525], line_94[523], line_93[521], line_92[519], line_91[517], line_90[515], line_89[513], line_88[511], line_87[509], line_86[507], line_85[505], line_84[503], line_83[501], line_82[499], line_81[497], line_80[495], line_79[493], line_78[491], line_77[489], line_76[487], line_75[485], line_74[483], line_73[481], line_72[479], line_71[477], line_70[475], line_69[473], line_68[471], line_67[469], line_66[467], line_65[465], line_64[463], line_63[461], line_62[459], line_61[457], line_60[455], line_59[453], line_58[451], line_57[449], line_56[447], line_55[445], line_54[443], line_53[441], line_52[439], line_51[437], line_50[435], line_49[433], line_48[431], line_47[429], line_46[427], line_45[425], line_44[423], line_43[421], line_42[419], line_41[417], line_40[415], line_39[413], line_38[411], line_37[409], line_36[407], line_35[405], line_34[403], line_33[401], line_32[399], line_31[397], line_30[395], line_29[393], line_28[391], line_27[389], line_26[387], line_25[385], line_24[383], line_23[381], line_22[379], line_21[377], line_20[375], line_19[373], line_18[371], line_17[369], line_16[367], line_15[365], line_14[363], line_13[361], line_12[359], line_11[357], line_10[355], line_9[353], line_8[351], line_7[349], line_6[347], line_5[345], line_4[343], line_3[341], line_2[339], line_1[337] };
assign col_592 = {line_128[592], line_127[590], line_126[588], line_125[586], line_124[584], line_123[582], line_122[580], line_121[578], line_120[576], line_119[574], line_118[572], line_117[570], line_116[568], line_115[566], line_114[564], line_113[562], line_112[560], line_111[558], line_110[556], line_109[554], line_108[552], line_107[550], line_106[548], line_105[546], line_104[544], line_103[542], line_102[540], line_101[538], line_100[536], line_99[534], line_98[532], line_97[530], line_96[528], line_95[526], line_94[524], line_93[522], line_92[520], line_91[518], line_90[516], line_89[514], line_88[512], line_87[510], line_86[508], line_85[506], line_84[504], line_83[502], line_82[500], line_81[498], line_80[496], line_79[494], line_78[492], line_77[490], line_76[488], line_75[486], line_74[484], line_73[482], line_72[480], line_71[478], line_70[476], line_69[474], line_68[472], line_67[470], line_66[468], line_65[466], line_64[464], line_63[462], line_62[460], line_61[458], line_60[456], line_59[454], line_58[452], line_57[450], line_56[448], line_55[446], line_54[444], line_53[442], line_52[440], line_51[438], line_50[436], line_49[434], line_48[432], line_47[430], line_46[428], line_45[426], line_44[424], line_43[422], line_42[420], line_41[418], line_40[416], line_39[414], line_38[412], line_37[410], line_36[408], line_35[406], line_34[404], line_33[402], line_32[400], line_31[398], line_30[396], line_29[394], line_28[392], line_27[390], line_26[388], line_25[386], line_24[384], line_23[382], line_22[380], line_21[378], line_20[376], line_19[374], line_18[372], line_17[370], line_16[368], line_15[366], line_14[364], line_13[362], line_12[360], line_11[358], line_10[356], line_9[354], line_8[352], line_7[350], line_6[348], line_5[346], line_4[344], line_3[342], line_2[340], line_1[338] };
assign col_593 = {line_128[593], line_127[591], line_126[589], line_125[587], line_124[585], line_123[583], line_122[581], line_121[579], line_120[577], line_119[575], line_118[573], line_117[571], line_116[569], line_115[567], line_114[565], line_113[563], line_112[561], line_111[559], line_110[557], line_109[555], line_108[553], line_107[551], line_106[549], line_105[547], line_104[545], line_103[543], line_102[541], line_101[539], line_100[537], line_99[535], line_98[533], line_97[531], line_96[529], line_95[527], line_94[525], line_93[523], line_92[521], line_91[519], line_90[517], line_89[515], line_88[513], line_87[511], line_86[509], line_85[507], line_84[505], line_83[503], line_82[501], line_81[499], line_80[497], line_79[495], line_78[493], line_77[491], line_76[489], line_75[487], line_74[485], line_73[483], line_72[481], line_71[479], line_70[477], line_69[475], line_68[473], line_67[471], line_66[469], line_65[467], line_64[465], line_63[463], line_62[461], line_61[459], line_60[457], line_59[455], line_58[453], line_57[451], line_56[449], line_55[447], line_54[445], line_53[443], line_52[441], line_51[439], line_50[437], line_49[435], line_48[433], line_47[431], line_46[429], line_45[427], line_44[425], line_43[423], line_42[421], line_41[419], line_40[417], line_39[415], line_38[413], line_37[411], line_36[409], line_35[407], line_34[405], line_33[403], line_32[401], line_31[399], line_30[397], line_29[395], line_28[393], line_27[391], line_26[389], line_25[387], line_24[385], line_23[383], line_22[381], line_21[379], line_20[377], line_19[375], line_18[373], line_17[371], line_16[369], line_15[367], line_14[365], line_13[363], line_12[361], line_11[359], line_10[357], line_9[355], line_8[353], line_7[351], line_6[349], line_5[347], line_4[345], line_3[343], line_2[341], line_1[339] };
assign col_594 = {line_128[594], line_127[592], line_126[590], line_125[588], line_124[586], line_123[584], line_122[582], line_121[580], line_120[578], line_119[576], line_118[574], line_117[572], line_116[570], line_115[568], line_114[566], line_113[564], line_112[562], line_111[560], line_110[558], line_109[556], line_108[554], line_107[552], line_106[550], line_105[548], line_104[546], line_103[544], line_102[542], line_101[540], line_100[538], line_99[536], line_98[534], line_97[532], line_96[530], line_95[528], line_94[526], line_93[524], line_92[522], line_91[520], line_90[518], line_89[516], line_88[514], line_87[512], line_86[510], line_85[508], line_84[506], line_83[504], line_82[502], line_81[500], line_80[498], line_79[496], line_78[494], line_77[492], line_76[490], line_75[488], line_74[486], line_73[484], line_72[482], line_71[480], line_70[478], line_69[476], line_68[474], line_67[472], line_66[470], line_65[468], line_64[466], line_63[464], line_62[462], line_61[460], line_60[458], line_59[456], line_58[454], line_57[452], line_56[450], line_55[448], line_54[446], line_53[444], line_52[442], line_51[440], line_50[438], line_49[436], line_48[434], line_47[432], line_46[430], line_45[428], line_44[426], line_43[424], line_42[422], line_41[420], line_40[418], line_39[416], line_38[414], line_37[412], line_36[410], line_35[408], line_34[406], line_33[404], line_32[402], line_31[400], line_30[398], line_29[396], line_28[394], line_27[392], line_26[390], line_25[388], line_24[386], line_23[384], line_22[382], line_21[380], line_20[378], line_19[376], line_18[374], line_17[372], line_16[370], line_15[368], line_14[366], line_13[364], line_12[362], line_11[360], line_10[358], line_9[356], line_8[354], line_7[352], line_6[350], line_5[348], line_4[346], line_3[344], line_2[342], line_1[340] };
assign col_595 = {line_128[595], line_127[593], line_126[591], line_125[589], line_124[587], line_123[585], line_122[583], line_121[581], line_120[579], line_119[577], line_118[575], line_117[573], line_116[571], line_115[569], line_114[567], line_113[565], line_112[563], line_111[561], line_110[559], line_109[557], line_108[555], line_107[553], line_106[551], line_105[549], line_104[547], line_103[545], line_102[543], line_101[541], line_100[539], line_99[537], line_98[535], line_97[533], line_96[531], line_95[529], line_94[527], line_93[525], line_92[523], line_91[521], line_90[519], line_89[517], line_88[515], line_87[513], line_86[511], line_85[509], line_84[507], line_83[505], line_82[503], line_81[501], line_80[499], line_79[497], line_78[495], line_77[493], line_76[491], line_75[489], line_74[487], line_73[485], line_72[483], line_71[481], line_70[479], line_69[477], line_68[475], line_67[473], line_66[471], line_65[469], line_64[467], line_63[465], line_62[463], line_61[461], line_60[459], line_59[457], line_58[455], line_57[453], line_56[451], line_55[449], line_54[447], line_53[445], line_52[443], line_51[441], line_50[439], line_49[437], line_48[435], line_47[433], line_46[431], line_45[429], line_44[427], line_43[425], line_42[423], line_41[421], line_40[419], line_39[417], line_38[415], line_37[413], line_36[411], line_35[409], line_34[407], line_33[405], line_32[403], line_31[401], line_30[399], line_29[397], line_28[395], line_27[393], line_26[391], line_25[389], line_24[387], line_23[385], line_22[383], line_21[381], line_20[379], line_19[377], line_18[375], line_17[373], line_16[371], line_15[369], line_14[367], line_13[365], line_12[363], line_11[361], line_10[359], line_9[357], line_8[355], line_7[353], line_6[351], line_5[349], line_4[347], line_3[345], line_2[343], line_1[341] };
assign col_596 = {line_128[596], line_127[594], line_126[592], line_125[590], line_124[588], line_123[586], line_122[584], line_121[582], line_120[580], line_119[578], line_118[576], line_117[574], line_116[572], line_115[570], line_114[568], line_113[566], line_112[564], line_111[562], line_110[560], line_109[558], line_108[556], line_107[554], line_106[552], line_105[550], line_104[548], line_103[546], line_102[544], line_101[542], line_100[540], line_99[538], line_98[536], line_97[534], line_96[532], line_95[530], line_94[528], line_93[526], line_92[524], line_91[522], line_90[520], line_89[518], line_88[516], line_87[514], line_86[512], line_85[510], line_84[508], line_83[506], line_82[504], line_81[502], line_80[500], line_79[498], line_78[496], line_77[494], line_76[492], line_75[490], line_74[488], line_73[486], line_72[484], line_71[482], line_70[480], line_69[478], line_68[476], line_67[474], line_66[472], line_65[470], line_64[468], line_63[466], line_62[464], line_61[462], line_60[460], line_59[458], line_58[456], line_57[454], line_56[452], line_55[450], line_54[448], line_53[446], line_52[444], line_51[442], line_50[440], line_49[438], line_48[436], line_47[434], line_46[432], line_45[430], line_44[428], line_43[426], line_42[424], line_41[422], line_40[420], line_39[418], line_38[416], line_37[414], line_36[412], line_35[410], line_34[408], line_33[406], line_32[404], line_31[402], line_30[400], line_29[398], line_28[396], line_27[394], line_26[392], line_25[390], line_24[388], line_23[386], line_22[384], line_21[382], line_20[380], line_19[378], line_18[376], line_17[374], line_16[372], line_15[370], line_14[368], line_13[366], line_12[364], line_11[362], line_10[360], line_9[358], line_8[356], line_7[354], line_6[352], line_5[350], line_4[348], line_3[346], line_2[344], line_1[342] };
assign col_597 = {line_128[597], line_127[595], line_126[593], line_125[591], line_124[589], line_123[587], line_122[585], line_121[583], line_120[581], line_119[579], line_118[577], line_117[575], line_116[573], line_115[571], line_114[569], line_113[567], line_112[565], line_111[563], line_110[561], line_109[559], line_108[557], line_107[555], line_106[553], line_105[551], line_104[549], line_103[547], line_102[545], line_101[543], line_100[541], line_99[539], line_98[537], line_97[535], line_96[533], line_95[531], line_94[529], line_93[527], line_92[525], line_91[523], line_90[521], line_89[519], line_88[517], line_87[515], line_86[513], line_85[511], line_84[509], line_83[507], line_82[505], line_81[503], line_80[501], line_79[499], line_78[497], line_77[495], line_76[493], line_75[491], line_74[489], line_73[487], line_72[485], line_71[483], line_70[481], line_69[479], line_68[477], line_67[475], line_66[473], line_65[471], line_64[469], line_63[467], line_62[465], line_61[463], line_60[461], line_59[459], line_58[457], line_57[455], line_56[453], line_55[451], line_54[449], line_53[447], line_52[445], line_51[443], line_50[441], line_49[439], line_48[437], line_47[435], line_46[433], line_45[431], line_44[429], line_43[427], line_42[425], line_41[423], line_40[421], line_39[419], line_38[417], line_37[415], line_36[413], line_35[411], line_34[409], line_33[407], line_32[405], line_31[403], line_30[401], line_29[399], line_28[397], line_27[395], line_26[393], line_25[391], line_24[389], line_23[387], line_22[385], line_21[383], line_20[381], line_19[379], line_18[377], line_17[375], line_16[373], line_15[371], line_14[369], line_13[367], line_12[365], line_11[363], line_10[361], line_9[359], line_8[357], line_7[355], line_6[353], line_5[351], line_4[349], line_3[347], line_2[345], line_1[343] };
assign col_598 = {line_128[598], line_127[596], line_126[594], line_125[592], line_124[590], line_123[588], line_122[586], line_121[584], line_120[582], line_119[580], line_118[578], line_117[576], line_116[574], line_115[572], line_114[570], line_113[568], line_112[566], line_111[564], line_110[562], line_109[560], line_108[558], line_107[556], line_106[554], line_105[552], line_104[550], line_103[548], line_102[546], line_101[544], line_100[542], line_99[540], line_98[538], line_97[536], line_96[534], line_95[532], line_94[530], line_93[528], line_92[526], line_91[524], line_90[522], line_89[520], line_88[518], line_87[516], line_86[514], line_85[512], line_84[510], line_83[508], line_82[506], line_81[504], line_80[502], line_79[500], line_78[498], line_77[496], line_76[494], line_75[492], line_74[490], line_73[488], line_72[486], line_71[484], line_70[482], line_69[480], line_68[478], line_67[476], line_66[474], line_65[472], line_64[470], line_63[468], line_62[466], line_61[464], line_60[462], line_59[460], line_58[458], line_57[456], line_56[454], line_55[452], line_54[450], line_53[448], line_52[446], line_51[444], line_50[442], line_49[440], line_48[438], line_47[436], line_46[434], line_45[432], line_44[430], line_43[428], line_42[426], line_41[424], line_40[422], line_39[420], line_38[418], line_37[416], line_36[414], line_35[412], line_34[410], line_33[408], line_32[406], line_31[404], line_30[402], line_29[400], line_28[398], line_27[396], line_26[394], line_25[392], line_24[390], line_23[388], line_22[386], line_21[384], line_20[382], line_19[380], line_18[378], line_17[376], line_16[374], line_15[372], line_14[370], line_13[368], line_12[366], line_11[364], line_10[362], line_9[360], line_8[358], line_7[356], line_6[354], line_5[352], line_4[350], line_3[348], line_2[346], line_1[344] };
assign col_599 = {line_128[599], line_127[597], line_126[595], line_125[593], line_124[591], line_123[589], line_122[587], line_121[585], line_120[583], line_119[581], line_118[579], line_117[577], line_116[575], line_115[573], line_114[571], line_113[569], line_112[567], line_111[565], line_110[563], line_109[561], line_108[559], line_107[557], line_106[555], line_105[553], line_104[551], line_103[549], line_102[547], line_101[545], line_100[543], line_99[541], line_98[539], line_97[537], line_96[535], line_95[533], line_94[531], line_93[529], line_92[527], line_91[525], line_90[523], line_89[521], line_88[519], line_87[517], line_86[515], line_85[513], line_84[511], line_83[509], line_82[507], line_81[505], line_80[503], line_79[501], line_78[499], line_77[497], line_76[495], line_75[493], line_74[491], line_73[489], line_72[487], line_71[485], line_70[483], line_69[481], line_68[479], line_67[477], line_66[475], line_65[473], line_64[471], line_63[469], line_62[467], line_61[465], line_60[463], line_59[461], line_58[459], line_57[457], line_56[455], line_55[453], line_54[451], line_53[449], line_52[447], line_51[445], line_50[443], line_49[441], line_48[439], line_47[437], line_46[435], line_45[433], line_44[431], line_43[429], line_42[427], line_41[425], line_40[423], line_39[421], line_38[419], line_37[417], line_36[415], line_35[413], line_34[411], line_33[409], line_32[407], line_31[405], line_30[403], line_29[401], line_28[399], line_27[397], line_26[395], line_25[393], line_24[391], line_23[389], line_22[387], line_21[385], line_20[383], line_19[381], line_18[379], line_17[377], line_16[375], line_15[373], line_14[371], line_13[369], line_12[367], line_11[365], line_10[363], line_9[361], line_8[359], line_7[357], line_6[355], line_5[353], line_4[351], line_3[349], line_2[347], line_1[345] };
assign col_600 = {line_128[600], line_127[598], line_126[596], line_125[594], line_124[592], line_123[590], line_122[588], line_121[586], line_120[584], line_119[582], line_118[580], line_117[578], line_116[576], line_115[574], line_114[572], line_113[570], line_112[568], line_111[566], line_110[564], line_109[562], line_108[560], line_107[558], line_106[556], line_105[554], line_104[552], line_103[550], line_102[548], line_101[546], line_100[544], line_99[542], line_98[540], line_97[538], line_96[536], line_95[534], line_94[532], line_93[530], line_92[528], line_91[526], line_90[524], line_89[522], line_88[520], line_87[518], line_86[516], line_85[514], line_84[512], line_83[510], line_82[508], line_81[506], line_80[504], line_79[502], line_78[500], line_77[498], line_76[496], line_75[494], line_74[492], line_73[490], line_72[488], line_71[486], line_70[484], line_69[482], line_68[480], line_67[478], line_66[476], line_65[474], line_64[472], line_63[470], line_62[468], line_61[466], line_60[464], line_59[462], line_58[460], line_57[458], line_56[456], line_55[454], line_54[452], line_53[450], line_52[448], line_51[446], line_50[444], line_49[442], line_48[440], line_47[438], line_46[436], line_45[434], line_44[432], line_43[430], line_42[428], line_41[426], line_40[424], line_39[422], line_38[420], line_37[418], line_36[416], line_35[414], line_34[412], line_33[410], line_32[408], line_31[406], line_30[404], line_29[402], line_28[400], line_27[398], line_26[396], line_25[394], line_24[392], line_23[390], line_22[388], line_21[386], line_20[384], line_19[382], line_18[380], line_17[378], line_16[376], line_15[374], line_14[372], line_13[370], line_12[368], line_11[366], line_10[364], line_9[362], line_8[360], line_7[358], line_6[356], line_5[354], line_4[352], line_3[350], line_2[348], line_1[346] };
assign col_601 = {line_128[601], line_127[599], line_126[597], line_125[595], line_124[593], line_123[591], line_122[589], line_121[587], line_120[585], line_119[583], line_118[581], line_117[579], line_116[577], line_115[575], line_114[573], line_113[571], line_112[569], line_111[567], line_110[565], line_109[563], line_108[561], line_107[559], line_106[557], line_105[555], line_104[553], line_103[551], line_102[549], line_101[547], line_100[545], line_99[543], line_98[541], line_97[539], line_96[537], line_95[535], line_94[533], line_93[531], line_92[529], line_91[527], line_90[525], line_89[523], line_88[521], line_87[519], line_86[517], line_85[515], line_84[513], line_83[511], line_82[509], line_81[507], line_80[505], line_79[503], line_78[501], line_77[499], line_76[497], line_75[495], line_74[493], line_73[491], line_72[489], line_71[487], line_70[485], line_69[483], line_68[481], line_67[479], line_66[477], line_65[475], line_64[473], line_63[471], line_62[469], line_61[467], line_60[465], line_59[463], line_58[461], line_57[459], line_56[457], line_55[455], line_54[453], line_53[451], line_52[449], line_51[447], line_50[445], line_49[443], line_48[441], line_47[439], line_46[437], line_45[435], line_44[433], line_43[431], line_42[429], line_41[427], line_40[425], line_39[423], line_38[421], line_37[419], line_36[417], line_35[415], line_34[413], line_33[411], line_32[409], line_31[407], line_30[405], line_29[403], line_28[401], line_27[399], line_26[397], line_25[395], line_24[393], line_23[391], line_22[389], line_21[387], line_20[385], line_19[383], line_18[381], line_17[379], line_16[377], line_15[375], line_14[373], line_13[371], line_12[369], line_11[367], line_10[365], line_9[363], line_8[361], line_7[359], line_6[357], line_5[355], line_4[353], line_3[351], line_2[349], line_1[347] };
assign col_602 = {line_128[602], line_127[600], line_126[598], line_125[596], line_124[594], line_123[592], line_122[590], line_121[588], line_120[586], line_119[584], line_118[582], line_117[580], line_116[578], line_115[576], line_114[574], line_113[572], line_112[570], line_111[568], line_110[566], line_109[564], line_108[562], line_107[560], line_106[558], line_105[556], line_104[554], line_103[552], line_102[550], line_101[548], line_100[546], line_99[544], line_98[542], line_97[540], line_96[538], line_95[536], line_94[534], line_93[532], line_92[530], line_91[528], line_90[526], line_89[524], line_88[522], line_87[520], line_86[518], line_85[516], line_84[514], line_83[512], line_82[510], line_81[508], line_80[506], line_79[504], line_78[502], line_77[500], line_76[498], line_75[496], line_74[494], line_73[492], line_72[490], line_71[488], line_70[486], line_69[484], line_68[482], line_67[480], line_66[478], line_65[476], line_64[474], line_63[472], line_62[470], line_61[468], line_60[466], line_59[464], line_58[462], line_57[460], line_56[458], line_55[456], line_54[454], line_53[452], line_52[450], line_51[448], line_50[446], line_49[444], line_48[442], line_47[440], line_46[438], line_45[436], line_44[434], line_43[432], line_42[430], line_41[428], line_40[426], line_39[424], line_38[422], line_37[420], line_36[418], line_35[416], line_34[414], line_33[412], line_32[410], line_31[408], line_30[406], line_29[404], line_28[402], line_27[400], line_26[398], line_25[396], line_24[394], line_23[392], line_22[390], line_21[388], line_20[386], line_19[384], line_18[382], line_17[380], line_16[378], line_15[376], line_14[374], line_13[372], line_12[370], line_11[368], line_10[366], line_9[364], line_8[362], line_7[360], line_6[358], line_5[356], line_4[354], line_3[352], line_2[350], line_1[348] };
assign col_603 = {line_128[603], line_127[601], line_126[599], line_125[597], line_124[595], line_123[593], line_122[591], line_121[589], line_120[587], line_119[585], line_118[583], line_117[581], line_116[579], line_115[577], line_114[575], line_113[573], line_112[571], line_111[569], line_110[567], line_109[565], line_108[563], line_107[561], line_106[559], line_105[557], line_104[555], line_103[553], line_102[551], line_101[549], line_100[547], line_99[545], line_98[543], line_97[541], line_96[539], line_95[537], line_94[535], line_93[533], line_92[531], line_91[529], line_90[527], line_89[525], line_88[523], line_87[521], line_86[519], line_85[517], line_84[515], line_83[513], line_82[511], line_81[509], line_80[507], line_79[505], line_78[503], line_77[501], line_76[499], line_75[497], line_74[495], line_73[493], line_72[491], line_71[489], line_70[487], line_69[485], line_68[483], line_67[481], line_66[479], line_65[477], line_64[475], line_63[473], line_62[471], line_61[469], line_60[467], line_59[465], line_58[463], line_57[461], line_56[459], line_55[457], line_54[455], line_53[453], line_52[451], line_51[449], line_50[447], line_49[445], line_48[443], line_47[441], line_46[439], line_45[437], line_44[435], line_43[433], line_42[431], line_41[429], line_40[427], line_39[425], line_38[423], line_37[421], line_36[419], line_35[417], line_34[415], line_33[413], line_32[411], line_31[409], line_30[407], line_29[405], line_28[403], line_27[401], line_26[399], line_25[397], line_24[395], line_23[393], line_22[391], line_21[389], line_20[387], line_19[385], line_18[383], line_17[381], line_16[379], line_15[377], line_14[375], line_13[373], line_12[371], line_11[369], line_10[367], line_9[365], line_8[363], line_7[361], line_6[359], line_5[357], line_4[355], line_3[353], line_2[351], line_1[349] };
assign col_604 = {line_128[604], line_127[602], line_126[600], line_125[598], line_124[596], line_123[594], line_122[592], line_121[590], line_120[588], line_119[586], line_118[584], line_117[582], line_116[580], line_115[578], line_114[576], line_113[574], line_112[572], line_111[570], line_110[568], line_109[566], line_108[564], line_107[562], line_106[560], line_105[558], line_104[556], line_103[554], line_102[552], line_101[550], line_100[548], line_99[546], line_98[544], line_97[542], line_96[540], line_95[538], line_94[536], line_93[534], line_92[532], line_91[530], line_90[528], line_89[526], line_88[524], line_87[522], line_86[520], line_85[518], line_84[516], line_83[514], line_82[512], line_81[510], line_80[508], line_79[506], line_78[504], line_77[502], line_76[500], line_75[498], line_74[496], line_73[494], line_72[492], line_71[490], line_70[488], line_69[486], line_68[484], line_67[482], line_66[480], line_65[478], line_64[476], line_63[474], line_62[472], line_61[470], line_60[468], line_59[466], line_58[464], line_57[462], line_56[460], line_55[458], line_54[456], line_53[454], line_52[452], line_51[450], line_50[448], line_49[446], line_48[444], line_47[442], line_46[440], line_45[438], line_44[436], line_43[434], line_42[432], line_41[430], line_40[428], line_39[426], line_38[424], line_37[422], line_36[420], line_35[418], line_34[416], line_33[414], line_32[412], line_31[410], line_30[408], line_29[406], line_28[404], line_27[402], line_26[400], line_25[398], line_24[396], line_23[394], line_22[392], line_21[390], line_20[388], line_19[386], line_18[384], line_17[382], line_16[380], line_15[378], line_14[376], line_13[374], line_12[372], line_11[370], line_10[368], line_9[366], line_8[364], line_7[362], line_6[360], line_5[358], line_4[356], line_3[354], line_2[352], line_1[350] };
assign col_605 = {line_128[605], line_127[603], line_126[601], line_125[599], line_124[597], line_123[595], line_122[593], line_121[591], line_120[589], line_119[587], line_118[585], line_117[583], line_116[581], line_115[579], line_114[577], line_113[575], line_112[573], line_111[571], line_110[569], line_109[567], line_108[565], line_107[563], line_106[561], line_105[559], line_104[557], line_103[555], line_102[553], line_101[551], line_100[549], line_99[547], line_98[545], line_97[543], line_96[541], line_95[539], line_94[537], line_93[535], line_92[533], line_91[531], line_90[529], line_89[527], line_88[525], line_87[523], line_86[521], line_85[519], line_84[517], line_83[515], line_82[513], line_81[511], line_80[509], line_79[507], line_78[505], line_77[503], line_76[501], line_75[499], line_74[497], line_73[495], line_72[493], line_71[491], line_70[489], line_69[487], line_68[485], line_67[483], line_66[481], line_65[479], line_64[477], line_63[475], line_62[473], line_61[471], line_60[469], line_59[467], line_58[465], line_57[463], line_56[461], line_55[459], line_54[457], line_53[455], line_52[453], line_51[451], line_50[449], line_49[447], line_48[445], line_47[443], line_46[441], line_45[439], line_44[437], line_43[435], line_42[433], line_41[431], line_40[429], line_39[427], line_38[425], line_37[423], line_36[421], line_35[419], line_34[417], line_33[415], line_32[413], line_31[411], line_30[409], line_29[407], line_28[405], line_27[403], line_26[401], line_25[399], line_24[397], line_23[395], line_22[393], line_21[391], line_20[389], line_19[387], line_18[385], line_17[383], line_16[381], line_15[379], line_14[377], line_13[375], line_12[373], line_11[371], line_10[369], line_9[367], line_8[365], line_7[363], line_6[361], line_5[359], line_4[357], line_3[355], line_2[353], line_1[351] };
assign col_606 = {line_128[606], line_127[604], line_126[602], line_125[600], line_124[598], line_123[596], line_122[594], line_121[592], line_120[590], line_119[588], line_118[586], line_117[584], line_116[582], line_115[580], line_114[578], line_113[576], line_112[574], line_111[572], line_110[570], line_109[568], line_108[566], line_107[564], line_106[562], line_105[560], line_104[558], line_103[556], line_102[554], line_101[552], line_100[550], line_99[548], line_98[546], line_97[544], line_96[542], line_95[540], line_94[538], line_93[536], line_92[534], line_91[532], line_90[530], line_89[528], line_88[526], line_87[524], line_86[522], line_85[520], line_84[518], line_83[516], line_82[514], line_81[512], line_80[510], line_79[508], line_78[506], line_77[504], line_76[502], line_75[500], line_74[498], line_73[496], line_72[494], line_71[492], line_70[490], line_69[488], line_68[486], line_67[484], line_66[482], line_65[480], line_64[478], line_63[476], line_62[474], line_61[472], line_60[470], line_59[468], line_58[466], line_57[464], line_56[462], line_55[460], line_54[458], line_53[456], line_52[454], line_51[452], line_50[450], line_49[448], line_48[446], line_47[444], line_46[442], line_45[440], line_44[438], line_43[436], line_42[434], line_41[432], line_40[430], line_39[428], line_38[426], line_37[424], line_36[422], line_35[420], line_34[418], line_33[416], line_32[414], line_31[412], line_30[410], line_29[408], line_28[406], line_27[404], line_26[402], line_25[400], line_24[398], line_23[396], line_22[394], line_21[392], line_20[390], line_19[388], line_18[386], line_17[384], line_16[382], line_15[380], line_14[378], line_13[376], line_12[374], line_11[372], line_10[370], line_9[368], line_8[366], line_7[364], line_6[362], line_5[360], line_4[358], line_3[356], line_2[354], line_1[352] };
assign col_607 = {line_128[607], line_127[605], line_126[603], line_125[601], line_124[599], line_123[597], line_122[595], line_121[593], line_120[591], line_119[589], line_118[587], line_117[585], line_116[583], line_115[581], line_114[579], line_113[577], line_112[575], line_111[573], line_110[571], line_109[569], line_108[567], line_107[565], line_106[563], line_105[561], line_104[559], line_103[557], line_102[555], line_101[553], line_100[551], line_99[549], line_98[547], line_97[545], line_96[543], line_95[541], line_94[539], line_93[537], line_92[535], line_91[533], line_90[531], line_89[529], line_88[527], line_87[525], line_86[523], line_85[521], line_84[519], line_83[517], line_82[515], line_81[513], line_80[511], line_79[509], line_78[507], line_77[505], line_76[503], line_75[501], line_74[499], line_73[497], line_72[495], line_71[493], line_70[491], line_69[489], line_68[487], line_67[485], line_66[483], line_65[481], line_64[479], line_63[477], line_62[475], line_61[473], line_60[471], line_59[469], line_58[467], line_57[465], line_56[463], line_55[461], line_54[459], line_53[457], line_52[455], line_51[453], line_50[451], line_49[449], line_48[447], line_47[445], line_46[443], line_45[441], line_44[439], line_43[437], line_42[435], line_41[433], line_40[431], line_39[429], line_38[427], line_37[425], line_36[423], line_35[421], line_34[419], line_33[417], line_32[415], line_31[413], line_30[411], line_29[409], line_28[407], line_27[405], line_26[403], line_25[401], line_24[399], line_23[397], line_22[395], line_21[393], line_20[391], line_19[389], line_18[387], line_17[385], line_16[383], line_15[381], line_14[379], line_13[377], line_12[375], line_11[373], line_10[371], line_9[369], line_8[367], line_7[365], line_6[363], line_5[361], line_4[359], line_3[357], line_2[355], line_1[353] };
assign col_608 = {line_128[608], line_127[606], line_126[604], line_125[602], line_124[600], line_123[598], line_122[596], line_121[594], line_120[592], line_119[590], line_118[588], line_117[586], line_116[584], line_115[582], line_114[580], line_113[578], line_112[576], line_111[574], line_110[572], line_109[570], line_108[568], line_107[566], line_106[564], line_105[562], line_104[560], line_103[558], line_102[556], line_101[554], line_100[552], line_99[550], line_98[548], line_97[546], line_96[544], line_95[542], line_94[540], line_93[538], line_92[536], line_91[534], line_90[532], line_89[530], line_88[528], line_87[526], line_86[524], line_85[522], line_84[520], line_83[518], line_82[516], line_81[514], line_80[512], line_79[510], line_78[508], line_77[506], line_76[504], line_75[502], line_74[500], line_73[498], line_72[496], line_71[494], line_70[492], line_69[490], line_68[488], line_67[486], line_66[484], line_65[482], line_64[480], line_63[478], line_62[476], line_61[474], line_60[472], line_59[470], line_58[468], line_57[466], line_56[464], line_55[462], line_54[460], line_53[458], line_52[456], line_51[454], line_50[452], line_49[450], line_48[448], line_47[446], line_46[444], line_45[442], line_44[440], line_43[438], line_42[436], line_41[434], line_40[432], line_39[430], line_38[428], line_37[426], line_36[424], line_35[422], line_34[420], line_33[418], line_32[416], line_31[414], line_30[412], line_29[410], line_28[408], line_27[406], line_26[404], line_25[402], line_24[400], line_23[398], line_22[396], line_21[394], line_20[392], line_19[390], line_18[388], line_17[386], line_16[384], line_15[382], line_14[380], line_13[378], line_12[376], line_11[374], line_10[372], line_9[370], line_8[368], line_7[366], line_6[364], line_5[362], line_4[360], line_3[358], line_2[356], line_1[354] };
assign col_609 = {line_128[609], line_127[607], line_126[605], line_125[603], line_124[601], line_123[599], line_122[597], line_121[595], line_120[593], line_119[591], line_118[589], line_117[587], line_116[585], line_115[583], line_114[581], line_113[579], line_112[577], line_111[575], line_110[573], line_109[571], line_108[569], line_107[567], line_106[565], line_105[563], line_104[561], line_103[559], line_102[557], line_101[555], line_100[553], line_99[551], line_98[549], line_97[547], line_96[545], line_95[543], line_94[541], line_93[539], line_92[537], line_91[535], line_90[533], line_89[531], line_88[529], line_87[527], line_86[525], line_85[523], line_84[521], line_83[519], line_82[517], line_81[515], line_80[513], line_79[511], line_78[509], line_77[507], line_76[505], line_75[503], line_74[501], line_73[499], line_72[497], line_71[495], line_70[493], line_69[491], line_68[489], line_67[487], line_66[485], line_65[483], line_64[481], line_63[479], line_62[477], line_61[475], line_60[473], line_59[471], line_58[469], line_57[467], line_56[465], line_55[463], line_54[461], line_53[459], line_52[457], line_51[455], line_50[453], line_49[451], line_48[449], line_47[447], line_46[445], line_45[443], line_44[441], line_43[439], line_42[437], line_41[435], line_40[433], line_39[431], line_38[429], line_37[427], line_36[425], line_35[423], line_34[421], line_33[419], line_32[417], line_31[415], line_30[413], line_29[411], line_28[409], line_27[407], line_26[405], line_25[403], line_24[401], line_23[399], line_22[397], line_21[395], line_20[393], line_19[391], line_18[389], line_17[387], line_16[385], line_15[383], line_14[381], line_13[379], line_12[377], line_11[375], line_10[373], line_9[371], line_8[369], line_7[367], line_6[365], line_5[363], line_4[361], line_3[359], line_2[357], line_1[355] };
assign col_610 = {line_128[610], line_127[608], line_126[606], line_125[604], line_124[602], line_123[600], line_122[598], line_121[596], line_120[594], line_119[592], line_118[590], line_117[588], line_116[586], line_115[584], line_114[582], line_113[580], line_112[578], line_111[576], line_110[574], line_109[572], line_108[570], line_107[568], line_106[566], line_105[564], line_104[562], line_103[560], line_102[558], line_101[556], line_100[554], line_99[552], line_98[550], line_97[548], line_96[546], line_95[544], line_94[542], line_93[540], line_92[538], line_91[536], line_90[534], line_89[532], line_88[530], line_87[528], line_86[526], line_85[524], line_84[522], line_83[520], line_82[518], line_81[516], line_80[514], line_79[512], line_78[510], line_77[508], line_76[506], line_75[504], line_74[502], line_73[500], line_72[498], line_71[496], line_70[494], line_69[492], line_68[490], line_67[488], line_66[486], line_65[484], line_64[482], line_63[480], line_62[478], line_61[476], line_60[474], line_59[472], line_58[470], line_57[468], line_56[466], line_55[464], line_54[462], line_53[460], line_52[458], line_51[456], line_50[454], line_49[452], line_48[450], line_47[448], line_46[446], line_45[444], line_44[442], line_43[440], line_42[438], line_41[436], line_40[434], line_39[432], line_38[430], line_37[428], line_36[426], line_35[424], line_34[422], line_33[420], line_32[418], line_31[416], line_30[414], line_29[412], line_28[410], line_27[408], line_26[406], line_25[404], line_24[402], line_23[400], line_22[398], line_21[396], line_20[394], line_19[392], line_18[390], line_17[388], line_16[386], line_15[384], line_14[382], line_13[380], line_12[378], line_11[376], line_10[374], line_9[372], line_8[370], line_7[368], line_6[366], line_5[364], line_4[362], line_3[360], line_2[358], line_1[356] };
assign col_611 = {line_128[611], line_127[609], line_126[607], line_125[605], line_124[603], line_123[601], line_122[599], line_121[597], line_120[595], line_119[593], line_118[591], line_117[589], line_116[587], line_115[585], line_114[583], line_113[581], line_112[579], line_111[577], line_110[575], line_109[573], line_108[571], line_107[569], line_106[567], line_105[565], line_104[563], line_103[561], line_102[559], line_101[557], line_100[555], line_99[553], line_98[551], line_97[549], line_96[547], line_95[545], line_94[543], line_93[541], line_92[539], line_91[537], line_90[535], line_89[533], line_88[531], line_87[529], line_86[527], line_85[525], line_84[523], line_83[521], line_82[519], line_81[517], line_80[515], line_79[513], line_78[511], line_77[509], line_76[507], line_75[505], line_74[503], line_73[501], line_72[499], line_71[497], line_70[495], line_69[493], line_68[491], line_67[489], line_66[487], line_65[485], line_64[483], line_63[481], line_62[479], line_61[477], line_60[475], line_59[473], line_58[471], line_57[469], line_56[467], line_55[465], line_54[463], line_53[461], line_52[459], line_51[457], line_50[455], line_49[453], line_48[451], line_47[449], line_46[447], line_45[445], line_44[443], line_43[441], line_42[439], line_41[437], line_40[435], line_39[433], line_38[431], line_37[429], line_36[427], line_35[425], line_34[423], line_33[421], line_32[419], line_31[417], line_30[415], line_29[413], line_28[411], line_27[409], line_26[407], line_25[405], line_24[403], line_23[401], line_22[399], line_21[397], line_20[395], line_19[393], line_18[391], line_17[389], line_16[387], line_15[385], line_14[383], line_13[381], line_12[379], line_11[377], line_10[375], line_9[373], line_8[371], line_7[369], line_6[367], line_5[365], line_4[363], line_3[361], line_2[359], line_1[357] };
assign col_612 = {line_128[612], line_127[610], line_126[608], line_125[606], line_124[604], line_123[602], line_122[600], line_121[598], line_120[596], line_119[594], line_118[592], line_117[590], line_116[588], line_115[586], line_114[584], line_113[582], line_112[580], line_111[578], line_110[576], line_109[574], line_108[572], line_107[570], line_106[568], line_105[566], line_104[564], line_103[562], line_102[560], line_101[558], line_100[556], line_99[554], line_98[552], line_97[550], line_96[548], line_95[546], line_94[544], line_93[542], line_92[540], line_91[538], line_90[536], line_89[534], line_88[532], line_87[530], line_86[528], line_85[526], line_84[524], line_83[522], line_82[520], line_81[518], line_80[516], line_79[514], line_78[512], line_77[510], line_76[508], line_75[506], line_74[504], line_73[502], line_72[500], line_71[498], line_70[496], line_69[494], line_68[492], line_67[490], line_66[488], line_65[486], line_64[484], line_63[482], line_62[480], line_61[478], line_60[476], line_59[474], line_58[472], line_57[470], line_56[468], line_55[466], line_54[464], line_53[462], line_52[460], line_51[458], line_50[456], line_49[454], line_48[452], line_47[450], line_46[448], line_45[446], line_44[444], line_43[442], line_42[440], line_41[438], line_40[436], line_39[434], line_38[432], line_37[430], line_36[428], line_35[426], line_34[424], line_33[422], line_32[420], line_31[418], line_30[416], line_29[414], line_28[412], line_27[410], line_26[408], line_25[406], line_24[404], line_23[402], line_22[400], line_21[398], line_20[396], line_19[394], line_18[392], line_17[390], line_16[388], line_15[386], line_14[384], line_13[382], line_12[380], line_11[378], line_10[376], line_9[374], line_8[372], line_7[370], line_6[368], line_5[366], line_4[364], line_3[362], line_2[360], line_1[358] };
assign col_613 = {line_128[613], line_127[611], line_126[609], line_125[607], line_124[605], line_123[603], line_122[601], line_121[599], line_120[597], line_119[595], line_118[593], line_117[591], line_116[589], line_115[587], line_114[585], line_113[583], line_112[581], line_111[579], line_110[577], line_109[575], line_108[573], line_107[571], line_106[569], line_105[567], line_104[565], line_103[563], line_102[561], line_101[559], line_100[557], line_99[555], line_98[553], line_97[551], line_96[549], line_95[547], line_94[545], line_93[543], line_92[541], line_91[539], line_90[537], line_89[535], line_88[533], line_87[531], line_86[529], line_85[527], line_84[525], line_83[523], line_82[521], line_81[519], line_80[517], line_79[515], line_78[513], line_77[511], line_76[509], line_75[507], line_74[505], line_73[503], line_72[501], line_71[499], line_70[497], line_69[495], line_68[493], line_67[491], line_66[489], line_65[487], line_64[485], line_63[483], line_62[481], line_61[479], line_60[477], line_59[475], line_58[473], line_57[471], line_56[469], line_55[467], line_54[465], line_53[463], line_52[461], line_51[459], line_50[457], line_49[455], line_48[453], line_47[451], line_46[449], line_45[447], line_44[445], line_43[443], line_42[441], line_41[439], line_40[437], line_39[435], line_38[433], line_37[431], line_36[429], line_35[427], line_34[425], line_33[423], line_32[421], line_31[419], line_30[417], line_29[415], line_28[413], line_27[411], line_26[409], line_25[407], line_24[405], line_23[403], line_22[401], line_21[399], line_20[397], line_19[395], line_18[393], line_17[391], line_16[389], line_15[387], line_14[385], line_13[383], line_12[381], line_11[379], line_10[377], line_9[375], line_8[373], line_7[371], line_6[369], line_5[367], line_4[365], line_3[363], line_2[361], line_1[359] };
assign col_614 = {line_128[614], line_127[612], line_126[610], line_125[608], line_124[606], line_123[604], line_122[602], line_121[600], line_120[598], line_119[596], line_118[594], line_117[592], line_116[590], line_115[588], line_114[586], line_113[584], line_112[582], line_111[580], line_110[578], line_109[576], line_108[574], line_107[572], line_106[570], line_105[568], line_104[566], line_103[564], line_102[562], line_101[560], line_100[558], line_99[556], line_98[554], line_97[552], line_96[550], line_95[548], line_94[546], line_93[544], line_92[542], line_91[540], line_90[538], line_89[536], line_88[534], line_87[532], line_86[530], line_85[528], line_84[526], line_83[524], line_82[522], line_81[520], line_80[518], line_79[516], line_78[514], line_77[512], line_76[510], line_75[508], line_74[506], line_73[504], line_72[502], line_71[500], line_70[498], line_69[496], line_68[494], line_67[492], line_66[490], line_65[488], line_64[486], line_63[484], line_62[482], line_61[480], line_60[478], line_59[476], line_58[474], line_57[472], line_56[470], line_55[468], line_54[466], line_53[464], line_52[462], line_51[460], line_50[458], line_49[456], line_48[454], line_47[452], line_46[450], line_45[448], line_44[446], line_43[444], line_42[442], line_41[440], line_40[438], line_39[436], line_38[434], line_37[432], line_36[430], line_35[428], line_34[426], line_33[424], line_32[422], line_31[420], line_30[418], line_29[416], line_28[414], line_27[412], line_26[410], line_25[408], line_24[406], line_23[404], line_22[402], line_21[400], line_20[398], line_19[396], line_18[394], line_17[392], line_16[390], line_15[388], line_14[386], line_13[384], line_12[382], line_11[380], line_10[378], line_9[376], line_8[374], line_7[372], line_6[370], line_5[368], line_4[366], line_3[364], line_2[362], line_1[360] };
assign col_615 = {line_128[615], line_127[613], line_126[611], line_125[609], line_124[607], line_123[605], line_122[603], line_121[601], line_120[599], line_119[597], line_118[595], line_117[593], line_116[591], line_115[589], line_114[587], line_113[585], line_112[583], line_111[581], line_110[579], line_109[577], line_108[575], line_107[573], line_106[571], line_105[569], line_104[567], line_103[565], line_102[563], line_101[561], line_100[559], line_99[557], line_98[555], line_97[553], line_96[551], line_95[549], line_94[547], line_93[545], line_92[543], line_91[541], line_90[539], line_89[537], line_88[535], line_87[533], line_86[531], line_85[529], line_84[527], line_83[525], line_82[523], line_81[521], line_80[519], line_79[517], line_78[515], line_77[513], line_76[511], line_75[509], line_74[507], line_73[505], line_72[503], line_71[501], line_70[499], line_69[497], line_68[495], line_67[493], line_66[491], line_65[489], line_64[487], line_63[485], line_62[483], line_61[481], line_60[479], line_59[477], line_58[475], line_57[473], line_56[471], line_55[469], line_54[467], line_53[465], line_52[463], line_51[461], line_50[459], line_49[457], line_48[455], line_47[453], line_46[451], line_45[449], line_44[447], line_43[445], line_42[443], line_41[441], line_40[439], line_39[437], line_38[435], line_37[433], line_36[431], line_35[429], line_34[427], line_33[425], line_32[423], line_31[421], line_30[419], line_29[417], line_28[415], line_27[413], line_26[411], line_25[409], line_24[407], line_23[405], line_22[403], line_21[401], line_20[399], line_19[397], line_18[395], line_17[393], line_16[391], line_15[389], line_14[387], line_13[385], line_12[383], line_11[381], line_10[379], line_9[377], line_8[375], line_7[373], line_6[371], line_5[369], line_4[367], line_3[365], line_2[363], line_1[361] };
assign col_616 = {line_128[616], line_127[614], line_126[612], line_125[610], line_124[608], line_123[606], line_122[604], line_121[602], line_120[600], line_119[598], line_118[596], line_117[594], line_116[592], line_115[590], line_114[588], line_113[586], line_112[584], line_111[582], line_110[580], line_109[578], line_108[576], line_107[574], line_106[572], line_105[570], line_104[568], line_103[566], line_102[564], line_101[562], line_100[560], line_99[558], line_98[556], line_97[554], line_96[552], line_95[550], line_94[548], line_93[546], line_92[544], line_91[542], line_90[540], line_89[538], line_88[536], line_87[534], line_86[532], line_85[530], line_84[528], line_83[526], line_82[524], line_81[522], line_80[520], line_79[518], line_78[516], line_77[514], line_76[512], line_75[510], line_74[508], line_73[506], line_72[504], line_71[502], line_70[500], line_69[498], line_68[496], line_67[494], line_66[492], line_65[490], line_64[488], line_63[486], line_62[484], line_61[482], line_60[480], line_59[478], line_58[476], line_57[474], line_56[472], line_55[470], line_54[468], line_53[466], line_52[464], line_51[462], line_50[460], line_49[458], line_48[456], line_47[454], line_46[452], line_45[450], line_44[448], line_43[446], line_42[444], line_41[442], line_40[440], line_39[438], line_38[436], line_37[434], line_36[432], line_35[430], line_34[428], line_33[426], line_32[424], line_31[422], line_30[420], line_29[418], line_28[416], line_27[414], line_26[412], line_25[410], line_24[408], line_23[406], line_22[404], line_21[402], line_20[400], line_19[398], line_18[396], line_17[394], line_16[392], line_15[390], line_14[388], line_13[386], line_12[384], line_11[382], line_10[380], line_9[378], line_8[376], line_7[374], line_6[372], line_5[370], line_4[368], line_3[366], line_2[364], line_1[362] };
assign col_617 = {line_128[617], line_127[615], line_126[613], line_125[611], line_124[609], line_123[607], line_122[605], line_121[603], line_120[601], line_119[599], line_118[597], line_117[595], line_116[593], line_115[591], line_114[589], line_113[587], line_112[585], line_111[583], line_110[581], line_109[579], line_108[577], line_107[575], line_106[573], line_105[571], line_104[569], line_103[567], line_102[565], line_101[563], line_100[561], line_99[559], line_98[557], line_97[555], line_96[553], line_95[551], line_94[549], line_93[547], line_92[545], line_91[543], line_90[541], line_89[539], line_88[537], line_87[535], line_86[533], line_85[531], line_84[529], line_83[527], line_82[525], line_81[523], line_80[521], line_79[519], line_78[517], line_77[515], line_76[513], line_75[511], line_74[509], line_73[507], line_72[505], line_71[503], line_70[501], line_69[499], line_68[497], line_67[495], line_66[493], line_65[491], line_64[489], line_63[487], line_62[485], line_61[483], line_60[481], line_59[479], line_58[477], line_57[475], line_56[473], line_55[471], line_54[469], line_53[467], line_52[465], line_51[463], line_50[461], line_49[459], line_48[457], line_47[455], line_46[453], line_45[451], line_44[449], line_43[447], line_42[445], line_41[443], line_40[441], line_39[439], line_38[437], line_37[435], line_36[433], line_35[431], line_34[429], line_33[427], line_32[425], line_31[423], line_30[421], line_29[419], line_28[417], line_27[415], line_26[413], line_25[411], line_24[409], line_23[407], line_22[405], line_21[403], line_20[401], line_19[399], line_18[397], line_17[395], line_16[393], line_15[391], line_14[389], line_13[387], line_12[385], line_11[383], line_10[381], line_9[379], line_8[377], line_7[375], line_6[373], line_5[371], line_4[369], line_3[367], line_2[365], line_1[363] };
assign col_618 = {line_128[618], line_127[616], line_126[614], line_125[612], line_124[610], line_123[608], line_122[606], line_121[604], line_120[602], line_119[600], line_118[598], line_117[596], line_116[594], line_115[592], line_114[590], line_113[588], line_112[586], line_111[584], line_110[582], line_109[580], line_108[578], line_107[576], line_106[574], line_105[572], line_104[570], line_103[568], line_102[566], line_101[564], line_100[562], line_99[560], line_98[558], line_97[556], line_96[554], line_95[552], line_94[550], line_93[548], line_92[546], line_91[544], line_90[542], line_89[540], line_88[538], line_87[536], line_86[534], line_85[532], line_84[530], line_83[528], line_82[526], line_81[524], line_80[522], line_79[520], line_78[518], line_77[516], line_76[514], line_75[512], line_74[510], line_73[508], line_72[506], line_71[504], line_70[502], line_69[500], line_68[498], line_67[496], line_66[494], line_65[492], line_64[490], line_63[488], line_62[486], line_61[484], line_60[482], line_59[480], line_58[478], line_57[476], line_56[474], line_55[472], line_54[470], line_53[468], line_52[466], line_51[464], line_50[462], line_49[460], line_48[458], line_47[456], line_46[454], line_45[452], line_44[450], line_43[448], line_42[446], line_41[444], line_40[442], line_39[440], line_38[438], line_37[436], line_36[434], line_35[432], line_34[430], line_33[428], line_32[426], line_31[424], line_30[422], line_29[420], line_28[418], line_27[416], line_26[414], line_25[412], line_24[410], line_23[408], line_22[406], line_21[404], line_20[402], line_19[400], line_18[398], line_17[396], line_16[394], line_15[392], line_14[390], line_13[388], line_12[386], line_11[384], line_10[382], line_9[380], line_8[378], line_7[376], line_6[374], line_5[372], line_4[370], line_3[368], line_2[366], line_1[364] };
assign col_619 = {line_128[619], line_127[617], line_126[615], line_125[613], line_124[611], line_123[609], line_122[607], line_121[605], line_120[603], line_119[601], line_118[599], line_117[597], line_116[595], line_115[593], line_114[591], line_113[589], line_112[587], line_111[585], line_110[583], line_109[581], line_108[579], line_107[577], line_106[575], line_105[573], line_104[571], line_103[569], line_102[567], line_101[565], line_100[563], line_99[561], line_98[559], line_97[557], line_96[555], line_95[553], line_94[551], line_93[549], line_92[547], line_91[545], line_90[543], line_89[541], line_88[539], line_87[537], line_86[535], line_85[533], line_84[531], line_83[529], line_82[527], line_81[525], line_80[523], line_79[521], line_78[519], line_77[517], line_76[515], line_75[513], line_74[511], line_73[509], line_72[507], line_71[505], line_70[503], line_69[501], line_68[499], line_67[497], line_66[495], line_65[493], line_64[491], line_63[489], line_62[487], line_61[485], line_60[483], line_59[481], line_58[479], line_57[477], line_56[475], line_55[473], line_54[471], line_53[469], line_52[467], line_51[465], line_50[463], line_49[461], line_48[459], line_47[457], line_46[455], line_45[453], line_44[451], line_43[449], line_42[447], line_41[445], line_40[443], line_39[441], line_38[439], line_37[437], line_36[435], line_35[433], line_34[431], line_33[429], line_32[427], line_31[425], line_30[423], line_29[421], line_28[419], line_27[417], line_26[415], line_25[413], line_24[411], line_23[409], line_22[407], line_21[405], line_20[403], line_19[401], line_18[399], line_17[397], line_16[395], line_15[393], line_14[391], line_13[389], line_12[387], line_11[385], line_10[383], line_9[381], line_8[379], line_7[377], line_6[375], line_5[373], line_4[371], line_3[369], line_2[367], line_1[365] };
assign col_620 = {line_128[620], line_127[618], line_126[616], line_125[614], line_124[612], line_123[610], line_122[608], line_121[606], line_120[604], line_119[602], line_118[600], line_117[598], line_116[596], line_115[594], line_114[592], line_113[590], line_112[588], line_111[586], line_110[584], line_109[582], line_108[580], line_107[578], line_106[576], line_105[574], line_104[572], line_103[570], line_102[568], line_101[566], line_100[564], line_99[562], line_98[560], line_97[558], line_96[556], line_95[554], line_94[552], line_93[550], line_92[548], line_91[546], line_90[544], line_89[542], line_88[540], line_87[538], line_86[536], line_85[534], line_84[532], line_83[530], line_82[528], line_81[526], line_80[524], line_79[522], line_78[520], line_77[518], line_76[516], line_75[514], line_74[512], line_73[510], line_72[508], line_71[506], line_70[504], line_69[502], line_68[500], line_67[498], line_66[496], line_65[494], line_64[492], line_63[490], line_62[488], line_61[486], line_60[484], line_59[482], line_58[480], line_57[478], line_56[476], line_55[474], line_54[472], line_53[470], line_52[468], line_51[466], line_50[464], line_49[462], line_48[460], line_47[458], line_46[456], line_45[454], line_44[452], line_43[450], line_42[448], line_41[446], line_40[444], line_39[442], line_38[440], line_37[438], line_36[436], line_35[434], line_34[432], line_33[430], line_32[428], line_31[426], line_30[424], line_29[422], line_28[420], line_27[418], line_26[416], line_25[414], line_24[412], line_23[410], line_22[408], line_21[406], line_20[404], line_19[402], line_18[400], line_17[398], line_16[396], line_15[394], line_14[392], line_13[390], line_12[388], line_11[386], line_10[384], line_9[382], line_8[380], line_7[378], line_6[376], line_5[374], line_4[372], line_3[370], line_2[368], line_1[366] };
assign col_621 = {line_128[621], line_127[619], line_126[617], line_125[615], line_124[613], line_123[611], line_122[609], line_121[607], line_120[605], line_119[603], line_118[601], line_117[599], line_116[597], line_115[595], line_114[593], line_113[591], line_112[589], line_111[587], line_110[585], line_109[583], line_108[581], line_107[579], line_106[577], line_105[575], line_104[573], line_103[571], line_102[569], line_101[567], line_100[565], line_99[563], line_98[561], line_97[559], line_96[557], line_95[555], line_94[553], line_93[551], line_92[549], line_91[547], line_90[545], line_89[543], line_88[541], line_87[539], line_86[537], line_85[535], line_84[533], line_83[531], line_82[529], line_81[527], line_80[525], line_79[523], line_78[521], line_77[519], line_76[517], line_75[515], line_74[513], line_73[511], line_72[509], line_71[507], line_70[505], line_69[503], line_68[501], line_67[499], line_66[497], line_65[495], line_64[493], line_63[491], line_62[489], line_61[487], line_60[485], line_59[483], line_58[481], line_57[479], line_56[477], line_55[475], line_54[473], line_53[471], line_52[469], line_51[467], line_50[465], line_49[463], line_48[461], line_47[459], line_46[457], line_45[455], line_44[453], line_43[451], line_42[449], line_41[447], line_40[445], line_39[443], line_38[441], line_37[439], line_36[437], line_35[435], line_34[433], line_33[431], line_32[429], line_31[427], line_30[425], line_29[423], line_28[421], line_27[419], line_26[417], line_25[415], line_24[413], line_23[411], line_22[409], line_21[407], line_20[405], line_19[403], line_18[401], line_17[399], line_16[397], line_15[395], line_14[393], line_13[391], line_12[389], line_11[387], line_10[385], line_9[383], line_8[381], line_7[379], line_6[377], line_5[375], line_4[373], line_3[371], line_2[369], line_1[367] };
assign col_622 = {line_128[622], line_127[620], line_126[618], line_125[616], line_124[614], line_123[612], line_122[610], line_121[608], line_120[606], line_119[604], line_118[602], line_117[600], line_116[598], line_115[596], line_114[594], line_113[592], line_112[590], line_111[588], line_110[586], line_109[584], line_108[582], line_107[580], line_106[578], line_105[576], line_104[574], line_103[572], line_102[570], line_101[568], line_100[566], line_99[564], line_98[562], line_97[560], line_96[558], line_95[556], line_94[554], line_93[552], line_92[550], line_91[548], line_90[546], line_89[544], line_88[542], line_87[540], line_86[538], line_85[536], line_84[534], line_83[532], line_82[530], line_81[528], line_80[526], line_79[524], line_78[522], line_77[520], line_76[518], line_75[516], line_74[514], line_73[512], line_72[510], line_71[508], line_70[506], line_69[504], line_68[502], line_67[500], line_66[498], line_65[496], line_64[494], line_63[492], line_62[490], line_61[488], line_60[486], line_59[484], line_58[482], line_57[480], line_56[478], line_55[476], line_54[474], line_53[472], line_52[470], line_51[468], line_50[466], line_49[464], line_48[462], line_47[460], line_46[458], line_45[456], line_44[454], line_43[452], line_42[450], line_41[448], line_40[446], line_39[444], line_38[442], line_37[440], line_36[438], line_35[436], line_34[434], line_33[432], line_32[430], line_31[428], line_30[426], line_29[424], line_28[422], line_27[420], line_26[418], line_25[416], line_24[414], line_23[412], line_22[410], line_21[408], line_20[406], line_19[404], line_18[402], line_17[400], line_16[398], line_15[396], line_14[394], line_13[392], line_12[390], line_11[388], line_10[386], line_9[384], line_8[382], line_7[380], line_6[378], line_5[376], line_4[374], line_3[372], line_2[370], line_1[368] };
assign col_623 = {line_128[623], line_127[621], line_126[619], line_125[617], line_124[615], line_123[613], line_122[611], line_121[609], line_120[607], line_119[605], line_118[603], line_117[601], line_116[599], line_115[597], line_114[595], line_113[593], line_112[591], line_111[589], line_110[587], line_109[585], line_108[583], line_107[581], line_106[579], line_105[577], line_104[575], line_103[573], line_102[571], line_101[569], line_100[567], line_99[565], line_98[563], line_97[561], line_96[559], line_95[557], line_94[555], line_93[553], line_92[551], line_91[549], line_90[547], line_89[545], line_88[543], line_87[541], line_86[539], line_85[537], line_84[535], line_83[533], line_82[531], line_81[529], line_80[527], line_79[525], line_78[523], line_77[521], line_76[519], line_75[517], line_74[515], line_73[513], line_72[511], line_71[509], line_70[507], line_69[505], line_68[503], line_67[501], line_66[499], line_65[497], line_64[495], line_63[493], line_62[491], line_61[489], line_60[487], line_59[485], line_58[483], line_57[481], line_56[479], line_55[477], line_54[475], line_53[473], line_52[471], line_51[469], line_50[467], line_49[465], line_48[463], line_47[461], line_46[459], line_45[457], line_44[455], line_43[453], line_42[451], line_41[449], line_40[447], line_39[445], line_38[443], line_37[441], line_36[439], line_35[437], line_34[435], line_33[433], line_32[431], line_31[429], line_30[427], line_29[425], line_28[423], line_27[421], line_26[419], line_25[417], line_24[415], line_23[413], line_22[411], line_21[409], line_20[407], line_19[405], line_18[403], line_17[401], line_16[399], line_15[397], line_14[395], line_13[393], line_12[391], line_11[389], line_10[387], line_9[385], line_8[383], line_7[381], line_6[379], line_5[377], line_4[375], line_3[373], line_2[371], line_1[369] };
assign col_624 = {line_128[624], line_127[622], line_126[620], line_125[618], line_124[616], line_123[614], line_122[612], line_121[610], line_120[608], line_119[606], line_118[604], line_117[602], line_116[600], line_115[598], line_114[596], line_113[594], line_112[592], line_111[590], line_110[588], line_109[586], line_108[584], line_107[582], line_106[580], line_105[578], line_104[576], line_103[574], line_102[572], line_101[570], line_100[568], line_99[566], line_98[564], line_97[562], line_96[560], line_95[558], line_94[556], line_93[554], line_92[552], line_91[550], line_90[548], line_89[546], line_88[544], line_87[542], line_86[540], line_85[538], line_84[536], line_83[534], line_82[532], line_81[530], line_80[528], line_79[526], line_78[524], line_77[522], line_76[520], line_75[518], line_74[516], line_73[514], line_72[512], line_71[510], line_70[508], line_69[506], line_68[504], line_67[502], line_66[500], line_65[498], line_64[496], line_63[494], line_62[492], line_61[490], line_60[488], line_59[486], line_58[484], line_57[482], line_56[480], line_55[478], line_54[476], line_53[474], line_52[472], line_51[470], line_50[468], line_49[466], line_48[464], line_47[462], line_46[460], line_45[458], line_44[456], line_43[454], line_42[452], line_41[450], line_40[448], line_39[446], line_38[444], line_37[442], line_36[440], line_35[438], line_34[436], line_33[434], line_32[432], line_31[430], line_30[428], line_29[426], line_28[424], line_27[422], line_26[420], line_25[418], line_24[416], line_23[414], line_22[412], line_21[410], line_20[408], line_19[406], line_18[404], line_17[402], line_16[400], line_15[398], line_14[396], line_13[394], line_12[392], line_11[390], line_10[388], line_9[386], line_8[384], line_7[382], line_6[380], line_5[378], line_4[376], line_3[374], line_2[372], line_1[370] };
assign col_625 = {line_128[625], line_127[623], line_126[621], line_125[619], line_124[617], line_123[615], line_122[613], line_121[611], line_120[609], line_119[607], line_118[605], line_117[603], line_116[601], line_115[599], line_114[597], line_113[595], line_112[593], line_111[591], line_110[589], line_109[587], line_108[585], line_107[583], line_106[581], line_105[579], line_104[577], line_103[575], line_102[573], line_101[571], line_100[569], line_99[567], line_98[565], line_97[563], line_96[561], line_95[559], line_94[557], line_93[555], line_92[553], line_91[551], line_90[549], line_89[547], line_88[545], line_87[543], line_86[541], line_85[539], line_84[537], line_83[535], line_82[533], line_81[531], line_80[529], line_79[527], line_78[525], line_77[523], line_76[521], line_75[519], line_74[517], line_73[515], line_72[513], line_71[511], line_70[509], line_69[507], line_68[505], line_67[503], line_66[501], line_65[499], line_64[497], line_63[495], line_62[493], line_61[491], line_60[489], line_59[487], line_58[485], line_57[483], line_56[481], line_55[479], line_54[477], line_53[475], line_52[473], line_51[471], line_50[469], line_49[467], line_48[465], line_47[463], line_46[461], line_45[459], line_44[457], line_43[455], line_42[453], line_41[451], line_40[449], line_39[447], line_38[445], line_37[443], line_36[441], line_35[439], line_34[437], line_33[435], line_32[433], line_31[431], line_30[429], line_29[427], line_28[425], line_27[423], line_26[421], line_25[419], line_24[417], line_23[415], line_22[413], line_21[411], line_20[409], line_19[407], line_18[405], line_17[403], line_16[401], line_15[399], line_14[397], line_13[395], line_12[393], line_11[391], line_10[389], line_9[387], line_8[385], line_7[383], line_6[381], line_5[379], line_4[377], line_3[375], line_2[373], line_1[371] };
assign col_626 = {line_128[626], line_127[624], line_126[622], line_125[620], line_124[618], line_123[616], line_122[614], line_121[612], line_120[610], line_119[608], line_118[606], line_117[604], line_116[602], line_115[600], line_114[598], line_113[596], line_112[594], line_111[592], line_110[590], line_109[588], line_108[586], line_107[584], line_106[582], line_105[580], line_104[578], line_103[576], line_102[574], line_101[572], line_100[570], line_99[568], line_98[566], line_97[564], line_96[562], line_95[560], line_94[558], line_93[556], line_92[554], line_91[552], line_90[550], line_89[548], line_88[546], line_87[544], line_86[542], line_85[540], line_84[538], line_83[536], line_82[534], line_81[532], line_80[530], line_79[528], line_78[526], line_77[524], line_76[522], line_75[520], line_74[518], line_73[516], line_72[514], line_71[512], line_70[510], line_69[508], line_68[506], line_67[504], line_66[502], line_65[500], line_64[498], line_63[496], line_62[494], line_61[492], line_60[490], line_59[488], line_58[486], line_57[484], line_56[482], line_55[480], line_54[478], line_53[476], line_52[474], line_51[472], line_50[470], line_49[468], line_48[466], line_47[464], line_46[462], line_45[460], line_44[458], line_43[456], line_42[454], line_41[452], line_40[450], line_39[448], line_38[446], line_37[444], line_36[442], line_35[440], line_34[438], line_33[436], line_32[434], line_31[432], line_30[430], line_29[428], line_28[426], line_27[424], line_26[422], line_25[420], line_24[418], line_23[416], line_22[414], line_21[412], line_20[410], line_19[408], line_18[406], line_17[404], line_16[402], line_15[400], line_14[398], line_13[396], line_12[394], line_11[392], line_10[390], line_9[388], line_8[386], line_7[384], line_6[382], line_5[380], line_4[378], line_3[376], line_2[374], line_1[372] };
assign col_627 = {line_128[627], line_127[625], line_126[623], line_125[621], line_124[619], line_123[617], line_122[615], line_121[613], line_120[611], line_119[609], line_118[607], line_117[605], line_116[603], line_115[601], line_114[599], line_113[597], line_112[595], line_111[593], line_110[591], line_109[589], line_108[587], line_107[585], line_106[583], line_105[581], line_104[579], line_103[577], line_102[575], line_101[573], line_100[571], line_99[569], line_98[567], line_97[565], line_96[563], line_95[561], line_94[559], line_93[557], line_92[555], line_91[553], line_90[551], line_89[549], line_88[547], line_87[545], line_86[543], line_85[541], line_84[539], line_83[537], line_82[535], line_81[533], line_80[531], line_79[529], line_78[527], line_77[525], line_76[523], line_75[521], line_74[519], line_73[517], line_72[515], line_71[513], line_70[511], line_69[509], line_68[507], line_67[505], line_66[503], line_65[501], line_64[499], line_63[497], line_62[495], line_61[493], line_60[491], line_59[489], line_58[487], line_57[485], line_56[483], line_55[481], line_54[479], line_53[477], line_52[475], line_51[473], line_50[471], line_49[469], line_48[467], line_47[465], line_46[463], line_45[461], line_44[459], line_43[457], line_42[455], line_41[453], line_40[451], line_39[449], line_38[447], line_37[445], line_36[443], line_35[441], line_34[439], line_33[437], line_32[435], line_31[433], line_30[431], line_29[429], line_28[427], line_27[425], line_26[423], line_25[421], line_24[419], line_23[417], line_22[415], line_21[413], line_20[411], line_19[409], line_18[407], line_17[405], line_16[403], line_15[401], line_14[399], line_13[397], line_12[395], line_11[393], line_10[391], line_9[389], line_8[387], line_7[385], line_6[383], line_5[381], line_4[379], line_3[377], line_2[375], line_1[373] };
assign col_628 = {line_128[628], line_127[626], line_126[624], line_125[622], line_124[620], line_123[618], line_122[616], line_121[614], line_120[612], line_119[610], line_118[608], line_117[606], line_116[604], line_115[602], line_114[600], line_113[598], line_112[596], line_111[594], line_110[592], line_109[590], line_108[588], line_107[586], line_106[584], line_105[582], line_104[580], line_103[578], line_102[576], line_101[574], line_100[572], line_99[570], line_98[568], line_97[566], line_96[564], line_95[562], line_94[560], line_93[558], line_92[556], line_91[554], line_90[552], line_89[550], line_88[548], line_87[546], line_86[544], line_85[542], line_84[540], line_83[538], line_82[536], line_81[534], line_80[532], line_79[530], line_78[528], line_77[526], line_76[524], line_75[522], line_74[520], line_73[518], line_72[516], line_71[514], line_70[512], line_69[510], line_68[508], line_67[506], line_66[504], line_65[502], line_64[500], line_63[498], line_62[496], line_61[494], line_60[492], line_59[490], line_58[488], line_57[486], line_56[484], line_55[482], line_54[480], line_53[478], line_52[476], line_51[474], line_50[472], line_49[470], line_48[468], line_47[466], line_46[464], line_45[462], line_44[460], line_43[458], line_42[456], line_41[454], line_40[452], line_39[450], line_38[448], line_37[446], line_36[444], line_35[442], line_34[440], line_33[438], line_32[436], line_31[434], line_30[432], line_29[430], line_28[428], line_27[426], line_26[424], line_25[422], line_24[420], line_23[418], line_22[416], line_21[414], line_20[412], line_19[410], line_18[408], line_17[406], line_16[404], line_15[402], line_14[400], line_13[398], line_12[396], line_11[394], line_10[392], line_9[390], line_8[388], line_7[386], line_6[384], line_5[382], line_4[380], line_3[378], line_2[376], line_1[374] };
assign col_629 = {line_128[629], line_127[627], line_126[625], line_125[623], line_124[621], line_123[619], line_122[617], line_121[615], line_120[613], line_119[611], line_118[609], line_117[607], line_116[605], line_115[603], line_114[601], line_113[599], line_112[597], line_111[595], line_110[593], line_109[591], line_108[589], line_107[587], line_106[585], line_105[583], line_104[581], line_103[579], line_102[577], line_101[575], line_100[573], line_99[571], line_98[569], line_97[567], line_96[565], line_95[563], line_94[561], line_93[559], line_92[557], line_91[555], line_90[553], line_89[551], line_88[549], line_87[547], line_86[545], line_85[543], line_84[541], line_83[539], line_82[537], line_81[535], line_80[533], line_79[531], line_78[529], line_77[527], line_76[525], line_75[523], line_74[521], line_73[519], line_72[517], line_71[515], line_70[513], line_69[511], line_68[509], line_67[507], line_66[505], line_65[503], line_64[501], line_63[499], line_62[497], line_61[495], line_60[493], line_59[491], line_58[489], line_57[487], line_56[485], line_55[483], line_54[481], line_53[479], line_52[477], line_51[475], line_50[473], line_49[471], line_48[469], line_47[467], line_46[465], line_45[463], line_44[461], line_43[459], line_42[457], line_41[455], line_40[453], line_39[451], line_38[449], line_37[447], line_36[445], line_35[443], line_34[441], line_33[439], line_32[437], line_31[435], line_30[433], line_29[431], line_28[429], line_27[427], line_26[425], line_25[423], line_24[421], line_23[419], line_22[417], line_21[415], line_20[413], line_19[411], line_18[409], line_17[407], line_16[405], line_15[403], line_14[401], line_13[399], line_12[397], line_11[395], line_10[393], line_9[391], line_8[389], line_7[387], line_6[385], line_5[383], line_4[381], line_3[379], line_2[377], line_1[375] };
assign col_630 = {line_128[630], line_127[628], line_126[626], line_125[624], line_124[622], line_123[620], line_122[618], line_121[616], line_120[614], line_119[612], line_118[610], line_117[608], line_116[606], line_115[604], line_114[602], line_113[600], line_112[598], line_111[596], line_110[594], line_109[592], line_108[590], line_107[588], line_106[586], line_105[584], line_104[582], line_103[580], line_102[578], line_101[576], line_100[574], line_99[572], line_98[570], line_97[568], line_96[566], line_95[564], line_94[562], line_93[560], line_92[558], line_91[556], line_90[554], line_89[552], line_88[550], line_87[548], line_86[546], line_85[544], line_84[542], line_83[540], line_82[538], line_81[536], line_80[534], line_79[532], line_78[530], line_77[528], line_76[526], line_75[524], line_74[522], line_73[520], line_72[518], line_71[516], line_70[514], line_69[512], line_68[510], line_67[508], line_66[506], line_65[504], line_64[502], line_63[500], line_62[498], line_61[496], line_60[494], line_59[492], line_58[490], line_57[488], line_56[486], line_55[484], line_54[482], line_53[480], line_52[478], line_51[476], line_50[474], line_49[472], line_48[470], line_47[468], line_46[466], line_45[464], line_44[462], line_43[460], line_42[458], line_41[456], line_40[454], line_39[452], line_38[450], line_37[448], line_36[446], line_35[444], line_34[442], line_33[440], line_32[438], line_31[436], line_30[434], line_29[432], line_28[430], line_27[428], line_26[426], line_25[424], line_24[422], line_23[420], line_22[418], line_21[416], line_20[414], line_19[412], line_18[410], line_17[408], line_16[406], line_15[404], line_14[402], line_13[400], line_12[398], line_11[396], line_10[394], line_9[392], line_8[390], line_7[388], line_6[386], line_5[384], line_4[382], line_3[380], line_2[378], line_1[376] };
assign col_631 = {line_128[631], line_127[629], line_126[627], line_125[625], line_124[623], line_123[621], line_122[619], line_121[617], line_120[615], line_119[613], line_118[611], line_117[609], line_116[607], line_115[605], line_114[603], line_113[601], line_112[599], line_111[597], line_110[595], line_109[593], line_108[591], line_107[589], line_106[587], line_105[585], line_104[583], line_103[581], line_102[579], line_101[577], line_100[575], line_99[573], line_98[571], line_97[569], line_96[567], line_95[565], line_94[563], line_93[561], line_92[559], line_91[557], line_90[555], line_89[553], line_88[551], line_87[549], line_86[547], line_85[545], line_84[543], line_83[541], line_82[539], line_81[537], line_80[535], line_79[533], line_78[531], line_77[529], line_76[527], line_75[525], line_74[523], line_73[521], line_72[519], line_71[517], line_70[515], line_69[513], line_68[511], line_67[509], line_66[507], line_65[505], line_64[503], line_63[501], line_62[499], line_61[497], line_60[495], line_59[493], line_58[491], line_57[489], line_56[487], line_55[485], line_54[483], line_53[481], line_52[479], line_51[477], line_50[475], line_49[473], line_48[471], line_47[469], line_46[467], line_45[465], line_44[463], line_43[461], line_42[459], line_41[457], line_40[455], line_39[453], line_38[451], line_37[449], line_36[447], line_35[445], line_34[443], line_33[441], line_32[439], line_31[437], line_30[435], line_29[433], line_28[431], line_27[429], line_26[427], line_25[425], line_24[423], line_23[421], line_22[419], line_21[417], line_20[415], line_19[413], line_18[411], line_17[409], line_16[407], line_15[405], line_14[403], line_13[401], line_12[399], line_11[397], line_10[395], line_9[393], line_8[391], line_7[389], line_6[387], line_5[385], line_4[383], line_3[381], line_2[379], line_1[377] };
assign col_632 = {line_128[632], line_127[630], line_126[628], line_125[626], line_124[624], line_123[622], line_122[620], line_121[618], line_120[616], line_119[614], line_118[612], line_117[610], line_116[608], line_115[606], line_114[604], line_113[602], line_112[600], line_111[598], line_110[596], line_109[594], line_108[592], line_107[590], line_106[588], line_105[586], line_104[584], line_103[582], line_102[580], line_101[578], line_100[576], line_99[574], line_98[572], line_97[570], line_96[568], line_95[566], line_94[564], line_93[562], line_92[560], line_91[558], line_90[556], line_89[554], line_88[552], line_87[550], line_86[548], line_85[546], line_84[544], line_83[542], line_82[540], line_81[538], line_80[536], line_79[534], line_78[532], line_77[530], line_76[528], line_75[526], line_74[524], line_73[522], line_72[520], line_71[518], line_70[516], line_69[514], line_68[512], line_67[510], line_66[508], line_65[506], line_64[504], line_63[502], line_62[500], line_61[498], line_60[496], line_59[494], line_58[492], line_57[490], line_56[488], line_55[486], line_54[484], line_53[482], line_52[480], line_51[478], line_50[476], line_49[474], line_48[472], line_47[470], line_46[468], line_45[466], line_44[464], line_43[462], line_42[460], line_41[458], line_40[456], line_39[454], line_38[452], line_37[450], line_36[448], line_35[446], line_34[444], line_33[442], line_32[440], line_31[438], line_30[436], line_29[434], line_28[432], line_27[430], line_26[428], line_25[426], line_24[424], line_23[422], line_22[420], line_21[418], line_20[416], line_19[414], line_18[412], line_17[410], line_16[408], line_15[406], line_14[404], line_13[402], line_12[400], line_11[398], line_10[396], line_9[394], line_8[392], line_7[390], line_6[388], line_5[386], line_4[384], line_3[382], line_2[380], line_1[378] };
assign col_633 = {line_128[633], line_127[631], line_126[629], line_125[627], line_124[625], line_123[623], line_122[621], line_121[619], line_120[617], line_119[615], line_118[613], line_117[611], line_116[609], line_115[607], line_114[605], line_113[603], line_112[601], line_111[599], line_110[597], line_109[595], line_108[593], line_107[591], line_106[589], line_105[587], line_104[585], line_103[583], line_102[581], line_101[579], line_100[577], line_99[575], line_98[573], line_97[571], line_96[569], line_95[567], line_94[565], line_93[563], line_92[561], line_91[559], line_90[557], line_89[555], line_88[553], line_87[551], line_86[549], line_85[547], line_84[545], line_83[543], line_82[541], line_81[539], line_80[537], line_79[535], line_78[533], line_77[531], line_76[529], line_75[527], line_74[525], line_73[523], line_72[521], line_71[519], line_70[517], line_69[515], line_68[513], line_67[511], line_66[509], line_65[507], line_64[505], line_63[503], line_62[501], line_61[499], line_60[497], line_59[495], line_58[493], line_57[491], line_56[489], line_55[487], line_54[485], line_53[483], line_52[481], line_51[479], line_50[477], line_49[475], line_48[473], line_47[471], line_46[469], line_45[467], line_44[465], line_43[463], line_42[461], line_41[459], line_40[457], line_39[455], line_38[453], line_37[451], line_36[449], line_35[447], line_34[445], line_33[443], line_32[441], line_31[439], line_30[437], line_29[435], line_28[433], line_27[431], line_26[429], line_25[427], line_24[425], line_23[423], line_22[421], line_21[419], line_20[417], line_19[415], line_18[413], line_17[411], line_16[409], line_15[407], line_14[405], line_13[403], line_12[401], line_11[399], line_10[397], line_9[395], line_8[393], line_7[391], line_6[389], line_5[387], line_4[385], line_3[383], line_2[381], line_1[379] };
assign col_634 = {line_128[634], line_127[632], line_126[630], line_125[628], line_124[626], line_123[624], line_122[622], line_121[620], line_120[618], line_119[616], line_118[614], line_117[612], line_116[610], line_115[608], line_114[606], line_113[604], line_112[602], line_111[600], line_110[598], line_109[596], line_108[594], line_107[592], line_106[590], line_105[588], line_104[586], line_103[584], line_102[582], line_101[580], line_100[578], line_99[576], line_98[574], line_97[572], line_96[570], line_95[568], line_94[566], line_93[564], line_92[562], line_91[560], line_90[558], line_89[556], line_88[554], line_87[552], line_86[550], line_85[548], line_84[546], line_83[544], line_82[542], line_81[540], line_80[538], line_79[536], line_78[534], line_77[532], line_76[530], line_75[528], line_74[526], line_73[524], line_72[522], line_71[520], line_70[518], line_69[516], line_68[514], line_67[512], line_66[510], line_65[508], line_64[506], line_63[504], line_62[502], line_61[500], line_60[498], line_59[496], line_58[494], line_57[492], line_56[490], line_55[488], line_54[486], line_53[484], line_52[482], line_51[480], line_50[478], line_49[476], line_48[474], line_47[472], line_46[470], line_45[468], line_44[466], line_43[464], line_42[462], line_41[460], line_40[458], line_39[456], line_38[454], line_37[452], line_36[450], line_35[448], line_34[446], line_33[444], line_32[442], line_31[440], line_30[438], line_29[436], line_28[434], line_27[432], line_26[430], line_25[428], line_24[426], line_23[424], line_22[422], line_21[420], line_20[418], line_19[416], line_18[414], line_17[412], line_16[410], line_15[408], line_14[406], line_13[404], line_12[402], line_11[400], line_10[398], line_9[396], line_8[394], line_7[392], line_6[390], line_5[388], line_4[386], line_3[384], line_2[382], line_1[380] };
assign col_635 = {line_128[635], line_127[633], line_126[631], line_125[629], line_124[627], line_123[625], line_122[623], line_121[621], line_120[619], line_119[617], line_118[615], line_117[613], line_116[611], line_115[609], line_114[607], line_113[605], line_112[603], line_111[601], line_110[599], line_109[597], line_108[595], line_107[593], line_106[591], line_105[589], line_104[587], line_103[585], line_102[583], line_101[581], line_100[579], line_99[577], line_98[575], line_97[573], line_96[571], line_95[569], line_94[567], line_93[565], line_92[563], line_91[561], line_90[559], line_89[557], line_88[555], line_87[553], line_86[551], line_85[549], line_84[547], line_83[545], line_82[543], line_81[541], line_80[539], line_79[537], line_78[535], line_77[533], line_76[531], line_75[529], line_74[527], line_73[525], line_72[523], line_71[521], line_70[519], line_69[517], line_68[515], line_67[513], line_66[511], line_65[509], line_64[507], line_63[505], line_62[503], line_61[501], line_60[499], line_59[497], line_58[495], line_57[493], line_56[491], line_55[489], line_54[487], line_53[485], line_52[483], line_51[481], line_50[479], line_49[477], line_48[475], line_47[473], line_46[471], line_45[469], line_44[467], line_43[465], line_42[463], line_41[461], line_40[459], line_39[457], line_38[455], line_37[453], line_36[451], line_35[449], line_34[447], line_33[445], line_32[443], line_31[441], line_30[439], line_29[437], line_28[435], line_27[433], line_26[431], line_25[429], line_24[427], line_23[425], line_22[423], line_21[421], line_20[419], line_19[417], line_18[415], line_17[413], line_16[411], line_15[409], line_14[407], line_13[405], line_12[403], line_11[401], line_10[399], line_9[397], line_8[395], line_7[393], line_6[391], line_5[389], line_4[387], line_3[385], line_2[383], line_1[381] };
assign col_636 = {line_128[636], line_127[634], line_126[632], line_125[630], line_124[628], line_123[626], line_122[624], line_121[622], line_120[620], line_119[618], line_118[616], line_117[614], line_116[612], line_115[610], line_114[608], line_113[606], line_112[604], line_111[602], line_110[600], line_109[598], line_108[596], line_107[594], line_106[592], line_105[590], line_104[588], line_103[586], line_102[584], line_101[582], line_100[580], line_99[578], line_98[576], line_97[574], line_96[572], line_95[570], line_94[568], line_93[566], line_92[564], line_91[562], line_90[560], line_89[558], line_88[556], line_87[554], line_86[552], line_85[550], line_84[548], line_83[546], line_82[544], line_81[542], line_80[540], line_79[538], line_78[536], line_77[534], line_76[532], line_75[530], line_74[528], line_73[526], line_72[524], line_71[522], line_70[520], line_69[518], line_68[516], line_67[514], line_66[512], line_65[510], line_64[508], line_63[506], line_62[504], line_61[502], line_60[500], line_59[498], line_58[496], line_57[494], line_56[492], line_55[490], line_54[488], line_53[486], line_52[484], line_51[482], line_50[480], line_49[478], line_48[476], line_47[474], line_46[472], line_45[470], line_44[468], line_43[466], line_42[464], line_41[462], line_40[460], line_39[458], line_38[456], line_37[454], line_36[452], line_35[450], line_34[448], line_33[446], line_32[444], line_31[442], line_30[440], line_29[438], line_28[436], line_27[434], line_26[432], line_25[430], line_24[428], line_23[426], line_22[424], line_21[422], line_20[420], line_19[418], line_18[416], line_17[414], line_16[412], line_15[410], line_14[408], line_13[406], line_12[404], line_11[402], line_10[400], line_9[398], line_8[396], line_7[394], line_6[392], line_5[390], line_4[388], line_3[386], line_2[384], line_1[382] };
assign col_637 = {line_128[637], line_127[635], line_126[633], line_125[631], line_124[629], line_123[627], line_122[625], line_121[623], line_120[621], line_119[619], line_118[617], line_117[615], line_116[613], line_115[611], line_114[609], line_113[607], line_112[605], line_111[603], line_110[601], line_109[599], line_108[597], line_107[595], line_106[593], line_105[591], line_104[589], line_103[587], line_102[585], line_101[583], line_100[581], line_99[579], line_98[577], line_97[575], line_96[573], line_95[571], line_94[569], line_93[567], line_92[565], line_91[563], line_90[561], line_89[559], line_88[557], line_87[555], line_86[553], line_85[551], line_84[549], line_83[547], line_82[545], line_81[543], line_80[541], line_79[539], line_78[537], line_77[535], line_76[533], line_75[531], line_74[529], line_73[527], line_72[525], line_71[523], line_70[521], line_69[519], line_68[517], line_67[515], line_66[513], line_65[511], line_64[509], line_63[507], line_62[505], line_61[503], line_60[501], line_59[499], line_58[497], line_57[495], line_56[493], line_55[491], line_54[489], line_53[487], line_52[485], line_51[483], line_50[481], line_49[479], line_48[477], line_47[475], line_46[473], line_45[471], line_44[469], line_43[467], line_42[465], line_41[463], line_40[461], line_39[459], line_38[457], line_37[455], line_36[453], line_35[451], line_34[449], line_33[447], line_32[445], line_31[443], line_30[441], line_29[439], line_28[437], line_27[435], line_26[433], line_25[431], line_24[429], line_23[427], line_22[425], line_21[423], line_20[421], line_19[419], line_18[417], line_17[415], line_16[413], line_15[411], line_14[409], line_13[407], line_12[405], line_11[403], line_10[401], line_9[399], line_8[397], line_7[395], line_6[393], line_5[391], line_4[389], line_3[387], line_2[385], line_1[383] };
assign col_638 = {line_128[638], line_127[636], line_126[634], line_125[632], line_124[630], line_123[628], line_122[626], line_121[624], line_120[622], line_119[620], line_118[618], line_117[616], line_116[614], line_115[612], line_114[610], line_113[608], line_112[606], line_111[604], line_110[602], line_109[600], line_108[598], line_107[596], line_106[594], line_105[592], line_104[590], line_103[588], line_102[586], line_101[584], line_100[582], line_99[580], line_98[578], line_97[576], line_96[574], line_95[572], line_94[570], line_93[568], line_92[566], line_91[564], line_90[562], line_89[560], line_88[558], line_87[556], line_86[554], line_85[552], line_84[550], line_83[548], line_82[546], line_81[544], line_80[542], line_79[540], line_78[538], line_77[536], line_76[534], line_75[532], line_74[530], line_73[528], line_72[526], line_71[524], line_70[522], line_69[520], line_68[518], line_67[516], line_66[514], line_65[512], line_64[510], line_63[508], line_62[506], line_61[504], line_60[502], line_59[500], line_58[498], line_57[496], line_56[494], line_55[492], line_54[490], line_53[488], line_52[486], line_51[484], line_50[482], line_49[480], line_48[478], line_47[476], line_46[474], line_45[472], line_44[470], line_43[468], line_42[466], line_41[464], line_40[462], line_39[460], line_38[458], line_37[456], line_36[454], line_35[452], line_34[450], line_33[448], line_32[446], line_31[444], line_30[442], line_29[440], line_28[438], line_27[436], line_26[434], line_25[432], line_24[430], line_23[428], line_22[426], line_21[424], line_20[422], line_19[420], line_18[418], line_17[416], line_16[414], line_15[412], line_14[410], line_13[408], line_12[406], line_11[404], line_10[402], line_9[400], line_8[398], line_7[396], line_6[394], line_5[392], line_4[390], line_3[388], line_2[386], line_1[384] };
assign col_639 = {line_128[639], line_127[637], line_126[635], line_125[633], line_124[631], line_123[629], line_122[627], line_121[625], line_120[623], line_119[621], line_118[619], line_117[617], line_116[615], line_115[613], line_114[611], line_113[609], line_112[607], line_111[605], line_110[603], line_109[601], line_108[599], line_107[597], line_106[595], line_105[593], line_104[591], line_103[589], line_102[587], line_101[585], line_100[583], line_99[581], line_98[579], line_97[577], line_96[575], line_95[573], line_94[571], line_93[569], line_92[567], line_91[565], line_90[563], line_89[561], line_88[559], line_87[557], line_86[555], line_85[553], line_84[551], line_83[549], line_82[547], line_81[545], line_80[543], line_79[541], line_78[539], line_77[537], line_76[535], line_75[533], line_74[531], line_73[529], line_72[527], line_71[525], line_70[523], line_69[521], line_68[519], line_67[517], line_66[515], line_65[513], line_64[511], line_63[509], line_62[507], line_61[505], line_60[503], line_59[501], line_58[499], line_57[497], line_56[495], line_55[493], line_54[491], line_53[489], line_52[487], line_51[485], line_50[483], line_49[481], line_48[479], line_47[477], line_46[475], line_45[473], line_44[471], line_43[469], line_42[467], line_41[465], line_40[463], line_39[461], line_38[459], line_37[457], line_36[455], line_35[453], line_34[451], line_33[449], line_32[447], line_31[445], line_30[443], line_29[441], line_28[439], line_27[437], line_26[435], line_25[433], line_24[431], line_23[429], line_22[427], line_21[425], line_20[423], line_19[421], line_18[419], line_17[417], line_16[415], line_15[413], line_14[411], line_13[409], line_12[407], line_11[405], line_10[403], line_9[401], line_8[399], line_7[397], line_6[395], line_5[393], line_4[391], line_3[389], line_2[387], line_1[385] };
assign col_640 = {line_128[640], line_127[638], line_126[636], line_125[634], line_124[632], line_123[630], line_122[628], line_121[626], line_120[624], line_119[622], line_118[620], line_117[618], line_116[616], line_115[614], line_114[612], line_113[610], line_112[608], line_111[606], line_110[604], line_109[602], line_108[600], line_107[598], line_106[596], line_105[594], line_104[592], line_103[590], line_102[588], line_101[586], line_100[584], line_99[582], line_98[580], line_97[578], line_96[576], line_95[574], line_94[572], line_93[570], line_92[568], line_91[566], line_90[564], line_89[562], line_88[560], line_87[558], line_86[556], line_85[554], line_84[552], line_83[550], line_82[548], line_81[546], line_80[544], line_79[542], line_78[540], line_77[538], line_76[536], line_75[534], line_74[532], line_73[530], line_72[528], line_71[526], line_70[524], line_69[522], line_68[520], line_67[518], line_66[516], line_65[514], line_64[512], line_63[510], line_62[508], line_61[506], line_60[504], line_59[502], line_58[500], line_57[498], line_56[496], line_55[494], line_54[492], line_53[490], line_52[488], line_51[486], line_50[484], line_49[482], line_48[480], line_47[478], line_46[476], line_45[474], line_44[472], line_43[470], line_42[468], line_41[466], line_40[464], line_39[462], line_38[460], line_37[458], line_36[456], line_35[454], line_34[452], line_33[450], line_32[448], line_31[446], line_30[444], line_29[442], line_28[440], line_27[438], line_26[436], line_25[434], line_24[432], line_23[430], line_22[428], line_21[426], line_20[424], line_19[422], line_18[420], line_17[418], line_16[416], line_15[414], line_14[412], line_13[410], line_12[408], line_11[406], line_10[404], line_9[402], line_8[400], line_7[398], line_6[396], line_5[394], line_4[392], line_3[390], line_2[388], line_1[386] };
assign col_641 = {line_128[641], line_127[639], line_126[637], line_125[635], line_124[633], line_123[631], line_122[629], line_121[627], line_120[625], line_119[623], line_118[621], line_117[619], line_116[617], line_115[615], line_114[613], line_113[611], line_112[609], line_111[607], line_110[605], line_109[603], line_108[601], line_107[599], line_106[597], line_105[595], line_104[593], line_103[591], line_102[589], line_101[587], line_100[585], line_99[583], line_98[581], line_97[579], line_96[577], line_95[575], line_94[573], line_93[571], line_92[569], line_91[567], line_90[565], line_89[563], line_88[561], line_87[559], line_86[557], line_85[555], line_84[553], line_83[551], line_82[549], line_81[547], line_80[545], line_79[543], line_78[541], line_77[539], line_76[537], line_75[535], line_74[533], line_73[531], line_72[529], line_71[527], line_70[525], line_69[523], line_68[521], line_67[519], line_66[517], line_65[515], line_64[513], line_63[511], line_62[509], line_61[507], line_60[505], line_59[503], line_58[501], line_57[499], line_56[497], line_55[495], line_54[493], line_53[491], line_52[489], line_51[487], line_50[485], line_49[483], line_48[481], line_47[479], line_46[477], line_45[475], line_44[473], line_43[471], line_42[469], line_41[467], line_40[465], line_39[463], line_38[461], line_37[459], line_36[457], line_35[455], line_34[453], line_33[451], line_32[449], line_31[447], line_30[445], line_29[443], line_28[441], line_27[439], line_26[437], line_25[435], line_24[433], line_23[431], line_22[429], line_21[427], line_20[425], line_19[423], line_18[421], line_17[419], line_16[417], line_15[415], line_14[413], line_13[411], line_12[409], line_11[407], line_10[405], line_9[403], line_8[401], line_7[399], line_6[397], line_5[395], line_4[393], line_3[391], line_2[389], line_1[387] };
assign col_642 = {line_128[642], line_127[640], line_126[638], line_125[636], line_124[634], line_123[632], line_122[630], line_121[628], line_120[626], line_119[624], line_118[622], line_117[620], line_116[618], line_115[616], line_114[614], line_113[612], line_112[610], line_111[608], line_110[606], line_109[604], line_108[602], line_107[600], line_106[598], line_105[596], line_104[594], line_103[592], line_102[590], line_101[588], line_100[586], line_99[584], line_98[582], line_97[580], line_96[578], line_95[576], line_94[574], line_93[572], line_92[570], line_91[568], line_90[566], line_89[564], line_88[562], line_87[560], line_86[558], line_85[556], line_84[554], line_83[552], line_82[550], line_81[548], line_80[546], line_79[544], line_78[542], line_77[540], line_76[538], line_75[536], line_74[534], line_73[532], line_72[530], line_71[528], line_70[526], line_69[524], line_68[522], line_67[520], line_66[518], line_65[516], line_64[514], line_63[512], line_62[510], line_61[508], line_60[506], line_59[504], line_58[502], line_57[500], line_56[498], line_55[496], line_54[494], line_53[492], line_52[490], line_51[488], line_50[486], line_49[484], line_48[482], line_47[480], line_46[478], line_45[476], line_44[474], line_43[472], line_42[470], line_41[468], line_40[466], line_39[464], line_38[462], line_37[460], line_36[458], line_35[456], line_34[454], line_33[452], line_32[450], line_31[448], line_30[446], line_29[444], line_28[442], line_27[440], line_26[438], line_25[436], line_24[434], line_23[432], line_22[430], line_21[428], line_20[426], line_19[424], line_18[422], line_17[420], line_16[418], line_15[416], line_14[414], line_13[412], line_12[410], line_11[408], line_10[406], line_9[404], line_8[402], line_7[400], line_6[398], line_5[396], line_4[394], line_3[392], line_2[390], line_1[388] };
assign col_643 = {line_128[643], line_127[641], line_126[639], line_125[637], line_124[635], line_123[633], line_122[631], line_121[629], line_120[627], line_119[625], line_118[623], line_117[621], line_116[619], line_115[617], line_114[615], line_113[613], line_112[611], line_111[609], line_110[607], line_109[605], line_108[603], line_107[601], line_106[599], line_105[597], line_104[595], line_103[593], line_102[591], line_101[589], line_100[587], line_99[585], line_98[583], line_97[581], line_96[579], line_95[577], line_94[575], line_93[573], line_92[571], line_91[569], line_90[567], line_89[565], line_88[563], line_87[561], line_86[559], line_85[557], line_84[555], line_83[553], line_82[551], line_81[549], line_80[547], line_79[545], line_78[543], line_77[541], line_76[539], line_75[537], line_74[535], line_73[533], line_72[531], line_71[529], line_70[527], line_69[525], line_68[523], line_67[521], line_66[519], line_65[517], line_64[515], line_63[513], line_62[511], line_61[509], line_60[507], line_59[505], line_58[503], line_57[501], line_56[499], line_55[497], line_54[495], line_53[493], line_52[491], line_51[489], line_50[487], line_49[485], line_48[483], line_47[481], line_46[479], line_45[477], line_44[475], line_43[473], line_42[471], line_41[469], line_40[467], line_39[465], line_38[463], line_37[461], line_36[459], line_35[457], line_34[455], line_33[453], line_32[451], line_31[449], line_30[447], line_29[445], line_28[443], line_27[441], line_26[439], line_25[437], line_24[435], line_23[433], line_22[431], line_21[429], line_20[427], line_19[425], line_18[423], line_17[421], line_16[419], line_15[417], line_14[415], line_13[413], line_12[411], line_11[409], line_10[407], line_9[405], line_8[403], line_7[401], line_6[399], line_5[397], line_4[395], line_3[393], line_2[391], line_1[389] };
assign col_644 = {line_128[644], line_127[642], line_126[640], line_125[638], line_124[636], line_123[634], line_122[632], line_121[630], line_120[628], line_119[626], line_118[624], line_117[622], line_116[620], line_115[618], line_114[616], line_113[614], line_112[612], line_111[610], line_110[608], line_109[606], line_108[604], line_107[602], line_106[600], line_105[598], line_104[596], line_103[594], line_102[592], line_101[590], line_100[588], line_99[586], line_98[584], line_97[582], line_96[580], line_95[578], line_94[576], line_93[574], line_92[572], line_91[570], line_90[568], line_89[566], line_88[564], line_87[562], line_86[560], line_85[558], line_84[556], line_83[554], line_82[552], line_81[550], line_80[548], line_79[546], line_78[544], line_77[542], line_76[540], line_75[538], line_74[536], line_73[534], line_72[532], line_71[530], line_70[528], line_69[526], line_68[524], line_67[522], line_66[520], line_65[518], line_64[516], line_63[514], line_62[512], line_61[510], line_60[508], line_59[506], line_58[504], line_57[502], line_56[500], line_55[498], line_54[496], line_53[494], line_52[492], line_51[490], line_50[488], line_49[486], line_48[484], line_47[482], line_46[480], line_45[478], line_44[476], line_43[474], line_42[472], line_41[470], line_40[468], line_39[466], line_38[464], line_37[462], line_36[460], line_35[458], line_34[456], line_33[454], line_32[452], line_31[450], line_30[448], line_29[446], line_28[444], line_27[442], line_26[440], line_25[438], line_24[436], line_23[434], line_22[432], line_21[430], line_20[428], line_19[426], line_18[424], line_17[422], line_16[420], line_15[418], line_14[416], line_13[414], line_12[412], line_11[410], line_10[408], line_9[406], line_8[404], line_7[402], line_6[400], line_5[398], line_4[396], line_3[394], line_2[392], line_1[390] };
assign col_645 = {line_128[645], line_127[643], line_126[641], line_125[639], line_124[637], line_123[635], line_122[633], line_121[631], line_120[629], line_119[627], line_118[625], line_117[623], line_116[621], line_115[619], line_114[617], line_113[615], line_112[613], line_111[611], line_110[609], line_109[607], line_108[605], line_107[603], line_106[601], line_105[599], line_104[597], line_103[595], line_102[593], line_101[591], line_100[589], line_99[587], line_98[585], line_97[583], line_96[581], line_95[579], line_94[577], line_93[575], line_92[573], line_91[571], line_90[569], line_89[567], line_88[565], line_87[563], line_86[561], line_85[559], line_84[557], line_83[555], line_82[553], line_81[551], line_80[549], line_79[547], line_78[545], line_77[543], line_76[541], line_75[539], line_74[537], line_73[535], line_72[533], line_71[531], line_70[529], line_69[527], line_68[525], line_67[523], line_66[521], line_65[519], line_64[517], line_63[515], line_62[513], line_61[511], line_60[509], line_59[507], line_58[505], line_57[503], line_56[501], line_55[499], line_54[497], line_53[495], line_52[493], line_51[491], line_50[489], line_49[487], line_48[485], line_47[483], line_46[481], line_45[479], line_44[477], line_43[475], line_42[473], line_41[471], line_40[469], line_39[467], line_38[465], line_37[463], line_36[461], line_35[459], line_34[457], line_33[455], line_32[453], line_31[451], line_30[449], line_29[447], line_28[445], line_27[443], line_26[441], line_25[439], line_24[437], line_23[435], line_22[433], line_21[431], line_20[429], line_19[427], line_18[425], line_17[423], line_16[421], line_15[419], line_14[417], line_13[415], line_12[413], line_11[411], line_10[409], line_9[407], line_8[405], line_7[403], line_6[401], line_5[399], line_4[397], line_3[395], line_2[393], line_1[391] };
assign col_646 = {line_128[646], line_127[644], line_126[642], line_125[640], line_124[638], line_123[636], line_122[634], line_121[632], line_120[630], line_119[628], line_118[626], line_117[624], line_116[622], line_115[620], line_114[618], line_113[616], line_112[614], line_111[612], line_110[610], line_109[608], line_108[606], line_107[604], line_106[602], line_105[600], line_104[598], line_103[596], line_102[594], line_101[592], line_100[590], line_99[588], line_98[586], line_97[584], line_96[582], line_95[580], line_94[578], line_93[576], line_92[574], line_91[572], line_90[570], line_89[568], line_88[566], line_87[564], line_86[562], line_85[560], line_84[558], line_83[556], line_82[554], line_81[552], line_80[550], line_79[548], line_78[546], line_77[544], line_76[542], line_75[540], line_74[538], line_73[536], line_72[534], line_71[532], line_70[530], line_69[528], line_68[526], line_67[524], line_66[522], line_65[520], line_64[518], line_63[516], line_62[514], line_61[512], line_60[510], line_59[508], line_58[506], line_57[504], line_56[502], line_55[500], line_54[498], line_53[496], line_52[494], line_51[492], line_50[490], line_49[488], line_48[486], line_47[484], line_46[482], line_45[480], line_44[478], line_43[476], line_42[474], line_41[472], line_40[470], line_39[468], line_38[466], line_37[464], line_36[462], line_35[460], line_34[458], line_33[456], line_32[454], line_31[452], line_30[450], line_29[448], line_28[446], line_27[444], line_26[442], line_25[440], line_24[438], line_23[436], line_22[434], line_21[432], line_20[430], line_19[428], line_18[426], line_17[424], line_16[422], line_15[420], line_14[418], line_13[416], line_12[414], line_11[412], line_10[410], line_9[408], line_8[406], line_7[404], line_6[402], line_5[400], line_4[398], line_3[396], line_2[394], line_1[392] };
assign col_647 = {line_128[647], line_127[645], line_126[643], line_125[641], line_124[639], line_123[637], line_122[635], line_121[633], line_120[631], line_119[629], line_118[627], line_117[625], line_116[623], line_115[621], line_114[619], line_113[617], line_112[615], line_111[613], line_110[611], line_109[609], line_108[607], line_107[605], line_106[603], line_105[601], line_104[599], line_103[597], line_102[595], line_101[593], line_100[591], line_99[589], line_98[587], line_97[585], line_96[583], line_95[581], line_94[579], line_93[577], line_92[575], line_91[573], line_90[571], line_89[569], line_88[567], line_87[565], line_86[563], line_85[561], line_84[559], line_83[557], line_82[555], line_81[553], line_80[551], line_79[549], line_78[547], line_77[545], line_76[543], line_75[541], line_74[539], line_73[537], line_72[535], line_71[533], line_70[531], line_69[529], line_68[527], line_67[525], line_66[523], line_65[521], line_64[519], line_63[517], line_62[515], line_61[513], line_60[511], line_59[509], line_58[507], line_57[505], line_56[503], line_55[501], line_54[499], line_53[497], line_52[495], line_51[493], line_50[491], line_49[489], line_48[487], line_47[485], line_46[483], line_45[481], line_44[479], line_43[477], line_42[475], line_41[473], line_40[471], line_39[469], line_38[467], line_37[465], line_36[463], line_35[461], line_34[459], line_33[457], line_32[455], line_31[453], line_30[451], line_29[449], line_28[447], line_27[445], line_26[443], line_25[441], line_24[439], line_23[437], line_22[435], line_21[433], line_20[431], line_19[429], line_18[427], line_17[425], line_16[423], line_15[421], line_14[419], line_13[417], line_12[415], line_11[413], line_10[411], line_9[409], line_8[407], line_7[405], line_6[403], line_5[401], line_4[399], line_3[397], line_2[395], line_1[393] };
assign col_648 = {line_128[648], line_127[646], line_126[644], line_125[642], line_124[640], line_123[638], line_122[636], line_121[634], line_120[632], line_119[630], line_118[628], line_117[626], line_116[624], line_115[622], line_114[620], line_113[618], line_112[616], line_111[614], line_110[612], line_109[610], line_108[608], line_107[606], line_106[604], line_105[602], line_104[600], line_103[598], line_102[596], line_101[594], line_100[592], line_99[590], line_98[588], line_97[586], line_96[584], line_95[582], line_94[580], line_93[578], line_92[576], line_91[574], line_90[572], line_89[570], line_88[568], line_87[566], line_86[564], line_85[562], line_84[560], line_83[558], line_82[556], line_81[554], line_80[552], line_79[550], line_78[548], line_77[546], line_76[544], line_75[542], line_74[540], line_73[538], line_72[536], line_71[534], line_70[532], line_69[530], line_68[528], line_67[526], line_66[524], line_65[522], line_64[520], line_63[518], line_62[516], line_61[514], line_60[512], line_59[510], line_58[508], line_57[506], line_56[504], line_55[502], line_54[500], line_53[498], line_52[496], line_51[494], line_50[492], line_49[490], line_48[488], line_47[486], line_46[484], line_45[482], line_44[480], line_43[478], line_42[476], line_41[474], line_40[472], line_39[470], line_38[468], line_37[466], line_36[464], line_35[462], line_34[460], line_33[458], line_32[456], line_31[454], line_30[452], line_29[450], line_28[448], line_27[446], line_26[444], line_25[442], line_24[440], line_23[438], line_22[436], line_21[434], line_20[432], line_19[430], line_18[428], line_17[426], line_16[424], line_15[422], line_14[420], line_13[418], line_12[416], line_11[414], line_10[412], line_9[410], line_8[408], line_7[406], line_6[404], line_5[402], line_4[400], line_3[398], line_2[396], line_1[394] };
assign col_649 = {line_128[649], line_127[647], line_126[645], line_125[643], line_124[641], line_123[639], line_122[637], line_121[635], line_120[633], line_119[631], line_118[629], line_117[627], line_116[625], line_115[623], line_114[621], line_113[619], line_112[617], line_111[615], line_110[613], line_109[611], line_108[609], line_107[607], line_106[605], line_105[603], line_104[601], line_103[599], line_102[597], line_101[595], line_100[593], line_99[591], line_98[589], line_97[587], line_96[585], line_95[583], line_94[581], line_93[579], line_92[577], line_91[575], line_90[573], line_89[571], line_88[569], line_87[567], line_86[565], line_85[563], line_84[561], line_83[559], line_82[557], line_81[555], line_80[553], line_79[551], line_78[549], line_77[547], line_76[545], line_75[543], line_74[541], line_73[539], line_72[537], line_71[535], line_70[533], line_69[531], line_68[529], line_67[527], line_66[525], line_65[523], line_64[521], line_63[519], line_62[517], line_61[515], line_60[513], line_59[511], line_58[509], line_57[507], line_56[505], line_55[503], line_54[501], line_53[499], line_52[497], line_51[495], line_50[493], line_49[491], line_48[489], line_47[487], line_46[485], line_45[483], line_44[481], line_43[479], line_42[477], line_41[475], line_40[473], line_39[471], line_38[469], line_37[467], line_36[465], line_35[463], line_34[461], line_33[459], line_32[457], line_31[455], line_30[453], line_29[451], line_28[449], line_27[447], line_26[445], line_25[443], line_24[441], line_23[439], line_22[437], line_21[435], line_20[433], line_19[431], line_18[429], line_17[427], line_16[425], line_15[423], line_14[421], line_13[419], line_12[417], line_11[415], line_10[413], line_9[411], line_8[409], line_7[407], line_6[405], line_5[403], line_4[401], line_3[399], line_2[397], line_1[395] };
assign col_650 = {line_128[650], line_127[648], line_126[646], line_125[644], line_124[642], line_123[640], line_122[638], line_121[636], line_120[634], line_119[632], line_118[630], line_117[628], line_116[626], line_115[624], line_114[622], line_113[620], line_112[618], line_111[616], line_110[614], line_109[612], line_108[610], line_107[608], line_106[606], line_105[604], line_104[602], line_103[600], line_102[598], line_101[596], line_100[594], line_99[592], line_98[590], line_97[588], line_96[586], line_95[584], line_94[582], line_93[580], line_92[578], line_91[576], line_90[574], line_89[572], line_88[570], line_87[568], line_86[566], line_85[564], line_84[562], line_83[560], line_82[558], line_81[556], line_80[554], line_79[552], line_78[550], line_77[548], line_76[546], line_75[544], line_74[542], line_73[540], line_72[538], line_71[536], line_70[534], line_69[532], line_68[530], line_67[528], line_66[526], line_65[524], line_64[522], line_63[520], line_62[518], line_61[516], line_60[514], line_59[512], line_58[510], line_57[508], line_56[506], line_55[504], line_54[502], line_53[500], line_52[498], line_51[496], line_50[494], line_49[492], line_48[490], line_47[488], line_46[486], line_45[484], line_44[482], line_43[480], line_42[478], line_41[476], line_40[474], line_39[472], line_38[470], line_37[468], line_36[466], line_35[464], line_34[462], line_33[460], line_32[458], line_31[456], line_30[454], line_29[452], line_28[450], line_27[448], line_26[446], line_25[444], line_24[442], line_23[440], line_22[438], line_21[436], line_20[434], line_19[432], line_18[430], line_17[428], line_16[426], line_15[424], line_14[422], line_13[420], line_12[418], line_11[416], line_10[414], line_9[412], line_8[410], line_7[408], line_6[406], line_5[404], line_4[402], line_3[400], line_2[398], line_1[396] };
assign col_651 = {line_128[651], line_127[649], line_126[647], line_125[645], line_124[643], line_123[641], line_122[639], line_121[637], line_120[635], line_119[633], line_118[631], line_117[629], line_116[627], line_115[625], line_114[623], line_113[621], line_112[619], line_111[617], line_110[615], line_109[613], line_108[611], line_107[609], line_106[607], line_105[605], line_104[603], line_103[601], line_102[599], line_101[597], line_100[595], line_99[593], line_98[591], line_97[589], line_96[587], line_95[585], line_94[583], line_93[581], line_92[579], line_91[577], line_90[575], line_89[573], line_88[571], line_87[569], line_86[567], line_85[565], line_84[563], line_83[561], line_82[559], line_81[557], line_80[555], line_79[553], line_78[551], line_77[549], line_76[547], line_75[545], line_74[543], line_73[541], line_72[539], line_71[537], line_70[535], line_69[533], line_68[531], line_67[529], line_66[527], line_65[525], line_64[523], line_63[521], line_62[519], line_61[517], line_60[515], line_59[513], line_58[511], line_57[509], line_56[507], line_55[505], line_54[503], line_53[501], line_52[499], line_51[497], line_50[495], line_49[493], line_48[491], line_47[489], line_46[487], line_45[485], line_44[483], line_43[481], line_42[479], line_41[477], line_40[475], line_39[473], line_38[471], line_37[469], line_36[467], line_35[465], line_34[463], line_33[461], line_32[459], line_31[457], line_30[455], line_29[453], line_28[451], line_27[449], line_26[447], line_25[445], line_24[443], line_23[441], line_22[439], line_21[437], line_20[435], line_19[433], line_18[431], line_17[429], line_16[427], line_15[425], line_14[423], line_13[421], line_12[419], line_11[417], line_10[415], line_9[413], line_8[411], line_7[409], line_6[407], line_5[405], line_4[403], line_3[401], line_2[399], line_1[397] };
assign col_652 = {line_128[652], line_127[650], line_126[648], line_125[646], line_124[644], line_123[642], line_122[640], line_121[638], line_120[636], line_119[634], line_118[632], line_117[630], line_116[628], line_115[626], line_114[624], line_113[622], line_112[620], line_111[618], line_110[616], line_109[614], line_108[612], line_107[610], line_106[608], line_105[606], line_104[604], line_103[602], line_102[600], line_101[598], line_100[596], line_99[594], line_98[592], line_97[590], line_96[588], line_95[586], line_94[584], line_93[582], line_92[580], line_91[578], line_90[576], line_89[574], line_88[572], line_87[570], line_86[568], line_85[566], line_84[564], line_83[562], line_82[560], line_81[558], line_80[556], line_79[554], line_78[552], line_77[550], line_76[548], line_75[546], line_74[544], line_73[542], line_72[540], line_71[538], line_70[536], line_69[534], line_68[532], line_67[530], line_66[528], line_65[526], line_64[524], line_63[522], line_62[520], line_61[518], line_60[516], line_59[514], line_58[512], line_57[510], line_56[508], line_55[506], line_54[504], line_53[502], line_52[500], line_51[498], line_50[496], line_49[494], line_48[492], line_47[490], line_46[488], line_45[486], line_44[484], line_43[482], line_42[480], line_41[478], line_40[476], line_39[474], line_38[472], line_37[470], line_36[468], line_35[466], line_34[464], line_33[462], line_32[460], line_31[458], line_30[456], line_29[454], line_28[452], line_27[450], line_26[448], line_25[446], line_24[444], line_23[442], line_22[440], line_21[438], line_20[436], line_19[434], line_18[432], line_17[430], line_16[428], line_15[426], line_14[424], line_13[422], line_12[420], line_11[418], line_10[416], line_9[414], line_8[412], line_7[410], line_6[408], line_5[406], line_4[404], line_3[402], line_2[400], line_1[398] };
assign col_653 = {line_128[653], line_127[651], line_126[649], line_125[647], line_124[645], line_123[643], line_122[641], line_121[639], line_120[637], line_119[635], line_118[633], line_117[631], line_116[629], line_115[627], line_114[625], line_113[623], line_112[621], line_111[619], line_110[617], line_109[615], line_108[613], line_107[611], line_106[609], line_105[607], line_104[605], line_103[603], line_102[601], line_101[599], line_100[597], line_99[595], line_98[593], line_97[591], line_96[589], line_95[587], line_94[585], line_93[583], line_92[581], line_91[579], line_90[577], line_89[575], line_88[573], line_87[571], line_86[569], line_85[567], line_84[565], line_83[563], line_82[561], line_81[559], line_80[557], line_79[555], line_78[553], line_77[551], line_76[549], line_75[547], line_74[545], line_73[543], line_72[541], line_71[539], line_70[537], line_69[535], line_68[533], line_67[531], line_66[529], line_65[527], line_64[525], line_63[523], line_62[521], line_61[519], line_60[517], line_59[515], line_58[513], line_57[511], line_56[509], line_55[507], line_54[505], line_53[503], line_52[501], line_51[499], line_50[497], line_49[495], line_48[493], line_47[491], line_46[489], line_45[487], line_44[485], line_43[483], line_42[481], line_41[479], line_40[477], line_39[475], line_38[473], line_37[471], line_36[469], line_35[467], line_34[465], line_33[463], line_32[461], line_31[459], line_30[457], line_29[455], line_28[453], line_27[451], line_26[449], line_25[447], line_24[445], line_23[443], line_22[441], line_21[439], line_20[437], line_19[435], line_18[433], line_17[431], line_16[429], line_15[427], line_14[425], line_13[423], line_12[421], line_11[419], line_10[417], line_9[415], line_8[413], line_7[411], line_6[409], line_5[407], line_4[405], line_3[403], line_2[401], line_1[399] };
assign col_654 = {line_128[654], line_127[652], line_126[650], line_125[648], line_124[646], line_123[644], line_122[642], line_121[640], line_120[638], line_119[636], line_118[634], line_117[632], line_116[630], line_115[628], line_114[626], line_113[624], line_112[622], line_111[620], line_110[618], line_109[616], line_108[614], line_107[612], line_106[610], line_105[608], line_104[606], line_103[604], line_102[602], line_101[600], line_100[598], line_99[596], line_98[594], line_97[592], line_96[590], line_95[588], line_94[586], line_93[584], line_92[582], line_91[580], line_90[578], line_89[576], line_88[574], line_87[572], line_86[570], line_85[568], line_84[566], line_83[564], line_82[562], line_81[560], line_80[558], line_79[556], line_78[554], line_77[552], line_76[550], line_75[548], line_74[546], line_73[544], line_72[542], line_71[540], line_70[538], line_69[536], line_68[534], line_67[532], line_66[530], line_65[528], line_64[526], line_63[524], line_62[522], line_61[520], line_60[518], line_59[516], line_58[514], line_57[512], line_56[510], line_55[508], line_54[506], line_53[504], line_52[502], line_51[500], line_50[498], line_49[496], line_48[494], line_47[492], line_46[490], line_45[488], line_44[486], line_43[484], line_42[482], line_41[480], line_40[478], line_39[476], line_38[474], line_37[472], line_36[470], line_35[468], line_34[466], line_33[464], line_32[462], line_31[460], line_30[458], line_29[456], line_28[454], line_27[452], line_26[450], line_25[448], line_24[446], line_23[444], line_22[442], line_21[440], line_20[438], line_19[436], line_18[434], line_17[432], line_16[430], line_15[428], line_14[426], line_13[424], line_12[422], line_11[420], line_10[418], line_9[416], line_8[414], line_7[412], line_6[410], line_5[408], line_4[406], line_3[404], line_2[402], line_1[400] };
assign col_655 = {line_128[655], line_127[653], line_126[651], line_125[649], line_124[647], line_123[645], line_122[643], line_121[641], line_120[639], line_119[637], line_118[635], line_117[633], line_116[631], line_115[629], line_114[627], line_113[625], line_112[623], line_111[621], line_110[619], line_109[617], line_108[615], line_107[613], line_106[611], line_105[609], line_104[607], line_103[605], line_102[603], line_101[601], line_100[599], line_99[597], line_98[595], line_97[593], line_96[591], line_95[589], line_94[587], line_93[585], line_92[583], line_91[581], line_90[579], line_89[577], line_88[575], line_87[573], line_86[571], line_85[569], line_84[567], line_83[565], line_82[563], line_81[561], line_80[559], line_79[557], line_78[555], line_77[553], line_76[551], line_75[549], line_74[547], line_73[545], line_72[543], line_71[541], line_70[539], line_69[537], line_68[535], line_67[533], line_66[531], line_65[529], line_64[527], line_63[525], line_62[523], line_61[521], line_60[519], line_59[517], line_58[515], line_57[513], line_56[511], line_55[509], line_54[507], line_53[505], line_52[503], line_51[501], line_50[499], line_49[497], line_48[495], line_47[493], line_46[491], line_45[489], line_44[487], line_43[485], line_42[483], line_41[481], line_40[479], line_39[477], line_38[475], line_37[473], line_36[471], line_35[469], line_34[467], line_33[465], line_32[463], line_31[461], line_30[459], line_29[457], line_28[455], line_27[453], line_26[451], line_25[449], line_24[447], line_23[445], line_22[443], line_21[441], line_20[439], line_19[437], line_18[435], line_17[433], line_16[431], line_15[429], line_14[427], line_13[425], line_12[423], line_11[421], line_10[419], line_9[417], line_8[415], line_7[413], line_6[411], line_5[409], line_4[407], line_3[405], line_2[403], line_1[401] };
assign col_656 = {line_128[656], line_127[654], line_126[652], line_125[650], line_124[648], line_123[646], line_122[644], line_121[642], line_120[640], line_119[638], line_118[636], line_117[634], line_116[632], line_115[630], line_114[628], line_113[626], line_112[624], line_111[622], line_110[620], line_109[618], line_108[616], line_107[614], line_106[612], line_105[610], line_104[608], line_103[606], line_102[604], line_101[602], line_100[600], line_99[598], line_98[596], line_97[594], line_96[592], line_95[590], line_94[588], line_93[586], line_92[584], line_91[582], line_90[580], line_89[578], line_88[576], line_87[574], line_86[572], line_85[570], line_84[568], line_83[566], line_82[564], line_81[562], line_80[560], line_79[558], line_78[556], line_77[554], line_76[552], line_75[550], line_74[548], line_73[546], line_72[544], line_71[542], line_70[540], line_69[538], line_68[536], line_67[534], line_66[532], line_65[530], line_64[528], line_63[526], line_62[524], line_61[522], line_60[520], line_59[518], line_58[516], line_57[514], line_56[512], line_55[510], line_54[508], line_53[506], line_52[504], line_51[502], line_50[500], line_49[498], line_48[496], line_47[494], line_46[492], line_45[490], line_44[488], line_43[486], line_42[484], line_41[482], line_40[480], line_39[478], line_38[476], line_37[474], line_36[472], line_35[470], line_34[468], line_33[466], line_32[464], line_31[462], line_30[460], line_29[458], line_28[456], line_27[454], line_26[452], line_25[450], line_24[448], line_23[446], line_22[444], line_21[442], line_20[440], line_19[438], line_18[436], line_17[434], line_16[432], line_15[430], line_14[428], line_13[426], line_12[424], line_11[422], line_10[420], line_9[418], line_8[416], line_7[414], line_6[412], line_5[410], line_4[408], line_3[406], line_2[404], line_1[402] };
assign col_657 = {line_128[657], line_127[655], line_126[653], line_125[651], line_124[649], line_123[647], line_122[645], line_121[643], line_120[641], line_119[639], line_118[637], line_117[635], line_116[633], line_115[631], line_114[629], line_113[627], line_112[625], line_111[623], line_110[621], line_109[619], line_108[617], line_107[615], line_106[613], line_105[611], line_104[609], line_103[607], line_102[605], line_101[603], line_100[601], line_99[599], line_98[597], line_97[595], line_96[593], line_95[591], line_94[589], line_93[587], line_92[585], line_91[583], line_90[581], line_89[579], line_88[577], line_87[575], line_86[573], line_85[571], line_84[569], line_83[567], line_82[565], line_81[563], line_80[561], line_79[559], line_78[557], line_77[555], line_76[553], line_75[551], line_74[549], line_73[547], line_72[545], line_71[543], line_70[541], line_69[539], line_68[537], line_67[535], line_66[533], line_65[531], line_64[529], line_63[527], line_62[525], line_61[523], line_60[521], line_59[519], line_58[517], line_57[515], line_56[513], line_55[511], line_54[509], line_53[507], line_52[505], line_51[503], line_50[501], line_49[499], line_48[497], line_47[495], line_46[493], line_45[491], line_44[489], line_43[487], line_42[485], line_41[483], line_40[481], line_39[479], line_38[477], line_37[475], line_36[473], line_35[471], line_34[469], line_33[467], line_32[465], line_31[463], line_30[461], line_29[459], line_28[457], line_27[455], line_26[453], line_25[451], line_24[449], line_23[447], line_22[445], line_21[443], line_20[441], line_19[439], line_18[437], line_17[435], line_16[433], line_15[431], line_14[429], line_13[427], line_12[425], line_11[423], line_10[421], line_9[419], line_8[417], line_7[415], line_6[413], line_5[411], line_4[409], line_3[407], line_2[405], line_1[403] };
assign col_658 = {line_128[658], line_127[656], line_126[654], line_125[652], line_124[650], line_123[648], line_122[646], line_121[644], line_120[642], line_119[640], line_118[638], line_117[636], line_116[634], line_115[632], line_114[630], line_113[628], line_112[626], line_111[624], line_110[622], line_109[620], line_108[618], line_107[616], line_106[614], line_105[612], line_104[610], line_103[608], line_102[606], line_101[604], line_100[602], line_99[600], line_98[598], line_97[596], line_96[594], line_95[592], line_94[590], line_93[588], line_92[586], line_91[584], line_90[582], line_89[580], line_88[578], line_87[576], line_86[574], line_85[572], line_84[570], line_83[568], line_82[566], line_81[564], line_80[562], line_79[560], line_78[558], line_77[556], line_76[554], line_75[552], line_74[550], line_73[548], line_72[546], line_71[544], line_70[542], line_69[540], line_68[538], line_67[536], line_66[534], line_65[532], line_64[530], line_63[528], line_62[526], line_61[524], line_60[522], line_59[520], line_58[518], line_57[516], line_56[514], line_55[512], line_54[510], line_53[508], line_52[506], line_51[504], line_50[502], line_49[500], line_48[498], line_47[496], line_46[494], line_45[492], line_44[490], line_43[488], line_42[486], line_41[484], line_40[482], line_39[480], line_38[478], line_37[476], line_36[474], line_35[472], line_34[470], line_33[468], line_32[466], line_31[464], line_30[462], line_29[460], line_28[458], line_27[456], line_26[454], line_25[452], line_24[450], line_23[448], line_22[446], line_21[444], line_20[442], line_19[440], line_18[438], line_17[436], line_16[434], line_15[432], line_14[430], line_13[428], line_12[426], line_11[424], line_10[422], line_9[420], line_8[418], line_7[416], line_6[414], line_5[412], line_4[410], line_3[408], line_2[406], line_1[404] };
assign col_659 = {line_128[659], line_127[657], line_126[655], line_125[653], line_124[651], line_123[649], line_122[647], line_121[645], line_120[643], line_119[641], line_118[639], line_117[637], line_116[635], line_115[633], line_114[631], line_113[629], line_112[627], line_111[625], line_110[623], line_109[621], line_108[619], line_107[617], line_106[615], line_105[613], line_104[611], line_103[609], line_102[607], line_101[605], line_100[603], line_99[601], line_98[599], line_97[597], line_96[595], line_95[593], line_94[591], line_93[589], line_92[587], line_91[585], line_90[583], line_89[581], line_88[579], line_87[577], line_86[575], line_85[573], line_84[571], line_83[569], line_82[567], line_81[565], line_80[563], line_79[561], line_78[559], line_77[557], line_76[555], line_75[553], line_74[551], line_73[549], line_72[547], line_71[545], line_70[543], line_69[541], line_68[539], line_67[537], line_66[535], line_65[533], line_64[531], line_63[529], line_62[527], line_61[525], line_60[523], line_59[521], line_58[519], line_57[517], line_56[515], line_55[513], line_54[511], line_53[509], line_52[507], line_51[505], line_50[503], line_49[501], line_48[499], line_47[497], line_46[495], line_45[493], line_44[491], line_43[489], line_42[487], line_41[485], line_40[483], line_39[481], line_38[479], line_37[477], line_36[475], line_35[473], line_34[471], line_33[469], line_32[467], line_31[465], line_30[463], line_29[461], line_28[459], line_27[457], line_26[455], line_25[453], line_24[451], line_23[449], line_22[447], line_21[445], line_20[443], line_19[441], line_18[439], line_17[437], line_16[435], line_15[433], line_14[431], line_13[429], line_12[427], line_11[425], line_10[423], line_9[421], line_8[419], line_7[417], line_6[415], line_5[413], line_4[411], line_3[409], line_2[407], line_1[405] };
assign col_660 = {line_128[660], line_127[658], line_126[656], line_125[654], line_124[652], line_123[650], line_122[648], line_121[646], line_120[644], line_119[642], line_118[640], line_117[638], line_116[636], line_115[634], line_114[632], line_113[630], line_112[628], line_111[626], line_110[624], line_109[622], line_108[620], line_107[618], line_106[616], line_105[614], line_104[612], line_103[610], line_102[608], line_101[606], line_100[604], line_99[602], line_98[600], line_97[598], line_96[596], line_95[594], line_94[592], line_93[590], line_92[588], line_91[586], line_90[584], line_89[582], line_88[580], line_87[578], line_86[576], line_85[574], line_84[572], line_83[570], line_82[568], line_81[566], line_80[564], line_79[562], line_78[560], line_77[558], line_76[556], line_75[554], line_74[552], line_73[550], line_72[548], line_71[546], line_70[544], line_69[542], line_68[540], line_67[538], line_66[536], line_65[534], line_64[532], line_63[530], line_62[528], line_61[526], line_60[524], line_59[522], line_58[520], line_57[518], line_56[516], line_55[514], line_54[512], line_53[510], line_52[508], line_51[506], line_50[504], line_49[502], line_48[500], line_47[498], line_46[496], line_45[494], line_44[492], line_43[490], line_42[488], line_41[486], line_40[484], line_39[482], line_38[480], line_37[478], line_36[476], line_35[474], line_34[472], line_33[470], line_32[468], line_31[466], line_30[464], line_29[462], line_28[460], line_27[458], line_26[456], line_25[454], line_24[452], line_23[450], line_22[448], line_21[446], line_20[444], line_19[442], line_18[440], line_17[438], line_16[436], line_15[434], line_14[432], line_13[430], line_12[428], line_11[426], line_10[424], line_9[422], line_8[420], line_7[418], line_6[416], line_5[414], line_4[412], line_3[410], line_2[408], line_1[406] };
assign col_661 = {line_128[661], line_127[659], line_126[657], line_125[655], line_124[653], line_123[651], line_122[649], line_121[647], line_120[645], line_119[643], line_118[641], line_117[639], line_116[637], line_115[635], line_114[633], line_113[631], line_112[629], line_111[627], line_110[625], line_109[623], line_108[621], line_107[619], line_106[617], line_105[615], line_104[613], line_103[611], line_102[609], line_101[607], line_100[605], line_99[603], line_98[601], line_97[599], line_96[597], line_95[595], line_94[593], line_93[591], line_92[589], line_91[587], line_90[585], line_89[583], line_88[581], line_87[579], line_86[577], line_85[575], line_84[573], line_83[571], line_82[569], line_81[567], line_80[565], line_79[563], line_78[561], line_77[559], line_76[557], line_75[555], line_74[553], line_73[551], line_72[549], line_71[547], line_70[545], line_69[543], line_68[541], line_67[539], line_66[537], line_65[535], line_64[533], line_63[531], line_62[529], line_61[527], line_60[525], line_59[523], line_58[521], line_57[519], line_56[517], line_55[515], line_54[513], line_53[511], line_52[509], line_51[507], line_50[505], line_49[503], line_48[501], line_47[499], line_46[497], line_45[495], line_44[493], line_43[491], line_42[489], line_41[487], line_40[485], line_39[483], line_38[481], line_37[479], line_36[477], line_35[475], line_34[473], line_33[471], line_32[469], line_31[467], line_30[465], line_29[463], line_28[461], line_27[459], line_26[457], line_25[455], line_24[453], line_23[451], line_22[449], line_21[447], line_20[445], line_19[443], line_18[441], line_17[439], line_16[437], line_15[435], line_14[433], line_13[431], line_12[429], line_11[427], line_10[425], line_9[423], line_8[421], line_7[419], line_6[417], line_5[415], line_4[413], line_3[411], line_2[409], line_1[407] };
assign col_662 = {line_128[662], line_127[660], line_126[658], line_125[656], line_124[654], line_123[652], line_122[650], line_121[648], line_120[646], line_119[644], line_118[642], line_117[640], line_116[638], line_115[636], line_114[634], line_113[632], line_112[630], line_111[628], line_110[626], line_109[624], line_108[622], line_107[620], line_106[618], line_105[616], line_104[614], line_103[612], line_102[610], line_101[608], line_100[606], line_99[604], line_98[602], line_97[600], line_96[598], line_95[596], line_94[594], line_93[592], line_92[590], line_91[588], line_90[586], line_89[584], line_88[582], line_87[580], line_86[578], line_85[576], line_84[574], line_83[572], line_82[570], line_81[568], line_80[566], line_79[564], line_78[562], line_77[560], line_76[558], line_75[556], line_74[554], line_73[552], line_72[550], line_71[548], line_70[546], line_69[544], line_68[542], line_67[540], line_66[538], line_65[536], line_64[534], line_63[532], line_62[530], line_61[528], line_60[526], line_59[524], line_58[522], line_57[520], line_56[518], line_55[516], line_54[514], line_53[512], line_52[510], line_51[508], line_50[506], line_49[504], line_48[502], line_47[500], line_46[498], line_45[496], line_44[494], line_43[492], line_42[490], line_41[488], line_40[486], line_39[484], line_38[482], line_37[480], line_36[478], line_35[476], line_34[474], line_33[472], line_32[470], line_31[468], line_30[466], line_29[464], line_28[462], line_27[460], line_26[458], line_25[456], line_24[454], line_23[452], line_22[450], line_21[448], line_20[446], line_19[444], line_18[442], line_17[440], line_16[438], line_15[436], line_14[434], line_13[432], line_12[430], line_11[428], line_10[426], line_9[424], line_8[422], line_7[420], line_6[418], line_5[416], line_4[414], line_3[412], line_2[410], line_1[408] };
assign col_663 = {line_128[663], line_127[661], line_126[659], line_125[657], line_124[655], line_123[653], line_122[651], line_121[649], line_120[647], line_119[645], line_118[643], line_117[641], line_116[639], line_115[637], line_114[635], line_113[633], line_112[631], line_111[629], line_110[627], line_109[625], line_108[623], line_107[621], line_106[619], line_105[617], line_104[615], line_103[613], line_102[611], line_101[609], line_100[607], line_99[605], line_98[603], line_97[601], line_96[599], line_95[597], line_94[595], line_93[593], line_92[591], line_91[589], line_90[587], line_89[585], line_88[583], line_87[581], line_86[579], line_85[577], line_84[575], line_83[573], line_82[571], line_81[569], line_80[567], line_79[565], line_78[563], line_77[561], line_76[559], line_75[557], line_74[555], line_73[553], line_72[551], line_71[549], line_70[547], line_69[545], line_68[543], line_67[541], line_66[539], line_65[537], line_64[535], line_63[533], line_62[531], line_61[529], line_60[527], line_59[525], line_58[523], line_57[521], line_56[519], line_55[517], line_54[515], line_53[513], line_52[511], line_51[509], line_50[507], line_49[505], line_48[503], line_47[501], line_46[499], line_45[497], line_44[495], line_43[493], line_42[491], line_41[489], line_40[487], line_39[485], line_38[483], line_37[481], line_36[479], line_35[477], line_34[475], line_33[473], line_32[471], line_31[469], line_30[467], line_29[465], line_28[463], line_27[461], line_26[459], line_25[457], line_24[455], line_23[453], line_22[451], line_21[449], line_20[447], line_19[445], line_18[443], line_17[441], line_16[439], line_15[437], line_14[435], line_13[433], line_12[431], line_11[429], line_10[427], line_9[425], line_8[423], line_7[421], line_6[419], line_5[417], line_4[415], line_3[413], line_2[411], line_1[409] };
assign col_664 = {line_128[664], line_127[662], line_126[660], line_125[658], line_124[656], line_123[654], line_122[652], line_121[650], line_120[648], line_119[646], line_118[644], line_117[642], line_116[640], line_115[638], line_114[636], line_113[634], line_112[632], line_111[630], line_110[628], line_109[626], line_108[624], line_107[622], line_106[620], line_105[618], line_104[616], line_103[614], line_102[612], line_101[610], line_100[608], line_99[606], line_98[604], line_97[602], line_96[600], line_95[598], line_94[596], line_93[594], line_92[592], line_91[590], line_90[588], line_89[586], line_88[584], line_87[582], line_86[580], line_85[578], line_84[576], line_83[574], line_82[572], line_81[570], line_80[568], line_79[566], line_78[564], line_77[562], line_76[560], line_75[558], line_74[556], line_73[554], line_72[552], line_71[550], line_70[548], line_69[546], line_68[544], line_67[542], line_66[540], line_65[538], line_64[536], line_63[534], line_62[532], line_61[530], line_60[528], line_59[526], line_58[524], line_57[522], line_56[520], line_55[518], line_54[516], line_53[514], line_52[512], line_51[510], line_50[508], line_49[506], line_48[504], line_47[502], line_46[500], line_45[498], line_44[496], line_43[494], line_42[492], line_41[490], line_40[488], line_39[486], line_38[484], line_37[482], line_36[480], line_35[478], line_34[476], line_33[474], line_32[472], line_31[470], line_30[468], line_29[466], line_28[464], line_27[462], line_26[460], line_25[458], line_24[456], line_23[454], line_22[452], line_21[450], line_20[448], line_19[446], line_18[444], line_17[442], line_16[440], line_15[438], line_14[436], line_13[434], line_12[432], line_11[430], line_10[428], line_9[426], line_8[424], line_7[422], line_6[420], line_5[418], line_4[416], line_3[414], line_2[412], line_1[410] };
assign col_665 = {line_128[665], line_127[663], line_126[661], line_125[659], line_124[657], line_123[655], line_122[653], line_121[651], line_120[649], line_119[647], line_118[645], line_117[643], line_116[641], line_115[639], line_114[637], line_113[635], line_112[633], line_111[631], line_110[629], line_109[627], line_108[625], line_107[623], line_106[621], line_105[619], line_104[617], line_103[615], line_102[613], line_101[611], line_100[609], line_99[607], line_98[605], line_97[603], line_96[601], line_95[599], line_94[597], line_93[595], line_92[593], line_91[591], line_90[589], line_89[587], line_88[585], line_87[583], line_86[581], line_85[579], line_84[577], line_83[575], line_82[573], line_81[571], line_80[569], line_79[567], line_78[565], line_77[563], line_76[561], line_75[559], line_74[557], line_73[555], line_72[553], line_71[551], line_70[549], line_69[547], line_68[545], line_67[543], line_66[541], line_65[539], line_64[537], line_63[535], line_62[533], line_61[531], line_60[529], line_59[527], line_58[525], line_57[523], line_56[521], line_55[519], line_54[517], line_53[515], line_52[513], line_51[511], line_50[509], line_49[507], line_48[505], line_47[503], line_46[501], line_45[499], line_44[497], line_43[495], line_42[493], line_41[491], line_40[489], line_39[487], line_38[485], line_37[483], line_36[481], line_35[479], line_34[477], line_33[475], line_32[473], line_31[471], line_30[469], line_29[467], line_28[465], line_27[463], line_26[461], line_25[459], line_24[457], line_23[455], line_22[453], line_21[451], line_20[449], line_19[447], line_18[445], line_17[443], line_16[441], line_15[439], line_14[437], line_13[435], line_12[433], line_11[431], line_10[429], line_9[427], line_8[425], line_7[423], line_6[421], line_5[419], line_4[417], line_3[415], line_2[413], line_1[411] };
assign col_666 = {line_128[666], line_127[664], line_126[662], line_125[660], line_124[658], line_123[656], line_122[654], line_121[652], line_120[650], line_119[648], line_118[646], line_117[644], line_116[642], line_115[640], line_114[638], line_113[636], line_112[634], line_111[632], line_110[630], line_109[628], line_108[626], line_107[624], line_106[622], line_105[620], line_104[618], line_103[616], line_102[614], line_101[612], line_100[610], line_99[608], line_98[606], line_97[604], line_96[602], line_95[600], line_94[598], line_93[596], line_92[594], line_91[592], line_90[590], line_89[588], line_88[586], line_87[584], line_86[582], line_85[580], line_84[578], line_83[576], line_82[574], line_81[572], line_80[570], line_79[568], line_78[566], line_77[564], line_76[562], line_75[560], line_74[558], line_73[556], line_72[554], line_71[552], line_70[550], line_69[548], line_68[546], line_67[544], line_66[542], line_65[540], line_64[538], line_63[536], line_62[534], line_61[532], line_60[530], line_59[528], line_58[526], line_57[524], line_56[522], line_55[520], line_54[518], line_53[516], line_52[514], line_51[512], line_50[510], line_49[508], line_48[506], line_47[504], line_46[502], line_45[500], line_44[498], line_43[496], line_42[494], line_41[492], line_40[490], line_39[488], line_38[486], line_37[484], line_36[482], line_35[480], line_34[478], line_33[476], line_32[474], line_31[472], line_30[470], line_29[468], line_28[466], line_27[464], line_26[462], line_25[460], line_24[458], line_23[456], line_22[454], line_21[452], line_20[450], line_19[448], line_18[446], line_17[444], line_16[442], line_15[440], line_14[438], line_13[436], line_12[434], line_11[432], line_10[430], line_9[428], line_8[426], line_7[424], line_6[422], line_5[420], line_4[418], line_3[416], line_2[414], line_1[412] };
assign col_667 = {line_128[667], line_127[665], line_126[663], line_125[661], line_124[659], line_123[657], line_122[655], line_121[653], line_120[651], line_119[649], line_118[647], line_117[645], line_116[643], line_115[641], line_114[639], line_113[637], line_112[635], line_111[633], line_110[631], line_109[629], line_108[627], line_107[625], line_106[623], line_105[621], line_104[619], line_103[617], line_102[615], line_101[613], line_100[611], line_99[609], line_98[607], line_97[605], line_96[603], line_95[601], line_94[599], line_93[597], line_92[595], line_91[593], line_90[591], line_89[589], line_88[587], line_87[585], line_86[583], line_85[581], line_84[579], line_83[577], line_82[575], line_81[573], line_80[571], line_79[569], line_78[567], line_77[565], line_76[563], line_75[561], line_74[559], line_73[557], line_72[555], line_71[553], line_70[551], line_69[549], line_68[547], line_67[545], line_66[543], line_65[541], line_64[539], line_63[537], line_62[535], line_61[533], line_60[531], line_59[529], line_58[527], line_57[525], line_56[523], line_55[521], line_54[519], line_53[517], line_52[515], line_51[513], line_50[511], line_49[509], line_48[507], line_47[505], line_46[503], line_45[501], line_44[499], line_43[497], line_42[495], line_41[493], line_40[491], line_39[489], line_38[487], line_37[485], line_36[483], line_35[481], line_34[479], line_33[477], line_32[475], line_31[473], line_30[471], line_29[469], line_28[467], line_27[465], line_26[463], line_25[461], line_24[459], line_23[457], line_22[455], line_21[453], line_20[451], line_19[449], line_18[447], line_17[445], line_16[443], line_15[441], line_14[439], line_13[437], line_12[435], line_11[433], line_10[431], line_9[429], line_8[427], line_7[425], line_6[423], line_5[421], line_4[419], line_3[417], line_2[415], line_1[413] };
assign col_668 = {line_128[668], line_127[666], line_126[664], line_125[662], line_124[660], line_123[658], line_122[656], line_121[654], line_120[652], line_119[650], line_118[648], line_117[646], line_116[644], line_115[642], line_114[640], line_113[638], line_112[636], line_111[634], line_110[632], line_109[630], line_108[628], line_107[626], line_106[624], line_105[622], line_104[620], line_103[618], line_102[616], line_101[614], line_100[612], line_99[610], line_98[608], line_97[606], line_96[604], line_95[602], line_94[600], line_93[598], line_92[596], line_91[594], line_90[592], line_89[590], line_88[588], line_87[586], line_86[584], line_85[582], line_84[580], line_83[578], line_82[576], line_81[574], line_80[572], line_79[570], line_78[568], line_77[566], line_76[564], line_75[562], line_74[560], line_73[558], line_72[556], line_71[554], line_70[552], line_69[550], line_68[548], line_67[546], line_66[544], line_65[542], line_64[540], line_63[538], line_62[536], line_61[534], line_60[532], line_59[530], line_58[528], line_57[526], line_56[524], line_55[522], line_54[520], line_53[518], line_52[516], line_51[514], line_50[512], line_49[510], line_48[508], line_47[506], line_46[504], line_45[502], line_44[500], line_43[498], line_42[496], line_41[494], line_40[492], line_39[490], line_38[488], line_37[486], line_36[484], line_35[482], line_34[480], line_33[478], line_32[476], line_31[474], line_30[472], line_29[470], line_28[468], line_27[466], line_26[464], line_25[462], line_24[460], line_23[458], line_22[456], line_21[454], line_20[452], line_19[450], line_18[448], line_17[446], line_16[444], line_15[442], line_14[440], line_13[438], line_12[436], line_11[434], line_10[432], line_9[430], line_8[428], line_7[426], line_6[424], line_5[422], line_4[420], line_3[418], line_2[416], line_1[414] };
assign col_669 = {line_128[669], line_127[667], line_126[665], line_125[663], line_124[661], line_123[659], line_122[657], line_121[655], line_120[653], line_119[651], line_118[649], line_117[647], line_116[645], line_115[643], line_114[641], line_113[639], line_112[637], line_111[635], line_110[633], line_109[631], line_108[629], line_107[627], line_106[625], line_105[623], line_104[621], line_103[619], line_102[617], line_101[615], line_100[613], line_99[611], line_98[609], line_97[607], line_96[605], line_95[603], line_94[601], line_93[599], line_92[597], line_91[595], line_90[593], line_89[591], line_88[589], line_87[587], line_86[585], line_85[583], line_84[581], line_83[579], line_82[577], line_81[575], line_80[573], line_79[571], line_78[569], line_77[567], line_76[565], line_75[563], line_74[561], line_73[559], line_72[557], line_71[555], line_70[553], line_69[551], line_68[549], line_67[547], line_66[545], line_65[543], line_64[541], line_63[539], line_62[537], line_61[535], line_60[533], line_59[531], line_58[529], line_57[527], line_56[525], line_55[523], line_54[521], line_53[519], line_52[517], line_51[515], line_50[513], line_49[511], line_48[509], line_47[507], line_46[505], line_45[503], line_44[501], line_43[499], line_42[497], line_41[495], line_40[493], line_39[491], line_38[489], line_37[487], line_36[485], line_35[483], line_34[481], line_33[479], line_32[477], line_31[475], line_30[473], line_29[471], line_28[469], line_27[467], line_26[465], line_25[463], line_24[461], line_23[459], line_22[457], line_21[455], line_20[453], line_19[451], line_18[449], line_17[447], line_16[445], line_15[443], line_14[441], line_13[439], line_12[437], line_11[435], line_10[433], line_9[431], line_8[429], line_7[427], line_6[425], line_5[423], line_4[421], line_3[419], line_2[417], line_1[415] };
assign col_670 = {line_128[670], line_127[668], line_126[666], line_125[664], line_124[662], line_123[660], line_122[658], line_121[656], line_120[654], line_119[652], line_118[650], line_117[648], line_116[646], line_115[644], line_114[642], line_113[640], line_112[638], line_111[636], line_110[634], line_109[632], line_108[630], line_107[628], line_106[626], line_105[624], line_104[622], line_103[620], line_102[618], line_101[616], line_100[614], line_99[612], line_98[610], line_97[608], line_96[606], line_95[604], line_94[602], line_93[600], line_92[598], line_91[596], line_90[594], line_89[592], line_88[590], line_87[588], line_86[586], line_85[584], line_84[582], line_83[580], line_82[578], line_81[576], line_80[574], line_79[572], line_78[570], line_77[568], line_76[566], line_75[564], line_74[562], line_73[560], line_72[558], line_71[556], line_70[554], line_69[552], line_68[550], line_67[548], line_66[546], line_65[544], line_64[542], line_63[540], line_62[538], line_61[536], line_60[534], line_59[532], line_58[530], line_57[528], line_56[526], line_55[524], line_54[522], line_53[520], line_52[518], line_51[516], line_50[514], line_49[512], line_48[510], line_47[508], line_46[506], line_45[504], line_44[502], line_43[500], line_42[498], line_41[496], line_40[494], line_39[492], line_38[490], line_37[488], line_36[486], line_35[484], line_34[482], line_33[480], line_32[478], line_31[476], line_30[474], line_29[472], line_28[470], line_27[468], line_26[466], line_25[464], line_24[462], line_23[460], line_22[458], line_21[456], line_20[454], line_19[452], line_18[450], line_17[448], line_16[446], line_15[444], line_14[442], line_13[440], line_12[438], line_11[436], line_10[434], line_9[432], line_8[430], line_7[428], line_6[426], line_5[424], line_4[422], line_3[420], line_2[418], line_1[416] };
assign col_671 = {line_128[671], line_127[669], line_126[667], line_125[665], line_124[663], line_123[661], line_122[659], line_121[657], line_120[655], line_119[653], line_118[651], line_117[649], line_116[647], line_115[645], line_114[643], line_113[641], line_112[639], line_111[637], line_110[635], line_109[633], line_108[631], line_107[629], line_106[627], line_105[625], line_104[623], line_103[621], line_102[619], line_101[617], line_100[615], line_99[613], line_98[611], line_97[609], line_96[607], line_95[605], line_94[603], line_93[601], line_92[599], line_91[597], line_90[595], line_89[593], line_88[591], line_87[589], line_86[587], line_85[585], line_84[583], line_83[581], line_82[579], line_81[577], line_80[575], line_79[573], line_78[571], line_77[569], line_76[567], line_75[565], line_74[563], line_73[561], line_72[559], line_71[557], line_70[555], line_69[553], line_68[551], line_67[549], line_66[547], line_65[545], line_64[543], line_63[541], line_62[539], line_61[537], line_60[535], line_59[533], line_58[531], line_57[529], line_56[527], line_55[525], line_54[523], line_53[521], line_52[519], line_51[517], line_50[515], line_49[513], line_48[511], line_47[509], line_46[507], line_45[505], line_44[503], line_43[501], line_42[499], line_41[497], line_40[495], line_39[493], line_38[491], line_37[489], line_36[487], line_35[485], line_34[483], line_33[481], line_32[479], line_31[477], line_30[475], line_29[473], line_28[471], line_27[469], line_26[467], line_25[465], line_24[463], line_23[461], line_22[459], line_21[457], line_20[455], line_19[453], line_18[451], line_17[449], line_16[447], line_15[445], line_14[443], line_13[441], line_12[439], line_11[437], line_10[435], line_9[433], line_8[431], line_7[429], line_6[427], line_5[425], line_4[423], line_3[421], line_2[419], line_1[417] };
assign col_672 = {line_128[672], line_127[670], line_126[668], line_125[666], line_124[664], line_123[662], line_122[660], line_121[658], line_120[656], line_119[654], line_118[652], line_117[650], line_116[648], line_115[646], line_114[644], line_113[642], line_112[640], line_111[638], line_110[636], line_109[634], line_108[632], line_107[630], line_106[628], line_105[626], line_104[624], line_103[622], line_102[620], line_101[618], line_100[616], line_99[614], line_98[612], line_97[610], line_96[608], line_95[606], line_94[604], line_93[602], line_92[600], line_91[598], line_90[596], line_89[594], line_88[592], line_87[590], line_86[588], line_85[586], line_84[584], line_83[582], line_82[580], line_81[578], line_80[576], line_79[574], line_78[572], line_77[570], line_76[568], line_75[566], line_74[564], line_73[562], line_72[560], line_71[558], line_70[556], line_69[554], line_68[552], line_67[550], line_66[548], line_65[546], line_64[544], line_63[542], line_62[540], line_61[538], line_60[536], line_59[534], line_58[532], line_57[530], line_56[528], line_55[526], line_54[524], line_53[522], line_52[520], line_51[518], line_50[516], line_49[514], line_48[512], line_47[510], line_46[508], line_45[506], line_44[504], line_43[502], line_42[500], line_41[498], line_40[496], line_39[494], line_38[492], line_37[490], line_36[488], line_35[486], line_34[484], line_33[482], line_32[480], line_31[478], line_30[476], line_29[474], line_28[472], line_27[470], line_26[468], line_25[466], line_24[464], line_23[462], line_22[460], line_21[458], line_20[456], line_19[454], line_18[452], line_17[450], line_16[448], line_15[446], line_14[444], line_13[442], line_12[440], line_11[438], line_10[436], line_9[434], line_8[432], line_7[430], line_6[428], line_5[426], line_4[424], line_3[422], line_2[420], line_1[418] };
assign col_673 = {line_128[673], line_127[671], line_126[669], line_125[667], line_124[665], line_123[663], line_122[661], line_121[659], line_120[657], line_119[655], line_118[653], line_117[651], line_116[649], line_115[647], line_114[645], line_113[643], line_112[641], line_111[639], line_110[637], line_109[635], line_108[633], line_107[631], line_106[629], line_105[627], line_104[625], line_103[623], line_102[621], line_101[619], line_100[617], line_99[615], line_98[613], line_97[611], line_96[609], line_95[607], line_94[605], line_93[603], line_92[601], line_91[599], line_90[597], line_89[595], line_88[593], line_87[591], line_86[589], line_85[587], line_84[585], line_83[583], line_82[581], line_81[579], line_80[577], line_79[575], line_78[573], line_77[571], line_76[569], line_75[567], line_74[565], line_73[563], line_72[561], line_71[559], line_70[557], line_69[555], line_68[553], line_67[551], line_66[549], line_65[547], line_64[545], line_63[543], line_62[541], line_61[539], line_60[537], line_59[535], line_58[533], line_57[531], line_56[529], line_55[527], line_54[525], line_53[523], line_52[521], line_51[519], line_50[517], line_49[515], line_48[513], line_47[511], line_46[509], line_45[507], line_44[505], line_43[503], line_42[501], line_41[499], line_40[497], line_39[495], line_38[493], line_37[491], line_36[489], line_35[487], line_34[485], line_33[483], line_32[481], line_31[479], line_30[477], line_29[475], line_28[473], line_27[471], line_26[469], line_25[467], line_24[465], line_23[463], line_22[461], line_21[459], line_20[457], line_19[455], line_18[453], line_17[451], line_16[449], line_15[447], line_14[445], line_13[443], line_12[441], line_11[439], line_10[437], line_9[435], line_8[433], line_7[431], line_6[429], line_5[427], line_4[425], line_3[423], line_2[421], line_1[419] };
assign col_674 = {line_128[674], line_127[672], line_126[670], line_125[668], line_124[666], line_123[664], line_122[662], line_121[660], line_120[658], line_119[656], line_118[654], line_117[652], line_116[650], line_115[648], line_114[646], line_113[644], line_112[642], line_111[640], line_110[638], line_109[636], line_108[634], line_107[632], line_106[630], line_105[628], line_104[626], line_103[624], line_102[622], line_101[620], line_100[618], line_99[616], line_98[614], line_97[612], line_96[610], line_95[608], line_94[606], line_93[604], line_92[602], line_91[600], line_90[598], line_89[596], line_88[594], line_87[592], line_86[590], line_85[588], line_84[586], line_83[584], line_82[582], line_81[580], line_80[578], line_79[576], line_78[574], line_77[572], line_76[570], line_75[568], line_74[566], line_73[564], line_72[562], line_71[560], line_70[558], line_69[556], line_68[554], line_67[552], line_66[550], line_65[548], line_64[546], line_63[544], line_62[542], line_61[540], line_60[538], line_59[536], line_58[534], line_57[532], line_56[530], line_55[528], line_54[526], line_53[524], line_52[522], line_51[520], line_50[518], line_49[516], line_48[514], line_47[512], line_46[510], line_45[508], line_44[506], line_43[504], line_42[502], line_41[500], line_40[498], line_39[496], line_38[494], line_37[492], line_36[490], line_35[488], line_34[486], line_33[484], line_32[482], line_31[480], line_30[478], line_29[476], line_28[474], line_27[472], line_26[470], line_25[468], line_24[466], line_23[464], line_22[462], line_21[460], line_20[458], line_19[456], line_18[454], line_17[452], line_16[450], line_15[448], line_14[446], line_13[444], line_12[442], line_11[440], line_10[438], line_9[436], line_8[434], line_7[432], line_6[430], line_5[428], line_4[426], line_3[424], line_2[422], line_1[420] };
assign col_675 = {line_128[675], line_127[673], line_126[671], line_125[669], line_124[667], line_123[665], line_122[663], line_121[661], line_120[659], line_119[657], line_118[655], line_117[653], line_116[651], line_115[649], line_114[647], line_113[645], line_112[643], line_111[641], line_110[639], line_109[637], line_108[635], line_107[633], line_106[631], line_105[629], line_104[627], line_103[625], line_102[623], line_101[621], line_100[619], line_99[617], line_98[615], line_97[613], line_96[611], line_95[609], line_94[607], line_93[605], line_92[603], line_91[601], line_90[599], line_89[597], line_88[595], line_87[593], line_86[591], line_85[589], line_84[587], line_83[585], line_82[583], line_81[581], line_80[579], line_79[577], line_78[575], line_77[573], line_76[571], line_75[569], line_74[567], line_73[565], line_72[563], line_71[561], line_70[559], line_69[557], line_68[555], line_67[553], line_66[551], line_65[549], line_64[547], line_63[545], line_62[543], line_61[541], line_60[539], line_59[537], line_58[535], line_57[533], line_56[531], line_55[529], line_54[527], line_53[525], line_52[523], line_51[521], line_50[519], line_49[517], line_48[515], line_47[513], line_46[511], line_45[509], line_44[507], line_43[505], line_42[503], line_41[501], line_40[499], line_39[497], line_38[495], line_37[493], line_36[491], line_35[489], line_34[487], line_33[485], line_32[483], line_31[481], line_30[479], line_29[477], line_28[475], line_27[473], line_26[471], line_25[469], line_24[467], line_23[465], line_22[463], line_21[461], line_20[459], line_19[457], line_18[455], line_17[453], line_16[451], line_15[449], line_14[447], line_13[445], line_12[443], line_11[441], line_10[439], line_9[437], line_8[435], line_7[433], line_6[431], line_5[429], line_4[427], line_3[425], line_2[423], line_1[421] };
assign col_676 = {line_128[676], line_127[674], line_126[672], line_125[670], line_124[668], line_123[666], line_122[664], line_121[662], line_120[660], line_119[658], line_118[656], line_117[654], line_116[652], line_115[650], line_114[648], line_113[646], line_112[644], line_111[642], line_110[640], line_109[638], line_108[636], line_107[634], line_106[632], line_105[630], line_104[628], line_103[626], line_102[624], line_101[622], line_100[620], line_99[618], line_98[616], line_97[614], line_96[612], line_95[610], line_94[608], line_93[606], line_92[604], line_91[602], line_90[600], line_89[598], line_88[596], line_87[594], line_86[592], line_85[590], line_84[588], line_83[586], line_82[584], line_81[582], line_80[580], line_79[578], line_78[576], line_77[574], line_76[572], line_75[570], line_74[568], line_73[566], line_72[564], line_71[562], line_70[560], line_69[558], line_68[556], line_67[554], line_66[552], line_65[550], line_64[548], line_63[546], line_62[544], line_61[542], line_60[540], line_59[538], line_58[536], line_57[534], line_56[532], line_55[530], line_54[528], line_53[526], line_52[524], line_51[522], line_50[520], line_49[518], line_48[516], line_47[514], line_46[512], line_45[510], line_44[508], line_43[506], line_42[504], line_41[502], line_40[500], line_39[498], line_38[496], line_37[494], line_36[492], line_35[490], line_34[488], line_33[486], line_32[484], line_31[482], line_30[480], line_29[478], line_28[476], line_27[474], line_26[472], line_25[470], line_24[468], line_23[466], line_22[464], line_21[462], line_20[460], line_19[458], line_18[456], line_17[454], line_16[452], line_15[450], line_14[448], line_13[446], line_12[444], line_11[442], line_10[440], line_9[438], line_8[436], line_7[434], line_6[432], line_5[430], line_4[428], line_3[426], line_2[424], line_1[422] };
assign col_677 = {line_128[677], line_127[675], line_126[673], line_125[671], line_124[669], line_123[667], line_122[665], line_121[663], line_120[661], line_119[659], line_118[657], line_117[655], line_116[653], line_115[651], line_114[649], line_113[647], line_112[645], line_111[643], line_110[641], line_109[639], line_108[637], line_107[635], line_106[633], line_105[631], line_104[629], line_103[627], line_102[625], line_101[623], line_100[621], line_99[619], line_98[617], line_97[615], line_96[613], line_95[611], line_94[609], line_93[607], line_92[605], line_91[603], line_90[601], line_89[599], line_88[597], line_87[595], line_86[593], line_85[591], line_84[589], line_83[587], line_82[585], line_81[583], line_80[581], line_79[579], line_78[577], line_77[575], line_76[573], line_75[571], line_74[569], line_73[567], line_72[565], line_71[563], line_70[561], line_69[559], line_68[557], line_67[555], line_66[553], line_65[551], line_64[549], line_63[547], line_62[545], line_61[543], line_60[541], line_59[539], line_58[537], line_57[535], line_56[533], line_55[531], line_54[529], line_53[527], line_52[525], line_51[523], line_50[521], line_49[519], line_48[517], line_47[515], line_46[513], line_45[511], line_44[509], line_43[507], line_42[505], line_41[503], line_40[501], line_39[499], line_38[497], line_37[495], line_36[493], line_35[491], line_34[489], line_33[487], line_32[485], line_31[483], line_30[481], line_29[479], line_28[477], line_27[475], line_26[473], line_25[471], line_24[469], line_23[467], line_22[465], line_21[463], line_20[461], line_19[459], line_18[457], line_17[455], line_16[453], line_15[451], line_14[449], line_13[447], line_12[445], line_11[443], line_10[441], line_9[439], line_8[437], line_7[435], line_6[433], line_5[431], line_4[429], line_3[427], line_2[425], line_1[423] };
assign col_678 = {line_128[678], line_127[676], line_126[674], line_125[672], line_124[670], line_123[668], line_122[666], line_121[664], line_120[662], line_119[660], line_118[658], line_117[656], line_116[654], line_115[652], line_114[650], line_113[648], line_112[646], line_111[644], line_110[642], line_109[640], line_108[638], line_107[636], line_106[634], line_105[632], line_104[630], line_103[628], line_102[626], line_101[624], line_100[622], line_99[620], line_98[618], line_97[616], line_96[614], line_95[612], line_94[610], line_93[608], line_92[606], line_91[604], line_90[602], line_89[600], line_88[598], line_87[596], line_86[594], line_85[592], line_84[590], line_83[588], line_82[586], line_81[584], line_80[582], line_79[580], line_78[578], line_77[576], line_76[574], line_75[572], line_74[570], line_73[568], line_72[566], line_71[564], line_70[562], line_69[560], line_68[558], line_67[556], line_66[554], line_65[552], line_64[550], line_63[548], line_62[546], line_61[544], line_60[542], line_59[540], line_58[538], line_57[536], line_56[534], line_55[532], line_54[530], line_53[528], line_52[526], line_51[524], line_50[522], line_49[520], line_48[518], line_47[516], line_46[514], line_45[512], line_44[510], line_43[508], line_42[506], line_41[504], line_40[502], line_39[500], line_38[498], line_37[496], line_36[494], line_35[492], line_34[490], line_33[488], line_32[486], line_31[484], line_30[482], line_29[480], line_28[478], line_27[476], line_26[474], line_25[472], line_24[470], line_23[468], line_22[466], line_21[464], line_20[462], line_19[460], line_18[458], line_17[456], line_16[454], line_15[452], line_14[450], line_13[448], line_12[446], line_11[444], line_10[442], line_9[440], line_8[438], line_7[436], line_6[434], line_5[432], line_4[430], line_3[428], line_2[426], line_1[424] };
assign col_679 = {line_128[679], line_127[677], line_126[675], line_125[673], line_124[671], line_123[669], line_122[667], line_121[665], line_120[663], line_119[661], line_118[659], line_117[657], line_116[655], line_115[653], line_114[651], line_113[649], line_112[647], line_111[645], line_110[643], line_109[641], line_108[639], line_107[637], line_106[635], line_105[633], line_104[631], line_103[629], line_102[627], line_101[625], line_100[623], line_99[621], line_98[619], line_97[617], line_96[615], line_95[613], line_94[611], line_93[609], line_92[607], line_91[605], line_90[603], line_89[601], line_88[599], line_87[597], line_86[595], line_85[593], line_84[591], line_83[589], line_82[587], line_81[585], line_80[583], line_79[581], line_78[579], line_77[577], line_76[575], line_75[573], line_74[571], line_73[569], line_72[567], line_71[565], line_70[563], line_69[561], line_68[559], line_67[557], line_66[555], line_65[553], line_64[551], line_63[549], line_62[547], line_61[545], line_60[543], line_59[541], line_58[539], line_57[537], line_56[535], line_55[533], line_54[531], line_53[529], line_52[527], line_51[525], line_50[523], line_49[521], line_48[519], line_47[517], line_46[515], line_45[513], line_44[511], line_43[509], line_42[507], line_41[505], line_40[503], line_39[501], line_38[499], line_37[497], line_36[495], line_35[493], line_34[491], line_33[489], line_32[487], line_31[485], line_30[483], line_29[481], line_28[479], line_27[477], line_26[475], line_25[473], line_24[471], line_23[469], line_22[467], line_21[465], line_20[463], line_19[461], line_18[459], line_17[457], line_16[455], line_15[453], line_14[451], line_13[449], line_12[447], line_11[445], line_10[443], line_9[441], line_8[439], line_7[437], line_6[435], line_5[433], line_4[431], line_3[429], line_2[427], line_1[425] };
assign col_680 = {line_128[680], line_127[678], line_126[676], line_125[674], line_124[672], line_123[670], line_122[668], line_121[666], line_120[664], line_119[662], line_118[660], line_117[658], line_116[656], line_115[654], line_114[652], line_113[650], line_112[648], line_111[646], line_110[644], line_109[642], line_108[640], line_107[638], line_106[636], line_105[634], line_104[632], line_103[630], line_102[628], line_101[626], line_100[624], line_99[622], line_98[620], line_97[618], line_96[616], line_95[614], line_94[612], line_93[610], line_92[608], line_91[606], line_90[604], line_89[602], line_88[600], line_87[598], line_86[596], line_85[594], line_84[592], line_83[590], line_82[588], line_81[586], line_80[584], line_79[582], line_78[580], line_77[578], line_76[576], line_75[574], line_74[572], line_73[570], line_72[568], line_71[566], line_70[564], line_69[562], line_68[560], line_67[558], line_66[556], line_65[554], line_64[552], line_63[550], line_62[548], line_61[546], line_60[544], line_59[542], line_58[540], line_57[538], line_56[536], line_55[534], line_54[532], line_53[530], line_52[528], line_51[526], line_50[524], line_49[522], line_48[520], line_47[518], line_46[516], line_45[514], line_44[512], line_43[510], line_42[508], line_41[506], line_40[504], line_39[502], line_38[500], line_37[498], line_36[496], line_35[494], line_34[492], line_33[490], line_32[488], line_31[486], line_30[484], line_29[482], line_28[480], line_27[478], line_26[476], line_25[474], line_24[472], line_23[470], line_22[468], line_21[466], line_20[464], line_19[462], line_18[460], line_17[458], line_16[456], line_15[454], line_14[452], line_13[450], line_12[448], line_11[446], line_10[444], line_9[442], line_8[440], line_7[438], line_6[436], line_5[434], line_4[432], line_3[430], line_2[428], line_1[426] };
assign col_681 = {line_128[681], line_127[679], line_126[677], line_125[675], line_124[673], line_123[671], line_122[669], line_121[667], line_120[665], line_119[663], line_118[661], line_117[659], line_116[657], line_115[655], line_114[653], line_113[651], line_112[649], line_111[647], line_110[645], line_109[643], line_108[641], line_107[639], line_106[637], line_105[635], line_104[633], line_103[631], line_102[629], line_101[627], line_100[625], line_99[623], line_98[621], line_97[619], line_96[617], line_95[615], line_94[613], line_93[611], line_92[609], line_91[607], line_90[605], line_89[603], line_88[601], line_87[599], line_86[597], line_85[595], line_84[593], line_83[591], line_82[589], line_81[587], line_80[585], line_79[583], line_78[581], line_77[579], line_76[577], line_75[575], line_74[573], line_73[571], line_72[569], line_71[567], line_70[565], line_69[563], line_68[561], line_67[559], line_66[557], line_65[555], line_64[553], line_63[551], line_62[549], line_61[547], line_60[545], line_59[543], line_58[541], line_57[539], line_56[537], line_55[535], line_54[533], line_53[531], line_52[529], line_51[527], line_50[525], line_49[523], line_48[521], line_47[519], line_46[517], line_45[515], line_44[513], line_43[511], line_42[509], line_41[507], line_40[505], line_39[503], line_38[501], line_37[499], line_36[497], line_35[495], line_34[493], line_33[491], line_32[489], line_31[487], line_30[485], line_29[483], line_28[481], line_27[479], line_26[477], line_25[475], line_24[473], line_23[471], line_22[469], line_21[467], line_20[465], line_19[463], line_18[461], line_17[459], line_16[457], line_15[455], line_14[453], line_13[451], line_12[449], line_11[447], line_10[445], line_9[443], line_8[441], line_7[439], line_6[437], line_5[435], line_4[433], line_3[431], line_2[429], line_1[427] };
assign col_682 = {line_128[682], line_127[680], line_126[678], line_125[676], line_124[674], line_123[672], line_122[670], line_121[668], line_120[666], line_119[664], line_118[662], line_117[660], line_116[658], line_115[656], line_114[654], line_113[652], line_112[650], line_111[648], line_110[646], line_109[644], line_108[642], line_107[640], line_106[638], line_105[636], line_104[634], line_103[632], line_102[630], line_101[628], line_100[626], line_99[624], line_98[622], line_97[620], line_96[618], line_95[616], line_94[614], line_93[612], line_92[610], line_91[608], line_90[606], line_89[604], line_88[602], line_87[600], line_86[598], line_85[596], line_84[594], line_83[592], line_82[590], line_81[588], line_80[586], line_79[584], line_78[582], line_77[580], line_76[578], line_75[576], line_74[574], line_73[572], line_72[570], line_71[568], line_70[566], line_69[564], line_68[562], line_67[560], line_66[558], line_65[556], line_64[554], line_63[552], line_62[550], line_61[548], line_60[546], line_59[544], line_58[542], line_57[540], line_56[538], line_55[536], line_54[534], line_53[532], line_52[530], line_51[528], line_50[526], line_49[524], line_48[522], line_47[520], line_46[518], line_45[516], line_44[514], line_43[512], line_42[510], line_41[508], line_40[506], line_39[504], line_38[502], line_37[500], line_36[498], line_35[496], line_34[494], line_33[492], line_32[490], line_31[488], line_30[486], line_29[484], line_28[482], line_27[480], line_26[478], line_25[476], line_24[474], line_23[472], line_22[470], line_21[468], line_20[466], line_19[464], line_18[462], line_17[460], line_16[458], line_15[456], line_14[454], line_13[452], line_12[450], line_11[448], line_10[446], line_9[444], line_8[442], line_7[440], line_6[438], line_5[436], line_4[434], line_3[432], line_2[430], line_1[428] };
assign col_683 = {line_128[683], line_127[681], line_126[679], line_125[677], line_124[675], line_123[673], line_122[671], line_121[669], line_120[667], line_119[665], line_118[663], line_117[661], line_116[659], line_115[657], line_114[655], line_113[653], line_112[651], line_111[649], line_110[647], line_109[645], line_108[643], line_107[641], line_106[639], line_105[637], line_104[635], line_103[633], line_102[631], line_101[629], line_100[627], line_99[625], line_98[623], line_97[621], line_96[619], line_95[617], line_94[615], line_93[613], line_92[611], line_91[609], line_90[607], line_89[605], line_88[603], line_87[601], line_86[599], line_85[597], line_84[595], line_83[593], line_82[591], line_81[589], line_80[587], line_79[585], line_78[583], line_77[581], line_76[579], line_75[577], line_74[575], line_73[573], line_72[571], line_71[569], line_70[567], line_69[565], line_68[563], line_67[561], line_66[559], line_65[557], line_64[555], line_63[553], line_62[551], line_61[549], line_60[547], line_59[545], line_58[543], line_57[541], line_56[539], line_55[537], line_54[535], line_53[533], line_52[531], line_51[529], line_50[527], line_49[525], line_48[523], line_47[521], line_46[519], line_45[517], line_44[515], line_43[513], line_42[511], line_41[509], line_40[507], line_39[505], line_38[503], line_37[501], line_36[499], line_35[497], line_34[495], line_33[493], line_32[491], line_31[489], line_30[487], line_29[485], line_28[483], line_27[481], line_26[479], line_25[477], line_24[475], line_23[473], line_22[471], line_21[469], line_20[467], line_19[465], line_18[463], line_17[461], line_16[459], line_15[457], line_14[455], line_13[453], line_12[451], line_11[449], line_10[447], line_9[445], line_8[443], line_7[441], line_6[439], line_5[437], line_4[435], line_3[433], line_2[431], line_1[429] };
assign col_684 = {line_128[684], line_127[682], line_126[680], line_125[678], line_124[676], line_123[674], line_122[672], line_121[670], line_120[668], line_119[666], line_118[664], line_117[662], line_116[660], line_115[658], line_114[656], line_113[654], line_112[652], line_111[650], line_110[648], line_109[646], line_108[644], line_107[642], line_106[640], line_105[638], line_104[636], line_103[634], line_102[632], line_101[630], line_100[628], line_99[626], line_98[624], line_97[622], line_96[620], line_95[618], line_94[616], line_93[614], line_92[612], line_91[610], line_90[608], line_89[606], line_88[604], line_87[602], line_86[600], line_85[598], line_84[596], line_83[594], line_82[592], line_81[590], line_80[588], line_79[586], line_78[584], line_77[582], line_76[580], line_75[578], line_74[576], line_73[574], line_72[572], line_71[570], line_70[568], line_69[566], line_68[564], line_67[562], line_66[560], line_65[558], line_64[556], line_63[554], line_62[552], line_61[550], line_60[548], line_59[546], line_58[544], line_57[542], line_56[540], line_55[538], line_54[536], line_53[534], line_52[532], line_51[530], line_50[528], line_49[526], line_48[524], line_47[522], line_46[520], line_45[518], line_44[516], line_43[514], line_42[512], line_41[510], line_40[508], line_39[506], line_38[504], line_37[502], line_36[500], line_35[498], line_34[496], line_33[494], line_32[492], line_31[490], line_30[488], line_29[486], line_28[484], line_27[482], line_26[480], line_25[478], line_24[476], line_23[474], line_22[472], line_21[470], line_20[468], line_19[466], line_18[464], line_17[462], line_16[460], line_15[458], line_14[456], line_13[454], line_12[452], line_11[450], line_10[448], line_9[446], line_8[444], line_7[442], line_6[440], line_5[438], line_4[436], line_3[434], line_2[432], line_1[430] };
assign col_685 = {line_128[685], line_127[683], line_126[681], line_125[679], line_124[677], line_123[675], line_122[673], line_121[671], line_120[669], line_119[667], line_118[665], line_117[663], line_116[661], line_115[659], line_114[657], line_113[655], line_112[653], line_111[651], line_110[649], line_109[647], line_108[645], line_107[643], line_106[641], line_105[639], line_104[637], line_103[635], line_102[633], line_101[631], line_100[629], line_99[627], line_98[625], line_97[623], line_96[621], line_95[619], line_94[617], line_93[615], line_92[613], line_91[611], line_90[609], line_89[607], line_88[605], line_87[603], line_86[601], line_85[599], line_84[597], line_83[595], line_82[593], line_81[591], line_80[589], line_79[587], line_78[585], line_77[583], line_76[581], line_75[579], line_74[577], line_73[575], line_72[573], line_71[571], line_70[569], line_69[567], line_68[565], line_67[563], line_66[561], line_65[559], line_64[557], line_63[555], line_62[553], line_61[551], line_60[549], line_59[547], line_58[545], line_57[543], line_56[541], line_55[539], line_54[537], line_53[535], line_52[533], line_51[531], line_50[529], line_49[527], line_48[525], line_47[523], line_46[521], line_45[519], line_44[517], line_43[515], line_42[513], line_41[511], line_40[509], line_39[507], line_38[505], line_37[503], line_36[501], line_35[499], line_34[497], line_33[495], line_32[493], line_31[491], line_30[489], line_29[487], line_28[485], line_27[483], line_26[481], line_25[479], line_24[477], line_23[475], line_22[473], line_21[471], line_20[469], line_19[467], line_18[465], line_17[463], line_16[461], line_15[459], line_14[457], line_13[455], line_12[453], line_11[451], line_10[449], line_9[447], line_8[445], line_7[443], line_6[441], line_5[439], line_4[437], line_3[435], line_2[433], line_1[431] };
assign col_686 = {line_128[686], line_127[684], line_126[682], line_125[680], line_124[678], line_123[676], line_122[674], line_121[672], line_120[670], line_119[668], line_118[666], line_117[664], line_116[662], line_115[660], line_114[658], line_113[656], line_112[654], line_111[652], line_110[650], line_109[648], line_108[646], line_107[644], line_106[642], line_105[640], line_104[638], line_103[636], line_102[634], line_101[632], line_100[630], line_99[628], line_98[626], line_97[624], line_96[622], line_95[620], line_94[618], line_93[616], line_92[614], line_91[612], line_90[610], line_89[608], line_88[606], line_87[604], line_86[602], line_85[600], line_84[598], line_83[596], line_82[594], line_81[592], line_80[590], line_79[588], line_78[586], line_77[584], line_76[582], line_75[580], line_74[578], line_73[576], line_72[574], line_71[572], line_70[570], line_69[568], line_68[566], line_67[564], line_66[562], line_65[560], line_64[558], line_63[556], line_62[554], line_61[552], line_60[550], line_59[548], line_58[546], line_57[544], line_56[542], line_55[540], line_54[538], line_53[536], line_52[534], line_51[532], line_50[530], line_49[528], line_48[526], line_47[524], line_46[522], line_45[520], line_44[518], line_43[516], line_42[514], line_41[512], line_40[510], line_39[508], line_38[506], line_37[504], line_36[502], line_35[500], line_34[498], line_33[496], line_32[494], line_31[492], line_30[490], line_29[488], line_28[486], line_27[484], line_26[482], line_25[480], line_24[478], line_23[476], line_22[474], line_21[472], line_20[470], line_19[468], line_18[466], line_17[464], line_16[462], line_15[460], line_14[458], line_13[456], line_12[454], line_11[452], line_10[450], line_9[448], line_8[446], line_7[444], line_6[442], line_5[440], line_4[438], line_3[436], line_2[434], line_1[432] };
assign col_687 = {line_128[687], line_127[685], line_126[683], line_125[681], line_124[679], line_123[677], line_122[675], line_121[673], line_120[671], line_119[669], line_118[667], line_117[665], line_116[663], line_115[661], line_114[659], line_113[657], line_112[655], line_111[653], line_110[651], line_109[649], line_108[647], line_107[645], line_106[643], line_105[641], line_104[639], line_103[637], line_102[635], line_101[633], line_100[631], line_99[629], line_98[627], line_97[625], line_96[623], line_95[621], line_94[619], line_93[617], line_92[615], line_91[613], line_90[611], line_89[609], line_88[607], line_87[605], line_86[603], line_85[601], line_84[599], line_83[597], line_82[595], line_81[593], line_80[591], line_79[589], line_78[587], line_77[585], line_76[583], line_75[581], line_74[579], line_73[577], line_72[575], line_71[573], line_70[571], line_69[569], line_68[567], line_67[565], line_66[563], line_65[561], line_64[559], line_63[557], line_62[555], line_61[553], line_60[551], line_59[549], line_58[547], line_57[545], line_56[543], line_55[541], line_54[539], line_53[537], line_52[535], line_51[533], line_50[531], line_49[529], line_48[527], line_47[525], line_46[523], line_45[521], line_44[519], line_43[517], line_42[515], line_41[513], line_40[511], line_39[509], line_38[507], line_37[505], line_36[503], line_35[501], line_34[499], line_33[497], line_32[495], line_31[493], line_30[491], line_29[489], line_28[487], line_27[485], line_26[483], line_25[481], line_24[479], line_23[477], line_22[475], line_21[473], line_20[471], line_19[469], line_18[467], line_17[465], line_16[463], line_15[461], line_14[459], line_13[457], line_12[455], line_11[453], line_10[451], line_9[449], line_8[447], line_7[445], line_6[443], line_5[441], line_4[439], line_3[437], line_2[435], line_1[433] };
assign col_688 = {line_128[688], line_127[686], line_126[684], line_125[682], line_124[680], line_123[678], line_122[676], line_121[674], line_120[672], line_119[670], line_118[668], line_117[666], line_116[664], line_115[662], line_114[660], line_113[658], line_112[656], line_111[654], line_110[652], line_109[650], line_108[648], line_107[646], line_106[644], line_105[642], line_104[640], line_103[638], line_102[636], line_101[634], line_100[632], line_99[630], line_98[628], line_97[626], line_96[624], line_95[622], line_94[620], line_93[618], line_92[616], line_91[614], line_90[612], line_89[610], line_88[608], line_87[606], line_86[604], line_85[602], line_84[600], line_83[598], line_82[596], line_81[594], line_80[592], line_79[590], line_78[588], line_77[586], line_76[584], line_75[582], line_74[580], line_73[578], line_72[576], line_71[574], line_70[572], line_69[570], line_68[568], line_67[566], line_66[564], line_65[562], line_64[560], line_63[558], line_62[556], line_61[554], line_60[552], line_59[550], line_58[548], line_57[546], line_56[544], line_55[542], line_54[540], line_53[538], line_52[536], line_51[534], line_50[532], line_49[530], line_48[528], line_47[526], line_46[524], line_45[522], line_44[520], line_43[518], line_42[516], line_41[514], line_40[512], line_39[510], line_38[508], line_37[506], line_36[504], line_35[502], line_34[500], line_33[498], line_32[496], line_31[494], line_30[492], line_29[490], line_28[488], line_27[486], line_26[484], line_25[482], line_24[480], line_23[478], line_22[476], line_21[474], line_20[472], line_19[470], line_18[468], line_17[466], line_16[464], line_15[462], line_14[460], line_13[458], line_12[456], line_11[454], line_10[452], line_9[450], line_8[448], line_7[446], line_6[444], line_5[442], line_4[440], line_3[438], line_2[436], line_1[434] };
assign col_689 = {line_128[689], line_127[687], line_126[685], line_125[683], line_124[681], line_123[679], line_122[677], line_121[675], line_120[673], line_119[671], line_118[669], line_117[667], line_116[665], line_115[663], line_114[661], line_113[659], line_112[657], line_111[655], line_110[653], line_109[651], line_108[649], line_107[647], line_106[645], line_105[643], line_104[641], line_103[639], line_102[637], line_101[635], line_100[633], line_99[631], line_98[629], line_97[627], line_96[625], line_95[623], line_94[621], line_93[619], line_92[617], line_91[615], line_90[613], line_89[611], line_88[609], line_87[607], line_86[605], line_85[603], line_84[601], line_83[599], line_82[597], line_81[595], line_80[593], line_79[591], line_78[589], line_77[587], line_76[585], line_75[583], line_74[581], line_73[579], line_72[577], line_71[575], line_70[573], line_69[571], line_68[569], line_67[567], line_66[565], line_65[563], line_64[561], line_63[559], line_62[557], line_61[555], line_60[553], line_59[551], line_58[549], line_57[547], line_56[545], line_55[543], line_54[541], line_53[539], line_52[537], line_51[535], line_50[533], line_49[531], line_48[529], line_47[527], line_46[525], line_45[523], line_44[521], line_43[519], line_42[517], line_41[515], line_40[513], line_39[511], line_38[509], line_37[507], line_36[505], line_35[503], line_34[501], line_33[499], line_32[497], line_31[495], line_30[493], line_29[491], line_28[489], line_27[487], line_26[485], line_25[483], line_24[481], line_23[479], line_22[477], line_21[475], line_20[473], line_19[471], line_18[469], line_17[467], line_16[465], line_15[463], line_14[461], line_13[459], line_12[457], line_11[455], line_10[453], line_9[451], line_8[449], line_7[447], line_6[445], line_5[443], line_4[441], line_3[439], line_2[437], line_1[435] };
assign col_690 = {line_128[690], line_127[688], line_126[686], line_125[684], line_124[682], line_123[680], line_122[678], line_121[676], line_120[674], line_119[672], line_118[670], line_117[668], line_116[666], line_115[664], line_114[662], line_113[660], line_112[658], line_111[656], line_110[654], line_109[652], line_108[650], line_107[648], line_106[646], line_105[644], line_104[642], line_103[640], line_102[638], line_101[636], line_100[634], line_99[632], line_98[630], line_97[628], line_96[626], line_95[624], line_94[622], line_93[620], line_92[618], line_91[616], line_90[614], line_89[612], line_88[610], line_87[608], line_86[606], line_85[604], line_84[602], line_83[600], line_82[598], line_81[596], line_80[594], line_79[592], line_78[590], line_77[588], line_76[586], line_75[584], line_74[582], line_73[580], line_72[578], line_71[576], line_70[574], line_69[572], line_68[570], line_67[568], line_66[566], line_65[564], line_64[562], line_63[560], line_62[558], line_61[556], line_60[554], line_59[552], line_58[550], line_57[548], line_56[546], line_55[544], line_54[542], line_53[540], line_52[538], line_51[536], line_50[534], line_49[532], line_48[530], line_47[528], line_46[526], line_45[524], line_44[522], line_43[520], line_42[518], line_41[516], line_40[514], line_39[512], line_38[510], line_37[508], line_36[506], line_35[504], line_34[502], line_33[500], line_32[498], line_31[496], line_30[494], line_29[492], line_28[490], line_27[488], line_26[486], line_25[484], line_24[482], line_23[480], line_22[478], line_21[476], line_20[474], line_19[472], line_18[470], line_17[468], line_16[466], line_15[464], line_14[462], line_13[460], line_12[458], line_11[456], line_10[454], line_9[452], line_8[450], line_7[448], line_6[446], line_5[444], line_4[442], line_3[440], line_2[438], line_1[436] };
assign col_691 = {line_128[691], line_127[689], line_126[687], line_125[685], line_124[683], line_123[681], line_122[679], line_121[677], line_120[675], line_119[673], line_118[671], line_117[669], line_116[667], line_115[665], line_114[663], line_113[661], line_112[659], line_111[657], line_110[655], line_109[653], line_108[651], line_107[649], line_106[647], line_105[645], line_104[643], line_103[641], line_102[639], line_101[637], line_100[635], line_99[633], line_98[631], line_97[629], line_96[627], line_95[625], line_94[623], line_93[621], line_92[619], line_91[617], line_90[615], line_89[613], line_88[611], line_87[609], line_86[607], line_85[605], line_84[603], line_83[601], line_82[599], line_81[597], line_80[595], line_79[593], line_78[591], line_77[589], line_76[587], line_75[585], line_74[583], line_73[581], line_72[579], line_71[577], line_70[575], line_69[573], line_68[571], line_67[569], line_66[567], line_65[565], line_64[563], line_63[561], line_62[559], line_61[557], line_60[555], line_59[553], line_58[551], line_57[549], line_56[547], line_55[545], line_54[543], line_53[541], line_52[539], line_51[537], line_50[535], line_49[533], line_48[531], line_47[529], line_46[527], line_45[525], line_44[523], line_43[521], line_42[519], line_41[517], line_40[515], line_39[513], line_38[511], line_37[509], line_36[507], line_35[505], line_34[503], line_33[501], line_32[499], line_31[497], line_30[495], line_29[493], line_28[491], line_27[489], line_26[487], line_25[485], line_24[483], line_23[481], line_22[479], line_21[477], line_20[475], line_19[473], line_18[471], line_17[469], line_16[467], line_15[465], line_14[463], line_13[461], line_12[459], line_11[457], line_10[455], line_9[453], line_8[451], line_7[449], line_6[447], line_5[445], line_4[443], line_3[441], line_2[439], line_1[437] };
assign col_692 = {line_128[692], line_127[690], line_126[688], line_125[686], line_124[684], line_123[682], line_122[680], line_121[678], line_120[676], line_119[674], line_118[672], line_117[670], line_116[668], line_115[666], line_114[664], line_113[662], line_112[660], line_111[658], line_110[656], line_109[654], line_108[652], line_107[650], line_106[648], line_105[646], line_104[644], line_103[642], line_102[640], line_101[638], line_100[636], line_99[634], line_98[632], line_97[630], line_96[628], line_95[626], line_94[624], line_93[622], line_92[620], line_91[618], line_90[616], line_89[614], line_88[612], line_87[610], line_86[608], line_85[606], line_84[604], line_83[602], line_82[600], line_81[598], line_80[596], line_79[594], line_78[592], line_77[590], line_76[588], line_75[586], line_74[584], line_73[582], line_72[580], line_71[578], line_70[576], line_69[574], line_68[572], line_67[570], line_66[568], line_65[566], line_64[564], line_63[562], line_62[560], line_61[558], line_60[556], line_59[554], line_58[552], line_57[550], line_56[548], line_55[546], line_54[544], line_53[542], line_52[540], line_51[538], line_50[536], line_49[534], line_48[532], line_47[530], line_46[528], line_45[526], line_44[524], line_43[522], line_42[520], line_41[518], line_40[516], line_39[514], line_38[512], line_37[510], line_36[508], line_35[506], line_34[504], line_33[502], line_32[500], line_31[498], line_30[496], line_29[494], line_28[492], line_27[490], line_26[488], line_25[486], line_24[484], line_23[482], line_22[480], line_21[478], line_20[476], line_19[474], line_18[472], line_17[470], line_16[468], line_15[466], line_14[464], line_13[462], line_12[460], line_11[458], line_10[456], line_9[454], line_8[452], line_7[450], line_6[448], line_5[446], line_4[444], line_3[442], line_2[440], line_1[438] };
assign col_693 = {line_128[693], line_127[691], line_126[689], line_125[687], line_124[685], line_123[683], line_122[681], line_121[679], line_120[677], line_119[675], line_118[673], line_117[671], line_116[669], line_115[667], line_114[665], line_113[663], line_112[661], line_111[659], line_110[657], line_109[655], line_108[653], line_107[651], line_106[649], line_105[647], line_104[645], line_103[643], line_102[641], line_101[639], line_100[637], line_99[635], line_98[633], line_97[631], line_96[629], line_95[627], line_94[625], line_93[623], line_92[621], line_91[619], line_90[617], line_89[615], line_88[613], line_87[611], line_86[609], line_85[607], line_84[605], line_83[603], line_82[601], line_81[599], line_80[597], line_79[595], line_78[593], line_77[591], line_76[589], line_75[587], line_74[585], line_73[583], line_72[581], line_71[579], line_70[577], line_69[575], line_68[573], line_67[571], line_66[569], line_65[567], line_64[565], line_63[563], line_62[561], line_61[559], line_60[557], line_59[555], line_58[553], line_57[551], line_56[549], line_55[547], line_54[545], line_53[543], line_52[541], line_51[539], line_50[537], line_49[535], line_48[533], line_47[531], line_46[529], line_45[527], line_44[525], line_43[523], line_42[521], line_41[519], line_40[517], line_39[515], line_38[513], line_37[511], line_36[509], line_35[507], line_34[505], line_33[503], line_32[501], line_31[499], line_30[497], line_29[495], line_28[493], line_27[491], line_26[489], line_25[487], line_24[485], line_23[483], line_22[481], line_21[479], line_20[477], line_19[475], line_18[473], line_17[471], line_16[469], line_15[467], line_14[465], line_13[463], line_12[461], line_11[459], line_10[457], line_9[455], line_8[453], line_7[451], line_6[449], line_5[447], line_4[445], line_3[443], line_2[441], line_1[439] };
assign col_694 = {line_128[694], line_127[692], line_126[690], line_125[688], line_124[686], line_123[684], line_122[682], line_121[680], line_120[678], line_119[676], line_118[674], line_117[672], line_116[670], line_115[668], line_114[666], line_113[664], line_112[662], line_111[660], line_110[658], line_109[656], line_108[654], line_107[652], line_106[650], line_105[648], line_104[646], line_103[644], line_102[642], line_101[640], line_100[638], line_99[636], line_98[634], line_97[632], line_96[630], line_95[628], line_94[626], line_93[624], line_92[622], line_91[620], line_90[618], line_89[616], line_88[614], line_87[612], line_86[610], line_85[608], line_84[606], line_83[604], line_82[602], line_81[600], line_80[598], line_79[596], line_78[594], line_77[592], line_76[590], line_75[588], line_74[586], line_73[584], line_72[582], line_71[580], line_70[578], line_69[576], line_68[574], line_67[572], line_66[570], line_65[568], line_64[566], line_63[564], line_62[562], line_61[560], line_60[558], line_59[556], line_58[554], line_57[552], line_56[550], line_55[548], line_54[546], line_53[544], line_52[542], line_51[540], line_50[538], line_49[536], line_48[534], line_47[532], line_46[530], line_45[528], line_44[526], line_43[524], line_42[522], line_41[520], line_40[518], line_39[516], line_38[514], line_37[512], line_36[510], line_35[508], line_34[506], line_33[504], line_32[502], line_31[500], line_30[498], line_29[496], line_28[494], line_27[492], line_26[490], line_25[488], line_24[486], line_23[484], line_22[482], line_21[480], line_20[478], line_19[476], line_18[474], line_17[472], line_16[470], line_15[468], line_14[466], line_13[464], line_12[462], line_11[460], line_10[458], line_9[456], line_8[454], line_7[452], line_6[450], line_5[448], line_4[446], line_3[444], line_2[442], line_1[440] };
assign col_695 = {line_128[695], line_127[693], line_126[691], line_125[689], line_124[687], line_123[685], line_122[683], line_121[681], line_120[679], line_119[677], line_118[675], line_117[673], line_116[671], line_115[669], line_114[667], line_113[665], line_112[663], line_111[661], line_110[659], line_109[657], line_108[655], line_107[653], line_106[651], line_105[649], line_104[647], line_103[645], line_102[643], line_101[641], line_100[639], line_99[637], line_98[635], line_97[633], line_96[631], line_95[629], line_94[627], line_93[625], line_92[623], line_91[621], line_90[619], line_89[617], line_88[615], line_87[613], line_86[611], line_85[609], line_84[607], line_83[605], line_82[603], line_81[601], line_80[599], line_79[597], line_78[595], line_77[593], line_76[591], line_75[589], line_74[587], line_73[585], line_72[583], line_71[581], line_70[579], line_69[577], line_68[575], line_67[573], line_66[571], line_65[569], line_64[567], line_63[565], line_62[563], line_61[561], line_60[559], line_59[557], line_58[555], line_57[553], line_56[551], line_55[549], line_54[547], line_53[545], line_52[543], line_51[541], line_50[539], line_49[537], line_48[535], line_47[533], line_46[531], line_45[529], line_44[527], line_43[525], line_42[523], line_41[521], line_40[519], line_39[517], line_38[515], line_37[513], line_36[511], line_35[509], line_34[507], line_33[505], line_32[503], line_31[501], line_30[499], line_29[497], line_28[495], line_27[493], line_26[491], line_25[489], line_24[487], line_23[485], line_22[483], line_21[481], line_20[479], line_19[477], line_18[475], line_17[473], line_16[471], line_15[469], line_14[467], line_13[465], line_12[463], line_11[461], line_10[459], line_9[457], line_8[455], line_7[453], line_6[451], line_5[449], line_4[447], line_3[445], line_2[443], line_1[441] };
assign col_696 = {line_128[696], line_127[694], line_126[692], line_125[690], line_124[688], line_123[686], line_122[684], line_121[682], line_120[680], line_119[678], line_118[676], line_117[674], line_116[672], line_115[670], line_114[668], line_113[666], line_112[664], line_111[662], line_110[660], line_109[658], line_108[656], line_107[654], line_106[652], line_105[650], line_104[648], line_103[646], line_102[644], line_101[642], line_100[640], line_99[638], line_98[636], line_97[634], line_96[632], line_95[630], line_94[628], line_93[626], line_92[624], line_91[622], line_90[620], line_89[618], line_88[616], line_87[614], line_86[612], line_85[610], line_84[608], line_83[606], line_82[604], line_81[602], line_80[600], line_79[598], line_78[596], line_77[594], line_76[592], line_75[590], line_74[588], line_73[586], line_72[584], line_71[582], line_70[580], line_69[578], line_68[576], line_67[574], line_66[572], line_65[570], line_64[568], line_63[566], line_62[564], line_61[562], line_60[560], line_59[558], line_58[556], line_57[554], line_56[552], line_55[550], line_54[548], line_53[546], line_52[544], line_51[542], line_50[540], line_49[538], line_48[536], line_47[534], line_46[532], line_45[530], line_44[528], line_43[526], line_42[524], line_41[522], line_40[520], line_39[518], line_38[516], line_37[514], line_36[512], line_35[510], line_34[508], line_33[506], line_32[504], line_31[502], line_30[500], line_29[498], line_28[496], line_27[494], line_26[492], line_25[490], line_24[488], line_23[486], line_22[484], line_21[482], line_20[480], line_19[478], line_18[476], line_17[474], line_16[472], line_15[470], line_14[468], line_13[466], line_12[464], line_11[462], line_10[460], line_9[458], line_8[456], line_7[454], line_6[452], line_5[450], line_4[448], line_3[446], line_2[444], line_1[442] };
assign col_697 = {line_128[697], line_127[695], line_126[693], line_125[691], line_124[689], line_123[687], line_122[685], line_121[683], line_120[681], line_119[679], line_118[677], line_117[675], line_116[673], line_115[671], line_114[669], line_113[667], line_112[665], line_111[663], line_110[661], line_109[659], line_108[657], line_107[655], line_106[653], line_105[651], line_104[649], line_103[647], line_102[645], line_101[643], line_100[641], line_99[639], line_98[637], line_97[635], line_96[633], line_95[631], line_94[629], line_93[627], line_92[625], line_91[623], line_90[621], line_89[619], line_88[617], line_87[615], line_86[613], line_85[611], line_84[609], line_83[607], line_82[605], line_81[603], line_80[601], line_79[599], line_78[597], line_77[595], line_76[593], line_75[591], line_74[589], line_73[587], line_72[585], line_71[583], line_70[581], line_69[579], line_68[577], line_67[575], line_66[573], line_65[571], line_64[569], line_63[567], line_62[565], line_61[563], line_60[561], line_59[559], line_58[557], line_57[555], line_56[553], line_55[551], line_54[549], line_53[547], line_52[545], line_51[543], line_50[541], line_49[539], line_48[537], line_47[535], line_46[533], line_45[531], line_44[529], line_43[527], line_42[525], line_41[523], line_40[521], line_39[519], line_38[517], line_37[515], line_36[513], line_35[511], line_34[509], line_33[507], line_32[505], line_31[503], line_30[501], line_29[499], line_28[497], line_27[495], line_26[493], line_25[491], line_24[489], line_23[487], line_22[485], line_21[483], line_20[481], line_19[479], line_18[477], line_17[475], line_16[473], line_15[471], line_14[469], line_13[467], line_12[465], line_11[463], line_10[461], line_9[459], line_8[457], line_7[455], line_6[453], line_5[451], line_4[449], line_3[447], line_2[445], line_1[443] };
assign col_698 = {line_128[698], line_127[696], line_126[694], line_125[692], line_124[690], line_123[688], line_122[686], line_121[684], line_120[682], line_119[680], line_118[678], line_117[676], line_116[674], line_115[672], line_114[670], line_113[668], line_112[666], line_111[664], line_110[662], line_109[660], line_108[658], line_107[656], line_106[654], line_105[652], line_104[650], line_103[648], line_102[646], line_101[644], line_100[642], line_99[640], line_98[638], line_97[636], line_96[634], line_95[632], line_94[630], line_93[628], line_92[626], line_91[624], line_90[622], line_89[620], line_88[618], line_87[616], line_86[614], line_85[612], line_84[610], line_83[608], line_82[606], line_81[604], line_80[602], line_79[600], line_78[598], line_77[596], line_76[594], line_75[592], line_74[590], line_73[588], line_72[586], line_71[584], line_70[582], line_69[580], line_68[578], line_67[576], line_66[574], line_65[572], line_64[570], line_63[568], line_62[566], line_61[564], line_60[562], line_59[560], line_58[558], line_57[556], line_56[554], line_55[552], line_54[550], line_53[548], line_52[546], line_51[544], line_50[542], line_49[540], line_48[538], line_47[536], line_46[534], line_45[532], line_44[530], line_43[528], line_42[526], line_41[524], line_40[522], line_39[520], line_38[518], line_37[516], line_36[514], line_35[512], line_34[510], line_33[508], line_32[506], line_31[504], line_30[502], line_29[500], line_28[498], line_27[496], line_26[494], line_25[492], line_24[490], line_23[488], line_22[486], line_21[484], line_20[482], line_19[480], line_18[478], line_17[476], line_16[474], line_15[472], line_14[470], line_13[468], line_12[466], line_11[464], line_10[462], line_9[460], line_8[458], line_7[456], line_6[454], line_5[452], line_4[450], line_3[448], line_2[446], line_1[444] };
assign col_699 = {line_128[699], line_127[697], line_126[695], line_125[693], line_124[691], line_123[689], line_122[687], line_121[685], line_120[683], line_119[681], line_118[679], line_117[677], line_116[675], line_115[673], line_114[671], line_113[669], line_112[667], line_111[665], line_110[663], line_109[661], line_108[659], line_107[657], line_106[655], line_105[653], line_104[651], line_103[649], line_102[647], line_101[645], line_100[643], line_99[641], line_98[639], line_97[637], line_96[635], line_95[633], line_94[631], line_93[629], line_92[627], line_91[625], line_90[623], line_89[621], line_88[619], line_87[617], line_86[615], line_85[613], line_84[611], line_83[609], line_82[607], line_81[605], line_80[603], line_79[601], line_78[599], line_77[597], line_76[595], line_75[593], line_74[591], line_73[589], line_72[587], line_71[585], line_70[583], line_69[581], line_68[579], line_67[577], line_66[575], line_65[573], line_64[571], line_63[569], line_62[567], line_61[565], line_60[563], line_59[561], line_58[559], line_57[557], line_56[555], line_55[553], line_54[551], line_53[549], line_52[547], line_51[545], line_50[543], line_49[541], line_48[539], line_47[537], line_46[535], line_45[533], line_44[531], line_43[529], line_42[527], line_41[525], line_40[523], line_39[521], line_38[519], line_37[517], line_36[515], line_35[513], line_34[511], line_33[509], line_32[507], line_31[505], line_30[503], line_29[501], line_28[499], line_27[497], line_26[495], line_25[493], line_24[491], line_23[489], line_22[487], line_21[485], line_20[483], line_19[481], line_18[479], line_17[477], line_16[475], line_15[473], line_14[471], line_13[469], line_12[467], line_11[465], line_10[463], line_9[461], line_8[459], line_7[457], line_6[455], line_5[453], line_4[451], line_3[449], line_2[447], line_1[445] };
assign col_700 = {line_128[700], line_127[698], line_126[696], line_125[694], line_124[692], line_123[690], line_122[688], line_121[686], line_120[684], line_119[682], line_118[680], line_117[678], line_116[676], line_115[674], line_114[672], line_113[670], line_112[668], line_111[666], line_110[664], line_109[662], line_108[660], line_107[658], line_106[656], line_105[654], line_104[652], line_103[650], line_102[648], line_101[646], line_100[644], line_99[642], line_98[640], line_97[638], line_96[636], line_95[634], line_94[632], line_93[630], line_92[628], line_91[626], line_90[624], line_89[622], line_88[620], line_87[618], line_86[616], line_85[614], line_84[612], line_83[610], line_82[608], line_81[606], line_80[604], line_79[602], line_78[600], line_77[598], line_76[596], line_75[594], line_74[592], line_73[590], line_72[588], line_71[586], line_70[584], line_69[582], line_68[580], line_67[578], line_66[576], line_65[574], line_64[572], line_63[570], line_62[568], line_61[566], line_60[564], line_59[562], line_58[560], line_57[558], line_56[556], line_55[554], line_54[552], line_53[550], line_52[548], line_51[546], line_50[544], line_49[542], line_48[540], line_47[538], line_46[536], line_45[534], line_44[532], line_43[530], line_42[528], line_41[526], line_40[524], line_39[522], line_38[520], line_37[518], line_36[516], line_35[514], line_34[512], line_33[510], line_32[508], line_31[506], line_30[504], line_29[502], line_28[500], line_27[498], line_26[496], line_25[494], line_24[492], line_23[490], line_22[488], line_21[486], line_20[484], line_19[482], line_18[480], line_17[478], line_16[476], line_15[474], line_14[472], line_13[470], line_12[468], line_11[466], line_10[464], line_9[462], line_8[460], line_7[458], line_6[456], line_5[454], line_4[452], line_3[450], line_2[448], line_1[446] };
assign col_701 = {line_128[701], line_127[699], line_126[697], line_125[695], line_124[693], line_123[691], line_122[689], line_121[687], line_120[685], line_119[683], line_118[681], line_117[679], line_116[677], line_115[675], line_114[673], line_113[671], line_112[669], line_111[667], line_110[665], line_109[663], line_108[661], line_107[659], line_106[657], line_105[655], line_104[653], line_103[651], line_102[649], line_101[647], line_100[645], line_99[643], line_98[641], line_97[639], line_96[637], line_95[635], line_94[633], line_93[631], line_92[629], line_91[627], line_90[625], line_89[623], line_88[621], line_87[619], line_86[617], line_85[615], line_84[613], line_83[611], line_82[609], line_81[607], line_80[605], line_79[603], line_78[601], line_77[599], line_76[597], line_75[595], line_74[593], line_73[591], line_72[589], line_71[587], line_70[585], line_69[583], line_68[581], line_67[579], line_66[577], line_65[575], line_64[573], line_63[571], line_62[569], line_61[567], line_60[565], line_59[563], line_58[561], line_57[559], line_56[557], line_55[555], line_54[553], line_53[551], line_52[549], line_51[547], line_50[545], line_49[543], line_48[541], line_47[539], line_46[537], line_45[535], line_44[533], line_43[531], line_42[529], line_41[527], line_40[525], line_39[523], line_38[521], line_37[519], line_36[517], line_35[515], line_34[513], line_33[511], line_32[509], line_31[507], line_30[505], line_29[503], line_28[501], line_27[499], line_26[497], line_25[495], line_24[493], line_23[491], line_22[489], line_21[487], line_20[485], line_19[483], line_18[481], line_17[479], line_16[477], line_15[475], line_14[473], line_13[471], line_12[469], line_11[467], line_10[465], line_9[463], line_8[461], line_7[459], line_6[457], line_5[455], line_4[453], line_3[451], line_2[449], line_1[447] };
assign col_702 = {line_128[702], line_127[700], line_126[698], line_125[696], line_124[694], line_123[692], line_122[690], line_121[688], line_120[686], line_119[684], line_118[682], line_117[680], line_116[678], line_115[676], line_114[674], line_113[672], line_112[670], line_111[668], line_110[666], line_109[664], line_108[662], line_107[660], line_106[658], line_105[656], line_104[654], line_103[652], line_102[650], line_101[648], line_100[646], line_99[644], line_98[642], line_97[640], line_96[638], line_95[636], line_94[634], line_93[632], line_92[630], line_91[628], line_90[626], line_89[624], line_88[622], line_87[620], line_86[618], line_85[616], line_84[614], line_83[612], line_82[610], line_81[608], line_80[606], line_79[604], line_78[602], line_77[600], line_76[598], line_75[596], line_74[594], line_73[592], line_72[590], line_71[588], line_70[586], line_69[584], line_68[582], line_67[580], line_66[578], line_65[576], line_64[574], line_63[572], line_62[570], line_61[568], line_60[566], line_59[564], line_58[562], line_57[560], line_56[558], line_55[556], line_54[554], line_53[552], line_52[550], line_51[548], line_50[546], line_49[544], line_48[542], line_47[540], line_46[538], line_45[536], line_44[534], line_43[532], line_42[530], line_41[528], line_40[526], line_39[524], line_38[522], line_37[520], line_36[518], line_35[516], line_34[514], line_33[512], line_32[510], line_31[508], line_30[506], line_29[504], line_28[502], line_27[500], line_26[498], line_25[496], line_24[494], line_23[492], line_22[490], line_21[488], line_20[486], line_19[484], line_18[482], line_17[480], line_16[478], line_15[476], line_14[474], line_13[472], line_12[470], line_11[468], line_10[466], line_9[464], line_8[462], line_7[460], line_6[458], line_5[456], line_4[454], line_3[452], line_2[450], line_1[448] };
assign col_703 = {line_128[703], line_127[701], line_126[699], line_125[697], line_124[695], line_123[693], line_122[691], line_121[689], line_120[687], line_119[685], line_118[683], line_117[681], line_116[679], line_115[677], line_114[675], line_113[673], line_112[671], line_111[669], line_110[667], line_109[665], line_108[663], line_107[661], line_106[659], line_105[657], line_104[655], line_103[653], line_102[651], line_101[649], line_100[647], line_99[645], line_98[643], line_97[641], line_96[639], line_95[637], line_94[635], line_93[633], line_92[631], line_91[629], line_90[627], line_89[625], line_88[623], line_87[621], line_86[619], line_85[617], line_84[615], line_83[613], line_82[611], line_81[609], line_80[607], line_79[605], line_78[603], line_77[601], line_76[599], line_75[597], line_74[595], line_73[593], line_72[591], line_71[589], line_70[587], line_69[585], line_68[583], line_67[581], line_66[579], line_65[577], line_64[575], line_63[573], line_62[571], line_61[569], line_60[567], line_59[565], line_58[563], line_57[561], line_56[559], line_55[557], line_54[555], line_53[553], line_52[551], line_51[549], line_50[547], line_49[545], line_48[543], line_47[541], line_46[539], line_45[537], line_44[535], line_43[533], line_42[531], line_41[529], line_40[527], line_39[525], line_38[523], line_37[521], line_36[519], line_35[517], line_34[515], line_33[513], line_32[511], line_31[509], line_30[507], line_29[505], line_28[503], line_27[501], line_26[499], line_25[497], line_24[495], line_23[493], line_22[491], line_21[489], line_20[487], line_19[485], line_18[483], line_17[481], line_16[479], line_15[477], line_14[475], line_13[473], line_12[471], line_11[469], line_10[467], line_9[465], line_8[463], line_7[461], line_6[459], line_5[457], line_4[455], line_3[453], line_2[451], line_1[449] };
assign col_704 = {line_128[704], line_127[702], line_126[700], line_125[698], line_124[696], line_123[694], line_122[692], line_121[690], line_120[688], line_119[686], line_118[684], line_117[682], line_116[680], line_115[678], line_114[676], line_113[674], line_112[672], line_111[670], line_110[668], line_109[666], line_108[664], line_107[662], line_106[660], line_105[658], line_104[656], line_103[654], line_102[652], line_101[650], line_100[648], line_99[646], line_98[644], line_97[642], line_96[640], line_95[638], line_94[636], line_93[634], line_92[632], line_91[630], line_90[628], line_89[626], line_88[624], line_87[622], line_86[620], line_85[618], line_84[616], line_83[614], line_82[612], line_81[610], line_80[608], line_79[606], line_78[604], line_77[602], line_76[600], line_75[598], line_74[596], line_73[594], line_72[592], line_71[590], line_70[588], line_69[586], line_68[584], line_67[582], line_66[580], line_65[578], line_64[576], line_63[574], line_62[572], line_61[570], line_60[568], line_59[566], line_58[564], line_57[562], line_56[560], line_55[558], line_54[556], line_53[554], line_52[552], line_51[550], line_50[548], line_49[546], line_48[544], line_47[542], line_46[540], line_45[538], line_44[536], line_43[534], line_42[532], line_41[530], line_40[528], line_39[526], line_38[524], line_37[522], line_36[520], line_35[518], line_34[516], line_33[514], line_32[512], line_31[510], line_30[508], line_29[506], line_28[504], line_27[502], line_26[500], line_25[498], line_24[496], line_23[494], line_22[492], line_21[490], line_20[488], line_19[486], line_18[484], line_17[482], line_16[480], line_15[478], line_14[476], line_13[474], line_12[472], line_11[470], line_10[468], line_9[466], line_8[464], line_7[462], line_6[460], line_5[458], line_4[456], line_3[454], line_2[452], line_1[450] };
assign col_705 = {line_128[705], line_127[703], line_126[701], line_125[699], line_124[697], line_123[695], line_122[693], line_121[691], line_120[689], line_119[687], line_118[685], line_117[683], line_116[681], line_115[679], line_114[677], line_113[675], line_112[673], line_111[671], line_110[669], line_109[667], line_108[665], line_107[663], line_106[661], line_105[659], line_104[657], line_103[655], line_102[653], line_101[651], line_100[649], line_99[647], line_98[645], line_97[643], line_96[641], line_95[639], line_94[637], line_93[635], line_92[633], line_91[631], line_90[629], line_89[627], line_88[625], line_87[623], line_86[621], line_85[619], line_84[617], line_83[615], line_82[613], line_81[611], line_80[609], line_79[607], line_78[605], line_77[603], line_76[601], line_75[599], line_74[597], line_73[595], line_72[593], line_71[591], line_70[589], line_69[587], line_68[585], line_67[583], line_66[581], line_65[579], line_64[577], line_63[575], line_62[573], line_61[571], line_60[569], line_59[567], line_58[565], line_57[563], line_56[561], line_55[559], line_54[557], line_53[555], line_52[553], line_51[551], line_50[549], line_49[547], line_48[545], line_47[543], line_46[541], line_45[539], line_44[537], line_43[535], line_42[533], line_41[531], line_40[529], line_39[527], line_38[525], line_37[523], line_36[521], line_35[519], line_34[517], line_33[515], line_32[513], line_31[511], line_30[509], line_29[507], line_28[505], line_27[503], line_26[501], line_25[499], line_24[497], line_23[495], line_22[493], line_21[491], line_20[489], line_19[487], line_18[485], line_17[483], line_16[481], line_15[479], line_14[477], line_13[475], line_12[473], line_11[471], line_10[469], line_9[467], line_8[465], line_7[463], line_6[461], line_5[459], line_4[457], line_3[455], line_2[453], line_1[451] };
assign col_706 = {line_128[706], line_127[704], line_126[702], line_125[700], line_124[698], line_123[696], line_122[694], line_121[692], line_120[690], line_119[688], line_118[686], line_117[684], line_116[682], line_115[680], line_114[678], line_113[676], line_112[674], line_111[672], line_110[670], line_109[668], line_108[666], line_107[664], line_106[662], line_105[660], line_104[658], line_103[656], line_102[654], line_101[652], line_100[650], line_99[648], line_98[646], line_97[644], line_96[642], line_95[640], line_94[638], line_93[636], line_92[634], line_91[632], line_90[630], line_89[628], line_88[626], line_87[624], line_86[622], line_85[620], line_84[618], line_83[616], line_82[614], line_81[612], line_80[610], line_79[608], line_78[606], line_77[604], line_76[602], line_75[600], line_74[598], line_73[596], line_72[594], line_71[592], line_70[590], line_69[588], line_68[586], line_67[584], line_66[582], line_65[580], line_64[578], line_63[576], line_62[574], line_61[572], line_60[570], line_59[568], line_58[566], line_57[564], line_56[562], line_55[560], line_54[558], line_53[556], line_52[554], line_51[552], line_50[550], line_49[548], line_48[546], line_47[544], line_46[542], line_45[540], line_44[538], line_43[536], line_42[534], line_41[532], line_40[530], line_39[528], line_38[526], line_37[524], line_36[522], line_35[520], line_34[518], line_33[516], line_32[514], line_31[512], line_30[510], line_29[508], line_28[506], line_27[504], line_26[502], line_25[500], line_24[498], line_23[496], line_22[494], line_21[492], line_20[490], line_19[488], line_18[486], line_17[484], line_16[482], line_15[480], line_14[478], line_13[476], line_12[474], line_11[472], line_10[470], line_9[468], line_8[466], line_7[464], line_6[462], line_5[460], line_4[458], line_3[456], line_2[454], line_1[452] };
assign col_707 = {line_128[707], line_127[705], line_126[703], line_125[701], line_124[699], line_123[697], line_122[695], line_121[693], line_120[691], line_119[689], line_118[687], line_117[685], line_116[683], line_115[681], line_114[679], line_113[677], line_112[675], line_111[673], line_110[671], line_109[669], line_108[667], line_107[665], line_106[663], line_105[661], line_104[659], line_103[657], line_102[655], line_101[653], line_100[651], line_99[649], line_98[647], line_97[645], line_96[643], line_95[641], line_94[639], line_93[637], line_92[635], line_91[633], line_90[631], line_89[629], line_88[627], line_87[625], line_86[623], line_85[621], line_84[619], line_83[617], line_82[615], line_81[613], line_80[611], line_79[609], line_78[607], line_77[605], line_76[603], line_75[601], line_74[599], line_73[597], line_72[595], line_71[593], line_70[591], line_69[589], line_68[587], line_67[585], line_66[583], line_65[581], line_64[579], line_63[577], line_62[575], line_61[573], line_60[571], line_59[569], line_58[567], line_57[565], line_56[563], line_55[561], line_54[559], line_53[557], line_52[555], line_51[553], line_50[551], line_49[549], line_48[547], line_47[545], line_46[543], line_45[541], line_44[539], line_43[537], line_42[535], line_41[533], line_40[531], line_39[529], line_38[527], line_37[525], line_36[523], line_35[521], line_34[519], line_33[517], line_32[515], line_31[513], line_30[511], line_29[509], line_28[507], line_27[505], line_26[503], line_25[501], line_24[499], line_23[497], line_22[495], line_21[493], line_20[491], line_19[489], line_18[487], line_17[485], line_16[483], line_15[481], line_14[479], line_13[477], line_12[475], line_11[473], line_10[471], line_9[469], line_8[467], line_7[465], line_6[463], line_5[461], line_4[459], line_3[457], line_2[455], line_1[453] };
assign col_708 = {line_128[708], line_127[706], line_126[704], line_125[702], line_124[700], line_123[698], line_122[696], line_121[694], line_120[692], line_119[690], line_118[688], line_117[686], line_116[684], line_115[682], line_114[680], line_113[678], line_112[676], line_111[674], line_110[672], line_109[670], line_108[668], line_107[666], line_106[664], line_105[662], line_104[660], line_103[658], line_102[656], line_101[654], line_100[652], line_99[650], line_98[648], line_97[646], line_96[644], line_95[642], line_94[640], line_93[638], line_92[636], line_91[634], line_90[632], line_89[630], line_88[628], line_87[626], line_86[624], line_85[622], line_84[620], line_83[618], line_82[616], line_81[614], line_80[612], line_79[610], line_78[608], line_77[606], line_76[604], line_75[602], line_74[600], line_73[598], line_72[596], line_71[594], line_70[592], line_69[590], line_68[588], line_67[586], line_66[584], line_65[582], line_64[580], line_63[578], line_62[576], line_61[574], line_60[572], line_59[570], line_58[568], line_57[566], line_56[564], line_55[562], line_54[560], line_53[558], line_52[556], line_51[554], line_50[552], line_49[550], line_48[548], line_47[546], line_46[544], line_45[542], line_44[540], line_43[538], line_42[536], line_41[534], line_40[532], line_39[530], line_38[528], line_37[526], line_36[524], line_35[522], line_34[520], line_33[518], line_32[516], line_31[514], line_30[512], line_29[510], line_28[508], line_27[506], line_26[504], line_25[502], line_24[500], line_23[498], line_22[496], line_21[494], line_20[492], line_19[490], line_18[488], line_17[486], line_16[484], line_15[482], line_14[480], line_13[478], line_12[476], line_11[474], line_10[472], line_9[470], line_8[468], line_7[466], line_6[464], line_5[462], line_4[460], line_3[458], line_2[456], line_1[454] };
assign col_709 = {line_128[709], line_127[707], line_126[705], line_125[703], line_124[701], line_123[699], line_122[697], line_121[695], line_120[693], line_119[691], line_118[689], line_117[687], line_116[685], line_115[683], line_114[681], line_113[679], line_112[677], line_111[675], line_110[673], line_109[671], line_108[669], line_107[667], line_106[665], line_105[663], line_104[661], line_103[659], line_102[657], line_101[655], line_100[653], line_99[651], line_98[649], line_97[647], line_96[645], line_95[643], line_94[641], line_93[639], line_92[637], line_91[635], line_90[633], line_89[631], line_88[629], line_87[627], line_86[625], line_85[623], line_84[621], line_83[619], line_82[617], line_81[615], line_80[613], line_79[611], line_78[609], line_77[607], line_76[605], line_75[603], line_74[601], line_73[599], line_72[597], line_71[595], line_70[593], line_69[591], line_68[589], line_67[587], line_66[585], line_65[583], line_64[581], line_63[579], line_62[577], line_61[575], line_60[573], line_59[571], line_58[569], line_57[567], line_56[565], line_55[563], line_54[561], line_53[559], line_52[557], line_51[555], line_50[553], line_49[551], line_48[549], line_47[547], line_46[545], line_45[543], line_44[541], line_43[539], line_42[537], line_41[535], line_40[533], line_39[531], line_38[529], line_37[527], line_36[525], line_35[523], line_34[521], line_33[519], line_32[517], line_31[515], line_30[513], line_29[511], line_28[509], line_27[507], line_26[505], line_25[503], line_24[501], line_23[499], line_22[497], line_21[495], line_20[493], line_19[491], line_18[489], line_17[487], line_16[485], line_15[483], line_14[481], line_13[479], line_12[477], line_11[475], line_10[473], line_9[471], line_8[469], line_7[467], line_6[465], line_5[463], line_4[461], line_3[459], line_2[457], line_1[455] };
assign col_710 = {line_128[710], line_127[708], line_126[706], line_125[704], line_124[702], line_123[700], line_122[698], line_121[696], line_120[694], line_119[692], line_118[690], line_117[688], line_116[686], line_115[684], line_114[682], line_113[680], line_112[678], line_111[676], line_110[674], line_109[672], line_108[670], line_107[668], line_106[666], line_105[664], line_104[662], line_103[660], line_102[658], line_101[656], line_100[654], line_99[652], line_98[650], line_97[648], line_96[646], line_95[644], line_94[642], line_93[640], line_92[638], line_91[636], line_90[634], line_89[632], line_88[630], line_87[628], line_86[626], line_85[624], line_84[622], line_83[620], line_82[618], line_81[616], line_80[614], line_79[612], line_78[610], line_77[608], line_76[606], line_75[604], line_74[602], line_73[600], line_72[598], line_71[596], line_70[594], line_69[592], line_68[590], line_67[588], line_66[586], line_65[584], line_64[582], line_63[580], line_62[578], line_61[576], line_60[574], line_59[572], line_58[570], line_57[568], line_56[566], line_55[564], line_54[562], line_53[560], line_52[558], line_51[556], line_50[554], line_49[552], line_48[550], line_47[548], line_46[546], line_45[544], line_44[542], line_43[540], line_42[538], line_41[536], line_40[534], line_39[532], line_38[530], line_37[528], line_36[526], line_35[524], line_34[522], line_33[520], line_32[518], line_31[516], line_30[514], line_29[512], line_28[510], line_27[508], line_26[506], line_25[504], line_24[502], line_23[500], line_22[498], line_21[496], line_20[494], line_19[492], line_18[490], line_17[488], line_16[486], line_15[484], line_14[482], line_13[480], line_12[478], line_11[476], line_10[474], line_9[472], line_8[470], line_7[468], line_6[466], line_5[464], line_4[462], line_3[460], line_2[458], line_1[456] };
assign col_711 = {line_128[711], line_127[709], line_126[707], line_125[705], line_124[703], line_123[701], line_122[699], line_121[697], line_120[695], line_119[693], line_118[691], line_117[689], line_116[687], line_115[685], line_114[683], line_113[681], line_112[679], line_111[677], line_110[675], line_109[673], line_108[671], line_107[669], line_106[667], line_105[665], line_104[663], line_103[661], line_102[659], line_101[657], line_100[655], line_99[653], line_98[651], line_97[649], line_96[647], line_95[645], line_94[643], line_93[641], line_92[639], line_91[637], line_90[635], line_89[633], line_88[631], line_87[629], line_86[627], line_85[625], line_84[623], line_83[621], line_82[619], line_81[617], line_80[615], line_79[613], line_78[611], line_77[609], line_76[607], line_75[605], line_74[603], line_73[601], line_72[599], line_71[597], line_70[595], line_69[593], line_68[591], line_67[589], line_66[587], line_65[585], line_64[583], line_63[581], line_62[579], line_61[577], line_60[575], line_59[573], line_58[571], line_57[569], line_56[567], line_55[565], line_54[563], line_53[561], line_52[559], line_51[557], line_50[555], line_49[553], line_48[551], line_47[549], line_46[547], line_45[545], line_44[543], line_43[541], line_42[539], line_41[537], line_40[535], line_39[533], line_38[531], line_37[529], line_36[527], line_35[525], line_34[523], line_33[521], line_32[519], line_31[517], line_30[515], line_29[513], line_28[511], line_27[509], line_26[507], line_25[505], line_24[503], line_23[501], line_22[499], line_21[497], line_20[495], line_19[493], line_18[491], line_17[489], line_16[487], line_15[485], line_14[483], line_13[481], line_12[479], line_11[477], line_10[475], line_9[473], line_8[471], line_7[469], line_6[467], line_5[465], line_4[463], line_3[461], line_2[459], line_1[457] };
assign col_712 = {line_128[712], line_127[710], line_126[708], line_125[706], line_124[704], line_123[702], line_122[700], line_121[698], line_120[696], line_119[694], line_118[692], line_117[690], line_116[688], line_115[686], line_114[684], line_113[682], line_112[680], line_111[678], line_110[676], line_109[674], line_108[672], line_107[670], line_106[668], line_105[666], line_104[664], line_103[662], line_102[660], line_101[658], line_100[656], line_99[654], line_98[652], line_97[650], line_96[648], line_95[646], line_94[644], line_93[642], line_92[640], line_91[638], line_90[636], line_89[634], line_88[632], line_87[630], line_86[628], line_85[626], line_84[624], line_83[622], line_82[620], line_81[618], line_80[616], line_79[614], line_78[612], line_77[610], line_76[608], line_75[606], line_74[604], line_73[602], line_72[600], line_71[598], line_70[596], line_69[594], line_68[592], line_67[590], line_66[588], line_65[586], line_64[584], line_63[582], line_62[580], line_61[578], line_60[576], line_59[574], line_58[572], line_57[570], line_56[568], line_55[566], line_54[564], line_53[562], line_52[560], line_51[558], line_50[556], line_49[554], line_48[552], line_47[550], line_46[548], line_45[546], line_44[544], line_43[542], line_42[540], line_41[538], line_40[536], line_39[534], line_38[532], line_37[530], line_36[528], line_35[526], line_34[524], line_33[522], line_32[520], line_31[518], line_30[516], line_29[514], line_28[512], line_27[510], line_26[508], line_25[506], line_24[504], line_23[502], line_22[500], line_21[498], line_20[496], line_19[494], line_18[492], line_17[490], line_16[488], line_15[486], line_14[484], line_13[482], line_12[480], line_11[478], line_10[476], line_9[474], line_8[472], line_7[470], line_6[468], line_5[466], line_4[464], line_3[462], line_2[460], line_1[458] };
assign col_713 = {line_128[713], line_127[711], line_126[709], line_125[707], line_124[705], line_123[703], line_122[701], line_121[699], line_120[697], line_119[695], line_118[693], line_117[691], line_116[689], line_115[687], line_114[685], line_113[683], line_112[681], line_111[679], line_110[677], line_109[675], line_108[673], line_107[671], line_106[669], line_105[667], line_104[665], line_103[663], line_102[661], line_101[659], line_100[657], line_99[655], line_98[653], line_97[651], line_96[649], line_95[647], line_94[645], line_93[643], line_92[641], line_91[639], line_90[637], line_89[635], line_88[633], line_87[631], line_86[629], line_85[627], line_84[625], line_83[623], line_82[621], line_81[619], line_80[617], line_79[615], line_78[613], line_77[611], line_76[609], line_75[607], line_74[605], line_73[603], line_72[601], line_71[599], line_70[597], line_69[595], line_68[593], line_67[591], line_66[589], line_65[587], line_64[585], line_63[583], line_62[581], line_61[579], line_60[577], line_59[575], line_58[573], line_57[571], line_56[569], line_55[567], line_54[565], line_53[563], line_52[561], line_51[559], line_50[557], line_49[555], line_48[553], line_47[551], line_46[549], line_45[547], line_44[545], line_43[543], line_42[541], line_41[539], line_40[537], line_39[535], line_38[533], line_37[531], line_36[529], line_35[527], line_34[525], line_33[523], line_32[521], line_31[519], line_30[517], line_29[515], line_28[513], line_27[511], line_26[509], line_25[507], line_24[505], line_23[503], line_22[501], line_21[499], line_20[497], line_19[495], line_18[493], line_17[491], line_16[489], line_15[487], line_14[485], line_13[483], line_12[481], line_11[479], line_10[477], line_9[475], line_8[473], line_7[471], line_6[469], line_5[467], line_4[465], line_3[463], line_2[461], line_1[459] };
assign col_714 = {line_128[714], line_127[712], line_126[710], line_125[708], line_124[706], line_123[704], line_122[702], line_121[700], line_120[698], line_119[696], line_118[694], line_117[692], line_116[690], line_115[688], line_114[686], line_113[684], line_112[682], line_111[680], line_110[678], line_109[676], line_108[674], line_107[672], line_106[670], line_105[668], line_104[666], line_103[664], line_102[662], line_101[660], line_100[658], line_99[656], line_98[654], line_97[652], line_96[650], line_95[648], line_94[646], line_93[644], line_92[642], line_91[640], line_90[638], line_89[636], line_88[634], line_87[632], line_86[630], line_85[628], line_84[626], line_83[624], line_82[622], line_81[620], line_80[618], line_79[616], line_78[614], line_77[612], line_76[610], line_75[608], line_74[606], line_73[604], line_72[602], line_71[600], line_70[598], line_69[596], line_68[594], line_67[592], line_66[590], line_65[588], line_64[586], line_63[584], line_62[582], line_61[580], line_60[578], line_59[576], line_58[574], line_57[572], line_56[570], line_55[568], line_54[566], line_53[564], line_52[562], line_51[560], line_50[558], line_49[556], line_48[554], line_47[552], line_46[550], line_45[548], line_44[546], line_43[544], line_42[542], line_41[540], line_40[538], line_39[536], line_38[534], line_37[532], line_36[530], line_35[528], line_34[526], line_33[524], line_32[522], line_31[520], line_30[518], line_29[516], line_28[514], line_27[512], line_26[510], line_25[508], line_24[506], line_23[504], line_22[502], line_21[500], line_20[498], line_19[496], line_18[494], line_17[492], line_16[490], line_15[488], line_14[486], line_13[484], line_12[482], line_11[480], line_10[478], line_9[476], line_8[474], line_7[472], line_6[470], line_5[468], line_4[466], line_3[464], line_2[462], line_1[460] };
assign col_715 = {line_128[715], line_127[713], line_126[711], line_125[709], line_124[707], line_123[705], line_122[703], line_121[701], line_120[699], line_119[697], line_118[695], line_117[693], line_116[691], line_115[689], line_114[687], line_113[685], line_112[683], line_111[681], line_110[679], line_109[677], line_108[675], line_107[673], line_106[671], line_105[669], line_104[667], line_103[665], line_102[663], line_101[661], line_100[659], line_99[657], line_98[655], line_97[653], line_96[651], line_95[649], line_94[647], line_93[645], line_92[643], line_91[641], line_90[639], line_89[637], line_88[635], line_87[633], line_86[631], line_85[629], line_84[627], line_83[625], line_82[623], line_81[621], line_80[619], line_79[617], line_78[615], line_77[613], line_76[611], line_75[609], line_74[607], line_73[605], line_72[603], line_71[601], line_70[599], line_69[597], line_68[595], line_67[593], line_66[591], line_65[589], line_64[587], line_63[585], line_62[583], line_61[581], line_60[579], line_59[577], line_58[575], line_57[573], line_56[571], line_55[569], line_54[567], line_53[565], line_52[563], line_51[561], line_50[559], line_49[557], line_48[555], line_47[553], line_46[551], line_45[549], line_44[547], line_43[545], line_42[543], line_41[541], line_40[539], line_39[537], line_38[535], line_37[533], line_36[531], line_35[529], line_34[527], line_33[525], line_32[523], line_31[521], line_30[519], line_29[517], line_28[515], line_27[513], line_26[511], line_25[509], line_24[507], line_23[505], line_22[503], line_21[501], line_20[499], line_19[497], line_18[495], line_17[493], line_16[491], line_15[489], line_14[487], line_13[485], line_12[483], line_11[481], line_10[479], line_9[477], line_8[475], line_7[473], line_6[471], line_5[469], line_4[467], line_3[465], line_2[463], line_1[461] };
assign col_716 = {line_128[716], line_127[714], line_126[712], line_125[710], line_124[708], line_123[706], line_122[704], line_121[702], line_120[700], line_119[698], line_118[696], line_117[694], line_116[692], line_115[690], line_114[688], line_113[686], line_112[684], line_111[682], line_110[680], line_109[678], line_108[676], line_107[674], line_106[672], line_105[670], line_104[668], line_103[666], line_102[664], line_101[662], line_100[660], line_99[658], line_98[656], line_97[654], line_96[652], line_95[650], line_94[648], line_93[646], line_92[644], line_91[642], line_90[640], line_89[638], line_88[636], line_87[634], line_86[632], line_85[630], line_84[628], line_83[626], line_82[624], line_81[622], line_80[620], line_79[618], line_78[616], line_77[614], line_76[612], line_75[610], line_74[608], line_73[606], line_72[604], line_71[602], line_70[600], line_69[598], line_68[596], line_67[594], line_66[592], line_65[590], line_64[588], line_63[586], line_62[584], line_61[582], line_60[580], line_59[578], line_58[576], line_57[574], line_56[572], line_55[570], line_54[568], line_53[566], line_52[564], line_51[562], line_50[560], line_49[558], line_48[556], line_47[554], line_46[552], line_45[550], line_44[548], line_43[546], line_42[544], line_41[542], line_40[540], line_39[538], line_38[536], line_37[534], line_36[532], line_35[530], line_34[528], line_33[526], line_32[524], line_31[522], line_30[520], line_29[518], line_28[516], line_27[514], line_26[512], line_25[510], line_24[508], line_23[506], line_22[504], line_21[502], line_20[500], line_19[498], line_18[496], line_17[494], line_16[492], line_15[490], line_14[488], line_13[486], line_12[484], line_11[482], line_10[480], line_9[478], line_8[476], line_7[474], line_6[472], line_5[470], line_4[468], line_3[466], line_2[464], line_1[462] };
assign col_717 = {line_128[717], line_127[715], line_126[713], line_125[711], line_124[709], line_123[707], line_122[705], line_121[703], line_120[701], line_119[699], line_118[697], line_117[695], line_116[693], line_115[691], line_114[689], line_113[687], line_112[685], line_111[683], line_110[681], line_109[679], line_108[677], line_107[675], line_106[673], line_105[671], line_104[669], line_103[667], line_102[665], line_101[663], line_100[661], line_99[659], line_98[657], line_97[655], line_96[653], line_95[651], line_94[649], line_93[647], line_92[645], line_91[643], line_90[641], line_89[639], line_88[637], line_87[635], line_86[633], line_85[631], line_84[629], line_83[627], line_82[625], line_81[623], line_80[621], line_79[619], line_78[617], line_77[615], line_76[613], line_75[611], line_74[609], line_73[607], line_72[605], line_71[603], line_70[601], line_69[599], line_68[597], line_67[595], line_66[593], line_65[591], line_64[589], line_63[587], line_62[585], line_61[583], line_60[581], line_59[579], line_58[577], line_57[575], line_56[573], line_55[571], line_54[569], line_53[567], line_52[565], line_51[563], line_50[561], line_49[559], line_48[557], line_47[555], line_46[553], line_45[551], line_44[549], line_43[547], line_42[545], line_41[543], line_40[541], line_39[539], line_38[537], line_37[535], line_36[533], line_35[531], line_34[529], line_33[527], line_32[525], line_31[523], line_30[521], line_29[519], line_28[517], line_27[515], line_26[513], line_25[511], line_24[509], line_23[507], line_22[505], line_21[503], line_20[501], line_19[499], line_18[497], line_17[495], line_16[493], line_15[491], line_14[489], line_13[487], line_12[485], line_11[483], line_10[481], line_9[479], line_8[477], line_7[475], line_6[473], line_5[471], line_4[469], line_3[467], line_2[465], line_1[463] };
assign col_718 = {line_128[718], line_127[716], line_126[714], line_125[712], line_124[710], line_123[708], line_122[706], line_121[704], line_120[702], line_119[700], line_118[698], line_117[696], line_116[694], line_115[692], line_114[690], line_113[688], line_112[686], line_111[684], line_110[682], line_109[680], line_108[678], line_107[676], line_106[674], line_105[672], line_104[670], line_103[668], line_102[666], line_101[664], line_100[662], line_99[660], line_98[658], line_97[656], line_96[654], line_95[652], line_94[650], line_93[648], line_92[646], line_91[644], line_90[642], line_89[640], line_88[638], line_87[636], line_86[634], line_85[632], line_84[630], line_83[628], line_82[626], line_81[624], line_80[622], line_79[620], line_78[618], line_77[616], line_76[614], line_75[612], line_74[610], line_73[608], line_72[606], line_71[604], line_70[602], line_69[600], line_68[598], line_67[596], line_66[594], line_65[592], line_64[590], line_63[588], line_62[586], line_61[584], line_60[582], line_59[580], line_58[578], line_57[576], line_56[574], line_55[572], line_54[570], line_53[568], line_52[566], line_51[564], line_50[562], line_49[560], line_48[558], line_47[556], line_46[554], line_45[552], line_44[550], line_43[548], line_42[546], line_41[544], line_40[542], line_39[540], line_38[538], line_37[536], line_36[534], line_35[532], line_34[530], line_33[528], line_32[526], line_31[524], line_30[522], line_29[520], line_28[518], line_27[516], line_26[514], line_25[512], line_24[510], line_23[508], line_22[506], line_21[504], line_20[502], line_19[500], line_18[498], line_17[496], line_16[494], line_15[492], line_14[490], line_13[488], line_12[486], line_11[484], line_10[482], line_9[480], line_8[478], line_7[476], line_6[474], line_5[472], line_4[470], line_3[468], line_2[466], line_1[464] };
assign col_719 = {line_128[719], line_127[717], line_126[715], line_125[713], line_124[711], line_123[709], line_122[707], line_121[705], line_120[703], line_119[701], line_118[699], line_117[697], line_116[695], line_115[693], line_114[691], line_113[689], line_112[687], line_111[685], line_110[683], line_109[681], line_108[679], line_107[677], line_106[675], line_105[673], line_104[671], line_103[669], line_102[667], line_101[665], line_100[663], line_99[661], line_98[659], line_97[657], line_96[655], line_95[653], line_94[651], line_93[649], line_92[647], line_91[645], line_90[643], line_89[641], line_88[639], line_87[637], line_86[635], line_85[633], line_84[631], line_83[629], line_82[627], line_81[625], line_80[623], line_79[621], line_78[619], line_77[617], line_76[615], line_75[613], line_74[611], line_73[609], line_72[607], line_71[605], line_70[603], line_69[601], line_68[599], line_67[597], line_66[595], line_65[593], line_64[591], line_63[589], line_62[587], line_61[585], line_60[583], line_59[581], line_58[579], line_57[577], line_56[575], line_55[573], line_54[571], line_53[569], line_52[567], line_51[565], line_50[563], line_49[561], line_48[559], line_47[557], line_46[555], line_45[553], line_44[551], line_43[549], line_42[547], line_41[545], line_40[543], line_39[541], line_38[539], line_37[537], line_36[535], line_35[533], line_34[531], line_33[529], line_32[527], line_31[525], line_30[523], line_29[521], line_28[519], line_27[517], line_26[515], line_25[513], line_24[511], line_23[509], line_22[507], line_21[505], line_20[503], line_19[501], line_18[499], line_17[497], line_16[495], line_15[493], line_14[491], line_13[489], line_12[487], line_11[485], line_10[483], line_9[481], line_8[479], line_7[477], line_6[475], line_5[473], line_4[471], line_3[469], line_2[467], line_1[465] };
assign col_720 = {line_128[720], line_127[718], line_126[716], line_125[714], line_124[712], line_123[710], line_122[708], line_121[706], line_120[704], line_119[702], line_118[700], line_117[698], line_116[696], line_115[694], line_114[692], line_113[690], line_112[688], line_111[686], line_110[684], line_109[682], line_108[680], line_107[678], line_106[676], line_105[674], line_104[672], line_103[670], line_102[668], line_101[666], line_100[664], line_99[662], line_98[660], line_97[658], line_96[656], line_95[654], line_94[652], line_93[650], line_92[648], line_91[646], line_90[644], line_89[642], line_88[640], line_87[638], line_86[636], line_85[634], line_84[632], line_83[630], line_82[628], line_81[626], line_80[624], line_79[622], line_78[620], line_77[618], line_76[616], line_75[614], line_74[612], line_73[610], line_72[608], line_71[606], line_70[604], line_69[602], line_68[600], line_67[598], line_66[596], line_65[594], line_64[592], line_63[590], line_62[588], line_61[586], line_60[584], line_59[582], line_58[580], line_57[578], line_56[576], line_55[574], line_54[572], line_53[570], line_52[568], line_51[566], line_50[564], line_49[562], line_48[560], line_47[558], line_46[556], line_45[554], line_44[552], line_43[550], line_42[548], line_41[546], line_40[544], line_39[542], line_38[540], line_37[538], line_36[536], line_35[534], line_34[532], line_33[530], line_32[528], line_31[526], line_30[524], line_29[522], line_28[520], line_27[518], line_26[516], line_25[514], line_24[512], line_23[510], line_22[508], line_21[506], line_20[504], line_19[502], line_18[500], line_17[498], line_16[496], line_15[494], line_14[492], line_13[490], line_12[488], line_11[486], line_10[484], line_9[482], line_8[480], line_7[478], line_6[476], line_5[474], line_4[472], line_3[470], line_2[468], line_1[466] };
assign col_721 = {line_128[721], line_127[719], line_126[717], line_125[715], line_124[713], line_123[711], line_122[709], line_121[707], line_120[705], line_119[703], line_118[701], line_117[699], line_116[697], line_115[695], line_114[693], line_113[691], line_112[689], line_111[687], line_110[685], line_109[683], line_108[681], line_107[679], line_106[677], line_105[675], line_104[673], line_103[671], line_102[669], line_101[667], line_100[665], line_99[663], line_98[661], line_97[659], line_96[657], line_95[655], line_94[653], line_93[651], line_92[649], line_91[647], line_90[645], line_89[643], line_88[641], line_87[639], line_86[637], line_85[635], line_84[633], line_83[631], line_82[629], line_81[627], line_80[625], line_79[623], line_78[621], line_77[619], line_76[617], line_75[615], line_74[613], line_73[611], line_72[609], line_71[607], line_70[605], line_69[603], line_68[601], line_67[599], line_66[597], line_65[595], line_64[593], line_63[591], line_62[589], line_61[587], line_60[585], line_59[583], line_58[581], line_57[579], line_56[577], line_55[575], line_54[573], line_53[571], line_52[569], line_51[567], line_50[565], line_49[563], line_48[561], line_47[559], line_46[557], line_45[555], line_44[553], line_43[551], line_42[549], line_41[547], line_40[545], line_39[543], line_38[541], line_37[539], line_36[537], line_35[535], line_34[533], line_33[531], line_32[529], line_31[527], line_30[525], line_29[523], line_28[521], line_27[519], line_26[517], line_25[515], line_24[513], line_23[511], line_22[509], line_21[507], line_20[505], line_19[503], line_18[501], line_17[499], line_16[497], line_15[495], line_14[493], line_13[491], line_12[489], line_11[487], line_10[485], line_9[483], line_8[481], line_7[479], line_6[477], line_5[475], line_4[473], line_3[471], line_2[469], line_1[467] };
assign col_722 = {line_128[722], line_127[720], line_126[718], line_125[716], line_124[714], line_123[712], line_122[710], line_121[708], line_120[706], line_119[704], line_118[702], line_117[700], line_116[698], line_115[696], line_114[694], line_113[692], line_112[690], line_111[688], line_110[686], line_109[684], line_108[682], line_107[680], line_106[678], line_105[676], line_104[674], line_103[672], line_102[670], line_101[668], line_100[666], line_99[664], line_98[662], line_97[660], line_96[658], line_95[656], line_94[654], line_93[652], line_92[650], line_91[648], line_90[646], line_89[644], line_88[642], line_87[640], line_86[638], line_85[636], line_84[634], line_83[632], line_82[630], line_81[628], line_80[626], line_79[624], line_78[622], line_77[620], line_76[618], line_75[616], line_74[614], line_73[612], line_72[610], line_71[608], line_70[606], line_69[604], line_68[602], line_67[600], line_66[598], line_65[596], line_64[594], line_63[592], line_62[590], line_61[588], line_60[586], line_59[584], line_58[582], line_57[580], line_56[578], line_55[576], line_54[574], line_53[572], line_52[570], line_51[568], line_50[566], line_49[564], line_48[562], line_47[560], line_46[558], line_45[556], line_44[554], line_43[552], line_42[550], line_41[548], line_40[546], line_39[544], line_38[542], line_37[540], line_36[538], line_35[536], line_34[534], line_33[532], line_32[530], line_31[528], line_30[526], line_29[524], line_28[522], line_27[520], line_26[518], line_25[516], line_24[514], line_23[512], line_22[510], line_21[508], line_20[506], line_19[504], line_18[502], line_17[500], line_16[498], line_15[496], line_14[494], line_13[492], line_12[490], line_11[488], line_10[486], line_9[484], line_8[482], line_7[480], line_6[478], line_5[476], line_4[474], line_3[472], line_2[470], line_1[468] };
assign col_723 = {line_128[723], line_127[721], line_126[719], line_125[717], line_124[715], line_123[713], line_122[711], line_121[709], line_120[707], line_119[705], line_118[703], line_117[701], line_116[699], line_115[697], line_114[695], line_113[693], line_112[691], line_111[689], line_110[687], line_109[685], line_108[683], line_107[681], line_106[679], line_105[677], line_104[675], line_103[673], line_102[671], line_101[669], line_100[667], line_99[665], line_98[663], line_97[661], line_96[659], line_95[657], line_94[655], line_93[653], line_92[651], line_91[649], line_90[647], line_89[645], line_88[643], line_87[641], line_86[639], line_85[637], line_84[635], line_83[633], line_82[631], line_81[629], line_80[627], line_79[625], line_78[623], line_77[621], line_76[619], line_75[617], line_74[615], line_73[613], line_72[611], line_71[609], line_70[607], line_69[605], line_68[603], line_67[601], line_66[599], line_65[597], line_64[595], line_63[593], line_62[591], line_61[589], line_60[587], line_59[585], line_58[583], line_57[581], line_56[579], line_55[577], line_54[575], line_53[573], line_52[571], line_51[569], line_50[567], line_49[565], line_48[563], line_47[561], line_46[559], line_45[557], line_44[555], line_43[553], line_42[551], line_41[549], line_40[547], line_39[545], line_38[543], line_37[541], line_36[539], line_35[537], line_34[535], line_33[533], line_32[531], line_31[529], line_30[527], line_29[525], line_28[523], line_27[521], line_26[519], line_25[517], line_24[515], line_23[513], line_22[511], line_21[509], line_20[507], line_19[505], line_18[503], line_17[501], line_16[499], line_15[497], line_14[495], line_13[493], line_12[491], line_11[489], line_10[487], line_9[485], line_8[483], line_7[481], line_6[479], line_5[477], line_4[475], line_3[473], line_2[471], line_1[469] };
assign col_724 = {line_128[724], line_127[722], line_126[720], line_125[718], line_124[716], line_123[714], line_122[712], line_121[710], line_120[708], line_119[706], line_118[704], line_117[702], line_116[700], line_115[698], line_114[696], line_113[694], line_112[692], line_111[690], line_110[688], line_109[686], line_108[684], line_107[682], line_106[680], line_105[678], line_104[676], line_103[674], line_102[672], line_101[670], line_100[668], line_99[666], line_98[664], line_97[662], line_96[660], line_95[658], line_94[656], line_93[654], line_92[652], line_91[650], line_90[648], line_89[646], line_88[644], line_87[642], line_86[640], line_85[638], line_84[636], line_83[634], line_82[632], line_81[630], line_80[628], line_79[626], line_78[624], line_77[622], line_76[620], line_75[618], line_74[616], line_73[614], line_72[612], line_71[610], line_70[608], line_69[606], line_68[604], line_67[602], line_66[600], line_65[598], line_64[596], line_63[594], line_62[592], line_61[590], line_60[588], line_59[586], line_58[584], line_57[582], line_56[580], line_55[578], line_54[576], line_53[574], line_52[572], line_51[570], line_50[568], line_49[566], line_48[564], line_47[562], line_46[560], line_45[558], line_44[556], line_43[554], line_42[552], line_41[550], line_40[548], line_39[546], line_38[544], line_37[542], line_36[540], line_35[538], line_34[536], line_33[534], line_32[532], line_31[530], line_30[528], line_29[526], line_28[524], line_27[522], line_26[520], line_25[518], line_24[516], line_23[514], line_22[512], line_21[510], line_20[508], line_19[506], line_18[504], line_17[502], line_16[500], line_15[498], line_14[496], line_13[494], line_12[492], line_11[490], line_10[488], line_9[486], line_8[484], line_7[482], line_6[480], line_5[478], line_4[476], line_3[474], line_2[472], line_1[470] };
assign col_725 = {line_128[725], line_127[723], line_126[721], line_125[719], line_124[717], line_123[715], line_122[713], line_121[711], line_120[709], line_119[707], line_118[705], line_117[703], line_116[701], line_115[699], line_114[697], line_113[695], line_112[693], line_111[691], line_110[689], line_109[687], line_108[685], line_107[683], line_106[681], line_105[679], line_104[677], line_103[675], line_102[673], line_101[671], line_100[669], line_99[667], line_98[665], line_97[663], line_96[661], line_95[659], line_94[657], line_93[655], line_92[653], line_91[651], line_90[649], line_89[647], line_88[645], line_87[643], line_86[641], line_85[639], line_84[637], line_83[635], line_82[633], line_81[631], line_80[629], line_79[627], line_78[625], line_77[623], line_76[621], line_75[619], line_74[617], line_73[615], line_72[613], line_71[611], line_70[609], line_69[607], line_68[605], line_67[603], line_66[601], line_65[599], line_64[597], line_63[595], line_62[593], line_61[591], line_60[589], line_59[587], line_58[585], line_57[583], line_56[581], line_55[579], line_54[577], line_53[575], line_52[573], line_51[571], line_50[569], line_49[567], line_48[565], line_47[563], line_46[561], line_45[559], line_44[557], line_43[555], line_42[553], line_41[551], line_40[549], line_39[547], line_38[545], line_37[543], line_36[541], line_35[539], line_34[537], line_33[535], line_32[533], line_31[531], line_30[529], line_29[527], line_28[525], line_27[523], line_26[521], line_25[519], line_24[517], line_23[515], line_22[513], line_21[511], line_20[509], line_19[507], line_18[505], line_17[503], line_16[501], line_15[499], line_14[497], line_13[495], line_12[493], line_11[491], line_10[489], line_9[487], line_8[485], line_7[483], line_6[481], line_5[479], line_4[477], line_3[475], line_2[473], line_1[471] };
assign col_726 = {line_128[726], line_127[724], line_126[722], line_125[720], line_124[718], line_123[716], line_122[714], line_121[712], line_120[710], line_119[708], line_118[706], line_117[704], line_116[702], line_115[700], line_114[698], line_113[696], line_112[694], line_111[692], line_110[690], line_109[688], line_108[686], line_107[684], line_106[682], line_105[680], line_104[678], line_103[676], line_102[674], line_101[672], line_100[670], line_99[668], line_98[666], line_97[664], line_96[662], line_95[660], line_94[658], line_93[656], line_92[654], line_91[652], line_90[650], line_89[648], line_88[646], line_87[644], line_86[642], line_85[640], line_84[638], line_83[636], line_82[634], line_81[632], line_80[630], line_79[628], line_78[626], line_77[624], line_76[622], line_75[620], line_74[618], line_73[616], line_72[614], line_71[612], line_70[610], line_69[608], line_68[606], line_67[604], line_66[602], line_65[600], line_64[598], line_63[596], line_62[594], line_61[592], line_60[590], line_59[588], line_58[586], line_57[584], line_56[582], line_55[580], line_54[578], line_53[576], line_52[574], line_51[572], line_50[570], line_49[568], line_48[566], line_47[564], line_46[562], line_45[560], line_44[558], line_43[556], line_42[554], line_41[552], line_40[550], line_39[548], line_38[546], line_37[544], line_36[542], line_35[540], line_34[538], line_33[536], line_32[534], line_31[532], line_30[530], line_29[528], line_28[526], line_27[524], line_26[522], line_25[520], line_24[518], line_23[516], line_22[514], line_21[512], line_20[510], line_19[508], line_18[506], line_17[504], line_16[502], line_15[500], line_14[498], line_13[496], line_12[494], line_11[492], line_10[490], line_9[488], line_8[486], line_7[484], line_6[482], line_5[480], line_4[478], line_3[476], line_2[474], line_1[472] };
assign col_727 = {line_128[727], line_127[725], line_126[723], line_125[721], line_124[719], line_123[717], line_122[715], line_121[713], line_120[711], line_119[709], line_118[707], line_117[705], line_116[703], line_115[701], line_114[699], line_113[697], line_112[695], line_111[693], line_110[691], line_109[689], line_108[687], line_107[685], line_106[683], line_105[681], line_104[679], line_103[677], line_102[675], line_101[673], line_100[671], line_99[669], line_98[667], line_97[665], line_96[663], line_95[661], line_94[659], line_93[657], line_92[655], line_91[653], line_90[651], line_89[649], line_88[647], line_87[645], line_86[643], line_85[641], line_84[639], line_83[637], line_82[635], line_81[633], line_80[631], line_79[629], line_78[627], line_77[625], line_76[623], line_75[621], line_74[619], line_73[617], line_72[615], line_71[613], line_70[611], line_69[609], line_68[607], line_67[605], line_66[603], line_65[601], line_64[599], line_63[597], line_62[595], line_61[593], line_60[591], line_59[589], line_58[587], line_57[585], line_56[583], line_55[581], line_54[579], line_53[577], line_52[575], line_51[573], line_50[571], line_49[569], line_48[567], line_47[565], line_46[563], line_45[561], line_44[559], line_43[557], line_42[555], line_41[553], line_40[551], line_39[549], line_38[547], line_37[545], line_36[543], line_35[541], line_34[539], line_33[537], line_32[535], line_31[533], line_30[531], line_29[529], line_28[527], line_27[525], line_26[523], line_25[521], line_24[519], line_23[517], line_22[515], line_21[513], line_20[511], line_19[509], line_18[507], line_17[505], line_16[503], line_15[501], line_14[499], line_13[497], line_12[495], line_11[493], line_10[491], line_9[489], line_8[487], line_7[485], line_6[483], line_5[481], line_4[479], line_3[477], line_2[475], line_1[473] };
assign col_728 = {line_128[728], line_127[726], line_126[724], line_125[722], line_124[720], line_123[718], line_122[716], line_121[714], line_120[712], line_119[710], line_118[708], line_117[706], line_116[704], line_115[702], line_114[700], line_113[698], line_112[696], line_111[694], line_110[692], line_109[690], line_108[688], line_107[686], line_106[684], line_105[682], line_104[680], line_103[678], line_102[676], line_101[674], line_100[672], line_99[670], line_98[668], line_97[666], line_96[664], line_95[662], line_94[660], line_93[658], line_92[656], line_91[654], line_90[652], line_89[650], line_88[648], line_87[646], line_86[644], line_85[642], line_84[640], line_83[638], line_82[636], line_81[634], line_80[632], line_79[630], line_78[628], line_77[626], line_76[624], line_75[622], line_74[620], line_73[618], line_72[616], line_71[614], line_70[612], line_69[610], line_68[608], line_67[606], line_66[604], line_65[602], line_64[600], line_63[598], line_62[596], line_61[594], line_60[592], line_59[590], line_58[588], line_57[586], line_56[584], line_55[582], line_54[580], line_53[578], line_52[576], line_51[574], line_50[572], line_49[570], line_48[568], line_47[566], line_46[564], line_45[562], line_44[560], line_43[558], line_42[556], line_41[554], line_40[552], line_39[550], line_38[548], line_37[546], line_36[544], line_35[542], line_34[540], line_33[538], line_32[536], line_31[534], line_30[532], line_29[530], line_28[528], line_27[526], line_26[524], line_25[522], line_24[520], line_23[518], line_22[516], line_21[514], line_20[512], line_19[510], line_18[508], line_17[506], line_16[504], line_15[502], line_14[500], line_13[498], line_12[496], line_11[494], line_10[492], line_9[490], line_8[488], line_7[486], line_6[484], line_5[482], line_4[480], line_3[478], line_2[476], line_1[474] };
assign col_729 = {line_128[729], line_127[727], line_126[725], line_125[723], line_124[721], line_123[719], line_122[717], line_121[715], line_120[713], line_119[711], line_118[709], line_117[707], line_116[705], line_115[703], line_114[701], line_113[699], line_112[697], line_111[695], line_110[693], line_109[691], line_108[689], line_107[687], line_106[685], line_105[683], line_104[681], line_103[679], line_102[677], line_101[675], line_100[673], line_99[671], line_98[669], line_97[667], line_96[665], line_95[663], line_94[661], line_93[659], line_92[657], line_91[655], line_90[653], line_89[651], line_88[649], line_87[647], line_86[645], line_85[643], line_84[641], line_83[639], line_82[637], line_81[635], line_80[633], line_79[631], line_78[629], line_77[627], line_76[625], line_75[623], line_74[621], line_73[619], line_72[617], line_71[615], line_70[613], line_69[611], line_68[609], line_67[607], line_66[605], line_65[603], line_64[601], line_63[599], line_62[597], line_61[595], line_60[593], line_59[591], line_58[589], line_57[587], line_56[585], line_55[583], line_54[581], line_53[579], line_52[577], line_51[575], line_50[573], line_49[571], line_48[569], line_47[567], line_46[565], line_45[563], line_44[561], line_43[559], line_42[557], line_41[555], line_40[553], line_39[551], line_38[549], line_37[547], line_36[545], line_35[543], line_34[541], line_33[539], line_32[537], line_31[535], line_30[533], line_29[531], line_28[529], line_27[527], line_26[525], line_25[523], line_24[521], line_23[519], line_22[517], line_21[515], line_20[513], line_19[511], line_18[509], line_17[507], line_16[505], line_15[503], line_14[501], line_13[499], line_12[497], line_11[495], line_10[493], line_9[491], line_8[489], line_7[487], line_6[485], line_5[483], line_4[481], line_3[479], line_2[477], line_1[475] };
assign col_730 = {line_128[730], line_127[728], line_126[726], line_125[724], line_124[722], line_123[720], line_122[718], line_121[716], line_120[714], line_119[712], line_118[710], line_117[708], line_116[706], line_115[704], line_114[702], line_113[700], line_112[698], line_111[696], line_110[694], line_109[692], line_108[690], line_107[688], line_106[686], line_105[684], line_104[682], line_103[680], line_102[678], line_101[676], line_100[674], line_99[672], line_98[670], line_97[668], line_96[666], line_95[664], line_94[662], line_93[660], line_92[658], line_91[656], line_90[654], line_89[652], line_88[650], line_87[648], line_86[646], line_85[644], line_84[642], line_83[640], line_82[638], line_81[636], line_80[634], line_79[632], line_78[630], line_77[628], line_76[626], line_75[624], line_74[622], line_73[620], line_72[618], line_71[616], line_70[614], line_69[612], line_68[610], line_67[608], line_66[606], line_65[604], line_64[602], line_63[600], line_62[598], line_61[596], line_60[594], line_59[592], line_58[590], line_57[588], line_56[586], line_55[584], line_54[582], line_53[580], line_52[578], line_51[576], line_50[574], line_49[572], line_48[570], line_47[568], line_46[566], line_45[564], line_44[562], line_43[560], line_42[558], line_41[556], line_40[554], line_39[552], line_38[550], line_37[548], line_36[546], line_35[544], line_34[542], line_33[540], line_32[538], line_31[536], line_30[534], line_29[532], line_28[530], line_27[528], line_26[526], line_25[524], line_24[522], line_23[520], line_22[518], line_21[516], line_20[514], line_19[512], line_18[510], line_17[508], line_16[506], line_15[504], line_14[502], line_13[500], line_12[498], line_11[496], line_10[494], line_9[492], line_8[490], line_7[488], line_6[486], line_5[484], line_4[482], line_3[480], line_2[478], line_1[476] };
assign col_731 = {line_128[731], line_127[729], line_126[727], line_125[725], line_124[723], line_123[721], line_122[719], line_121[717], line_120[715], line_119[713], line_118[711], line_117[709], line_116[707], line_115[705], line_114[703], line_113[701], line_112[699], line_111[697], line_110[695], line_109[693], line_108[691], line_107[689], line_106[687], line_105[685], line_104[683], line_103[681], line_102[679], line_101[677], line_100[675], line_99[673], line_98[671], line_97[669], line_96[667], line_95[665], line_94[663], line_93[661], line_92[659], line_91[657], line_90[655], line_89[653], line_88[651], line_87[649], line_86[647], line_85[645], line_84[643], line_83[641], line_82[639], line_81[637], line_80[635], line_79[633], line_78[631], line_77[629], line_76[627], line_75[625], line_74[623], line_73[621], line_72[619], line_71[617], line_70[615], line_69[613], line_68[611], line_67[609], line_66[607], line_65[605], line_64[603], line_63[601], line_62[599], line_61[597], line_60[595], line_59[593], line_58[591], line_57[589], line_56[587], line_55[585], line_54[583], line_53[581], line_52[579], line_51[577], line_50[575], line_49[573], line_48[571], line_47[569], line_46[567], line_45[565], line_44[563], line_43[561], line_42[559], line_41[557], line_40[555], line_39[553], line_38[551], line_37[549], line_36[547], line_35[545], line_34[543], line_33[541], line_32[539], line_31[537], line_30[535], line_29[533], line_28[531], line_27[529], line_26[527], line_25[525], line_24[523], line_23[521], line_22[519], line_21[517], line_20[515], line_19[513], line_18[511], line_17[509], line_16[507], line_15[505], line_14[503], line_13[501], line_12[499], line_11[497], line_10[495], line_9[493], line_8[491], line_7[489], line_6[487], line_5[485], line_4[483], line_3[481], line_2[479], line_1[477] };
assign col_732 = {line_128[732], line_127[730], line_126[728], line_125[726], line_124[724], line_123[722], line_122[720], line_121[718], line_120[716], line_119[714], line_118[712], line_117[710], line_116[708], line_115[706], line_114[704], line_113[702], line_112[700], line_111[698], line_110[696], line_109[694], line_108[692], line_107[690], line_106[688], line_105[686], line_104[684], line_103[682], line_102[680], line_101[678], line_100[676], line_99[674], line_98[672], line_97[670], line_96[668], line_95[666], line_94[664], line_93[662], line_92[660], line_91[658], line_90[656], line_89[654], line_88[652], line_87[650], line_86[648], line_85[646], line_84[644], line_83[642], line_82[640], line_81[638], line_80[636], line_79[634], line_78[632], line_77[630], line_76[628], line_75[626], line_74[624], line_73[622], line_72[620], line_71[618], line_70[616], line_69[614], line_68[612], line_67[610], line_66[608], line_65[606], line_64[604], line_63[602], line_62[600], line_61[598], line_60[596], line_59[594], line_58[592], line_57[590], line_56[588], line_55[586], line_54[584], line_53[582], line_52[580], line_51[578], line_50[576], line_49[574], line_48[572], line_47[570], line_46[568], line_45[566], line_44[564], line_43[562], line_42[560], line_41[558], line_40[556], line_39[554], line_38[552], line_37[550], line_36[548], line_35[546], line_34[544], line_33[542], line_32[540], line_31[538], line_30[536], line_29[534], line_28[532], line_27[530], line_26[528], line_25[526], line_24[524], line_23[522], line_22[520], line_21[518], line_20[516], line_19[514], line_18[512], line_17[510], line_16[508], line_15[506], line_14[504], line_13[502], line_12[500], line_11[498], line_10[496], line_9[494], line_8[492], line_7[490], line_6[488], line_5[486], line_4[484], line_3[482], line_2[480], line_1[478] };
assign col_733 = {line_128[733], line_127[731], line_126[729], line_125[727], line_124[725], line_123[723], line_122[721], line_121[719], line_120[717], line_119[715], line_118[713], line_117[711], line_116[709], line_115[707], line_114[705], line_113[703], line_112[701], line_111[699], line_110[697], line_109[695], line_108[693], line_107[691], line_106[689], line_105[687], line_104[685], line_103[683], line_102[681], line_101[679], line_100[677], line_99[675], line_98[673], line_97[671], line_96[669], line_95[667], line_94[665], line_93[663], line_92[661], line_91[659], line_90[657], line_89[655], line_88[653], line_87[651], line_86[649], line_85[647], line_84[645], line_83[643], line_82[641], line_81[639], line_80[637], line_79[635], line_78[633], line_77[631], line_76[629], line_75[627], line_74[625], line_73[623], line_72[621], line_71[619], line_70[617], line_69[615], line_68[613], line_67[611], line_66[609], line_65[607], line_64[605], line_63[603], line_62[601], line_61[599], line_60[597], line_59[595], line_58[593], line_57[591], line_56[589], line_55[587], line_54[585], line_53[583], line_52[581], line_51[579], line_50[577], line_49[575], line_48[573], line_47[571], line_46[569], line_45[567], line_44[565], line_43[563], line_42[561], line_41[559], line_40[557], line_39[555], line_38[553], line_37[551], line_36[549], line_35[547], line_34[545], line_33[543], line_32[541], line_31[539], line_30[537], line_29[535], line_28[533], line_27[531], line_26[529], line_25[527], line_24[525], line_23[523], line_22[521], line_21[519], line_20[517], line_19[515], line_18[513], line_17[511], line_16[509], line_15[507], line_14[505], line_13[503], line_12[501], line_11[499], line_10[497], line_9[495], line_8[493], line_7[491], line_6[489], line_5[487], line_4[485], line_3[483], line_2[481], line_1[479] };
assign col_734 = {line_128[734], line_127[732], line_126[730], line_125[728], line_124[726], line_123[724], line_122[722], line_121[720], line_120[718], line_119[716], line_118[714], line_117[712], line_116[710], line_115[708], line_114[706], line_113[704], line_112[702], line_111[700], line_110[698], line_109[696], line_108[694], line_107[692], line_106[690], line_105[688], line_104[686], line_103[684], line_102[682], line_101[680], line_100[678], line_99[676], line_98[674], line_97[672], line_96[670], line_95[668], line_94[666], line_93[664], line_92[662], line_91[660], line_90[658], line_89[656], line_88[654], line_87[652], line_86[650], line_85[648], line_84[646], line_83[644], line_82[642], line_81[640], line_80[638], line_79[636], line_78[634], line_77[632], line_76[630], line_75[628], line_74[626], line_73[624], line_72[622], line_71[620], line_70[618], line_69[616], line_68[614], line_67[612], line_66[610], line_65[608], line_64[606], line_63[604], line_62[602], line_61[600], line_60[598], line_59[596], line_58[594], line_57[592], line_56[590], line_55[588], line_54[586], line_53[584], line_52[582], line_51[580], line_50[578], line_49[576], line_48[574], line_47[572], line_46[570], line_45[568], line_44[566], line_43[564], line_42[562], line_41[560], line_40[558], line_39[556], line_38[554], line_37[552], line_36[550], line_35[548], line_34[546], line_33[544], line_32[542], line_31[540], line_30[538], line_29[536], line_28[534], line_27[532], line_26[530], line_25[528], line_24[526], line_23[524], line_22[522], line_21[520], line_20[518], line_19[516], line_18[514], line_17[512], line_16[510], line_15[508], line_14[506], line_13[504], line_12[502], line_11[500], line_10[498], line_9[496], line_8[494], line_7[492], line_6[490], line_5[488], line_4[486], line_3[484], line_2[482], line_1[480] };
assign col_735 = {line_128[735], line_127[733], line_126[731], line_125[729], line_124[727], line_123[725], line_122[723], line_121[721], line_120[719], line_119[717], line_118[715], line_117[713], line_116[711], line_115[709], line_114[707], line_113[705], line_112[703], line_111[701], line_110[699], line_109[697], line_108[695], line_107[693], line_106[691], line_105[689], line_104[687], line_103[685], line_102[683], line_101[681], line_100[679], line_99[677], line_98[675], line_97[673], line_96[671], line_95[669], line_94[667], line_93[665], line_92[663], line_91[661], line_90[659], line_89[657], line_88[655], line_87[653], line_86[651], line_85[649], line_84[647], line_83[645], line_82[643], line_81[641], line_80[639], line_79[637], line_78[635], line_77[633], line_76[631], line_75[629], line_74[627], line_73[625], line_72[623], line_71[621], line_70[619], line_69[617], line_68[615], line_67[613], line_66[611], line_65[609], line_64[607], line_63[605], line_62[603], line_61[601], line_60[599], line_59[597], line_58[595], line_57[593], line_56[591], line_55[589], line_54[587], line_53[585], line_52[583], line_51[581], line_50[579], line_49[577], line_48[575], line_47[573], line_46[571], line_45[569], line_44[567], line_43[565], line_42[563], line_41[561], line_40[559], line_39[557], line_38[555], line_37[553], line_36[551], line_35[549], line_34[547], line_33[545], line_32[543], line_31[541], line_30[539], line_29[537], line_28[535], line_27[533], line_26[531], line_25[529], line_24[527], line_23[525], line_22[523], line_21[521], line_20[519], line_19[517], line_18[515], line_17[513], line_16[511], line_15[509], line_14[507], line_13[505], line_12[503], line_11[501], line_10[499], line_9[497], line_8[495], line_7[493], line_6[491], line_5[489], line_4[487], line_3[485], line_2[483], line_1[481] };
assign col_736 = {line_128[736], line_127[734], line_126[732], line_125[730], line_124[728], line_123[726], line_122[724], line_121[722], line_120[720], line_119[718], line_118[716], line_117[714], line_116[712], line_115[710], line_114[708], line_113[706], line_112[704], line_111[702], line_110[700], line_109[698], line_108[696], line_107[694], line_106[692], line_105[690], line_104[688], line_103[686], line_102[684], line_101[682], line_100[680], line_99[678], line_98[676], line_97[674], line_96[672], line_95[670], line_94[668], line_93[666], line_92[664], line_91[662], line_90[660], line_89[658], line_88[656], line_87[654], line_86[652], line_85[650], line_84[648], line_83[646], line_82[644], line_81[642], line_80[640], line_79[638], line_78[636], line_77[634], line_76[632], line_75[630], line_74[628], line_73[626], line_72[624], line_71[622], line_70[620], line_69[618], line_68[616], line_67[614], line_66[612], line_65[610], line_64[608], line_63[606], line_62[604], line_61[602], line_60[600], line_59[598], line_58[596], line_57[594], line_56[592], line_55[590], line_54[588], line_53[586], line_52[584], line_51[582], line_50[580], line_49[578], line_48[576], line_47[574], line_46[572], line_45[570], line_44[568], line_43[566], line_42[564], line_41[562], line_40[560], line_39[558], line_38[556], line_37[554], line_36[552], line_35[550], line_34[548], line_33[546], line_32[544], line_31[542], line_30[540], line_29[538], line_28[536], line_27[534], line_26[532], line_25[530], line_24[528], line_23[526], line_22[524], line_21[522], line_20[520], line_19[518], line_18[516], line_17[514], line_16[512], line_15[510], line_14[508], line_13[506], line_12[504], line_11[502], line_10[500], line_9[498], line_8[496], line_7[494], line_6[492], line_5[490], line_4[488], line_3[486], line_2[484], line_1[482] };
assign col_737 = {line_128[737], line_127[735], line_126[733], line_125[731], line_124[729], line_123[727], line_122[725], line_121[723], line_120[721], line_119[719], line_118[717], line_117[715], line_116[713], line_115[711], line_114[709], line_113[707], line_112[705], line_111[703], line_110[701], line_109[699], line_108[697], line_107[695], line_106[693], line_105[691], line_104[689], line_103[687], line_102[685], line_101[683], line_100[681], line_99[679], line_98[677], line_97[675], line_96[673], line_95[671], line_94[669], line_93[667], line_92[665], line_91[663], line_90[661], line_89[659], line_88[657], line_87[655], line_86[653], line_85[651], line_84[649], line_83[647], line_82[645], line_81[643], line_80[641], line_79[639], line_78[637], line_77[635], line_76[633], line_75[631], line_74[629], line_73[627], line_72[625], line_71[623], line_70[621], line_69[619], line_68[617], line_67[615], line_66[613], line_65[611], line_64[609], line_63[607], line_62[605], line_61[603], line_60[601], line_59[599], line_58[597], line_57[595], line_56[593], line_55[591], line_54[589], line_53[587], line_52[585], line_51[583], line_50[581], line_49[579], line_48[577], line_47[575], line_46[573], line_45[571], line_44[569], line_43[567], line_42[565], line_41[563], line_40[561], line_39[559], line_38[557], line_37[555], line_36[553], line_35[551], line_34[549], line_33[547], line_32[545], line_31[543], line_30[541], line_29[539], line_28[537], line_27[535], line_26[533], line_25[531], line_24[529], line_23[527], line_22[525], line_21[523], line_20[521], line_19[519], line_18[517], line_17[515], line_16[513], line_15[511], line_14[509], line_13[507], line_12[505], line_11[503], line_10[501], line_9[499], line_8[497], line_7[495], line_6[493], line_5[491], line_4[489], line_3[487], line_2[485], line_1[483] };
assign col_738 = {line_128[738], line_127[736], line_126[734], line_125[732], line_124[730], line_123[728], line_122[726], line_121[724], line_120[722], line_119[720], line_118[718], line_117[716], line_116[714], line_115[712], line_114[710], line_113[708], line_112[706], line_111[704], line_110[702], line_109[700], line_108[698], line_107[696], line_106[694], line_105[692], line_104[690], line_103[688], line_102[686], line_101[684], line_100[682], line_99[680], line_98[678], line_97[676], line_96[674], line_95[672], line_94[670], line_93[668], line_92[666], line_91[664], line_90[662], line_89[660], line_88[658], line_87[656], line_86[654], line_85[652], line_84[650], line_83[648], line_82[646], line_81[644], line_80[642], line_79[640], line_78[638], line_77[636], line_76[634], line_75[632], line_74[630], line_73[628], line_72[626], line_71[624], line_70[622], line_69[620], line_68[618], line_67[616], line_66[614], line_65[612], line_64[610], line_63[608], line_62[606], line_61[604], line_60[602], line_59[600], line_58[598], line_57[596], line_56[594], line_55[592], line_54[590], line_53[588], line_52[586], line_51[584], line_50[582], line_49[580], line_48[578], line_47[576], line_46[574], line_45[572], line_44[570], line_43[568], line_42[566], line_41[564], line_40[562], line_39[560], line_38[558], line_37[556], line_36[554], line_35[552], line_34[550], line_33[548], line_32[546], line_31[544], line_30[542], line_29[540], line_28[538], line_27[536], line_26[534], line_25[532], line_24[530], line_23[528], line_22[526], line_21[524], line_20[522], line_19[520], line_18[518], line_17[516], line_16[514], line_15[512], line_14[510], line_13[508], line_12[506], line_11[504], line_10[502], line_9[500], line_8[498], line_7[496], line_6[494], line_5[492], line_4[490], line_3[488], line_2[486], line_1[484] };
assign col_739 = {line_128[739], line_127[737], line_126[735], line_125[733], line_124[731], line_123[729], line_122[727], line_121[725], line_120[723], line_119[721], line_118[719], line_117[717], line_116[715], line_115[713], line_114[711], line_113[709], line_112[707], line_111[705], line_110[703], line_109[701], line_108[699], line_107[697], line_106[695], line_105[693], line_104[691], line_103[689], line_102[687], line_101[685], line_100[683], line_99[681], line_98[679], line_97[677], line_96[675], line_95[673], line_94[671], line_93[669], line_92[667], line_91[665], line_90[663], line_89[661], line_88[659], line_87[657], line_86[655], line_85[653], line_84[651], line_83[649], line_82[647], line_81[645], line_80[643], line_79[641], line_78[639], line_77[637], line_76[635], line_75[633], line_74[631], line_73[629], line_72[627], line_71[625], line_70[623], line_69[621], line_68[619], line_67[617], line_66[615], line_65[613], line_64[611], line_63[609], line_62[607], line_61[605], line_60[603], line_59[601], line_58[599], line_57[597], line_56[595], line_55[593], line_54[591], line_53[589], line_52[587], line_51[585], line_50[583], line_49[581], line_48[579], line_47[577], line_46[575], line_45[573], line_44[571], line_43[569], line_42[567], line_41[565], line_40[563], line_39[561], line_38[559], line_37[557], line_36[555], line_35[553], line_34[551], line_33[549], line_32[547], line_31[545], line_30[543], line_29[541], line_28[539], line_27[537], line_26[535], line_25[533], line_24[531], line_23[529], line_22[527], line_21[525], line_20[523], line_19[521], line_18[519], line_17[517], line_16[515], line_15[513], line_14[511], line_13[509], line_12[507], line_11[505], line_10[503], line_9[501], line_8[499], line_7[497], line_6[495], line_5[493], line_4[491], line_3[489], line_2[487], line_1[485] };
assign col_740 = {line_128[740], line_127[738], line_126[736], line_125[734], line_124[732], line_123[730], line_122[728], line_121[726], line_120[724], line_119[722], line_118[720], line_117[718], line_116[716], line_115[714], line_114[712], line_113[710], line_112[708], line_111[706], line_110[704], line_109[702], line_108[700], line_107[698], line_106[696], line_105[694], line_104[692], line_103[690], line_102[688], line_101[686], line_100[684], line_99[682], line_98[680], line_97[678], line_96[676], line_95[674], line_94[672], line_93[670], line_92[668], line_91[666], line_90[664], line_89[662], line_88[660], line_87[658], line_86[656], line_85[654], line_84[652], line_83[650], line_82[648], line_81[646], line_80[644], line_79[642], line_78[640], line_77[638], line_76[636], line_75[634], line_74[632], line_73[630], line_72[628], line_71[626], line_70[624], line_69[622], line_68[620], line_67[618], line_66[616], line_65[614], line_64[612], line_63[610], line_62[608], line_61[606], line_60[604], line_59[602], line_58[600], line_57[598], line_56[596], line_55[594], line_54[592], line_53[590], line_52[588], line_51[586], line_50[584], line_49[582], line_48[580], line_47[578], line_46[576], line_45[574], line_44[572], line_43[570], line_42[568], line_41[566], line_40[564], line_39[562], line_38[560], line_37[558], line_36[556], line_35[554], line_34[552], line_33[550], line_32[548], line_31[546], line_30[544], line_29[542], line_28[540], line_27[538], line_26[536], line_25[534], line_24[532], line_23[530], line_22[528], line_21[526], line_20[524], line_19[522], line_18[520], line_17[518], line_16[516], line_15[514], line_14[512], line_13[510], line_12[508], line_11[506], line_10[504], line_9[502], line_8[500], line_7[498], line_6[496], line_5[494], line_4[492], line_3[490], line_2[488], line_1[486] };
assign col_741 = {line_128[741], line_127[739], line_126[737], line_125[735], line_124[733], line_123[731], line_122[729], line_121[727], line_120[725], line_119[723], line_118[721], line_117[719], line_116[717], line_115[715], line_114[713], line_113[711], line_112[709], line_111[707], line_110[705], line_109[703], line_108[701], line_107[699], line_106[697], line_105[695], line_104[693], line_103[691], line_102[689], line_101[687], line_100[685], line_99[683], line_98[681], line_97[679], line_96[677], line_95[675], line_94[673], line_93[671], line_92[669], line_91[667], line_90[665], line_89[663], line_88[661], line_87[659], line_86[657], line_85[655], line_84[653], line_83[651], line_82[649], line_81[647], line_80[645], line_79[643], line_78[641], line_77[639], line_76[637], line_75[635], line_74[633], line_73[631], line_72[629], line_71[627], line_70[625], line_69[623], line_68[621], line_67[619], line_66[617], line_65[615], line_64[613], line_63[611], line_62[609], line_61[607], line_60[605], line_59[603], line_58[601], line_57[599], line_56[597], line_55[595], line_54[593], line_53[591], line_52[589], line_51[587], line_50[585], line_49[583], line_48[581], line_47[579], line_46[577], line_45[575], line_44[573], line_43[571], line_42[569], line_41[567], line_40[565], line_39[563], line_38[561], line_37[559], line_36[557], line_35[555], line_34[553], line_33[551], line_32[549], line_31[547], line_30[545], line_29[543], line_28[541], line_27[539], line_26[537], line_25[535], line_24[533], line_23[531], line_22[529], line_21[527], line_20[525], line_19[523], line_18[521], line_17[519], line_16[517], line_15[515], line_14[513], line_13[511], line_12[509], line_11[507], line_10[505], line_9[503], line_8[501], line_7[499], line_6[497], line_5[495], line_4[493], line_3[491], line_2[489], line_1[487] };
assign col_742 = {line_128[742], line_127[740], line_126[738], line_125[736], line_124[734], line_123[732], line_122[730], line_121[728], line_120[726], line_119[724], line_118[722], line_117[720], line_116[718], line_115[716], line_114[714], line_113[712], line_112[710], line_111[708], line_110[706], line_109[704], line_108[702], line_107[700], line_106[698], line_105[696], line_104[694], line_103[692], line_102[690], line_101[688], line_100[686], line_99[684], line_98[682], line_97[680], line_96[678], line_95[676], line_94[674], line_93[672], line_92[670], line_91[668], line_90[666], line_89[664], line_88[662], line_87[660], line_86[658], line_85[656], line_84[654], line_83[652], line_82[650], line_81[648], line_80[646], line_79[644], line_78[642], line_77[640], line_76[638], line_75[636], line_74[634], line_73[632], line_72[630], line_71[628], line_70[626], line_69[624], line_68[622], line_67[620], line_66[618], line_65[616], line_64[614], line_63[612], line_62[610], line_61[608], line_60[606], line_59[604], line_58[602], line_57[600], line_56[598], line_55[596], line_54[594], line_53[592], line_52[590], line_51[588], line_50[586], line_49[584], line_48[582], line_47[580], line_46[578], line_45[576], line_44[574], line_43[572], line_42[570], line_41[568], line_40[566], line_39[564], line_38[562], line_37[560], line_36[558], line_35[556], line_34[554], line_33[552], line_32[550], line_31[548], line_30[546], line_29[544], line_28[542], line_27[540], line_26[538], line_25[536], line_24[534], line_23[532], line_22[530], line_21[528], line_20[526], line_19[524], line_18[522], line_17[520], line_16[518], line_15[516], line_14[514], line_13[512], line_12[510], line_11[508], line_10[506], line_9[504], line_8[502], line_7[500], line_6[498], line_5[496], line_4[494], line_3[492], line_2[490], line_1[488] };
assign col_743 = {line_128[743], line_127[741], line_126[739], line_125[737], line_124[735], line_123[733], line_122[731], line_121[729], line_120[727], line_119[725], line_118[723], line_117[721], line_116[719], line_115[717], line_114[715], line_113[713], line_112[711], line_111[709], line_110[707], line_109[705], line_108[703], line_107[701], line_106[699], line_105[697], line_104[695], line_103[693], line_102[691], line_101[689], line_100[687], line_99[685], line_98[683], line_97[681], line_96[679], line_95[677], line_94[675], line_93[673], line_92[671], line_91[669], line_90[667], line_89[665], line_88[663], line_87[661], line_86[659], line_85[657], line_84[655], line_83[653], line_82[651], line_81[649], line_80[647], line_79[645], line_78[643], line_77[641], line_76[639], line_75[637], line_74[635], line_73[633], line_72[631], line_71[629], line_70[627], line_69[625], line_68[623], line_67[621], line_66[619], line_65[617], line_64[615], line_63[613], line_62[611], line_61[609], line_60[607], line_59[605], line_58[603], line_57[601], line_56[599], line_55[597], line_54[595], line_53[593], line_52[591], line_51[589], line_50[587], line_49[585], line_48[583], line_47[581], line_46[579], line_45[577], line_44[575], line_43[573], line_42[571], line_41[569], line_40[567], line_39[565], line_38[563], line_37[561], line_36[559], line_35[557], line_34[555], line_33[553], line_32[551], line_31[549], line_30[547], line_29[545], line_28[543], line_27[541], line_26[539], line_25[537], line_24[535], line_23[533], line_22[531], line_21[529], line_20[527], line_19[525], line_18[523], line_17[521], line_16[519], line_15[517], line_14[515], line_13[513], line_12[511], line_11[509], line_10[507], line_9[505], line_8[503], line_7[501], line_6[499], line_5[497], line_4[495], line_3[493], line_2[491], line_1[489] };
assign col_744 = {line_128[744], line_127[742], line_126[740], line_125[738], line_124[736], line_123[734], line_122[732], line_121[730], line_120[728], line_119[726], line_118[724], line_117[722], line_116[720], line_115[718], line_114[716], line_113[714], line_112[712], line_111[710], line_110[708], line_109[706], line_108[704], line_107[702], line_106[700], line_105[698], line_104[696], line_103[694], line_102[692], line_101[690], line_100[688], line_99[686], line_98[684], line_97[682], line_96[680], line_95[678], line_94[676], line_93[674], line_92[672], line_91[670], line_90[668], line_89[666], line_88[664], line_87[662], line_86[660], line_85[658], line_84[656], line_83[654], line_82[652], line_81[650], line_80[648], line_79[646], line_78[644], line_77[642], line_76[640], line_75[638], line_74[636], line_73[634], line_72[632], line_71[630], line_70[628], line_69[626], line_68[624], line_67[622], line_66[620], line_65[618], line_64[616], line_63[614], line_62[612], line_61[610], line_60[608], line_59[606], line_58[604], line_57[602], line_56[600], line_55[598], line_54[596], line_53[594], line_52[592], line_51[590], line_50[588], line_49[586], line_48[584], line_47[582], line_46[580], line_45[578], line_44[576], line_43[574], line_42[572], line_41[570], line_40[568], line_39[566], line_38[564], line_37[562], line_36[560], line_35[558], line_34[556], line_33[554], line_32[552], line_31[550], line_30[548], line_29[546], line_28[544], line_27[542], line_26[540], line_25[538], line_24[536], line_23[534], line_22[532], line_21[530], line_20[528], line_19[526], line_18[524], line_17[522], line_16[520], line_15[518], line_14[516], line_13[514], line_12[512], line_11[510], line_10[508], line_9[506], line_8[504], line_7[502], line_6[500], line_5[498], line_4[496], line_3[494], line_2[492], line_1[490] };
assign col_745 = {line_128[745], line_127[743], line_126[741], line_125[739], line_124[737], line_123[735], line_122[733], line_121[731], line_120[729], line_119[727], line_118[725], line_117[723], line_116[721], line_115[719], line_114[717], line_113[715], line_112[713], line_111[711], line_110[709], line_109[707], line_108[705], line_107[703], line_106[701], line_105[699], line_104[697], line_103[695], line_102[693], line_101[691], line_100[689], line_99[687], line_98[685], line_97[683], line_96[681], line_95[679], line_94[677], line_93[675], line_92[673], line_91[671], line_90[669], line_89[667], line_88[665], line_87[663], line_86[661], line_85[659], line_84[657], line_83[655], line_82[653], line_81[651], line_80[649], line_79[647], line_78[645], line_77[643], line_76[641], line_75[639], line_74[637], line_73[635], line_72[633], line_71[631], line_70[629], line_69[627], line_68[625], line_67[623], line_66[621], line_65[619], line_64[617], line_63[615], line_62[613], line_61[611], line_60[609], line_59[607], line_58[605], line_57[603], line_56[601], line_55[599], line_54[597], line_53[595], line_52[593], line_51[591], line_50[589], line_49[587], line_48[585], line_47[583], line_46[581], line_45[579], line_44[577], line_43[575], line_42[573], line_41[571], line_40[569], line_39[567], line_38[565], line_37[563], line_36[561], line_35[559], line_34[557], line_33[555], line_32[553], line_31[551], line_30[549], line_29[547], line_28[545], line_27[543], line_26[541], line_25[539], line_24[537], line_23[535], line_22[533], line_21[531], line_20[529], line_19[527], line_18[525], line_17[523], line_16[521], line_15[519], line_14[517], line_13[515], line_12[513], line_11[511], line_10[509], line_9[507], line_8[505], line_7[503], line_6[501], line_5[499], line_4[497], line_3[495], line_2[493], line_1[491] };
assign col_746 = {line_128[746], line_127[744], line_126[742], line_125[740], line_124[738], line_123[736], line_122[734], line_121[732], line_120[730], line_119[728], line_118[726], line_117[724], line_116[722], line_115[720], line_114[718], line_113[716], line_112[714], line_111[712], line_110[710], line_109[708], line_108[706], line_107[704], line_106[702], line_105[700], line_104[698], line_103[696], line_102[694], line_101[692], line_100[690], line_99[688], line_98[686], line_97[684], line_96[682], line_95[680], line_94[678], line_93[676], line_92[674], line_91[672], line_90[670], line_89[668], line_88[666], line_87[664], line_86[662], line_85[660], line_84[658], line_83[656], line_82[654], line_81[652], line_80[650], line_79[648], line_78[646], line_77[644], line_76[642], line_75[640], line_74[638], line_73[636], line_72[634], line_71[632], line_70[630], line_69[628], line_68[626], line_67[624], line_66[622], line_65[620], line_64[618], line_63[616], line_62[614], line_61[612], line_60[610], line_59[608], line_58[606], line_57[604], line_56[602], line_55[600], line_54[598], line_53[596], line_52[594], line_51[592], line_50[590], line_49[588], line_48[586], line_47[584], line_46[582], line_45[580], line_44[578], line_43[576], line_42[574], line_41[572], line_40[570], line_39[568], line_38[566], line_37[564], line_36[562], line_35[560], line_34[558], line_33[556], line_32[554], line_31[552], line_30[550], line_29[548], line_28[546], line_27[544], line_26[542], line_25[540], line_24[538], line_23[536], line_22[534], line_21[532], line_20[530], line_19[528], line_18[526], line_17[524], line_16[522], line_15[520], line_14[518], line_13[516], line_12[514], line_11[512], line_10[510], line_9[508], line_8[506], line_7[504], line_6[502], line_5[500], line_4[498], line_3[496], line_2[494], line_1[492] };
assign col_747 = {line_128[747], line_127[745], line_126[743], line_125[741], line_124[739], line_123[737], line_122[735], line_121[733], line_120[731], line_119[729], line_118[727], line_117[725], line_116[723], line_115[721], line_114[719], line_113[717], line_112[715], line_111[713], line_110[711], line_109[709], line_108[707], line_107[705], line_106[703], line_105[701], line_104[699], line_103[697], line_102[695], line_101[693], line_100[691], line_99[689], line_98[687], line_97[685], line_96[683], line_95[681], line_94[679], line_93[677], line_92[675], line_91[673], line_90[671], line_89[669], line_88[667], line_87[665], line_86[663], line_85[661], line_84[659], line_83[657], line_82[655], line_81[653], line_80[651], line_79[649], line_78[647], line_77[645], line_76[643], line_75[641], line_74[639], line_73[637], line_72[635], line_71[633], line_70[631], line_69[629], line_68[627], line_67[625], line_66[623], line_65[621], line_64[619], line_63[617], line_62[615], line_61[613], line_60[611], line_59[609], line_58[607], line_57[605], line_56[603], line_55[601], line_54[599], line_53[597], line_52[595], line_51[593], line_50[591], line_49[589], line_48[587], line_47[585], line_46[583], line_45[581], line_44[579], line_43[577], line_42[575], line_41[573], line_40[571], line_39[569], line_38[567], line_37[565], line_36[563], line_35[561], line_34[559], line_33[557], line_32[555], line_31[553], line_30[551], line_29[549], line_28[547], line_27[545], line_26[543], line_25[541], line_24[539], line_23[537], line_22[535], line_21[533], line_20[531], line_19[529], line_18[527], line_17[525], line_16[523], line_15[521], line_14[519], line_13[517], line_12[515], line_11[513], line_10[511], line_9[509], line_8[507], line_7[505], line_6[503], line_5[501], line_4[499], line_3[497], line_2[495], line_1[493] };
assign col_748 = {line_128[748], line_127[746], line_126[744], line_125[742], line_124[740], line_123[738], line_122[736], line_121[734], line_120[732], line_119[730], line_118[728], line_117[726], line_116[724], line_115[722], line_114[720], line_113[718], line_112[716], line_111[714], line_110[712], line_109[710], line_108[708], line_107[706], line_106[704], line_105[702], line_104[700], line_103[698], line_102[696], line_101[694], line_100[692], line_99[690], line_98[688], line_97[686], line_96[684], line_95[682], line_94[680], line_93[678], line_92[676], line_91[674], line_90[672], line_89[670], line_88[668], line_87[666], line_86[664], line_85[662], line_84[660], line_83[658], line_82[656], line_81[654], line_80[652], line_79[650], line_78[648], line_77[646], line_76[644], line_75[642], line_74[640], line_73[638], line_72[636], line_71[634], line_70[632], line_69[630], line_68[628], line_67[626], line_66[624], line_65[622], line_64[620], line_63[618], line_62[616], line_61[614], line_60[612], line_59[610], line_58[608], line_57[606], line_56[604], line_55[602], line_54[600], line_53[598], line_52[596], line_51[594], line_50[592], line_49[590], line_48[588], line_47[586], line_46[584], line_45[582], line_44[580], line_43[578], line_42[576], line_41[574], line_40[572], line_39[570], line_38[568], line_37[566], line_36[564], line_35[562], line_34[560], line_33[558], line_32[556], line_31[554], line_30[552], line_29[550], line_28[548], line_27[546], line_26[544], line_25[542], line_24[540], line_23[538], line_22[536], line_21[534], line_20[532], line_19[530], line_18[528], line_17[526], line_16[524], line_15[522], line_14[520], line_13[518], line_12[516], line_11[514], line_10[512], line_9[510], line_8[508], line_7[506], line_6[504], line_5[502], line_4[500], line_3[498], line_2[496], line_1[494] };
assign col_749 = {line_128[749], line_127[747], line_126[745], line_125[743], line_124[741], line_123[739], line_122[737], line_121[735], line_120[733], line_119[731], line_118[729], line_117[727], line_116[725], line_115[723], line_114[721], line_113[719], line_112[717], line_111[715], line_110[713], line_109[711], line_108[709], line_107[707], line_106[705], line_105[703], line_104[701], line_103[699], line_102[697], line_101[695], line_100[693], line_99[691], line_98[689], line_97[687], line_96[685], line_95[683], line_94[681], line_93[679], line_92[677], line_91[675], line_90[673], line_89[671], line_88[669], line_87[667], line_86[665], line_85[663], line_84[661], line_83[659], line_82[657], line_81[655], line_80[653], line_79[651], line_78[649], line_77[647], line_76[645], line_75[643], line_74[641], line_73[639], line_72[637], line_71[635], line_70[633], line_69[631], line_68[629], line_67[627], line_66[625], line_65[623], line_64[621], line_63[619], line_62[617], line_61[615], line_60[613], line_59[611], line_58[609], line_57[607], line_56[605], line_55[603], line_54[601], line_53[599], line_52[597], line_51[595], line_50[593], line_49[591], line_48[589], line_47[587], line_46[585], line_45[583], line_44[581], line_43[579], line_42[577], line_41[575], line_40[573], line_39[571], line_38[569], line_37[567], line_36[565], line_35[563], line_34[561], line_33[559], line_32[557], line_31[555], line_30[553], line_29[551], line_28[549], line_27[547], line_26[545], line_25[543], line_24[541], line_23[539], line_22[537], line_21[535], line_20[533], line_19[531], line_18[529], line_17[527], line_16[525], line_15[523], line_14[521], line_13[519], line_12[517], line_11[515], line_10[513], line_9[511], line_8[509], line_7[507], line_6[505], line_5[503], line_4[501], line_3[499], line_2[497], line_1[495] };
assign col_750 = {line_128[750], line_127[748], line_126[746], line_125[744], line_124[742], line_123[740], line_122[738], line_121[736], line_120[734], line_119[732], line_118[730], line_117[728], line_116[726], line_115[724], line_114[722], line_113[720], line_112[718], line_111[716], line_110[714], line_109[712], line_108[710], line_107[708], line_106[706], line_105[704], line_104[702], line_103[700], line_102[698], line_101[696], line_100[694], line_99[692], line_98[690], line_97[688], line_96[686], line_95[684], line_94[682], line_93[680], line_92[678], line_91[676], line_90[674], line_89[672], line_88[670], line_87[668], line_86[666], line_85[664], line_84[662], line_83[660], line_82[658], line_81[656], line_80[654], line_79[652], line_78[650], line_77[648], line_76[646], line_75[644], line_74[642], line_73[640], line_72[638], line_71[636], line_70[634], line_69[632], line_68[630], line_67[628], line_66[626], line_65[624], line_64[622], line_63[620], line_62[618], line_61[616], line_60[614], line_59[612], line_58[610], line_57[608], line_56[606], line_55[604], line_54[602], line_53[600], line_52[598], line_51[596], line_50[594], line_49[592], line_48[590], line_47[588], line_46[586], line_45[584], line_44[582], line_43[580], line_42[578], line_41[576], line_40[574], line_39[572], line_38[570], line_37[568], line_36[566], line_35[564], line_34[562], line_33[560], line_32[558], line_31[556], line_30[554], line_29[552], line_28[550], line_27[548], line_26[546], line_25[544], line_24[542], line_23[540], line_22[538], line_21[536], line_20[534], line_19[532], line_18[530], line_17[528], line_16[526], line_15[524], line_14[522], line_13[520], line_12[518], line_11[516], line_10[514], line_9[512], line_8[510], line_7[508], line_6[506], line_5[504], line_4[502], line_3[500], line_2[498], line_1[496] };
assign col_751 = {line_128[751], line_127[749], line_126[747], line_125[745], line_124[743], line_123[741], line_122[739], line_121[737], line_120[735], line_119[733], line_118[731], line_117[729], line_116[727], line_115[725], line_114[723], line_113[721], line_112[719], line_111[717], line_110[715], line_109[713], line_108[711], line_107[709], line_106[707], line_105[705], line_104[703], line_103[701], line_102[699], line_101[697], line_100[695], line_99[693], line_98[691], line_97[689], line_96[687], line_95[685], line_94[683], line_93[681], line_92[679], line_91[677], line_90[675], line_89[673], line_88[671], line_87[669], line_86[667], line_85[665], line_84[663], line_83[661], line_82[659], line_81[657], line_80[655], line_79[653], line_78[651], line_77[649], line_76[647], line_75[645], line_74[643], line_73[641], line_72[639], line_71[637], line_70[635], line_69[633], line_68[631], line_67[629], line_66[627], line_65[625], line_64[623], line_63[621], line_62[619], line_61[617], line_60[615], line_59[613], line_58[611], line_57[609], line_56[607], line_55[605], line_54[603], line_53[601], line_52[599], line_51[597], line_50[595], line_49[593], line_48[591], line_47[589], line_46[587], line_45[585], line_44[583], line_43[581], line_42[579], line_41[577], line_40[575], line_39[573], line_38[571], line_37[569], line_36[567], line_35[565], line_34[563], line_33[561], line_32[559], line_31[557], line_30[555], line_29[553], line_28[551], line_27[549], line_26[547], line_25[545], line_24[543], line_23[541], line_22[539], line_21[537], line_20[535], line_19[533], line_18[531], line_17[529], line_16[527], line_15[525], line_14[523], line_13[521], line_12[519], line_11[517], line_10[515], line_9[513], line_8[511], line_7[509], line_6[507], line_5[505], line_4[503], line_3[501], line_2[499], line_1[497] };
assign col_752 = {line_128[752], line_127[750], line_126[748], line_125[746], line_124[744], line_123[742], line_122[740], line_121[738], line_120[736], line_119[734], line_118[732], line_117[730], line_116[728], line_115[726], line_114[724], line_113[722], line_112[720], line_111[718], line_110[716], line_109[714], line_108[712], line_107[710], line_106[708], line_105[706], line_104[704], line_103[702], line_102[700], line_101[698], line_100[696], line_99[694], line_98[692], line_97[690], line_96[688], line_95[686], line_94[684], line_93[682], line_92[680], line_91[678], line_90[676], line_89[674], line_88[672], line_87[670], line_86[668], line_85[666], line_84[664], line_83[662], line_82[660], line_81[658], line_80[656], line_79[654], line_78[652], line_77[650], line_76[648], line_75[646], line_74[644], line_73[642], line_72[640], line_71[638], line_70[636], line_69[634], line_68[632], line_67[630], line_66[628], line_65[626], line_64[624], line_63[622], line_62[620], line_61[618], line_60[616], line_59[614], line_58[612], line_57[610], line_56[608], line_55[606], line_54[604], line_53[602], line_52[600], line_51[598], line_50[596], line_49[594], line_48[592], line_47[590], line_46[588], line_45[586], line_44[584], line_43[582], line_42[580], line_41[578], line_40[576], line_39[574], line_38[572], line_37[570], line_36[568], line_35[566], line_34[564], line_33[562], line_32[560], line_31[558], line_30[556], line_29[554], line_28[552], line_27[550], line_26[548], line_25[546], line_24[544], line_23[542], line_22[540], line_21[538], line_20[536], line_19[534], line_18[532], line_17[530], line_16[528], line_15[526], line_14[524], line_13[522], line_12[520], line_11[518], line_10[516], line_9[514], line_8[512], line_7[510], line_6[508], line_5[506], line_4[504], line_3[502], line_2[500], line_1[498] };
assign col_753 = {line_128[753], line_127[751], line_126[749], line_125[747], line_124[745], line_123[743], line_122[741], line_121[739], line_120[737], line_119[735], line_118[733], line_117[731], line_116[729], line_115[727], line_114[725], line_113[723], line_112[721], line_111[719], line_110[717], line_109[715], line_108[713], line_107[711], line_106[709], line_105[707], line_104[705], line_103[703], line_102[701], line_101[699], line_100[697], line_99[695], line_98[693], line_97[691], line_96[689], line_95[687], line_94[685], line_93[683], line_92[681], line_91[679], line_90[677], line_89[675], line_88[673], line_87[671], line_86[669], line_85[667], line_84[665], line_83[663], line_82[661], line_81[659], line_80[657], line_79[655], line_78[653], line_77[651], line_76[649], line_75[647], line_74[645], line_73[643], line_72[641], line_71[639], line_70[637], line_69[635], line_68[633], line_67[631], line_66[629], line_65[627], line_64[625], line_63[623], line_62[621], line_61[619], line_60[617], line_59[615], line_58[613], line_57[611], line_56[609], line_55[607], line_54[605], line_53[603], line_52[601], line_51[599], line_50[597], line_49[595], line_48[593], line_47[591], line_46[589], line_45[587], line_44[585], line_43[583], line_42[581], line_41[579], line_40[577], line_39[575], line_38[573], line_37[571], line_36[569], line_35[567], line_34[565], line_33[563], line_32[561], line_31[559], line_30[557], line_29[555], line_28[553], line_27[551], line_26[549], line_25[547], line_24[545], line_23[543], line_22[541], line_21[539], line_20[537], line_19[535], line_18[533], line_17[531], line_16[529], line_15[527], line_14[525], line_13[523], line_12[521], line_11[519], line_10[517], line_9[515], line_8[513], line_7[511], line_6[509], line_5[507], line_4[505], line_3[503], line_2[501], line_1[499] };
assign col_754 = {line_128[754], line_127[752], line_126[750], line_125[748], line_124[746], line_123[744], line_122[742], line_121[740], line_120[738], line_119[736], line_118[734], line_117[732], line_116[730], line_115[728], line_114[726], line_113[724], line_112[722], line_111[720], line_110[718], line_109[716], line_108[714], line_107[712], line_106[710], line_105[708], line_104[706], line_103[704], line_102[702], line_101[700], line_100[698], line_99[696], line_98[694], line_97[692], line_96[690], line_95[688], line_94[686], line_93[684], line_92[682], line_91[680], line_90[678], line_89[676], line_88[674], line_87[672], line_86[670], line_85[668], line_84[666], line_83[664], line_82[662], line_81[660], line_80[658], line_79[656], line_78[654], line_77[652], line_76[650], line_75[648], line_74[646], line_73[644], line_72[642], line_71[640], line_70[638], line_69[636], line_68[634], line_67[632], line_66[630], line_65[628], line_64[626], line_63[624], line_62[622], line_61[620], line_60[618], line_59[616], line_58[614], line_57[612], line_56[610], line_55[608], line_54[606], line_53[604], line_52[602], line_51[600], line_50[598], line_49[596], line_48[594], line_47[592], line_46[590], line_45[588], line_44[586], line_43[584], line_42[582], line_41[580], line_40[578], line_39[576], line_38[574], line_37[572], line_36[570], line_35[568], line_34[566], line_33[564], line_32[562], line_31[560], line_30[558], line_29[556], line_28[554], line_27[552], line_26[550], line_25[548], line_24[546], line_23[544], line_22[542], line_21[540], line_20[538], line_19[536], line_18[534], line_17[532], line_16[530], line_15[528], line_14[526], line_13[524], line_12[522], line_11[520], line_10[518], line_9[516], line_8[514], line_7[512], line_6[510], line_5[508], line_4[506], line_3[504], line_2[502], line_1[500] };
assign col_755 = {line_128[755], line_127[753], line_126[751], line_125[749], line_124[747], line_123[745], line_122[743], line_121[741], line_120[739], line_119[737], line_118[735], line_117[733], line_116[731], line_115[729], line_114[727], line_113[725], line_112[723], line_111[721], line_110[719], line_109[717], line_108[715], line_107[713], line_106[711], line_105[709], line_104[707], line_103[705], line_102[703], line_101[701], line_100[699], line_99[697], line_98[695], line_97[693], line_96[691], line_95[689], line_94[687], line_93[685], line_92[683], line_91[681], line_90[679], line_89[677], line_88[675], line_87[673], line_86[671], line_85[669], line_84[667], line_83[665], line_82[663], line_81[661], line_80[659], line_79[657], line_78[655], line_77[653], line_76[651], line_75[649], line_74[647], line_73[645], line_72[643], line_71[641], line_70[639], line_69[637], line_68[635], line_67[633], line_66[631], line_65[629], line_64[627], line_63[625], line_62[623], line_61[621], line_60[619], line_59[617], line_58[615], line_57[613], line_56[611], line_55[609], line_54[607], line_53[605], line_52[603], line_51[601], line_50[599], line_49[597], line_48[595], line_47[593], line_46[591], line_45[589], line_44[587], line_43[585], line_42[583], line_41[581], line_40[579], line_39[577], line_38[575], line_37[573], line_36[571], line_35[569], line_34[567], line_33[565], line_32[563], line_31[561], line_30[559], line_29[557], line_28[555], line_27[553], line_26[551], line_25[549], line_24[547], line_23[545], line_22[543], line_21[541], line_20[539], line_19[537], line_18[535], line_17[533], line_16[531], line_15[529], line_14[527], line_13[525], line_12[523], line_11[521], line_10[519], line_9[517], line_8[515], line_7[513], line_6[511], line_5[509], line_4[507], line_3[505], line_2[503], line_1[501] };
assign col_756 = {line_128[756], line_127[754], line_126[752], line_125[750], line_124[748], line_123[746], line_122[744], line_121[742], line_120[740], line_119[738], line_118[736], line_117[734], line_116[732], line_115[730], line_114[728], line_113[726], line_112[724], line_111[722], line_110[720], line_109[718], line_108[716], line_107[714], line_106[712], line_105[710], line_104[708], line_103[706], line_102[704], line_101[702], line_100[700], line_99[698], line_98[696], line_97[694], line_96[692], line_95[690], line_94[688], line_93[686], line_92[684], line_91[682], line_90[680], line_89[678], line_88[676], line_87[674], line_86[672], line_85[670], line_84[668], line_83[666], line_82[664], line_81[662], line_80[660], line_79[658], line_78[656], line_77[654], line_76[652], line_75[650], line_74[648], line_73[646], line_72[644], line_71[642], line_70[640], line_69[638], line_68[636], line_67[634], line_66[632], line_65[630], line_64[628], line_63[626], line_62[624], line_61[622], line_60[620], line_59[618], line_58[616], line_57[614], line_56[612], line_55[610], line_54[608], line_53[606], line_52[604], line_51[602], line_50[600], line_49[598], line_48[596], line_47[594], line_46[592], line_45[590], line_44[588], line_43[586], line_42[584], line_41[582], line_40[580], line_39[578], line_38[576], line_37[574], line_36[572], line_35[570], line_34[568], line_33[566], line_32[564], line_31[562], line_30[560], line_29[558], line_28[556], line_27[554], line_26[552], line_25[550], line_24[548], line_23[546], line_22[544], line_21[542], line_20[540], line_19[538], line_18[536], line_17[534], line_16[532], line_15[530], line_14[528], line_13[526], line_12[524], line_11[522], line_10[520], line_9[518], line_8[516], line_7[514], line_6[512], line_5[510], line_4[508], line_3[506], line_2[504], line_1[502] };
assign col_757 = {line_128[757], line_127[755], line_126[753], line_125[751], line_124[749], line_123[747], line_122[745], line_121[743], line_120[741], line_119[739], line_118[737], line_117[735], line_116[733], line_115[731], line_114[729], line_113[727], line_112[725], line_111[723], line_110[721], line_109[719], line_108[717], line_107[715], line_106[713], line_105[711], line_104[709], line_103[707], line_102[705], line_101[703], line_100[701], line_99[699], line_98[697], line_97[695], line_96[693], line_95[691], line_94[689], line_93[687], line_92[685], line_91[683], line_90[681], line_89[679], line_88[677], line_87[675], line_86[673], line_85[671], line_84[669], line_83[667], line_82[665], line_81[663], line_80[661], line_79[659], line_78[657], line_77[655], line_76[653], line_75[651], line_74[649], line_73[647], line_72[645], line_71[643], line_70[641], line_69[639], line_68[637], line_67[635], line_66[633], line_65[631], line_64[629], line_63[627], line_62[625], line_61[623], line_60[621], line_59[619], line_58[617], line_57[615], line_56[613], line_55[611], line_54[609], line_53[607], line_52[605], line_51[603], line_50[601], line_49[599], line_48[597], line_47[595], line_46[593], line_45[591], line_44[589], line_43[587], line_42[585], line_41[583], line_40[581], line_39[579], line_38[577], line_37[575], line_36[573], line_35[571], line_34[569], line_33[567], line_32[565], line_31[563], line_30[561], line_29[559], line_28[557], line_27[555], line_26[553], line_25[551], line_24[549], line_23[547], line_22[545], line_21[543], line_20[541], line_19[539], line_18[537], line_17[535], line_16[533], line_15[531], line_14[529], line_13[527], line_12[525], line_11[523], line_10[521], line_9[519], line_8[517], line_7[515], line_6[513], line_5[511], line_4[509], line_3[507], line_2[505], line_1[503] };
assign col_758 = {line_128[758], line_127[756], line_126[754], line_125[752], line_124[750], line_123[748], line_122[746], line_121[744], line_120[742], line_119[740], line_118[738], line_117[736], line_116[734], line_115[732], line_114[730], line_113[728], line_112[726], line_111[724], line_110[722], line_109[720], line_108[718], line_107[716], line_106[714], line_105[712], line_104[710], line_103[708], line_102[706], line_101[704], line_100[702], line_99[700], line_98[698], line_97[696], line_96[694], line_95[692], line_94[690], line_93[688], line_92[686], line_91[684], line_90[682], line_89[680], line_88[678], line_87[676], line_86[674], line_85[672], line_84[670], line_83[668], line_82[666], line_81[664], line_80[662], line_79[660], line_78[658], line_77[656], line_76[654], line_75[652], line_74[650], line_73[648], line_72[646], line_71[644], line_70[642], line_69[640], line_68[638], line_67[636], line_66[634], line_65[632], line_64[630], line_63[628], line_62[626], line_61[624], line_60[622], line_59[620], line_58[618], line_57[616], line_56[614], line_55[612], line_54[610], line_53[608], line_52[606], line_51[604], line_50[602], line_49[600], line_48[598], line_47[596], line_46[594], line_45[592], line_44[590], line_43[588], line_42[586], line_41[584], line_40[582], line_39[580], line_38[578], line_37[576], line_36[574], line_35[572], line_34[570], line_33[568], line_32[566], line_31[564], line_30[562], line_29[560], line_28[558], line_27[556], line_26[554], line_25[552], line_24[550], line_23[548], line_22[546], line_21[544], line_20[542], line_19[540], line_18[538], line_17[536], line_16[534], line_15[532], line_14[530], line_13[528], line_12[526], line_11[524], line_10[522], line_9[520], line_8[518], line_7[516], line_6[514], line_5[512], line_4[510], line_3[508], line_2[506], line_1[504] };
assign col_759 = {line_128[759], line_127[757], line_126[755], line_125[753], line_124[751], line_123[749], line_122[747], line_121[745], line_120[743], line_119[741], line_118[739], line_117[737], line_116[735], line_115[733], line_114[731], line_113[729], line_112[727], line_111[725], line_110[723], line_109[721], line_108[719], line_107[717], line_106[715], line_105[713], line_104[711], line_103[709], line_102[707], line_101[705], line_100[703], line_99[701], line_98[699], line_97[697], line_96[695], line_95[693], line_94[691], line_93[689], line_92[687], line_91[685], line_90[683], line_89[681], line_88[679], line_87[677], line_86[675], line_85[673], line_84[671], line_83[669], line_82[667], line_81[665], line_80[663], line_79[661], line_78[659], line_77[657], line_76[655], line_75[653], line_74[651], line_73[649], line_72[647], line_71[645], line_70[643], line_69[641], line_68[639], line_67[637], line_66[635], line_65[633], line_64[631], line_63[629], line_62[627], line_61[625], line_60[623], line_59[621], line_58[619], line_57[617], line_56[615], line_55[613], line_54[611], line_53[609], line_52[607], line_51[605], line_50[603], line_49[601], line_48[599], line_47[597], line_46[595], line_45[593], line_44[591], line_43[589], line_42[587], line_41[585], line_40[583], line_39[581], line_38[579], line_37[577], line_36[575], line_35[573], line_34[571], line_33[569], line_32[567], line_31[565], line_30[563], line_29[561], line_28[559], line_27[557], line_26[555], line_25[553], line_24[551], line_23[549], line_22[547], line_21[545], line_20[543], line_19[541], line_18[539], line_17[537], line_16[535], line_15[533], line_14[531], line_13[529], line_12[527], line_11[525], line_10[523], line_9[521], line_8[519], line_7[517], line_6[515], line_5[513], line_4[511], line_3[509], line_2[507], line_1[505] };
assign col_760 = {line_128[760], line_127[758], line_126[756], line_125[754], line_124[752], line_123[750], line_122[748], line_121[746], line_120[744], line_119[742], line_118[740], line_117[738], line_116[736], line_115[734], line_114[732], line_113[730], line_112[728], line_111[726], line_110[724], line_109[722], line_108[720], line_107[718], line_106[716], line_105[714], line_104[712], line_103[710], line_102[708], line_101[706], line_100[704], line_99[702], line_98[700], line_97[698], line_96[696], line_95[694], line_94[692], line_93[690], line_92[688], line_91[686], line_90[684], line_89[682], line_88[680], line_87[678], line_86[676], line_85[674], line_84[672], line_83[670], line_82[668], line_81[666], line_80[664], line_79[662], line_78[660], line_77[658], line_76[656], line_75[654], line_74[652], line_73[650], line_72[648], line_71[646], line_70[644], line_69[642], line_68[640], line_67[638], line_66[636], line_65[634], line_64[632], line_63[630], line_62[628], line_61[626], line_60[624], line_59[622], line_58[620], line_57[618], line_56[616], line_55[614], line_54[612], line_53[610], line_52[608], line_51[606], line_50[604], line_49[602], line_48[600], line_47[598], line_46[596], line_45[594], line_44[592], line_43[590], line_42[588], line_41[586], line_40[584], line_39[582], line_38[580], line_37[578], line_36[576], line_35[574], line_34[572], line_33[570], line_32[568], line_31[566], line_30[564], line_29[562], line_28[560], line_27[558], line_26[556], line_25[554], line_24[552], line_23[550], line_22[548], line_21[546], line_20[544], line_19[542], line_18[540], line_17[538], line_16[536], line_15[534], line_14[532], line_13[530], line_12[528], line_11[526], line_10[524], line_9[522], line_8[520], line_7[518], line_6[516], line_5[514], line_4[512], line_3[510], line_2[508], line_1[506] };
assign col_761 = {line_128[761], line_127[759], line_126[757], line_125[755], line_124[753], line_123[751], line_122[749], line_121[747], line_120[745], line_119[743], line_118[741], line_117[739], line_116[737], line_115[735], line_114[733], line_113[731], line_112[729], line_111[727], line_110[725], line_109[723], line_108[721], line_107[719], line_106[717], line_105[715], line_104[713], line_103[711], line_102[709], line_101[707], line_100[705], line_99[703], line_98[701], line_97[699], line_96[697], line_95[695], line_94[693], line_93[691], line_92[689], line_91[687], line_90[685], line_89[683], line_88[681], line_87[679], line_86[677], line_85[675], line_84[673], line_83[671], line_82[669], line_81[667], line_80[665], line_79[663], line_78[661], line_77[659], line_76[657], line_75[655], line_74[653], line_73[651], line_72[649], line_71[647], line_70[645], line_69[643], line_68[641], line_67[639], line_66[637], line_65[635], line_64[633], line_63[631], line_62[629], line_61[627], line_60[625], line_59[623], line_58[621], line_57[619], line_56[617], line_55[615], line_54[613], line_53[611], line_52[609], line_51[607], line_50[605], line_49[603], line_48[601], line_47[599], line_46[597], line_45[595], line_44[593], line_43[591], line_42[589], line_41[587], line_40[585], line_39[583], line_38[581], line_37[579], line_36[577], line_35[575], line_34[573], line_33[571], line_32[569], line_31[567], line_30[565], line_29[563], line_28[561], line_27[559], line_26[557], line_25[555], line_24[553], line_23[551], line_22[549], line_21[547], line_20[545], line_19[543], line_18[541], line_17[539], line_16[537], line_15[535], line_14[533], line_13[531], line_12[529], line_11[527], line_10[525], line_9[523], line_8[521], line_7[519], line_6[517], line_5[515], line_4[513], line_3[511], line_2[509], line_1[507] };
assign col_762 = {line_128[762], line_127[760], line_126[758], line_125[756], line_124[754], line_123[752], line_122[750], line_121[748], line_120[746], line_119[744], line_118[742], line_117[740], line_116[738], line_115[736], line_114[734], line_113[732], line_112[730], line_111[728], line_110[726], line_109[724], line_108[722], line_107[720], line_106[718], line_105[716], line_104[714], line_103[712], line_102[710], line_101[708], line_100[706], line_99[704], line_98[702], line_97[700], line_96[698], line_95[696], line_94[694], line_93[692], line_92[690], line_91[688], line_90[686], line_89[684], line_88[682], line_87[680], line_86[678], line_85[676], line_84[674], line_83[672], line_82[670], line_81[668], line_80[666], line_79[664], line_78[662], line_77[660], line_76[658], line_75[656], line_74[654], line_73[652], line_72[650], line_71[648], line_70[646], line_69[644], line_68[642], line_67[640], line_66[638], line_65[636], line_64[634], line_63[632], line_62[630], line_61[628], line_60[626], line_59[624], line_58[622], line_57[620], line_56[618], line_55[616], line_54[614], line_53[612], line_52[610], line_51[608], line_50[606], line_49[604], line_48[602], line_47[600], line_46[598], line_45[596], line_44[594], line_43[592], line_42[590], line_41[588], line_40[586], line_39[584], line_38[582], line_37[580], line_36[578], line_35[576], line_34[574], line_33[572], line_32[570], line_31[568], line_30[566], line_29[564], line_28[562], line_27[560], line_26[558], line_25[556], line_24[554], line_23[552], line_22[550], line_21[548], line_20[546], line_19[544], line_18[542], line_17[540], line_16[538], line_15[536], line_14[534], line_13[532], line_12[530], line_11[528], line_10[526], line_9[524], line_8[522], line_7[520], line_6[518], line_5[516], line_4[514], line_3[512], line_2[510], line_1[508] };
assign col_763 = {line_128[763], line_127[761], line_126[759], line_125[757], line_124[755], line_123[753], line_122[751], line_121[749], line_120[747], line_119[745], line_118[743], line_117[741], line_116[739], line_115[737], line_114[735], line_113[733], line_112[731], line_111[729], line_110[727], line_109[725], line_108[723], line_107[721], line_106[719], line_105[717], line_104[715], line_103[713], line_102[711], line_101[709], line_100[707], line_99[705], line_98[703], line_97[701], line_96[699], line_95[697], line_94[695], line_93[693], line_92[691], line_91[689], line_90[687], line_89[685], line_88[683], line_87[681], line_86[679], line_85[677], line_84[675], line_83[673], line_82[671], line_81[669], line_80[667], line_79[665], line_78[663], line_77[661], line_76[659], line_75[657], line_74[655], line_73[653], line_72[651], line_71[649], line_70[647], line_69[645], line_68[643], line_67[641], line_66[639], line_65[637], line_64[635], line_63[633], line_62[631], line_61[629], line_60[627], line_59[625], line_58[623], line_57[621], line_56[619], line_55[617], line_54[615], line_53[613], line_52[611], line_51[609], line_50[607], line_49[605], line_48[603], line_47[601], line_46[599], line_45[597], line_44[595], line_43[593], line_42[591], line_41[589], line_40[587], line_39[585], line_38[583], line_37[581], line_36[579], line_35[577], line_34[575], line_33[573], line_32[571], line_31[569], line_30[567], line_29[565], line_28[563], line_27[561], line_26[559], line_25[557], line_24[555], line_23[553], line_22[551], line_21[549], line_20[547], line_19[545], line_18[543], line_17[541], line_16[539], line_15[537], line_14[535], line_13[533], line_12[531], line_11[529], line_10[527], line_9[525], line_8[523], line_7[521], line_6[519], line_5[517], line_4[515], line_3[513], line_2[511], line_1[509] };
assign col_764 = {line_128[764], line_127[762], line_126[760], line_125[758], line_124[756], line_123[754], line_122[752], line_121[750], line_120[748], line_119[746], line_118[744], line_117[742], line_116[740], line_115[738], line_114[736], line_113[734], line_112[732], line_111[730], line_110[728], line_109[726], line_108[724], line_107[722], line_106[720], line_105[718], line_104[716], line_103[714], line_102[712], line_101[710], line_100[708], line_99[706], line_98[704], line_97[702], line_96[700], line_95[698], line_94[696], line_93[694], line_92[692], line_91[690], line_90[688], line_89[686], line_88[684], line_87[682], line_86[680], line_85[678], line_84[676], line_83[674], line_82[672], line_81[670], line_80[668], line_79[666], line_78[664], line_77[662], line_76[660], line_75[658], line_74[656], line_73[654], line_72[652], line_71[650], line_70[648], line_69[646], line_68[644], line_67[642], line_66[640], line_65[638], line_64[636], line_63[634], line_62[632], line_61[630], line_60[628], line_59[626], line_58[624], line_57[622], line_56[620], line_55[618], line_54[616], line_53[614], line_52[612], line_51[610], line_50[608], line_49[606], line_48[604], line_47[602], line_46[600], line_45[598], line_44[596], line_43[594], line_42[592], line_41[590], line_40[588], line_39[586], line_38[584], line_37[582], line_36[580], line_35[578], line_34[576], line_33[574], line_32[572], line_31[570], line_30[568], line_29[566], line_28[564], line_27[562], line_26[560], line_25[558], line_24[556], line_23[554], line_22[552], line_21[550], line_20[548], line_19[546], line_18[544], line_17[542], line_16[540], line_15[538], line_14[536], line_13[534], line_12[532], line_11[530], line_10[528], line_9[526], line_8[524], line_7[522], line_6[520], line_5[518], line_4[516], line_3[514], line_2[512], line_1[510] };
assign col_765 = {line_128[765], line_127[763], line_126[761], line_125[759], line_124[757], line_123[755], line_122[753], line_121[751], line_120[749], line_119[747], line_118[745], line_117[743], line_116[741], line_115[739], line_114[737], line_113[735], line_112[733], line_111[731], line_110[729], line_109[727], line_108[725], line_107[723], line_106[721], line_105[719], line_104[717], line_103[715], line_102[713], line_101[711], line_100[709], line_99[707], line_98[705], line_97[703], line_96[701], line_95[699], line_94[697], line_93[695], line_92[693], line_91[691], line_90[689], line_89[687], line_88[685], line_87[683], line_86[681], line_85[679], line_84[677], line_83[675], line_82[673], line_81[671], line_80[669], line_79[667], line_78[665], line_77[663], line_76[661], line_75[659], line_74[657], line_73[655], line_72[653], line_71[651], line_70[649], line_69[647], line_68[645], line_67[643], line_66[641], line_65[639], line_64[637], line_63[635], line_62[633], line_61[631], line_60[629], line_59[627], line_58[625], line_57[623], line_56[621], line_55[619], line_54[617], line_53[615], line_52[613], line_51[611], line_50[609], line_49[607], line_48[605], line_47[603], line_46[601], line_45[599], line_44[597], line_43[595], line_42[593], line_41[591], line_40[589], line_39[587], line_38[585], line_37[583], line_36[581], line_35[579], line_34[577], line_33[575], line_32[573], line_31[571], line_30[569], line_29[567], line_28[565], line_27[563], line_26[561], line_25[559], line_24[557], line_23[555], line_22[553], line_21[551], line_20[549], line_19[547], line_18[545], line_17[543], line_16[541], line_15[539], line_14[537], line_13[535], line_12[533], line_11[531], line_10[529], line_9[527], line_8[525], line_7[523], line_6[521], line_5[519], line_4[517], line_3[515], line_2[513], line_1[511] };
assign col_766 = {line_128[766], line_127[764], line_126[762], line_125[760], line_124[758], line_123[756], line_122[754], line_121[752], line_120[750], line_119[748], line_118[746], line_117[744], line_116[742], line_115[740], line_114[738], line_113[736], line_112[734], line_111[732], line_110[730], line_109[728], line_108[726], line_107[724], line_106[722], line_105[720], line_104[718], line_103[716], line_102[714], line_101[712], line_100[710], line_99[708], line_98[706], line_97[704], line_96[702], line_95[700], line_94[698], line_93[696], line_92[694], line_91[692], line_90[690], line_89[688], line_88[686], line_87[684], line_86[682], line_85[680], line_84[678], line_83[676], line_82[674], line_81[672], line_80[670], line_79[668], line_78[666], line_77[664], line_76[662], line_75[660], line_74[658], line_73[656], line_72[654], line_71[652], line_70[650], line_69[648], line_68[646], line_67[644], line_66[642], line_65[640], line_64[638], line_63[636], line_62[634], line_61[632], line_60[630], line_59[628], line_58[626], line_57[624], line_56[622], line_55[620], line_54[618], line_53[616], line_52[614], line_51[612], line_50[610], line_49[608], line_48[606], line_47[604], line_46[602], line_45[600], line_44[598], line_43[596], line_42[594], line_41[592], line_40[590], line_39[588], line_38[586], line_37[584], line_36[582], line_35[580], line_34[578], line_33[576], line_32[574], line_31[572], line_30[570], line_29[568], line_28[566], line_27[564], line_26[562], line_25[560], line_24[558], line_23[556], line_22[554], line_21[552], line_20[550], line_19[548], line_18[546], line_17[544], line_16[542], line_15[540], line_14[538], line_13[536], line_12[534], line_11[532], line_10[530], line_9[528], line_8[526], line_7[524], line_6[522], line_5[520], line_4[518], line_3[516], line_2[514], line_1[512] };
assign col_767 = {line_128[767], line_127[765], line_126[763], line_125[761], line_124[759], line_123[757], line_122[755], line_121[753], line_120[751], line_119[749], line_118[747], line_117[745], line_116[743], line_115[741], line_114[739], line_113[737], line_112[735], line_111[733], line_110[731], line_109[729], line_108[727], line_107[725], line_106[723], line_105[721], line_104[719], line_103[717], line_102[715], line_101[713], line_100[711], line_99[709], line_98[707], line_97[705], line_96[703], line_95[701], line_94[699], line_93[697], line_92[695], line_91[693], line_90[691], line_89[689], line_88[687], line_87[685], line_86[683], line_85[681], line_84[679], line_83[677], line_82[675], line_81[673], line_80[671], line_79[669], line_78[667], line_77[665], line_76[663], line_75[661], line_74[659], line_73[657], line_72[655], line_71[653], line_70[651], line_69[649], line_68[647], line_67[645], line_66[643], line_65[641], line_64[639], line_63[637], line_62[635], line_61[633], line_60[631], line_59[629], line_58[627], line_57[625], line_56[623], line_55[621], line_54[619], line_53[617], line_52[615], line_51[613], line_50[611], line_49[609], line_48[607], line_47[605], line_46[603], line_45[601], line_44[599], line_43[597], line_42[595], line_41[593], line_40[591], line_39[589], line_38[587], line_37[585], line_36[583], line_35[581], line_34[579], line_33[577], line_32[575], line_31[573], line_30[571], line_29[569], line_28[567], line_27[565], line_26[563], line_25[561], line_24[559], line_23[557], line_22[555], line_21[553], line_20[551], line_19[549], line_18[547], line_17[545], line_16[543], line_15[541], line_14[539], line_13[537], line_12[535], line_11[533], line_10[531], line_9[529], line_8[527], line_7[525], line_6[523], line_5[521], line_4[519], line_3[517], line_2[515], line_1[513] };
assign col_768 = {line_128[768], line_127[766], line_126[764], line_125[762], line_124[760], line_123[758], line_122[756], line_121[754], line_120[752], line_119[750], line_118[748], line_117[746], line_116[744], line_115[742], line_114[740], line_113[738], line_112[736], line_111[734], line_110[732], line_109[730], line_108[728], line_107[726], line_106[724], line_105[722], line_104[720], line_103[718], line_102[716], line_101[714], line_100[712], line_99[710], line_98[708], line_97[706], line_96[704], line_95[702], line_94[700], line_93[698], line_92[696], line_91[694], line_90[692], line_89[690], line_88[688], line_87[686], line_86[684], line_85[682], line_84[680], line_83[678], line_82[676], line_81[674], line_80[672], line_79[670], line_78[668], line_77[666], line_76[664], line_75[662], line_74[660], line_73[658], line_72[656], line_71[654], line_70[652], line_69[650], line_68[648], line_67[646], line_66[644], line_65[642], line_64[640], line_63[638], line_62[636], line_61[634], line_60[632], line_59[630], line_58[628], line_57[626], line_56[624], line_55[622], line_54[620], line_53[618], line_52[616], line_51[614], line_50[612], line_49[610], line_48[608], line_47[606], line_46[604], line_45[602], line_44[600], line_43[598], line_42[596], line_41[594], line_40[592], line_39[590], line_38[588], line_37[586], line_36[584], line_35[582], line_34[580], line_33[578], line_32[576], line_31[574], line_30[572], line_29[570], line_28[568], line_27[566], line_26[564], line_25[562], line_24[560], line_23[558], line_22[556], line_21[554], line_20[552], line_19[550], line_18[548], line_17[546], line_16[544], line_15[542], line_14[540], line_13[538], line_12[536], line_11[534], line_10[532], line_9[530], line_8[528], line_7[526], line_6[524], line_5[522], line_4[520], line_3[518], line_2[516], line_1[514] };
assign col_769 = {line_128[769], line_127[767], line_126[765], line_125[763], line_124[761], line_123[759], line_122[757], line_121[755], line_120[753], line_119[751], line_118[749], line_117[747], line_116[745], line_115[743], line_114[741], line_113[739], line_112[737], line_111[735], line_110[733], line_109[731], line_108[729], line_107[727], line_106[725], line_105[723], line_104[721], line_103[719], line_102[717], line_101[715], line_100[713], line_99[711], line_98[709], line_97[707], line_96[705], line_95[703], line_94[701], line_93[699], line_92[697], line_91[695], line_90[693], line_89[691], line_88[689], line_87[687], line_86[685], line_85[683], line_84[681], line_83[679], line_82[677], line_81[675], line_80[673], line_79[671], line_78[669], line_77[667], line_76[665], line_75[663], line_74[661], line_73[659], line_72[657], line_71[655], line_70[653], line_69[651], line_68[649], line_67[647], line_66[645], line_65[643], line_64[641], line_63[639], line_62[637], line_61[635], line_60[633], line_59[631], line_58[629], line_57[627], line_56[625], line_55[623], line_54[621], line_53[619], line_52[617], line_51[615], line_50[613], line_49[611], line_48[609], line_47[607], line_46[605], line_45[603], line_44[601], line_43[599], line_42[597], line_41[595], line_40[593], line_39[591], line_38[589], line_37[587], line_36[585], line_35[583], line_34[581], line_33[579], line_32[577], line_31[575], line_30[573], line_29[571], line_28[569], line_27[567], line_26[565], line_25[563], line_24[561], line_23[559], line_22[557], line_21[555], line_20[553], line_19[551], line_18[549], line_17[547], line_16[545], line_15[543], line_14[541], line_13[539], line_12[537], line_11[535], line_10[533], line_9[531], line_8[529], line_7[527], line_6[525], line_5[523], line_4[521], line_3[519], line_2[517], line_1[515] };
assign col_770 = {line_128[770], line_127[768], line_126[766], line_125[764], line_124[762], line_123[760], line_122[758], line_121[756], line_120[754], line_119[752], line_118[750], line_117[748], line_116[746], line_115[744], line_114[742], line_113[740], line_112[738], line_111[736], line_110[734], line_109[732], line_108[730], line_107[728], line_106[726], line_105[724], line_104[722], line_103[720], line_102[718], line_101[716], line_100[714], line_99[712], line_98[710], line_97[708], line_96[706], line_95[704], line_94[702], line_93[700], line_92[698], line_91[696], line_90[694], line_89[692], line_88[690], line_87[688], line_86[686], line_85[684], line_84[682], line_83[680], line_82[678], line_81[676], line_80[674], line_79[672], line_78[670], line_77[668], line_76[666], line_75[664], line_74[662], line_73[660], line_72[658], line_71[656], line_70[654], line_69[652], line_68[650], line_67[648], line_66[646], line_65[644], line_64[642], line_63[640], line_62[638], line_61[636], line_60[634], line_59[632], line_58[630], line_57[628], line_56[626], line_55[624], line_54[622], line_53[620], line_52[618], line_51[616], line_50[614], line_49[612], line_48[610], line_47[608], line_46[606], line_45[604], line_44[602], line_43[600], line_42[598], line_41[596], line_40[594], line_39[592], line_38[590], line_37[588], line_36[586], line_35[584], line_34[582], line_33[580], line_32[578], line_31[576], line_30[574], line_29[572], line_28[570], line_27[568], line_26[566], line_25[564], line_24[562], line_23[560], line_22[558], line_21[556], line_20[554], line_19[552], line_18[550], line_17[548], line_16[546], line_15[544], line_14[542], line_13[540], line_12[538], line_11[536], line_10[534], line_9[532], line_8[530], line_7[528], line_6[526], line_5[524], line_4[522], line_3[520], line_2[518], line_1[516] };
assign col_771 = {line_128[771], line_127[769], line_126[767], line_125[765], line_124[763], line_123[761], line_122[759], line_121[757], line_120[755], line_119[753], line_118[751], line_117[749], line_116[747], line_115[745], line_114[743], line_113[741], line_112[739], line_111[737], line_110[735], line_109[733], line_108[731], line_107[729], line_106[727], line_105[725], line_104[723], line_103[721], line_102[719], line_101[717], line_100[715], line_99[713], line_98[711], line_97[709], line_96[707], line_95[705], line_94[703], line_93[701], line_92[699], line_91[697], line_90[695], line_89[693], line_88[691], line_87[689], line_86[687], line_85[685], line_84[683], line_83[681], line_82[679], line_81[677], line_80[675], line_79[673], line_78[671], line_77[669], line_76[667], line_75[665], line_74[663], line_73[661], line_72[659], line_71[657], line_70[655], line_69[653], line_68[651], line_67[649], line_66[647], line_65[645], line_64[643], line_63[641], line_62[639], line_61[637], line_60[635], line_59[633], line_58[631], line_57[629], line_56[627], line_55[625], line_54[623], line_53[621], line_52[619], line_51[617], line_50[615], line_49[613], line_48[611], line_47[609], line_46[607], line_45[605], line_44[603], line_43[601], line_42[599], line_41[597], line_40[595], line_39[593], line_38[591], line_37[589], line_36[587], line_35[585], line_34[583], line_33[581], line_32[579], line_31[577], line_30[575], line_29[573], line_28[571], line_27[569], line_26[567], line_25[565], line_24[563], line_23[561], line_22[559], line_21[557], line_20[555], line_19[553], line_18[551], line_17[549], line_16[547], line_15[545], line_14[543], line_13[541], line_12[539], line_11[537], line_10[535], line_9[533], line_8[531], line_7[529], line_6[527], line_5[525], line_4[523], line_3[521], line_2[519], line_1[517] };
assign col_772 = {line_128[772], line_127[770], line_126[768], line_125[766], line_124[764], line_123[762], line_122[760], line_121[758], line_120[756], line_119[754], line_118[752], line_117[750], line_116[748], line_115[746], line_114[744], line_113[742], line_112[740], line_111[738], line_110[736], line_109[734], line_108[732], line_107[730], line_106[728], line_105[726], line_104[724], line_103[722], line_102[720], line_101[718], line_100[716], line_99[714], line_98[712], line_97[710], line_96[708], line_95[706], line_94[704], line_93[702], line_92[700], line_91[698], line_90[696], line_89[694], line_88[692], line_87[690], line_86[688], line_85[686], line_84[684], line_83[682], line_82[680], line_81[678], line_80[676], line_79[674], line_78[672], line_77[670], line_76[668], line_75[666], line_74[664], line_73[662], line_72[660], line_71[658], line_70[656], line_69[654], line_68[652], line_67[650], line_66[648], line_65[646], line_64[644], line_63[642], line_62[640], line_61[638], line_60[636], line_59[634], line_58[632], line_57[630], line_56[628], line_55[626], line_54[624], line_53[622], line_52[620], line_51[618], line_50[616], line_49[614], line_48[612], line_47[610], line_46[608], line_45[606], line_44[604], line_43[602], line_42[600], line_41[598], line_40[596], line_39[594], line_38[592], line_37[590], line_36[588], line_35[586], line_34[584], line_33[582], line_32[580], line_31[578], line_30[576], line_29[574], line_28[572], line_27[570], line_26[568], line_25[566], line_24[564], line_23[562], line_22[560], line_21[558], line_20[556], line_19[554], line_18[552], line_17[550], line_16[548], line_15[546], line_14[544], line_13[542], line_12[540], line_11[538], line_10[536], line_9[534], line_8[532], line_7[530], line_6[528], line_5[526], line_4[524], line_3[522], line_2[520], line_1[518] };
assign col_773 = {line_128[773], line_127[771], line_126[769], line_125[767], line_124[765], line_123[763], line_122[761], line_121[759], line_120[757], line_119[755], line_118[753], line_117[751], line_116[749], line_115[747], line_114[745], line_113[743], line_112[741], line_111[739], line_110[737], line_109[735], line_108[733], line_107[731], line_106[729], line_105[727], line_104[725], line_103[723], line_102[721], line_101[719], line_100[717], line_99[715], line_98[713], line_97[711], line_96[709], line_95[707], line_94[705], line_93[703], line_92[701], line_91[699], line_90[697], line_89[695], line_88[693], line_87[691], line_86[689], line_85[687], line_84[685], line_83[683], line_82[681], line_81[679], line_80[677], line_79[675], line_78[673], line_77[671], line_76[669], line_75[667], line_74[665], line_73[663], line_72[661], line_71[659], line_70[657], line_69[655], line_68[653], line_67[651], line_66[649], line_65[647], line_64[645], line_63[643], line_62[641], line_61[639], line_60[637], line_59[635], line_58[633], line_57[631], line_56[629], line_55[627], line_54[625], line_53[623], line_52[621], line_51[619], line_50[617], line_49[615], line_48[613], line_47[611], line_46[609], line_45[607], line_44[605], line_43[603], line_42[601], line_41[599], line_40[597], line_39[595], line_38[593], line_37[591], line_36[589], line_35[587], line_34[585], line_33[583], line_32[581], line_31[579], line_30[577], line_29[575], line_28[573], line_27[571], line_26[569], line_25[567], line_24[565], line_23[563], line_22[561], line_21[559], line_20[557], line_19[555], line_18[553], line_17[551], line_16[549], line_15[547], line_14[545], line_13[543], line_12[541], line_11[539], line_10[537], line_9[535], line_8[533], line_7[531], line_6[529], line_5[527], line_4[525], line_3[523], line_2[521], line_1[519] };
assign col_774 = {line_128[774], line_127[772], line_126[770], line_125[768], line_124[766], line_123[764], line_122[762], line_121[760], line_120[758], line_119[756], line_118[754], line_117[752], line_116[750], line_115[748], line_114[746], line_113[744], line_112[742], line_111[740], line_110[738], line_109[736], line_108[734], line_107[732], line_106[730], line_105[728], line_104[726], line_103[724], line_102[722], line_101[720], line_100[718], line_99[716], line_98[714], line_97[712], line_96[710], line_95[708], line_94[706], line_93[704], line_92[702], line_91[700], line_90[698], line_89[696], line_88[694], line_87[692], line_86[690], line_85[688], line_84[686], line_83[684], line_82[682], line_81[680], line_80[678], line_79[676], line_78[674], line_77[672], line_76[670], line_75[668], line_74[666], line_73[664], line_72[662], line_71[660], line_70[658], line_69[656], line_68[654], line_67[652], line_66[650], line_65[648], line_64[646], line_63[644], line_62[642], line_61[640], line_60[638], line_59[636], line_58[634], line_57[632], line_56[630], line_55[628], line_54[626], line_53[624], line_52[622], line_51[620], line_50[618], line_49[616], line_48[614], line_47[612], line_46[610], line_45[608], line_44[606], line_43[604], line_42[602], line_41[600], line_40[598], line_39[596], line_38[594], line_37[592], line_36[590], line_35[588], line_34[586], line_33[584], line_32[582], line_31[580], line_30[578], line_29[576], line_28[574], line_27[572], line_26[570], line_25[568], line_24[566], line_23[564], line_22[562], line_21[560], line_20[558], line_19[556], line_18[554], line_17[552], line_16[550], line_15[548], line_14[546], line_13[544], line_12[542], line_11[540], line_10[538], line_9[536], line_8[534], line_7[532], line_6[530], line_5[528], line_4[526], line_3[524], line_2[522], line_1[520] };
assign col_775 = {line_128[775], line_127[773], line_126[771], line_125[769], line_124[767], line_123[765], line_122[763], line_121[761], line_120[759], line_119[757], line_118[755], line_117[753], line_116[751], line_115[749], line_114[747], line_113[745], line_112[743], line_111[741], line_110[739], line_109[737], line_108[735], line_107[733], line_106[731], line_105[729], line_104[727], line_103[725], line_102[723], line_101[721], line_100[719], line_99[717], line_98[715], line_97[713], line_96[711], line_95[709], line_94[707], line_93[705], line_92[703], line_91[701], line_90[699], line_89[697], line_88[695], line_87[693], line_86[691], line_85[689], line_84[687], line_83[685], line_82[683], line_81[681], line_80[679], line_79[677], line_78[675], line_77[673], line_76[671], line_75[669], line_74[667], line_73[665], line_72[663], line_71[661], line_70[659], line_69[657], line_68[655], line_67[653], line_66[651], line_65[649], line_64[647], line_63[645], line_62[643], line_61[641], line_60[639], line_59[637], line_58[635], line_57[633], line_56[631], line_55[629], line_54[627], line_53[625], line_52[623], line_51[621], line_50[619], line_49[617], line_48[615], line_47[613], line_46[611], line_45[609], line_44[607], line_43[605], line_42[603], line_41[601], line_40[599], line_39[597], line_38[595], line_37[593], line_36[591], line_35[589], line_34[587], line_33[585], line_32[583], line_31[581], line_30[579], line_29[577], line_28[575], line_27[573], line_26[571], line_25[569], line_24[567], line_23[565], line_22[563], line_21[561], line_20[559], line_19[557], line_18[555], line_17[553], line_16[551], line_15[549], line_14[547], line_13[545], line_12[543], line_11[541], line_10[539], line_9[537], line_8[535], line_7[533], line_6[531], line_5[529], line_4[527], line_3[525], line_2[523], line_1[521] };
assign col_776 = {line_128[776], line_127[774], line_126[772], line_125[770], line_124[768], line_123[766], line_122[764], line_121[762], line_120[760], line_119[758], line_118[756], line_117[754], line_116[752], line_115[750], line_114[748], line_113[746], line_112[744], line_111[742], line_110[740], line_109[738], line_108[736], line_107[734], line_106[732], line_105[730], line_104[728], line_103[726], line_102[724], line_101[722], line_100[720], line_99[718], line_98[716], line_97[714], line_96[712], line_95[710], line_94[708], line_93[706], line_92[704], line_91[702], line_90[700], line_89[698], line_88[696], line_87[694], line_86[692], line_85[690], line_84[688], line_83[686], line_82[684], line_81[682], line_80[680], line_79[678], line_78[676], line_77[674], line_76[672], line_75[670], line_74[668], line_73[666], line_72[664], line_71[662], line_70[660], line_69[658], line_68[656], line_67[654], line_66[652], line_65[650], line_64[648], line_63[646], line_62[644], line_61[642], line_60[640], line_59[638], line_58[636], line_57[634], line_56[632], line_55[630], line_54[628], line_53[626], line_52[624], line_51[622], line_50[620], line_49[618], line_48[616], line_47[614], line_46[612], line_45[610], line_44[608], line_43[606], line_42[604], line_41[602], line_40[600], line_39[598], line_38[596], line_37[594], line_36[592], line_35[590], line_34[588], line_33[586], line_32[584], line_31[582], line_30[580], line_29[578], line_28[576], line_27[574], line_26[572], line_25[570], line_24[568], line_23[566], line_22[564], line_21[562], line_20[560], line_19[558], line_18[556], line_17[554], line_16[552], line_15[550], line_14[548], line_13[546], line_12[544], line_11[542], line_10[540], line_9[538], line_8[536], line_7[534], line_6[532], line_5[530], line_4[528], line_3[526], line_2[524], line_1[522] };
assign col_777 = {line_128[777], line_127[775], line_126[773], line_125[771], line_124[769], line_123[767], line_122[765], line_121[763], line_120[761], line_119[759], line_118[757], line_117[755], line_116[753], line_115[751], line_114[749], line_113[747], line_112[745], line_111[743], line_110[741], line_109[739], line_108[737], line_107[735], line_106[733], line_105[731], line_104[729], line_103[727], line_102[725], line_101[723], line_100[721], line_99[719], line_98[717], line_97[715], line_96[713], line_95[711], line_94[709], line_93[707], line_92[705], line_91[703], line_90[701], line_89[699], line_88[697], line_87[695], line_86[693], line_85[691], line_84[689], line_83[687], line_82[685], line_81[683], line_80[681], line_79[679], line_78[677], line_77[675], line_76[673], line_75[671], line_74[669], line_73[667], line_72[665], line_71[663], line_70[661], line_69[659], line_68[657], line_67[655], line_66[653], line_65[651], line_64[649], line_63[647], line_62[645], line_61[643], line_60[641], line_59[639], line_58[637], line_57[635], line_56[633], line_55[631], line_54[629], line_53[627], line_52[625], line_51[623], line_50[621], line_49[619], line_48[617], line_47[615], line_46[613], line_45[611], line_44[609], line_43[607], line_42[605], line_41[603], line_40[601], line_39[599], line_38[597], line_37[595], line_36[593], line_35[591], line_34[589], line_33[587], line_32[585], line_31[583], line_30[581], line_29[579], line_28[577], line_27[575], line_26[573], line_25[571], line_24[569], line_23[567], line_22[565], line_21[563], line_20[561], line_19[559], line_18[557], line_17[555], line_16[553], line_15[551], line_14[549], line_13[547], line_12[545], line_11[543], line_10[541], line_9[539], line_8[537], line_7[535], line_6[533], line_5[531], line_4[529], line_3[527], line_2[525], line_1[523] };
assign col_778 = {line_128[778], line_127[776], line_126[774], line_125[772], line_124[770], line_123[768], line_122[766], line_121[764], line_120[762], line_119[760], line_118[758], line_117[756], line_116[754], line_115[752], line_114[750], line_113[748], line_112[746], line_111[744], line_110[742], line_109[740], line_108[738], line_107[736], line_106[734], line_105[732], line_104[730], line_103[728], line_102[726], line_101[724], line_100[722], line_99[720], line_98[718], line_97[716], line_96[714], line_95[712], line_94[710], line_93[708], line_92[706], line_91[704], line_90[702], line_89[700], line_88[698], line_87[696], line_86[694], line_85[692], line_84[690], line_83[688], line_82[686], line_81[684], line_80[682], line_79[680], line_78[678], line_77[676], line_76[674], line_75[672], line_74[670], line_73[668], line_72[666], line_71[664], line_70[662], line_69[660], line_68[658], line_67[656], line_66[654], line_65[652], line_64[650], line_63[648], line_62[646], line_61[644], line_60[642], line_59[640], line_58[638], line_57[636], line_56[634], line_55[632], line_54[630], line_53[628], line_52[626], line_51[624], line_50[622], line_49[620], line_48[618], line_47[616], line_46[614], line_45[612], line_44[610], line_43[608], line_42[606], line_41[604], line_40[602], line_39[600], line_38[598], line_37[596], line_36[594], line_35[592], line_34[590], line_33[588], line_32[586], line_31[584], line_30[582], line_29[580], line_28[578], line_27[576], line_26[574], line_25[572], line_24[570], line_23[568], line_22[566], line_21[564], line_20[562], line_19[560], line_18[558], line_17[556], line_16[554], line_15[552], line_14[550], line_13[548], line_12[546], line_11[544], line_10[542], line_9[540], line_8[538], line_7[536], line_6[534], line_5[532], line_4[530], line_3[528], line_2[526], line_1[524] };
assign col_779 = {line_128[779], line_127[777], line_126[775], line_125[773], line_124[771], line_123[769], line_122[767], line_121[765], line_120[763], line_119[761], line_118[759], line_117[757], line_116[755], line_115[753], line_114[751], line_113[749], line_112[747], line_111[745], line_110[743], line_109[741], line_108[739], line_107[737], line_106[735], line_105[733], line_104[731], line_103[729], line_102[727], line_101[725], line_100[723], line_99[721], line_98[719], line_97[717], line_96[715], line_95[713], line_94[711], line_93[709], line_92[707], line_91[705], line_90[703], line_89[701], line_88[699], line_87[697], line_86[695], line_85[693], line_84[691], line_83[689], line_82[687], line_81[685], line_80[683], line_79[681], line_78[679], line_77[677], line_76[675], line_75[673], line_74[671], line_73[669], line_72[667], line_71[665], line_70[663], line_69[661], line_68[659], line_67[657], line_66[655], line_65[653], line_64[651], line_63[649], line_62[647], line_61[645], line_60[643], line_59[641], line_58[639], line_57[637], line_56[635], line_55[633], line_54[631], line_53[629], line_52[627], line_51[625], line_50[623], line_49[621], line_48[619], line_47[617], line_46[615], line_45[613], line_44[611], line_43[609], line_42[607], line_41[605], line_40[603], line_39[601], line_38[599], line_37[597], line_36[595], line_35[593], line_34[591], line_33[589], line_32[587], line_31[585], line_30[583], line_29[581], line_28[579], line_27[577], line_26[575], line_25[573], line_24[571], line_23[569], line_22[567], line_21[565], line_20[563], line_19[561], line_18[559], line_17[557], line_16[555], line_15[553], line_14[551], line_13[549], line_12[547], line_11[545], line_10[543], line_9[541], line_8[539], line_7[537], line_6[535], line_5[533], line_4[531], line_3[529], line_2[527], line_1[525] };
assign col_780 = {line_128[780], line_127[778], line_126[776], line_125[774], line_124[772], line_123[770], line_122[768], line_121[766], line_120[764], line_119[762], line_118[760], line_117[758], line_116[756], line_115[754], line_114[752], line_113[750], line_112[748], line_111[746], line_110[744], line_109[742], line_108[740], line_107[738], line_106[736], line_105[734], line_104[732], line_103[730], line_102[728], line_101[726], line_100[724], line_99[722], line_98[720], line_97[718], line_96[716], line_95[714], line_94[712], line_93[710], line_92[708], line_91[706], line_90[704], line_89[702], line_88[700], line_87[698], line_86[696], line_85[694], line_84[692], line_83[690], line_82[688], line_81[686], line_80[684], line_79[682], line_78[680], line_77[678], line_76[676], line_75[674], line_74[672], line_73[670], line_72[668], line_71[666], line_70[664], line_69[662], line_68[660], line_67[658], line_66[656], line_65[654], line_64[652], line_63[650], line_62[648], line_61[646], line_60[644], line_59[642], line_58[640], line_57[638], line_56[636], line_55[634], line_54[632], line_53[630], line_52[628], line_51[626], line_50[624], line_49[622], line_48[620], line_47[618], line_46[616], line_45[614], line_44[612], line_43[610], line_42[608], line_41[606], line_40[604], line_39[602], line_38[600], line_37[598], line_36[596], line_35[594], line_34[592], line_33[590], line_32[588], line_31[586], line_30[584], line_29[582], line_28[580], line_27[578], line_26[576], line_25[574], line_24[572], line_23[570], line_22[568], line_21[566], line_20[564], line_19[562], line_18[560], line_17[558], line_16[556], line_15[554], line_14[552], line_13[550], line_12[548], line_11[546], line_10[544], line_9[542], line_8[540], line_7[538], line_6[536], line_5[534], line_4[532], line_3[530], line_2[528], line_1[526] };
assign col_781 = {line_128[781], line_127[779], line_126[777], line_125[775], line_124[773], line_123[771], line_122[769], line_121[767], line_120[765], line_119[763], line_118[761], line_117[759], line_116[757], line_115[755], line_114[753], line_113[751], line_112[749], line_111[747], line_110[745], line_109[743], line_108[741], line_107[739], line_106[737], line_105[735], line_104[733], line_103[731], line_102[729], line_101[727], line_100[725], line_99[723], line_98[721], line_97[719], line_96[717], line_95[715], line_94[713], line_93[711], line_92[709], line_91[707], line_90[705], line_89[703], line_88[701], line_87[699], line_86[697], line_85[695], line_84[693], line_83[691], line_82[689], line_81[687], line_80[685], line_79[683], line_78[681], line_77[679], line_76[677], line_75[675], line_74[673], line_73[671], line_72[669], line_71[667], line_70[665], line_69[663], line_68[661], line_67[659], line_66[657], line_65[655], line_64[653], line_63[651], line_62[649], line_61[647], line_60[645], line_59[643], line_58[641], line_57[639], line_56[637], line_55[635], line_54[633], line_53[631], line_52[629], line_51[627], line_50[625], line_49[623], line_48[621], line_47[619], line_46[617], line_45[615], line_44[613], line_43[611], line_42[609], line_41[607], line_40[605], line_39[603], line_38[601], line_37[599], line_36[597], line_35[595], line_34[593], line_33[591], line_32[589], line_31[587], line_30[585], line_29[583], line_28[581], line_27[579], line_26[577], line_25[575], line_24[573], line_23[571], line_22[569], line_21[567], line_20[565], line_19[563], line_18[561], line_17[559], line_16[557], line_15[555], line_14[553], line_13[551], line_12[549], line_11[547], line_10[545], line_9[543], line_8[541], line_7[539], line_6[537], line_5[535], line_4[533], line_3[531], line_2[529], line_1[527] };
assign col_782 = {line_128[782], line_127[780], line_126[778], line_125[776], line_124[774], line_123[772], line_122[770], line_121[768], line_120[766], line_119[764], line_118[762], line_117[760], line_116[758], line_115[756], line_114[754], line_113[752], line_112[750], line_111[748], line_110[746], line_109[744], line_108[742], line_107[740], line_106[738], line_105[736], line_104[734], line_103[732], line_102[730], line_101[728], line_100[726], line_99[724], line_98[722], line_97[720], line_96[718], line_95[716], line_94[714], line_93[712], line_92[710], line_91[708], line_90[706], line_89[704], line_88[702], line_87[700], line_86[698], line_85[696], line_84[694], line_83[692], line_82[690], line_81[688], line_80[686], line_79[684], line_78[682], line_77[680], line_76[678], line_75[676], line_74[674], line_73[672], line_72[670], line_71[668], line_70[666], line_69[664], line_68[662], line_67[660], line_66[658], line_65[656], line_64[654], line_63[652], line_62[650], line_61[648], line_60[646], line_59[644], line_58[642], line_57[640], line_56[638], line_55[636], line_54[634], line_53[632], line_52[630], line_51[628], line_50[626], line_49[624], line_48[622], line_47[620], line_46[618], line_45[616], line_44[614], line_43[612], line_42[610], line_41[608], line_40[606], line_39[604], line_38[602], line_37[600], line_36[598], line_35[596], line_34[594], line_33[592], line_32[590], line_31[588], line_30[586], line_29[584], line_28[582], line_27[580], line_26[578], line_25[576], line_24[574], line_23[572], line_22[570], line_21[568], line_20[566], line_19[564], line_18[562], line_17[560], line_16[558], line_15[556], line_14[554], line_13[552], line_12[550], line_11[548], line_10[546], line_9[544], line_8[542], line_7[540], line_6[538], line_5[536], line_4[534], line_3[532], line_2[530], line_1[528] };
assign col_783 = {line_128[783], line_127[781], line_126[779], line_125[777], line_124[775], line_123[773], line_122[771], line_121[769], line_120[767], line_119[765], line_118[763], line_117[761], line_116[759], line_115[757], line_114[755], line_113[753], line_112[751], line_111[749], line_110[747], line_109[745], line_108[743], line_107[741], line_106[739], line_105[737], line_104[735], line_103[733], line_102[731], line_101[729], line_100[727], line_99[725], line_98[723], line_97[721], line_96[719], line_95[717], line_94[715], line_93[713], line_92[711], line_91[709], line_90[707], line_89[705], line_88[703], line_87[701], line_86[699], line_85[697], line_84[695], line_83[693], line_82[691], line_81[689], line_80[687], line_79[685], line_78[683], line_77[681], line_76[679], line_75[677], line_74[675], line_73[673], line_72[671], line_71[669], line_70[667], line_69[665], line_68[663], line_67[661], line_66[659], line_65[657], line_64[655], line_63[653], line_62[651], line_61[649], line_60[647], line_59[645], line_58[643], line_57[641], line_56[639], line_55[637], line_54[635], line_53[633], line_52[631], line_51[629], line_50[627], line_49[625], line_48[623], line_47[621], line_46[619], line_45[617], line_44[615], line_43[613], line_42[611], line_41[609], line_40[607], line_39[605], line_38[603], line_37[601], line_36[599], line_35[597], line_34[595], line_33[593], line_32[591], line_31[589], line_30[587], line_29[585], line_28[583], line_27[581], line_26[579], line_25[577], line_24[575], line_23[573], line_22[571], line_21[569], line_20[567], line_19[565], line_18[563], line_17[561], line_16[559], line_15[557], line_14[555], line_13[553], line_12[551], line_11[549], line_10[547], line_9[545], line_8[543], line_7[541], line_6[539], line_5[537], line_4[535], line_3[533], line_2[531], line_1[529] };
assign col_784 = {line_128[784], line_127[782], line_126[780], line_125[778], line_124[776], line_123[774], line_122[772], line_121[770], line_120[768], line_119[766], line_118[764], line_117[762], line_116[760], line_115[758], line_114[756], line_113[754], line_112[752], line_111[750], line_110[748], line_109[746], line_108[744], line_107[742], line_106[740], line_105[738], line_104[736], line_103[734], line_102[732], line_101[730], line_100[728], line_99[726], line_98[724], line_97[722], line_96[720], line_95[718], line_94[716], line_93[714], line_92[712], line_91[710], line_90[708], line_89[706], line_88[704], line_87[702], line_86[700], line_85[698], line_84[696], line_83[694], line_82[692], line_81[690], line_80[688], line_79[686], line_78[684], line_77[682], line_76[680], line_75[678], line_74[676], line_73[674], line_72[672], line_71[670], line_70[668], line_69[666], line_68[664], line_67[662], line_66[660], line_65[658], line_64[656], line_63[654], line_62[652], line_61[650], line_60[648], line_59[646], line_58[644], line_57[642], line_56[640], line_55[638], line_54[636], line_53[634], line_52[632], line_51[630], line_50[628], line_49[626], line_48[624], line_47[622], line_46[620], line_45[618], line_44[616], line_43[614], line_42[612], line_41[610], line_40[608], line_39[606], line_38[604], line_37[602], line_36[600], line_35[598], line_34[596], line_33[594], line_32[592], line_31[590], line_30[588], line_29[586], line_28[584], line_27[582], line_26[580], line_25[578], line_24[576], line_23[574], line_22[572], line_21[570], line_20[568], line_19[566], line_18[564], line_17[562], line_16[560], line_15[558], line_14[556], line_13[554], line_12[552], line_11[550], line_10[548], line_9[546], line_8[544], line_7[542], line_6[540], line_5[538], line_4[536], line_3[534], line_2[532], line_1[530] };
assign col_785 = {line_128[785], line_127[783], line_126[781], line_125[779], line_124[777], line_123[775], line_122[773], line_121[771], line_120[769], line_119[767], line_118[765], line_117[763], line_116[761], line_115[759], line_114[757], line_113[755], line_112[753], line_111[751], line_110[749], line_109[747], line_108[745], line_107[743], line_106[741], line_105[739], line_104[737], line_103[735], line_102[733], line_101[731], line_100[729], line_99[727], line_98[725], line_97[723], line_96[721], line_95[719], line_94[717], line_93[715], line_92[713], line_91[711], line_90[709], line_89[707], line_88[705], line_87[703], line_86[701], line_85[699], line_84[697], line_83[695], line_82[693], line_81[691], line_80[689], line_79[687], line_78[685], line_77[683], line_76[681], line_75[679], line_74[677], line_73[675], line_72[673], line_71[671], line_70[669], line_69[667], line_68[665], line_67[663], line_66[661], line_65[659], line_64[657], line_63[655], line_62[653], line_61[651], line_60[649], line_59[647], line_58[645], line_57[643], line_56[641], line_55[639], line_54[637], line_53[635], line_52[633], line_51[631], line_50[629], line_49[627], line_48[625], line_47[623], line_46[621], line_45[619], line_44[617], line_43[615], line_42[613], line_41[611], line_40[609], line_39[607], line_38[605], line_37[603], line_36[601], line_35[599], line_34[597], line_33[595], line_32[593], line_31[591], line_30[589], line_29[587], line_28[585], line_27[583], line_26[581], line_25[579], line_24[577], line_23[575], line_22[573], line_21[571], line_20[569], line_19[567], line_18[565], line_17[563], line_16[561], line_15[559], line_14[557], line_13[555], line_12[553], line_11[551], line_10[549], line_9[547], line_8[545], line_7[543], line_6[541], line_5[539], line_4[537], line_3[535], line_2[533], line_1[531] };
assign col_786 = {line_128[786], line_127[784], line_126[782], line_125[780], line_124[778], line_123[776], line_122[774], line_121[772], line_120[770], line_119[768], line_118[766], line_117[764], line_116[762], line_115[760], line_114[758], line_113[756], line_112[754], line_111[752], line_110[750], line_109[748], line_108[746], line_107[744], line_106[742], line_105[740], line_104[738], line_103[736], line_102[734], line_101[732], line_100[730], line_99[728], line_98[726], line_97[724], line_96[722], line_95[720], line_94[718], line_93[716], line_92[714], line_91[712], line_90[710], line_89[708], line_88[706], line_87[704], line_86[702], line_85[700], line_84[698], line_83[696], line_82[694], line_81[692], line_80[690], line_79[688], line_78[686], line_77[684], line_76[682], line_75[680], line_74[678], line_73[676], line_72[674], line_71[672], line_70[670], line_69[668], line_68[666], line_67[664], line_66[662], line_65[660], line_64[658], line_63[656], line_62[654], line_61[652], line_60[650], line_59[648], line_58[646], line_57[644], line_56[642], line_55[640], line_54[638], line_53[636], line_52[634], line_51[632], line_50[630], line_49[628], line_48[626], line_47[624], line_46[622], line_45[620], line_44[618], line_43[616], line_42[614], line_41[612], line_40[610], line_39[608], line_38[606], line_37[604], line_36[602], line_35[600], line_34[598], line_33[596], line_32[594], line_31[592], line_30[590], line_29[588], line_28[586], line_27[584], line_26[582], line_25[580], line_24[578], line_23[576], line_22[574], line_21[572], line_20[570], line_19[568], line_18[566], line_17[564], line_16[562], line_15[560], line_14[558], line_13[556], line_12[554], line_11[552], line_10[550], line_9[548], line_8[546], line_7[544], line_6[542], line_5[540], line_4[538], line_3[536], line_2[534], line_1[532] };
assign col_787 = {line_128[787], line_127[785], line_126[783], line_125[781], line_124[779], line_123[777], line_122[775], line_121[773], line_120[771], line_119[769], line_118[767], line_117[765], line_116[763], line_115[761], line_114[759], line_113[757], line_112[755], line_111[753], line_110[751], line_109[749], line_108[747], line_107[745], line_106[743], line_105[741], line_104[739], line_103[737], line_102[735], line_101[733], line_100[731], line_99[729], line_98[727], line_97[725], line_96[723], line_95[721], line_94[719], line_93[717], line_92[715], line_91[713], line_90[711], line_89[709], line_88[707], line_87[705], line_86[703], line_85[701], line_84[699], line_83[697], line_82[695], line_81[693], line_80[691], line_79[689], line_78[687], line_77[685], line_76[683], line_75[681], line_74[679], line_73[677], line_72[675], line_71[673], line_70[671], line_69[669], line_68[667], line_67[665], line_66[663], line_65[661], line_64[659], line_63[657], line_62[655], line_61[653], line_60[651], line_59[649], line_58[647], line_57[645], line_56[643], line_55[641], line_54[639], line_53[637], line_52[635], line_51[633], line_50[631], line_49[629], line_48[627], line_47[625], line_46[623], line_45[621], line_44[619], line_43[617], line_42[615], line_41[613], line_40[611], line_39[609], line_38[607], line_37[605], line_36[603], line_35[601], line_34[599], line_33[597], line_32[595], line_31[593], line_30[591], line_29[589], line_28[587], line_27[585], line_26[583], line_25[581], line_24[579], line_23[577], line_22[575], line_21[573], line_20[571], line_19[569], line_18[567], line_17[565], line_16[563], line_15[561], line_14[559], line_13[557], line_12[555], line_11[553], line_10[551], line_9[549], line_8[547], line_7[545], line_6[543], line_5[541], line_4[539], line_3[537], line_2[535], line_1[533] };
assign col_788 = {line_128[788], line_127[786], line_126[784], line_125[782], line_124[780], line_123[778], line_122[776], line_121[774], line_120[772], line_119[770], line_118[768], line_117[766], line_116[764], line_115[762], line_114[760], line_113[758], line_112[756], line_111[754], line_110[752], line_109[750], line_108[748], line_107[746], line_106[744], line_105[742], line_104[740], line_103[738], line_102[736], line_101[734], line_100[732], line_99[730], line_98[728], line_97[726], line_96[724], line_95[722], line_94[720], line_93[718], line_92[716], line_91[714], line_90[712], line_89[710], line_88[708], line_87[706], line_86[704], line_85[702], line_84[700], line_83[698], line_82[696], line_81[694], line_80[692], line_79[690], line_78[688], line_77[686], line_76[684], line_75[682], line_74[680], line_73[678], line_72[676], line_71[674], line_70[672], line_69[670], line_68[668], line_67[666], line_66[664], line_65[662], line_64[660], line_63[658], line_62[656], line_61[654], line_60[652], line_59[650], line_58[648], line_57[646], line_56[644], line_55[642], line_54[640], line_53[638], line_52[636], line_51[634], line_50[632], line_49[630], line_48[628], line_47[626], line_46[624], line_45[622], line_44[620], line_43[618], line_42[616], line_41[614], line_40[612], line_39[610], line_38[608], line_37[606], line_36[604], line_35[602], line_34[600], line_33[598], line_32[596], line_31[594], line_30[592], line_29[590], line_28[588], line_27[586], line_26[584], line_25[582], line_24[580], line_23[578], line_22[576], line_21[574], line_20[572], line_19[570], line_18[568], line_17[566], line_16[564], line_15[562], line_14[560], line_13[558], line_12[556], line_11[554], line_10[552], line_9[550], line_8[548], line_7[546], line_6[544], line_5[542], line_4[540], line_3[538], line_2[536], line_1[534] };
assign col_789 = {line_128[789], line_127[787], line_126[785], line_125[783], line_124[781], line_123[779], line_122[777], line_121[775], line_120[773], line_119[771], line_118[769], line_117[767], line_116[765], line_115[763], line_114[761], line_113[759], line_112[757], line_111[755], line_110[753], line_109[751], line_108[749], line_107[747], line_106[745], line_105[743], line_104[741], line_103[739], line_102[737], line_101[735], line_100[733], line_99[731], line_98[729], line_97[727], line_96[725], line_95[723], line_94[721], line_93[719], line_92[717], line_91[715], line_90[713], line_89[711], line_88[709], line_87[707], line_86[705], line_85[703], line_84[701], line_83[699], line_82[697], line_81[695], line_80[693], line_79[691], line_78[689], line_77[687], line_76[685], line_75[683], line_74[681], line_73[679], line_72[677], line_71[675], line_70[673], line_69[671], line_68[669], line_67[667], line_66[665], line_65[663], line_64[661], line_63[659], line_62[657], line_61[655], line_60[653], line_59[651], line_58[649], line_57[647], line_56[645], line_55[643], line_54[641], line_53[639], line_52[637], line_51[635], line_50[633], line_49[631], line_48[629], line_47[627], line_46[625], line_45[623], line_44[621], line_43[619], line_42[617], line_41[615], line_40[613], line_39[611], line_38[609], line_37[607], line_36[605], line_35[603], line_34[601], line_33[599], line_32[597], line_31[595], line_30[593], line_29[591], line_28[589], line_27[587], line_26[585], line_25[583], line_24[581], line_23[579], line_22[577], line_21[575], line_20[573], line_19[571], line_18[569], line_17[567], line_16[565], line_15[563], line_14[561], line_13[559], line_12[557], line_11[555], line_10[553], line_9[551], line_8[549], line_7[547], line_6[545], line_5[543], line_4[541], line_3[539], line_2[537], line_1[535] };
assign col_790 = {line_128[790], line_127[788], line_126[786], line_125[784], line_124[782], line_123[780], line_122[778], line_121[776], line_120[774], line_119[772], line_118[770], line_117[768], line_116[766], line_115[764], line_114[762], line_113[760], line_112[758], line_111[756], line_110[754], line_109[752], line_108[750], line_107[748], line_106[746], line_105[744], line_104[742], line_103[740], line_102[738], line_101[736], line_100[734], line_99[732], line_98[730], line_97[728], line_96[726], line_95[724], line_94[722], line_93[720], line_92[718], line_91[716], line_90[714], line_89[712], line_88[710], line_87[708], line_86[706], line_85[704], line_84[702], line_83[700], line_82[698], line_81[696], line_80[694], line_79[692], line_78[690], line_77[688], line_76[686], line_75[684], line_74[682], line_73[680], line_72[678], line_71[676], line_70[674], line_69[672], line_68[670], line_67[668], line_66[666], line_65[664], line_64[662], line_63[660], line_62[658], line_61[656], line_60[654], line_59[652], line_58[650], line_57[648], line_56[646], line_55[644], line_54[642], line_53[640], line_52[638], line_51[636], line_50[634], line_49[632], line_48[630], line_47[628], line_46[626], line_45[624], line_44[622], line_43[620], line_42[618], line_41[616], line_40[614], line_39[612], line_38[610], line_37[608], line_36[606], line_35[604], line_34[602], line_33[600], line_32[598], line_31[596], line_30[594], line_29[592], line_28[590], line_27[588], line_26[586], line_25[584], line_24[582], line_23[580], line_22[578], line_21[576], line_20[574], line_19[572], line_18[570], line_17[568], line_16[566], line_15[564], line_14[562], line_13[560], line_12[558], line_11[556], line_10[554], line_9[552], line_8[550], line_7[548], line_6[546], line_5[544], line_4[542], line_3[540], line_2[538], line_1[536] };
assign col_791 = {line_128[791], line_127[789], line_126[787], line_125[785], line_124[783], line_123[781], line_122[779], line_121[777], line_120[775], line_119[773], line_118[771], line_117[769], line_116[767], line_115[765], line_114[763], line_113[761], line_112[759], line_111[757], line_110[755], line_109[753], line_108[751], line_107[749], line_106[747], line_105[745], line_104[743], line_103[741], line_102[739], line_101[737], line_100[735], line_99[733], line_98[731], line_97[729], line_96[727], line_95[725], line_94[723], line_93[721], line_92[719], line_91[717], line_90[715], line_89[713], line_88[711], line_87[709], line_86[707], line_85[705], line_84[703], line_83[701], line_82[699], line_81[697], line_80[695], line_79[693], line_78[691], line_77[689], line_76[687], line_75[685], line_74[683], line_73[681], line_72[679], line_71[677], line_70[675], line_69[673], line_68[671], line_67[669], line_66[667], line_65[665], line_64[663], line_63[661], line_62[659], line_61[657], line_60[655], line_59[653], line_58[651], line_57[649], line_56[647], line_55[645], line_54[643], line_53[641], line_52[639], line_51[637], line_50[635], line_49[633], line_48[631], line_47[629], line_46[627], line_45[625], line_44[623], line_43[621], line_42[619], line_41[617], line_40[615], line_39[613], line_38[611], line_37[609], line_36[607], line_35[605], line_34[603], line_33[601], line_32[599], line_31[597], line_30[595], line_29[593], line_28[591], line_27[589], line_26[587], line_25[585], line_24[583], line_23[581], line_22[579], line_21[577], line_20[575], line_19[573], line_18[571], line_17[569], line_16[567], line_15[565], line_14[563], line_13[561], line_12[559], line_11[557], line_10[555], line_9[553], line_8[551], line_7[549], line_6[547], line_5[545], line_4[543], line_3[541], line_2[539], line_1[537] };
assign col_792 = {line_128[792], line_127[790], line_126[788], line_125[786], line_124[784], line_123[782], line_122[780], line_121[778], line_120[776], line_119[774], line_118[772], line_117[770], line_116[768], line_115[766], line_114[764], line_113[762], line_112[760], line_111[758], line_110[756], line_109[754], line_108[752], line_107[750], line_106[748], line_105[746], line_104[744], line_103[742], line_102[740], line_101[738], line_100[736], line_99[734], line_98[732], line_97[730], line_96[728], line_95[726], line_94[724], line_93[722], line_92[720], line_91[718], line_90[716], line_89[714], line_88[712], line_87[710], line_86[708], line_85[706], line_84[704], line_83[702], line_82[700], line_81[698], line_80[696], line_79[694], line_78[692], line_77[690], line_76[688], line_75[686], line_74[684], line_73[682], line_72[680], line_71[678], line_70[676], line_69[674], line_68[672], line_67[670], line_66[668], line_65[666], line_64[664], line_63[662], line_62[660], line_61[658], line_60[656], line_59[654], line_58[652], line_57[650], line_56[648], line_55[646], line_54[644], line_53[642], line_52[640], line_51[638], line_50[636], line_49[634], line_48[632], line_47[630], line_46[628], line_45[626], line_44[624], line_43[622], line_42[620], line_41[618], line_40[616], line_39[614], line_38[612], line_37[610], line_36[608], line_35[606], line_34[604], line_33[602], line_32[600], line_31[598], line_30[596], line_29[594], line_28[592], line_27[590], line_26[588], line_25[586], line_24[584], line_23[582], line_22[580], line_21[578], line_20[576], line_19[574], line_18[572], line_17[570], line_16[568], line_15[566], line_14[564], line_13[562], line_12[560], line_11[558], line_10[556], line_9[554], line_8[552], line_7[550], line_6[548], line_5[546], line_4[544], line_3[542], line_2[540], line_1[538] };
assign col_793 = {line_128[793], line_127[791], line_126[789], line_125[787], line_124[785], line_123[783], line_122[781], line_121[779], line_120[777], line_119[775], line_118[773], line_117[771], line_116[769], line_115[767], line_114[765], line_113[763], line_112[761], line_111[759], line_110[757], line_109[755], line_108[753], line_107[751], line_106[749], line_105[747], line_104[745], line_103[743], line_102[741], line_101[739], line_100[737], line_99[735], line_98[733], line_97[731], line_96[729], line_95[727], line_94[725], line_93[723], line_92[721], line_91[719], line_90[717], line_89[715], line_88[713], line_87[711], line_86[709], line_85[707], line_84[705], line_83[703], line_82[701], line_81[699], line_80[697], line_79[695], line_78[693], line_77[691], line_76[689], line_75[687], line_74[685], line_73[683], line_72[681], line_71[679], line_70[677], line_69[675], line_68[673], line_67[671], line_66[669], line_65[667], line_64[665], line_63[663], line_62[661], line_61[659], line_60[657], line_59[655], line_58[653], line_57[651], line_56[649], line_55[647], line_54[645], line_53[643], line_52[641], line_51[639], line_50[637], line_49[635], line_48[633], line_47[631], line_46[629], line_45[627], line_44[625], line_43[623], line_42[621], line_41[619], line_40[617], line_39[615], line_38[613], line_37[611], line_36[609], line_35[607], line_34[605], line_33[603], line_32[601], line_31[599], line_30[597], line_29[595], line_28[593], line_27[591], line_26[589], line_25[587], line_24[585], line_23[583], line_22[581], line_21[579], line_20[577], line_19[575], line_18[573], line_17[571], line_16[569], line_15[567], line_14[565], line_13[563], line_12[561], line_11[559], line_10[557], line_9[555], line_8[553], line_7[551], line_6[549], line_5[547], line_4[545], line_3[543], line_2[541], line_1[539] };
assign col_794 = {line_128[794], line_127[792], line_126[790], line_125[788], line_124[786], line_123[784], line_122[782], line_121[780], line_120[778], line_119[776], line_118[774], line_117[772], line_116[770], line_115[768], line_114[766], line_113[764], line_112[762], line_111[760], line_110[758], line_109[756], line_108[754], line_107[752], line_106[750], line_105[748], line_104[746], line_103[744], line_102[742], line_101[740], line_100[738], line_99[736], line_98[734], line_97[732], line_96[730], line_95[728], line_94[726], line_93[724], line_92[722], line_91[720], line_90[718], line_89[716], line_88[714], line_87[712], line_86[710], line_85[708], line_84[706], line_83[704], line_82[702], line_81[700], line_80[698], line_79[696], line_78[694], line_77[692], line_76[690], line_75[688], line_74[686], line_73[684], line_72[682], line_71[680], line_70[678], line_69[676], line_68[674], line_67[672], line_66[670], line_65[668], line_64[666], line_63[664], line_62[662], line_61[660], line_60[658], line_59[656], line_58[654], line_57[652], line_56[650], line_55[648], line_54[646], line_53[644], line_52[642], line_51[640], line_50[638], line_49[636], line_48[634], line_47[632], line_46[630], line_45[628], line_44[626], line_43[624], line_42[622], line_41[620], line_40[618], line_39[616], line_38[614], line_37[612], line_36[610], line_35[608], line_34[606], line_33[604], line_32[602], line_31[600], line_30[598], line_29[596], line_28[594], line_27[592], line_26[590], line_25[588], line_24[586], line_23[584], line_22[582], line_21[580], line_20[578], line_19[576], line_18[574], line_17[572], line_16[570], line_15[568], line_14[566], line_13[564], line_12[562], line_11[560], line_10[558], line_9[556], line_8[554], line_7[552], line_6[550], line_5[548], line_4[546], line_3[544], line_2[542], line_1[540] };
assign col_795 = {line_128[795], line_127[793], line_126[791], line_125[789], line_124[787], line_123[785], line_122[783], line_121[781], line_120[779], line_119[777], line_118[775], line_117[773], line_116[771], line_115[769], line_114[767], line_113[765], line_112[763], line_111[761], line_110[759], line_109[757], line_108[755], line_107[753], line_106[751], line_105[749], line_104[747], line_103[745], line_102[743], line_101[741], line_100[739], line_99[737], line_98[735], line_97[733], line_96[731], line_95[729], line_94[727], line_93[725], line_92[723], line_91[721], line_90[719], line_89[717], line_88[715], line_87[713], line_86[711], line_85[709], line_84[707], line_83[705], line_82[703], line_81[701], line_80[699], line_79[697], line_78[695], line_77[693], line_76[691], line_75[689], line_74[687], line_73[685], line_72[683], line_71[681], line_70[679], line_69[677], line_68[675], line_67[673], line_66[671], line_65[669], line_64[667], line_63[665], line_62[663], line_61[661], line_60[659], line_59[657], line_58[655], line_57[653], line_56[651], line_55[649], line_54[647], line_53[645], line_52[643], line_51[641], line_50[639], line_49[637], line_48[635], line_47[633], line_46[631], line_45[629], line_44[627], line_43[625], line_42[623], line_41[621], line_40[619], line_39[617], line_38[615], line_37[613], line_36[611], line_35[609], line_34[607], line_33[605], line_32[603], line_31[601], line_30[599], line_29[597], line_28[595], line_27[593], line_26[591], line_25[589], line_24[587], line_23[585], line_22[583], line_21[581], line_20[579], line_19[577], line_18[575], line_17[573], line_16[571], line_15[569], line_14[567], line_13[565], line_12[563], line_11[561], line_10[559], line_9[557], line_8[555], line_7[553], line_6[551], line_5[549], line_4[547], line_3[545], line_2[543], line_1[541] };
assign col_796 = {line_128[796], line_127[794], line_126[792], line_125[790], line_124[788], line_123[786], line_122[784], line_121[782], line_120[780], line_119[778], line_118[776], line_117[774], line_116[772], line_115[770], line_114[768], line_113[766], line_112[764], line_111[762], line_110[760], line_109[758], line_108[756], line_107[754], line_106[752], line_105[750], line_104[748], line_103[746], line_102[744], line_101[742], line_100[740], line_99[738], line_98[736], line_97[734], line_96[732], line_95[730], line_94[728], line_93[726], line_92[724], line_91[722], line_90[720], line_89[718], line_88[716], line_87[714], line_86[712], line_85[710], line_84[708], line_83[706], line_82[704], line_81[702], line_80[700], line_79[698], line_78[696], line_77[694], line_76[692], line_75[690], line_74[688], line_73[686], line_72[684], line_71[682], line_70[680], line_69[678], line_68[676], line_67[674], line_66[672], line_65[670], line_64[668], line_63[666], line_62[664], line_61[662], line_60[660], line_59[658], line_58[656], line_57[654], line_56[652], line_55[650], line_54[648], line_53[646], line_52[644], line_51[642], line_50[640], line_49[638], line_48[636], line_47[634], line_46[632], line_45[630], line_44[628], line_43[626], line_42[624], line_41[622], line_40[620], line_39[618], line_38[616], line_37[614], line_36[612], line_35[610], line_34[608], line_33[606], line_32[604], line_31[602], line_30[600], line_29[598], line_28[596], line_27[594], line_26[592], line_25[590], line_24[588], line_23[586], line_22[584], line_21[582], line_20[580], line_19[578], line_18[576], line_17[574], line_16[572], line_15[570], line_14[568], line_13[566], line_12[564], line_11[562], line_10[560], line_9[558], line_8[556], line_7[554], line_6[552], line_5[550], line_4[548], line_3[546], line_2[544], line_1[542] };
assign col_797 = {line_128[797], line_127[795], line_126[793], line_125[791], line_124[789], line_123[787], line_122[785], line_121[783], line_120[781], line_119[779], line_118[777], line_117[775], line_116[773], line_115[771], line_114[769], line_113[767], line_112[765], line_111[763], line_110[761], line_109[759], line_108[757], line_107[755], line_106[753], line_105[751], line_104[749], line_103[747], line_102[745], line_101[743], line_100[741], line_99[739], line_98[737], line_97[735], line_96[733], line_95[731], line_94[729], line_93[727], line_92[725], line_91[723], line_90[721], line_89[719], line_88[717], line_87[715], line_86[713], line_85[711], line_84[709], line_83[707], line_82[705], line_81[703], line_80[701], line_79[699], line_78[697], line_77[695], line_76[693], line_75[691], line_74[689], line_73[687], line_72[685], line_71[683], line_70[681], line_69[679], line_68[677], line_67[675], line_66[673], line_65[671], line_64[669], line_63[667], line_62[665], line_61[663], line_60[661], line_59[659], line_58[657], line_57[655], line_56[653], line_55[651], line_54[649], line_53[647], line_52[645], line_51[643], line_50[641], line_49[639], line_48[637], line_47[635], line_46[633], line_45[631], line_44[629], line_43[627], line_42[625], line_41[623], line_40[621], line_39[619], line_38[617], line_37[615], line_36[613], line_35[611], line_34[609], line_33[607], line_32[605], line_31[603], line_30[601], line_29[599], line_28[597], line_27[595], line_26[593], line_25[591], line_24[589], line_23[587], line_22[585], line_21[583], line_20[581], line_19[579], line_18[577], line_17[575], line_16[573], line_15[571], line_14[569], line_13[567], line_12[565], line_11[563], line_10[561], line_9[559], line_8[557], line_7[555], line_6[553], line_5[551], line_4[549], line_3[547], line_2[545], line_1[543] };
assign col_798 = {line_128[798], line_127[796], line_126[794], line_125[792], line_124[790], line_123[788], line_122[786], line_121[784], line_120[782], line_119[780], line_118[778], line_117[776], line_116[774], line_115[772], line_114[770], line_113[768], line_112[766], line_111[764], line_110[762], line_109[760], line_108[758], line_107[756], line_106[754], line_105[752], line_104[750], line_103[748], line_102[746], line_101[744], line_100[742], line_99[740], line_98[738], line_97[736], line_96[734], line_95[732], line_94[730], line_93[728], line_92[726], line_91[724], line_90[722], line_89[720], line_88[718], line_87[716], line_86[714], line_85[712], line_84[710], line_83[708], line_82[706], line_81[704], line_80[702], line_79[700], line_78[698], line_77[696], line_76[694], line_75[692], line_74[690], line_73[688], line_72[686], line_71[684], line_70[682], line_69[680], line_68[678], line_67[676], line_66[674], line_65[672], line_64[670], line_63[668], line_62[666], line_61[664], line_60[662], line_59[660], line_58[658], line_57[656], line_56[654], line_55[652], line_54[650], line_53[648], line_52[646], line_51[644], line_50[642], line_49[640], line_48[638], line_47[636], line_46[634], line_45[632], line_44[630], line_43[628], line_42[626], line_41[624], line_40[622], line_39[620], line_38[618], line_37[616], line_36[614], line_35[612], line_34[610], line_33[608], line_32[606], line_31[604], line_30[602], line_29[600], line_28[598], line_27[596], line_26[594], line_25[592], line_24[590], line_23[588], line_22[586], line_21[584], line_20[582], line_19[580], line_18[578], line_17[576], line_16[574], line_15[572], line_14[570], line_13[568], line_12[566], line_11[564], line_10[562], line_9[560], line_8[558], line_7[556], line_6[554], line_5[552], line_4[550], line_3[548], line_2[546], line_1[544] };
assign col_799 = {line_128[799], line_127[797], line_126[795], line_125[793], line_124[791], line_123[789], line_122[787], line_121[785], line_120[783], line_119[781], line_118[779], line_117[777], line_116[775], line_115[773], line_114[771], line_113[769], line_112[767], line_111[765], line_110[763], line_109[761], line_108[759], line_107[757], line_106[755], line_105[753], line_104[751], line_103[749], line_102[747], line_101[745], line_100[743], line_99[741], line_98[739], line_97[737], line_96[735], line_95[733], line_94[731], line_93[729], line_92[727], line_91[725], line_90[723], line_89[721], line_88[719], line_87[717], line_86[715], line_85[713], line_84[711], line_83[709], line_82[707], line_81[705], line_80[703], line_79[701], line_78[699], line_77[697], line_76[695], line_75[693], line_74[691], line_73[689], line_72[687], line_71[685], line_70[683], line_69[681], line_68[679], line_67[677], line_66[675], line_65[673], line_64[671], line_63[669], line_62[667], line_61[665], line_60[663], line_59[661], line_58[659], line_57[657], line_56[655], line_55[653], line_54[651], line_53[649], line_52[647], line_51[645], line_50[643], line_49[641], line_48[639], line_47[637], line_46[635], line_45[633], line_44[631], line_43[629], line_42[627], line_41[625], line_40[623], line_39[621], line_38[619], line_37[617], line_36[615], line_35[613], line_34[611], line_33[609], line_32[607], line_31[605], line_30[603], line_29[601], line_28[599], line_27[597], line_26[595], line_25[593], line_24[591], line_23[589], line_22[587], line_21[585], line_20[583], line_19[581], line_18[579], line_17[577], line_16[575], line_15[573], line_14[571], line_13[569], line_12[567], line_11[565], line_10[563], line_9[561], line_8[559], line_7[557], line_6[555], line_5[553], line_4[551], line_3[549], line_2[547], line_1[545] };
assign col_800 = {line_128[800], line_127[798], line_126[796], line_125[794], line_124[792], line_123[790], line_122[788], line_121[786], line_120[784], line_119[782], line_118[780], line_117[778], line_116[776], line_115[774], line_114[772], line_113[770], line_112[768], line_111[766], line_110[764], line_109[762], line_108[760], line_107[758], line_106[756], line_105[754], line_104[752], line_103[750], line_102[748], line_101[746], line_100[744], line_99[742], line_98[740], line_97[738], line_96[736], line_95[734], line_94[732], line_93[730], line_92[728], line_91[726], line_90[724], line_89[722], line_88[720], line_87[718], line_86[716], line_85[714], line_84[712], line_83[710], line_82[708], line_81[706], line_80[704], line_79[702], line_78[700], line_77[698], line_76[696], line_75[694], line_74[692], line_73[690], line_72[688], line_71[686], line_70[684], line_69[682], line_68[680], line_67[678], line_66[676], line_65[674], line_64[672], line_63[670], line_62[668], line_61[666], line_60[664], line_59[662], line_58[660], line_57[658], line_56[656], line_55[654], line_54[652], line_53[650], line_52[648], line_51[646], line_50[644], line_49[642], line_48[640], line_47[638], line_46[636], line_45[634], line_44[632], line_43[630], line_42[628], line_41[626], line_40[624], line_39[622], line_38[620], line_37[618], line_36[616], line_35[614], line_34[612], line_33[610], line_32[608], line_31[606], line_30[604], line_29[602], line_28[600], line_27[598], line_26[596], line_25[594], line_24[592], line_23[590], line_22[588], line_21[586], line_20[584], line_19[582], line_18[580], line_17[578], line_16[576], line_15[574], line_14[572], line_13[570], line_12[568], line_11[566], line_10[564], line_9[562], line_8[560], line_7[558], line_6[556], line_5[554], line_4[552], line_3[550], line_2[548], line_1[546] };
assign col_801 = {line_128[801], line_127[799], line_126[797], line_125[795], line_124[793], line_123[791], line_122[789], line_121[787], line_120[785], line_119[783], line_118[781], line_117[779], line_116[777], line_115[775], line_114[773], line_113[771], line_112[769], line_111[767], line_110[765], line_109[763], line_108[761], line_107[759], line_106[757], line_105[755], line_104[753], line_103[751], line_102[749], line_101[747], line_100[745], line_99[743], line_98[741], line_97[739], line_96[737], line_95[735], line_94[733], line_93[731], line_92[729], line_91[727], line_90[725], line_89[723], line_88[721], line_87[719], line_86[717], line_85[715], line_84[713], line_83[711], line_82[709], line_81[707], line_80[705], line_79[703], line_78[701], line_77[699], line_76[697], line_75[695], line_74[693], line_73[691], line_72[689], line_71[687], line_70[685], line_69[683], line_68[681], line_67[679], line_66[677], line_65[675], line_64[673], line_63[671], line_62[669], line_61[667], line_60[665], line_59[663], line_58[661], line_57[659], line_56[657], line_55[655], line_54[653], line_53[651], line_52[649], line_51[647], line_50[645], line_49[643], line_48[641], line_47[639], line_46[637], line_45[635], line_44[633], line_43[631], line_42[629], line_41[627], line_40[625], line_39[623], line_38[621], line_37[619], line_36[617], line_35[615], line_34[613], line_33[611], line_32[609], line_31[607], line_30[605], line_29[603], line_28[601], line_27[599], line_26[597], line_25[595], line_24[593], line_23[591], line_22[589], line_21[587], line_20[585], line_19[583], line_18[581], line_17[579], line_16[577], line_15[575], line_14[573], line_13[571], line_12[569], line_11[567], line_10[565], line_9[563], line_8[561], line_7[559], line_6[557], line_5[555], line_4[553], line_3[551], line_2[549], line_1[547] };
assign col_802 = {line_128[802], line_127[800], line_126[798], line_125[796], line_124[794], line_123[792], line_122[790], line_121[788], line_120[786], line_119[784], line_118[782], line_117[780], line_116[778], line_115[776], line_114[774], line_113[772], line_112[770], line_111[768], line_110[766], line_109[764], line_108[762], line_107[760], line_106[758], line_105[756], line_104[754], line_103[752], line_102[750], line_101[748], line_100[746], line_99[744], line_98[742], line_97[740], line_96[738], line_95[736], line_94[734], line_93[732], line_92[730], line_91[728], line_90[726], line_89[724], line_88[722], line_87[720], line_86[718], line_85[716], line_84[714], line_83[712], line_82[710], line_81[708], line_80[706], line_79[704], line_78[702], line_77[700], line_76[698], line_75[696], line_74[694], line_73[692], line_72[690], line_71[688], line_70[686], line_69[684], line_68[682], line_67[680], line_66[678], line_65[676], line_64[674], line_63[672], line_62[670], line_61[668], line_60[666], line_59[664], line_58[662], line_57[660], line_56[658], line_55[656], line_54[654], line_53[652], line_52[650], line_51[648], line_50[646], line_49[644], line_48[642], line_47[640], line_46[638], line_45[636], line_44[634], line_43[632], line_42[630], line_41[628], line_40[626], line_39[624], line_38[622], line_37[620], line_36[618], line_35[616], line_34[614], line_33[612], line_32[610], line_31[608], line_30[606], line_29[604], line_28[602], line_27[600], line_26[598], line_25[596], line_24[594], line_23[592], line_22[590], line_21[588], line_20[586], line_19[584], line_18[582], line_17[580], line_16[578], line_15[576], line_14[574], line_13[572], line_12[570], line_11[568], line_10[566], line_9[564], line_8[562], line_7[560], line_6[558], line_5[556], line_4[554], line_3[552], line_2[550], line_1[548] };
assign col_803 = {line_128[803], line_127[801], line_126[799], line_125[797], line_124[795], line_123[793], line_122[791], line_121[789], line_120[787], line_119[785], line_118[783], line_117[781], line_116[779], line_115[777], line_114[775], line_113[773], line_112[771], line_111[769], line_110[767], line_109[765], line_108[763], line_107[761], line_106[759], line_105[757], line_104[755], line_103[753], line_102[751], line_101[749], line_100[747], line_99[745], line_98[743], line_97[741], line_96[739], line_95[737], line_94[735], line_93[733], line_92[731], line_91[729], line_90[727], line_89[725], line_88[723], line_87[721], line_86[719], line_85[717], line_84[715], line_83[713], line_82[711], line_81[709], line_80[707], line_79[705], line_78[703], line_77[701], line_76[699], line_75[697], line_74[695], line_73[693], line_72[691], line_71[689], line_70[687], line_69[685], line_68[683], line_67[681], line_66[679], line_65[677], line_64[675], line_63[673], line_62[671], line_61[669], line_60[667], line_59[665], line_58[663], line_57[661], line_56[659], line_55[657], line_54[655], line_53[653], line_52[651], line_51[649], line_50[647], line_49[645], line_48[643], line_47[641], line_46[639], line_45[637], line_44[635], line_43[633], line_42[631], line_41[629], line_40[627], line_39[625], line_38[623], line_37[621], line_36[619], line_35[617], line_34[615], line_33[613], line_32[611], line_31[609], line_30[607], line_29[605], line_28[603], line_27[601], line_26[599], line_25[597], line_24[595], line_23[593], line_22[591], line_21[589], line_20[587], line_19[585], line_18[583], line_17[581], line_16[579], line_15[577], line_14[575], line_13[573], line_12[571], line_11[569], line_10[567], line_9[565], line_8[563], line_7[561], line_6[559], line_5[557], line_4[555], line_3[553], line_2[551], line_1[549] };
assign col_804 = {line_128[804], line_127[802], line_126[800], line_125[798], line_124[796], line_123[794], line_122[792], line_121[790], line_120[788], line_119[786], line_118[784], line_117[782], line_116[780], line_115[778], line_114[776], line_113[774], line_112[772], line_111[770], line_110[768], line_109[766], line_108[764], line_107[762], line_106[760], line_105[758], line_104[756], line_103[754], line_102[752], line_101[750], line_100[748], line_99[746], line_98[744], line_97[742], line_96[740], line_95[738], line_94[736], line_93[734], line_92[732], line_91[730], line_90[728], line_89[726], line_88[724], line_87[722], line_86[720], line_85[718], line_84[716], line_83[714], line_82[712], line_81[710], line_80[708], line_79[706], line_78[704], line_77[702], line_76[700], line_75[698], line_74[696], line_73[694], line_72[692], line_71[690], line_70[688], line_69[686], line_68[684], line_67[682], line_66[680], line_65[678], line_64[676], line_63[674], line_62[672], line_61[670], line_60[668], line_59[666], line_58[664], line_57[662], line_56[660], line_55[658], line_54[656], line_53[654], line_52[652], line_51[650], line_50[648], line_49[646], line_48[644], line_47[642], line_46[640], line_45[638], line_44[636], line_43[634], line_42[632], line_41[630], line_40[628], line_39[626], line_38[624], line_37[622], line_36[620], line_35[618], line_34[616], line_33[614], line_32[612], line_31[610], line_30[608], line_29[606], line_28[604], line_27[602], line_26[600], line_25[598], line_24[596], line_23[594], line_22[592], line_21[590], line_20[588], line_19[586], line_18[584], line_17[582], line_16[580], line_15[578], line_14[576], line_13[574], line_12[572], line_11[570], line_10[568], line_9[566], line_8[564], line_7[562], line_6[560], line_5[558], line_4[556], line_3[554], line_2[552], line_1[550] };
assign col_805 = {line_128[805], line_127[803], line_126[801], line_125[799], line_124[797], line_123[795], line_122[793], line_121[791], line_120[789], line_119[787], line_118[785], line_117[783], line_116[781], line_115[779], line_114[777], line_113[775], line_112[773], line_111[771], line_110[769], line_109[767], line_108[765], line_107[763], line_106[761], line_105[759], line_104[757], line_103[755], line_102[753], line_101[751], line_100[749], line_99[747], line_98[745], line_97[743], line_96[741], line_95[739], line_94[737], line_93[735], line_92[733], line_91[731], line_90[729], line_89[727], line_88[725], line_87[723], line_86[721], line_85[719], line_84[717], line_83[715], line_82[713], line_81[711], line_80[709], line_79[707], line_78[705], line_77[703], line_76[701], line_75[699], line_74[697], line_73[695], line_72[693], line_71[691], line_70[689], line_69[687], line_68[685], line_67[683], line_66[681], line_65[679], line_64[677], line_63[675], line_62[673], line_61[671], line_60[669], line_59[667], line_58[665], line_57[663], line_56[661], line_55[659], line_54[657], line_53[655], line_52[653], line_51[651], line_50[649], line_49[647], line_48[645], line_47[643], line_46[641], line_45[639], line_44[637], line_43[635], line_42[633], line_41[631], line_40[629], line_39[627], line_38[625], line_37[623], line_36[621], line_35[619], line_34[617], line_33[615], line_32[613], line_31[611], line_30[609], line_29[607], line_28[605], line_27[603], line_26[601], line_25[599], line_24[597], line_23[595], line_22[593], line_21[591], line_20[589], line_19[587], line_18[585], line_17[583], line_16[581], line_15[579], line_14[577], line_13[575], line_12[573], line_11[571], line_10[569], line_9[567], line_8[565], line_7[563], line_6[561], line_5[559], line_4[557], line_3[555], line_2[553], line_1[551] };
assign col_806 = {line_128[806], line_127[804], line_126[802], line_125[800], line_124[798], line_123[796], line_122[794], line_121[792], line_120[790], line_119[788], line_118[786], line_117[784], line_116[782], line_115[780], line_114[778], line_113[776], line_112[774], line_111[772], line_110[770], line_109[768], line_108[766], line_107[764], line_106[762], line_105[760], line_104[758], line_103[756], line_102[754], line_101[752], line_100[750], line_99[748], line_98[746], line_97[744], line_96[742], line_95[740], line_94[738], line_93[736], line_92[734], line_91[732], line_90[730], line_89[728], line_88[726], line_87[724], line_86[722], line_85[720], line_84[718], line_83[716], line_82[714], line_81[712], line_80[710], line_79[708], line_78[706], line_77[704], line_76[702], line_75[700], line_74[698], line_73[696], line_72[694], line_71[692], line_70[690], line_69[688], line_68[686], line_67[684], line_66[682], line_65[680], line_64[678], line_63[676], line_62[674], line_61[672], line_60[670], line_59[668], line_58[666], line_57[664], line_56[662], line_55[660], line_54[658], line_53[656], line_52[654], line_51[652], line_50[650], line_49[648], line_48[646], line_47[644], line_46[642], line_45[640], line_44[638], line_43[636], line_42[634], line_41[632], line_40[630], line_39[628], line_38[626], line_37[624], line_36[622], line_35[620], line_34[618], line_33[616], line_32[614], line_31[612], line_30[610], line_29[608], line_28[606], line_27[604], line_26[602], line_25[600], line_24[598], line_23[596], line_22[594], line_21[592], line_20[590], line_19[588], line_18[586], line_17[584], line_16[582], line_15[580], line_14[578], line_13[576], line_12[574], line_11[572], line_10[570], line_9[568], line_8[566], line_7[564], line_6[562], line_5[560], line_4[558], line_3[556], line_2[554], line_1[552] };
assign col_807 = {line_128[807], line_127[805], line_126[803], line_125[801], line_124[799], line_123[797], line_122[795], line_121[793], line_120[791], line_119[789], line_118[787], line_117[785], line_116[783], line_115[781], line_114[779], line_113[777], line_112[775], line_111[773], line_110[771], line_109[769], line_108[767], line_107[765], line_106[763], line_105[761], line_104[759], line_103[757], line_102[755], line_101[753], line_100[751], line_99[749], line_98[747], line_97[745], line_96[743], line_95[741], line_94[739], line_93[737], line_92[735], line_91[733], line_90[731], line_89[729], line_88[727], line_87[725], line_86[723], line_85[721], line_84[719], line_83[717], line_82[715], line_81[713], line_80[711], line_79[709], line_78[707], line_77[705], line_76[703], line_75[701], line_74[699], line_73[697], line_72[695], line_71[693], line_70[691], line_69[689], line_68[687], line_67[685], line_66[683], line_65[681], line_64[679], line_63[677], line_62[675], line_61[673], line_60[671], line_59[669], line_58[667], line_57[665], line_56[663], line_55[661], line_54[659], line_53[657], line_52[655], line_51[653], line_50[651], line_49[649], line_48[647], line_47[645], line_46[643], line_45[641], line_44[639], line_43[637], line_42[635], line_41[633], line_40[631], line_39[629], line_38[627], line_37[625], line_36[623], line_35[621], line_34[619], line_33[617], line_32[615], line_31[613], line_30[611], line_29[609], line_28[607], line_27[605], line_26[603], line_25[601], line_24[599], line_23[597], line_22[595], line_21[593], line_20[591], line_19[589], line_18[587], line_17[585], line_16[583], line_15[581], line_14[579], line_13[577], line_12[575], line_11[573], line_10[571], line_9[569], line_8[567], line_7[565], line_6[563], line_5[561], line_4[559], line_3[557], line_2[555], line_1[553] };
assign col_808 = {line_128[808], line_127[806], line_126[804], line_125[802], line_124[800], line_123[798], line_122[796], line_121[794], line_120[792], line_119[790], line_118[788], line_117[786], line_116[784], line_115[782], line_114[780], line_113[778], line_112[776], line_111[774], line_110[772], line_109[770], line_108[768], line_107[766], line_106[764], line_105[762], line_104[760], line_103[758], line_102[756], line_101[754], line_100[752], line_99[750], line_98[748], line_97[746], line_96[744], line_95[742], line_94[740], line_93[738], line_92[736], line_91[734], line_90[732], line_89[730], line_88[728], line_87[726], line_86[724], line_85[722], line_84[720], line_83[718], line_82[716], line_81[714], line_80[712], line_79[710], line_78[708], line_77[706], line_76[704], line_75[702], line_74[700], line_73[698], line_72[696], line_71[694], line_70[692], line_69[690], line_68[688], line_67[686], line_66[684], line_65[682], line_64[680], line_63[678], line_62[676], line_61[674], line_60[672], line_59[670], line_58[668], line_57[666], line_56[664], line_55[662], line_54[660], line_53[658], line_52[656], line_51[654], line_50[652], line_49[650], line_48[648], line_47[646], line_46[644], line_45[642], line_44[640], line_43[638], line_42[636], line_41[634], line_40[632], line_39[630], line_38[628], line_37[626], line_36[624], line_35[622], line_34[620], line_33[618], line_32[616], line_31[614], line_30[612], line_29[610], line_28[608], line_27[606], line_26[604], line_25[602], line_24[600], line_23[598], line_22[596], line_21[594], line_20[592], line_19[590], line_18[588], line_17[586], line_16[584], line_15[582], line_14[580], line_13[578], line_12[576], line_11[574], line_10[572], line_9[570], line_8[568], line_7[566], line_6[564], line_5[562], line_4[560], line_3[558], line_2[556], line_1[554] };
assign col_809 = {line_128[809], line_127[807], line_126[805], line_125[803], line_124[801], line_123[799], line_122[797], line_121[795], line_120[793], line_119[791], line_118[789], line_117[787], line_116[785], line_115[783], line_114[781], line_113[779], line_112[777], line_111[775], line_110[773], line_109[771], line_108[769], line_107[767], line_106[765], line_105[763], line_104[761], line_103[759], line_102[757], line_101[755], line_100[753], line_99[751], line_98[749], line_97[747], line_96[745], line_95[743], line_94[741], line_93[739], line_92[737], line_91[735], line_90[733], line_89[731], line_88[729], line_87[727], line_86[725], line_85[723], line_84[721], line_83[719], line_82[717], line_81[715], line_80[713], line_79[711], line_78[709], line_77[707], line_76[705], line_75[703], line_74[701], line_73[699], line_72[697], line_71[695], line_70[693], line_69[691], line_68[689], line_67[687], line_66[685], line_65[683], line_64[681], line_63[679], line_62[677], line_61[675], line_60[673], line_59[671], line_58[669], line_57[667], line_56[665], line_55[663], line_54[661], line_53[659], line_52[657], line_51[655], line_50[653], line_49[651], line_48[649], line_47[647], line_46[645], line_45[643], line_44[641], line_43[639], line_42[637], line_41[635], line_40[633], line_39[631], line_38[629], line_37[627], line_36[625], line_35[623], line_34[621], line_33[619], line_32[617], line_31[615], line_30[613], line_29[611], line_28[609], line_27[607], line_26[605], line_25[603], line_24[601], line_23[599], line_22[597], line_21[595], line_20[593], line_19[591], line_18[589], line_17[587], line_16[585], line_15[583], line_14[581], line_13[579], line_12[577], line_11[575], line_10[573], line_9[571], line_8[569], line_7[567], line_6[565], line_5[563], line_4[561], line_3[559], line_2[557], line_1[555] };
assign col_810 = {line_128[810], line_127[808], line_126[806], line_125[804], line_124[802], line_123[800], line_122[798], line_121[796], line_120[794], line_119[792], line_118[790], line_117[788], line_116[786], line_115[784], line_114[782], line_113[780], line_112[778], line_111[776], line_110[774], line_109[772], line_108[770], line_107[768], line_106[766], line_105[764], line_104[762], line_103[760], line_102[758], line_101[756], line_100[754], line_99[752], line_98[750], line_97[748], line_96[746], line_95[744], line_94[742], line_93[740], line_92[738], line_91[736], line_90[734], line_89[732], line_88[730], line_87[728], line_86[726], line_85[724], line_84[722], line_83[720], line_82[718], line_81[716], line_80[714], line_79[712], line_78[710], line_77[708], line_76[706], line_75[704], line_74[702], line_73[700], line_72[698], line_71[696], line_70[694], line_69[692], line_68[690], line_67[688], line_66[686], line_65[684], line_64[682], line_63[680], line_62[678], line_61[676], line_60[674], line_59[672], line_58[670], line_57[668], line_56[666], line_55[664], line_54[662], line_53[660], line_52[658], line_51[656], line_50[654], line_49[652], line_48[650], line_47[648], line_46[646], line_45[644], line_44[642], line_43[640], line_42[638], line_41[636], line_40[634], line_39[632], line_38[630], line_37[628], line_36[626], line_35[624], line_34[622], line_33[620], line_32[618], line_31[616], line_30[614], line_29[612], line_28[610], line_27[608], line_26[606], line_25[604], line_24[602], line_23[600], line_22[598], line_21[596], line_20[594], line_19[592], line_18[590], line_17[588], line_16[586], line_15[584], line_14[582], line_13[580], line_12[578], line_11[576], line_10[574], line_9[572], line_8[570], line_7[568], line_6[566], line_5[564], line_4[562], line_3[560], line_2[558], line_1[556] };
assign col_811 = {line_128[811], line_127[809], line_126[807], line_125[805], line_124[803], line_123[801], line_122[799], line_121[797], line_120[795], line_119[793], line_118[791], line_117[789], line_116[787], line_115[785], line_114[783], line_113[781], line_112[779], line_111[777], line_110[775], line_109[773], line_108[771], line_107[769], line_106[767], line_105[765], line_104[763], line_103[761], line_102[759], line_101[757], line_100[755], line_99[753], line_98[751], line_97[749], line_96[747], line_95[745], line_94[743], line_93[741], line_92[739], line_91[737], line_90[735], line_89[733], line_88[731], line_87[729], line_86[727], line_85[725], line_84[723], line_83[721], line_82[719], line_81[717], line_80[715], line_79[713], line_78[711], line_77[709], line_76[707], line_75[705], line_74[703], line_73[701], line_72[699], line_71[697], line_70[695], line_69[693], line_68[691], line_67[689], line_66[687], line_65[685], line_64[683], line_63[681], line_62[679], line_61[677], line_60[675], line_59[673], line_58[671], line_57[669], line_56[667], line_55[665], line_54[663], line_53[661], line_52[659], line_51[657], line_50[655], line_49[653], line_48[651], line_47[649], line_46[647], line_45[645], line_44[643], line_43[641], line_42[639], line_41[637], line_40[635], line_39[633], line_38[631], line_37[629], line_36[627], line_35[625], line_34[623], line_33[621], line_32[619], line_31[617], line_30[615], line_29[613], line_28[611], line_27[609], line_26[607], line_25[605], line_24[603], line_23[601], line_22[599], line_21[597], line_20[595], line_19[593], line_18[591], line_17[589], line_16[587], line_15[585], line_14[583], line_13[581], line_12[579], line_11[577], line_10[575], line_9[573], line_8[571], line_7[569], line_6[567], line_5[565], line_4[563], line_3[561], line_2[559], line_1[557] };
assign col_812 = {line_128[812], line_127[810], line_126[808], line_125[806], line_124[804], line_123[802], line_122[800], line_121[798], line_120[796], line_119[794], line_118[792], line_117[790], line_116[788], line_115[786], line_114[784], line_113[782], line_112[780], line_111[778], line_110[776], line_109[774], line_108[772], line_107[770], line_106[768], line_105[766], line_104[764], line_103[762], line_102[760], line_101[758], line_100[756], line_99[754], line_98[752], line_97[750], line_96[748], line_95[746], line_94[744], line_93[742], line_92[740], line_91[738], line_90[736], line_89[734], line_88[732], line_87[730], line_86[728], line_85[726], line_84[724], line_83[722], line_82[720], line_81[718], line_80[716], line_79[714], line_78[712], line_77[710], line_76[708], line_75[706], line_74[704], line_73[702], line_72[700], line_71[698], line_70[696], line_69[694], line_68[692], line_67[690], line_66[688], line_65[686], line_64[684], line_63[682], line_62[680], line_61[678], line_60[676], line_59[674], line_58[672], line_57[670], line_56[668], line_55[666], line_54[664], line_53[662], line_52[660], line_51[658], line_50[656], line_49[654], line_48[652], line_47[650], line_46[648], line_45[646], line_44[644], line_43[642], line_42[640], line_41[638], line_40[636], line_39[634], line_38[632], line_37[630], line_36[628], line_35[626], line_34[624], line_33[622], line_32[620], line_31[618], line_30[616], line_29[614], line_28[612], line_27[610], line_26[608], line_25[606], line_24[604], line_23[602], line_22[600], line_21[598], line_20[596], line_19[594], line_18[592], line_17[590], line_16[588], line_15[586], line_14[584], line_13[582], line_12[580], line_11[578], line_10[576], line_9[574], line_8[572], line_7[570], line_6[568], line_5[566], line_4[564], line_3[562], line_2[560], line_1[558] };
assign col_813 = {line_128[813], line_127[811], line_126[809], line_125[807], line_124[805], line_123[803], line_122[801], line_121[799], line_120[797], line_119[795], line_118[793], line_117[791], line_116[789], line_115[787], line_114[785], line_113[783], line_112[781], line_111[779], line_110[777], line_109[775], line_108[773], line_107[771], line_106[769], line_105[767], line_104[765], line_103[763], line_102[761], line_101[759], line_100[757], line_99[755], line_98[753], line_97[751], line_96[749], line_95[747], line_94[745], line_93[743], line_92[741], line_91[739], line_90[737], line_89[735], line_88[733], line_87[731], line_86[729], line_85[727], line_84[725], line_83[723], line_82[721], line_81[719], line_80[717], line_79[715], line_78[713], line_77[711], line_76[709], line_75[707], line_74[705], line_73[703], line_72[701], line_71[699], line_70[697], line_69[695], line_68[693], line_67[691], line_66[689], line_65[687], line_64[685], line_63[683], line_62[681], line_61[679], line_60[677], line_59[675], line_58[673], line_57[671], line_56[669], line_55[667], line_54[665], line_53[663], line_52[661], line_51[659], line_50[657], line_49[655], line_48[653], line_47[651], line_46[649], line_45[647], line_44[645], line_43[643], line_42[641], line_41[639], line_40[637], line_39[635], line_38[633], line_37[631], line_36[629], line_35[627], line_34[625], line_33[623], line_32[621], line_31[619], line_30[617], line_29[615], line_28[613], line_27[611], line_26[609], line_25[607], line_24[605], line_23[603], line_22[601], line_21[599], line_20[597], line_19[595], line_18[593], line_17[591], line_16[589], line_15[587], line_14[585], line_13[583], line_12[581], line_11[579], line_10[577], line_9[575], line_8[573], line_7[571], line_6[569], line_5[567], line_4[565], line_3[563], line_2[561], line_1[559] };
assign col_814 = {line_128[814], line_127[812], line_126[810], line_125[808], line_124[806], line_123[804], line_122[802], line_121[800], line_120[798], line_119[796], line_118[794], line_117[792], line_116[790], line_115[788], line_114[786], line_113[784], line_112[782], line_111[780], line_110[778], line_109[776], line_108[774], line_107[772], line_106[770], line_105[768], line_104[766], line_103[764], line_102[762], line_101[760], line_100[758], line_99[756], line_98[754], line_97[752], line_96[750], line_95[748], line_94[746], line_93[744], line_92[742], line_91[740], line_90[738], line_89[736], line_88[734], line_87[732], line_86[730], line_85[728], line_84[726], line_83[724], line_82[722], line_81[720], line_80[718], line_79[716], line_78[714], line_77[712], line_76[710], line_75[708], line_74[706], line_73[704], line_72[702], line_71[700], line_70[698], line_69[696], line_68[694], line_67[692], line_66[690], line_65[688], line_64[686], line_63[684], line_62[682], line_61[680], line_60[678], line_59[676], line_58[674], line_57[672], line_56[670], line_55[668], line_54[666], line_53[664], line_52[662], line_51[660], line_50[658], line_49[656], line_48[654], line_47[652], line_46[650], line_45[648], line_44[646], line_43[644], line_42[642], line_41[640], line_40[638], line_39[636], line_38[634], line_37[632], line_36[630], line_35[628], line_34[626], line_33[624], line_32[622], line_31[620], line_30[618], line_29[616], line_28[614], line_27[612], line_26[610], line_25[608], line_24[606], line_23[604], line_22[602], line_21[600], line_20[598], line_19[596], line_18[594], line_17[592], line_16[590], line_15[588], line_14[586], line_13[584], line_12[582], line_11[580], line_10[578], line_9[576], line_8[574], line_7[572], line_6[570], line_5[568], line_4[566], line_3[564], line_2[562], line_1[560] };
assign col_815 = {line_128[815], line_127[813], line_126[811], line_125[809], line_124[807], line_123[805], line_122[803], line_121[801], line_120[799], line_119[797], line_118[795], line_117[793], line_116[791], line_115[789], line_114[787], line_113[785], line_112[783], line_111[781], line_110[779], line_109[777], line_108[775], line_107[773], line_106[771], line_105[769], line_104[767], line_103[765], line_102[763], line_101[761], line_100[759], line_99[757], line_98[755], line_97[753], line_96[751], line_95[749], line_94[747], line_93[745], line_92[743], line_91[741], line_90[739], line_89[737], line_88[735], line_87[733], line_86[731], line_85[729], line_84[727], line_83[725], line_82[723], line_81[721], line_80[719], line_79[717], line_78[715], line_77[713], line_76[711], line_75[709], line_74[707], line_73[705], line_72[703], line_71[701], line_70[699], line_69[697], line_68[695], line_67[693], line_66[691], line_65[689], line_64[687], line_63[685], line_62[683], line_61[681], line_60[679], line_59[677], line_58[675], line_57[673], line_56[671], line_55[669], line_54[667], line_53[665], line_52[663], line_51[661], line_50[659], line_49[657], line_48[655], line_47[653], line_46[651], line_45[649], line_44[647], line_43[645], line_42[643], line_41[641], line_40[639], line_39[637], line_38[635], line_37[633], line_36[631], line_35[629], line_34[627], line_33[625], line_32[623], line_31[621], line_30[619], line_29[617], line_28[615], line_27[613], line_26[611], line_25[609], line_24[607], line_23[605], line_22[603], line_21[601], line_20[599], line_19[597], line_18[595], line_17[593], line_16[591], line_15[589], line_14[587], line_13[585], line_12[583], line_11[581], line_10[579], line_9[577], line_8[575], line_7[573], line_6[571], line_5[569], line_4[567], line_3[565], line_2[563], line_1[561] };
assign col_816 = {line_128[816], line_127[814], line_126[812], line_125[810], line_124[808], line_123[806], line_122[804], line_121[802], line_120[800], line_119[798], line_118[796], line_117[794], line_116[792], line_115[790], line_114[788], line_113[786], line_112[784], line_111[782], line_110[780], line_109[778], line_108[776], line_107[774], line_106[772], line_105[770], line_104[768], line_103[766], line_102[764], line_101[762], line_100[760], line_99[758], line_98[756], line_97[754], line_96[752], line_95[750], line_94[748], line_93[746], line_92[744], line_91[742], line_90[740], line_89[738], line_88[736], line_87[734], line_86[732], line_85[730], line_84[728], line_83[726], line_82[724], line_81[722], line_80[720], line_79[718], line_78[716], line_77[714], line_76[712], line_75[710], line_74[708], line_73[706], line_72[704], line_71[702], line_70[700], line_69[698], line_68[696], line_67[694], line_66[692], line_65[690], line_64[688], line_63[686], line_62[684], line_61[682], line_60[680], line_59[678], line_58[676], line_57[674], line_56[672], line_55[670], line_54[668], line_53[666], line_52[664], line_51[662], line_50[660], line_49[658], line_48[656], line_47[654], line_46[652], line_45[650], line_44[648], line_43[646], line_42[644], line_41[642], line_40[640], line_39[638], line_38[636], line_37[634], line_36[632], line_35[630], line_34[628], line_33[626], line_32[624], line_31[622], line_30[620], line_29[618], line_28[616], line_27[614], line_26[612], line_25[610], line_24[608], line_23[606], line_22[604], line_21[602], line_20[600], line_19[598], line_18[596], line_17[594], line_16[592], line_15[590], line_14[588], line_13[586], line_12[584], line_11[582], line_10[580], line_9[578], line_8[576], line_7[574], line_6[572], line_5[570], line_4[568], line_3[566], line_2[564], line_1[562] };
assign col_817 = {line_128[817], line_127[815], line_126[813], line_125[811], line_124[809], line_123[807], line_122[805], line_121[803], line_120[801], line_119[799], line_118[797], line_117[795], line_116[793], line_115[791], line_114[789], line_113[787], line_112[785], line_111[783], line_110[781], line_109[779], line_108[777], line_107[775], line_106[773], line_105[771], line_104[769], line_103[767], line_102[765], line_101[763], line_100[761], line_99[759], line_98[757], line_97[755], line_96[753], line_95[751], line_94[749], line_93[747], line_92[745], line_91[743], line_90[741], line_89[739], line_88[737], line_87[735], line_86[733], line_85[731], line_84[729], line_83[727], line_82[725], line_81[723], line_80[721], line_79[719], line_78[717], line_77[715], line_76[713], line_75[711], line_74[709], line_73[707], line_72[705], line_71[703], line_70[701], line_69[699], line_68[697], line_67[695], line_66[693], line_65[691], line_64[689], line_63[687], line_62[685], line_61[683], line_60[681], line_59[679], line_58[677], line_57[675], line_56[673], line_55[671], line_54[669], line_53[667], line_52[665], line_51[663], line_50[661], line_49[659], line_48[657], line_47[655], line_46[653], line_45[651], line_44[649], line_43[647], line_42[645], line_41[643], line_40[641], line_39[639], line_38[637], line_37[635], line_36[633], line_35[631], line_34[629], line_33[627], line_32[625], line_31[623], line_30[621], line_29[619], line_28[617], line_27[615], line_26[613], line_25[611], line_24[609], line_23[607], line_22[605], line_21[603], line_20[601], line_19[599], line_18[597], line_17[595], line_16[593], line_15[591], line_14[589], line_13[587], line_12[585], line_11[583], line_10[581], line_9[579], line_8[577], line_7[575], line_6[573], line_5[571], line_4[569], line_3[567], line_2[565], line_1[563] };
assign col_818 = {line_128[818], line_127[816], line_126[814], line_125[812], line_124[810], line_123[808], line_122[806], line_121[804], line_120[802], line_119[800], line_118[798], line_117[796], line_116[794], line_115[792], line_114[790], line_113[788], line_112[786], line_111[784], line_110[782], line_109[780], line_108[778], line_107[776], line_106[774], line_105[772], line_104[770], line_103[768], line_102[766], line_101[764], line_100[762], line_99[760], line_98[758], line_97[756], line_96[754], line_95[752], line_94[750], line_93[748], line_92[746], line_91[744], line_90[742], line_89[740], line_88[738], line_87[736], line_86[734], line_85[732], line_84[730], line_83[728], line_82[726], line_81[724], line_80[722], line_79[720], line_78[718], line_77[716], line_76[714], line_75[712], line_74[710], line_73[708], line_72[706], line_71[704], line_70[702], line_69[700], line_68[698], line_67[696], line_66[694], line_65[692], line_64[690], line_63[688], line_62[686], line_61[684], line_60[682], line_59[680], line_58[678], line_57[676], line_56[674], line_55[672], line_54[670], line_53[668], line_52[666], line_51[664], line_50[662], line_49[660], line_48[658], line_47[656], line_46[654], line_45[652], line_44[650], line_43[648], line_42[646], line_41[644], line_40[642], line_39[640], line_38[638], line_37[636], line_36[634], line_35[632], line_34[630], line_33[628], line_32[626], line_31[624], line_30[622], line_29[620], line_28[618], line_27[616], line_26[614], line_25[612], line_24[610], line_23[608], line_22[606], line_21[604], line_20[602], line_19[600], line_18[598], line_17[596], line_16[594], line_15[592], line_14[590], line_13[588], line_12[586], line_11[584], line_10[582], line_9[580], line_8[578], line_7[576], line_6[574], line_5[572], line_4[570], line_3[568], line_2[566], line_1[564] };
assign col_819 = {line_128[819], line_127[817], line_126[815], line_125[813], line_124[811], line_123[809], line_122[807], line_121[805], line_120[803], line_119[801], line_118[799], line_117[797], line_116[795], line_115[793], line_114[791], line_113[789], line_112[787], line_111[785], line_110[783], line_109[781], line_108[779], line_107[777], line_106[775], line_105[773], line_104[771], line_103[769], line_102[767], line_101[765], line_100[763], line_99[761], line_98[759], line_97[757], line_96[755], line_95[753], line_94[751], line_93[749], line_92[747], line_91[745], line_90[743], line_89[741], line_88[739], line_87[737], line_86[735], line_85[733], line_84[731], line_83[729], line_82[727], line_81[725], line_80[723], line_79[721], line_78[719], line_77[717], line_76[715], line_75[713], line_74[711], line_73[709], line_72[707], line_71[705], line_70[703], line_69[701], line_68[699], line_67[697], line_66[695], line_65[693], line_64[691], line_63[689], line_62[687], line_61[685], line_60[683], line_59[681], line_58[679], line_57[677], line_56[675], line_55[673], line_54[671], line_53[669], line_52[667], line_51[665], line_50[663], line_49[661], line_48[659], line_47[657], line_46[655], line_45[653], line_44[651], line_43[649], line_42[647], line_41[645], line_40[643], line_39[641], line_38[639], line_37[637], line_36[635], line_35[633], line_34[631], line_33[629], line_32[627], line_31[625], line_30[623], line_29[621], line_28[619], line_27[617], line_26[615], line_25[613], line_24[611], line_23[609], line_22[607], line_21[605], line_20[603], line_19[601], line_18[599], line_17[597], line_16[595], line_15[593], line_14[591], line_13[589], line_12[587], line_11[585], line_10[583], line_9[581], line_8[579], line_7[577], line_6[575], line_5[573], line_4[571], line_3[569], line_2[567], line_1[565] };
assign col_820 = {line_128[820], line_127[818], line_126[816], line_125[814], line_124[812], line_123[810], line_122[808], line_121[806], line_120[804], line_119[802], line_118[800], line_117[798], line_116[796], line_115[794], line_114[792], line_113[790], line_112[788], line_111[786], line_110[784], line_109[782], line_108[780], line_107[778], line_106[776], line_105[774], line_104[772], line_103[770], line_102[768], line_101[766], line_100[764], line_99[762], line_98[760], line_97[758], line_96[756], line_95[754], line_94[752], line_93[750], line_92[748], line_91[746], line_90[744], line_89[742], line_88[740], line_87[738], line_86[736], line_85[734], line_84[732], line_83[730], line_82[728], line_81[726], line_80[724], line_79[722], line_78[720], line_77[718], line_76[716], line_75[714], line_74[712], line_73[710], line_72[708], line_71[706], line_70[704], line_69[702], line_68[700], line_67[698], line_66[696], line_65[694], line_64[692], line_63[690], line_62[688], line_61[686], line_60[684], line_59[682], line_58[680], line_57[678], line_56[676], line_55[674], line_54[672], line_53[670], line_52[668], line_51[666], line_50[664], line_49[662], line_48[660], line_47[658], line_46[656], line_45[654], line_44[652], line_43[650], line_42[648], line_41[646], line_40[644], line_39[642], line_38[640], line_37[638], line_36[636], line_35[634], line_34[632], line_33[630], line_32[628], line_31[626], line_30[624], line_29[622], line_28[620], line_27[618], line_26[616], line_25[614], line_24[612], line_23[610], line_22[608], line_21[606], line_20[604], line_19[602], line_18[600], line_17[598], line_16[596], line_15[594], line_14[592], line_13[590], line_12[588], line_11[586], line_10[584], line_9[582], line_8[580], line_7[578], line_6[576], line_5[574], line_4[572], line_3[570], line_2[568], line_1[566] };
assign col_821 = {line_128[821], line_127[819], line_126[817], line_125[815], line_124[813], line_123[811], line_122[809], line_121[807], line_120[805], line_119[803], line_118[801], line_117[799], line_116[797], line_115[795], line_114[793], line_113[791], line_112[789], line_111[787], line_110[785], line_109[783], line_108[781], line_107[779], line_106[777], line_105[775], line_104[773], line_103[771], line_102[769], line_101[767], line_100[765], line_99[763], line_98[761], line_97[759], line_96[757], line_95[755], line_94[753], line_93[751], line_92[749], line_91[747], line_90[745], line_89[743], line_88[741], line_87[739], line_86[737], line_85[735], line_84[733], line_83[731], line_82[729], line_81[727], line_80[725], line_79[723], line_78[721], line_77[719], line_76[717], line_75[715], line_74[713], line_73[711], line_72[709], line_71[707], line_70[705], line_69[703], line_68[701], line_67[699], line_66[697], line_65[695], line_64[693], line_63[691], line_62[689], line_61[687], line_60[685], line_59[683], line_58[681], line_57[679], line_56[677], line_55[675], line_54[673], line_53[671], line_52[669], line_51[667], line_50[665], line_49[663], line_48[661], line_47[659], line_46[657], line_45[655], line_44[653], line_43[651], line_42[649], line_41[647], line_40[645], line_39[643], line_38[641], line_37[639], line_36[637], line_35[635], line_34[633], line_33[631], line_32[629], line_31[627], line_30[625], line_29[623], line_28[621], line_27[619], line_26[617], line_25[615], line_24[613], line_23[611], line_22[609], line_21[607], line_20[605], line_19[603], line_18[601], line_17[599], line_16[597], line_15[595], line_14[593], line_13[591], line_12[589], line_11[587], line_10[585], line_9[583], line_8[581], line_7[579], line_6[577], line_5[575], line_4[573], line_3[571], line_2[569], line_1[567] };
assign col_822 = {line_128[822], line_127[820], line_126[818], line_125[816], line_124[814], line_123[812], line_122[810], line_121[808], line_120[806], line_119[804], line_118[802], line_117[800], line_116[798], line_115[796], line_114[794], line_113[792], line_112[790], line_111[788], line_110[786], line_109[784], line_108[782], line_107[780], line_106[778], line_105[776], line_104[774], line_103[772], line_102[770], line_101[768], line_100[766], line_99[764], line_98[762], line_97[760], line_96[758], line_95[756], line_94[754], line_93[752], line_92[750], line_91[748], line_90[746], line_89[744], line_88[742], line_87[740], line_86[738], line_85[736], line_84[734], line_83[732], line_82[730], line_81[728], line_80[726], line_79[724], line_78[722], line_77[720], line_76[718], line_75[716], line_74[714], line_73[712], line_72[710], line_71[708], line_70[706], line_69[704], line_68[702], line_67[700], line_66[698], line_65[696], line_64[694], line_63[692], line_62[690], line_61[688], line_60[686], line_59[684], line_58[682], line_57[680], line_56[678], line_55[676], line_54[674], line_53[672], line_52[670], line_51[668], line_50[666], line_49[664], line_48[662], line_47[660], line_46[658], line_45[656], line_44[654], line_43[652], line_42[650], line_41[648], line_40[646], line_39[644], line_38[642], line_37[640], line_36[638], line_35[636], line_34[634], line_33[632], line_32[630], line_31[628], line_30[626], line_29[624], line_28[622], line_27[620], line_26[618], line_25[616], line_24[614], line_23[612], line_22[610], line_21[608], line_20[606], line_19[604], line_18[602], line_17[600], line_16[598], line_15[596], line_14[594], line_13[592], line_12[590], line_11[588], line_10[586], line_9[584], line_8[582], line_7[580], line_6[578], line_5[576], line_4[574], line_3[572], line_2[570], line_1[568] };
assign col_823 = {line_128[823], line_127[821], line_126[819], line_125[817], line_124[815], line_123[813], line_122[811], line_121[809], line_120[807], line_119[805], line_118[803], line_117[801], line_116[799], line_115[797], line_114[795], line_113[793], line_112[791], line_111[789], line_110[787], line_109[785], line_108[783], line_107[781], line_106[779], line_105[777], line_104[775], line_103[773], line_102[771], line_101[769], line_100[767], line_99[765], line_98[763], line_97[761], line_96[759], line_95[757], line_94[755], line_93[753], line_92[751], line_91[749], line_90[747], line_89[745], line_88[743], line_87[741], line_86[739], line_85[737], line_84[735], line_83[733], line_82[731], line_81[729], line_80[727], line_79[725], line_78[723], line_77[721], line_76[719], line_75[717], line_74[715], line_73[713], line_72[711], line_71[709], line_70[707], line_69[705], line_68[703], line_67[701], line_66[699], line_65[697], line_64[695], line_63[693], line_62[691], line_61[689], line_60[687], line_59[685], line_58[683], line_57[681], line_56[679], line_55[677], line_54[675], line_53[673], line_52[671], line_51[669], line_50[667], line_49[665], line_48[663], line_47[661], line_46[659], line_45[657], line_44[655], line_43[653], line_42[651], line_41[649], line_40[647], line_39[645], line_38[643], line_37[641], line_36[639], line_35[637], line_34[635], line_33[633], line_32[631], line_31[629], line_30[627], line_29[625], line_28[623], line_27[621], line_26[619], line_25[617], line_24[615], line_23[613], line_22[611], line_21[609], line_20[607], line_19[605], line_18[603], line_17[601], line_16[599], line_15[597], line_14[595], line_13[593], line_12[591], line_11[589], line_10[587], line_9[585], line_8[583], line_7[581], line_6[579], line_5[577], line_4[575], line_3[573], line_2[571], line_1[569] };
assign col_824 = {line_128[824], line_127[822], line_126[820], line_125[818], line_124[816], line_123[814], line_122[812], line_121[810], line_120[808], line_119[806], line_118[804], line_117[802], line_116[800], line_115[798], line_114[796], line_113[794], line_112[792], line_111[790], line_110[788], line_109[786], line_108[784], line_107[782], line_106[780], line_105[778], line_104[776], line_103[774], line_102[772], line_101[770], line_100[768], line_99[766], line_98[764], line_97[762], line_96[760], line_95[758], line_94[756], line_93[754], line_92[752], line_91[750], line_90[748], line_89[746], line_88[744], line_87[742], line_86[740], line_85[738], line_84[736], line_83[734], line_82[732], line_81[730], line_80[728], line_79[726], line_78[724], line_77[722], line_76[720], line_75[718], line_74[716], line_73[714], line_72[712], line_71[710], line_70[708], line_69[706], line_68[704], line_67[702], line_66[700], line_65[698], line_64[696], line_63[694], line_62[692], line_61[690], line_60[688], line_59[686], line_58[684], line_57[682], line_56[680], line_55[678], line_54[676], line_53[674], line_52[672], line_51[670], line_50[668], line_49[666], line_48[664], line_47[662], line_46[660], line_45[658], line_44[656], line_43[654], line_42[652], line_41[650], line_40[648], line_39[646], line_38[644], line_37[642], line_36[640], line_35[638], line_34[636], line_33[634], line_32[632], line_31[630], line_30[628], line_29[626], line_28[624], line_27[622], line_26[620], line_25[618], line_24[616], line_23[614], line_22[612], line_21[610], line_20[608], line_19[606], line_18[604], line_17[602], line_16[600], line_15[598], line_14[596], line_13[594], line_12[592], line_11[590], line_10[588], line_9[586], line_8[584], line_7[582], line_6[580], line_5[578], line_4[576], line_3[574], line_2[572], line_1[570] };
assign col_825 = {line_128[825], line_127[823], line_126[821], line_125[819], line_124[817], line_123[815], line_122[813], line_121[811], line_120[809], line_119[807], line_118[805], line_117[803], line_116[801], line_115[799], line_114[797], line_113[795], line_112[793], line_111[791], line_110[789], line_109[787], line_108[785], line_107[783], line_106[781], line_105[779], line_104[777], line_103[775], line_102[773], line_101[771], line_100[769], line_99[767], line_98[765], line_97[763], line_96[761], line_95[759], line_94[757], line_93[755], line_92[753], line_91[751], line_90[749], line_89[747], line_88[745], line_87[743], line_86[741], line_85[739], line_84[737], line_83[735], line_82[733], line_81[731], line_80[729], line_79[727], line_78[725], line_77[723], line_76[721], line_75[719], line_74[717], line_73[715], line_72[713], line_71[711], line_70[709], line_69[707], line_68[705], line_67[703], line_66[701], line_65[699], line_64[697], line_63[695], line_62[693], line_61[691], line_60[689], line_59[687], line_58[685], line_57[683], line_56[681], line_55[679], line_54[677], line_53[675], line_52[673], line_51[671], line_50[669], line_49[667], line_48[665], line_47[663], line_46[661], line_45[659], line_44[657], line_43[655], line_42[653], line_41[651], line_40[649], line_39[647], line_38[645], line_37[643], line_36[641], line_35[639], line_34[637], line_33[635], line_32[633], line_31[631], line_30[629], line_29[627], line_28[625], line_27[623], line_26[621], line_25[619], line_24[617], line_23[615], line_22[613], line_21[611], line_20[609], line_19[607], line_18[605], line_17[603], line_16[601], line_15[599], line_14[597], line_13[595], line_12[593], line_11[591], line_10[589], line_9[587], line_8[585], line_7[583], line_6[581], line_5[579], line_4[577], line_3[575], line_2[573], line_1[571] };
assign col_826 = {line_128[826], line_127[824], line_126[822], line_125[820], line_124[818], line_123[816], line_122[814], line_121[812], line_120[810], line_119[808], line_118[806], line_117[804], line_116[802], line_115[800], line_114[798], line_113[796], line_112[794], line_111[792], line_110[790], line_109[788], line_108[786], line_107[784], line_106[782], line_105[780], line_104[778], line_103[776], line_102[774], line_101[772], line_100[770], line_99[768], line_98[766], line_97[764], line_96[762], line_95[760], line_94[758], line_93[756], line_92[754], line_91[752], line_90[750], line_89[748], line_88[746], line_87[744], line_86[742], line_85[740], line_84[738], line_83[736], line_82[734], line_81[732], line_80[730], line_79[728], line_78[726], line_77[724], line_76[722], line_75[720], line_74[718], line_73[716], line_72[714], line_71[712], line_70[710], line_69[708], line_68[706], line_67[704], line_66[702], line_65[700], line_64[698], line_63[696], line_62[694], line_61[692], line_60[690], line_59[688], line_58[686], line_57[684], line_56[682], line_55[680], line_54[678], line_53[676], line_52[674], line_51[672], line_50[670], line_49[668], line_48[666], line_47[664], line_46[662], line_45[660], line_44[658], line_43[656], line_42[654], line_41[652], line_40[650], line_39[648], line_38[646], line_37[644], line_36[642], line_35[640], line_34[638], line_33[636], line_32[634], line_31[632], line_30[630], line_29[628], line_28[626], line_27[624], line_26[622], line_25[620], line_24[618], line_23[616], line_22[614], line_21[612], line_20[610], line_19[608], line_18[606], line_17[604], line_16[602], line_15[600], line_14[598], line_13[596], line_12[594], line_11[592], line_10[590], line_9[588], line_8[586], line_7[584], line_6[582], line_5[580], line_4[578], line_3[576], line_2[574], line_1[572] };
assign col_827 = {line_128[827], line_127[825], line_126[823], line_125[821], line_124[819], line_123[817], line_122[815], line_121[813], line_120[811], line_119[809], line_118[807], line_117[805], line_116[803], line_115[801], line_114[799], line_113[797], line_112[795], line_111[793], line_110[791], line_109[789], line_108[787], line_107[785], line_106[783], line_105[781], line_104[779], line_103[777], line_102[775], line_101[773], line_100[771], line_99[769], line_98[767], line_97[765], line_96[763], line_95[761], line_94[759], line_93[757], line_92[755], line_91[753], line_90[751], line_89[749], line_88[747], line_87[745], line_86[743], line_85[741], line_84[739], line_83[737], line_82[735], line_81[733], line_80[731], line_79[729], line_78[727], line_77[725], line_76[723], line_75[721], line_74[719], line_73[717], line_72[715], line_71[713], line_70[711], line_69[709], line_68[707], line_67[705], line_66[703], line_65[701], line_64[699], line_63[697], line_62[695], line_61[693], line_60[691], line_59[689], line_58[687], line_57[685], line_56[683], line_55[681], line_54[679], line_53[677], line_52[675], line_51[673], line_50[671], line_49[669], line_48[667], line_47[665], line_46[663], line_45[661], line_44[659], line_43[657], line_42[655], line_41[653], line_40[651], line_39[649], line_38[647], line_37[645], line_36[643], line_35[641], line_34[639], line_33[637], line_32[635], line_31[633], line_30[631], line_29[629], line_28[627], line_27[625], line_26[623], line_25[621], line_24[619], line_23[617], line_22[615], line_21[613], line_20[611], line_19[609], line_18[607], line_17[605], line_16[603], line_15[601], line_14[599], line_13[597], line_12[595], line_11[593], line_10[591], line_9[589], line_8[587], line_7[585], line_6[583], line_5[581], line_4[579], line_3[577], line_2[575], line_1[573] };
assign col_828 = {line_128[828], line_127[826], line_126[824], line_125[822], line_124[820], line_123[818], line_122[816], line_121[814], line_120[812], line_119[810], line_118[808], line_117[806], line_116[804], line_115[802], line_114[800], line_113[798], line_112[796], line_111[794], line_110[792], line_109[790], line_108[788], line_107[786], line_106[784], line_105[782], line_104[780], line_103[778], line_102[776], line_101[774], line_100[772], line_99[770], line_98[768], line_97[766], line_96[764], line_95[762], line_94[760], line_93[758], line_92[756], line_91[754], line_90[752], line_89[750], line_88[748], line_87[746], line_86[744], line_85[742], line_84[740], line_83[738], line_82[736], line_81[734], line_80[732], line_79[730], line_78[728], line_77[726], line_76[724], line_75[722], line_74[720], line_73[718], line_72[716], line_71[714], line_70[712], line_69[710], line_68[708], line_67[706], line_66[704], line_65[702], line_64[700], line_63[698], line_62[696], line_61[694], line_60[692], line_59[690], line_58[688], line_57[686], line_56[684], line_55[682], line_54[680], line_53[678], line_52[676], line_51[674], line_50[672], line_49[670], line_48[668], line_47[666], line_46[664], line_45[662], line_44[660], line_43[658], line_42[656], line_41[654], line_40[652], line_39[650], line_38[648], line_37[646], line_36[644], line_35[642], line_34[640], line_33[638], line_32[636], line_31[634], line_30[632], line_29[630], line_28[628], line_27[626], line_26[624], line_25[622], line_24[620], line_23[618], line_22[616], line_21[614], line_20[612], line_19[610], line_18[608], line_17[606], line_16[604], line_15[602], line_14[600], line_13[598], line_12[596], line_11[594], line_10[592], line_9[590], line_8[588], line_7[586], line_6[584], line_5[582], line_4[580], line_3[578], line_2[576], line_1[574] };
assign col_829 = {line_128[829], line_127[827], line_126[825], line_125[823], line_124[821], line_123[819], line_122[817], line_121[815], line_120[813], line_119[811], line_118[809], line_117[807], line_116[805], line_115[803], line_114[801], line_113[799], line_112[797], line_111[795], line_110[793], line_109[791], line_108[789], line_107[787], line_106[785], line_105[783], line_104[781], line_103[779], line_102[777], line_101[775], line_100[773], line_99[771], line_98[769], line_97[767], line_96[765], line_95[763], line_94[761], line_93[759], line_92[757], line_91[755], line_90[753], line_89[751], line_88[749], line_87[747], line_86[745], line_85[743], line_84[741], line_83[739], line_82[737], line_81[735], line_80[733], line_79[731], line_78[729], line_77[727], line_76[725], line_75[723], line_74[721], line_73[719], line_72[717], line_71[715], line_70[713], line_69[711], line_68[709], line_67[707], line_66[705], line_65[703], line_64[701], line_63[699], line_62[697], line_61[695], line_60[693], line_59[691], line_58[689], line_57[687], line_56[685], line_55[683], line_54[681], line_53[679], line_52[677], line_51[675], line_50[673], line_49[671], line_48[669], line_47[667], line_46[665], line_45[663], line_44[661], line_43[659], line_42[657], line_41[655], line_40[653], line_39[651], line_38[649], line_37[647], line_36[645], line_35[643], line_34[641], line_33[639], line_32[637], line_31[635], line_30[633], line_29[631], line_28[629], line_27[627], line_26[625], line_25[623], line_24[621], line_23[619], line_22[617], line_21[615], line_20[613], line_19[611], line_18[609], line_17[607], line_16[605], line_15[603], line_14[601], line_13[599], line_12[597], line_11[595], line_10[593], line_9[591], line_8[589], line_7[587], line_6[585], line_5[583], line_4[581], line_3[579], line_2[577], line_1[575] };
assign col_830 = {line_128[830], line_127[828], line_126[826], line_125[824], line_124[822], line_123[820], line_122[818], line_121[816], line_120[814], line_119[812], line_118[810], line_117[808], line_116[806], line_115[804], line_114[802], line_113[800], line_112[798], line_111[796], line_110[794], line_109[792], line_108[790], line_107[788], line_106[786], line_105[784], line_104[782], line_103[780], line_102[778], line_101[776], line_100[774], line_99[772], line_98[770], line_97[768], line_96[766], line_95[764], line_94[762], line_93[760], line_92[758], line_91[756], line_90[754], line_89[752], line_88[750], line_87[748], line_86[746], line_85[744], line_84[742], line_83[740], line_82[738], line_81[736], line_80[734], line_79[732], line_78[730], line_77[728], line_76[726], line_75[724], line_74[722], line_73[720], line_72[718], line_71[716], line_70[714], line_69[712], line_68[710], line_67[708], line_66[706], line_65[704], line_64[702], line_63[700], line_62[698], line_61[696], line_60[694], line_59[692], line_58[690], line_57[688], line_56[686], line_55[684], line_54[682], line_53[680], line_52[678], line_51[676], line_50[674], line_49[672], line_48[670], line_47[668], line_46[666], line_45[664], line_44[662], line_43[660], line_42[658], line_41[656], line_40[654], line_39[652], line_38[650], line_37[648], line_36[646], line_35[644], line_34[642], line_33[640], line_32[638], line_31[636], line_30[634], line_29[632], line_28[630], line_27[628], line_26[626], line_25[624], line_24[622], line_23[620], line_22[618], line_21[616], line_20[614], line_19[612], line_18[610], line_17[608], line_16[606], line_15[604], line_14[602], line_13[600], line_12[598], line_11[596], line_10[594], line_9[592], line_8[590], line_7[588], line_6[586], line_5[584], line_4[582], line_3[580], line_2[578], line_1[576] };
assign col_831 = {line_128[831], line_127[829], line_126[827], line_125[825], line_124[823], line_123[821], line_122[819], line_121[817], line_120[815], line_119[813], line_118[811], line_117[809], line_116[807], line_115[805], line_114[803], line_113[801], line_112[799], line_111[797], line_110[795], line_109[793], line_108[791], line_107[789], line_106[787], line_105[785], line_104[783], line_103[781], line_102[779], line_101[777], line_100[775], line_99[773], line_98[771], line_97[769], line_96[767], line_95[765], line_94[763], line_93[761], line_92[759], line_91[757], line_90[755], line_89[753], line_88[751], line_87[749], line_86[747], line_85[745], line_84[743], line_83[741], line_82[739], line_81[737], line_80[735], line_79[733], line_78[731], line_77[729], line_76[727], line_75[725], line_74[723], line_73[721], line_72[719], line_71[717], line_70[715], line_69[713], line_68[711], line_67[709], line_66[707], line_65[705], line_64[703], line_63[701], line_62[699], line_61[697], line_60[695], line_59[693], line_58[691], line_57[689], line_56[687], line_55[685], line_54[683], line_53[681], line_52[679], line_51[677], line_50[675], line_49[673], line_48[671], line_47[669], line_46[667], line_45[665], line_44[663], line_43[661], line_42[659], line_41[657], line_40[655], line_39[653], line_38[651], line_37[649], line_36[647], line_35[645], line_34[643], line_33[641], line_32[639], line_31[637], line_30[635], line_29[633], line_28[631], line_27[629], line_26[627], line_25[625], line_24[623], line_23[621], line_22[619], line_21[617], line_20[615], line_19[613], line_18[611], line_17[609], line_16[607], line_15[605], line_14[603], line_13[601], line_12[599], line_11[597], line_10[595], line_9[593], line_8[591], line_7[589], line_6[587], line_5[585], line_4[583], line_3[581], line_2[579], line_1[577] };
assign col_832 = {line_128[832], line_127[830], line_126[828], line_125[826], line_124[824], line_123[822], line_122[820], line_121[818], line_120[816], line_119[814], line_118[812], line_117[810], line_116[808], line_115[806], line_114[804], line_113[802], line_112[800], line_111[798], line_110[796], line_109[794], line_108[792], line_107[790], line_106[788], line_105[786], line_104[784], line_103[782], line_102[780], line_101[778], line_100[776], line_99[774], line_98[772], line_97[770], line_96[768], line_95[766], line_94[764], line_93[762], line_92[760], line_91[758], line_90[756], line_89[754], line_88[752], line_87[750], line_86[748], line_85[746], line_84[744], line_83[742], line_82[740], line_81[738], line_80[736], line_79[734], line_78[732], line_77[730], line_76[728], line_75[726], line_74[724], line_73[722], line_72[720], line_71[718], line_70[716], line_69[714], line_68[712], line_67[710], line_66[708], line_65[706], line_64[704], line_63[702], line_62[700], line_61[698], line_60[696], line_59[694], line_58[692], line_57[690], line_56[688], line_55[686], line_54[684], line_53[682], line_52[680], line_51[678], line_50[676], line_49[674], line_48[672], line_47[670], line_46[668], line_45[666], line_44[664], line_43[662], line_42[660], line_41[658], line_40[656], line_39[654], line_38[652], line_37[650], line_36[648], line_35[646], line_34[644], line_33[642], line_32[640], line_31[638], line_30[636], line_29[634], line_28[632], line_27[630], line_26[628], line_25[626], line_24[624], line_23[622], line_22[620], line_21[618], line_20[616], line_19[614], line_18[612], line_17[610], line_16[608], line_15[606], line_14[604], line_13[602], line_12[600], line_11[598], line_10[596], line_9[594], line_8[592], line_7[590], line_6[588], line_5[586], line_4[584], line_3[582], line_2[580], line_1[578] };
assign col_833 = {line_128[833], line_127[831], line_126[829], line_125[827], line_124[825], line_123[823], line_122[821], line_121[819], line_120[817], line_119[815], line_118[813], line_117[811], line_116[809], line_115[807], line_114[805], line_113[803], line_112[801], line_111[799], line_110[797], line_109[795], line_108[793], line_107[791], line_106[789], line_105[787], line_104[785], line_103[783], line_102[781], line_101[779], line_100[777], line_99[775], line_98[773], line_97[771], line_96[769], line_95[767], line_94[765], line_93[763], line_92[761], line_91[759], line_90[757], line_89[755], line_88[753], line_87[751], line_86[749], line_85[747], line_84[745], line_83[743], line_82[741], line_81[739], line_80[737], line_79[735], line_78[733], line_77[731], line_76[729], line_75[727], line_74[725], line_73[723], line_72[721], line_71[719], line_70[717], line_69[715], line_68[713], line_67[711], line_66[709], line_65[707], line_64[705], line_63[703], line_62[701], line_61[699], line_60[697], line_59[695], line_58[693], line_57[691], line_56[689], line_55[687], line_54[685], line_53[683], line_52[681], line_51[679], line_50[677], line_49[675], line_48[673], line_47[671], line_46[669], line_45[667], line_44[665], line_43[663], line_42[661], line_41[659], line_40[657], line_39[655], line_38[653], line_37[651], line_36[649], line_35[647], line_34[645], line_33[643], line_32[641], line_31[639], line_30[637], line_29[635], line_28[633], line_27[631], line_26[629], line_25[627], line_24[625], line_23[623], line_22[621], line_21[619], line_20[617], line_19[615], line_18[613], line_17[611], line_16[609], line_15[607], line_14[605], line_13[603], line_12[601], line_11[599], line_10[597], line_9[595], line_8[593], line_7[591], line_6[589], line_5[587], line_4[585], line_3[583], line_2[581], line_1[579] };
assign col_834 = {line_128[834], line_127[832], line_126[830], line_125[828], line_124[826], line_123[824], line_122[822], line_121[820], line_120[818], line_119[816], line_118[814], line_117[812], line_116[810], line_115[808], line_114[806], line_113[804], line_112[802], line_111[800], line_110[798], line_109[796], line_108[794], line_107[792], line_106[790], line_105[788], line_104[786], line_103[784], line_102[782], line_101[780], line_100[778], line_99[776], line_98[774], line_97[772], line_96[770], line_95[768], line_94[766], line_93[764], line_92[762], line_91[760], line_90[758], line_89[756], line_88[754], line_87[752], line_86[750], line_85[748], line_84[746], line_83[744], line_82[742], line_81[740], line_80[738], line_79[736], line_78[734], line_77[732], line_76[730], line_75[728], line_74[726], line_73[724], line_72[722], line_71[720], line_70[718], line_69[716], line_68[714], line_67[712], line_66[710], line_65[708], line_64[706], line_63[704], line_62[702], line_61[700], line_60[698], line_59[696], line_58[694], line_57[692], line_56[690], line_55[688], line_54[686], line_53[684], line_52[682], line_51[680], line_50[678], line_49[676], line_48[674], line_47[672], line_46[670], line_45[668], line_44[666], line_43[664], line_42[662], line_41[660], line_40[658], line_39[656], line_38[654], line_37[652], line_36[650], line_35[648], line_34[646], line_33[644], line_32[642], line_31[640], line_30[638], line_29[636], line_28[634], line_27[632], line_26[630], line_25[628], line_24[626], line_23[624], line_22[622], line_21[620], line_20[618], line_19[616], line_18[614], line_17[612], line_16[610], line_15[608], line_14[606], line_13[604], line_12[602], line_11[600], line_10[598], line_9[596], line_8[594], line_7[592], line_6[590], line_5[588], line_4[586], line_3[584], line_2[582], line_1[580] };
assign col_835 = {line_128[835], line_127[833], line_126[831], line_125[829], line_124[827], line_123[825], line_122[823], line_121[821], line_120[819], line_119[817], line_118[815], line_117[813], line_116[811], line_115[809], line_114[807], line_113[805], line_112[803], line_111[801], line_110[799], line_109[797], line_108[795], line_107[793], line_106[791], line_105[789], line_104[787], line_103[785], line_102[783], line_101[781], line_100[779], line_99[777], line_98[775], line_97[773], line_96[771], line_95[769], line_94[767], line_93[765], line_92[763], line_91[761], line_90[759], line_89[757], line_88[755], line_87[753], line_86[751], line_85[749], line_84[747], line_83[745], line_82[743], line_81[741], line_80[739], line_79[737], line_78[735], line_77[733], line_76[731], line_75[729], line_74[727], line_73[725], line_72[723], line_71[721], line_70[719], line_69[717], line_68[715], line_67[713], line_66[711], line_65[709], line_64[707], line_63[705], line_62[703], line_61[701], line_60[699], line_59[697], line_58[695], line_57[693], line_56[691], line_55[689], line_54[687], line_53[685], line_52[683], line_51[681], line_50[679], line_49[677], line_48[675], line_47[673], line_46[671], line_45[669], line_44[667], line_43[665], line_42[663], line_41[661], line_40[659], line_39[657], line_38[655], line_37[653], line_36[651], line_35[649], line_34[647], line_33[645], line_32[643], line_31[641], line_30[639], line_29[637], line_28[635], line_27[633], line_26[631], line_25[629], line_24[627], line_23[625], line_22[623], line_21[621], line_20[619], line_19[617], line_18[615], line_17[613], line_16[611], line_15[609], line_14[607], line_13[605], line_12[603], line_11[601], line_10[599], line_9[597], line_8[595], line_7[593], line_6[591], line_5[589], line_4[587], line_3[585], line_2[583], line_1[581] };
assign col_836 = {line_128[836], line_127[834], line_126[832], line_125[830], line_124[828], line_123[826], line_122[824], line_121[822], line_120[820], line_119[818], line_118[816], line_117[814], line_116[812], line_115[810], line_114[808], line_113[806], line_112[804], line_111[802], line_110[800], line_109[798], line_108[796], line_107[794], line_106[792], line_105[790], line_104[788], line_103[786], line_102[784], line_101[782], line_100[780], line_99[778], line_98[776], line_97[774], line_96[772], line_95[770], line_94[768], line_93[766], line_92[764], line_91[762], line_90[760], line_89[758], line_88[756], line_87[754], line_86[752], line_85[750], line_84[748], line_83[746], line_82[744], line_81[742], line_80[740], line_79[738], line_78[736], line_77[734], line_76[732], line_75[730], line_74[728], line_73[726], line_72[724], line_71[722], line_70[720], line_69[718], line_68[716], line_67[714], line_66[712], line_65[710], line_64[708], line_63[706], line_62[704], line_61[702], line_60[700], line_59[698], line_58[696], line_57[694], line_56[692], line_55[690], line_54[688], line_53[686], line_52[684], line_51[682], line_50[680], line_49[678], line_48[676], line_47[674], line_46[672], line_45[670], line_44[668], line_43[666], line_42[664], line_41[662], line_40[660], line_39[658], line_38[656], line_37[654], line_36[652], line_35[650], line_34[648], line_33[646], line_32[644], line_31[642], line_30[640], line_29[638], line_28[636], line_27[634], line_26[632], line_25[630], line_24[628], line_23[626], line_22[624], line_21[622], line_20[620], line_19[618], line_18[616], line_17[614], line_16[612], line_15[610], line_14[608], line_13[606], line_12[604], line_11[602], line_10[600], line_9[598], line_8[596], line_7[594], line_6[592], line_5[590], line_4[588], line_3[586], line_2[584], line_1[582] };
assign col_837 = {line_128[837], line_127[835], line_126[833], line_125[831], line_124[829], line_123[827], line_122[825], line_121[823], line_120[821], line_119[819], line_118[817], line_117[815], line_116[813], line_115[811], line_114[809], line_113[807], line_112[805], line_111[803], line_110[801], line_109[799], line_108[797], line_107[795], line_106[793], line_105[791], line_104[789], line_103[787], line_102[785], line_101[783], line_100[781], line_99[779], line_98[777], line_97[775], line_96[773], line_95[771], line_94[769], line_93[767], line_92[765], line_91[763], line_90[761], line_89[759], line_88[757], line_87[755], line_86[753], line_85[751], line_84[749], line_83[747], line_82[745], line_81[743], line_80[741], line_79[739], line_78[737], line_77[735], line_76[733], line_75[731], line_74[729], line_73[727], line_72[725], line_71[723], line_70[721], line_69[719], line_68[717], line_67[715], line_66[713], line_65[711], line_64[709], line_63[707], line_62[705], line_61[703], line_60[701], line_59[699], line_58[697], line_57[695], line_56[693], line_55[691], line_54[689], line_53[687], line_52[685], line_51[683], line_50[681], line_49[679], line_48[677], line_47[675], line_46[673], line_45[671], line_44[669], line_43[667], line_42[665], line_41[663], line_40[661], line_39[659], line_38[657], line_37[655], line_36[653], line_35[651], line_34[649], line_33[647], line_32[645], line_31[643], line_30[641], line_29[639], line_28[637], line_27[635], line_26[633], line_25[631], line_24[629], line_23[627], line_22[625], line_21[623], line_20[621], line_19[619], line_18[617], line_17[615], line_16[613], line_15[611], line_14[609], line_13[607], line_12[605], line_11[603], line_10[601], line_9[599], line_8[597], line_7[595], line_6[593], line_5[591], line_4[589], line_3[587], line_2[585], line_1[583] };
assign col_838 = {line_128[838], line_127[836], line_126[834], line_125[832], line_124[830], line_123[828], line_122[826], line_121[824], line_120[822], line_119[820], line_118[818], line_117[816], line_116[814], line_115[812], line_114[810], line_113[808], line_112[806], line_111[804], line_110[802], line_109[800], line_108[798], line_107[796], line_106[794], line_105[792], line_104[790], line_103[788], line_102[786], line_101[784], line_100[782], line_99[780], line_98[778], line_97[776], line_96[774], line_95[772], line_94[770], line_93[768], line_92[766], line_91[764], line_90[762], line_89[760], line_88[758], line_87[756], line_86[754], line_85[752], line_84[750], line_83[748], line_82[746], line_81[744], line_80[742], line_79[740], line_78[738], line_77[736], line_76[734], line_75[732], line_74[730], line_73[728], line_72[726], line_71[724], line_70[722], line_69[720], line_68[718], line_67[716], line_66[714], line_65[712], line_64[710], line_63[708], line_62[706], line_61[704], line_60[702], line_59[700], line_58[698], line_57[696], line_56[694], line_55[692], line_54[690], line_53[688], line_52[686], line_51[684], line_50[682], line_49[680], line_48[678], line_47[676], line_46[674], line_45[672], line_44[670], line_43[668], line_42[666], line_41[664], line_40[662], line_39[660], line_38[658], line_37[656], line_36[654], line_35[652], line_34[650], line_33[648], line_32[646], line_31[644], line_30[642], line_29[640], line_28[638], line_27[636], line_26[634], line_25[632], line_24[630], line_23[628], line_22[626], line_21[624], line_20[622], line_19[620], line_18[618], line_17[616], line_16[614], line_15[612], line_14[610], line_13[608], line_12[606], line_11[604], line_10[602], line_9[600], line_8[598], line_7[596], line_6[594], line_5[592], line_4[590], line_3[588], line_2[586], line_1[584] };
assign col_839 = {line_128[839], line_127[837], line_126[835], line_125[833], line_124[831], line_123[829], line_122[827], line_121[825], line_120[823], line_119[821], line_118[819], line_117[817], line_116[815], line_115[813], line_114[811], line_113[809], line_112[807], line_111[805], line_110[803], line_109[801], line_108[799], line_107[797], line_106[795], line_105[793], line_104[791], line_103[789], line_102[787], line_101[785], line_100[783], line_99[781], line_98[779], line_97[777], line_96[775], line_95[773], line_94[771], line_93[769], line_92[767], line_91[765], line_90[763], line_89[761], line_88[759], line_87[757], line_86[755], line_85[753], line_84[751], line_83[749], line_82[747], line_81[745], line_80[743], line_79[741], line_78[739], line_77[737], line_76[735], line_75[733], line_74[731], line_73[729], line_72[727], line_71[725], line_70[723], line_69[721], line_68[719], line_67[717], line_66[715], line_65[713], line_64[711], line_63[709], line_62[707], line_61[705], line_60[703], line_59[701], line_58[699], line_57[697], line_56[695], line_55[693], line_54[691], line_53[689], line_52[687], line_51[685], line_50[683], line_49[681], line_48[679], line_47[677], line_46[675], line_45[673], line_44[671], line_43[669], line_42[667], line_41[665], line_40[663], line_39[661], line_38[659], line_37[657], line_36[655], line_35[653], line_34[651], line_33[649], line_32[647], line_31[645], line_30[643], line_29[641], line_28[639], line_27[637], line_26[635], line_25[633], line_24[631], line_23[629], line_22[627], line_21[625], line_20[623], line_19[621], line_18[619], line_17[617], line_16[615], line_15[613], line_14[611], line_13[609], line_12[607], line_11[605], line_10[603], line_9[601], line_8[599], line_7[597], line_6[595], line_5[593], line_4[591], line_3[589], line_2[587], line_1[585] };
assign col_840 = {line_128[840], line_127[838], line_126[836], line_125[834], line_124[832], line_123[830], line_122[828], line_121[826], line_120[824], line_119[822], line_118[820], line_117[818], line_116[816], line_115[814], line_114[812], line_113[810], line_112[808], line_111[806], line_110[804], line_109[802], line_108[800], line_107[798], line_106[796], line_105[794], line_104[792], line_103[790], line_102[788], line_101[786], line_100[784], line_99[782], line_98[780], line_97[778], line_96[776], line_95[774], line_94[772], line_93[770], line_92[768], line_91[766], line_90[764], line_89[762], line_88[760], line_87[758], line_86[756], line_85[754], line_84[752], line_83[750], line_82[748], line_81[746], line_80[744], line_79[742], line_78[740], line_77[738], line_76[736], line_75[734], line_74[732], line_73[730], line_72[728], line_71[726], line_70[724], line_69[722], line_68[720], line_67[718], line_66[716], line_65[714], line_64[712], line_63[710], line_62[708], line_61[706], line_60[704], line_59[702], line_58[700], line_57[698], line_56[696], line_55[694], line_54[692], line_53[690], line_52[688], line_51[686], line_50[684], line_49[682], line_48[680], line_47[678], line_46[676], line_45[674], line_44[672], line_43[670], line_42[668], line_41[666], line_40[664], line_39[662], line_38[660], line_37[658], line_36[656], line_35[654], line_34[652], line_33[650], line_32[648], line_31[646], line_30[644], line_29[642], line_28[640], line_27[638], line_26[636], line_25[634], line_24[632], line_23[630], line_22[628], line_21[626], line_20[624], line_19[622], line_18[620], line_17[618], line_16[616], line_15[614], line_14[612], line_13[610], line_12[608], line_11[606], line_10[604], line_9[602], line_8[600], line_7[598], line_6[596], line_5[594], line_4[592], line_3[590], line_2[588], line_1[586] };
assign col_841 = {line_128[841], line_127[839], line_126[837], line_125[835], line_124[833], line_123[831], line_122[829], line_121[827], line_120[825], line_119[823], line_118[821], line_117[819], line_116[817], line_115[815], line_114[813], line_113[811], line_112[809], line_111[807], line_110[805], line_109[803], line_108[801], line_107[799], line_106[797], line_105[795], line_104[793], line_103[791], line_102[789], line_101[787], line_100[785], line_99[783], line_98[781], line_97[779], line_96[777], line_95[775], line_94[773], line_93[771], line_92[769], line_91[767], line_90[765], line_89[763], line_88[761], line_87[759], line_86[757], line_85[755], line_84[753], line_83[751], line_82[749], line_81[747], line_80[745], line_79[743], line_78[741], line_77[739], line_76[737], line_75[735], line_74[733], line_73[731], line_72[729], line_71[727], line_70[725], line_69[723], line_68[721], line_67[719], line_66[717], line_65[715], line_64[713], line_63[711], line_62[709], line_61[707], line_60[705], line_59[703], line_58[701], line_57[699], line_56[697], line_55[695], line_54[693], line_53[691], line_52[689], line_51[687], line_50[685], line_49[683], line_48[681], line_47[679], line_46[677], line_45[675], line_44[673], line_43[671], line_42[669], line_41[667], line_40[665], line_39[663], line_38[661], line_37[659], line_36[657], line_35[655], line_34[653], line_33[651], line_32[649], line_31[647], line_30[645], line_29[643], line_28[641], line_27[639], line_26[637], line_25[635], line_24[633], line_23[631], line_22[629], line_21[627], line_20[625], line_19[623], line_18[621], line_17[619], line_16[617], line_15[615], line_14[613], line_13[611], line_12[609], line_11[607], line_10[605], line_9[603], line_8[601], line_7[599], line_6[597], line_5[595], line_4[593], line_3[591], line_2[589], line_1[587] };
assign col_842 = {line_128[842], line_127[840], line_126[838], line_125[836], line_124[834], line_123[832], line_122[830], line_121[828], line_120[826], line_119[824], line_118[822], line_117[820], line_116[818], line_115[816], line_114[814], line_113[812], line_112[810], line_111[808], line_110[806], line_109[804], line_108[802], line_107[800], line_106[798], line_105[796], line_104[794], line_103[792], line_102[790], line_101[788], line_100[786], line_99[784], line_98[782], line_97[780], line_96[778], line_95[776], line_94[774], line_93[772], line_92[770], line_91[768], line_90[766], line_89[764], line_88[762], line_87[760], line_86[758], line_85[756], line_84[754], line_83[752], line_82[750], line_81[748], line_80[746], line_79[744], line_78[742], line_77[740], line_76[738], line_75[736], line_74[734], line_73[732], line_72[730], line_71[728], line_70[726], line_69[724], line_68[722], line_67[720], line_66[718], line_65[716], line_64[714], line_63[712], line_62[710], line_61[708], line_60[706], line_59[704], line_58[702], line_57[700], line_56[698], line_55[696], line_54[694], line_53[692], line_52[690], line_51[688], line_50[686], line_49[684], line_48[682], line_47[680], line_46[678], line_45[676], line_44[674], line_43[672], line_42[670], line_41[668], line_40[666], line_39[664], line_38[662], line_37[660], line_36[658], line_35[656], line_34[654], line_33[652], line_32[650], line_31[648], line_30[646], line_29[644], line_28[642], line_27[640], line_26[638], line_25[636], line_24[634], line_23[632], line_22[630], line_21[628], line_20[626], line_19[624], line_18[622], line_17[620], line_16[618], line_15[616], line_14[614], line_13[612], line_12[610], line_11[608], line_10[606], line_9[604], line_8[602], line_7[600], line_6[598], line_5[596], line_4[594], line_3[592], line_2[590], line_1[588] };
assign col_843 = {line_128[843], line_127[841], line_126[839], line_125[837], line_124[835], line_123[833], line_122[831], line_121[829], line_120[827], line_119[825], line_118[823], line_117[821], line_116[819], line_115[817], line_114[815], line_113[813], line_112[811], line_111[809], line_110[807], line_109[805], line_108[803], line_107[801], line_106[799], line_105[797], line_104[795], line_103[793], line_102[791], line_101[789], line_100[787], line_99[785], line_98[783], line_97[781], line_96[779], line_95[777], line_94[775], line_93[773], line_92[771], line_91[769], line_90[767], line_89[765], line_88[763], line_87[761], line_86[759], line_85[757], line_84[755], line_83[753], line_82[751], line_81[749], line_80[747], line_79[745], line_78[743], line_77[741], line_76[739], line_75[737], line_74[735], line_73[733], line_72[731], line_71[729], line_70[727], line_69[725], line_68[723], line_67[721], line_66[719], line_65[717], line_64[715], line_63[713], line_62[711], line_61[709], line_60[707], line_59[705], line_58[703], line_57[701], line_56[699], line_55[697], line_54[695], line_53[693], line_52[691], line_51[689], line_50[687], line_49[685], line_48[683], line_47[681], line_46[679], line_45[677], line_44[675], line_43[673], line_42[671], line_41[669], line_40[667], line_39[665], line_38[663], line_37[661], line_36[659], line_35[657], line_34[655], line_33[653], line_32[651], line_31[649], line_30[647], line_29[645], line_28[643], line_27[641], line_26[639], line_25[637], line_24[635], line_23[633], line_22[631], line_21[629], line_20[627], line_19[625], line_18[623], line_17[621], line_16[619], line_15[617], line_14[615], line_13[613], line_12[611], line_11[609], line_10[607], line_9[605], line_8[603], line_7[601], line_6[599], line_5[597], line_4[595], line_3[593], line_2[591], line_1[589] };
assign col_844 = {line_128[844], line_127[842], line_126[840], line_125[838], line_124[836], line_123[834], line_122[832], line_121[830], line_120[828], line_119[826], line_118[824], line_117[822], line_116[820], line_115[818], line_114[816], line_113[814], line_112[812], line_111[810], line_110[808], line_109[806], line_108[804], line_107[802], line_106[800], line_105[798], line_104[796], line_103[794], line_102[792], line_101[790], line_100[788], line_99[786], line_98[784], line_97[782], line_96[780], line_95[778], line_94[776], line_93[774], line_92[772], line_91[770], line_90[768], line_89[766], line_88[764], line_87[762], line_86[760], line_85[758], line_84[756], line_83[754], line_82[752], line_81[750], line_80[748], line_79[746], line_78[744], line_77[742], line_76[740], line_75[738], line_74[736], line_73[734], line_72[732], line_71[730], line_70[728], line_69[726], line_68[724], line_67[722], line_66[720], line_65[718], line_64[716], line_63[714], line_62[712], line_61[710], line_60[708], line_59[706], line_58[704], line_57[702], line_56[700], line_55[698], line_54[696], line_53[694], line_52[692], line_51[690], line_50[688], line_49[686], line_48[684], line_47[682], line_46[680], line_45[678], line_44[676], line_43[674], line_42[672], line_41[670], line_40[668], line_39[666], line_38[664], line_37[662], line_36[660], line_35[658], line_34[656], line_33[654], line_32[652], line_31[650], line_30[648], line_29[646], line_28[644], line_27[642], line_26[640], line_25[638], line_24[636], line_23[634], line_22[632], line_21[630], line_20[628], line_19[626], line_18[624], line_17[622], line_16[620], line_15[618], line_14[616], line_13[614], line_12[612], line_11[610], line_10[608], line_9[606], line_8[604], line_7[602], line_6[600], line_5[598], line_4[596], line_3[594], line_2[592], line_1[590] };
assign col_845 = {line_128[845], line_127[843], line_126[841], line_125[839], line_124[837], line_123[835], line_122[833], line_121[831], line_120[829], line_119[827], line_118[825], line_117[823], line_116[821], line_115[819], line_114[817], line_113[815], line_112[813], line_111[811], line_110[809], line_109[807], line_108[805], line_107[803], line_106[801], line_105[799], line_104[797], line_103[795], line_102[793], line_101[791], line_100[789], line_99[787], line_98[785], line_97[783], line_96[781], line_95[779], line_94[777], line_93[775], line_92[773], line_91[771], line_90[769], line_89[767], line_88[765], line_87[763], line_86[761], line_85[759], line_84[757], line_83[755], line_82[753], line_81[751], line_80[749], line_79[747], line_78[745], line_77[743], line_76[741], line_75[739], line_74[737], line_73[735], line_72[733], line_71[731], line_70[729], line_69[727], line_68[725], line_67[723], line_66[721], line_65[719], line_64[717], line_63[715], line_62[713], line_61[711], line_60[709], line_59[707], line_58[705], line_57[703], line_56[701], line_55[699], line_54[697], line_53[695], line_52[693], line_51[691], line_50[689], line_49[687], line_48[685], line_47[683], line_46[681], line_45[679], line_44[677], line_43[675], line_42[673], line_41[671], line_40[669], line_39[667], line_38[665], line_37[663], line_36[661], line_35[659], line_34[657], line_33[655], line_32[653], line_31[651], line_30[649], line_29[647], line_28[645], line_27[643], line_26[641], line_25[639], line_24[637], line_23[635], line_22[633], line_21[631], line_20[629], line_19[627], line_18[625], line_17[623], line_16[621], line_15[619], line_14[617], line_13[615], line_12[613], line_11[611], line_10[609], line_9[607], line_8[605], line_7[603], line_6[601], line_5[599], line_4[597], line_3[595], line_2[593], line_1[591] };
assign col_846 = {line_128[846], line_127[844], line_126[842], line_125[840], line_124[838], line_123[836], line_122[834], line_121[832], line_120[830], line_119[828], line_118[826], line_117[824], line_116[822], line_115[820], line_114[818], line_113[816], line_112[814], line_111[812], line_110[810], line_109[808], line_108[806], line_107[804], line_106[802], line_105[800], line_104[798], line_103[796], line_102[794], line_101[792], line_100[790], line_99[788], line_98[786], line_97[784], line_96[782], line_95[780], line_94[778], line_93[776], line_92[774], line_91[772], line_90[770], line_89[768], line_88[766], line_87[764], line_86[762], line_85[760], line_84[758], line_83[756], line_82[754], line_81[752], line_80[750], line_79[748], line_78[746], line_77[744], line_76[742], line_75[740], line_74[738], line_73[736], line_72[734], line_71[732], line_70[730], line_69[728], line_68[726], line_67[724], line_66[722], line_65[720], line_64[718], line_63[716], line_62[714], line_61[712], line_60[710], line_59[708], line_58[706], line_57[704], line_56[702], line_55[700], line_54[698], line_53[696], line_52[694], line_51[692], line_50[690], line_49[688], line_48[686], line_47[684], line_46[682], line_45[680], line_44[678], line_43[676], line_42[674], line_41[672], line_40[670], line_39[668], line_38[666], line_37[664], line_36[662], line_35[660], line_34[658], line_33[656], line_32[654], line_31[652], line_30[650], line_29[648], line_28[646], line_27[644], line_26[642], line_25[640], line_24[638], line_23[636], line_22[634], line_21[632], line_20[630], line_19[628], line_18[626], line_17[624], line_16[622], line_15[620], line_14[618], line_13[616], line_12[614], line_11[612], line_10[610], line_9[608], line_8[606], line_7[604], line_6[602], line_5[600], line_4[598], line_3[596], line_2[594], line_1[592] };
assign col_847 = {line_128[847], line_127[845], line_126[843], line_125[841], line_124[839], line_123[837], line_122[835], line_121[833], line_120[831], line_119[829], line_118[827], line_117[825], line_116[823], line_115[821], line_114[819], line_113[817], line_112[815], line_111[813], line_110[811], line_109[809], line_108[807], line_107[805], line_106[803], line_105[801], line_104[799], line_103[797], line_102[795], line_101[793], line_100[791], line_99[789], line_98[787], line_97[785], line_96[783], line_95[781], line_94[779], line_93[777], line_92[775], line_91[773], line_90[771], line_89[769], line_88[767], line_87[765], line_86[763], line_85[761], line_84[759], line_83[757], line_82[755], line_81[753], line_80[751], line_79[749], line_78[747], line_77[745], line_76[743], line_75[741], line_74[739], line_73[737], line_72[735], line_71[733], line_70[731], line_69[729], line_68[727], line_67[725], line_66[723], line_65[721], line_64[719], line_63[717], line_62[715], line_61[713], line_60[711], line_59[709], line_58[707], line_57[705], line_56[703], line_55[701], line_54[699], line_53[697], line_52[695], line_51[693], line_50[691], line_49[689], line_48[687], line_47[685], line_46[683], line_45[681], line_44[679], line_43[677], line_42[675], line_41[673], line_40[671], line_39[669], line_38[667], line_37[665], line_36[663], line_35[661], line_34[659], line_33[657], line_32[655], line_31[653], line_30[651], line_29[649], line_28[647], line_27[645], line_26[643], line_25[641], line_24[639], line_23[637], line_22[635], line_21[633], line_20[631], line_19[629], line_18[627], line_17[625], line_16[623], line_15[621], line_14[619], line_13[617], line_12[615], line_11[613], line_10[611], line_9[609], line_8[607], line_7[605], line_6[603], line_5[601], line_4[599], line_3[597], line_2[595], line_1[593] };
assign col_848 = {line_128[848], line_127[846], line_126[844], line_125[842], line_124[840], line_123[838], line_122[836], line_121[834], line_120[832], line_119[830], line_118[828], line_117[826], line_116[824], line_115[822], line_114[820], line_113[818], line_112[816], line_111[814], line_110[812], line_109[810], line_108[808], line_107[806], line_106[804], line_105[802], line_104[800], line_103[798], line_102[796], line_101[794], line_100[792], line_99[790], line_98[788], line_97[786], line_96[784], line_95[782], line_94[780], line_93[778], line_92[776], line_91[774], line_90[772], line_89[770], line_88[768], line_87[766], line_86[764], line_85[762], line_84[760], line_83[758], line_82[756], line_81[754], line_80[752], line_79[750], line_78[748], line_77[746], line_76[744], line_75[742], line_74[740], line_73[738], line_72[736], line_71[734], line_70[732], line_69[730], line_68[728], line_67[726], line_66[724], line_65[722], line_64[720], line_63[718], line_62[716], line_61[714], line_60[712], line_59[710], line_58[708], line_57[706], line_56[704], line_55[702], line_54[700], line_53[698], line_52[696], line_51[694], line_50[692], line_49[690], line_48[688], line_47[686], line_46[684], line_45[682], line_44[680], line_43[678], line_42[676], line_41[674], line_40[672], line_39[670], line_38[668], line_37[666], line_36[664], line_35[662], line_34[660], line_33[658], line_32[656], line_31[654], line_30[652], line_29[650], line_28[648], line_27[646], line_26[644], line_25[642], line_24[640], line_23[638], line_22[636], line_21[634], line_20[632], line_19[630], line_18[628], line_17[626], line_16[624], line_15[622], line_14[620], line_13[618], line_12[616], line_11[614], line_10[612], line_9[610], line_8[608], line_7[606], line_6[604], line_5[602], line_4[600], line_3[598], line_2[596], line_1[594] };
assign col_849 = {line_128[849], line_127[847], line_126[845], line_125[843], line_124[841], line_123[839], line_122[837], line_121[835], line_120[833], line_119[831], line_118[829], line_117[827], line_116[825], line_115[823], line_114[821], line_113[819], line_112[817], line_111[815], line_110[813], line_109[811], line_108[809], line_107[807], line_106[805], line_105[803], line_104[801], line_103[799], line_102[797], line_101[795], line_100[793], line_99[791], line_98[789], line_97[787], line_96[785], line_95[783], line_94[781], line_93[779], line_92[777], line_91[775], line_90[773], line_89[771], line_88[769], line_87[767], line_86[765], line_85[763], line_84[761], line_83[759], line_82[757], line_81[755], line_80[753], line_79[751], line_78[749], line_77[747], line_76[745], line_75[743], line_74[741], line_73[739], line_72[737], line_71[735], line_70[733], line_69[731], line_68[729], line_67[727], line_66[725], line_65[723], line_64[721], line_63[719], line_62[717], line_61[715], line_60[713], line_59[711], line_58[709], line_57[707], line_56[705], line_55[703], line_54[701], line_53[699], line_52[697], line_51[695], line_50[693], line_49[691], line_48[689], line_47[687], line_46[685], line_45[683], line_44[681], line_43[679], line_42[677], line_41[675], line_40[673], line_39[671], line_38[669], line_37[667], line_36[665], line_35[663], line_34[661], line_33[659], line_32[657], line_31[655], line_30[653], line_29[651], line_28[649], line_27[647], line_26[645], line_25[643], line_24[641], line_23[639], line_22[637], line_21[635], line_20[633], line_19[631], line_18[629], line_17[627], line_16[625], line_15[623], line_14[621], line_13[619], line_12[617], line_11[615], line_10[613], line_9[611], line_8[609], line_7[607], line_6[605], line_5[603], line_4[601], line_3[599], line_2[597], line_1[595] };
assign col_850 = {line_128[850], line_127[848], line_126[846], line_125[844], line_124[842], line_123[840], line_122[838], line_121[836], line_120[834], line_119[832], line_118[830], line_117[828], line_116[826], line_115[824], line_114[822], line_113[820], line_112[818], line_111[816], line_110[814], line_109[812], line_108[810], line_107[808], line_106[806], line_105[804], line_104[802], line_103[800], line_102[798], line_101[796], line_100[794], line_99[792], line_98[790], line_97[788], line_96[786], line_95[784], line_94[782], line_93[780], line_92[778], line_91[776], line_90[774], line_89[772], line_88[770], line_87[768], line_86[766], line_85[764], line_84[762], line_83[760], line_82[758], line_81[756], line_80[754], line_79[752], line_78[750], line_77[748], line_76[746], line_75[744], line_74[742], line_73[740], line_72[738], line_71[736], line_70[734], line_69[732], line_68[730], line_67[728], line_66[726], line_65[724], line_64[722], line_63[720], line_62[718], line_61[716], line_60[714], line_59[712], line_58[710], line_57[708], line_56[706], line_55[704], line_54[702], line_53[700], line_52[698], line_51[696], line_50[694], line_49[692], line_48[690], line_47[688], line_46[686], line_45[684], line_44[682], line_43[680], line_42[678], line_41[676], line_40[674], line_39[672], line_38[670], line_37[668], line_36[666], line_35[664], line_34[662], line_33[660], line_32[658], line_31[656], line_30[654], line_29[652], line_28[650], line_27[648], line_26[646], line_25[644], line_24[642], line_23[640], line_22[638], line_21[636], line_20[634], line_19[632], line_18[630], line_17[628], line_16[626], line_15[624], line_14[622], line_13[620], line_12[618], line_11[616], line_10[614], line_9[612], line_8[610], line_7[608], line_6[606], line_5[604], line_4[602], line_3[600], line_2[598], line_1[596] };
assign col_851 = {line_128[851], line_127[849], line_126[847], line_125[845], line_124[843], line_123[841], line_122[839], line_121[837], line_120[835], line_119[833], line_118[831], line_117[829], line_116[827], line_115[825], line_114[823], line_113[821], line_112[819], line_111[817], line_110[815], line_109[813], line_108[811], line_107[809], line_106[807], line_105[805], line_104[803], line_103[801], line_102[799], line_101[797], line_100[795], line_99[793], line_98[791], line_97[789], line_96[787], line_95[785], line_94[783], line_93[781], line_92[779], line_91[777], line_90[775], line_89[773], line_88[771], line_87[769], line_86[767], line_85[765], line_84[763], line_83[761], line_82[759], line_81[757], line_80[755], line_79[753], line_78[751], line_77[749], line_76[747], line_75[745], line_74[743], line_73[741], line_72[739], line_71[737], line_70[735], line_69[733], line_68[731], line_67[729], line_66[727], line_65[725], line_64[723], line_63[721], line_62[719], line_61[717], line_60[715], line_59[713], line_58[711], line_57[709], line_56[707], line_55[705], line_54[703], line_53[701], line_52[699], line_51[697], line_50[695], line_49[693], line_48[691], line_47[689], line_46[687], line_45[685], line_44[683], line_43[681], line_42[679], line_41[677], line_40[675], line_39[673], line_38[671], line_37[669], line_36[667], line_35[665], line_34[663], line_33[661], line_32[659], line_31[657], line_30[655], line_29[653], line_28[651], line_27[649], line_26[647], line_25[645], line_24[643], line_23[641], line_22[639], line_21[637], line_20[635], line_19[633], line_18[631], line_17[629], line_16[627], line_15[625], line_14[623], line_13[621], line_12[619], line_11[617], line_10[615], line_9[613], line_8[611], line_7[609], line_6[607], line_5[605], line_4[603], line_3[601], line_2[599], line_1[597] };
assign col_852 = {line_128[852], line_127[850], line_126[848], line_125[846], line_124[844], line_123[842], line_122[840], line_121[838], line_120[836], line_119[834], line_118[832], line_117[830], line_116[828], line_115[826], line_114[824], line_113[822], line_112[820], line_111[818], line_110[816], line_109[814], line_108[812], line_107[810], line_106[808], line_105[806], line_104[804], line_103[802], line_102[800], line_101[798], line_100[796], line_99[794], line_98[792], line_97[790], line_96[788], line_95[786], line_94[784], line_93[782], line_92[780], line_91[778], line_90[776], line_89[774], line_88[772], line_87[770], line_86[768], line_85[766], line_84[764], line_83[762], line_82[760], line_81[758], line_80[756], line_79[754], line_78[752], line_77[750], line_76[748], line_75[746], line_74[744], line_73[742], line_72[740], line_71[738], line_70[736], line_69[734], line_68[732], line_67[730], line_66[728], line_65[726], line_64[724], line_63[722], line_62[720], line_61[718], line_60[716], line_59[714], line_58[712], line_57[710], line_56[708], line_55[706], line_54[704], line_53[702], line_52[700], line_51[698], line_50[696], line_49[694], line_48[692], line_47[690], line_46[688], line_45[686], line_44[684], line_43[682], line_42[680], line_41[678], line_40[676], line_39[674], line_38[672], line_37[670], line_36[668], line_35[666], line_34[664], line_33[662], line_32[660], line_31[658], line_30[656], line_29[654], line_28[652], line_27[650], line_26[648], line_25[646], line_24[644], line_23[642], line_22[640], line_21[638], line_20[636], line_19[634], line_18[632], line_17[630], line_16[628], line_15[626], line_14[624], line_13[622], line_12[620], line_11[618], line_10[616], line_9[614], line_8[612], line_7[610], line_6[608], line_5[606], line_4[604], line_3[602], line_2[600], line_1[598] };
assign col_853 = {line_128[853], line_127[851], line_126[849], line_125[847], line_124[845], line_123[843], line_122[841], line_121[839], line_120[837], line_119[835], line_118[833], line_117[831], line_116[829], line_115[827], line_114[825], line_113[823], line_112[821], line_111[819], line_110[817], line_109[815], line_108[813], line_107[811], line_106[809], line_105[807], line_104[805], line_103[803], line_102[801], line_101[799], line_100[797], line_99[795], line_98[793], line_97[791], line_96[789], line_95[787], line_94[785], line_93[783], line_92[781], line_91[779], line_90[777], line_89[775], line_88[773], line_87[771], line_86[769], line_85[767], line_84[765], line_83[763], line_82[761], line_81[759], line_80[757], line_79[755], line_78[753], line_77[751], line_76[749], line_75[747], line_74[745], line_73[743], line_72[741], line_71[739], line_70[737], line_69[735], line_68[733], line_67[731], line_66[729], line_65[727], line_64[725], line_63[723], line_62[721], line_61[719], line_60[717], line_59[715], line_58[713], line_57[711], line_56[709], line_55[707], line_54[705], line_53[703], line_52[701], line_51[699], line_50[697], line_49[695], line_48[693], line_47[691], line_46[689], line_45[687], line_44[685], line_43[683], line_42[681], line_41[679], line_40[677], line_39[675], line_38[673], line_37[671], line_36[669], line_35[667], line_34[665], line_33[663], line_32[661], line_31[659], line_30[657], line_29[655], line_28[653], line_27[651], line_26[649], line_25[647], line_24[645], line_23[643], line_22[641], line_21[639], line_20[637], line_19[635], line_18[633], line_17[631], line_16[629], line_15[627], line_14[625], line_13[623], line_12[621], line_11[619], line_10[617], line_9[615], line_8[613], line_7[611], line_6[609], line_5[607], line_4[605], line_3[603], line_2[601], line_1[599] };
assign col_854 = {line_128[854], line_127[852], line_126[850], line_125[848], line_124[846], line_123[844], line_122[842], line_121[840], line_120[838], line_119[836], line_118[834], line_117[832], line_116[830], line_115[828], line_114[826], line_113[824], line_112[822], line_111[820], line_110[818], line_109[816], line_108[814], line_107[812], line_106[810], line_105[808], line_104[806], line_103[804], line_102[802], line_101[800], line_100[798], line_99[796], line_98[794], line_97[792], line_96[790], line_95[788], line_94[786], line_93[784], line_92[782], line_91[780], line_90[778], line_89[776], line_88[774], line_87[772], line_86[770], line_85[768], line_84[766], line_83[764], line_82[762], line_81[760], line_80[758], line_79[756], line_78[754], line_77[752], line_76[750], line_75[748], line_74[746], line_73[744], line_72[742], line_71[740], line_70[738], line_69[736], line_68[734], line_67[732], line_66[730], line_65[728], line_64[726], line_63[724], line_62[722], line_61[720], line_60[718], line_59[716], line_58[714], line_57[712], line_56[710], line_55[708], line_54[706], line_53[704], line_52[702], line_51[700], line_50[698], line_49[696], line_48[694], line_47[692], line_46[690], line_45[688], line_44[686], line_43[684], line_42[682], line_41[680], line_40[678], line_39[676], line_38[674], line_37[672], line_36[670], line_35[668], line_34[666], line_33[664], line_32[662], line_31[660], line_30[658], line_29[656], line_28[654], line_27[652], line_26[650], line_25[648], line_24[646], line_23[644], line_22[642], line_21[640], line_20[638], line_19[636], line_18[634], line_17[632], line_16[630], line_15[628], line_14[626], line_13[624], line_12[622], line_11[620], line_10[618], line_9[616], line_8[614], line_7[612], line_6[610], line_5[608], line_4[606], line_3[604], line_2[602], line_1[600] };
assign col_855 = {line_128[855], line_127[853], line_126[851], line_125[849], line_124[847], line_123[845], line_122[843], line_121[841], line_120[839], line_119[837], line_118[835], line_117[833], line_116[831], line_115[829], line_114[827], line_113[825], line_112[823], line_111[821], line_110[819], line_109[817], line_108[815], line_107[813], line_106[811], line_105[809], line_104[807], line_103[805], line_102[803], line_101[801], line_100[799], line_99[797], line_98[795], line_97[793], line_96[791], line_95[789], line_94[787], line_93[785], line_92[783], line_91[781], line_90[779], line_89[777], line_88[775], line_87[773], line_86[771], line_85[769], line_84[767], line_83[765], line_82[763], line_81[761], line_80[759], line_79[757], line_78[755], line_77[753], line_76[751], line_75[749], line_74[747], line_73[745], line_72[743], line_71[741], line_70[739], line_69[737], line_68[735], line_67[733], line_66[731], line_65[729], line_64[727], line_63[725], line_62[723], line_61[721], line_60[719], line_59[717], line_58[715], line_57[713], line_56[711], line_55[709], line_54[707], line_53[705], line_52[703], line_51[701], line_50[699], line_49[697], line_48[695], line_47[693], line_46[691], line_45[689], line_44[687], line_43[685], line_42[683], line_41[681], line_40[679], line_39[677], line_38[675], line_37[673], line_36[671], line_35[669], line_34[667], line_33[665], line_32[663], line_31[661], line_30[659], line_29[657], line_28[655], line_27[653], line_26[651], line_25[649], line_24[647], line_23[645], line_22[643], line_21[641], line_20[639], line_19[637], line_18[635], line_17[633], line_16[631], line_15[629], line_14[627], line_13[625], line_12[623], line_11[621], line_10[619], line_9[617], line_8[615], line_7[613], line_6[611], line_5[609], line_4[607], line_3[605], line_2[603], line_1[601] };
assign col_856 = {line_128[856], line_127[854], line_126[852], line_125[850], line_124[848], line_123[846], line_122[844], line_121[842], line_120[840], line_119[838], line_118[836], line_117[834], line_116[832], line_115[830], line_114[828], line_113[826], line_112[824], line_111[822], line_110[820], line_109[818], line_108[816], line_107[814], line_106[812], line_105[810], line_104[808], line_103[806], line_102[804], line_101[802], line_100[800], line_99[798], line_98[796], line_97[794], line_96[792], line_95[790], line_94[788], line_93[786], line_92[784], line_91[782], line_90[780], line_89[778], line_88[776], line_87[774], line_86[772], line_85[770], line_84[768], line_83[766], line_82[764], line_81[762], line_80[760], line_79[758], line_78[756], line_77[754], line_76[752], line_75[750], line_74[748], line_73[746], line_72[744], line_71[742], line_70[740], line_69[738], line_68[736], line_67[734], line_66[732], line_65[730], line_64[728], line_63[726], line_62[724], line_61[722], line_60[720], line_59[718], line_58[716], line_57[714], line_56[712], line_55[710], line_54[708], line_53[706], line_52[704], line_51[702], line_50[700], line_49[698], line_48[696], line_47[694], line_46[692], line_45[690], line_44[688], line_43[686], line_42[684], line_41[682], line_40[680], line_39[678], line_38[676], line_37[674], line_36[672], line_35[670], line_34[668], line_33[666], line_32[664], line_31[662], line_30[660], line_29[658], line_28[656], line_27[654], line_26[652], line_25[650], line_24[648], line_23[646], line_22[644], line_21[642], line_20[640], line_19[638], line_18[636], line_17[634], line_16[632], line_15[630], line_14[628], line_13[626], line_12[624], line_11[622], line_10[620], line_9[618], line_8[616], line_7[614], line_6[612], line_5[610], line_4[608], line_3[606], line_2[604], line_1[602] };
assign col_857 = {line_128[857], line_127[855], line_126[853], line_125[851], line_124[849], line_123[847], line_122[845], line_121[843], line_120[841], line_119[839], line_118[837], line_117[835], line_116[833], line_115[831], line_114[829], line_113[827], line_112[825], line_111[823], line_110[821], line_109[819], line_108[817], line_107[815], line_106[813], line_105[811], line_104[809], line_103[807], line_102[805], line_101[803], line_100[801], line_99[799], line_98[797], line_97[795], line_96[793], line_95[791], line_94[789], line_93[787], line_92[785], line_91[783], line_90[781], line_89[779], line_88[777], line_87[775], line_86[773], line_85[771], line_84[769], line_83[767], line_82[765], line_81[763], line_80[761], line_79[759], line_78[757], line_77[755], line_76[753], line_75[751], line_74[749], line_73[747], line_72[745], line_71[743], line_70[741], line_69[739], line_68[737], line_67[735], line_66[733], line_65[731], line_64[729], line_63[727], line_62[725], line_61[723], line_60[721], line_59[719], line_58[717], line_57[715], line_56[713], line_55[711], line_54[709], line_53[707], line_52[705], line_51[703], line_50[701], line_49[699], line_48[697], line_47[695], line_46[693], line_45[691], line_44[689], line_43[687], line_42[685], line_41[683], line_40[681], line_39[679], line_38[677], line_37[675], line_36[673], line_35[671], line_34[669], line_33[667], line_32[665], line_31[663], line_30[661], line_29[659], line_28[657], line_27[655], line_26[653], line_25[651], line_24[649], line_23[647], line_22[645], line_21[643], line_20[641], line_19[639], line_18[637], line_17[635], line_16[633], line_15[631], line_14[629], line_13[627], line_12[625], line_11[623], line_10[621], line_9[619], line_8[617], line_7[615], line_6[613], line_5[611], line_4[609], line_3[607], line_2[605], line_1[603] };
assign col_858 = {line_128[858], line_127[856], line_126[854], line_125[852], line_124[850], line_123[848], line_122[846], line_121[844], line_120[842], line_119[840], line_118[838], line_117[836], line_116[834], line_115[832], line_114[830], line_113[828], line_112[826], line_111[824], line_110[822], line_109[820], line_108[818], line_107[816], line_106[814], line_105[812], line_104[810], line_103[808], line_102[806], line_101[804], line_100[802], line_99[800], line_98[798], line_97[796], line_96[794], line_95[792], line_94[790], line_93[788], line_92[786], line_91[784], line_90[782], line_89[780], line_88[778], line_87[776], line_86[774], line_85[772], line_84[770], line_83[768], line_82[766], line_81[764], line_80[762], line_79[760], line_78[758], line_77[756], line_76[754], line_75[752], line_74[750], line_73[748], line_72[746], line_71[744], line_70[742], line_69[740], line_68[738], line_67[736], line_66[734], line_65[732], line_64[730], line_63[728], line_62[726], line_61[724], line_60[722], line_59[720], line_58[718], line_57[716], line_56[714], line_55[712], line_54[710], line_53[708], line_52[706], line_51[704], line_50[702], line_49[700], line_48[698], line_47[696], line_46[694], line_45[692], line_44[690], line_43[688], line_42[686], line_41[684], line_40[682], line_39[680], line_38[678], line_37[676], line_36[674], line_35[672], line_34[670], line_33[668], line_32[666], line_31[664], line_30[662], line_29[660], line_28[658], line_27[656], line_26[654], line_25[652], line_24[650], line_23[648], line_22[646], line_21[644], line_20[642], line_19[640], line_18[638], line_17[636], line_16[634], line_15[632], line_14[630], line_13[628], line_12[626], line_11[624], line_10[622], line_9[620], line_8[618], line_7[616], line_6[614], line_5[612], line_4[610], line_3[608], line_2[606], line_1[604] };
assign col_859 = {line_128[859], line_127[857], line_126[855], line_125[853], line_124[851], line_123[849], line_122[847], line_121[845], line_120[843], line_119[841], line_118[839], line_117[837], line_116[835], line_115[833], line_114[831], line_113[829], line_112[827], line_111[825], line_110[823], line_109[821], line_108[819], line_107[817], line_106[815], line_105[813], line_104[811], line_103[809], line_102[807], line_101[805], line_100[803], line_99[801], line_98[799], line_97[797], line_96[795], line_95[793], line_94[791], line_93[789], line_92[787], line_91[785], line_90[783], line_89[781], line_88[779], line_87[777], line_86[775], line_85[773], line_84[771], line_83[769], line_82[767], line_81[765], line_80[763], line_79[761], line_78[759], line_77[757], line_76[755], line_75[753], line_74[751], line_73[749], line_72[747], line_71[745], line_70[743], line_69[741], line_68[739], line_67[737], line_66[735], line_65[733], line_64[731], line_63[729], line_62[727], line_61[725], line_60[723], line_59[721], line_58[719], line_57[717], line_56[715], line_55[713], line_54[711], line_53[709], line_52[707], line_51[705], line_50[703], line_49[701], line_48[699], line_47[697], line_46[695], line_45[693], line_44[691], line_43[689], line_42[687], line_41[685], line_40[683], line_39[681], line_38[679], line_37[677], line_36[675], line_35[673], line_34[671], line_33[669], line_32[667], line_31[665], line_30[663], line_29[661], line_28[659], line_27[657], line_26[655], line_25[653], line_24[651], line_23[649], line_22[647], line_21[645], line_20[643], line_19[641], line_18[639], line_17[637], line_16[635], line_15[633], line_14[631], line_13[629], line_12[627], line_11[625], line_10[623], line_9[621], line_8[619], line_7[617], line_6[615], line_5[613], line_4[611], line_3[609], line_2[607], line_1[605] };
assign col_860 = {line_128[860], line_127[858], line_126[856], line_125[854], line_124[852], line_123[850], line_122[848], line_121[846], line_120[844], line_119[842], line_118[840], line_117[838], line_116[836], line_115[834], line_114[832], line_113[830], line_112[828], line_111[826], line_110[824], line_109[822], line_108[820], line_107[818], line_106[816], line_105[814], line_104[812], line_103[810], line_102[808], line_101[806], line_100[804], line_99[802], line_98[800], line_97[798], line_96[796], line_95[794], line_94[792], line_93[790], line_92[788], line_91[786], line_90[784], line_89[782], line_88[780], line_87[778], line_86[776], line_85[774], line_84[772], line_83[770], line_82[768], line_81[766], line_80[764], line_79[762], line_78[760], line_77[758], line_76[756], line_75[754], line_74[752], line_73[750], line_72[748], line_71[746], line_70[744], line_69[742], line_68[740], line_67[738], line_66[736], line_65[734], line_64[732], line_63[730], line_62[728], line_61[726], line_60[724], line_59[722], line_58[720], line_57[718], line_56[716], line_55[714], line_54[712], line_53[710], line_52[708], line_51[706], line_50[704], line_49[702], line_48[700], line_47[698], line_46[696], line_45[694], line_44[692], line_43[690], line_42[688], line_41[686], line_40[684], line_39[682], line_38[680], line_37[678], line_36[676], line_35[674], line_34[672], line_33[670], line_32[668], line_31[666], line_30[664], line_29[662], line_28[660], line_27[658], line_26[656], line_25[654], line_24[652], line_23[650], line_22[648], line_21[646], line_20[644], line_19[642], line_18[640], line_17[638], line_16[636], line_15[634], line_14[632], line_13[630], line_12[628], line_11[626], line_10[624], line_9[622], line_8[620], line_7[618], line_6[616], line_5[614], line_4[612], line_3[610], line_2[608], line_1[606] };
assign col_861 = {line_128[861], line_127[859], line_126[857], line_125[855], line_124[853], line_123[851], line_122[849], line_121[847], line_120[845], line_119[843], line_118[841], line_117[839], line_116[837], line_115[835], line_114[833], line_113[831], line_112[829], line_111[827], line_110[825], line_109[823], line_108[821], line_107[819], line_106[817], line_105[815], line_104[813], line_103[811], line_102[809], line_101[807], line_100[805], line_99[803], line_98[801], line_97[799], line_96[797], line_95[795], line_94[793], line_93[791], line_92[789], line_91[787], line_90[785], line_89[783], line_88[781], line_87[779], line_86[777], line_85[775], line_84[773], line_83[771], line_82[769], line_81[767], line_80[765], line_79[763], line_78[761], line_77[759], line_76[757], line_75[755], line_74[753], line_73[751], line_72[749], line_71[747], line_70[745], line_69[743], line_68[741], line_67[739], line_66[737], line_65[735], line_64[733], line_63[731], line_62[729], line_61[727], line_60[725], line_59[723], line_58[721], line_57[719], line_56[717], line_55[715], line_54[713], line_53[711], line_52[709], line_51[707], line_50[705], line_49[703], line_48[701], line_47[699], line_46[697], line_45[695], line_44[693], line_43[691], line_42[689], line_41[687], line_40[685], line_39[683], line_38[681], line_37[679], line_36[677], line_35[675], line_34[673], line_33[671], line_32[669], line_31[667], line_30[665], line_29[663], line_28[661], line_27[659], line_26[657], line_25[655], line_24[653], line_23[651], line_22[649], line_21[647], line_20[645], line_19[643], line_18[641], line_17[639], line_16[637], line_15[635], line_14[633], line_13[631], line_12[629], line_11[627], line_10[625], line_9[623], line_8[621], line_7[619], line_6[617], line_5[615], line_4[613], line_3[611], line_2[609], line_1[607] };
assign col_862 = {line_128[862], line_127[860], line_126[858], line_125[856], line_124[854], line_123[852], line_122[850], line_121[848], line_120[846], line_119[844], line_118[842], line_117[840], line_116[838], line_115[836], line_114[834], line_113[832], line_112[830], line_111[828], line_110[826], line_109[824], line_108[822], line_107[820], line_106[818], line_105[816], line_104[814], line_103[812], line_102[810], line_101[808], line_100[806], line_99[804], line_98[802], line_97[800], line_96[798], line_95[796], line_94[794], line_93[792], line_92[790], line_91[788], line_90[786], line_89[784], line_88[782], line_87[780], line_86[778], line_85[776], line_84[774], line_83[772], line_82[770], line_81[768], line_80[766], line_79[764], line_78[762], line_77[760], line_76[758], line_75[756], line_74[754], line_73[752], line_72[750], line_71[748], line_70[746], line_69[744], line_68[742], line_67[740], line_66[738], line_65[736], line_64[734], line_63[732], line_62[730], line_61[728], line_60[726], line_59[724], line_58[722], line_57[720], line_56[718], line_55[716], line_54[714], line_53[712], line_52[710], line_51[708], line_50[706], line_49[704], line_48[702], line_47[700], line_46[698], line_45[696], line_44[694], line_43[692], line_42[690], line_41[688], line_40[686], line_39[684], line_38[682], line_37[680], line_36[678], line_35[676], line_34[674], line_33[672], line_32[670], line_31[668], line_30[666], line_29[664], line_28[662], line_27[660], line_26[658], line_25[656], line_24[654], line_23[652], line_22[650], line_21[648], line_20[646], line_19[644], line_18[642], line_17[640], line_16[638], line_15[636], line_14[634], line_13[632], line_12[630], line_11[628], line_10[626], line_9[624], line_8[622], line_7[620], line_6[618], line_5[616], line_4[614], line_3[612], line_2[610], line_1[608] };
assign col_863 = {line_128[863], line_127[861], line_126[859], line_125[857], line_124[855], line_123[853], line_122[851], line_121[849], line_120[847], line_119[845], line_118[843], line_117[841], line_116[839], line_115[837], line_114[835], line_113[833], line_112[831], line_111[829], line_110[827], line_109[825], line_108[823], line_107[821], line_106[819], line_105[817], line_104[815], line_103[813], line_102[811], line_101[809], line_100[807], line_99[805], line_98[803], line_97[801], line_96[799], line_95[797], line_94[795], line_93[793], line_92[791], line_91[789], line_90[787], line_89[785], line_88[783], line_87[781], line_86[779], line_85[777], line_84[775], line_83[773], line_82[771], line_81[769], line_80[767], line_79[765], line_78[763], line_77[761], line_76[759], line_75[757], line_74[755], line_73[753], line_72[751], line_71[749], line_70[747], line_69[745], line_68[743], line_67[741], line_66[739], line_65[737], line_64[735], line_63[733], line_62[731], line_61[729], line_60[727], line_59[725], line_58[723], line_57[721], line_56[719], line_55[717], line_54[715], line_53[713], line_52[711], line_51[709], line_50[707], line_49[705], line_48[703], line_47[701], line_46[699], line_45[697], line_44[695], line_43[693], line_42[691], line_41[689], line_40[687], line_39[685], line_38[683], line_37[681], line_36[679], line_35[677], line_34[675], line_33[673], line_32[671], line_31[669], line_30[667], line_29[665], line_28[663], line_27[661], line_26[659], line_25[657], line_24[655], line_23[653], line_22[651], line_21[649], line_20[647], line_19[645], line_18[643], line_17[641], line_16[639], line_15[637], line_14[635], line_13[633], line_12[631], line_11[629], line_10[627], line_9[625], line_8[623], line_7[621], line_6[619], line_5[617], line_4[615], line_3[613], line_2[611], line_1[609] };
assign col_864 = {line_128[864], line_127[862], line_126[860], line_125[858], line_124[856], line_123[854], line_122[852], line_121[850], line_120[848], line_119[846], line_118[844], line_117[842], line_116[840], line_115[838], line_114[836], line_113[834], line_112[832], line_111[830], line_110[828], line_109[826], line_108[824], line_107[822], line_106[820], line_105[818], line_104[816], line_103[814], line_102[812], line_101[810], line_100[808], line_99[806], line_98[804], line_97[802], line_96[800], line_95[798], line_94[796], line_93[794], line_92[792], line_91[790], line_90[788], line_89[786], line_88[784], line_87[782], line_86[780], line_85[778], line_84[776], line_83[774], line_82[772], line_81[770], line_80[768], line_79[766], line_78[764], line_77[762], line_76[760], line_75[758], line_74[756], line_73[754], line_72[752], line_71[750], line_70[748], line_69[746], line_68[744], line_67[742], line_66[740], line_65[738], line_64[736], line_63[734], line_62[732], line_61[730], line_60[728], line_59[726], line_58[724], line_57[722], line_56[720], line_55[718], line_54[716], line_53[714], line_52[712], line_51[710], line_50[708], line_49[706], line_48[704], line_47[702], line_46[700], line_45[698], line_44[696], line_43[694], line_42[692], line_41[690], line_40[688], line_39[686], line_38[684], line_37[682], line_36[680], line_35[678], line_34[676], line_33[674], line_32[672], line_31[670], line_30[668], line_29[666], line_28[664], line_27[662], line_26[660], line_25[658], line_24[656], line_23[654], line_22[652], line_21[650], line_20[648], line_19[646], line_18[644], line_17[642], line_16[640], line_15[638], line_14[636], line_13[634], line_12[632], line_11[630], line_10[628], line_9[626], line_8[624], line_7[622], line_6[620], line_5[618], line_4[616], line_3[614], line_2[612], line_1[610] };
assign col_865 = {line_128[865], line_127[863], line_126[861], line_125[859], line_124[857], line_123[855], line_122[853], line_121[851], line_120[849], line_119[847], line_118[845], line_117[843], line_116[841], line_115[839], line_114[837], line_113[835], line_112[833], line_111[831], line_110[829], line_109[827], line_108[825], line_107[823], line_106[821], line_105[819], line_104[817], line_103[815], line_102[813], line_101[811], line_100[809], line_99[807], line_98[805], line_97[803], line_96[801], line_95[799], line_94[797], line_93[795], line_92[793], line_91[791], line_90[789], line_89[787], line_88[785], line_87[783], line_86[781], line_85[779], line_84[777], line_83[775], line_82[773], line_81[771], line_80[769], line_79[767], line_78[765], line_77[763], line_76[761], line_75[759], line_74[757], line_73[755], line_72[753], line_71[751], line_70[749], line_69[747], line_68[745], line_67[743], line_66[741], line_65[739], line_64[737], line_63[735], line_62[733], line_61[731], line_60[729], line_59[727], line_58[725], line_57[723], line_56[721], line_55[719], line_54[717], line_53[715], line_52[713], line_51[711], line_50[709], line_49[707], line_48[705], line_47[703], line_46[701], line_45[699], line_44[697], line_43[695], line_42[693], line_41[691], line_40[689], line_39[687], line_38[685], line_37[683], line_36[681], line_35[679], line_34[677], line_33[675], line_32[673], line_31[671], line_30[669], line_29[667], line_28[665], line_27[663], line_26[661], line_25[659], line_24[657], line_23[655], line_22[653], line_21[651], line_20[649], line_19[647], line_18[645], line_17[643], line_16[641], line_15[639], line_14[637], line_13[635], line_12[633], line_11[631], line_10[629], line_9[627], line_8[625], line_7[623], line_6[621], line_5[619], line_4[617], line_3[615], line_2[613], line_1[611] };
assign col_866 = {line_128[866], line_127[864], line_126[862], line_125[860], line_124[858], line_123[856], line_122[854], line_121[852], line_120[850], line_119[848], line_118[846], line_117[844], line_116[842], line_115[840], line_114[838], line_113[836], line_112[834], line_111[832], line_110[830], line_109[828], line_108[826], line_107[824], line_106[822], line_105[820], line_104[818], line_103[816], line_102[814], line_101[812], line_100[810], line_99[808], line_98[806], line_97[804], line_96[802], line_95[800], line_94[798], line_93[796], line_92[794], line_91[792], line_90[790], line_89[788], line_88[786], line_87[784], line_86[782], line_85[780], line_84[778], line_83[776], line_82[774], line_81[772], line_80[770], line_79[768], line_78[766], line_77[764], line_76[762], line_75[760], line_74[758], line_73[756], line_72[754], line_71[752], line_70[750], line_69[748], line_68[746], line_67[744], line_66[742], line_65[740], line_64[738], line_63[736], line_62[734], line_61[732], line_60[730], line_59[728], line_58[726], line_57[724], line_56[722], line_55[720], line_54[718], line_53[716], line_52[714], line_51[712], line_50[710], line_49[708], line_48[706], line_47[704], line_46[702], line_45[700], line_44[698], line_43[696], line_42[694], line_41[692], line_40[690], line_39[688], line_38[686], line_37[684], line_36[682], line_35[680], line_34[678], line_33[676], line_32[674], line_31[672], line_30[670], line_29[668], line_28[666], line_27[664], line_26[662], line_25[660], line_24[658], line_23[656], line_22[654], line_21[652], line_20[650], line_19[648], line_18[646], line_17[644], line_16[642], line_15[640], line_14[638], line_13[636], line_12[634], line_11[632], line_10[630], line_9[628], line_8[626], line_7[624], line_6[622], line_5[620], line_4[618], line_3[616], line_2[614], line_1[612] };
assign col_867 = {line_128[867], line_127[865], line_126[863], line_125[861], line_124[859], line_123[857], line_122[855], line_121[853], line_120[851], line_119[849], line_118[847], line_117[845], line_116[843], line_115[841], line_114[839], line_113[837], line_112[835], line_111[833], line_110[831], line_109[829], line_108[827], line_107[825], line_106[823], line_105[821], line_104[819], line_103[817], line_102[815], line_101[813], line_100[811], line_99[809], line_98[807], line_97[805], line_96[803], line_95[801], line_94[799], line_93[797], line_92[795], line_91[793], line_90[791], line_89[789], line_88[787], line_87[785], line_86[783], line_85[781], line_84[779], line_83[777], line_82[775], line_81[773], line_80[771], line_79[769], line_78[767], line_77[765], line_76[763], line_75[761], line_74[759], line_73[757], line_72[755], line_71[753], line_70[751], line_69[749], line_68[747], line_67[745], line_66[743], line_65[741], line_64[739], line_63[737], line_62[735], line_61[733], line_60[731], line_59[729], line_58[727], line_57[725], line_56[723], line_55[721], line_54[719], line_53[717], line_52[715], line_51[713], line_50[711], line_49[709], line_48[707], line_47[705], line_46[703], line_45[701], line_44[699], line_43[697], line_42[695], line_41[693], line_40[691], line_39[689], line_38[687], line_37[685], line_36[683], line_35[681], line_34[679], line_33[677], line_32[675], line_31[673], line_30[671], line_29[669], line_28[667], line_27[665], line_26[663], line_25[661], line_24[659], line_23[657], line_22[655], line_21[653], line_20[651], line_19[649], line_18[647], line_17[645], line_16[643], line_15[641], line_14[639], line_13[637], line_12[635], line_11[633], line_10[631], line_9[629], line_8[627], line_7[625], line_6[623], line_5[621], line_4[619], line_3[617], line_2[615], line_1[613] };
assign col_868 = {line_128[868], line_127[866], line_126[864], line_125[862], line_124[860], line_123[858], line_122[856], line_121[854], line_120[852], line_119[850], line_118[848], line_117[846], line_116[844], line_115[842], line_114[840], line_113[838], line_112[836], line_111[834], line_110[832], line_109[830], line_108[828], line_107[826], line_106[824], line_105[822], line_104[820], line_103[818], line_102[816], line_101[814], line_100[812], line_99[810], line_98[808], line_97[806], line_96[804], line_95[802], line_94[800], line_93[798], line_92[796], line_91[794], line_90[792], line_89[790], line_88[788], line_87[786], line_86[784], line_85[782], line_84[780], line_83[778], line_82[776], line_81[774], line_80[772], line_79[770], line_78[768], line_77[766], line_76[764], line_75[762], line_74[760], line_73[758], line_72[756], line_71[754], line_70[752], line_69[750], line_68[748], line_67[746], line_66[744], line_65[742], line_64[740], line_63[738], line_62[736], line_61[734], line_60[732], line_59[730], line_58[728], line_57[726], line_56[724], line_55[722], line_54[720], line_53[718], line_52[716], line_51[714], line_50[712], line_49[710], line_48[708], line_47[706], line_46[704], line_45[702], line_44[700], line_43[698], line_42[696], line_41[694], line_40[692], line_39[690], line_38[688], line_37[686], line_36[684], line_35[682], line_34[680], line_33[678], line_32[676], line_31[674], line_30[672], line_29[670], line_28[668], line_27[666], line_26[664], line_25[662], line_24[660], line_23[658], line_22[656], line_21[654], line_20[652], line_19[650], line_18[648], line_17[646], line_16[644], line_15[642], line_14[640], line_13[638], line_12[636], line_11[634], line_10[632], line_9[630], line_8[628], line_7[626], line_6[624], line_5[622], line_4[620], line_3[618], line_2[616], line_1[614] };
assign col_869 = {line_128[869], line_127[867], line_126[865], line_125[863], line_124[861], line_123[859], line_122[857], line_121[855], line_120[853], line_119[851], line_118[849], line_117[847], line_116[845], line_115[843], line_114[841], line_113[839], line_112[837], line_111[835], line_110[833], line_109[831], line_108[829], line_107[827], line_106[825], line_105[823], line_104[821], line_103[819], line_102[817], line_101[815], line_100[813], line_99[811], line_98[809], line_97[807], line_96[805], line_95[803], line_94[801], line_93[799], line_92[797], line_91[795], line_90[793], line_89[791], line_88[789], line_87[787], line_86[785], line_85[783], line_84[781], line_83[779], line_82[777], line_81[775], line_80[773], line_79[771], line_78[769], line_77[767], line_76[765], line_75[763], line_74[761], line_73[759], line_72[757], line_71[755], line_70[753], line_69[751], line_68[749], line_67[747], line_66[745], line_65[743], line_64[741], line_63[739], line_62[737], line_61[735], line_60[733], line_59[731], line_58[729], line_57[727], line_56[725], line_55[723], line_54[721], line_53[719], line_52[717], line_51[715], line_50[713], line_49[711], line_48[709], line_47[707], line_46[705], line_45[703], line_44[701], line_43[699], line_42[697], line_41[695], line_40[693], line_39[691], line_38[689], line_37[687], line_36[685], line_35[683], line_34[681], line_33[679], line_32[677], line_31[675], line_30[673], line_29[671], line_28[669], line_27[667], line_26[665], line_25[663], line_24[661], line_23[659], line_22[657], line_21[655], line_20[653], line_19[651], line_18[649], line_17[647], line_16[645], line_15[643], line_14[641], line_13[639], line_12[637], line_11[635], line_10[633], line_9[631], line_8[629], line_7[627], line_6[625], line_5[623], line_4[621], line_3[619], line_2[617], line_1[615] };
assign col_870 = {line_128[870], line_127[868], line_126[866], line_125[864], line_124[862], line_123[860], line_122[858], line_121[856], line_120[854], line_119[852], line_118[850], line_117[848], line_116[846], line_115[844], line_114[842], line_113[840], line_112[838], line_111[836], line_110[834], line_109[832], line_108[830], line_107[828], line_106[826], line_105[824], line_104[822], line_103[820], line_102[818], line_101[816], line_100[814], line_99[812], line_98[810], line_97[808], line_96[806], line_95[804], line_94[802], line_93[800], line_92[798], line_91[796], line_90[794], line_89[792], line_88[790], line_87[788], line_86[786], line_85[784], line_84[782], line_83[780], line_82[778], line_81[776], line_80[774], line_79[772], line_78[770], line_77[768], line_76[766], line_75[764], line_74[762], line_73[760], line_72[758], line_71[756], line_70[754], line_69[752], line_68[750], line_67[748], line_66[746], line_65[744], line_64[742], line_63[740], line_62[738], line_61[736], line_60[734], line_59[732], line_58[730], line_57[728], line_56[726], line_55[724], line_54[722], line_53[720], line_52[718], line_51[716], line_50[714], line_49[712], line_48[710], line_47[708], line_46[706], line_45[704], line_44[702], line_43[700], line_42[698], line_41[696], line_40[694], line_39[692], line_38[690], line_37[688], line_36[686], line_35[684], line_34[682], line_33[680], line_32[678], line_31[676], line_30[674], line_29[672], line_28[670], line_27[668], line_26[666], line_25[664], line_24[662], line_23[660], line_22[658], line_21[656], line_20[654], line_19[652], line_18[650], line_17[648], line_16[646], line_15[644], line_14[642], line_13[640], line_12[638], line_11[636], line_10[634], line_9[632], line_8[630], line_7[628], line_6[626], line_5[624], line_4[622], line_3[620], line_2[618], line_1[616] };
assign col_871 = {line_128[871], line_127[869], line_126[867], line_125[865], line_124[863], line_123[861], line_122[859], line_121[857], line_120[855], line_119[853], line_118[851], line_117[849], line_116[847], line_115[845], line_114[843], line_113[841], line_112[839], line_111[837], line_110[835], line_109[833], line_108[831], line_107[829], line_106[827], line_105[825], line_104[823], line_103[821], line_102[819], line_101[817], line_100[815], line_99[813], line_98[811], line_97[809], line_96[807], line_95[805], line_94[803], line_93[801], line_92[799], line_91[797], line_90[795], line_89[793], line_88[791], line_87[789], line_86[787], line_85[785], line_84[783], line_83[781], line_82[779], line_81[777], line_80[775], line_79[773], line_78[771], line_77[769], line_76[767], line_75[765], line_74[763], line_73[761], line_72[759], line_71[757], line_70[755], line_69[753], line_68[751], line_67[749], line_66[747], line_65[745], line_64[743], line_63[741], line_62[739], line_61[737], line_60[735], line_59[733], line_58[731], line_57[729], line_56[727], line_55[725], line_54[723], line_53[721], line_52[719], line_51[717], line_50[715], line_49[713], line_48[711], line_47[709], line_46[707], line_45[705], line_44[703], line_43[701], line_42[699], line_41[697], line_40[695], line_39[693], line_38[691], line_37[689], line_36[687], line_35[685], line_34[683], line_33[681], line_32[679], line_31[677], line_30[675], line_29[673], line_28[671], line_27[669], line_26[667], line_25[665], line_24[663], line_23[661], line_22[659], line_21[657], line_20[655], line_19[653], line_18[651], line_17[649], line_16[647], line_15[645], line_14[643], line_13[641], line_12[639], line_11[637], line_10[635], line_9[633], line_8[631], line_7[629], line_6[627], line_5[625], line_4[623], line_3[621], line_2[619], line_1[617] };
assign col_872 = {line_128[872], line_127[870], line_126[868], line_125[866], line_124[864], line_123[862], line_122[860], line_121[858], line_120[856], line_119[854], line_118[852], line_117[850], line_116[848], line_115[846], line_114[844], line_113[842], line_112[840], line_111[838], line_110[836], line_109[834], line_108[832], line_107[830], line_106[828], line_105[826], line_104[824], line_103[822], line_102[820], line_101[818], line_100[816], line_99[814], line_98[812], line_97[810], line_96[808], line_95[806], line_94[804], line_93[802], line_92[800], line_91[798], line_90[796], line_89[794], line_88[792], line_87[790], line_86[788], line_85[786], line_84[784], line_83[782], line_82[780], line_81[778], line_80[776], line_79[774], line_78[772], line_77[770], line_76[768], line_75[766], line_74[764], line_73[762], line_72[760], line_71[758], line_70[756], line_69[754], line_68[752], line_67[750], line_66[748], line_65[746], line_64[744], line_63[742], line_62[740], line_61[738], line_60[736], line_59[734], line_58[732], line_57[730], line_56[728], line_55[726], line_54[724], line_53[722], line_52[720], line_51[718], line_50[716], line_49[714], line_48[712], line_47[710], line_46[708], line_45[706], line_44[704], line_43[702], line_42[700], line_41[698], line_40[696], line_39[694], line_38[692], line_37[690], line_36[688], line_35[686], line_34[684], line_33[682], line_32[680], line_31[678], line_30[676], line_29[674], line_28[672], line_27[670], line_26[668], line_25[666], line_24[664], line_23[662], line_22[660], line_21[658], line_20[656], line_19[654], line_18[652], line_17[650], line_16[648], line_15[646], line_14[644], line_13[642], line_12[640], line_11[638], line_10[636], line_9[634], line_8[632], line_7[630], line_6[628], line_5[626], line_4[624], line_3[622], line_2[620], line_1[618] };
assign col_873 = {line_128[873], line_127[871], line_126[869], line_125[867], line_124[865], line_123[863], line_122[861], line_121[859], line_120[857], line_119[855], line_118[853], line_117[851], line_116[849], line_115[847], line_114[845], line_113[843], line_112[841], line_111[839], line_110[837], line_109[835], line_108[833], line_107[831], line_106[829], line_105[827], line_104[825], line_103[823], line_102[821], line_101[819], line_100[817], line_99[815], line_98[813], line_97[811], line_96[809], line_95[807], line_94[805], line_93[803], line_92[801], line_91[799], line_90[797], line_89[795], line_88[793], line_87[791], line_86[789], line_85[787], line_84[785], line_83[783], line_82[781], line_81[779], line_80[777], line_79[775], line_78[773], line_77[771], line_76[769], line_75[767], line_74[765], line_73[763], line_72[761], line_71[759], line_70[757], line_69[755], line_68[753], line_67[751], line_66[749], line_65[747], line_64[745], line_63[743], line_62[741], line_61[739], line_60[737], line_59[735], line_58[733], line_57[731], line_56[729], line_55[727], line_54[725], line_53[723], line_52[721], line_51[719], line_50[717], line_49[715], line_48[713], line_47[711], line_46[709], line_45[707], line_44[705], line_43[703], line_42[701], line_41[699], line_40[697], line_39[695], line_38[693], line_37[691], line_36[689], line_35[687], line_34[685], line_33[683], line_32[681], line_31[679], line_30[677], line_29[675], line_28[673], line_27[671], line_26[669], line_25[667], line_24[665], line_23[663], line_22[661], line_21[659], line_20[657], line_19[655], line_18[653], line_17[651], line_16[649], line_15[647], line_14[645], line_13[643], line_12[641], line_11[639], line_10[637], line_9[635], line_8[633], line_7[631], line_6[629], line_5[627], line_4[625], line_3[623], line_2[621], line_1[619] };
assign col_874 = {line_128[874], line_127[872], line_126[870], line_125[868], line_124[866], line_123[864], line_122[862], line_121[860], line_120[858], line_119[856], line_118[854], line_117[852], line_116[850], line_115[848], line_114[846], line_113[844], line_112[842], line_111[840], line_110[838], line_109[836], line_108[834], line_107[832], line_106[830], line_105[828], line_104[826], line_103[824], line_102[822], line_101[820], line_100[818], line_99[816], line_98[814], line_97[812], line_96[810], line_95[808], line_94[806], line_93[804], line_92[802], line_91[800], line_90[798], line_89[796], line_88[794], line_87[792], line_86[790], line_85[788], line_84[786], line_83[784], line_82[782], line_81[780], line_80[778], line_79[776], line_78[774], line_77[772], line_76[770], line_75[768], line_74[766], line_73[764], line_72[762], line_71[760], line_70[758], line_69[756], line_68[754], line_67[752], line_66[750], line_65[748], line_64[746], line_63[744], line_62[742], line_61[740], line_60[738], line_59[736], line_58[734], line_57[732], line_56[730], line_55[728], line_54[726], line_53[724], line_52[722], line_51[720], line_50[718], line_49[716], line_48[714], line_47[712], line_46[710], line_45[708], line_44[706], line_43[704], line_42[702], line_41[700], line_40[698], line_39[696], line_38[694], line_37[692], line_36[690], line_35[688], line_34[686], line_33[684], line_32[682], line_31[680], line_30[678], line_29[676], line_28[674], line_27[672], line_26[670], line_25[668], line_24[666], line_23[664], line_22[662], line_21[660], line_20[658], line_19[656], line_18[654], line_17[652], line_16[650], line_15[648], line_14[646], line_13[644], line_12[642], line_11[640], line_10[638], line_9[636], line_8[634], line_7[632], line_6[630], line_5[628], line_4[626], line_3[624], line_2[622], line_1[620] };
assign col_875 = {line_128[875], line_127[873], line_126[871], line_125[869], line_124[867], line_123[865], line_122[863], line_121[861], line_120[859], line_119[857], line_118[855], line_117[853], line_116[851], line_115[849], line_114[847], line_113[845], line_112[843], line_111[841], line_110[839], line_109[837], line_108[835], line_107[833], line_106[831], line_105[829], line_104[827], line_103[825], line_102[823], line_101[821], line_100[819], line_99[817], line_98[815], line_97[813], line_96[811], line_95[809], line_94[807], line_93[805], line_92[803], line_91[801], line_90[799], line_89[797], line_88[795], line_87[793], line_86[791], line_85[789], line_84[787], line_83[785], line_82[783], line_81[781], line_80[779], line_79[777], line_78[775], line_77[773], line_76[771], line_75[769], line_74[767], line_73[765], line_72[763], line_71[761], line_70[759], line_69[757], line_68[755], line_67[753], line_66[751], line_65[749], line_64[747], line_63[745], line_62[743], line_61[741], line_60[739], line_59[737], line_58[735], line_57[733], line_56[731], line_55[729], line_54[727], line_53[725], line_52[723], line_51[721], line_50[719], line_49[717], line_48[715], line_47[713], line_46[711], line_45[709], line_44[707], line_43[705], line_42[703], line_41[701], line_40[699], line_39[697], line_38[695], line_37[693], line_36[691], line_35[689], line_34[687], line_33[685], line_32[683], line_31[681], line_30[679], line_29[677], line_28[675], line_27[673], line_26[671], line_25[669], line_24[667], line_23[665], line_22[663], line_21[661], line_20[659], line_19[657], line_18[655], line_17[653], line_16[651], line_15[649], line_14[647], line_13[645], line_12[643], line_11[641], line_10[639], line_9[637], line_8[635], line_7[633], line_6[631], line_5[629], line_4[627], line_3[625], line_2[623], line_1[621] };
assign col_876 = {line_128[876], line_127[874], line_126[872], line_125[870], line_124[868], line_123[866], line_122[864], line_121[862], line_120[860], line_119[858], line_118[856], line_117[854], line_116[852], line_115[850], line_114[848], line_113[846], line_112[844], line_111[842], line_110[840], line_109[838], line_108[836], line_107[834], line_106[832], line_105[830], line_104[828], line_103[826], line_102[824], line_101[822], line_100[820], line_99[818], line_98[816], line_97[814], line_96[812], line_95[810], line_94[808], line_93[806], line_92[804], line_91[802], line_90[800], line_89[798], line_88[796], line_87[794], line_86[792], line_85[790], line_84[788], line_83[786], line_82[784], line_81[782], line_80[780], line_79[778], line_78[776], line_77[774], line_76[772], line_75[770], line_74[768], line_73[766], line_72[764], line_71[762], line_70[760], line_69[758], line_68[756], line_67[754], line_66[752], line_65[750], line_64[748], line_63[746], line_62[744], line_61[742], line_60[740], line_59[738], line_58[736], line_57[734], line_56[732], line_55[730], line_54[728], line_53[726], line_52[724], line_51[722], line_50[720], line_49[718], line_48[716], line_47[714], line_46[712], line_45[710], line_44[708], line_43[706], line_42[704], line_41[702], line_40[700], line_39[698], line_38[696], line_37[694], line_36[692], line_35[690], line_34[688], line_33[686], line_32[684], line_31[682], line_30[680], line_29[678], line_28[676], line_27[674], line_26[672], line_25[670], line_24[668], line_23[666], line_22[664], line_21[662], line_20[660], line_19[658], line_18[656], line_17[654], line_16[652], line_15[650], line_14[648], line_13[646], line_12[644], line_11[642], line_10[640], line_9[638], line_8[636], line_7[634], line_6[632], line_5[630], line_4[628], line_3[626], line_2[624], line_1[622] };
assign col_877 = {line_128[877], line_127[875], line_126[873], line_125[871], line_124[869], line_123[867], line_122[865], line_121[863], line_120[861], line_119[859], line_118[857], line_117[855], line_116[853], line_115[851], line_114[849], line_113[847], line_112[845], line_111[843], line_110[841], line_109[839], line_108[837], line_107[835], line_106[833], line_105[831], line_104[829], line_103[827], line_102[825], line_101[823], line_100[821], line_99[819], line_98[817], line_97[815], line_96[813], line_95[811], line_94[809], line_93[807], line_92[805], line_91[803], line_90[801], line_89[799], line_88[797], line_87[795], line_86[793], line_85[791], line_84[789], line_83[787], line_82[785], line_81[783], line_80[781], line_79[779], line_78[777], line_77[775], line_76[773], line_75[771], line_74[769], line_73[767], line_72[765], line_71[763], line_70[761], line_69[759], line_68[757], line_67[755], line_66[753], line_65[751], line_64[749], line_63[747], line_62[745], line_61[743], line_60[741], line_59[739], line_58[737], line_57[735], line_56[733], line_55[731], line_54[729], line_53[727], line_52[725], line_51[723], line_50[721], line_49[719], line_48[717], line_47[715], line_46[713], line_45[711], line_44[709], line_43[707], line_42[705], line_41[703], line_40[701], line_39[699], line_38[697], line_37[695], line_36[693], line_35[691], line_34[689], line_33[687], line_32[685], line_31[683], line_30[681], line_29[679], line_28[677], line_27[675], line_26[673], line_25[671], line_24[669], line_23[667], line_22[665], line_21[663], line_20[661], line_19[659], line_18[657], line_17[655], line_16[653], line_15[651], line_14[649], line_13[647], line_12[645], line_11[643], line_10[641], line_9[639], line_8[637], line_7[635], line_6[633], line_5[631], line_4[629], line_3[627], line_2[625], line_1[623] };
assign col_878 = {line_128[878], line_127[876], line_126[874], line_125[872], line_124[870], line_123[868], line_122[866], line_121[864], line_120[862], line_119[860], line_118[858], line_117[856], line_116[854], line_115[852], line_114[850], line_113[848], line_112[846], line_111[844], line_110[842], line_109[840], line_108[838], line_107[836], line_106[834], line_105[832], line_104[830], line_103[828], line_102[826], line_101[824], line_100[822], line_99[820], line_98[818], line_97[816], line_96[814], line_95[812], line_94[810], line_93[808], line_92[806], line_91[804], line_90[802], line_89[800], line_88[798], line_87[796], line_86[794], line_85[792], line_84[790], line_83[788], line_82[786], line_81[784], line_80[782], line_79[780], line_78[778], line_77[776], line_76[774], line_75[772], line_74[770], line_73[768], line_72[766], line_71[764], line_70[762], line_69[760], line_68[758], line_67[756], line_66[754], line_65[752], line_64[750], line_63[748], line_62[746], line_61[744], line_60[742], line_59[740], line_58[738], line_57[736], line_56[734], line_55[732], line_54[730], line_53[728], line_52[726], line_51[724], line_50[722], line_49[720], line_48[718], line_47[716], line_46[714], line_45[712], line_44[710], line_43[708], line_42[706], line_41[704], line_40[702], line_39[700], line_38[698], line_37[696], line_36[694], line_35[692], line_34[690], line_33[688], line_32[686], line_31[684], line_30[682], line_29[680], line_28[678], line_27[676], line_26[674], line_25[672], line_24[670], line_23[668], line_22[666], line_21[664], line_20[662], line_19[660], line_18[658], line_17[656], line_16[654], line_15[652], line_14[650], line_13[648], line_12[646], line_11[644], line_10[642], line_9[640], line_8[638], line_7[636], line_6[634], line_5[632], line_4[630], line_3[628], line_2[626], line_1[624] };
assign col_879 = {line_128[879], line_127[877], line_126[875], line_125[873], line_124[871], line_123[869], line_122[867], line_121[865], line_120[863], line_119[861], line_118[859], line_117[857], line_116[855], line_115[853], line_114[851], line_113[849], line_112[847], line_111[845], line_110[843], line_109[841], line_108[839], line_107[837], line_106[835], line_105[833], line_104[831], line_103[829], line_102[827], line_101[825], line_100[823], line_99[821], line_98[819], line_97[817], line_96[815], line_95[813], line_94[811], line_93[809], line_92[807], line_91[805], line_90[803], line_89[801], line_88[799], line_87[797], line_86[795], line_85[793], line_84[791], line_83[789], line_82[787], line_81[785], line_80[783], line_79[781], line_78[779], line_77[777], line_76[775], line_75[773], line_74[771], line_73[769], line_72[767], line_71[765], line_70[763], line_69[761], line_68[759], line_67[757], line_66[755], line_65[753], line_64[751], line_63[749], line_62[747], line_61[745], line_60[743], line_59[741], line_58[739], line_57[737], line_56[735], line_55[733], line_54[731], line_53[729], line_52[727], line_51[725], line_50[723], line_49[721], line_48[719], line_47[717], line_46[715], line_45[713], line_44[711], line_43[709], line_42[707], line_41[705], line_40[703], line_39[701], line_38[699], line_37[697], line_36[695], line_35[693], line_34[691], line_33[689], line_32[687], line_31[685], line_30[683], line_29[681], line_28[679], line_27[677], line_26[675], line_25[673], line_24[671], line_23[669], line_22[667], line_21[665], line_20[663], line_19[661], line_18[659], line_17[657], line_16[655], line_15[653], line_14[651], line_13[649], line_12[647], line_11[645], line_10[643], line_9[641], line_8[639], line_7[637], line_6[635], line_5[633], line_4[631], line_3[629], line_2[627], line_1[625] };
assign col_880 = {line_128[880], line_127[878], line_126[876], line_125[874], line_124[872], line_123[870], line_122[868], line_121[866], line_120[864], line_119[862], line_118[860], line_117[858], line_116[856], line_115[854], line_114[852], line_113[850], line_112[848], line_111[846], line_110[844], line_109[842], line_108[840], line_107[838], line_106[836], line_105[834], line_104[832], line_103[830], line_102[828], line_101[826], line_100[824], line_99[822], line_98[820], line_97[818], line_96[816], line_95[814], line_94[812], line_93[810], line_92[808], line_91[806], line_90[804], line_89[802], line_88[800], line_87[798], line_86[796], line_85[794], line_84[792], line_83[790], line_82[788], line_81[786], line_80[784], line_79[782], line_78[780], line_77[778], line_76[776], line_75[774], line_74[772], line_73[770], line_72[768], line_71[766], line_70[764], line_69[762], line_68[760], line_67[758], line_66[756], line_65[754], line_64[752], line_63[750], line_62[748], line_61[746], line_60[744], line_59[742], line_58[740], line_57[738], line_56[736], line_55[734], line_54[732], line_53[730], line_52[728], line_51[726], line_50[724], line_49[722], line_48[720], line_47[718], line_46[716], line_45[714], line_44[712], line_43[710], line_42[708], line_41[706], line_40[704], line_39[702], line_38[700], line_37[698], line_36[696], line_35[694], line_34[692], line_33[690], line_32[688], line_31[686], line_30[684], line_29[682], line_28[680], line_27[678], line_26[676], line_25[674], line_24[672], line_23[670], line_22[668], line_21[666], line_20[664], line_19[662], line_18[660], line_17[658], line_16[656], line_15[654], line_14[652], line_13[650], line_12[648], line_11[646], line_10[644], line_9[642], line_8[640], line_7[638], line_6[636], line_5[634], line_4[632], line_3[630], line_2[628], line_1[626] };
assign col_881 = {line_128[881], line_127[879], line_126[877], line_125[875], line_124[873], line_123[871], line_122[869], line_121[867], line_120[865], line_119[863], line_118[861], line_117[859], line_116[857], line_115[855], line_114[853], line_113[851], line_112[849], line_111[847], line_110[845], line_109[843], line_108[841], line_107[839], line_106[837], line_105[835], line_104[833], line_103[831], line_102[829], line_101[827], line_100[825], line_99[823], line_98[821], line_97[819], line_96[817], line_95[815], line_94[813], line_93[811], line_92[809], line_91[807], line_90[805], line_89[803], line_88[801], line_87[799], line_86[797], line_85[795], line_84[793], line_83[791], line_82[789], line_81[787], line_80[785], line_79[783], line_78[781], line_77[779], line_76[777], line_75[775], line_74[773], line_73[771], line_72[769], line_71[767], line_70[765], line_69[763], line_68[761], line_67[759], line_66[757], line_65[755], line_64[753], line_63[751], line_62[749], line_61[747], line_60[745], line_59[743], line_58[741], line_57[739], line_56[737], line_55[735], line_54[733], line_53[731], line_52[729], line_51[727], line_50[725], line_49[723], line_48[721], line_47[719], line_46[717], line_45[715], line_44[713], line_43[711], line_42[709], line_41[707], line_40[705], line_39[703], line_38[701], line_37[699], line_36[697], line_35[695], line_34[693], line_33[691], line_32[689], line_31[687], line_30[685], line_29[683], line_28[681], line_27[679], line_26[677], line_25[675], line_24[673], line_23[671], line_22[669], line_21[667], line_20[665], line_19[663], line_18[661], line_17[659], line_16[657], line_15[655], line_14[653], line_13[651], line_12[649], line_11[647], line_10[645], line_9[643], line_8[641], line_7[639], line_6[637], line_5[635], line_4[633], line_3[631], line_2[629], line_1[627] };
assign col_882 = {line_128[882], line_127[880], line_126[878], line_125[876], line_124[874], line_123[872], line_122[870], line_121[868], line_120[866], line_119[864], line_118[862], line_117[860], line_116[858], line_115[856], line_114[854], line_113[852], line_112[850], line_111[848], line_110[846], line_109[844], line_108[842], line_107[840], line_106[838], line_105[836], line_104[834], line_103[832], line_102[830], line_101[828], line_100[826], line_99[824], line_98[822], line_97[820], line_96[818], line_95[816], line_94[814], line_93[812], line_92[810], line_91[808], line_90[806], line_89[804], line_88[802], line_87[800], line_86[798], line_85[796], line_84[794], line_83[792], line_82[790], line_81[788], line_80[786], line_79[784], line_78[782], line_77[780], line_76[778], line_75[776], line_74[774], line_73[772], line_72[770], line_71[768], line_70[766], line_69[764], line_68[762], line_67[760], line_66[758], line_65[756], line_64[754], line_63[752], line_62[750], line_61[748], line_60[746], line_59[744], line_58[742], line_57[740], line_56[738], line_55[736], line_54[734], line_53[732], line_52[730], line_51[728], line_50[726], line_49[724], line_48[722], line_47[720], line_46[718], line_45[716], line_44[714], line_43[712], line_42[710], line_41[708], line_40[706], line_39[704], line_38[702], line_37[700], line_36[698], line_35[696], line_34[694], line_33[692], line_32[690], line_31[688], line_30[686], line_29[684], line_28[682], line_27[680], line_26[678], line_25[676], line_24[674], line_23[672], line_22[670], line_21[668], line_20[666], line_19[664], line_18[662], line_17[660], line_16[658], line_15[656], line_14[654], line_13[652], line_12[650], line_11[648], line_10[646], line_9[644], line_8[642], line_7[640], line_6[638], line_5[636], line_4[634], line_3[632], line_2[630], line_1[628] };
assign col_883 = {line_128[883], line_127[881], line_126[879], line_125[877], line_124[875], line_123[873], line_122[871], line_121[869], line_120[867], line_119[865], line_118[863], line_117[861], line_116[859], line_115[857], line_114[855], line_113[853], line_112[851], line_111[849], line_110[847], line_109[845], line_108[843], line_107[841], line_106[839], line_105[837], line_104[835], line_103[833], line_102[831], line_101[829], line_100[827], line_99[825], line_98[823], line_97[821], line_96[819], line_95[817], line_94[815], line_93[813], line_92[811], line_91[809], line_90[807], line_89[805], line_88[803], line_87[801], line_86[799], line_85[797], line_84[795], line_83[793], line_82[791], line_81[789], line_80[787], line_79[785], line_78[783], line_77[781], line_76[779], line_75[777], line_74[775], line_73[773], line_72[771], line_71[769], line_70[767], line_69[765], line_68[763], line_67[761], line_66[759], line_65[757], line_64[755], line_63[753], line_62[751], line_61[749], line_60[747], line_59[745], line_58[743], line_57[741], line_56[739], line_55[737], line_54[735], line_53[733], line_52[731], line_51[729], line_50[727], line_49[725], line_48[723], line_47[721], line_46[719], line_45[717], line_44[715], line_43[713], line_42[711], line_41[709], line_40[707], line_39[705], line_38[703], line_37[701], line_36[699], line_35[697], line_34[695], line_33[693], line_32[691], line_31[689], line_30[687], line_29[685], line_28[683], line_27[681], line_26[679], line_25[677], line_24[675], line_23[673], line_22[671], line_21[669], line_20[667], line_19[665], line_18[663], line_17[661], line_16[659], line_15[657], line_14[655], line_13[653], line_12[651], line_11[649], line_10[647], line_9[645], line_8[643], line_7[641], line_6[639], line_5[637], line_4[635], line_3[633], line_2[631], line_1[629] };
assign col_884 = {line_128[884], line_127[882], line_126[880], line_125[878], line_124[876], line_123[874], line_122[872], line_121[870], line_120[868], line_119[866], line_118[864], line_117[862], line_116[860], line_115[858], line_114[856], line_113[854], line_112[852], line_111[850], line_110[848], line_109[846], line_108[844], line_107[842], line_106[840], line_105[838], line_104[836], line_103[834], line_102[832], line_101[830], line_100[828], line_99[826], line_98[824], line_97[822], line_96[820], line_95[818], line_94[816], line_93[814], line_92[812], line_91[810], line_90[808], line_89[806], line_88[804], line_87[802], line_86[800], line_85[798], line_84[796], line_83[794], line_82[792], line_81[790], line_80[788], line_79[786], line_78[784], line_77[782], line_76[780], line_75[778], line_74[776], line_73[774], line_72[772], line_71[770], line_70[768], line_69[766], line_68[764], line_67[762], line_66[760], line_65[758], line_64[756], line_63[754], line_62[752], line_61[750], line_60[748], line_59[746], line_58[744], line_57[742], line_56[740], line_55[738], line_54[736], line_53[734], line_52[732], line_51[730], line_50[728], line_49[726], line_48[724], line_47[722], line_46[720], line_45[718], line_44[716], line_43[714], line_42[712], line_41[710], line_40[708], line_39[706], line_38[704], line_37[702], line_36[700], line_35[698], line_34[696], line_33[694], line_32[692], line_31[690], line_30[688], line_29[686], line_28[684], line_27[682], line_26[680], line_25[678], line_24[676], line_23[674], line_22[672], line_21[670], line_20[668], line_19[666], line_18[664], line_17[662], line_16[660], line_15[658], line_14[656], line_13[654], line_12[652], line_11[650], line_10[648], line_9[646], line_8[644], line_7[642], line_6[640], line_5[638], line_4[636], line_3[634], line_2[632], line_1[630] };
assign col_885 = {line_128[885], line_127[883], line_126[881], line_125[879], line_124[877], line_123[875], line_122[873], line_121[871], line_120[869], line_119[867], line_118[865], line_117[863], line_116[861], line_115[859], line_114[857], line_113[855], line_112[853], line_111[851], line_110[849], line_109[847], line_108[845], line_107[843], line_106[841], line_105[839], line_104[837], line_103[835], line_102[833], line_101[831], line_100[829], line_99[827], line_98[825], line_97[823], line_96[821], line_95[819], line_94[817], line_93[815], line_92[813], line_91[811], line_90[809], line_89[807], line_88[805], line_87[803], line_86[801], line_85[799], line_84[797], line_83[795], line_82[793], line_81[791], line_80[789], line_79[787], line_78[785], line_77[783], line_76[781], line_75[779], line_74[777], line_73[775], line_72[773], line_71[771], line_70[769], line_69[767], line_68[765], line_67[763], line_66[761], line_65[759], line_64[757], line_63[755], line_62[753], line_61[751], line_60[749], line_59[747], line_58[745], line_57[743], line_56[741], line_55[739], line_54[737], line_53[735], line_52[733], line_51[731], line_50[729], line_49[727], line_48[725], line_47[723], line_46[721], line_45[719], line_44[717], line_43[715], line_42[713], line_41[711], line_40[709], line_39[707], line_38[705], line_37[703], line_36[701], line_35[699], line_34[697], line_33[695], line_32[693], line_31[691], line_30[689], line_29[687], line_28[685], line_27[683], line_26[681], line_25[679], line_24[677], line_23[675], line_22[673], line_21[671], line_20[669], line_19[667], line_18[665], line_17[663], line_16[661], line_15[659], line_14[657], line_13[655], line_12[653], line_11[651], line_10[649], line_9[647], line_8[645], line_7[643], line_6[641], line_5[639], line_4[637], line_3[635], line_2[633], line_1[631] };
assign col_886 = {line_128[886], line_127[884], line_126[882], line_125[880], line_124[878], line_123[876], line_122[874], line_121[872], line_120[870], line_119[868], line_118[866], line_117[864], line_116[862], line_115[860], line_114[858], line_113[856], line_112[854], line_111[852], line_110[850], line_109[848], line_108[846], line_107[844], line_106[842], line_105[840], line_104[838], line_103[836], line_102[834], line_101[832], line_100[830], line_99[828], line_98[826], line_97[824], line_96[822], line_95[820], line_94[818], line_93[816], line_92[814], line_91[812], line_90[810], line_89[808], line_88[806], line_87[804], line_86[802], line_85[800], line_84[798], line_83[796], line_82[794], line_81[792], line_80[790], line_79[788], line_78[786], line_77[784], line_76[782], line_75[780], line_74[778], line_73[776], line_72[774], line_71[772], line_70[770], line_69[768], line_68[766], line_67[764], line_66[762], line_65[760], line_64[758], line_63[756], line_62[754], line_61[752], line_60[750], line_59[748], line_58[746], line_57[744], line_56[742], line_55[740], line_54[738], line_53[736], line_52[734], line_51[732], line_50[730], line_49[728], line_48[726], line_47[724], line_46[722], line_45[720], line_44[718], line_43[716], line_42[714], line_41[712], line_40[710], line_39[708], line_38[706], line_37[704], line_36[702], line_35[700], line_34[698], line_33[696], line_32[694], line_31[692], line_30[690], line_29[688], line_28[686], line_27[684], line_26[682], line_25[680], line_24[678], line_23[676], line_22[674], line_21[672], line_20[670], line_19[668], line_18[666], line_17[664], line_16[662], line_15[660], line_14[658], line_13[656], line_12[654], line_11[652], line_10[650], line_9[648], line_8[646], line_7[644], line_6[642], line_5[640], line_4[638], line_3[636], line_2[634], line_1[632] };
assign col_887 = {line_128[887], line_127[885], line_126[883], line_125[881], line_124[879], line_123[877], line_122[875], line_121[873], line_120[871], line_119[869], line_118[867], line_117[865], line_116[863], line_115[861], line_114[859], line_113[857], line_112[855], line_111[853], line_110[851], line_109[849], line_108[847], line_107[845], line_106[843], line_105[841], line_104[839], line_103[837], line_102[835], line_101[833], line_100[831], line_99[829], line_98[827], line_97[825], line_96[823], line_95[821], line_94[819], line_93[817], line_92[815], line_91[813], line_90[811], line_89[809], line_88[807], line_87[805], line_86[803], line_85[801], line_84[799], line_83[797], line_82[795], line_81[793], line_80[791], line_79[789], line_78[787], line_77[785], line_76[783], line_75[781], line_74[779], line_73[777], line_72[775], line_71[773], line_70[771], line_69[769], line_68[767], line_67[765], line_66[763], line_65[761], line_64[759], line_63[757], line_62[755], line_61[753], line_60[751], line_59[749], line_58[747], line_57[745], line_56[743], line_55[741], line_54[739], line_53[737], line_52[735], line_51[733], line_50[731], line_49[729], line_48[727], line_47[725], line_46[723], line_45[721], line_44[719], line_43[717], line_42[715], line_41[713], line_40[711], line_39[709], line_38[707], line_37[705], line_36[703], line_35[701], line_34[699], line_33[697], line_32[695], line_31[693], line_30[691], line_29[689], line_28[687], line_27[685], line_26[683], line_25[681], line_24[679], line_23[677], line_22[675], line_21[673], line_20[671], line_19[669], line_18[667], line_17[665], line_16[663], line_15[661], line_14[659], line_13[657], line_12[655], line_11[653], line_10[651], line_9[649], line_8[647], line_7[645], line_6[643], line_5[641], line_4[639], line_3[637], line_2[635], line_1[633] };
assign col_888 = {line_128[888], line_127[886], line_126[884], line_125[882], line_124[880], line_123[878], line_122[876], line_121[874], line_120[872], line_119[870], line_118[868], line_117[866], line_116[864], line_115[862], line_114[860], line_113[858], line_112[856], line_111[854], line_110[852], line_109[850], line_108[848], line_107[846], line_106[844], line_105[842], line_104[840], line_103[838], line_102[836], line_101[834], line_100[832], line_99[830], line_98[828], line_97[826], line_96[824], line_95[822], line_94[820], line_93[818], line_92[816], line_91[814], line_90[812], line_89[810], line_88[808], line_87[806], line_86[804], line_85[802], line_84[800], line_83[798], line_82[796], line_81[794], line_80[792], line_79[790], line_78[788], line_77[786], line_76[784], line_75[782], line_74[780], line_73[778], line_72[776], line_71[774], line_70[772], line_69[770], line_68[768], line_67[766], line_66[764], line_65[762], line_64[760], line_63[758], line_62[756], line_61[754], line_60[752], line_59[750], line_58[748], line_57[746], line_56[744], line_55[742], line_54[740], line_53[738], line_52[736], line_51[734], line_50[732], line_49[730], line_48[728], line_47[726], line_46[724], line_45[722], line_44[720], line_43[718], line_42[716], line_41[714], line_40[712], line_39[710], line_38[708], line_37[706], line_36[704], line_35[702], line_34[700], line_33[698], line_32[696], line_31[694], line_30[692], line_29[690], line_28[688], line_27[686], line_26[684], line_25[682], line_24[680], line_23[678], line_22[676], line_21[674], line_20[672], line_19[670], line_18[668], line_17[666], line_16[664], line_15[662], line_14[660], line_13[658], line_12[656], line_11[654], line_10[652], line_9[650], line_8[648], line_7[646], line_6[644], line_5[642], line_4[640], line_3[638], line_2[636], line_1[634] };
assign col_889 = {line_128[889], line_127[887], line_126[885], line_125[883], line_124[881], line_123[879], line_122[877], line_121[875], line_120[873], line_119[871], line_118[869], line_117[867], line_116[865], line_115[863], line_114[861], line_113[859], line_112[857], line_111[855], line_110[853], line_109[851], line_108[849], line_107[847], line_106[845], line_105[843], line_104[841], line_103[839], line_102[837], line_101[835], line_100[833], line_99[831], line_98[829], line_97[827], line_96[825], line_95[823], line_94[821], line_93[819], line_92[817], line_91[815], line_90[813], line_89[811], line_88[809], line_87[807], line_86[805], line_85[803], line_84[801], line_83[799], line_82[797], line_81[795], line_80[793], line_79[791], line_78[789], line_77[787], line_76[785], line_75[783], line_74[781], line_73[779], line_72[777], line_71[775], line_70[773], line_69[771], line_68[769], line_67[767], line_66[765], line_65[763], line_64[761], line_63[759], line_62[757], line_61[755], line_60[753], line_59[751], line_58[749], line_57[747], line_56[745], line_55[743], line_54[741], line_53[739], line_52[737], line_51[735], line_50[733], line_49[731], line_48[729], line_47[727], line_46[725], line_45[723], line_44[721], line_43[719], line_42[717], line_41[715], line_40[713], line_39[711], line_38[709], line_37[707], line_36[705], line_35[703], line_34[701], line_33[699], line_32[697], line_31[695], line_30[693], line_29[691], line_28[689], line_27[687], line_26[685], line_25[683], line_24[681], line_23[679], line_22[677], line_21[675], line_20[673], line_19[671], line_18[669], line_17[667], line_16[665], line_15[663], line_14[661], line_13[659], line_12[657], line_11[655], line_10[653], line_9[651], line_8[649], line_7[647], line_6[645], line_5[643], line_4[641], line_3[639], line_2[637], line_1[635] };
assign col_890 = {line_128[890], line_127[888], line_126[886], line_125[884], line_124[882], line_123[880], line_122[878], line_121[876], line_120[874], line_119[872], line_118[870], line_117[868], line_116[866], line_115[864], line_114[862], line_113[860], line_112[858], line_111[856], line_110[854], line_109[852], line_108[850], line_107[848], line_106[846], line_105[844], line_104[842], line_103[840], line_102[838], line_101[836], line_100[834], line_99[832], line_98[830], line_97[828], line_96[826], line_95[824], line_94[822], line_93[820], line_92[818], line_91[816], line_90[814], line_89[812], line_88[810], line_87[808], line_86[806], line_85[804], line_84[802], line_83[800], line_82[798], line_81[796], line_80[794], line_79[792], line_78[790], line_77[788], line_76[786], line_75[784], line_74[782], line_73[780], line_72[778], line_71[776], line_70[774], line_69[772], line_68[770], line_67[768], line_66[766], line_65[764], line_64[762], line_63[760], line_62[758], line_61[756], line_60[754], line_59[752], line_58[750], line_57[748], line_56[746], line_55[744], line_54[742], line_53[740], line_52[738], line_51[736], line_50[734], line_49[732], line_48[730], line_47[728], line_46[726], line_45[724], line_44[722], line_43[720], line_42[718], line_41[716], line_40[714], line_39[712], line_38[710], line_37[708], line_36[706], line_35[704], line_34[702], line_33[700], line_32[698], line_31[696], line_30[694], line_29[692], line_28[690], line_27[688], line_26[686], line_25[684], line_24[682], line_23[680], line_22[678], line_21[676], line_20[674], line_19[672], line_18[670], line_17[668], line_16[666], line_15[664], line_14[662], line_13[660], line_12[658], line_11[656], line_10[654], line_9[652], line_8[650], line_7[648], line_6[646], line_5[644], line_4[642], line_3[640], line_2[638], line_1[636] };
assign col_891 = {line_128[891], line_127[889], line_126[887], line_125[885], line_124[883], line_123[881], line_122[879], line_121[877], line_120[875], line_119[873], line_118[871], line_117[869], line_116[867], line_115[865], line_114[863], line_113[861], line_112[859], line_111[857], line_110[855], line_109[853], line_108[851], line_107[849], line_106[847], line_105[845], line_104[843], line_103[841], line_102[839], line_101[837], line_100[835], line_99[833], line_98[831], line_97[829], line_96[827], line_95[825], line_94[823], line_93[821], line_92[819], line_91[817], line_90[815], line_89[813], line_88[811], line_87[809], line_86[807], line_85[805], line_84[803], line_83[801], line_82[799], line_81[797], line_80[795], line_79[793], line_78[791], line_77[789], line_76[787], line_75[785], line_74[783], line_73[781], line_72[779], line_71[777], line_70[775], line_69[773], line_68[771], line_67[769], line_66[767], line_65[765], line_64[763], line_63[761], line_62[759], line_61[757], line_60[755], line_59[753], line_58[751], line_57[749], line_56[747], line_55[745], line_54[743], line_53[741], line_52[739], line_51[737], line_50[735], line_49[733], line_48[731], line_47[729], line_46[727], line_45[725], line_44[723], line_43[721], line_42[719], line_41[717], line_40[715], line_39[713], line_38[711], line_37[709], line_36[707], line_35[705], line_34[703], line_33[701], line_32[699], line_31[697], line_30[695], line_29[693], line_28[691], line_27[689], line_26[687], line_25[685], line_24[683], line_23[681], line_22[679], line_21[677], line_20[675], line_19[673], line_18[671], line_17[669], line_16[667], line_15[665], line_14[663], line_13[661], line_12[659], line_11[657], line_10[655], line_9[653], line_8[651], line_7[649], line_6[647], line_5[645], line_4[643], line_3[641], line_2[639], line_1[637] };
assign col_892 = {line_128[892], line_127[890], line_126[888], line_125[886], line_124[884], line_123[882], line_122[880], line_121[878], line_120[876], line_119[874], line_118[872], line_117[870], line_116[868], line_115[866], line_114[864], line_113[862], line_112[860], line_111[858], line_110[856], line_109[854], line_108[852], line_107[850], line_106[848], line_105[846], line_104[844], line_103[842], line_102[840], line_101[838], line_100[836], line_99[834], line_98[832], line_97[830], line_96[828], line_95[826], line_94[824], line_93[822], line_92[820], line_91[818], line_90[816], line_89[814], line_88[812], line_87[810], line_86[808], line_85[806], line_84[804], line_83[802], line_82[800], line_81[798], line_80[796], line_79[794], line_78[792], line_77[790], line_76[788], line_75[786], line_74[784], line_73[782], line_72[780], line_71[778], line_70[776], line_69[774], line_68[772], line_67[770], line_66[768], line_65[766], line_64[764], line_63[762], line_62[760], line_61[758], line_60[756], line_59[754], line_58[752], line_57[750], line_56[748], line_55[746], line_54[744], line_53[742], line_52[740], line_51[738], line_50[736], line_49[734], line_48[732], line_47[730], line_46[728], line_45[726], line_44[724], line_43[722], line_42[720], line_41[718], line_40[716], line_39[714], line_38[712], line_37[710], line_36[708], line_35[706], line_34[704], line_33[702], line_32[700], line_31[698], line_30[696], line_29[694], line_28[692], line_27[690], line_26[688], line_25[686], line_24[684], line_23[682], line_22[680], line_21[678], line_20[676], line_19[674], line_18[672], line_17[670], line_16[668], line_15[666], line_14[664], line_13[662], line_12[660], line_11[658], line_10[656], line_9[654], line_8[652], line_7[650], line_6[648], line_5[646], line_4[644], line_3[642], line_2[640], line_1[638] };
assign col_893 = {line_128[893], line_127[891], line_126[889], line_125[887], line_124[885], line_123[883], line_122[881], line_121[879], line_120[877], line_119[875], line_118[873], line_117[871], line_116[869], line_115[867], line_114[865], line_113[863], line_112[861], line_111[859], line_110[857], line_109[855], line_108[853], line_107[851], line_106[849], line_105[847], line_104[845], line_103[843], line_102[841], line_101[839], line_100[837], line_99[835], line_98[833], line_97[831], line_96[829], line_95[827], line_94[825], line_93[823], line_92[821], line_91[819], line_90[817], line_89[815], line_88[813], line_87[811], line_86[809], line_85[807], line_84[805], line_83[803], line_82[801], line_81[799], line_80[797], line_79[795], line_78[793], line_77[791], line_76[789], line_75[787], line_74[785], line_73[783], line_72[781], line_71[779], line_70[777], line_69[775], line_68[773], line_67[771], line_66[769], line_65[767], line_64[765], line_63[763], line_62[761], line_61[759], line_60[757], line_59[755], line_58[753], line_57[751], line_56[749], line_55[747], line_54[745], line_53[743], line_52[741], line_51[739], line_50[737], line_49[735], line_48[733], line_47[731], line_46[729], line_45[727], line_44[725], line_43[723], line_42[721], line_41[719], line_40[717], line_39[715], line_38[713], line_37[711], line_36[709], line_35[707], line_34[705], line_33[703], line_32[701], line_31[699], line_30[697], line_29[695], line_28[693], line_27[691], line_26[689], line_25[687], line_24[685], line_23[683], line_22[681], line_21[679], line_20[677], line_19[675], line_18[673], line_17[671], line_16[669], line_15[667], line_14[665], line_13[663], line_12[661], line_11[659], line_10[657], line_9[655], line_8[653], line_7[651], line_6[649], line_5[647], line_4[645], line_3[643], line_2[641], line_1[639] };
assign col_894 = {line_128[894], line_127[892], line_126[890], line_125[888], line_124[886], line_123[884], line_122[882], line_121[880], line_120[878], line_119[876], line_118[874], line_117[872], line_116[870], line_115[868], line_114[866], line_113[864], line_112[862], line_111[860], line_110[858], line_109[856], line_108[854], line_107[852], line_106[850], line_105[848], line_104[846], line_103[844], line_102[842], line_101[840], line_100[838], line_99[836], line_98[834], line_97[832], line_96[830], line_95[828], line_94[826], line_93[824], line_92[822], line_91[820], line_90[818], line_89[816], line_88[814], line_87[812], line_86[810], line_85[808], line_84[806], line_83[804], line_82[802], line_81[800], line_80[798], line_79[796], line_78[794], line_77[792], line_76[790], line_75[788], line_74[786], line_73[784], line_72[782], line_71[780], line_70[778], line_69[776], line_68[774], line_67[772], line_66[770], line_65[768], line_64[766], line_63[764], line_62[762], line_61[760], line_60[758], line_59[756], line_58[754], line_57[752], line_56[750], line_55[748], line_54[746], line_53[744], line_52[742], line_51[740], line_50[738], line_49[736], line_48[734], line_47[732], line_46[730], line_45[728], line_44[726], line_43[724], line_42[722], line_41[720], line_40[718], line_39[716], line_38[714], line_37[712], line_36[710], line_35[708], line_34[706], line_33[704], line_32[702], line_31[700], line_30[698], line_29[696], line_28[694], line_27[692], line_26[690], line_25[688], line_24[686], line_23[684], line_22[682], line_21[680], line_20[678], line_19[676], line_18[674], line_17[672], line_16[670], line_15[668], line_14[666], line_13[664], line_12[662], line_11[660], line_10[658], line_9[656], line_8[654], line_7[652], line_6[650], line_5[648], line_4[646], line_3[644], line_2[642], line_1[640] };
assign col_895 = {line_128[895], line_127[893], line_126[891], line_125[889], line_124[887], line_123[885], line_122[883], line_121[881], line_120[879], line_119[877], line_118[875], line_117[873], line_116[871], line_115[869], line_114[867], line_113[865], line_112[863], line_111[861], line_110[859], line_109[857], line_108[855], line_107[853], line_106[851], line_105[849], line_104[847], line_103[845], line_102[843], line_101[841], line_100[839], line_99[837], line_98[835], line_97[833], line_96[831], line_95[829], line_94[827], line_93[825], line_92[823], line_91[821], line_90[819], line_89[817], line_88[815], line_87[813], line_86[811], line_85[809], line_84[807], line_83[805], line_82[803], line_81[801], line_80[799], line_79[797], line_78[795], line_77[793], line_76[791], line_75[789], line_74[787], line_73[785], line_72[783], line_71[781], line_70[779], line_69[777], line_68[775], line_67[773], line_66[771], line_65[769], line_64[767], line_63[765], line_62[763], line_61[761], line_60[759], line_59[757], line_58[755], line_57[753], line_56[751], line_55[749], line_54[747], line_53[745], line_52[743], line_51[741], line_50[739], line_49[737], line_48[735], line_47[733], line_46[731], line_45[729], line_44[727], line_43[725], line_42[723], line_41[721], line_40[719], line_39[717], line_38[715], line_37[713], line_36[711], line_35[709], line_34[707], line_33[705], line_32[703], line_31[701], line_30[699], line_29[697], line_28[695], line_27[693], line_26[691], line_25[689], line_24[687], line_23[685], line_22[683], line_21[681], line_20[679], line_19[677], line_18[675], line_17[673], line_16[671], line_15[669], line_14[667], line_13[665], line_12[663], line_11[661], line_10[659], line_9[657], line_8[655], line_7[653], line_6[651], line_5[649], line_4[647], line_3[645], line_2[643], line_1[641] };
assign col_896 = {line_128[896], line_127[894], line_126[892], line_125[890], line_124[888], line_123[886], line_122[884], line_121[882], line_120[880], line_119[878], line_118[876], line_117[874], line_116[872], line_115[870], line_114[868], line_113[866], line_112[864], line_111[862], line_110[860], line_109[858], line_108[856], line_107[854], line_106[852], line_105[850], line_104[848], line_103[846], line_102[844], line_101[842], line_100[840], line_99[838], line_98[836], line_97[834], line_96[832], line_95[830], line_94[828], line_93[826], line_92[824], line_91[822], line_90[820], line_89[818], line_88[816], line_87[814], line_86[812], line_85[810], line_84[808], line_83[806], line_82[804], line_81[802], line_80[800], line_79[798], line_78[796], line_77[794], line_76[792], line_75[790], line_74[788], line_73[786], line_72[784], line_71[782], line_70[780], line_69[778], line_68[776], line_67[774], line_66[772], line_65[770], line_64[768], line_63[766], line_62[764], line_61[762], line_60[760], line_59[758], line_58[756], line_57[754], line_56[752], line_55[750], line_54[748], line_53[746], line_52[744], line_51[742], line_50[740], line_49[738], line_48[736], line_47[734], line_46[732], line_45[730], line_44[728], line_43[726], line_42[724], line_41[722], line_40[720], line_39[718], line_38[716], line_37[714], line_36[712], line_35[710], line_34[708], line_33[706], line_32[704], line_31[702], line_30[700], line_29[698], line_28[696], line_27[694], line_26[692], line_25[690], line_24[688], line_23[686], line_22[684], line_21[682], line_20[680], line_19[678], line_18[676], line_17[674], line_16[672], line_15[670], line_14[668], line_13[666], line_12[664], line_11[662], line_10[660], line_9[658], line_8[656], line_7[654], line_6[652], line_5[650], line_4[648], line_3[646], line_2[644], line_1[642] };
assign col_897 = {line_128[897], line_127[895], line_126[893], line_125[891], line_124[889], line_123[887], line_122[885], line_121[883], line_120[881], line_119[879], line_118[877], line_117[875], line_116[873], line_115[871], line_114[869], line_113[867], line_112[865], line_111[863], line_110[861], line_109[859], line_108[857], line_107[855], line_106[853], line_105[851], line_104[849], line_103[847], line_102[845], line_101[843], line_100[841], line_99[839], line_98[837], line_97[835], line_96[833], line_95[831], line_94[829], line_93[827], line_92[825], line_91[823], line_90[821], line_89[819], line_88[817], line_87[815], line_86[813], line_85[811], line_84[809], line_83[807], line_82[805], line_81[803], line_80[801], line_79[799], line_78[797], line_77[795], line_76[793], line_75[791], line_74[789], line_73[787], line_72[785], line_71[783], line_70[781], line_69[779], line_68[777], line_67[775], line_66[773], line_65[771], line_64[769], line_63[767], line_62[765], line_61[763], line_60[761], line_59[759], line_58[757], line_57[755], line_56[753], line_55[751], line_54[749], line_53[747], line_52[745], line_51[743], line_50[741], line_49[739], line_48[737], line_47[735], line_46[733], line_45[731], line_44[729], line_43[727], line_42[725], line_41[723], line_40[721], line_39[719], line_38[717], line_37[715], line_36[713], line_35[711], line_34[709], line_33[707], line_32[705], line_31[703], line_30[701], line_29[699], line_28[697], line_27[695], line_26[693], line_25[691], line_24[689], line_23[687], line_22[685], line_21[683], line_20[681], line_19[679], line_18[677], line_17[675], line_16[673], line_15[671], line_14[669], line_13[667], line_12[665], line_11[663], line_10[661], line_9[659], line_8[657], line_7[655], line_6[653], line_5[651], line_4[649], line_3[647], line_2[645], line_1[643] };
assign col_898 = {line_128[898], line_127[896], line_126[894], line_125[892], line_124[890], line_123[888], line_122[886], line_121[884], line_120[882], line_119[880], line_118[878], line_117[876], line_116[874], line_115[872], line_114[870], line_113[868], line_112[866], line_111[864], line_110[862], line_109[860], line_108[858], line_107[856], line_106[854], line_105[852], line_104[850], line_103[848], line_102[846], line_101[844], line_100[842], line_99[840], line_98[838], line_97[836], line_96[834], line_95[832], line_94[830], line_93[828], line_92[826], line_91[824], line_90[822], line_89[820], line_88[818], line_87[816], line_86[814], line_85[812], line_84[810], line_83[808], line_82[806], line_81[804], line_80[802], line_79[800], line_78[798], line_77[796], line_76[794], line_75[792], line_74[790], line_73[788], line_72[786], line_71[784], line_70[782], line_69[780], line_68[778], line_67[776], line_66[774], line_65[772], line_64[770], line_63[768], line_62[766], line_61[764], line_60[762], line_59[760], line_58[758], line_57[756], line_56[754], line_55[752], line_54[750], line_53[748], line_52[746], line_51[744], line_50[742], line_49[740], line_48[738], line_47[736], line_46[734], line_45[732], line_44[730], line_43[728], line_42[726], line_41[724], line_40[722], line_39[720], line_38[718], line_37[716], line_36[714], line_35[712], line_34[710], line_33[708], line_32[706], line_31[704], line_30[702], line_29[700], line_28[698], line_27[696], line_26[694], line_25[692], line_24[690], line_23[688], line_22[686], line_21[684], line_20[682], line_19[680], line_18[678], line_17[676], line_16[674], line_15[672], line_14[670], line_13[668], line_12[666], line_11[664], line_10[662], line_9[660], line_8[658], line_7[656], line_6[654], line_5[652], line_4[650], line_3[648], line_2[646], line_1[644] };
assign col_899 = {line_128[899], line_127[897], line_126[895], line_125[893], line_124[891], line_123[889], line_122[887], line_121[885], line_120[883], line_119[881], line_118[879], line_117[877], line_116[875], line_115[873], line_114[871], line_113[869], line_112[867], line_111[865], line_110[863], line_109[861], line_108[859], line_107[857], line_106[855], line_105[853], line_104[851], line_103[849], line_102[847], line_101[845], line_100[843], line_99[841], line_98[839], line_97[837], line_96[835], line_95[833], line_94[831], line_93[829], line_92[827], line_91[825], line_90[823], line_89[821], line_88[819], line_87[817], line_86[815], line_85[813], line_84[811], line_83[809], line_82[807], line_81[805], line_80[803], line_79[801], line_78[799], line_77[797], line_76[795], line_75[793], line_74[791], line_73[789], line_72[787], line_71[785], line_70[783], line_69[781], line_68[779], line_67[777], line_66[775], line_65[773], line_64[771], line_63[769], line_62[767], line_61[765], line_60[763], line_59[761], line_58[759], line_57[757], line_56[755], line_55[753], line_54[751], line_53[749], line_52[747], line_51[745], line_50[743], line_49[741], line_48[739], line_47[737], line_46[735], line_45[733], line_44[731], line_43[729], line_42[727], line_41[725], line_40[723], line_39[721], line_38[719], line_37[717], line_36[715], line_35[713], line_34[711], line_33[709], line_32[707], line_31[705], line_30[703], line_29[701], line_28[699], line_27[697], line_26[695], line_25[693], line_24[691], line_23[689], line_22[687], line_21[685], line_20[683], line_19[681], line_18[679], line_17[677], line_16[675], line_15[673], line_14[671], line_13[669], line_12[667], line_11[665], line_10[663], line_9[661], line_8[659], line_7[657], line_6[655], line_5[653], line_4[651], line_3[649], line_2[647], line_1[645] };
assign col_900 = {line_128[900], line_127[898], line_126[896], line_125[894], line_124[892], line_123[890], line_122[888], line_121[886], line_120[884], line_119[882], line_118[880], line_117[878], line_116[876], line_115[874], line_114[872], line_113[870], line_112[868], line_111[866], line_110[864], line_109[862], line_108[860], line_107[858], line_106[856], line_105[854], line_104[852], line_103[850], line_102[848], line_101[846], line_100[844], line_99[842], line_98[840], line_97[838], line_96[836], line_95[834], line_94[832], line_93[830], line_92[828], line_91[826], line_90[824], line_89[822], line_88[820], line_87[818], line_86[816], line_85[814], line_84[812], line_83[810], line_82[808], line_81[806], line_80[804], line_79[802], line_78[800], line_77[798], line_76[796], line_75[794], line_74[792], line_73[790], line_72[788], line_71[786], line_70[784], line_69[782], line_68[780], line_67[778], line_66[776], line_65[774], line_64[772], line_63[770], line_62[768], line_61[766], line_60[764], line_59[762], line_58[760], line_57[758], line_56[756], line_55[754], line_54[752], line_53[750], line_52[748], line_51[746], line_50[744], line_49[742], line_48[740], line_47[738], line_46[736], line_45[734], line_44[732], line_43[730], line_42[728], line_41[726], line_40[724], line_39[722], line_38[720], line_37[718], line_36[716], line_35[714], line_34[712], line_33[710], line_32[708], line_31[706], line_30[704], line_29[702], line_28[700], line_27[698], line_26[696], line_25[694], line_24[692], line_23[690], line_22[688], line_21[686], line_20[684], line_19[682], line_18[680], line_17[678], line_16[676], line_15[674], line_14[672], line_13[670], line_12[668], line_11[666], line_10[664], line_9[662], line_8[660], line_7[658], line_6[656], line_5[654], line_4[652], line_3[650], line_2[648], line_1[646] };
assign col_901 = {line_128[901], line_127[899], line_126[897], line_125[895], line_124[893], line_123[891], line_122[889], line_121[887], line_120[885], line_119[883], line_118[881], line_117[879], line_116[877], line_115[875], line_114[873], line_113[871], line_112[869], line_111[867], line_110[865], line_109[863], line_108[861], line_107[859], line_106[857], line_105[855], line_104[853], line_103[851], line_102[849], line_101[847], line_100[845], line_99[843], line_98[841], line_97[839], line_96[837], line_95[835], line_94[833], line_93[831], line_92[829], line_91[827], line_90[825], line_89[823], line_88[821], line_87[819], line_86[817], line_85[815], line_84[813], line_83[811], line_82[809], line_81[807], line_80[805], line_79[803], line_78[801], line_77[799], line_76[797], line_75[795], line_74[793], line_73[791], line_72[789], line_71[787], line_70[785], line_69[783], line_68[781], line_67[779], line_66[777], line_65[775], line_64[773], line_63[771], line_62[769], line_61[767], line_60[765], line_59[763], line_58[761], line_57[759], line_56[757], line_55[755], line_54[753], line_53[751], line_52[749], line_51[747], line_50[745], line_49[743], line_48[741], line_47[739], line_46[737], line_45[735], line_44[733], line_43[731], line_42[729], line_41[727], line_40[725], line_39[723], line_38[721], line_37[719], line_36[717], line_35[715], line_34[713], line_33[711], line_32[709], line_31[707], line_30[705], line_29[703], line_28[701], line_27[699], line_26[697], line_25[695], line_24[693], line_23[691], line_22[689], line_21[687], line_20[685], line_19[683], line_18[681], line_17[679], line_16[677], line_15[675], line_14[673], line_13[671], line_12[669], line_11[667], line_10[665], line_9[663], line_8[661], line_7[659], line_6[657], line_5[655], line_4[653], line_3[651], line_2[649], line_1[647] };
assign col_902 = {line_128[902], line_127[900], line_126[898], line_125[896], line_124[894], line_123[892], line_122[890], line_121[888], line_120[886], line_119[884], line_118[882], line_117[880], line_116[878], line_115[876], line_114[874], line_113[872], line_112[870], line_111[868], line_110[866], line_109[864], line_108[862], line_107[860], line_106[858], line_105[856], line_104[854], line_103[852], line_102[850], line_101[848], line_100[846], line_99[844], line_98[842], line_97[840], line_96[838], line_95[836], line_94[834], line_93[832], line_92[830], line_91[828], line_90[826], line_89[824], line_88[822], line_87[820], line_86[818], line_85[816], line_84[814], line_83[812], line_82[810], line_81[808], line_80[806], line_79[804], line_78[802], line_77[800], line_76[798], line_75[796], line_74[794], line_73[792], line_72[790], line_71[788], line_70[786], line_69[784], line_68[782], line_67[780], line_66[778], line_65[776], line_64[774], line_63[772], line_62[770], line_61[768], line_60[766], line_59[764], line_58[762], line_57[760], line_56[758], line_55[756], line_54[754], line_53[752], line_52[750], line_51[748], line_50[746], line_49[744], line_48[742], line_47[740], line_46[738], line_45[736], line_44[734], line_43[732], line_42[730], line_41[728], line_40[726], line_39[724], line_38[722], line_37[720], line_36[718], line_35[716], line_34[714], line_33[712], line_32[710], line_31[708], line_30[706], line_29[704], line_28[702], line_27[700], line_26[698], line_25[696], line_24[694], line_23[692], line_22[690], line_21[688], line_20[686], line_19[684], line_18[682], line_17[680], line_16[678], line_15[676], line_14[674], line_13[672], line_12[670], line_11[668], line_10[666], line_9[664], line_8[662], line_7[660], line_6[658], line_5[656], line_4[654], line_3[652], line_2[650], line_1[648] };
assign col_903 = {line_128[903], line_127[901], line_126[899], line_125[897], line_124[895], line_123[893], line_122[891], line_121[889], line_120[887], line_119[885], line_118[883], line_117[881], line_116[879], line_115[877], line_114[875], line_113[873], line_112[871], line_111[869], line_110[867], line_109[865], line_108[863], line_107[861], line_106[859], line_105[857], line_104[855], line_103[853], line_102[851], line_101[849], line_100[847], line_99[845], line_98[843], line_97[841], line_96[839], line_95[837], line_94[835], line_93[833], line_92[831], line_91[829], line_90[827], line_89[825], line_88[823], line_87[821], line_86[819], line_85[817], line_84[815], line_83[813], line_82[811], line_81[809], line_80[807], line_79[805], line_78[803], line_77[801], line_76[799], line_75[797], line_74[795], line_73[793], line_72[791], line_71[789], line_70[787], line_69[785], line_68[783], line_67[781], line_66[779], line_65[777], line_64[775], line_63[773], line_62[771], line_61[769], line_60[767], line_59[765], line_58[763], line_57[761], line_56[759], line_55[757], line_54[755], line_53[753], line_52[751], line_51[749], line_50[747], line_49[745], line_48[743], line_47[741], line_46[739], line_45[737], line_44[735], line_43[733], line_42[731], line_41[729], line_40[727], line_39[725], line_38[723], line_37[721], line_36[719], line_35[717], line_34[715], line_33[713], line_32[711], line_31[709], line_30[707], line_29[705], line_28[703], line_27[701], line_26[699], line_25[697], line_24[695], line_23[693], line_22[691], line_21[689], line_20[687], line_19[685], line_18[683], line_17[681], line_16[679], line_15[677], line_14[675], line_13[673], line_12[671], line_11[669], line_10[667], line_9[665], line_8[663], line_7[661], line_6[659], line_5[657], line_4[655], line_3[653], line_2[651], line_1[649] };
assign col_904 = {line_128[904], line_127[902], line_126[900], line_125[898], line_124[896], line_123[894], line_122[892], line_121[890], line_120[888], line_119[886], line_118[884], line_117[882], line_116[880], line_115[878], line_114[876], line_113[874], line_112[872], line_111[870], line_110[868], line_109[866], line_108[864], line_107[862], line_106[860], line_105[858], line_104[856], line_103[854], line_102[852], line_101[850], line_100[848], line_99[846], line_98[844], line_97[842], line_96[840], line_95[838], line_94[836], line_93[834], line_92[832], line_91[830], line_90[828], line_89[826], line_88[824], line_87[822], line_86[820], line_85[818], line_84[816], line_83[814], line_82[812], line_81[810], line_80[808], line_79[806], line_78[804], line_77[802], line_76[800], line_75[798], line_74[796], line_73[794], line_72[792], line_71[790], line_70[788], line_69[786], line_68[784], line_67[782], line_66[780], line_65[778], line_64[776], line_63[774], line_62[772], line_61[770], line_60[768], line_59[766], line_58[764], line_57[762], line_56[760], line_55[758], line_54[756], line_53[754], line_52[752], line_51[750], line_50[748], line_49[746], line_48[744], line_47[742], line_46[740], line_45[738], line_44[736], line_43[734], line_42[732], line_41[730], line_40[728], line_39[726], line_38[724], line_37[722], line_36[720], line_35[718], line_34[716], line_33[714], line_32[712], line_31[710], line_30[708], line_29[706], line_28[704], line_27[702], line_26[700], line_25[698], line_24[696], line_23[694], line_22[692], line_21[690], line_20[688], line_19[686], line_18[684], line_17[682], line_16[680], line_15[678], line_14[676], line_13[674], line_12[672], line_11[670], line_10[668], line_9[666], line_8[664], line_7[662], line_6[660], line_5[658], line_4[656], line_3[654], line_2[652], line_1[650] };
assign col_905 = {line_128[905], line_127[903], line_126[901], line_125[899], line_124[897], line_123[895], line_122[893], line_121[891], line_120[889], line_119[887], line_118[885], line_117[883], line_116[881], line_115[879], line_114[877], line_113[875], line_112[873], line_111[871], line_110[869], line_109[867], line_108[865], line_107[863], line_106[861], line_105[859], line_104[857], line_103[855], line_102[853], line_101[851], line_100[849], line_99[847], line_98[845], line_97[843], line_96[841], line_95[839], line_94[837], line_93[835], line_92[833], line_91[831], line_90[829], line_89[827], line_88[825], line_87[823], line_86[821], line_85[819], line_84[817], line_83[815], line_82[813], line_81[811], line_80[809], line_79[807], line_78[805], line_77[803], line_76[801], line_75[799], line_74[797], line_73[795], line_72[793], line_71[791], line_70[789], line_69[787], line_68[785], line_67[783], line_66[781], line_65[779], line_64[777], line_63[775], line_62[773], line_61[771], line_60[769], line_59[767], line_58[765], line_57[763], line_56[761], line_55[759], line_54[757], line_53[755], line_52[753], line_51[751], line_50[749], line_49[747], line_48[745], line_47[743], line_46[741], line_45[739], line_44[737], line_43[735], line_42[733], line_41[731], line_40[729], line_39[727], line_38[725], line_37[723], line_36[721], line_35[719], line_34[717], line_33[715], line_32[713], line_31[711], line_30[709], line_29[707], line_28[705], line_27[703], line_26[701], line_25[699], line_24[697], line_23[695], line_22[693], line_21[691], line_20[689], line_19[687], line_18[685], line_17[683], line_16[681], line_15[679], line_14[677], line_13[675], line_12[673], line_11[671], line_10[669], line_9[667], line_8[665], line_7[663], line_6[661], line_5[659], line_4[657], line_3[655], line_2[653], line_1[651] };
assign col_906 = {line_128[906], line_127[904], line_126[902], line_125[900], line_124[898], line_123[896], line_122[894], line_121[892], line_120[890], line_119[888], line_118[886], line_117[884], line_116[882], line_115[880], line_114[878], line_113[876], line_112[874], line_111[872], line_110[870], line_109[868], line_108[866], line_107[864], line_106[862], line_105[860], line_104[858], line_103[856], line_102[854], line_101[852], line_100[850], line_99[848], line_98[846], line_97[844], line_96[842], line_95[840], line_94[838], line_93[836], line_92[834], line_91[832], line_90[830], line_89[828], line_88[826], line_87[824], line_86[822], line_85[820], line_84[818], line_83[816], line_82[814], line_81[812], line_80[810], line_79[808], line_78[806], line_77[804], line_76[802], line_75[800], line_74[798], line_73[796], line_72[794], line_71[792], line_70[790], line_69[788], line_68[786], line_67[784], line_66[782], line_65[780], line_64[778], line_63[776], line_62[774], line_61[772], line_60[770], line_59[768], line_58[766], line_57[764], line_56[762], line_55[760], line_54[758], line_53[756], line_52[754], line_51[752], line_50[750], line_49[748], line_48[746], line_47[744], line_46[742], line_45[740], line_44[738], line_43[736], line_42[734], line_41[732], line_40[730], line_39[728], line_38[726], line_37[724], line_36[722], line_35[720], line_34[718], line_33[716], line_32[714], line_31[712], line_30[710], line_29[708], line_28[706], line_27[704], line_26[702], line_25[700], line_24[698], line_23[696], line_22[694], line_21[692], line_20[690], line_19[688], line_18[686], line_17[684], line_16[682], line_15[680], line_14[678], line_13[676], line_12[674], line_11[672], line_10[670], line_9[668], line_8[666], line_7[664], line_6[662], line_5[660], line_4[658], line_3[656], line_2[654], line_1[652] };
assign col_907 = {line_128[907], line_127[905], line_126[903], line_125[901], line_124[899], line_123[897], line_122[895], line_121[893], line_120[891], line_119[889], line_118[887], line_117[885], line_116[883], line_115[881], line_114[879], line_113[877], line_112[875], line_111[873], line_110[871], line_109[869], line_108[867], line_107[865], line_106[863], line_105[861], line_104[859], line_103[857], line_102[855], line_101[853], line_100[851], line_99[849], line_98[847], line_97[845], line_96[843], line_95[841], line_94[839], line_93[837], line_92[835], line_91[833], line_90[831], line_89[829], line_88[827], line_87[825], line_86[823], line_85[821], line_84[819], line_83[817], line_82[815], line_81[813], line_80[811], line_79[809], line_78[807], line_77[805], line_76[803], line_75[801], line_74[799], line_73[797], line_72[795], line_71[793], line_70[791], line_69[789], line_68[787], line_67[785], line_66[783], line_65[781], line_64[779], line_63[777], line_62[775], line_61[773], line_60[771], line_59[769], line_58[767], line_57[765], line_56[763], line_55[761], line_54[759], line_53[757], line_52[755], line_51[753], line_50[751], line_49[749], line_48[747], line_47[745], line_46[743], line_45[741], line_44[739], line_43[737], line_42[735], line_41[733], line_40[731], line_39[729], line_38[727], line_37[725], line_36[723], line_35[721], line_34[719], line_33[717], line_32[715], line_31[713], line_30[711], line_29[709], line_28[707], line_27[705], line_26[703], line_25[701], line_24[699], line_23[697], line_22[695], line_21[693], line_20[691], line_19[689], line_18[687], line_17[685], line_16[683], line_15[681], line_14[679], line_13[677], line_12[675], line_11[673], line_10[671], line_9[669], line_8[667], line_7[665], line_6[663], line_5[661], line_4[659], line_3[657], line_2[655], line_1[653] };
assign col_908 = {line_128[908], line_127[906], line_126[904], line_125[902], line_124[900], line_123[898], line_122[896], line_121[894], line_120[892], line_119[890], line_118[888], line_117[886], line_116[884], line_115[882], line_114[880], line_113[878], line_112[876], line_111[874], line_110[872], line_109[870], line_108[868], line_107[866], line_106[864], line_105[862], line_104[860], line_103[858], line_102[856], line_101[854], line_100[852], line_99[850], line_98[848], line_97[846], line_96[844], line_95[842], line_94[840], line_93[838], line_92[836], line_91[834], line_90[832], line_89[830], line_88[828], line_87[826], line_86[824], line_85[822], line_84[820], line_83[818], line_82[816], line_81[814], line_80[812], line_79[810], line_78[808], line_77[806], line_76[804], line_75[802], line_74[800], line_73[798], line_72[796], line_71[794], line_70[792], line_69[790], line_68[788], line_67[786], line_66[784], line_65[782], line_64[780], line_63[778], line_62[776], line_61[774], line_60[772], line_59[770], line_58[768], line_57[766], line_56[764], line_55[762], line_54[760], line_53[758], line_52[756], line_51[754], line_50[752], line_49[750], line_48[748], line_47[746], line_46[744], line_45[742], line_44[740], line_43[738], line_42[736], line_41[734], line_40[732], line_39[730], line_38[728], line_37[726], line_36[724], line_35[722], line_34[720], line_33[718], line_32[716], line_31[714], line_30[712], line_29[710], line_28[708], line_27[706], line_26[704], line_25[702], line_24[700], line_23[698], line_22[696], line_21[694], line_20[692], line_19[690], line_18[688], line_17[686], line_16[684], line_15[682], line_14[680], line_13[678], line_12[676], line_11[674], line_10[672], line_9[670], line_8[668], line_7[666], line_6[664], line_5[662], line_4[660], line_3[658], line_2[656], line_1[654] };
assign col_909 = {line_128[909], line_127[907], line_126[905], line_125[903], line_124[901], line_123[899], line_122[897], line_121[895], line_120[893], line_119[891], line_118[889], line_117[887], line_116[885], line_115[883], line_114[881], line_113[879], line_112[877], line_111[875], line_110[873], line_109[871], line_108[869], line_107[867], line_106[865], line_105[863], line_104[861], line_103[859], line_102[857], line_101[855], line_100[853], line_99[851], line_98[849], line_97[847], line_96[845], line_95[843], line_94[841], line_93[839], line_92[837], line_91[835], line_90[833], line_89[831], line_88[829], line_87[827], line_86[825], line_85[823], line_84[821], line_83[819], line_82[817], line_81[815], line_80[813], line_79[811], line_78[809], line_77[807], line_76[805], line_75[803], line_74[801], line_73[799], line_72[797], line_71[795], line_70[793], line_69[791], line_68[789], line_67[787], line_66[785], line_65[783], line_64[781], line_63[779], line_62[777], line_61[775], line_60[773], line_59[771], line_58[769], line_57[767], line_56[765], line_55[763], line_54[761], line_53[759], line_52[757], line_51[755], line_50[753], line_49[751], line_48[749], line_47[747], line_46[745], line_45[743], line_44[741], line_43[739], line_42[737], line_41[735], line_40[733], line_39[731], line_38[729], line_37[727], line_36[725], line_35[723], line_34[721], line_33[719], line_32[717], line_31[715], line_30[713], line_29[711], line_28[709], line_27[707], line_26[705], line_25[703], line_24[701], line_23[699], line_22[697], line_21[695], line_20[693], line_19[691], line_18[689], line_17[687], line_16[685], line_15[683], line_14[681], line_13[679], line_12[677], line_11[675], line_10[673], line_9[671], line_8[669], line_7[667], line_6[665], line_5[663], line_4[661], line_3[659], line_2[657], line_1[655] };
assign col_910 = {line_128[910], line_127[908], line_126[906], line_125[904], line_124[902], line_123[900], line_122[898], line_121[896], line_120[894], line_119[892], line_118[890], line_117[888], line_116[886], line_115[884], line_114[882], line_113[880], line_112[878], line_111[876], line_110[874], line_109[872], line_108[870], line_107[868], line_106[866], line_105[864], line_104[862], line_103[860], line_102[858], line_101[856], line_100[854], line_99[852], line_98[850], line_97[848], line_96[846], line_95[844], line_94[842], line_93[840], line_92[838], line_91[836], line_90[834], line_89[832], line_88[830], line_87[828], line_86[826], line_85[824], line_84[822], line_83[820], line_82[818], line_81[816], line_80[814], line_79[812], line_78[810], line_77[808], line_76[806], line_75[804], line_74[802], line_73[800], line_72[798], line_71[796], line_70[794], line_69[792], line_68[790], line_67[788], line_66[786], line_65[784], line_64[782], line_63[780], line_62[778], line_61[776], line_60[774], line_59[772], line_58[770], line_57[768], line_56[766], line_55[764], line_54[762], line_53[760], line_52[758], line_51[756], line_50[754], line_49[752], line_48[750], line_47[748], line_46[746], line_45[744], line_44[742], line_43[740], line_42[738], line_41[736], line_40[734], line_39[732], line_38[730], line_37[728], line_36[726], line_35[724], line_34[722], line_33[720], line_32[718], line_31[716], line_30[714], line_29[712], line_28[710], line_27[708], line_26[706], line_25[704], line_24[702], line_23[700], line_22[698], line_21[696], line_20[694], line_19[692], line_18[690], line_17[688], line_16[686], line_15[684], line_14[682], line_13[680], line_12[678], line_11[676], line_10[674], line_9[672], line_8[670], line_7[668], line_6[666], line_5[664], line_4[662], line_3[660], line_2[658], line_1[656] };
assign col_911 = {line_128[911], line_127[909], line_126[907], line_125[905], line_124[903], line_123[901], line_122[899], line_121[897], line_120[895], line_119[893], line_118[891], line_117[889], line_116[887], line_115[885], line_114[883], line_113[881], line_112[879], line_111[877], line_110[875], line_109[873], line_108[871], line_107[869], line_106[867], line_105[865], line_104[863], line_103[861], line_102[859], line_101[857], line_100[855], line_99[853], line_98[851], line_97[849], line_96[847], line_95[845], line_94[843], line_93[841], line_92[839], line_91[837], line_90[835], line_89[833], line_88[831], line_87[829], line_86[827], line_85[825], line_84[823], line_83[821], line_82[819], line_81[817], line_80[815], line_79[813], line_78[811], line_77[809], line_76[807], line_75[805], line_74[803], line_73[801], line_72[799], line_71[797], line_70[795], line_69[793], line_68[791], line_67[789], line_66[787], line_65[785], line_64[783], line_63[781], line_62[779], line_61[777], line_60[775], line_59[773], line_58[771], line_57[769], line_56[767], line_55[765], line_54[763], line_53[761], line_52[759], line_51[757], line_50[755], line_49[753], line_48[751], line_47[749], line_46[747], line_45[745], line_44[743], line_43[741], line_42[739], line_41[737], line_40[735], line_39[733], line_38[731], line_37[729], line_36[727], line_35[725], line_34[723], line_33[721], line_32[719], line_31[717], line_30[715], line_29[713], line_28[711], line_27[709], line_26[707], line_25[705], line_24[703], line_23[701], line_22[699], line_21[697], line_20[695], line_19[693], line_18[691], line_17[689], line_16[687], line_15[685], line_14[683], line_13[681], line_12[679], line_11[677], line_10[675], line_9[673], line_8[671], line_7[669], line_6[667], line_5[665], line_4[663], line_3[661], line_2[659], line_1[657] };
assign col_912 = {line_128[912], line_127[910], line_126[908], line_125[906], line_124[904], line_123[902], line_122[900], line_121[898], line_120[896], line_119[894], line_118[892], line_117[890], line_116[888], line_115[886], line_114[884], line_113[882], line_112[880], line_111[878], line_110[876], line_109[874], line_108[872], line_107[870], line_106[868], line_105[866], line_104[864], line_103[862], line_102[860], line_101[858], line_100[856], line_99[854], line_98[852], line_97[850], line_96[848], line_95[846], line_94[844], line_93[842], line_92[840], line_91[838], line_90[836], line_89[834], line_88[832], line_87[830], line_86[828], line_85[826], line_84[824], line_83[822], line_82[820], line_81[818], line_80[816], line_79[814], line_78[812], line_77[810], line_76[808], line_75[806], line_74[804], line_73[802], line_72[800], line_71[798], line_70[796], line_69[794], line_68[792], line_67[790], line_66[788], line_65[786], line_64[784], line_63[782], line_62[780], line_61[778], line_60[776], line_59[774], line_58[772], line_57[770], line_56[768], line_55[766], line_54[764], line_53[762], line_52[760], line_51[758], line_50[756], line_49[754], line_48[752], line_47[750], line_46[748], line_45[746], line_44[744], line_43[742], line_42[740], line_41[738], line_40[736], line_39[734], line_38[732], line_37[730], line_36[728], line_35[726], line_34[724], line_33[722], line_32[720], line_31[718], line_30[716], line_29[714], line_28[712], line_27[710], line_26[708], line_25[706], line_24[704], line_23[702], line_22[700], line_21[698], line_20[696], line_19[694], line_18[692], line_17[690], line_16[688], line_15[686], line_14[684], line_13[682], line_12[680], line_11[678], line_10[676], line_9[674], line_8[672], line_7[670], line_6[668], line_5[666], line_4[664], line_3[662], line_2[660], line_1[658] };
assign col_913 = {line_128[913], line_127[911], line_126[909], line_125[907], line_124[905], line_123[903], line_122[901], line_121[899], line_120[897], line_119[895], line_118[893], line_117[891], line_116[889], line_115[887], line_114[885], line_113[883], line_112[881], line_111[879], line_110[877], line_109[875], line_108[873], line_107[871], line_106[869], line_105[867], line_104[865], line_103[863], line_102[861], line_101[859], line_100[857], line_99[855], line_98[853], line_97[851], line_96[849], line_95[847], line_94[845], line_93[843], line_92[841], line_91[839], line_90[837], line_89[835], line_88[833], line_87[831], line_86[829], line_85[827], line_84[825], line_83[823], line_82[821], line_81[819], line_80[817], line_79[815], line_78[813], line_77[811], line_76[809], line_75[807], line_74[805], line_73[803], line_72[801], line_71[799], line_70[797], line_69[795], line_68[793], line_67[791], line_66[789], line_65[787], line_64[785], line_63[783], line_62[781], line_61[779], line_60[777], line_59[775], line_58[773], line_57[771], line_56[769], line_55[767], line_54[765], line_53[763], line_52[761], line_51[759], line_50[757], line_49[755], line_48[753], line_47[751], line_46[749], line_45[747], line_44[745], line_43[743], line_42[741], line_41[739], line_40[737], line_39[735], line_38[733], line_37[731], line_36[729], line_35[727], line_34[725], line_33[723], line_32[721], line_31[719], line_30[717], line_29[715], line_28[713], line_27[711], line_26[709], line_25[707], line_24[705], line_23[703], line_22[701], line_21[699], line_20[697], line_19[695], line_18[693], line_17[691], line_16[689], line_15[687], line_14[685], line_13[683], line_12[681], line_11[679], line_10[677], line_9[675], line_8[673], line_7[671], line_6[669], line_5[667], line_4[665], line_3[663], line_2[661], line_1[659] };
assign col_914 = {line_128[914], line_127[912], line_126[910], line_125[908], line_124[906], line_123[904], line_122[902], line_121[900], line_120[898], line_119[896], line_118[894], line_117[892], line_116[890], line_115[888], line_114[886], line_113[884], line_112[882], line_111[880], line_110[878], line_109[876], line_108[874], line_107[872], line_106[870], line_105[868], line_104[866], line_103[864], line_102[862], line_101[860], line_100[858], line_99[856], line_98[854], line_97[852], line_96[850], line_95[848], line_94[846], line_93[844], line_92[842], line_91[840], line_90[838], line_89[836], line_88[834], line_87[832], line_86[830], line_85[828], line_84[826], line_83[824], line_82[822], line_81[820], line_80[818], line_79[816], line_78[814], line_77[812], line_76[810], line_75[808], line_74[806], line_73[804], line_72[802], line_71[800], line_70[798], line_69[796], line_68[794], line_67[792], line_66[790], line_65[788], line_64[786], line_63[784], line_62[782], line_61[780], line_60[778], line_59[776], line_58[774], line_57[772], line_56[770], line_55[768], line_54[766], line_53[764], line_52[762], line_51[760], line_50[758], line_49[756], line_48[754], line_47[752], line_46[750], line_45[748], line_44[746], line_43[744], line_42[742], line_41[740], line_40[738], line_39[736], line_38[734], line_37[732], line_36[730], line_35[728], line_34[726], line_33[724], line_32[722], line_31[720], line_30[718], line_29[716], line_28[714], line_27[712], line_26[710], line_25[708], line_24[706], line_23[704], line_22[702], line_21[700], line_20[698], line_19[696], line_18[694], line_17[692], line_16[690], line_15[688], line_14[686], line_13[684], line_12[682], line_11[680], line_10[678], line_9[676], line_8[674], line_7[672], line_6[670], line_5[668], line_4[666], line_3[664], line_2[662], line_1[660] };
assign col_915 = {line_128[915], line_127[913], line_126[911], line_125[909], line_124[907], line_123[905], line_122[903], line_121[901], line_120[899], line_119[897], line_118[895], line_117[893], line_116[891], line_115[889], line_114[887], line_113[885], line_112[883], line_111[881], line_110[879], line_109[877], line_108[875], line_107[873], line_106[871], line_105[869], line_104[867], line_103[865], line_102[863], line_101[861], line_100[859], line_99[857], line_98[855], line_97[853], line_96[851], line_95[849], line_94[847], line_93[845], line_92[843], line_91[841], line_90[839], line_89[837], line_88[835], line_87[833], line_86[831], line_85[829], line_84[827], line_83[825], line_82[823], line_81[821], line_80[819], line_79[817], line_78[815], line_77[813], line_76[811], line_75[809], line_74[807], line_73[805], line_72[803], line_71[801], line_70[799], line_69[797], line_68[795], line_67[793], line_66[791], line_65[789], line_64[787], line_63[785], line_62[783], line_61[781], line_60[779], line_59[777], line_58[775], line_57[773], line_56[771], line_55[769], line_54[767], line_53[765], line_52[763], line_51[761], line_50[759], line_49[757], line_48[755], line_47[753], line_46[751], line_45[749], line_44[747], line_43[745], line_42[743], line_41[741], line_40[739], line_39[737], line_38[735], line_37[733], line_36[731], line_35[729], line_34[727], line_33[725], line_32[723], line_31[721], line_30[719], line_29[717], line_28[715], line_27[713], line_26[711], line_25[709], line_24[707], line_23[705], line_22[703], line_21[701], line_20[699], line_19[697], line_18[695], line_17[693], line_16[691], line_15[689], line_14[687], line_13[685], line_12[683], line_11[681], line_10[679], line_9[677], line_8[675], line_7[673], line_6[671], line_5[669], line_4[667], line_3[665], line_2[663], line_1[661] };
assign col_916 = {line_128[916], line_127[914], line_126[912], line_125[910], line_124[908], line_123[906], line_122[904], line_121[902], line_120[900], line_119[898], line_118[896], line_117[894], line_116[892], line_115[890], line_114[888], line_113[886], line_112[884], line_111[882], line_110[880], line_109[878], line_108[876], line_107[874], line_106[872], line_105[870], line_104[868], line_103[866], line_102[864], line_101[862], line_100[860], line_99[858], line_98[856], line_97[854], line_96[852], line_95[850], line_94[848], line_93[846], line_92[844], line_91[842], line_90[840], line_89[838], line_88[836], line_87[834], line_86[832], line_85[830], line_84[828], line_83[826], line_82[824], line_81[822], line_80[820], line_79[818], line_78[816], line_77[814], line_76[812], line_75[810], line_74[808], line_73[806], line_72[804], line_71[802], line_70[800], line_69[798], line_68[796], line_67[794], line_66[792], line_65[790], line_64[788], line_63[786], line_62[784], line_61[782], line_60[780], line_59[778], line_58[776], line_57[774], line_56[772], line_55[770], line_54[768], line_53[766], line_52[764], line_51[762], line_50[760], line_49[758], line_48[756], line_47[754], line_46[752], line_45[750], line_44[748], line_43[746], line_42[744], line_41[742], line_40[740], line_39[738], line_38[736], line_37[734], line_36[732], line_35[730], line_34[728], line_33[726], line_32[724], line_31[722], line_30[720], line_29[718], line_28[716], line_27[714], line_26[712], line_25[710], line_24[708], line_23[706], line_22[704], line_21[702], line_20[700], line_19[698], line_18[696], line_17[694], line_16[692], line_15[690], line_14[688], line_13[686], line_12[684], line_11[682], line_10[680], line_9[678], line_8[676], line_7[674], line_6[672], line_5[670], line_4[668], line_3[666], line_2[664], line_1[662] };
assign col_917 = {line_128[917], line_127[915], line_126[913], line_125[911], line_124[909], line_123[907], line_122[905], line_121[903], line_120[901], line_119[899], line_118[897], line_117[895], line_116[893], line_115[891], line_114[889], line_113[887], line_112[885], line_111[883], line_110[881], line_109[879], line_108[877], line_107[875], line_106[873], line_105[871], line_104[869], line_103[867], line_102[865], line_101[863], line_100[861], line_99[859], line_98[857], line_97[855], line_96[853], line_95[851], line_94[849], line_93[847], line_92[845], line_91[843], line_90[841], line_89[839], line_88[837], line_87[835], line_86[833], line_85[831], line_84[829], line_83[827], line_82[825], line_81[823], line_80[821], line_79[819], line_78[817], line_77[815], line_76[813], line_75[811], line_74[809], line_73[807], line_72[805], line_71[803], line_70[801], line_69[799], line_68[797], line_67[795], line_66[793], line_65[791], line_64[789], line_63[787], line_62[785], line_61[783], line_60[781], line_59[779], line_58[777], line_57[775], line_56[773], line_55[771], line_54[769], line_53[767], line_52[765], line_51[763], line_50[761], line_49[759], line_48[757], line_47[755], line_46[753], line_45[751], line_44[749], line_43[747], line_42[745], line_41[743], line_40[741], line_39[739], line_38[737], line_37[735], line_36[733], line_35[731], line_34[729], line_33[727], line_32[725], line_31[723], line_30[721], line_29[719], line_28[717], line_27[715], line_26[713], line_25[711], line_24[709], line_23[707], line_22[705], line_21[703], line_20[701], line_19[699], line_18[697], line_17[695], line_16[693], line_15[691], line_14[689], line_13[687], line_12[685], line_11[683], line_10[681], line_9[679], line_8[677], line_7[675], line_6[673], line_5[671], line_4[669], line_3[667], line_2[665], line_1[663] };
assign col_918 = {line_128[918], line_127[916], line_126[914], line_125[912], line_124[910], line_123[908], line_122[906], line_121[904], line_120[902], line_119[900], line_118[898], line_117[896], line_116[894], line_115[892], line_114[890], line_113[888], line_112[886], line_111[884], line_110[882], line_109[880], line_108[878], line_107[876], line_106[874], line_105[872], line_104[870], line_103[868], line_102[866], line_101[864], line_100[862], line_99[860], line_98[858], line_97[856], line_96[854], line_95[852], line_94[850], line_93[848], line_92[846], line_91[844], line_90[842], line_89[840], line_88[838], line_87[836], line_86[834], line_85[832], line_84[830], line_83[828], line_82[826], line_81[824], line_80[822], line_79[820], line_78[818], line_77[816], line_76[814], line_75[812], line_74[810], line_73[808], line_72[806], line_71[804], line_70[802], line_69[800], line_68[798], line_67[796], line_66[794], line_65[792], line_64[790], line_63[788], line_62[786], line_61[784], line_60[782], line_59[780], line_58[778], line_57[776], line_56[774], line_55[772], line_54[770], line_53[768], line_52[766], line_51[764], line_50[762], line_49[760], line_48[758], line_47[756], line_46[754], line_45[752], line_44[750], line_43[748], line_42[746], line_41[744], line_40[742], line_39[740], line_38[738], line_37[736], line_36[734], line_35[732], line_34[730], line_33[728], line_32[726], line_31[724], line_30[722], line_29[720], line_28[718], line_27[716], line_26[714], line_25[712], line_24[710], line_23[708], line_22[706], line_21[704], line_20[702], line_19[700], line_18[698], line_17[696], line_16[694], line_15[692], line_14[690], line_13[688], line_12[686], line_11[684], line_10[682], line_9[680], line_8[678], line_7[676], line_6[674], line_5[672], line_4[670], line_3[668], line_2[666], line_1[664] };
assign col_919 = {line_128[919], line_127[917], line_126[915], line_125[913], line_124[911], line_123[909], line_122[907], line_121[905], line_120[903], line_119[901], line_118[899], line_117[897], line_116[895], line_115[893], line_114[891], line_113[889], line_112[887], line_111[885], line_110[883], line_109[881], line_108[879], line_107[877], line_106[875], line_105[873], line_104[871], line_103[869], line_102[867], line_101[865], line_100[863], line_99[861], line_98[859], line_97[857], line_96[855], line_95[853], line_94[851], line_93[849], line_92[847], line_91[845], line_90[843], line_89[841], line_88[839], line_87[837], line_86[835], line_85[833], line_84[831], line_83[829], line_82[827], line_81[825], line_80[823], line_79[821], line_78[819], line_77[817], line_76[815], line_75[813], line_74[811], line_73[809], line_72[807], line_71[805], line_70[803], line_69[801], line_68[799], line_67[797], line_66[795], line_65[793], line_64[791], line_63[789], line_62[787], line_61[785], line_60[783], line_59[781], line_58[779], line_57[777], line_56[775], line_55[773], line_54[771], line_53[769], line_52[767], line_51[765], line_50[763], line_49[761], line_48[759], line_47[757], line_46[755], line_45[753], line_44[751], line_43[749], line_42[747], line_41[745], line_40[743], line_39[741], line_38[739], line_37[737], line_36[735], line_35[733], line_34[731], line_33[729], line_32[727], line_31[725], line_30[723], line_29[721], line_28[719], line_27[717], line_26[715], line_25[713], line_24[711], line_23[709], line_22[707], line_21[705], line_20[703], line_19[701], line_18[699], line_17[697], line_16[695], line_15[693], line_14[691], line_13[689], line_12[687], line_11[685], line_10[683], line_9[681], line_8[679], line_7[677], line_6[675], line_5[673], line_4[671], line_3[669], line_2[667], line_1[665] };
assign col_920 = {line_128[920], line_127[918], line_126[916], line_125[914], line_124[912], line_123[910], line_122[908], line_121[906], line_120[904], line_119[902], line_118[900], line_117[898], line_116[896], line_115[894], line_114[892], line_113[890], line_112[888], line_111[886], line_110[884], line_109[882], line_108[880], line_107[878], line_106[876], line_105[874], line_104[872], line_103[870], line_102[868], line_101[866], line_100[864], line_99[862], line_98[860], line_97[858], line_96[856], line_95[854], line_94[852], line_93[850], line_92[848], line_91[846], line_90[844], line_89[842], line_88[840], line_87[838], line_86[836], line_85[834], line_84[832], line_83[830], line_82[828], line_81[826], line_80[824], line_79[822], line_78[820], line_77[818], line_76[816], line_75[814], line_74[812], line_73[810], line_72[808], line_71[806], line_70[804], line_69[802], line_68[800], line_67[798], line_66[796], line_65[794], line_64[792], line_63[790], line_62[788], line_61[786], line_60[784], line_59[782], line_58[780], line_57[778], line_56[776], line_55[774], line_54[772], line_53[770], line_52[768], line_51[766], line_50[764], line_49[762], line_48[760], line_47[758], line_46[756], line_45[754], line_44[752], line_43[750], line_42[748], line_41[746], line_40[744], line_39[742], line_38[740], line_37[738], line_36[736], line_35[734], line_34[732], line_33[730], line_32[728], line_31[726], line_30[724], line_29[722], line_28[720], line_27[718], line_26[716], line_25[714], line_24[712], line_23[710], line_22[708], line_21[706], line_20[704], line_19[702], line_18[700], line_17[698], line_16[696], line_15[694], line_14[692], line_13[690], line_12[688], line_11[686], line_10[684], line_9[682], line_8[680], line_7[678], line_6[676], line_5[674], line_4[672], line_3[670], line_2[668], line_1[666] };
assign col_921 = {line_128[921], line_127[919], line_126[917], line_125[915], line_124[913], line_123[911], line_122[909], line_121[907], line_120[905], line_119[903], line_118[901], line_117[899], line_116[897], line_115[895], line_114[893], line_113[891], line_112[889], line_111[887], line_110[885], line_109[883], line_108[881], line_107[879], line_106[877], line_105[875], line_104[873], line_103[871], line_102[869], line_101[867], line_100[865], line_99[863], line_98[861], line_97[859], line_96[857], line_95[855], line_94[853], line_93[851], line_92[849], line_91[847], line_90[845], line_89[843], line_88[841], line_87[839], line_86[837], line_85[835], line_84[833], line_83[831], line_82[829], line_81[827], line_80[825], line_79[823], line_78[821], line_77[819], line_76[817], line_75[815], line_74[813], line_73[811], line_72[809], line_71[807], line_70[805], line_69[803], line_68[801], line_67[799], line_66[797], line_65[795], line_64[793], line_63[791], line_62[789], line_61[787], line_60[785], line_59[783], line_58[781], line_57[779], line_56[777], line_55[775], line_54[773], line_53[771], line_52[769], line_51[767], line_50[765], line_49[763], line_48[761], line_47[759], line_46[757], line_45[755], line_44[753], line_43[751], line_42[749], line_41[747], line_40[745], line_39[743], line_38[741], line_37[739], line_36[737], line_35[735], line_34[733], line_33[731], line_32[729], line_31[727], line_30[725], line_29[723], line_28[721], line_27[719], line_26[717], line_25[715], line_24[713], line_23[711], line_22[709], line_21[707], line_20[705], line_19[703], line_18[701], line_17[699], line_16[697], line_15[695], line_14[693], line_13[691], line_12[689], line_11[687], line_10[685], line_9[683], line_8[681], line_7[679], line_6[677], line_5[675], line_4[673], line_3[671], line_2[669], line_1[667] };
assign col_922 = {line_128[922], line_127[920], line_126[918], line_125[916], line_124[914], line_123[912], line_122[910], line_121[908], line_120[906], line_119[904], line_118[902], line_117[900], line_116[898], line_115[896], line_114[894], line_113[892], line_112[890], line_111[888], line_110[886], line_109[884], line_108[882], line_107[880], line_106[878], line_105[876], line_104[874], line_103[872], line_102[870], line_101[868], line_100[866], line_99[864], line_98[862], line_97[860], line_96[858], line_95[856], line_94[854], line_93[852], line_92[850], line_91[848], line_90[846], line_89[844], line_88[842], line_87[840], line_86[838], line_85[836], line_84[834], line_83[832], line_82[830], line_81[828], line_80[826], line_79[824], line_78[822], line_77[820], line_76[818], line_75[816], line_74[814], line_73[812], line_72[810], line_71[808], line_70[806], line_69[804], line_68[802], line_67[800], line_66[798], line_65[796], line_64[794], line_63[792], line_62[790], line_61[788], line_60[786], line_59[784], line_58[782], line_57[780], line_56[778], line_55[776], line_54[774], line_53[772], line_52[770], line_51[768], line_50[766], line_49[764], line_48[762], line_47[760], line_46[758], line_45[756], line_44[754], line_43[752], line_42[750], line_41[748], line_40[746], line_39[744], line_38[742], line_37[740], line_36[738], line_35[736], line_34[734], line_33[732], line_32[730], line_31[728], line_30[726], line_29[724], line_28[722], line_27[720], line_26[718], line_25[716], line_24[714], line_23[712], line_22[710], line_21[708], line_20[706], line_19[704], line_18[702], line_17[700], line_16[698], line_15[696], line_14[694], line_13[692], line_12[690], line_11[688], line_10[686], line_9[684], line_8[682], line_7[680], line_6[678], line_5[676], line_4[674], line_3[672], line_2[670], line_1[668] };
assign col_923 = {line_128[923], line_127[921], line_126[919], line_125[917], line_124[915], line_123[913], line_122[911], line_121[909], line_120[907], line_119[905], line_118[903], line_117[901], line_116[899], line_115[897], line_114[895], line_113[893], line_112[891], line_111[889], line_110[887], line_109[885], line_108[883], line_107[881], line_106[879], line_105[877], line_104[875], line_103[873], line_102[871], line_101[869], line_100[867], line_99[865], line_98[863], line_97[861], line_96[859], line_95[857], line_94[855], line_93[853], line_92[851], line_91[849], line_90[847], line_89[845], line_88[843], line_87[841], line_86[839], line_85[837], line_84[835], line_83[833], line_82[831], line_81[829], line_80[827], line_79[825], line_78[823], line_77[821], line_76[819], line_75[817], line_74[815], line_73[813], line_72[811], line_71[809], line_70[807], line_69[805], line_68[803], line_67[801], line_66[799], line_65[797], line_64[795], line_63[793], line_62[791], line_61[789], line_60[787], line_59[785], line_58[783], line_57[781], line_56[779], line_55[777], line_54[775], line_53[773], line_52[771], line_51[769], line_50[767], line_49[765], line_48[763], line_47[761], line_46[759], line_45[757], line_44[755], line_43[753], line_42[751], line_41[749], line_40[747], line_39[745], line_38[743], line_37[741], line_36[739], line_35[737], line_34[735], line_33[733], line_32[731], line_31[729], line_30[727], line_29[725], line_28[723], line_27[721], line_26[719], line_25[717], line_24[715], line_23[713], line_22[711], line_21[709], line_20[707], line_19[705], line_18[703], line_17[701], line_16[699], line_15[697], line_14[695], line_13[693], line_12[691], line_11[689], line_10[687], line_9[685], line_8[683], line_7[681], line_6[679], line_5[677], line_4[675], line_3[673], line_2[671], line_1[669] };
assign col_924 = {line_128[924], line_127[922], line_126[920], line_125[918], line_124[916], line_123[914], line_122[912], line_121[910], line_120[908], line_119[906], line_118[904], line_117[902], line_116[900], line_115[898], line_114[896], line_113[894], line_112[892], line_111[890], line_110[888], line_109[886], line_108[884], line_107[882], line_106[880], line_105[878], line_104[876], line_103[874], line_102[872], line_101[870], line_100[868], line_99[866], line_98[864], line_97[862], line_96[860], line_95[858], line_94[856], line_93[854], line_92[852], line_91[850], line_90[848], line_89[846], line_88[844], line_87[842], line_86[840], line_85[838], line_84[836], line_83[834], line_82[832], line_81[830], line_80[828], line_79[826], line_78[824], line_77[822], line_76[820], line_75[818], line_74[816], line_73[814], line_72[812], line_71[810], line_70[808], line_69[806], line_68[804], line_67[802], line_66[800], line_65[798], line_64[796], line_63[794], line_62[792], line_61[790], line_60[788], line_59[786], line_58[784], line_57[782], line_56[780], line_55[778], line_54[776], line_53[774], line_52[772], line_51[770], line_50[768], line_49[766], line_48[764], line_47[762], line_46[760], line_45[758], line_44[756], line_43[754], line_42[752], line_41[750], line_40[748], line_39[746], line_38[744], line_37[742], line_36[740], line_35[738], line_34[736], line_33[734], line_32[732], line_31[730], line_30[728], line_29[726], line_28[724], line_27[722], line_26[720], line_25[718], line_24[716], line_23[714], line_22[712], line_21[710], line_20[708], line_19[706], line_18[704], line_17[702], line_16[700], line_15[698], line_14[696], line_13[694], line_12[692], line_11[690], line_10[688], line_9[686], line_8[684], line_7[682], line_6[680], line_5[678], line_4[676], line_3[674], line_2[672], line_1[670] };
assign col_925 = {line_128[925], line_127[923], line_126[921], line_125[919], line_124[917], line_123[915], line_122[913], line_121[911], line_120[909], line_119[907], line_118[905], line_117[903], line_116[901], line_115[899], line_114[897], line_113[895], line_112[893], line_111[891], line_110[889], line_109[887], line_108[885], line_107[883], line_106[881], line_105[879], line_104[877], line_103[875], line_102[873], line_101[871], line_100[869], line_99[867], line_98[865], line_97[863], line_96[861], line_95[859], line_94[857], line_93[855], line_92[853], line_91[851], line_90[849], line_89[847], line_88[845], line_87[843], line_86[841], line_85[839], line_84[837], line_83[835], line_82[833], line_81[831], line_80[829], line_79[827], line_78[825], line_77[823], line_76[821], line_75[819], line_74[817], line_73[815], line_72[813], line_71[811], line_70[809], line_69[807], line_68[805], line_67[803], line_66[801], line_65[799], line_64[797], line_63[795], line_62[793], line_61[791], line_60[789], line_59[787], line_58[785], line_57[783], line_56[781], line_55[779], line_54[777], line_53[775], line_52[773], line_51[771], line_50[769], line_49[767], line_48[765], line_47[763], line_46[761], line_45[759], line_44[757], line_43[755], line_42[753], line_41[751], line_40[749], line_39[747], line_38[745], line_37[743], line_36[741], line_35[739], line_34[737], line_33[735], line_32[733], line_31[731], line_30[729], line_29[727], line_28[725], line_27[723], line_26[721], line_25[719], line_24[717], line_23[715], line_22[713], line_21[711], line_20[709], line_19[707], line_18[705], line_17[703], line_16[701], line_15[699], line_14[697], line_13[695], line_12[693], line_11[691], line_10[689], line_9[687], line_8[685], line_7[683], line_6[681], line_5[679], line_4[677], line_3[675], line_2[673], line_1[671] };
assign col_926 = {line_128[926], line_127[924], line_126[922], line_125[920], line_124[918], line_123[916], line_122[914], line_121[912], line_120[910], line_119[908], line_118[906], line_117[904], line_116[902], line_115[900], line_114[898], line_113[896], line_112[894], line_111[892], line_110[890], line_109[888], line_108[886], line_107[884], line_106[882], line_105[880], line_104[878], line_103[876], line_102[874], line_101[872], line_100[870], line_99[868], line_98[866], line_97[864], line_96[862], line_95[860], line_94[858], line_93[856], line_92[854], line_91[852], line_90[850], line_89[848], line_88[846], line_87[844], line_86[842], line_85[840], line_84[838], line_83[836], line_82[834], line_81[832], line_80[830], line_79[828], line_78[826], line_77[824], line_76[822], line_75[820], line_74[818], line_73[816], line_72[814], line_71[812], line_70[810], line_69[808], line_68[806], line_67[804], line_66[802], line_65[800], line_64[798], line_63[796], line_62[794], line_61[792], line_60[790], line_59[788], line_58[786], line_57[784], line_56[782], line_55[780], line_54[778], line_53[776], line_52[774], line_51[772], line_50[770], line_49[768], line_48[766], line_47[764], line_46[762], line_45[760], line_44[758], line_43[756], line_42[754], line_41[752], line_40[750], line_39[748], line_38[746], line_37[744], line_36[742], line_35[740], line_34[738], line_33[736], line_32[734], line_31[732], line_30[730], line_29[728], line_28[726], line_27[724], line_26[722], line_25[720], line_24[718], line_23[716], line_22[714], line_21[712], line_20[710], line_19[708], line_18[706], line_17[704], line_16[702], line_15[700], line_14[698], line_13[696], line_12[694], line_11[692], line_10[690], line_9[688], line_8[686], line_7[684], line_6[682], line_5[680], line_4[678], line_3[676], line_2[674], line_1[672] };
assign col_927 = {line_128[927], line_127[925], line_126[923], line_125[921], line_124[919], line_123[917], line_122[915], line_121[913], line_120[911], line_119[909], line_118[907], line_117[905], line_116[903], line_115[901], line_114[899], line_113[897], line_112[895], line_111[893], line_110[891], line_109[889], line_108[887], line_107[885], line_106[883], line_105[881], line_104[879], line_103[877], line_102[875], line_101[873], line_100[871], line_99[869], line_98[867], line_97[865], line_96[863], line_95[861], line_94[859], line_93[857], line_92[855], line_91[853], line_90[851], line_89[849], line_88[847], line_87[845], line_86[843], line_85[841], line_84[839], line_83[837], line_82[835], line_81[833], line_80[831], line_79[829], line_78[827], line_77[825], line_76[823], line_75[821], line_74[819], line_73[817], line_72[815], line_71[813], line_70[811], line_69[809], line_68[807], line_67[805], line_66[803], line_65[801], line_64[799], line_63[797], line_62[795], line_61[793], line_60[791], line_59[789], line_58[787], line_57[785], line_56[783], line_55[781], line_54[779], line_53[777], line_52[775], line_51[773], line_50[771], line_49[769], line_48[767], line_47[765], line_46[763], line_45[761], line_44[759], line_43[757], line_42[755], line_41[753], line_40[751], line_39[749], line_38[747], line_37[745], line_36[743], line_35[741], line_34[739], line_33[737], line_32[735], line_31[733], line_30[731], line_29[729], line_28[727], line_27[725], line_26[723], line_25[721], line_24[719], line_23[717], line_22[715], line_21[713], line_20[711], line_19[709], line_18[707], line_17[705], line_16[703], line_15[701], line_14[699], line_13[697], line_12[695], line_11[693], line_10[691], line_9[689], line_8[687], line_7[685], line_6[683], line_5[681], line_4[679], line_3[677], line_2[675], line_1[673] };
assign col_928 = {line_128[928], line_127[926], line_126[924], line_125[922], line_124[920], line_123[918], line_122[916], line_121[914], line_120[912], line_119[910], line_118[908], line_117[906], line_116[904], line_115[902], line_114[900], line_113[898], line_112[896], line_111[894], line_110[892], line_109[890], line_108[888], line_107[886], line_106[884], line_105[882], line_104[880], line_103[878], line_102[876], line_101[874], line_100[872], line_99[870], line_98[868], line_97[866], line_96[864], line_95[862], line_94[860], line_93[858], line_92[856], line_91[854], line_90[852], line_89[850], line_88[848], line_87[846], line_86[844], line_85[842], line_84[840], line_83[838], line_82[836], line_81[834], line_80[832], line_79[830], line_78[828], line_77[826], line_76[824], line_75[822], line_74[820], line_73[818], line_72[816], line_71[814], line_70[812], line_69[810], line_68[808], line_67[806], line_66[804], line_65[802], line_64[800], line_63[798], line_62[796], line_61[794], line_60[792], line_59[790], line_58[788], line_57[786], line_56[784], line_55[782], line_54[780], line_53[778], line_52[776], line_51[774], line_50[772], line_49[770], line_48[768], line_47[766], line_46[764], line_45[762], line_44[760], line_43[758], line_42[756], line_41[754], line_40[752], line_39[750], line_38[748], line_37[746], line_36[744], line_35[742], line_34[740], line_33[738], line_32[736], line_31[734], line_30[732], line_29[730], line_28[728], line_27[726], line_26[724], line_25[722], line_24[720], line_23[718], line_22[716], line_21[714], line_20[712], line_19[710], line_18[708], line_17[706], line_16[704], line_15[702], line_14[700], line_13[698], line_12[696], line_11[694], line_10[692], line_9[690], line_8[688], line_7[686], line_6[684], line_5[682], line_4[680], line_3[678], line_2[676], line_1[674] };
assign col_929 = {line_128[929], line_127[927], line_126[925], line_125[923], line_124[921], line_123[919], line_122[917], line_121[915], line_120[913], line_119[911], line_118[909], line_117[907], line_116[905], line_115[903], line_114[901], line_113[899], line_112[897], line_111[895], line_110[893], line_109[891], line_108[889], line_107[887], line_106[885], line_105[883], line_104[881], line_103[879], line_102[877], line_101[875], line_100[873], line_99[871], line_98[869], line_97[867], line_96[865], line_95[863], line_94[861], line_93[859], line_92[857], line_91[855], line_90[853], line_89[851], line_88[849], line_87[847], line_86[845], line_85[843], line_84[841], line_83[839], line_82[837], line_81[835], line_80[833], line_79[831], line_78[829], line_77[827], line_76[825], line_75[823], line_74[821], line_73[819], line_72[817], line_71[815], line_70[813], line_69[811], line_68[809], line_67[807], line_66[805], line_65[803], line_64[801], line_63[799], line_62[797], line_61[795], line_60[793], line_59[791], line_58[789], line_57[787], line_56[785], line_55[783], line_54[781], line_53[779], line_52[777], line_51[775], line_50[773], line_49[771], line_48[769], line_47[767], line_46[765], line_45[763], line_44[761], line_43[759], line_42[757], line_41[755], line_40[753], line_39[751], line_38[749], line_37[747], line_36[745], line_35[743], line_34[741], line_33[739], line_32[737], line_31[735], line_30[733], line_29[731], line_28[729], line_27[727], line_26[725], line_25[723], line_24[721], line_23[719], line_22[717], line_21[715], line_20[713], line_19[711], line_18[709], line_17[707], line_16[705], line_15[703], line_14[701], line_13[699], line_12[697], line_11[695], line_10[693], line_9[691], line_8[689], line_7[687], line_6[685], line_5[683], line_4[681], line_3[679], line_2[677], line_1[675] };
assign col_930 = {line_128[930], line_127[928], line_126[926], line_125[924], line_124[922], line_123[920], line_122[918], line_121[916], line_120[914], line_119[912], line_118[910], line_117[908], line_116[906], line_115[904], line_114[902], line_113[900], line_112[898], line_111[896], line_110[894], line_109[892], line_108[890], line_107[888], line_106[886], line_105[884], line_104[882], line_103[880], line_102[878], line_101[876], line_100[874], line_99[872], line_98[870], line_97[868], line_96[866], line_95[864], line_94[862], line_93[860], line_92[858], line_91[856], line_90[854], line_89[852], line_88[850], line_87[848], line_86[846], line_85[844], line_84[842], line_83[840], line_82[838], line_81[836], line_80[834], line_79[832], line_78[830], line_77[828], line_76[826], line_75[824], line_74[822], line_73[820], line_72[818], line_71[816], line_70[814], line_69[812], line_68[810], line_67[808], line_66[806], line_65[804], line_64[802], line_63[800], line_62[798], line_61[796], line_60[794], line_59[792], line_58[790], line_57[788], line_56[786], line_55[784], line_54[782], line_53[780], line_52[778], line_51[776], line_50[774], line_49[772], line_48[770], line_47[768], line_46[766], line_45[764], line_44[762], line_43[760], line_42[758], line_41[756], line_40[754], line_39[752], line_38[750], line_37[748], line_36[746], line_35[744], line_34[742], line_33[740], line_32[738], line_31[736], line_30[734], line_29[732], line_28[730], line_27[728], line_26[726], line_25[724], line_24[722], line_23[720], line_22[718], line_21[716], line_20[714], line_19[712], line_18[710], line_17[708], line_16[706], line_15[704], line_14[702], line_13[700], line_12[698], line_11[696], line_10[694], line_9[692], line_8[690], line_7[688], line_6[686], line_5[684], line_4[682], line_3[680], line_2[678], line_1[676] };
assign col_931 = {line_128[931], line_127[929], line_126[927], line_125[925], line_124[923], line_123[921], line_122[919], line_121[917], line_120[915], line_119[913], line_118[911], line_117[909], line_116[907], line_115[905], line_114[903], line_113[901], line_112[899], line_111[897], line_110[895], line_109[893], line_108[891], line_107[889], line_106[887], line_105[885], line_104[883], line_103[881], line_102[879], line_101[877], line_100[875], line_99[873], line_98[871], line_97[869], line_96[867], line_95[865], line_94[863], line_93[861], line_92[859], line_91[857], line_90[855], line_89[853], line_88[851], line_87[849], line_86[847], line_85[845], line_84[843], line_83[841], line_82[839], line_81[837], line_80[835], line_79[833], line_78[831], line_77[829], line_76[827], line_75[825], line_74[823], line_73[821], line_72[819], line_71[817], line_70[815], line_69[813], line_68[811], line_67[809], line_66[807], line_65[805], line_64[803], line_63[801], line_62[799], line_61[797], line_60[795], line_59[793], line_58[791], line_57[789], line_56[787], line_55[785], line_54[783], line_53[781], line_52[779], line_51[777], line_50[775], line_49[773], line_48[771], line_47[769], line_46[767], line_45[765], line_44[763], line_43[761], line_42[759], line_41[757], line_40[755], line_39[753], line_38[751], line_37[749], line_36[747], line_35[745], line_34[743], line_33[741], line_32[739], line_31[737], line_30[735], line_29[733], line_28[731], line_27[729], line_26[727], line_25[725], line_24[723], line_23[721], line_22[719], line_21[717], line_20[715], line_19[713], line_18[711], line_17[709], line_16[707], line_15[705], line_14[703], line_13[701], line_12[699], line_11[697], line_10[695], line_9[693], line_8[691], line_7[689], line_6[687], line_5[685], line_4[683], line_3[681], line_2[679], line_1[677] };
assign col_932 = {line_128[932], line_127[930], line_126[928], line_125[926], line_124[924], line_123[922], line_122[920], line_121[918], line_120[916], line_119[914], line_118[912], line_117[910], line_116[908], line_115[906], line_114[904], line_113[902], line_112[900], line_111[898], line_110[896], line_109[894], line_108[892], line_107[890], line_106[888], line_105[886], line_104[884], line_103[882], line_102[880], line_101[878], line_100[876], line_99[874], line_98[872], line_97[870], line_96[868], line_95[866], line_94[864], line_93[862], line_92[860], line_91[858], line_90[856], line_89[854], line_88[852], line_87[850], line_86[848], line_85[846], line_84[844], line_83[842], line_82[840], line_81[838], line_80[836], line_79[834], line_78[832], line_77[830], line_76[828], line_75[826], line_74[824], line_73[822], line_72[820], line_71[818], line_70[816], line_69[814], line_68[812], line_67[810], line_66[808], line_65[806], line_64[804], line_63[802], line_62[800], line_61[798], line_60[796], line_59[794], line_58[792], line_57[790], line_56[788], line_55[786], line_54[784], line_53[782], line_52[780], line_51[778], line_50[776], line_49[774], line_48[772], line_47[770], line_46[768], line_45[766], line_44[764], line_43[762], line_42[760], line_41[758], line_40[756], line_39[754], line_38[752], line_37[750], line_36[748], line_35[746], line_34[744], line_33[742], line_32[740], line_31[738], line_30[736], line_29[734], line_28[732], line_27[730], line_26[728], line_25[726], line_24[724], line_23[722], line_22[720], line_21[718], line_20[716], line_19[714], line_18[712], line_17[710], line_16[708], line_15[706], line_14[704], line_13[702], line_12[700], line_11[698], line_10[696], line_9[694], line_8[692], line_7[690], line_6[688], line_5[686], line_4[684], line_3[682], line_2[680], line_1[678] };
assign col_933 = {line_128[933], line_127[931], line_126[929], line_125[927], line_124[925], line_123[923], line_122[921], line_121[919], line_120[917], line_119[915], line_118[913], line_117[911], line_116[909], line_115[907], line_114[905], line_113[903], line_112[901], line_111[899], line_110[897], line_109[895], line_108[893], line_107[891], line_106[889], line_105[887], line_104[885], line_103[883], line_102[881], line_101[879], line_100[877], line_99[875], line_98[873], line_97[871], line_96[869], line_95[867], line_94[865], line_93[863], line_92[861], line_91[859], line_90[857], line_89[855], line_88[853], line_87[851], line_86[849], line_85[847], line_84[845], line_83[843], line_82[841], line_81[839], line_80[837], line_79[835], line_78[833], line_77[831], line_76[829], line_75[827], line_74[825], line_73[823], line_72[821], line_71[819], line_70[817], line_69[815], line_68[813], line_67[811], line_66[809], line_65[807], line_64[805], line_63[803], line_62[801], line_61[799], line_60[797], line_59[795], line_58[793], line_57[791], line_56[789], line_55[787], line_54[785], line_53[783], line_52[781], line_51[779], line_50[777], line_49[775], line_48[773], line_47[771], line_46[769], line_45[767], line_44[765], line_43[763], line_42[761], line_41[759], line_40[757], line_39[755], line_38[753], line_37[751], line_36[749], line_35[747], line_34[745], line_33[743], line_32[741], line_31[739], line_30[737], line_29[735], line_28[733], line_27[731], line_26[729], line_25[727], line_24[725], line_23[723], line_22[721], line_21[719], line_20[717], line_19[715], line_18[713], line_17[711], line_16[709], line_15[707], line_14[705], line_13[703], line_12[701], line_11[699], line_10[697], line_9[695], line_8[693], line_7[691], line_6[689], line_5[687], line_4[685], line_3[683], line_2[681], line_1[679] };
assign col_934 = {line_128[934], line_127[932], line_126[930], line_125[928], line_124[926], line_123[924], line_122[922], line_121[920], line_120[918], line_119[916], line_118[914], line_117[912], line_116[910], line_115[908], line_114[906], line_113[904], line_112[902], line_111[900], line_110[898], line_109[896], line_108[894], line_107[892], line_106[890], line_105[888], line_104[886], line_103[884], line_102[882], line_101[880], line_100[878], line_99[876], line_98[874], line_97[872], line_96[870], line_95[868], line_94[866], line_93[864], line_92[862], line_91[860], line_90[858], line_89[856], line_88[854], line_87[852], line_86[850], line_85[848], line_84[846], line_83[844], line_82[842], line_81[840], line_80[838], line_79[836], line_78[834], line_77[832], line_76[830], line_75[828], line_74[826], line_73[824], line_72[822], line_71[820], line_70[818], line_69[816], line_68[814], line_67[812], line_66[810], line_65[808], line_64[806], line_63[804], line_62[802], line_61[800], line_60[798], line_59[796], line_58[794], line_57[792], line_56[790], line_55[788], line_54[786], line_53[784], line_52[782], line_51[780], line_50[778], line_49[776], line_48[774], line_47[772], line_46[770], line_45[768], line_44[766], line_43[764], line_42[762], line_41[760], line_40[758], line_39[756], line_38[754], line_37[752], line_36[750], line_35[748], line_34[746], line_33[744], line_32[742], line_31[740], line_30[738], line_29[736], line_28[734], line_27[732], line_26[730], line_25[728], line_24[726], line_23[724], line_22[722], line_21[720], line_20[718], line_19[716], line_18[714], line_17[712], line_16[710], line_15[708], line_14[706], line_13[704], line_12[702], line_11[700], line_10[698], line_9[696], line_8[694], line_7[692], line_6[690], line_5[688], line_4[686], line_3[684], line_2[682], line_1[680] };
assign col_935 = {line_128[935], line_127[933], line_126[931], line_125[929], line_124[927], line_123[925], line_122[923], line_121[921], line_120[919], line_119[917], line_118[915], line_117[913], line_116[911], line_115[909], line_114[907], line_113[905], line_112[903], line_111[901], line_110[899], line_109[897], line_108[895], line_107[893], line_106[891], line_105[889], line_104[887], line_103[885], line_102[883], line_101[881], line_100[879], line_99[877], line_98[875], line_97[873], line_96[871], line_95[869], line_94[867], line_93[865], line_92[863], line_91[861], line_90[859], line_89[857], line_88[855], line_87[853], line_86[851], line_85[849], line_84[847], line_83[845], line_82[843], line_81[841], line_80[839], line_79[837], line_78[835], line_77[833], line_76[831], line_75[829], line_74[827], line_73[825], line_72[823], line_71[821], line_70[819], line_69[817], line_68[815], line_67[813], line_66[811], line_65[809], line_64[807], line_63[805], line_62[803], line_61[801], line_60[799], line_59[797], line_58[795], line_57[793], line_56[791], line_55[789], line_54[787], line_53[785], line_52[783], line_51[781], line_50[779], line_49[777], line_48[775], line_47[773], line_46[771], line_45[769], line_44[767], line_43[765], line_42[763], line_41[761], line_40[759], line_39[757], line_38[755], line_37[753], line_36[751], line_35[749], line_34[747], line_33[745], line_32[743], line_31[741], line_30[739], line_29[737], line_28[735], line_27[733], line_26[731], line_25[729], line_24[727], line_23[725], line_22[723], line_21[721], line_20[719], line_19[717], line_18[715], line_17[713], line_16[711], line_15[709], line_14[707], line_13[705], line_12[703], line_11[701], line_10[699], line_9[697], line_8[695], line_7[693], line_6[691], line_5[689], line_4[687], line_3[685], line_2[683], line_1[681] };
assign col_936 = {line_128[936], line_127[934], line_126[932], line_125[930], line_124[928], line_123[926], line_122[924], line_121[922], line_120[920], line_119[918], line_118[916], line_117[914], line_116[912], line_115[910], line_114[908], line_113[906], line_112[904], line_111[902], line_110[900], line_109[898], line_108[896], line_107[894], line_106[892], line_105[890], line_104[888], line_103[886], line_102[884], line_101[882], line_100[880], line_99[878], line_98[876], line_97[874], line_96[872], line_95[870], line_94[868], line_93[866], line_92[864], line_91[862], line_90[860], line_89[858], line_88[856], line_87[854], line_86[852], line_85[850], line_84[848], line_83[846], line_82[844], line_81[842], line_80[840], line_79[838], line_78[836], line_77[834], line_76[832], line_75[830], line_74[828], line_73[826], line_72[824], line_71[822], line_70[820], line_69[818], line_68[816], line_67[814], line_66[812], line_65[810], line_64[808], line_63[806], line_62[804], line_61[802], line_60[800], line_59[798], line_58[796], line_57[794], line_56[792], line_55[790], line_54[788], line_53[786], line_52[784], line_51[782], line_50[780], line_49[778], line_48[776], line_47[774], line_46[772], line_45[770], line_44[768], line_43[766], line_42[764], line_41[762], line_40[760], line_39[758], line_38[756], line_37[754], line_36[752], line_35[750], line_34[748], line_33[746], line_32[744], line_31[742], line_30[740], line_29[738], line_28[736], line_27[734], line_26[732], line_25[730], line_24[728], line_23[726], line_22[724], line_21[722], line_20[720], line_19[718], line_18[716], line_17[714], line_16[712], line_15[710], line_14[708], line_13[706], line_12[704], line_11[702], line_10[700], line_9[698], line_8[696], line_7[694], line_6[692], line_5[690], line_4[688], line_3[686], line_2[684], line_1[682] };
assign col_937 = {line_128[937], line_127[935], line_126[933], line_125[931], line_124[929], line_123[927], line_122[925], line_121[923], line_120[921], line_119[919], line_118[917], line_117[915], line_116[913], line_115[911], line_114[909], line_113[907], line_112[905], line_111[903], line_110[901], line_109[899], line_108[897], line_107[895], line_106[893], line_105[891], line_104[889], line_103[887], line_102[885], line_101[883], line_100[881], line_99[879], line_98[877], line_97[875], line_96[873], line_95[871], line_94[869], line_93[867], line_92[865], line_91[863], line_90[861], line_89[859], line_88[857], line_87[855], line_86[853], line_85[851], line_84[849], line_83[847], line_82[845], line_81[843], line_80[841], line_79[839], line_78[837], line_77[835], line_76[833], line_75[831], line_74[829], line_73[827], line_72[825], line_71[823], line_70[821], line_69[819], line_68[817], line_67[815], line_66[813], line_65[811], line_64[809], line_63[807], line_62[805], line_61[803], line_60[801], line_59[799], line_58[797], line_57[795], line_56[793], line_55[791], line_54[789], line_53[787], line_52[785], line_51[783], line_50[781], line_49[779], line_48[777], line_47[775], line_46[773], line_45[771], line_44[769], line_43[767], line_42[765], line_41[763], line_40[761], line_39[759], line_38[757], line_37[755], line_36[753], line_35[751], line_34[749], line_33[747], line_32[745], line_31[743], line_30[741], line_29[739], line_28[737], line_27[735], line_26[733], line_25[731], line_24[729], line_23[727], line_22[725], line_21[723], line_20[721], line_19[719], line_18[717], line_17[715], line_16[713], line_15[711], line_14[709], line_13[707], line_12[705], line_11[703], line_10[701], line_9[699], line_8[697], line_7[695], line_6[693], line_5[691], line_4[689], line_3[687], line_2[685], line_1[683] };
assign col_938 = {line_128[938], line_127[936], line_126[934], line_125[932], line_124[930], line_123[928], line_122[926], line_121[924], line_120[922], line_119[920], line_118[918], line_117[916], line_116[914], line_115[912], line_114[910], line_113[908], line_112[906], line_111[904], line_110[902], line_109[900], line_108[898], line_107[896], line_106[894], line_105[892], line_104[890], line_103[888], line_102[886], line_101[884], line_100[882], line_99[880], line_98[878], line_97[876], line_96[874], line_95[872], line_94[870], line_93[868], line_92[866], line_91[864], line_90[862], line_89[860], line_88[858], line_87[856], line_86[854], line_85[852], line_84[850], line_83[848], line_82[846], line_81[844], line_80[842], line_79[840], line_78[838], line_77[836], line_76[834], line_75[832], line_74[830], line_73[828], line_72[826], line_71[824], line_70[822], line_69[820], line_68[818], line_67[816], line_66[814], line_65[812], line_64[810], line_63[808], line_62[806], line_61[804], line_60[802], line_59[800], line_58[798], line_57[796], line_56[794], line_55[792], line_54[790], line_53[788], line_52[786], line_51[784], line_50[782], line_49[780], line_48[778], line_47[776], line_46[774], line_45[772], line_44[770], line_43[768], line_42[766], line_41[764], line_40[762], line_39[760], line_38[758], line_37[756], line_36[754], line_35[752], line_34[750], line_33[748], line_32[746], line_31[744], line_30[742], line_29[740], line_28[738], line_27[736], line_26[734], line_25[732], line_24[730], line_23[728], line_22[726], line_21[724], line_20[722], line_19[720], line_18[718], line_17[716], line_16[714], line_15[712], line_14[710], line_13[708], line_12[706], line_11[704], line_10[702], line_9[700], line_8[698], line_7[696], line_6[694], line_5[692], line_4[690], line_3[688], line_2[686], line_1[684] };
assign col_939 = {line_128[939], line_127[937], line_126[935], line_125[933], line_124[931], line_123[929], line_122[927], line_121[925], line_120[923], line_119[921], line_118[919], line_117[917], line_116[915], line_115[913], line_114[911], line_113[909], line_112[907], line_111[905], line_110[903], line_109[901], line_108[899], line_107[897], line_106[895], line_105[893], line_104[891], line_103[889], line_102[887], line_101[885], line_100[883], line_99[881], line_98[879], line_97[877], line_96[875], line_95[873], line_94[871], line_93[869], line_92[867], line_91[865], line_90[863], line_89[861], line_88[859], line_87[857], line_86[855], line_85[853], line_84[851], line_83[849], line_82[847], line_81[845], line_80[843], line_79[841], line_78[839], line_77[837], line_76[835], line_75[833], line_74[831], line_73[829], line_72[827], line_71[825], line_70[823], line_69[821], line_68[819], line_67[817], line_66[815], line_65[813], line_64[811], line_63[809], line_62[807], line_61[805], line_60[803], line_59[801], line_58[799], line_57[797], line_56[795], line_55[793], line_54[791], line_53[789], line_52[787], line_51[785], line_50[783], line_49[781], line_48[779], line_47[777], line_46[775], line_45[773], line_44[771], line_43[769], line_42[767], line_41[765], line_40[763], line_39[761], line_38[759], line_37[757], line_36[755], line_35[753], line_34[751], line_33[749], line_32[747], line_31[745], line_30[743], line_29[741], line_28[739], line_27[737], line_26[735], line_25[733], line_24[731], line_23[729], line_22[727], line_21[725], line_20[723], line_19[721], line_18[719], line_17[717], line_16[715], line_15[713], line_14[711], line_13[709], line_12[707], line_11[705], line_10[703], line_9[701], line_8[699], line_7[697], line_6[695], line_5[693], line_4[691], line_3[689], line_2[687], line_1[685] };
assign col_940 = {line_128[940], line_127[938], line_126[936], line_125[934], line_124[932], line_123[930], line_122[928], line_121[926], line_120[924], line_119[922], line_118[920], line_117[918], line_116[916], line_115[914], line_114[912], line_113[910], line_112[908], line_111[906], line_110[904], line_109[902], line_108[900], line_107[898], line_106[896], line_105[894], line_104[892], line_103[890], line_102[888], line_101[886], line_100[884], line_99[882], line_98[880], line_97[878], line_96[876], line_95[874], line_94[872], line_93[870], line_92[868], line_91[866], line_90[864], line_89[862], line_88[860], line_87[858], line_86[856], line_85[854], line_84[852], line_83[850], line_82[848], line_81[846], line_80[844], line_79[842], line_78[840], line_77[838], line_76[836], line_75[834], line_74[832], line_73[830], line_72[828], line_71[826], line_70[824], line_69[822], line_68[820], line_67[818], line_66[816], line_65[814], line_64[812], line_63[810], line_62[808], line_61[806], line_60[804], line_59[802], line_58[800], line_57[798], line_56[796], line_55[794], line_54[792], line_53[790], line_52[788], line_51[786], line_50[784], line_49[782], line_48[780], line_47[778], line_46[776], line_45[774], line_44[772], line_43[770], line_42[768], line_41[766], line_40[764], line_39[762], line_38[760], line_37[758], line_36[756], line_35[754], line_34[752], line_33[750], line_32[748], line_31[746], line_30[744], line_29[742], line_28[740], line_27[738], line_26[736], line_25[734], line_24[732], line_23[730], line_22[728], line_21[726], line_20[724], line_19[722], line_18[720], line_17[718], line_16[716], line_15[714], line_14[712], line_13[710], line_12[708], line_11[706], line_10[704], line_9[702], line_8[700], line_7[698], line_6[696], line_5[694], line_4[692], line_3[690], line_2[688], line_1[686] };
assign col_941 = {line_128[941], line_127[939], line_126[937], line_125[935], line_124[933], line_123[931], line_122[929], line_121[927], line_120[925], line_119[923], line_118[921], line_117[919], line_116[917], line_115[915], line_114[913], line_113[911], line_112[909], line_111[907], line_110[905], line_109[903], line_108[901], line_107[899], line_106[897], line_105[895], line_104[893], line_103[891], line_102[889], line_101[887], line_100[885], line_99[883], line_98[881], line_97[879], line_96[877], line_95[875], line_94[873], line_93[871], line_92[869], line_91[867], line_90[865], line_89[863], line_88[861], line_87[859], line_86[857], line_85[855], line_84[853], line_83[851], line_82[849], line_81[847], line_80[845], line_79[843], line_78[841], line_77[839], line_76[837], line_75[835], line_74[833], line_73[831], line_72[829], line_71[827], line_70[825], line_69[823], line_68[821], line_67[819], line_66[817], line_65[815], line_64[813], line_63[811], line_62[809], line_61[807], line_60[805], line_59[803], line_58[801], line_57[799], line_56[797], line_55[795], line_54[793], line_53[791], line_52[789], line_51[787], line_50[785], line_49[783], line_48[781], line_47[779], line_46[777], line_45[775], line_44[773], line_43[771], line_42[769], line_41[767], line_40[765], line_39[763], line_38[761], line_37[759], line_36[757], line_35[755], line_34[753], line_33[751], line_32[749], line_31[747], line_30[745], line_29[743], line_28[741], line_27[739], line_26[737], line_25[735], line_24[733], line_23[731], line_22[729], line_21[727], line_20[725], line_19[723], line_18[721], line_17[719], line_16[717], line_15[715], line_14[713], line_13[711], line_12[709], line_11[707], line_10[705], line_9[703], line_8[701], line_7[699], line_6[697], line_5[695], line_4[693], line_3[691], line_2[689], line_1[687] };
assign col_942 = {line_128[942], line_127[940], line_126[938], line_125[936], line_124[934], line_123[932], line_122[930], line_121[928], line_120[926], line_119[924], line_118[922], line_117[920], line_116[918], line_115[916], line_114[914], line_113[912], line_112[910], line_111[908], line_110[906], line_109[904], line_108[902], line_107[900], line_106[898], line_105[896], line_104[894], line_103[892], line_102[890], line_101[888], line_100[886], line_99[884], line_98[882], line_97[880], line_96[878], line_95[876], line_94[874], line_93[872], line_92[870], line_91[868], line_90[866], line_89[864], line_88[862], line_87[860], line_86[858], line_85[856], line_84[854], line_83[852], line_82[850], line_81[848], line_80[846], line_79[844], line_78[842], line_77[840], line_76[838], line_75[836], line_74[834], line_73[832], line_72[830], line_71[828], line_70[826], line_69[824], line_68[822], line_67[820], line_66[818], line_65[816], line_64[814], line_63[812], line_62[810], line_61[808], line_60[806], line_59[804], line_58[802], line_57[800], line_56[798], line_55[796], line_54[794], line_53[792], line_52[790], line_51[788], line_50[786], line_49[784], line_48[782], line_47[780], line_46[778], line_45[776], line_44[774], line_43[772], line_42[770], line_41[768], line_40[766], line_39[764], line_38[762], line_37[760], line_36[758], line_35[756], line_34[754], line_33[752], line_32[750], line_31[748], line_30[746], line_29[744], line_28[742], line_27[740], line_26[738], line_25[736], line_24[734], line_23[732], line_22[730], line_21[728], line_20[726], line_19[724], line_18[722], line_17[720], line_16[718], line_15[716], line_14[714], line_13[712], line_12[710], line_11[708], line_10[706], line_9[704], line_8[702], line_7[700], line_6[698], line_5[696], line_4[694], line_3[692], line_2[690], line_1[688] };
assign col_943 = {line_128[943], line_127[941], line_126[939], line_125[937], line_124[935], line_123[933], line_122[931], line_121[929], line_120[927], line_119[925], line_118[923], line_117[921], line_116[919], line_115[917], line_114[915], line_113[913], line_112[911], line_111[909], line_110[907], line_109[905], line_108[903], line_107[901], line_106[899], line_105[897], line_104[895], line_103[893], line_102[891], line_101[889], line_100[887], line_99[885], line_98[883], line_97[881], line_96[879], line_95[877], line_94[875], line_93[873], line_92[871], line_91[869], line_90[867], line_89[865], line_88[863], line_87[861], line_86[859], line_85[857], line_84[855], line_83[853], line_82[851], line_81[849], line_80[847], line_79[845], line_78[843], line_77[841], line_76[839], line_75[837], line_74[835], line_73[833], line_72[831], line_71[829], line_70[827], line_69[825], line_68[823], line_67[821], line_66[819], line_65[817], line_64[815], line_63[813], line_62[811], line_61[809], line_60[807], line_59[805], line_58[803], line_57[801], line_56[799], line_55[797], line_54[795], line_53[793], line_52[791], line_51[789], line_50[787], line_49[785], line_48[783], line_47[781], line_46[779], line_45[777], line_44[775], line_43[773], line_42[771], line_41[769], line_40[767], line_39[765], line_38[763], line_37[761], line_36[759], line_35[757], line_34[755], line_33[753], line_32[751], line_31[749], line_30[747], line_29[745], line_28[743], line_27[741], line_26[739], line_25[737], line_24[735], line_23[733], line_22[731], line_21[729], line_20[727], line_19[725], line_18[723], line_17[721], line_16[719], line_15[717], line_14[715], line_13[713], line_12[711], line_11[709], line_10[707], line_9[705], line_8[703], line_7[701], line_6[699], line_5[697], line_4[695], line_3[693], line_2[691], line_1[689] };
assign col_944 = {line_128[944], line_127[942], line_126[940], line_125[938], line_124[936], line_123[934], line_122[932], line_121[930], line_120[928], line_119[926], line_118[924], line_117[922], line_116[920], line_115[918], line_114[916], line_113[914], line_112[912], line_111[910], line_110[908], line_109[906], line_108[904], line_107[902], line_106[900], line_105[898], line_104[896], line_103[894], line_102[892], line_101[890], line_100[888], line_99[886], line_98[884], line_97[882], line_96[880], line_95[878], line_94[876], line_93[874], line_92[872], line_91[870], line_90[868], line_89[866], line_88[864], line_87[862], line_86[860], line_85[858], line_84[856], line_83[854], line_82[852], line_81[850], line_80[848], line_79[846], line_78[844], line_77[842], line_76[840], line_75[838], line_74[836], line_73[834], line_72[832], line_71[830], line_70[828], line_69[826], line_68[824], line_67[822], line_66[820], line_65[818], line_64[816], line_63[814], line_62[812], line_61[810], line_60[808], line_59[806], line_58[804], line_57[802], line_56[800], line_55[798], line_54[796], line_53[794], line_52[792], line_51[790], line_50[788], line_49[786], line_48[784], line_47[782], line_46[780], line_45[778], line_44[776], line_43[774], line_42[772], line_41[770], line_40[768], line_39[766], line_38[764], line_37[762], line_36[760], line_35[758], line_34[756], line_33[754], line_32[752], line_31[750], line_30[748], line_29[746], line_28[744], line_27[742], line_26[740], line_25[738], line_24[736], line_23[734], line_22[732], line_21[730], line_20[728], line_19[726], line_18[724], line_17[722], line_16[720], line_15[718], line_14[716], line_13[714], line_12[712], line_11[710], line_10[708], line_9[706], line_8[704], line_7[702], line_6[700], line_5[698], line_4[696], line_3[694], line_2[692], line_1[690] };
assign col_945 = {line_128[945], line_127[943], line_126[941], line_125[939], line_124[937], line_123[935], line_122[933], line_121[931], line_120[929], line_119[927], line_118[925], line_117[923], line_116[921], line_115[919], line_114[917], line_113[915], line_112[913], line_111[911], line_110[909], line_109[907], line_108[905], line_107[903], line_106[901], line_105[899], line_104[897], line_103[895], line_102[893], line_101[891], line_100[889], line_99[887], line_98[885], line_97[883], line_96[881], line_95[879], line_94[877], line_93[875], line_92[873], line_91[871], line_90[869], line_89[867], line_88[865], line_87[863], line_86[861], line_85[859], line_84[857], line_83[855], line_82[853], line_81[851], line_80[849], line_79[847], line_78[845], line_77[843], line_76[841], line_75[839], line_74[837], line_73[835], line_72[833], line_71[831], line_70[829], line_69[827], line_68[825], line_67[823], line_66[821], line_65[819], line_64[817], line_63[815], line_62[813], line_61[811], line_60[809], line_59[807], line_58[805], line_57[803], line_56[801], line_55[799], line_54[797], line_53[795], line_52[793], line_51[791], line_50[789], line_49[787], line_48[785], line_47[783], line_46[781], line_45[779], line_44[777], line_43[775], line_42[773], line_41[771], line_40[769], line_39[767], line_38[765], line_37[763], line_36[761], line_35[759], line_34[757], line_33[755], line_32[753], line_31[751], line_30[749], line_29[747], line_28[745], line_27[743], line_26[741], line_25[739], line_24[737], line_23[735], line_22[733], line_21[731], line_20[729], line_19[727], line_18[725], line_17[723], line_16[721], line_15[719], line_14[717], line_13[715], line_12[713], line_11[711], line_10[709], line_9[707], line_8[705], line_7[703], line_6[701], line_5[699], line_4[697], line_3[695], line_2[693], line_1[691] };
assign col_946 = {line_128[946], line_127[944], line_126[942], line_125[940], line_124[938], line_123[936], line_122[934], line_121[932], line_120[930], line_119[928], line_118[926], line_117[924], line_116[922], line_115[920], line_114[918], line_113[916], line_112[914], line_111[912], line_110[910], line_109[908], line_108[906], line_107[904], line_106[902], line_105[900], line_104[898], line_103[896], line_102[894], line_101[892], line_100[890], line_99[888], line_98[886], line_97[884], line_96[882], line_95[880], line_94[878], line_93[876], line_92[874], line_91[872], line_90[870], line_89[868], line_88[866], line_87[864], line_86[862], line_85[860], line_84[858], line_83[856], line_82[854], line_81[852], line_80[850], line_79[848], line_78[846], line_77[844], line_76[842], line_75[840], line_74[838], line_73[836], line_72[834], line_71[832], line_70[830], line_69[828], line_68[826], line_67[824], line_66[822], line_65[820], line_64[818], line_63[816], line_62[814], line_61[812], line_60[810], line_59[808], line_58[806], line_57[804], line_56[802], line_55[800], line_54[798], line_53[796], line_52[794], line_51[792], line_50[790], line_49[788], line_48[786], line_47[784], line_46[782], line_45[780], line_44[778], line_43[776], line_42[774], line_41[772], line_40[770], line_39[768], line_38[766], line_37[764], line_36[762], line_35[760], line_34[758], line_33[756], line_32[754], line_31[752], line_30[750], line_29[748], line_28[746], line_27[744], line_26[742], line_25[740], line_24[738], line_23[736], line_22[734], line_21[732], line_20[730], line_19[728], line_18[726], line_17[724], line_16[722], line_15[720], line_14[718], line_13[716], line_12[714], line_11[712], line_10[710], line_9[708], line_8[706], line_7[704], line_6[702], line_5[700], line_4[698], line_3[696], line_2[694], line_1[692] };
assign col_947 = {line_128[947], line_127[945], line_126[943], line_125[941], line_124[939], line_123[937], line_122[935], line_121[933], line_120[931], line_119[929], line_118[927], line_117[925], line_116[923], line_115[921], line_114[919], line_113[917], line_112[915], line_111[913], line_110[911], line_109[909], line_108[907], line_107[905], line_106[903], line_105[901], line_104[899], line_103[897], line_102[895], line_101[893], line_100[891], line_99[889], line_98[887], line_97[885], line_96[883], line_95[881], line_94[879], line_93[877], line_92[875], line_91[873], line_90[871], line_89[869], line_88[867], line_87[865], line_86[863], line_85[861], line_84[859], line_83[857], line_82[855], line_81[853], line_80[851], line_79[849], line_78[847], line_77[845], line_76[843], line_75[841], line_74[839], line_73[837], line_72[835], line_71[833], line_70[831], line_69[829], line_68[827], line_67[825], line_66[823], line_65[821], line_64[819], line_63[817], line_62[815], line_61[813], line_60[811], line_59[809], line_58[807], line_57[805], line_56[803], line_55[801], line_54[799], line_53[797], line_52[795], line_51[793], line_50[791], line_49[789], line_48[787], line_47[785], line_46[783], line_45[781], line_44[779], line_43[777], line_42[775], line_41[773], line_40[771], line_39[769], line_38[767], line_37[765], line_36[763], line_35[761], line_34[759], line_33[757], line_32[755], line_31[753], line_30[751], line_29[749], line_28[747], line_27[745], line_26[743], line_25[741], line_24[739], line_23[737], line_22[735], line_21[733], line_20[731], line_19[729], line_18[727], line_17[725], line_16[723], line_15[721], line_14[719], line_13[717], line_12[715], line_11[713], line_10[711], line_9[709], line_8[707], line_7[705], line_6[703], line_5[701], line_4[699], line_3[697], line_2[695], line_1[693] };
assign col_948 = {line_128[948], line_127[946], line_126[944], line_125[942], line_124[940], line_123[938], line_122[936], line_121[934], line_120[932], line_119[930], line_118[928], line_117[926], line_116[924], line_115[922], line_114[920], line_113[918], line_112[916], line_111[914], line_110[912], line_109[910], line_108[908], line_107[906], line_106[904], line_105[902], line_104[900], line_103[898], line_102[896], line_101[894], line_100[892], line_99[890], line_98[888], line_97[886], line_96[884], line_95[882], line_94[880], line_93[878], line_92[876], line_91[874], line_90[872], line_89[870], line_88[868], line_87[866], line_86[864], line_85[862], line_84[860], line_83[858], line_82[856], line_81[854], line_80[852], line_79[850], line_78[848], line_77[846], line_76[844], line_75[842], line_74[840], line_73[838], line_72[836], line_71[834], line_70[832], line_69[830], line_68[828], line_67[826], line_66[824], line_65[822], line_64[820], line_63[818], line_62[816], line_61[814], line_60[812], line_59[810], line_58[808], line_57[806], line_56[804], line_55[802], line_54[800], line_53[798], line_52[796], line_51[794], line_50[792], line_49[790], line_48[788], line_47[786], line_46[784], line_45[782], line_44[780], line_43[778], line_42[776], line_41[774], line_40[772], line_39[770], line_38[768], line_37[766], line_36[764], line_35[762], line_34[760], line_33[758], line_32[756], line_31[754], line_30[752], line_29[750], line_28[748], line_27[746], line_26[744], line_25[742], line_24[740], line_23[738], line_22[736], line_21[734], line_20[732], line_19[730], line_18[728], line_17[726], line_16[724], line_15[722], line_14[720], line_13[718], line_12[716], line_11[714], line_10[712], line_9[710], line_8[708], line_7[706], line_6[704], line_5[702], line_4[700], line_3[698], line_2[696], line_1[694] };
assign col_949 = {line_128[949], line_127[947], line_126[945], line_125[943], line_124[941], line_123[939], line_122[937], line_121[935], line_120[933], line_119[931], line_118[929], line_117[927], line_116[925], line_115[923], line_114[921], line_113[919], line_112[917], line_111[915], line_110[913], line_109[911], line_108[909], line_107[907], line_106[905], line_105[903], line_104[901], line_103[899], line_102[897], line_101[895], line_100[893], line_99[891], line_98[889], line_97[887], line_96[885], line_95[883], line_94[881], line_93[879], line_92[877], line_91[875], line_90[873], line_89[871], line_88[869], line_87[867], line_86[865], line_85[863], line_84[861], line_83[859], line_82[857], line_81[855], line_80[853], line_79[851], line_78[849], line_77[847], line_76[845], line_75[843], line_74[841], line_73[839], line_72[837], line_71[835], line_70[833], line_69[831], line_68[829], line_67[827], line_66[825], line_65[823], line_64[821], line_63[819], line_62[817], line_61[815], line_60[813], line_59[811], line_58[809], line_57[807], line_56[805], line_55[803], line_54[801], line_53[799], line_52[797], line_51[795], line_50[793], line_49[791], line_48[789], line_47[787], line_46[785], line_45[783], line_44[781], line_43[779], line_42[777], line_41[775], line_40[773], line_39[771], line_38[769], line_37[767], line_36[765], line_35[763], line_34[761], line_33[759], line_32[757], line_31[755], line_30[753], line_29[751], line_28[749], line_27[747], line_26[745], line_25[743], line_24[741], line_23[739], line_22[737], line_21[735], line_20[733], line_19[731], line_18[729], line_17[727], line_16[725], line_15[723], line_14[721], line_13[719], line_12[717], line_11[715], line_10[713], line_9[711], line_8[709], line_7[707], line_6[705], line_5[703], line_4[701], line_3[699], line_2[697], line_1[695] };
assign col_950 = {line_128[950], line_127[948], line_126[946], line_125[944], line_124[942], line_123[940], line_122[938], line_121[936], line_120[934], line_119[932], line_118[930], line_117[928], line_116[926], line_115[924], line_114[922], line_113[920], line_112[918], line_111[916], line_110[914], line_109[912], line_108[910], line_107[908], line_106[906], line_105[904], line_104[902], line_103[900], line_102[898], line_101[896], line_100[894], line_99[892], line_98[890], line_97[888], line_96[886], line_95[884], line_94[882], line_93[880], line_92[878], line_91[876], line_90[874], line_89[872], line_88[870], line_87[868], line_86[866], line_85[864], line_84[862], line_83[860], line_82[858], line_81[856], line_80[854], line_79[852], line_78[850], line_77[848], line_76[846], line_75[844], line_74[842], line_73[840], line_72[838], line_71[836], line_70[834], line_69[832], line_68[830], line_67[828], line_66[826], line_65[824], line_64[822], line_63[820], line_62[818], line_61[816], line_60[814], line_59[812], line_58[810], line_57[808], line_56[806], line_55[804], line_54[802], line_53[800], line_52[798], line_51[796], line_50[794], line_49[792], line_48[790], line_47[788], line_46[786], line_45[784], line_44[782], line_43[780], line_42[778], line_41[776], line_40[774], line_39[772], line_38[770], line_37[768], line_36[766], line_35[764], line_34[762], line_33[760], line_32[758], line_31[756], line_30[754], line_29[752], line_28[750], line_27[748], line_26[746], line_25[744], line_24[742], line_23[740], line_22[738], line_21[736], line_20[734], line_19[732], line_18[730], line_17[728], line_16[726], line_15[724], line_14[722], line_13[720], line_12[718], line_11[716], line_10[714], line_9[712], line_8[710], line_7[708], line_6[706], line_5[704], line_4[702], line_3[700], line_2[698], line_1[696] };
assign col_951 = {line_128[951], line_127[949], line_126[947], line_125[945], line_124[943], line_123[941], line_122[939], line_121[937], line_120[935], line_119[933], line_118[931], line_117[929], line_116[927], line_115[925], line_114[923], line_113[921], line_112[919], line_111[917], line_110[915], line_109[913], line_108[911], line_107[909], line_106[907], line_105[905], line_104[903], line_103[901], line_102[899], line_101[897], line_100[895], line_99[893], line_98[891], line_97[889], line_96[887], line_95[885], line_94[883], line_93[881], line_92[879], line_91[877], line_90[875], line_89[873], line_88[871], line_87[869], line_86[867], line_85[865], line_84[863], line_83[861], line_82[859], line_81[857], line_80[855], line_79[853], line_78[851], line_77[849], line_76[847], line_75[845], line_74[843], line_73[841], line_72[839], line_71[837], line_70[835], line_69[833], line_68[831], line_67[829], line_66[827], line_65[825], line_64[823], line_63[821], line_62[819], line_61[817], line_60[815], line_59[813], line_58[811], line_57[809], line_56[807], line_55[805], line_54[803], line_53[801], line_52[799], line_51[797], line_50[795], line_49[793], line_48[791], line_47[789], line_46[787], line_45[785], line_44[783], line_43[781], line_42[779], line_41[777], line_40[775], line_39[773], line_38[771], line_37[769], line_36[767], line_35[765], line_34[763], line_33[761], line_32[759], line_31[757], line_30[755], line_29[753], line_28[751], line_27[749], line_26[747], line_25[745], line_24[743], line_23[741], line_22[739], line_21[737], line_20[735], line_19[733], line_18[731], line_17[729], line_16[727], line_15[725], line_14[723], line_13[721], line_12[719], line_11[717], line_10[715], line_9[713], line_8[711], line_7[709], line_6[707], line_5[705], line_4[703], line_3[701], line_2[699], line_1[697] };
assign col_952 = {line_128[952], line_127[950], line_126[948], line_125[946], line_124[944], line_123[942], line_122[940], line_121[938], line_120[936], line_119[934], line_118[932], line_117[930], line_116[928], line_115[926], line_114[924], line_113[922], line_112[920], line_111[918], line_110[916], line_109[914], line_108[912], line_107[910], line_106[908], line_105[906], line_104[904], line_103[902], line_102[900], line_101[898], line_100[896], line_99[894], line_98[892], line_97[890], line_96[888], line_95[886], line_94[884], line_93[882], line_92[880], line_91[878], line_90[876], line_89[874], line_88[872], line_87[870], line_86[868], line_85[866], line_84[864], line_83[862], line_82[860], line_81[858], line_80[856], line_79[854], line_78[852], line_77[850], line_76[848], line_75[846], line_74[844], line_73[842], line_72[840], line_71[838], line_70[836], line_69[834], line_68[832], line_67[830], line_66[828], line_65[826], line_64[824], line_63[822], line_62[820], line_61[818], line_60[816], line_59[814], line_58[812], line_57[810], line_56[808], line_55[806], line_54[804], line_53[802], line_52[800], line_51[798], line_50[796], line_49[794], line_48[792], line_47[790], line_46[788], line_45[786], line_44[784], line_43[782], line_42[780], line_41[778], line_40[776], line_39[774], line_38[772], line_37[770], line_36[768], line_35[766], line_34[764], line_33[762], line_32[760], line_31[758], line_30[756], line_29[754], line_28[752], line_27[750], line_26[748], line_25[746], line_24[744], line_23[742], line_22[740], line_21[738], line_20[736], line_19[734], line_18[732], line_17[730], line_16[728], line_15[726], line_14[724], line_13[722], line_12[720], line_11[718], line_10[716], line_9[714], line_8[712], line_7[710], line_6[708], line_5[706], line_4[704], line_3[702], line_2[700], line_1[698] };
assign col_953 = {line_128[953], line_127[951], line_126[949], line_125[947], line_124[945], line_123[943], line_122[941], line_121[939], line_120[937], line_119[935], line_118[933], line_117[931], line_116[929], line_115[927], line_114[925], line_113[923], line_112[921], line_111[919], line_110[917], line_109[915], line_108[913], line_107[911], line_106[909], line_105[907], line_104[905], line_103[903], line_102[901], line_101[899], line_100[897], line_99[895], line_98[893], line_97[891], line_96[889], line_95[887], line_94[885], line_93[883], line_92[881], line_91[879], line_90[877], line_89[875], line_88[873], line_87[871], line_86[869], line_85[867], line_84[865], line_83[863], line_82[861], line_81[859], line_80[857], line_79[855], line_78[853], line_77[851], line_76[849], line_75[847], line_74[845], line_73[843], line_72[841], line_71[839], line_70[837], line_69[835], line_68[833], line_67[831], line_66[829], line_65[827], line_64[825], line_63[823], line_62[821], line_61[819], line_60[817], line_59[815], line_58[813], line_57[811], line_56[809], line_55[807], line_54[805], line_53[803], line_52[801], line_51[799], line_50[797], line_49[795], line_48[793], line_47[791], line_46[789], line_45[787], line_44[785], line_43[783], line_42[781], line_41[779], line_40[777], line_39[775], line_38[773], line_37[771], line_36[769], line_35[767], line_34[765], line_33[763], line_32[761], line_31[759], line_30[757], line_29[755], line_28[753], line_27[751], line_26[749], line_25[747], line_24[745], line_23[743], line_22[741], line_21[739], line_20[737], line_19[735], line_18[733], line_17[731], line_16[729], line_15[727], line_14[725], line_13[723], line_12[721], line_11[719], line_10[717], line_9[715], line_8[713], line_7[711], line_6[709], line_5[707], line_4[705], line_3[703], line_2[701], line_1[699] };
assign col_954 = {line_128[954], line_127[952], line_126[950], line_125[948], line_124[946], line_123[944], line_122[942], line_121[940], line_120[938], line_119[936], line_118[934], line_117[932], line_116[930], line_115[928], line_114[926], line_113[924], line_112[922], line_111[920], line_110[918], line_109[916], line_108[914], line_107[912], line_106[910], line_105[908], line_104[906], line_103[904], line_102[902], line_101[900], line_100[898], line_99[896], line_98[894], line_97[892], line_96[890], line_95[888], line_94[886], line_93[884], line_92[882], line_91[880], line_90[878], line_89[876], line_88[874], line_87[872], line_86[870], line_85[868], line_84[866], line_83[864], line_82[862], line_81[860], line_80[858], line_79[856], line_78[854], line_77[852], line_76[850], line_75[848], line_74[846], line_73[844], line_72[842], line_71[840], line_70[838], line_69[836], line_68[834], line_67[832], line_66[830], line_65[828], line_64[826], line_63[824], line_62[822], line_61[820], line_60[818], line_59[816], line_58[814], line_57[812], line_56[810], line_55[808], line_54[806], line_53[804], line_52[802], line_51[800], line_50[798], line_49[796], line_48[794], line_47[792], line_46[790], line_45[788], line_44[786], line_43[784], line_42[782], line_41[780], line_40[778], line_39[776], line_38[774], line_37[772], line_36[770], line_35[768], line_34[766], line_33[764], line_32[762], line_31[760], line_30[758], line_29[756], line_28[754], line_27[752], line_26[750], line_25[748], line_24[746], line_23[744], line_22[742], line_21[740], line_20[738], line_19[736], line_18[734], line_17[732], line_16[730], line_15[728], line_14[726], line_13[724], line_12[722], line_11[720], line_10[718], line_9[716], line_8[714], line_7[712], line_6[710], line_5[708], line_4[706], line_3[704], line_2[702], line_1[700] };
assign col_955 = {line_128[955], line_127[953], line_126[951], line_125[949], line_124[947], line_123[945], line_122[943], line_121[941], line_120[939], line_119[937], line_118[935], line_117[933], line_116[931], line_115[929], line_114[927], line_113[925], line_112[923], line_111[921], line_110[919], line_109[917], line_108[915], line_107[913], line_106[911], line_105[909], line_104[907], line_103[905], line_102[903], line_101[901], line_100[899], line_99[897], line_98[895], line_97[893], line_96[891], line_95[889], line_94[887], line_93[885], line_92[883], line_91[881], line_90[879], line_89[877], line_88[875], line_87[873], line_86[871], line_85[869], line_84[867], line_83[865], line_82[863], line_81[861], line_80[859], line_79[857], line_78[855], line_77[853], line_76[851], line_75[849], line_74[847], line_73[845], line_72[843], line_71[841], line_70[839], line_69[837], line_68[835], line_67[833], line_66[831], line_65[829], line_64[827], line_63[825], line_62[823], line_61[821], line_60[819], line_59[817], line_58[815], line_57[813], line_56[811], line_55[809], line_54[807], line_53[805], line_52[803], line_51[801], line_50[799], line_49[797], line_48[795], line_47[793], line_46[791], line_45[789], line_44[787], line_43[785], line_42[783], line_41[781], line_40[779], line_39[777], line_38[775], line_37[773], line_36[771], line_35[769], line_34[767], line_33[765], line_32[763], line_31[761], line_30[759], line_29[757], line_28[755], line_27[753], line_26[751], line_25[749], line_24[747], line_23[745], line_22[743], line_21[741], line_20[739], line_19[737], line_18[735], line_17[733], line_16[731], line_15[729], line_14[727], line_13[725], line_12[723], line_11[721], line_10[719], line_9[717], line_8[715], line_7[713], line_6[711], line_5[709], line_4[707], line_3[705], line_2[703], line_1[701] };
assign col_956 = {line_128[956], line_127[954], line_126[952], line_125[950], line_124[948], line_123[946], line_122[944], line_121[942], line_120[940], line_119[938], line_118[936], line_117[934], line_116[932], line_115[930], line_114[928], line_113[926], line_112[924], line_111[922], line_110[920], line_109[918], line_108[916], line_107[914], line_106[912], line_105[910], line_104[908], line_103[906], line_102[904], line_101[902], line_100[900], line_99[898], line_98[896], line_97[894], line_96[892], line_95[890], line_94[888], line_93[886], line_92[884], line_91[882], line_90[880], line_89[878], line_88[876], line_87[874], line_86[872], line_85[870], line_84[868], line_83[866], line_82[864], line_81[862], line_80[860], line_79[858], line_78[856], line_77[854], line_76[852], line_75[850], line_74[848], line_73[846], line_72[844], line_71[842], line_70[840], line_69[838], line_68[836], line_67[834], line_66[832], line_65[830], line_64[828], line_63[826], line_62[824], line_61[822], line_60[820], line_59[818], line_58[816], line_57[814], line_56[812], line_55[810], line_54[808], line_53[806], line_52[804], line_51[802], line_50[800], line_49[798], line_48[796], line_47[794], line_46[792], line_45[790], line_44[788], line_43[786], line_42[784], line_41[782], line_40[780], line_39[778], line_38[776], line_37[774], line_36[772], line_35[770], line_34[768], line_33[766], line_32[764], line_31[762], line_30[760], line_29[758], line_28[756], line_27[754], line_26[752], line_25[750], line_24[748], line_23[746], line_22[744], line_21[742], line_20[740], line_19[738], line_18[736], line_17[734], line_16[732], line_15[730], line_14[728], line_13[726], line_12[724], line_11[722], line_10[720], line_9[718], line_8[716], line_7[714], line_6[712], line_5[710], line_4[708], line_3[706], line_2[704], line_1[702] };
assign col_957 = {line_128[957], line_127[955], line_126[953], line_125[951], line_124[949], line_123[947], line_122[945], line_121[943], line_120[941], line_119[939], line_118[937], line_117[935], line_116[933], line_115[931], line_114[929], line_113[927], line_112[925], line_111[923], line_110[921], line_109[919], line_108[917], line_107[915], line_106[913], line_105[911], line_104[909], line_103[907], line_102[905], line_101[903], line_100[901], line_99[899], line_98[897], line_97[895], line_96[893], line_95[891], line_94[889], line_93[887], line_92[885], line_91[883], line_90[881], line_89[879], line_88[877], line_87[875], line_86[873], line_85[871], line_84[869], line_83[867], line_82[865], line_81[863], line_80[861], line_79[859], line_78[857], line_77[855], line_76[853], line_75[851], line_74[849], line_73[847], line_72[845], line_71[843], line_70[841], line_69[839], line_68[837], line_67[835], line_66[833], line_65[831], line_64[829], line_63[827], line_62[825], line_61[823], line_60[821], line_59[819], line_58[817], line_57[815], line_56[813], line_55[811], line_54[809], line_53[807], line_52[805], line_51[803], line_50[801], line_49[799], line_48[797], line_47[795], line_46[793], line_45[791], line_44[789], line_43[787], line_42[785], line_41[783], line_40[781], line_39[779], line_38[777], line_37[775], line_36[773], line_35[771], line_34[769], line_33[767], line_32[765], line_31[763], line_30[761], line_29[759], line_28[757], line_27[755], line_26[753], line_25[751], line_24[749], line_23[747], line_22[745], line_21[743], line_20[741], line_19[739], line_18[737], line_17[735], line_16[733], line_15[731], line_14[729], line_13[727], line_12[725], line_11[723], line_10[721], line_9[719], line_8[717], line_7[715], line_6[713], line_5[711], line_4[709], line_3[707], line_2[705], line_1[703] };
assign col_958 = {line_128[958], line_127[956], line_126[954], line_125[952], line_124[950], line_123[948], line_122[946], line_121[944], line_120[942], line_119[940], line_118[938], line_117[936], line_116[934], line_115[932], line_114[930], line_113[928], line_112[926], line_111[924], line_110[922], line_109[920], line_108[918], line_107[916], line_106[914], line_105[912], line_104[910], line_103[908], line_102[906], line_101[904], line_100[902], line_99[900], line_98[898], line_97[896], line_96[894], line_95[892], line_94[890], line_93[888], line_92[886], line_91[884], line_90[882], line_89[880], line_88[878], line_87[876], line_86[874], line_85[872], line_84[870], line_83[868], line_82[866], line_81[864], line_80[862], line_79[860], line_78[858], line_77[856], line_76[854], line_75[852], line_74[850], line_73[848], line_72[846], line_71[844], line_70[842], line_69[840], line_68[838], line_67[836], line_66[834], line_65[832], line_64[830], line_63[828], line_62[826], line_61[824], line_60[822], line_59[820], line_58[818], line_57[816], line_56[814], line_55[812], line_54[810], line_53[808], line_52[806], line_51[804], line_50[802], line_49[800], line_48[798], line_47[796], line_46[794], line_45[792], line_44[790], line_43[788], line_42[786], line_41[784], line_40[782], line_39[780], line_38[778], line_37[776], line_36[774], line_35[772], line_34[770], line_33[768], line_32[766], line_31[764], line_30[762], line_29[760], line_28[758], line_27[756], line_26[754], line_25[752], line_24[750], line_23[748], line_22[746], line_21[744], line_20[742], line_19[740], line_18[738], line_17[736], line_16[734], line_15[732], line_14[730], line_13[728], line_12[726], line_11[724], line_10[722], line_9[720], line_8[718], line_7[716], line_6[714], line_5[712], line_4[710], line_3[708], line_2[706], line_1[704] };
assign col_959 = {line_128[959], line_127[957], line_126[955], line_125[953], line_124[951], line_123[949], line_122[947], line_121[945], line_120[943], line_119[941], line_118[939], line_117[937], line_116[935], line_115[933], line_114[931], line_113[929], line_112[927], line_111[925], line_110[923], line_109[921], line_108[919], line_107[917], line_106[915], line_105[913], line_104[911], line_103[909], line_102[907], line_101[905], line_100[903], line_99[901], line_98[899], line_97[897], line_96[895], line_95[893], line_94[891], line_93[889], line_92[887], line_91[885], line_90[883], line_89[881], line_88[879], line_87[877], line_86[875], line_85[873], line_84[871], line_83[869], line_82[867], line_81[865], line_80[863], line_79[861], line_78[859], line_77[857], line_76[855], line_75[853], line_74[851], line_73[849], line_72[847], line_71[845], line_70[843], line_69[841], line_68[839], line_67[837], line_66[835], line_65[833], line_64[831], line_63[829], line_62[827], line_61[825], line_60[823], line_59[821], line_58[819], line_57[817], line_56[815], line_55[813], line_54[811], line_53[809], line_52[807], line_51[805], line_50[803], line_49[801], line_48[799], line_47[797], line_46[795], line_45[793], line_44[791], line_43[789], line_42[787], line_41[785], line_40[783], line_39[781], line_38[779], line_37[777], line_36[775], line_35[773], line_34[771], line_33[769], line_32[767], line_31[765], line_30[763], line_29[761], line_28[759], line_27[757], line_26[755], line_25[753], line_24[751], line_23[749], line_22[747], line_21[745], line_20[743], line_19[741], line_18[739], line_17[737], line_16[735], line_15[733], line_14[731], line_13[729], line_12[727], line_11[725], line_10[723], line_9[721], line_8[719], line_7[717], line_6[715], line_5[713], line_4[711], line_3[709], line_2[707], line_1[705] };
assign col_960 = {line_128[960], line_127[958], line_126[956], line_125[954], line_124[952], line_123[950], line_122[948], line_121[946], line_120[944], line_119[942], line_118[940], line_117[938], line_116[936], line_115[934], line_114[932], line_113[930], line_112[928], line_111[926], line_110[924], line_109[922], line_108[920], line_107[918], line_106[916], line_105[914], line_104[912], line_103[910], line_102[908], line_101[906], line_100[904], line_99[902], line_98[900], line_97[898], line_96[896], line_95[894], line_94[892], line_93[890], line_92[888], line_91[886], line_90[884], line_89[882], line_88[880], line_87[878], line_86[876], line_85[874], line_84[872], line_83[870], line_82[868], line_81[866], line_80[864], line_79[862], line_78[860], line_77[858], line_76[856], line_75[854], line_74[852], line_73[850], line_72[848], line_71[846], line_70[844], line_69[842], line_68[840], line_67[838], line_66[836], line_65[834], line_64[832], line_63[830], line_62[828], line_61[826], line_60[824], line_59[822], line_58[820], line_57[818], line_56[816], line_55[814], line_54[812], line_53[810], line_52[808], line_51[806], line_50[804], line_49[802], line_48[800], line_47[798], line_46[796], line_45[794], line_44[792], line_43[790], line_42[788], line_41[786], line_40[784], line_39[782], line_38[780], line_37[778], line_36[776], line_35[774], line_34[772], line_33[770], line_32[768], line_31[766], line_30[764], line_29[762], line_28[760], line_27[758], line_26[756], line_25[754], line_24[752], line_23[750], line_22[748], line_21[746], line_20[744], line_19[742], line_18[740], line_17[738], line_16[736], line_15[734], line_14[732], line_13[730], line_12[728], line_11[726], line_10[724], line_9[722], line_8[720], line_7[718], line_6[716], line_5[714], line_4[712], line_3[710], line_2[708], line_1[706] };
assign col_961 = {line_128[961], line_127[959], line_126[957], line_125[955], line_124[953], line_123[951], line_122[949], line_121[947], line_120[945], line_119[943], line_118[941], line_117[939], line_116[937], line_115[935], line_114[933], line_113[931], line_112[929], line_111[927], line_110[925], line_109[923], line_108[921], line_107[919], line_106[917], line_105[915], line_104[913], line_103[911], line_102[909], line_101[907], line_100[905], line_99[903], line_98[901], line_97[899], line_96[897], line_95[895], line_94[893], line_93[891], line_92[889], line_91[887], line_90[885], line_89[883], line_88[881], line_87[879], line_86[877], line_85[875], line_84[873], line_83[871], line_82[869], line_81[867], line_80[865], line_79[863], line_78[861], line_77[859], line_76[857], line_75[855], line_74[853], line_73[851], line_72[849], line_71[847], line_70[845], line_69[843], line_68[841], line_67[839], line_66[837], line_65[835], line_64[833], line_63[831], line_62[829], line_61[827], line_60[825], line_59[823], line_58[821], line_57[819], line_56[817], line_55[815], line_54[813], line_53[811], line_52[809], line_51[807], line_50[805], line_49[803], line_48[801], line_47[799], line_46[797], line_45[795], line_44[793], line_43[791], line_42[789], line_41[787], line_40[785], line_39[783], line_38[781], line_37[779], line_36[777], line_35[775], line_34[773], line_33[771], line_32[769], line_31[767], line_30[765], line_29[763], line_28[761], line_27[759], line_26[757], line_25[755], line_24[753], line_23[751], line_22[749], line_21[747], line_20[745], line_19[743], line_18[741], line_17[739], line_16[737], line_15[735], line_14[733], line_13[731], line_12[729], line_11[727], line_10[725], line_9[723], line_8[721], line_7[719], line_6[717], line_5[715], line_4[713], line_3[711], line_2[709], line_1[707] };
assign col_962 = {line_128[962], line_127[960], line_126[958], line_125[956], line_124[954], line_123[952], line_122[950], line_121[948], line_120[946], line_119[944], line_118[942], line_117[940], line_116[938], line_115[936], line_114[934], line_113[932], line_112[930], line_111[928], line_110[926], line_109[924], line_108[922], line_107[920], line_106[918], line_105[916], line_104[914], line_103[912], line_102[910], line_101[908], line_100[906], line_99[904], line_98[902], line_97[900], line_96[898], line_95[896], line_94[894], line_93[892], line_92[890], line_91[888], line_90[886], line_89[884], line_88[882], line_87[880], line_86[878], line_85[876], line_84[874], line_83[872], line_82[870], line_81[868], line_80[866], line_79[864], line_78[862], line_77[860], line_76[858], line_75[856], line_74[854], line_73[852], line_72[850], line_71[848], line_70[846], line_69[844], line_68[842], line_67[840], line_66[838], line_65[836], line_64[834], line_63[832], line_62[830], line_61[828], line_60[826], line_59[824], line_58[822], line_57[820], line_56[818], line_55[816], line_54[814], line_53[812], line_52[810], line_51[808], line_50[806], line_49[804], line_48[802], line_47[800], line_46[798], line_45[796], line_44[794], line_43[792], line_42[790], line_41[788], line_40[786], line_39[784], line_38[782], line_37[780], line_36[778], line_35[776], line_34[774], line_33[772], line_32[770], line_31[768], line_30[766], line_29[764], line_28[762], line_27[760], line_26[758], line_25[756], line_24[754], line_23[752], line_22[750], line_21[748], line_20[746], line_19[744], line_18[742], line_17[740], line_16[738], line_15[736], line_14[734], line_13[732], line_12[730], line_11[728], line_10[726], line_9[724], line_8[722], line_7[720], line_6[718], line_5[716], line_4[714], line_3[712], line_2[710], line_1[708] };
assign col_963 = {line_128[963], line_127[961], line_126[959], line_125[957], line_124[955], line_123[953], line_122[951], line_121[949], line_120[947], line_119[945], line_118[943], line_117[941], line_116[939], line_115[937], line_114[935], line_113[933], line_112[931], line_111[929], line_110[927], line_109[925], line_108[923], line_107[921], line_106[919], line_105[917], line_104[915], line_103[913], line_102[911], line_101[909], line_100[907], line_99[905], line_98[903], line_97[901], line_96[899], line_95[897], line_94[895], line_93[893], line_92[891], line_91[889], line_90[887], line_89[885], line_88[883], line_87[881], line_86[879], line_85[877], line_84[875], line_83[873], line_82[871], line_81[869], line_80[867], line_79[865], line_78[863], line_77[861], line_76[859], line_75[857], line_74[855], line_73[853], line_72[851], line_71[849], line_70[847], line_69[845], line_68[843], line_67[841], line_66[839], line_65[837], line_64[835], line_63[833], line_62[831], line_61[829], line_60[827], line_59[825], line_58[823], line_57[821], line_56[819], line_55[817], line_54[815], line_53[813], line_52[811], line_51[809], line_50[807], line_49[805], line_48[803], line_47[801], line_46[799], line_45[797], line_44[795], line_43[793], line_42[791], line_41[789], line_40[787], line_39[785], line_38[783], line_37[781], line_36[779], line_35[777], line_34[775], line_33[773], line_32[771], line_31[769], line_30[767], line_29[765], line_28[763], line_27[761], line_26[759], line_25[757], line_24[755], line_23[753], line_22[751], line_21[749], line_20[747], line_19[745], line_18[743], line_17[741], line_16[739], line_15[737], line_14[735], line_13[733], line_12[731], line_11[729], line_10[727], line_9[725], line_8[723], line_7[721], line_6[719], line_5[717], line_4[715], line_3[713], line_2[711], line_1[709] };
assign col_964 = {line_128[964], line_127[962], line_126[960], line_125[958], line_124[956], line_123[954], line_122[952], line_121[950], line_120[948], line_119[946], line_118[944], line_117[942], line_116[940], line_115[938], line_114[936], line_113[934], line_112[932], line_111[930], line_110[928], line_109[926], line_108[924], line_107[922], line_106[920], line_105[918], line_104[916], line_103[914], line_102[912], line_101[910], line_100[908], line_99[906], line_98[904], line_97[902], line_96[900], line_95[898], line_94[896], line_93[894], line_92[892], line_91[890], line_90[888], line_89[886], line_88[884], line_87[882], line_86[880], line_85[878], line_84[876], line_83[874], line_82[872], line_81[870], line_80[868], line_79[866], line_78[864], line_77[862], line_76[860], line_75[858], line_74[856], line_73[854], line_72[852], line_71[850], line_70[848], line_69[846], line_68[844], line_67[842], line_66[840], line_65[838], line_64[836], line_63[834], line_62[832], line_61[830], line_60[828], line_59[826], line_58[824], line_57[822], line_56[820], line_55[818], line_54[816], line_53[814], line_52[812], line_51[810], line_50[808], line_49[806], line_48[804], line_47[802], line_46[800], line_45[798], line_44[796], line_43[794], line_42[792], line_41[790], line_40[788], line_39[786], line_38[784], line_37[782], line_36[780], line_35[778], line_34[776], line_33[774], line_32[772], line_31[770], line_30[768], line_29[766], line_28[764], line_27[762], line_26[760], line_25[758], line_24[756], line_23[754], line_22[752], line_21[750], line_20[748], line_19[746], line_18[744], line_17[742], line_16[740], line_15[738], line_14[736], line_13[734], line_12[732], line_11[730], line_10[728], line_9[726], line_8[724], line_7[722], line_6[720], line_5[718], line_4[716], line_3[714], line_2[712], line_1[710] };
assign col_965 = {line_128[965], line_127[963], line_126[961], line_125[959], line_124[957], line_123[955], line_122[953], line_121[951], line_120[949], line_119[947], line_118[945], line_117[943], line_116[941], line_115[939], line_114[937], line_113[935], line_112[933], line_111[931], line_110[929], line_109[927], line_108[925], line_107[923], line_106[921], line_105[919], line_104[917], line_103[915], line_102[913], line_101[911], line_100[909], line_99[907], line_98[905], line_97[903], line_96[901], line_95[899], line_94[897], line_93[895], line_92[893], line_91[891], line_90[889], line_89[887], line_88[885], line_87[883], line_86[881], line_85[879], line_84[877], line_83[875], line_82[873], line_81[871], line_80[869], line_79[867], line_78[865], line_77[863], line_76[861], line_75[859], line_74[857], line_73[855], line_72[853], line_71[851], line_70[849], line_69[847], line_68[845], line_67[843], line_66[841], line_65[839], line_64[837], line_63[835], line_62[833], line_61[831], line_60[829], line_59[827], line_58[825], line_57[823], line_56[821], line_55[819], line_54[817], line_53[815], line_52[813], line_51[811], line_50[809], line_49[807], line_48[805], line_47[803], line_46[801], line_45[799], line_44[797], line_43[795], line_42[793], line_41[791], line_40[789], line_39[787], line_38[785], line_37[783], line_36[781], line_35[779], line_34[777], line_33[775], line_32[773], line_31[771], line_30[769], line_29[767], line_28[765], line_27[763], line_26[761], line_25[759], line_24[757], line_23[755], line_22[753], line_21[751], line_20[749], line_19[747], line_18[745], line_17[743], line_16[741], line_15[739], line_14[737], line_13[735], line_12[733], line_11[731], line_10[729], line_9[727], line_8[725], line_7[723], line_6[721], line_5[719], line_4[717], line_3[715], line_2[713], line_1[711] };
assign col_966 = {line_128[966], line_127[964], line_126[962], line_125[960], line_124[958], line_123[956], line_122[954], line_121[952], line_120[950], line_119[948], line_118[946], line_117[944], line_116[942], line_115[940], line_114[938], line_113[936], line_112[934], line_111[932], line_110[930], line_109[928], line_108[926], line_107[924], line_106[922], line_105[920], line_104[918], line_103[916], line_102[914], line_101[912], line_100[910], line_99[908], line_98[906], line_97[904], line_96[902], line_95[900], line_94[898], line_93[896], line_92[894], line_91[892], line_90[890], line_89[888], line_88[886], line_87[884], line_86[882], line_85[880], line_84[878], line_83[876], line_82[874], line_81[872], line_80[870], line_79[868], line_78[866], line_77[864], line_76[862], line_75[860], line_74[858], line_73[856], line_72[854], line_71[852], line_70[850], line_69[848], line_68[846], line_67[844], line_66[842], line_65[840], line_64[838], line_63[836], line_62[834], line_61[832], line_60[830], line_59[828], line_58[826], line_57[824], line_56[822], line_55[820], line_54[818], line_53[816], line_52[814], line_51[812], line_50[810], line_49[808], line_48[806], line_47[804], line_46[802], line_45[800], line_44[798], line_43[796], line_42[794], line_41[792], line_40[790], line_39[788], line_38[786], line_37[784], line_36[782], line_35[780], line_34[778], line_33[776], line_32[774], line_31[772], line_30[770], line_29[768], line_28[766], line_27[764], line_26[762], line_25[760], line_24[758], line_23[756], line_22[754], line_21[752], line_20[750], line_19[748], line_18[746], line_17[744], line_16[742], line_15[740], line_14[738], line_13[736], line_12[734], line_11[732], line_10[730], line_9[728], line_8[726], line_7[724], line_6[722], line_5[720], line_4[718], line_3[716], line_2[714], line_1[712] };
assign col_967 = {line_128[967], line_127[965], line_126[963], line_125[961], line_124[959], line_123[957], line_122[955], line_121[953], line_120[951], line_119[949], line_118[947], line_117[945], line_116[943], line_115[941], line_114[939], line_113[937], line_112[935], line_111[933], line_110[931], line_109[929], line_108[927], line_107[925], line_106[923], line_105[921], line_104[919], line_103[917], line_102[915], line_101[913], line_100[911], line_99[909], line_98[907], line_97[905], line_96[903], line_95[901], line_94[899], line_93[897], line_92[895], line_91[893], line_90[891], line_89[889], line_88[887], line_87[885], line_86[883], line_85[881], line_84[879], line_83[877], line_82[875], line_81[873], line_80[871], line_79[869], line_78[867], line_77[865], line_76[863], line_75[861], line_74[859], line_73[857], line_72[855], line_71[853], line_70[851], line_69[849], line_68[847], line_67[845], line_66[843], line_65[841], line_64[839], line_63[837], line_62[835], line_61[833], line_60[831], line_59[829], line_58[827], line_57[825], line_56[823], line_55[821], line_54[819], line_53[817], line_52[815], line_51[813], line_50[811], line_49[809], line_48[807], line_47[805], line_46[803], line_45[801], line_44[799], line_43[797], line_42[795], line_41[793], line_40[791], line_39[789], line_38[787], line_37[785], line_36[783], line_35[781], line_34[779], line_33[777], line_32[775], line_31[773], line_30[771], line_29[769], line_28[767], line_27[765], line_26[763], line_25[761], line_24[759], line_23[757], line_22[755], line_21[753], line_20[751], line_19[749], line_18[747], line_17[745], line_16[743], line_15[741], line_14[739], line_13[737], line_12[735], line_11[733], line_10[731], line_9[729], line_8[727], line_7[725], line_6[723], line_5[721], line_4[719], line_3[717], line_2[715], line_1[713] };
assign col_968 = {line_128[968], line_127[966], line_126[964], line_125[962], line_124[960], line_123[958], line_122[956], line_121[954], line_120[952], line_119[950], line_118[948], line_117[946], line_116[944], line_115[942], line_114[940], line_113[938], line_112[936], line_111[934], line_110[932], line_109[930], line_108[928], line_107[926], line_106[924], line_105[922], line_104[920], line_103[918], line_102[916], line_101[914], line_100[912], line_99[910], line_98[908], line_97[906], line_96[904], line_95[902], line_94[900], line_93[898], line_92[896], line_91[894], line_90[892], line_89[890], line_88[888], line_87[886], line_86[884], line_85[882], line_84[880], line_83[878], line_82[876], line_81[874], line_80[872], line_79[870], line_78[868], line_77[866], line_76[864], line_75[862], line_74[860], line_73[858], line_72[856], line_71[854], line_70[852], line_69[850], line_68[848], line_67[846], line_66[844], line_65[842], line_64[840], line_63[838], line_62[836], line_61[834], line_60[832], line_59[830], line_58[828], line_57[826], line_56[824], line_55[822], line_54[820], line_53[818], line_52[816], line_51[814], line_50[812], line_49[810], line_48[808], line_47[806], line_46[804], line_45[802], line_44[800], line_43[798], line_42[796], line_41[794], line_40[792], line_39[790], line_38[788], line_37[786], line_36[784], line_35[782], line_34[780], line_33[778], line_32[776], line_31[774], line_30[772], line_29[770], line_28[768], line_27[766], line_26[764], line_25[762], line_24[760], line_23[758], line_22[756], line_21[754], line_20[752], line_19[750], line_18[748], line_17[746], line_16[744], line_15[742], line_14[740], line_13[738], line_12[736], line_11[734], line_10[732], line_9[730], line_8[728], line_7[726], line_6[724], line_5[722], line_4[720], line_3[718], line_2[716], line_1[714] };
assign col_969 = {line_128[969], line_127[967], line_126[965], line_125[963], line_124[961], line_123[959], line_122[957], line_121[955], line_120[953], line_119[951], line_118[949], line_117[947], line_116[945], line_115[943], line_114[941], line_113[939], line_112[937], line_111[935], line_110[933], line_109[931], line_108[929], line_107[927], line_106[925], line_105[923], line_104[921], line_103[919], line_102[917], line_101[915], line_100[913], line_99[911], line_98[909], line_97[907], line_96[905], line_95[903], line_94[901], line_93[899], line_92[897], line_91[895], line_90[893], line_89[891], line_88[889], line_87[887], line_86[885], line_85[883], line_84[881], line_83[879], line_82[877], line_81[875], line_80[873], line_79[871], line_78[869], line_77[867], line_76[865], line_75[863], line_74[861], line_73[859], line_72[857], line_71[855], line_70[853], line_69[851], line_68[849], line_67[847], line_66[845], line_65[843], line_64[841], line_63[839], line_62[837], line_61[835], line_60[833], line_59[831], line_58[829], line_57[827], line_56[825], line_55[823], line_54[821], line_53[819], line_52[817], line_51[815], line_50[813], line_49[811], line_48[809], line_47[807], line_46[805], line_45[803], line_44[801], line_43[799], line_42[797], line_41[795], line_40[793], line_39[791], line_38[789], line_37[787], line_36[785], line_35[783], line_34[781], line_33[779], line_32[777], line_31[775], line_30[773], line_29[771], line_28[769], line_27[767], line_26[765], line_25[763], line_24[761], line_23[759], line_22[757], line_21[755], line_20[753], line_19[751], line_18[749], line_17[747], line_16[745], line_15[743], line_14[741], line_13[739], line_12[737], line_11[735], line_10[733], line_9[731], line_8[729], line_7[727], line_6[725], line_5[723], line_4[721], line_3[719], line_2[717], line_1[715] };
assign col_970 = {line_128[970], line_127[968], line_126[966], line_125[964], line_124[962], line_123[960], line_122[958], line_121[956], line_120[954], line_119[952], line_118[950], line_117[948], line_116[946], line_115[944], line_114[942], line_113[940], line_112[938], line_111[936], line_110[934], line_109[932], line_108[930], line_107[928], line_106[926], line_105[924], line_104[922], line_103[920], line_102[918], line_101[916], line_100[914], line_99[912], line_98[910], line_97[908], line_96[906], line_95[904], line_94[902], line_93[900], line_92[898], line_91[896], line_90[894], line_89[892], line_88[890], line_87[888], line_86[886], line_85[884], line_84[882], line_83[880], line_82[878], line_81[876], line_80[874], line_79[872], line_78[870], line_77[868], line_76[866], line_75[864], line_74[862], line_73[860], line_72[858], line_71[856], line_70[854], line_69[852], line_68[850], line_67[848], line_66[846], line_65[844], line_64[842], line_63[840], line_62[838], line_61[836], line_60[834], line_59[832], line_58[830], line_57[828], line_56[826], line_55[824], line_54[822], line_53[820], line_52[818], line_51[816], line_50[814], line_49[812], line_48[810], line_47[808], line_46[806], line_45[804], line_44[802], line_43[800], line_42[798], line_41[796], line_40[794], line_39[792], line_38[790], line_37[788], line_36[786], line_35[784], line_34[782], line_33[780], line_32[778], line_31[776], line_30[774], line_29[772], line_28[770], line_27[768], line_26[766], line_25[764], line_24[762], line_23[760], line_22[758], line_21[756], line_20[754], line_19[752], line_18[750], line_17[748], line_16[746], line_15[744], line_14[742], line_13[740], line_12[738], line_11[736], line_10[734], line_9[732], line_8[730], line_7[728], line_6[726], line_5[724], line_4[722], line_3[720], line_2[718], line_1[716] };
assign col_971 = {line_128[971], line_127[969], line_126[967], line_125[965], line_124[963], line_123[961], line_122[959], line_121[957], line_120[955], line_119[953], line_118[951], line_117[949], line_116[947], line_115[945], line_114[943], line_113[941], line_112[939], line_111[937], line_110[935], line_109[933], line_108[931], line_107[929], line_106[927], line_105[925], line_104[923], line_103[921], line_102[919], line_101[917], line_100[915], line_99[913], line_98[911], line_97[909], line_96[907], line_95[905], line_94[903], line_93[901], line_92[899], line_91[897], line_90[895], line_89[893], line_88[891], line_87[889], line_86[887], line_85[885], line_84[883], line_83[881], line_82[879], line_81[877], line_80[875], line_79[873], line_78[871], line_77[869], line_76[867], line_75[865], line_74[863], line_73[861], line_72[859], line_71[857], line_70[855], line_69[853], line_68[851], line_67[849], line_66[847], line_65[845], line_64[843], line_63[841], line_62[839], line_61[837], line_60[835], line_59[833], line_58[831], line_57[829], line_56[827], line_55[825], line_54[823], line_53[821], line_52[819], line_51[817], line_50[815], line_49[813], line_48[811], line_47[809], line_46[807], line_45[805], line_44[803], line_43[801], line_42[799], line_41[797], line_40[795], line_39[793], line_38[791], line_37[789], line_36[787], line_35[785], line_34[783], line_33[781], line_32[779], line_31[777], line_30[775], line_29[773], line_28[771], line_27[769], line_26[767], line_25[765], line_24[763], line_23[761], line_22[759], line_21[757], line_20[755], line_19[753], line_18[751], line_17[749], line_16[747], line_15[745], line_14[743], line_13[741], line_12[739], line_11[737], line_10[735], line_9[733], line_8[731], line_7[729], line_6[727], line_5[725], line_4[723], line_3[721], line_2[719], line_1[717] };
assign col_972 = {line_128[972], line_127[970], line_126[968], line_125[966], line_124[964], line_123[962], line_122[960], line_121[958], line_120[956], line_119[954], line_118[952], line_117[950], line_116[948], line_115[946], line_114[944], line_113[942], line_112[940], line_111[938], line_110[936], line_109[934], line_108[932], line_107[930], line_106[928], line_105[926], line_104[924], line_103[922], line_102[920], line_101[918], line_100[916], line_99[914], line_98[912], line_97[910], line_96[908], line_95[906], line_94[904], line_93[902], line_92[900], line_91[898], line_90[896], line_89[894], line_88[892], line_87[890], line_86[888], line_85[886], line_84[884], line_83[882], line_82[880], line_81[878], line_80[876], line_79[874], line_78[872], line_77[870], line_76[868], line_75[866], line_74[864], line_73[862], line_72[860], line_71[858], line_70[856], line_69[854], line_68[852], line_67[850], line_66[848], line_65[846], line_64[844], line_63[842], line_62[840], line_61[838], line_60[836], line_59[834], line_58[832], line_57[830], line_56[828], line_55[826], line_54[824], line_53[822], line_52[820], line_51[818], line_50[816], line_49[814], line_48[812], line_47[810], line_46[808], line_45[806], line_44[804], line_43[802], line_42[800], line_41[798], line_40[796], line_39[794], line_38[792], line_37[790], line_36[788], line_35[786], line_34[784], line_33[782], line_32[780], line_31[778], line_30[776], line_29[774], line_28[772], line_27[770], line_26[768], line_25[766], line_24[764], line_23[762], line_22[760], line_21[758], line_20[756], line_19[754], line_18[752], line_17[750], line_16[748], line_15[746], line_14[744], line_13[742], line_12[740], line_11[738], line_10[736], line_9[734], line_8[732], line_7[730], line_6[728], line_5[726], line_4[724], line_3[722], line_2[720], line_1[718] };
assign col_973 = {line_128[973], line_127[971], line_126[969], line_125[967], line_124[965], line_123[963], line_122[961], line_121[959], line_120[957], line_119[955], line_118[953], line_117[951], line_116[949], line_115[947], line_114[945], line_113[943], line_112[941], line_111[939], line_110[937], line_109[935], line_108[933], line_107[931], line_106[929], line_105[927], line_104[925], line_103[923], line_102[921], line_101[919], line_100[917], line_99[915], line_98[913], line_97[911], line_96[909], line_95[907], line_94[905], line_93[903], line_92[901], line_91[899], line_90[897], line_89[895], line_88[893], line_87[891], line_86[889], line_85[887], line_84[885], line_83[883], line_82[881], line_81[879], line_80[877], line_79[875], line_78[873], line_77[871], line_76[869], line_75[867], line_74[865], line_73[863], line_72[861], line_71[859], line_70[857], line_69[855], line_68[853], line_67[851], line_66[849], line_65[847], line_64[845], line_63[843], line_62[841], line_61[839], line_60[837], line_59[835], line_58[833], line_57[831], line_56[829], line_55[827], line_54[825], line_53[823], line_52[821], line_51[819], line_50[817], line_49[815], line_48[813], line_47[811], line_46[809], line_45[807], line_44[805], line_43[803], line_42[801], line_41[799], line_40[797], line_39[795], line_38[793], line_37[791], line_36[789], line_35[787], line_34[785], line_33[783], line_32[781], line_31[779], line_30[777], line_29[775], line_28[773], line_27[771], line_26[769], line_25[767], line_24[765], line_23[763], line_22[761], line_21[759], line_20[757], line_19[755], line_18[753], line_17[751], line_16[749], line_15[747], line_14[745], line_13[743], line_12[741], line_11[739], line_10[737], line_9[735], line_8[733], line_7[731], line_6[729], line_5[727], line_4[725], line_3[723], line_2[721], line_1[719] };
assign col_974 = {line_128[974], line_127[972], line_126[970], line_125[968], line_124[966], line_123[964], line_122[962], line_121[960], line_120[958], line_119[956], line_118[954], line_117[952], line_116[950], line_115[948], line_114[946], line_113[944], line_112[942], line_111[940], line_110[938], line_109[936], line_108[934], line_107[932], line_106[930], line_105[928], line_104[926], line_103[924], line_102[922], line_101[920], line_100[918], line_99[916], line_98[914], line_97[912], line_96[910], line_95[908], line_94[906], line_93[904], line_92[902], line_91[900], line_90[898], line_89[896], line_88[894], line_87[892], line_86[890], line_85[888], line_84[886], line_83[884], line_82[882], line_81[880], line_80[878], line_79[876], line_78[874], line_77[872], line_76[870], line_75[868], line_74[866], line_73[864], line_72[862], line_71[860], line_70[858], line_69[856], line_68[854], line_67[852], line_66[850], line_65[848], line_64[846], line_63[844], line_62[842], line_61[840], line_60[838], line_59[836], line_58[834], line_57[832], line_56[830], line_55[828], line_54[826], line_53[824], line_52[822], line_51[820], line_50[818], line_49[816], line_48[814], line_47[812], line_46[810], line_45[808], line_44[806], line_43[804], line_42[802], line_41[800], line_40[798], line_39[796], line_38[794], line_37[792], line_36[790], line_35[788], line_34[786], line_33[784], line_32[782], line_31[780], line_30[778], line_29[776], line_28[774], line_27[772], line_26[770], line_25[768], line_24[766], line_23[764], line_22[762], line_21[760], line_20[758], line_19[756], line_18[754], line_17[752], line_16[750], line_15[748], line_14[746], line_13[744], line_12[742], line_11[740], line_10[738], line_9[736], line_8[734], line_7[732], line_6[730], line_5[728], line_4[726], line_3[724], line_2[722], line_1[720] };
assign col_975 = {line_128[975], line_127[973], line_126[971], line_125[969], line_124[967], line_123[965], line_122[963], line_121[961], line_120[959], line_119[957], line_118[955], line_117[953], line_116[951], line_115[949], line_114[947], line_113[945], line_112[943], line_111[941], line_110[939], line_109[937], line_108[935], line_107[933], line_106[931], line_105[929], line_104[927], line_103[925], line_102[923], line_101[921], line_100[919], line_99[917], line_98[915], line_97[913], line_96[911], line_95[909], line_94[907], line_93[905], line_92[903], line_91[901], line_90[899], line_89[897], line_88[895], line_87[893], line_86[891], line_85[889], line_84[887], line_83[885], line_82[883], line_81[881], line_80[879], line_79[877], line_78[875], line_77[873], line_76[871], line_75[869], line_74[867], line_73[865], line_72[863], line_71[861], line_70[859], line_69[857], line_68[855], line_67[853], line_66[851], line_65[849], line_64[847], line_63[845], line_62[843], line_61[841], line_60[839], line_59[837], line_58[835], line_57[833], line_56[831], line_55[829], line_54[827], line_53[825], line_52[823], line_51[821], line_50[819], line_49[817], line_48[815], line_47[813], line_46[811], line_45[809], line_44[807], line_43[805], line_42[803], line_41[801], line_40[799], line_39[797], line_38[795], line_37[793], line_36[791], line_35[789], line_34[787], line_33[785], line_32[783], line_31[781], line_30[779], line_29[777], line_28[775], line_27[773], line_26[771], line_25[769], line_24[767], line_23[765], line_22[763], line_21[761], line_20[759], line_19[757], line_18[755], line_17[753], line_16[751], line_15[749], line_14[747], line_13[745], line_12[743], line_11[741], line_10[739], line_9[737], line_8[735], line_7[733], line_6[731], line_5[729], line_4[727], line_3[725], line_2[723], line_1[721] };
assign col_976 = {line_128[976], line_127[974], line_126[972], line_125[970], line_124[968], line_123[966], line_122[964], line_121[962], line_120[960], line_119[958], line_118[956], line_117[954], line_116[952], line_115[950], line_114[948], line_113[946], line_112[944], line_111[942], line_110[940], line_109[938], line_108[936], line_107[934], line_106[932], line_105[930], line_104[928], line_103[926], line_102[924], line_101[922], line_100[920], line_99[918], line_98[916], line_97[914], line_96[912], line_95[910], line_94[908], line_93[906], line_92[904], line_91[902], line_90[900], line_89[898], line_88[896], line_87[894], line_86[892], line_85[890], line_84[888], line_83[886], line_82[884], line_81[882], line_80[880], line_79[878], line_78[876], line_77[874], line_76[872], line_75[870], line_74[868], line_73[866], line_72[864], line_71[862], line_70[860], line_69[858], line_68[856], line_67[854], line_66[852], line_65[850], line_64[848], line_63[846], line_62[844], line_61[842], line_60[840], line_59[838], line_58[836], line_57[834], line_56[832], line_55[830], line_54[828], line_53[826], line_52[824], line_51[822], line_50[820], line_49[818], line_48[816], line_47[814], line_46[812], line_45[810], line_44[808], line_43[806], line_42[804], line_41[802], line_40[800], line_39[798], line_38[796], line_37[794], line_36[792], line_35[790], line_34[788], line_33[786], line_32[784], line_31[782], line_30[780], line_29[778], line_28[776], line_27[774], line_26[772], line_25[770], line_24[768], line_23[766], line_22[764], line_21[762], line_20[760], line_19[758], line_18[756], line_17[754], line_16[752], line_15[750], line_14[748], line_13[746], line_12[744], line_11[742], line_10[740], line_9[738], line_8[736], line_7[734], line_6[732], line_5[730], line_4[728], line_3[726], line_2[724], line_1[722] };
assign col_977 = {line_128[977], line_127[975], line_126[973], line_125[971], line_124[969], line_123[967], line_122[965], line_121[963], line_120[961], line_119[959], line_118[957], line_117[955], line_116[953], line_115[951], line_114[949], line_113[947], line_112[945], line_111[943], line_110[941], line_109[939], line_108[937], line_107[935], line_106[933], line_105[931], line_104[929], line_103[927], line_102[925], line_101[923], line_100[921], line_99[919], line_98[917], line_97[915], line_96[913], line_95[911], line_94[909], line_93[907], line_92[905], line_91[903], line_90[901], line_89[899], line_88[897], line_87[895], line_86[893], line_85[891], line_84[889], line_83[887], line_82[885], line_81[883], line_80[881], line_79[879], line_78[877], line_77[875], line_76[873], line_75[871], line_74[869], line_73[867], line_72[865], line_71[863], line_70[861], line_69[859], line_68[857], line_67[855], line_66[853], line_65[851], line_64[849], line_63[847], line_62[845], line_61[843], line_60[841], line_59[839], line_58[837], line_57[835], line_56[833], line_55[831], line_54[829], line_53[827], line_52[825], line_51[823], line_50[821], line_49[819], line_48[817], line_47[815], line_46[813], line_45[811], line_44[809], line_43[807], line_42[805], line_41[803], line_40[801], line_39[799], line_38[797], line_37[795], line_36[793], line_35[791], line_34[789], line_33[787], line_32[785], line_31[783], line_30[781], line_29[779], line_28[777], line_27[775], line_26[773], line_25[771], line_24[769], line_23[767], line_22[765], line_21[763], line_20[761], line_19[759], line_18[757], line_17[755], line_16[753], line_15[751], line_14[749], line_13[747], line_12[745], line_11[743], line_10[741], line_9[739], line_8[737], line_7[735], line_6[733], line_5[731], line_4[729], line_3[727], line_2[725], line_1[723] };
assign col_978 = {line_128[978], line_127[976], line_126[974], line_125[972], line_124[970], line_123[968], line_122[966], line_121[964], line_120[962], line_119[960], line_118[958], line_117[956], line_116[954], line_115[952], line_114[950], line_113[948], line_112[946], line_111[944], line_110[942], line_109[940], line_108[938], line_107[936], line_106[934], line_105[932], line_104[930], line_103[928], line_102[926], line_101[924], line_100[922], line_99[920], line_98[918], line_97[916], line_96[914], line_95[912], line_94[910], line_93[908], line_92[906], line_91[904], line_90[902], line_89[900], line_88[898], line_87[896], line_86[894], line_85[892], line_84[890], line_83[888], line_82[886], line_81[884], line_80[882], line_79[880], line_78[878], line_77[876], line_76[874], line_75[872], line_74[870], line_73[868], line_72[866], line_71[864], line_70[862], line_69[860], line_68[858], line_67[856], line_66[854], line_65[852], line_64[850], line_63[848], line_62[846], line_61[844], line_60[842], line_59[840], line_58[838], line_57[836], line_56[834], line_55[832], line_54[830], line_53[828], line_52[826], line_51[824], line_50[822], line_49[820], line_48[818], line_47[816], line_46[814], line_45[812], line_44[810], line_43[808], line_42[806], line_41[804], line_40[802], line_39[800], line_38[798], line_37[796], line_36[794], line_35[792], line_34[790], line_33[788], line_32[786], line_31[784], line_30[782], line_29[780], line_28[778], line_27[776], line_26[774], line_25[772], line_24[770], line_23[768], line_22[766], line_21[764], line_20[762], line_19[760], line_18[758], line_17[756], line_16[754], line_15[752], line_14[750], line_13[748], line_12[746], line_11[744], line_10[742], line_9[740], line_8[738], line_7[736], line_6[734], line_5[732], line_4[730], line_3[728], line_2[726], line_1[724] };
assign col_979 = {line_128[979], line_127[977], line_126[975], line_125[973], line_124[971], line_123[969], line_122[967], line_121[965], line_120[963], line_119[961], line_118[959], line_117[957], line_116[955], line_115[953], line_114[951], line_113[949], line_112[947], line_111[945], line_110[943], line_109[941], line_108[939], line_107[937], line_106[935], line_105[933], line_104[931], line_103[929], line_102[927], line_101[925], line_100[923], line_99[921], line_98[919], line_97[917], line_96[915], line_95[913], line_94[911], line_93[909], line_92[907], line_91[905], line_90[903], line_89[901], line_88[899], line_87[897], line_86[895], line_85[893], line_84[891], line_83[889], line_82[887], line_81[885], line_80[883], line_79[881], line_78[879], line_77[877], line_76[875], line_75[873], line_74[871], line_73[869], line_72[867], line_71[865], line_70[863], line_69[861], line_68[859], line_67[857], line_66[855], line_65[853], line_64[851], line_63[849], line_62[847], line_61[845], line_60[843], line_59[841], line_58[839], line_57[837], line_56[835], line_55[833], line_54[831], line_53[829], line_52[827], line_51[825], line_50[823], line_49[821], line_48[819], line_47[817], line_46[815], line_45[813], line_44[811], line_43[809], line_42[807], line_41[805], line_40[803], line_39[801], line_38[799], line_37[797], line_36[795], line_35[793], line_34[791], line_33[789], line_32[787], line_31[785], line_30[783], line_29[781], line_28[779], line_27[777], line_26[775], line_25[773], line_24[771], line_23[769], line_22[767], line_21[765], line_20[763], line_19[761], line_18[759], line_17[757], line_16[755], line_15[753], line_14[751], line_13[749], line_12[747], line_11[745], line_10[743], line_9[741], line_8[739], line_7[737], line_6[735], line_5[733], line_4[731], line_3[729], line_2[727], line_1[725] };
assign col_980 = {line_128[980], line_127[978], line_126[976], line_125[974], line_124[972], line_123[970], line_122[968], line_121[966], line_120[964], line_119[962], line_118[960], line_117[958], line_116[956], line_115[954], line_114[952], line_113[950], line_112[948], line_111[946], line_110[944], line_109[942], line_108[940], line_107[938], line_106[936], line_105[934], line_104[932], line_103[930], line_102[928], line_101[926], line_100[924], line_99[922], line_98[920], line_97[918], line_96[916], line_95[914], line_94[912], line_93[910], line_92[908], line_91[906], line_90[904], line_89[902], line_88[900], line_87[898], line_86[896], line_85[894], line_84[892], line_83[890], line_82[888], line_81[886], line_80[884], line_79[882], line_78[880], line_77[878], line_76[876], line_75[874], line_74[872], line_73[870], line_72[868], line_71[866], line_70[864], line_69[862], line_68[860], line_67[858], line_66[856], line_65[854], line_64[852], line_63[850], line_62[848], line_61[846], line_60[844], line_59[842], line_58[840], line_57[838], line_56[836], line_55[834], line_54[832], line_53[830], line_52[828], line_51[826], line_50[824], line_49[822], line_48[820], line_47[818], line_46[816], line_45[814], line_44[812], line_43[810], line_42[808], line_41[806], line_40[804], line_39[802], line_38[800], line_37[798], line_36[796], line_35[794], line_34[792], line_33[790], line_32[788], line_31[786], line_30[784], line_29[782], line_28[780], line_27[778], line_26[776], line_25[774], line_24[772], line_23[770], line_22[768], line_21[766], line_20[764], line_19[762], line_18[760], line_17[758], line_16[756], line_15[754], line_14[752], line_13[750], line_12[748], line_11[746], line_10[744], line_9[742], line_8[740], line_7[738], line_6[736], line_5[734], line_4[732], line_3[730], line_2[728], line_1[726] };
assign col_981 = {line_128[981], line_127[979], line_126[977], line_125[975], line_124[973], line_123[971], line_122[969], line_121[967], line_120[965], line_119[963], line_118[961], line_117[959], line_116[957], line_115[955], line_114[953], line_113[951], line_112[949], line_111[947], line_110[945], line_109[943], line_108[941], line_107[939], line_106[937], line_105[935], line_104[933], line_103[931], line_102[929], line_101[927], line_100[925], line_99[923], line_98[921], line_97[919], line_96[917], line_95[915], line_94[913], line_93[911], line_92[909], line_91[907], line_90[905], line_89[903], line_88[901], line_87[899], line_86[897], line_85[895], line_84[893], line_83[891], line_82[889], line_81[887], line_80[885], line_79[883], line_78[881], line_77[879], line_76[877], line_75[875], line_74[873], line_73[871], line_72[869], line_71[867], line_70[865], line_69[863], line_68[861], line_67[859], line_66[857], line_65[855], line_64[853], line_63[851], line_62[849], line_61[847], line_60[845], line_59[843], line_58[841], line_57[839], line_56[837], line_55[835], line_54[833], line_53[831], line_52[829], line_51[827], line_50[825], line_49[823], line_48[821], line_47[819], line_46[817], line_45[815], line_44[813], line_43[811], line_42[809], line_41[807], line_40[805], line_39[803], line_38[801], line_37[799], line_36[797], line_35[795], line_34[793], line_33[791], line_32[789], line_31[787], line_30[785], line_29[783], line_28[781], line_27[779], line_26[777], line_25[775], line_24[773], line_23[771], line_22[769], line_21[767], line_20[765], line_19[763], line_18[761], line_17[759], line_16[757], line_15[755], line_14[753], line_13[751], line_12[749], line_11[747], line_10[745], line_9[743], line_8[741], line_7[739], line_6[737], line_5[735], line_4[733], line_3[731], line_2[729], line_1[727] };
assign col_982 = {line_128[982], line_127[980], line_126[978], line_125[976], line_124[974], line_123[972], line_122[970], line_121[968], line_120[966], line_119[964], line_118[962], line_117[960], line_116[958], line_115[956], line_114[954], line_113[952], line_112[950], line_111[948], line_110[946], line_109[944], line_108[942], line_107[940], line_106[938], line_105[936], line_104[934], line_103[932], line_102[930], line_101[928], line_100[926], line_99[924], line_98[922], line_97[920], line_96[918], line_95[916], line_94[914], line_93[912], line_92[910], line_91[908], line_90[906], line_89[904], line_88[902], line_87[900], line_86[898], line_85[896], line_84[894], line_83[892], line_82[890], line_81[888], line_80[886], line_79[884], line_78[882], line_77[880], line_76[878], line_75[876], line_74[874], line_73[872], line_72[870], line_71[868], line_70[866], line_69[864], line_68[862], line_67[860], line_66[858], line_65[856], line_64[854], line_63[852], line_62[850], line_61[848], line_60[846], line_59[844], line_58[842], line_57[840], line_56[838], line_55[836], line_54[834], line_53[832], line_52[830], line_51[828], line_50[826], line_49[824], line_48[822], line_47[820], line_46[818], line_45[816], line_44[814], line_43[812], line_42[810], line_41[808], line_40[806], line_39[804], line_38[802], line_37[800], line_36[798], line_35[796], line_34[794], line_33[792], line_32[790], line_31[788], line_30[786], line_29[784], line_28[782], line_27[780], line_26[778], line_25[776], line_24[774], line_23[772], line_22[770], line_21[768], line_20[766], line_19[764], line_18[762], line_17[760], line_16[758], line_15[756], line_14[754], line_13[752], line_12[750], line_11[748], line_10[746], line_9[744], line_8[742], line_7[740], line_6[738], line_5[736], line_4[734], line_3[732], line_2[730], line_1[728] };
assign col_983 = {line_128[983], line_127[981], line_126[979], line_125[977], line_124[975], line_123[973], line_122[971], line_121[969], line_120[967], line_119[965], line_118[963], line_117[961], line_116[959], line_115[957], line_114[955], line_113[953], line_112[951], line_111[949], line_110[947], line_109[945], line_108[943], line_107[941], line_106[939], line_105[937], line_104[935], line_103[933], line_102[931], line_101[929], line_100[927], line_99[925], line_98[923], line_97[921], line_96[919], line_95[917], line_94[915], line_93[913], line_92[911], line_91[909], line_90[907], line_89[905], line_88[903], line_87[901], line_86[899], line_85[897], line_84[895], line_83[893], line_82[891], line_81[889], line_80[887], line_79[885], line_78[883], line_77[881], line_76[879], line_75[877], line_74[875], line_73[873], line_72[871], line_71[869], line_70[867], line_69[865], line_68[863], line_67[861], line_66[859], line_65[857], line_64[855], line_63[853], line_62[851], line_61[849], line_60[847], line_59[845], line_58[843], line_57[841], line_56[839], line_55[837], line_54[835], line_53[833], line_52[831], line_51[829], line_50[827], line_49[825], line_48[823], line_47[821], line_46[819], line_45[817], line_44[815], line_43[813], line_42[811], line_41[809], line_40[807], line_39[805], line_38[803], line_37[801], line_36[799], line_35[797], line_34[795], line_33[793], line_32[791], line_31[789], line_30[787], line_29[785], line_28[783], line_27[781], line_26[779], line_25[777], line_24[775], line_23[773], line_22[771], line_21[769], line_20[767], line_19[765], line_18[763], line_17[761], line_16[759], line_15[757], line_14[755], line_13[753], line_12[751], line_11[749], line_10[747], line_9[745], line_8[743], line_7[741], line_6[739], line_5[737], line_4[735], line_3[733], line_2[731], line_1[729] };
assign col_984 = {line_128[984], line_127[982], line_126[980], line_125[978], line_124[976], line_123[974], line_122[972], line_121[970], line_120[968], line_119[966], line_118[964], line_117[962], line_116[960], line_115[958], line_114[956], line_113[954], line_112[952], line_111[950], line_110[948], line_109[946], line_108[944], line_107[942], line_106[940], line_105[938], line_104[936], line_103[934], line_102[932], line_101[930], line_100[928], line_99[926], line_98[924], line_97[922], line_96[920], line_95[918], line_94[916], line_93[914], line_92[912], line_91[910], line_90[908], line_89[906], line_88[904], line_87[902], line_86[900], line_85[898], line_84[896], line_83[894], line_82[892], line_81[890], line_80[888], line_79[886], line_78[884], line_77[882], line_76[880], line_75[878], line_74[876], line_73[874], line_72[872], line_71[870], line_70[868], line_69[866], line_68[864], line_67[862], line_66[860], line_65[858], line_64[856], line_63[854], line_62[852], line_61[850], line_60[848], line_59[846], line_58[844], line_57[842], line_56[840], line_55[838], line_54[836], line_53[834], line_52[832], line_51[830], line_50[828], line_49[826], line_48[824], line_47[822], line_46[820], line_45[818], line_44[816], line_43[814], line_42[812], line_41[810], line_40[808], line_39[806], line_38[804], line_37[802], line_36[800], line_35[798], line_34[796], line_33[794], line_32[792], line_31[790], line_30[788], line_29[786], line_28[784], line_27[782], line_26[780], line_25[778], line_24[776], line_23[774], line_22[772], line_21[770], line_20[768], line_19[766], line_18[764], line_17[762], line_16[760], line_15[758], line_14[756], line_13[754], line_12[752], line_11[750], line_10[748], line_9[746], line_8[744], line_7[742], line_6[740], line_5[738], line_4[736], line_3[734], line_2[732], line_1[730] };
assign col_985 = {line_128[985], line_127[983], line_126[981], line_125[979], line_124[977], line_123[975], line_122[973], line_121[971], line_120[969], line_119[967], line_118[965], line_117[963], line_116[961], line_115[959], line_114[957], line_113[955], line_112[953], line_111[951], line_110[949], line_109[947], line_108[945], line_107[943], line_106[941], line_105[939], line_104[937], line_103[935], line_102[933], line_101[931], line_100[929], line_99[927], line_98[925], line_97[923], line_96[921], line_95[919], line_94[917], line_93[915], line_92[913], line_91[911], line_90[909], line_89[907], line_88[905], line_87[903], line_86[901], line_85[899], line_84[897], line_83[895], line_82[893], line_81[891], line_80[889], line_79[887], line_78[885], line_77[883], line_76[881], line_75[879], line_74[877], line_73[875], line_72[873], line_71[871], line_70[869], line_69[867], line_68[865], line_67[863], line_66[861], line_65[859], line_64[857], line_63[855], line_62[853], line_61[851], line_60[849], line_59[847], line_58[845], line_57[843], line_56[841], line_55[839], line_54[837], line_53[835], line_52[833], line_51[831], line_50[829], line_49[827], line_48[825], line_47[823], line_46[821], line_45[819], line_44[817], line_43[815], line_42[813], line_41[811], line_40[809], line_39[807], line_38[805], line_37[803], line_36[801], line_35[799], line_34[797], line_33[795], line_32[793], line_31[791], line_30[789], line_29[787], line_28[785], line_27[783], line_26[781], line_25[779], line_24[777], line_23[775], line_22[773], line_21[771], line_20[769], line_19[767], line_18[765], line_17[763], line_16[761], line_15[759], line_14[757], line_13[755], line_12[753], line_11[751], line_10[749], line_9[747], line_8[745], line_7[743], line_6[741], line_5[739], line_4[737], line_3[735], line_2[733], line_1[731] };
assign col_986 = {line_128[986], line_127[984], line_126[982], line_125[980], line_124[978], line_123[976], line_122[974], line_121[972], line_120[970], line_119[968], line_118[966], line_117[964], line_116[962], line_115[960], line_114[958], line_113[956], line_112[954], line_111[952], line_110[950], line_109[948], line_108[946], line_107[944], line_106[942], line_105[940], line_104[938], line_103[936], line_102[934], line_101[932], line_100[930], line_99[928], line_98[926], line_97[924], line_96[922], line_95[920], line_94[918], line_93[916], line_92[914], line_91[912], line_90[910], line_89[908], line_88[906], line_87[904], line_86[902], line_85[900], line_84[898], line_83[896], line_82[894], line_81[892], line_80[890], line_79[888], line_78[886], line_77[884], line_76[882], line_75[880], line_74[878], line_73[876], line_72[874], line_71[872], line_70[870], line_69[868], line_68[866], line_67[864], line_66[862], line_65[860], line_64[858], line_63[856], line_62[854], line_61[852], line_60[850], line_59[848], line_58[846], line_57[844], line_56[842], line_55[840], line_54[838], line_53[836], line_52[834], line_51[832], line_50[830], line_49[828], line_48[826], line_47[824], line_46[822], line_45[820], line_44[818], line_43[816], line_42[814], line_41[812], line_40[810], line_39[808], line_38[806], line_37[804], line_36[802], line_35[800], line_34[798], line_33[796], line_32[794], line_31[792], line_30[790], line_29[788], line_28[786], line_27[784], line_26[782], line_25[780], line_24[778], line_23[776], line_22[774], line_21[772], line_20[770], line_19[768], line_18[766], line_17[764], line_16[762], line_15[760], line_14[758], line_13[756], line_12[754], line_11[752], line_10[750], line_9[748], line_8[746], line_7[744], line_6[742], line_5[740], line_4[738], line_3[736], line_2[734], line_1[732] };
assign col_987 = {line_128[987], line_127[985], line_126[983], line_125[981], line_124[979], line_123[977], line_122[975], line_121[973], line_120[971], line_119[969], line_118[967], line_117[965], line_116[963], line_115[961], line_114[959], line_113[957], line_112[955], line_111[953], line_110[951], line_109[949], line_108[947], line_107[945], line_106[943], line_105[941], line_104[939], line_103[937], line_102[935], line_101[933], line_100[931], line_99[929], line_98[927], line_97[925], line_96[923], line_95[921], line_94[919], line_93[917], line_92[915], line_91[913], line_90[911], line_89[909], line_88[907], line_87[905], line_86[903], line_85[901], line_84[899], line_83[897], line_82[895], line_81[893], line_80[891], line_79[889], line_78[887], line_77[885], line_76[883], line_75[881], line_74[879], line_73[877], line_72[875], line_71[873], line_70[871], line_69[869], line_68[867], line_67[865], line_66[863], line_65[861], line_64[859], line_63[857], line_62[855], line_61[853], line_60[851], line_59[849], line_58[847], line_57[845], line_56[843], line_55[841], line_54[839], line_53[837], line_52[835], line_51[833], line_50[831], line_49[829], line_48[827], line_47[825], line_46[823], line_45[821], line_44[819], line_43[817], line_42[815], line_41[813], line_40[811], line_39[809], line_38[807], line_37[805], line_36[803], line_35[801], line_34[799], line_33[797], line_32[795], line_31[793], line_30[791], line_29[789], line_28[787], line_27[785], line_26[783], line_25[781], line_24[779], line_23[777], line_22[775], line_21[773], line_20[771], line_19[769], line_18[767], line_17[765], line_16[763], line_15[761], line_14[759], line_13[757], line_12[755], line_11[753], line_10[751], line_9[749], line_8[747], line_7[745], line_6[743], line_5[741], line_4[739], line_3[737], line_2[735], line_1[733] };
assign col_988 = {line_128[988], line_127[986], line_126[984], line_125[982], line_124[980], line_123[978], line_122[976], line_121[974], line_120[972], line_119[970], line_118[968], line_117[966], line_116[964], line_115[962], line_114[960], line_113[958], line_112[956], line_111[954], line_110[952], line_109[950], line_108[948], line_107[946], line_106[944], line_105[942], line_104[940], line_103[938], line_102[936], line_101[934], line_100[932], line_99[930], line_98[928], line_97[926], line_96[924], line_95[922], line_94[920], line_93[918], line_92[916], line_91[914], line_90[912], line_89[910], line_88[908], line_87[906], line_86[904], line_85[902], line_84[900], line_83[898], line_82[896], line_81[894], line_80[892], line_79[890], line_78[888], line_77[886], line_76[884], line_75[882], line_74[880], line_73[878], line_72[876], line_71[874], line_70[872], line_69[870], line_68[868], line_67[866], line_66[864], line_65[862], line_64[860], line_63[858], line_62[856], line_61[854], line_60[852], line_59[850], line_58[848], line_57[846], line_56[844], line_55[842], line_54[840], line_53[838], line_52[836], line_51[834], line_50[832], line_49[830], line_48[828], line_47[826], line_46[824], line_45[822], line_44[820], line_43[818], line_42[816], line_41[814], line_40[812], line_39[810], line_38[808], line_37[806], line_36[804], line_35[802], line_34[800], line_33[798], line_32[796], line_31[794], line_30[792], line_29[790], line_28[788], line_27[786], line_26[784], line_25[782], line_24[780], line_23[778], line_22[776], line_21[774], line_20[772], line_19[770], line_18[768], line_17[766], line_16[764], line_15[762], line_14[760], line_13[758], line_12[756], line_11[754], line_10[752], line_9[750], line_8[748], line_7[746], line_6[744], line_5[742], line_4[740], line_3[738], line_2[736], line_1[734] };
assign col_989 = {line_128[989], line_127[987], line_126[985], line_125[983], line_124[981], line_123[979], line_122[977], line_121[975], line_120[973], line_119[971], line_118[969], line_117[967], line_116[965], line_115[963], line_114[961], line_113[959], line_112[957], line_111[955], line_110[953], line_109[951], line_108[949], line_107[947], line_106[945], line_105[943], line_104[941], line_103[939], line_102[937], line_101[935], line_100[933], line_99[931], line_98[929], line_97[927], line_96[925], line_95[923], line_94[921], line_93[919], line_92[917], line_91[915], line_90[913], line_89[911], line_88[909], line_87[907], line_86[905], line_85[903], line_84[901], line_83[899], line_82[897], line_81[895], line_80[893], line_79[891], line_78[889], line_77[887], line_76[885], line_75[883], line_74[881], line_73[879], line_72[877], line_71[875], line_70[873], line_69[871], line_68[869], line_67[867], line_66[865], line_65[863], line_64[861], line_63[859], line_62[857], line_61[855], line_60[853], line_59[851], line_58[849], line_57[847], line_56[845], line_55[843], line_54[841], line_53[839], line_52[837], line_51[835], line_50[833], line_49[831], line_48[829], line_47[827], line_46[825], line_45[823], line_44[821], line_43[819], line_42[817], line_41[815], line_40[813], line_39[811], line_38[809], line_37[807], line_36[805], line_35[803], line_34[801], line_33[799], line_32[797], line_31[795], line_30[793], line_29[791], line_28[789], line_27[787], line_26[785], line_25[783], line_24[781], line_23[779], line_22[777], line_21[775], line_20[773], line_19[771], line_18[769], line_17[767], line_16[765], line_15[763], line_14[761], line_13[759], line_12[757], line_11[755], line_10[753], line_9[751], line_8[749], line_7[747], line_6[745], line_5[743], line_4[741], line_3[739], line_2[737], line_1[735] };
assign col_990 = {line_128[990], line_127[988], line_126[986], line_125[984], line_124[982], line_123[980], line_122[978], line_121[976], line_120[974], line_119[972], line_118[970], line_117[968], line_116[966], line_115[964], line_114[962], line_113[960], line_112[958], line_111[956], line_110[954], line_109[952], line_108[950], line_107[948], line_106[946], line_105[944], line_104[942], line_103[940], line_102[938], line_101[936], line_100[934], line_99[932], line_98[930], line_97[928], line_96[926], line_95[924], line_94[922], line_93[920], line_92[918], line_91[916], line_90[914], line_89[912], line_88[910], line_87[908], line_86[906], line_85[904], line_84[902], line_83[900], line_82[898], line_81[896], line_80[894], line_79[892], line_78[890], line_77[888], line_76[886], line_75[884], line_74[882], line_73[880], line_72[878], line_71[876], line_70[874], line_69[872], line_68[870], line_67[868], line_66[866], line_65[864], line_64[862], line_63[860], line_62[858], line_61[856], line_60[854], line_59[852], line_58[850], line_57[848], line_56[846], line_55[844], line_54[842], line_53[840], line_52[838], line_51[836], line_50[834], line_49[832], line_48[830], line_47[828], line_46[826], line_45[824], line_44[822], line_43[820], line_42[818], line_41[816], line_40[814], line_39[812], line_38[810], line_37[808], line_36[806], line_35[804], line_34[802], line_33[800], line_32[798], line_31[796], line_30[794], line_29[792], line_28[790], line_27[788], line_26[786], line_25[784], line_24[782], line_23[780], line_22[778], line_21[776], line_20[774], line_19[772], line_18[770], line_17[768], line_16[766], line_15[764], line_14[762], line_13[760], line_12[758], line_11[756], line_10[754], line_9[752], line_8[750], line_7[748], line_6[746], line_5[744], line_4[742], line_3[740], line_2[738], line_1[736] };
assign col_991 = {line_128[991], line_127[989], line_126[987], line_125[985], line_124[983], line_123[981], line_122[979], line_121[977], line_120[975], line_119[973], line_118[971], line_117[969], line_116[967], line_115[965], line_114[963], line_113[961], line_112[959], line_111[957], line_110[955], line_109[953], line_108[951], line_107[949], line_106[947], line_105[945], line_104[943], line_103[941], line_102[939], line_101[937], line_100[935], line_99[933], line_98[931], line_97[929], line_96[927], line_95[925], line_94[923], line_93[921], line_92[919], line_91[917], line_90[915], line_89[913], line_88[911], line_87[909], line_86[907], line_85[905], line_84[903], line_83[901], line_82[899], line_81[897], line_80[895], line_79[893], line_78[891], line_77[889], line_76[887], line_75[885], line_74[883], line_73[881], line_72[879], line_71[877], line_70[875], line_69[873], line_68[871], line_67[869], line_66[867], line_65[865], line_64[863], line_63[861], line_62[859], line_61[857], line_60[855], line_59[853], line_58[851], line_57[849], line_56[847], line_55[845], line_54[843], line_53[841], line_52[839], line_51[837], line_50[835], line_49[833], line_48[831], line_47[829], line_46[827], line_45[825], line_44[823], line_43[821], line_42[819], line_41[817], line_40[815], line_39[813], line_38[811], line_37[809], line_36[807], line_35[805], line_34[803], line_33[801], line_32[799], line_31[797], line_30[795], line_29[793], line_28[791], line_27[789], line_26[787], line_25[785], line_24[783], line_23[781], line_22[779], line_21[777], line_20[775], line_19[773], line_18[771], line_17[769], line_16[767], line_15[765], line_14[763], line_13[761], line_12[759], line_11[757], line_10[755], line_9[753], line_8[751], line_7[749], line_6[747], line_5[745], line_4[743], line_3[741], line_2[739], line_1[737] };
assign col_992 = {line_128[992], line_127[990], line_126[988], line_125[986], line_124[984], line_123[982], line_122[980], line_121[978], line_120[976], line_119[974], line_118[972], line_117[970], line_116[968], line_115[966], line_114[964], line_113[962], line_112[960], line_111[958], line_110[956], line_109[954], line_108[952], line_107[950], line_106[948], line_105[946], line_104[944], line_103[942], line_102[940], line_101[938], line_100[936], line_99[934], line_98[932], line_97[930], line_96[928], line_95[926], line_94[924], line_93[922], line_92[920], line_91[918], line_90[916], line_89[914], line_88[912], line_87[910], line_86[908], line_85[906], line_84[904], line_83[902], line_82[900], line_81[898], line_80[896], line_79[894], line_78[892], line_77[890], line_76[888], line_75[886], line_74[884], line_73[882], line_72[880], line_71[878], line_70[876], line_69[874], line_68[872], line_67[870], line_66[868], line_65[866], line_64[864], line_63[862], line_62[860], line_61[858], line_60[856], line_59[854], line_58[852], line_57[850], line_56[848], line_55[846], line_54[844], line_53[842], line_52[840], line_51[838], line_50[836], line_49[834], line_48[832], line_47[830], line_46[828], line_45[826], line_44[824], line_43[822], line_42[820], line_41[818], line_40[816], line_39[814], line_38[812], line_37[810], line_36[808], line_35[806], line_34[804], line_33[802], line_32[800], line_31[798], line_30[796], line_29[794], line_28[792], line_27[790], line_26[788], line_25[786], line_24[784], line_23[782], line_22[780], line_21[778], line_20[776], line_19[774], line_18[772], line_17[770], line_16[768], line_15[766], line_14[764], line_13[762], line_12[760], line_11[758], line_10[756], line_9[754], line_8[752], line_7[750], line_6[748], line_5[746], line_4[744], line_3[742], line_2[740], line_1[738] };
assign col_993 = {line_128[993], line_127[991], line_126[989], line_125[987], line_124[985], line_123[983], line_122[981], line_121[979], line_120[977], line_119[975], line_118[973], line_117[971], line_116[969], line_115[967], line_114[965], line_113[963], line_112[961], line_111[959], line_110[957], line_109[955], line_108[953], line_107[951], line_106[949], line_105[947], line_104[945], line_103[943], line_102[941], line_101[939], line_100[937], line_99[935], line_98[933], line_97[931], line_96[929], line_95[927], line_94[925], line_93[923], line_92[921], line_91[919], line_90[917], line_89[915], line_88[913], line_87[911], line_86[909], line_85[907], line_84[905], line_83[903], line_82[901], line_81[899], line_80[897], line_79[895], line_78[893], line_77[891], line_76[889], line_75[887], line_74[885], line_73[883], line_72[881], line_71[879], line_70[877], line_69[875], line_68[873], line_67[871], line_66[869], line_65[867], line_64[865], line_63[863], line_62[861], line_61[859], line_60[857], line_59[855], line_58[853], line_57[851], line_56[849], line_55[847], line_54[845], line_53[843], line_52[841], line_51[839], line_50[837], line_49[835], line_48[833], line_47[831], line_46[829], line_45[827], line_44[825], line_43[823], line_42[821], line_41[819], line_40[817], line_39[815], line_38[813], line_37[811], line_36[809], line_35[807], line_34[805], line_33[803], line_32[801], line_31[799], line_30[797], line_29[795], line_28[793], line_27[791], line_26[789], line_25[787], line_24[785], line_23[783], line_22[781], line_21[779], line_20[777], line_19[775], line_18[773], line_17[771], line_16[769], line_15[767], line_14[765], line_13[763], line_12[761], line_11[759], line_10[757], line_9[755], line_8[753], line_7[751], line_6[749], line_5[747], line_4[745], line_3[743], line_2[741], line_1[739] };
assign col_994 = {line_128[994], line_127[992], line_126[990], line_125[988], line_124[986], line_123[984], line_122[982], line_121[980], line_120[978], line_119[976], line_118[974], line_117[972], line_116[970], line_115[968], line_114[966], line_113[964], line_112[962], line_111[960], line_110[958], line_109[956], line_108[954], line_107[952], line_106[950], line_105[948], line_104[946], line_103[944], line_102[942], line_101[940], line_100[938], line_99[936], line_98[934], line_97[932], line_96[930], line_95[928], line_94[926], line_93[924], line_92[922], line_91[920], line_90[918], line_89[916], line_88[914], line_87[912], line_86[910], line_85[908], line_84[906], line_83[904], line_82[902], line_81[900], line_80[898], line_79[896], line_78[894], line_77[892], line_76[890], line_75[888], line_74[886], line_73[884], line_72[882], line_71[880], line_70[878], line_69[876], line_68[874], line_67[872], line_66[870], line_65[868], line_64[866], line_63[864], line_62[862], line_61[860], line_60[858], line_59[856], line_58[854], line_57[852], line_56[850], line_55[848], line_54[846], line_53[844], line_52[842], line_51[840], line_50[838], line_49[836], line_48[834], line_47[832], line_46[830], line_45[828], line_44[826], line_43[824], line_42[822], line_41[820], line_40[818], line_39[816], line_38[814], line_37[812], line_36[810], line_35[808], line_34[806], line_33[804], line_32[802], line_31[800], line_30[798], line_29[796], line_28[794], line_27[792], line_26[790], line_25[788], line_24[786], line_23[784], line_22[782], line_21[780], line_20[778], line_19[776], line_18[774], line_17[772], line_16[770], line_15[768], line_14[766], line_13[764], line_12[762], line_11[760], line_10[758], line_9[756], line_8[754], line_7[752], line_6[750], line_5[748], line_4[746], line_3[744], line_2[742], line_1[740] };
assign col_995 = {line_128[995], line_127[993], line_126[991], line_125[989], line_124[987], line_123[985], line_122[983], line_121[981], line_120[979], line_119[977], line_118[975], line_117[973], line_116[971], line_115[969], line_114[967], line_113[965], line_112[963], line_111[961], line_110[959], line_109[957], line_108[955], line_107[953], line_106[951], line_105[949], line_104[947], line_103[945], line_102[943], line_101[941], line_100[939], line_99[937], line_98[935], line_97[933], line_96[931], line_95[929], line_94[927], line_93[925], line_92[923], line_91[921], line_90[919], line_89[917], line_88[915], line_87[913], line_86[911], line_85[909], line_84[907], line_83[905], line_82[903], line_81[901], line_80[899], line_79[897], line_78[895], line_77[893], line_76[891], line_75[889], line_74[887], line_73[885], line_72[883], line_71[881], line_70[879], line_69[877], line_68[875], line_67[873], line_66[871], line_65[869], line_64[867], line_63[865], line_62[863], line_61[861], line_60[859], line_59[857], line_58[855], line_57[853], line_56[851], line_55[849], line_54[847], line_53[845], line_52[843], line_51[841], line_50[839], line_49[837], line_48[835], line_47[833], line_46[831], line_45[829], line_44[827], line_43[825], line_42[823], line_41[821], line_40[819], line_39[817], line_38[815], line_37[813], line_36[811], line_35[809], line_34[807], line_33[805], line_32[803], line_31[801], line_30[799], line_29[797], line_28[795], line_27[793], line_26[791], line_25[789], line_24[787], line_23[785], line_22[783], line_21[781], line_20[779], line_19[777], line_18[775], line_17[773], line_16[771], line_15[769], line_14[767], line_13[765], line_12[763], line_11[761], line_10[759], line_9[757], line_8[755], line_7[753], line_6[751], line_5[749], line_4[747], line_3[745], line_2[743], line_1[741] };
assign col_996 = {line_128[996], line_127[994], line_126[992], line_125[990], line_124[988], line_123[986], line_122[984], line_121[982], line_120[980], line_119[978], line_118[976], line_117[974], line_116[972], line_115[970], line_114[968], line_113[966], line_112[964], line_111[962], line_110[960], line_109[958], line_108[956], line_107[954], line_106[952], line_105[950], line_104[948], line_103[946], line_102[944], line_101[942], line_100[940], line_99[938], line_98[936], line_97[934], line_96[932], line_95[930], line_94[928], line_93[926], line_92[924], line_91[922], line_90[920], line_89[918], line_88[916], line_87[914], line_86[912], line_85[910], line_84[908], line_83[906], line_82[904], line_81[902], line_80[900], line_79[898], line_78[896], line_77[894], line_76[892], line_75[890], line_74[888], line_73[886], line_72[884], line_71[882], line_70[880], line_69[878], line_68[876], line_67[874], line_66[872], line_65[870], line_64[868], line_63[866], line_62[864], line_61[862], line_60[860], line_59[858], line_58[856], line_57[854], line_56[852], line_55[850], line_54[848], line_53[846], line_52[844], line_51[842], line_50[840], line_49[838], line_48[836], line_47[834], line_46[832], line_45[830], line_44[828], line_43[826], line_42[824], line_41[822], line_40[820], line_39[818], line_38[816], line_37[814], line_36[812], line_35[810], line_34[808], line_33[806], line_32[804], line_31[802], line_30[800], line_29[798], line_28[796], line_27[794], line_26[792], line_25[790], line_24[788], line_23[786], line_22[784], line_21[782], line_20[780], line_19[778], line_18[776], line_17[774], line_16[772], line_15[770], line_14[768], line_13[766], line_12[764], line_11[762], line_10[760], line_9[758], line_8[756], line_7[754], line_6[752], line_5[750], line_4[748], line_3[746], line_2[744], line_1[742] };
assign col_997 = {line_128[997], line_127[995], line_126[993], line_125[991], line_124[989], line_123[987], line_122[985], line_121[983], line_120[981], line_119[979], line_118[977], line_117[975], line_116[973], line_115[971], line_114[969], line_113[967], line_112[965], line_111[963], line_110[961], line_109[959], line_108[957], line_107[955], line_106[953], line_105[951], line_104[949], line_103[947], line_102[945], line_101[943], line_100[941], line_99[939], line_98[937], line_97[935], line_96[933], line_95[931], line_94[929], line_93[927], line_92[925], line_91[923], line_90[921], line_89[919], line_88[917], line_87[915], line_86[913], line_85[911], line_84[909], line_83[907], line_82[905], line_81[903], line_80[901], line_79[899], line_78[897], line_77[895], line_76[893], line_75[891], line_74[889], line_73[887], line_72[885], line_71[883], line_70[881], line_69[879], line_68[877], line_67[875], line_66[873], line_65[871], line_64[869], line_63[867], line_62[865], line_61[863], line_60[861], line_59[859], line_58[857], line_57[855], line_56[853], line_55[851], line_54[849], line_53[847], line_52[845], line_51[843], line_50[841], line_49[839], line_48[837], line_47[835], line_46[833], line_45[831], line_44[829], line_43[827], line_42[825], line_41[823], line_40[821], line_39[819], line_38[817], line_37[815], line_36[813], line_35[811], line_34[809], line_33[807], line_32[805], line_31[803], line_30[801], line_29[799], line_28[797], line_27[795], line_26[793], line_25[791], line_24[789], line_23[787], line_22[785], line_21[783], line_20[781], line_19[779], line_18[777], line_17[775], line_16[773], line_15[771], line_14[769], line_13[767], line_12[765], line_11[763], line_10[761], line_9[759], line_8[757], line_7[755], line_6[753], line_5[751], line_4[749], line_3[747], line_2[745], line_1[743] };
assign col_998 = {line_128[998], line_127[996], line_126[994], line_125[992], line_124[990], line_123[988], line_122[986], line_121[984], line_120[982], line_119[980], line_118[978], line_117[976], line_116[974], line_115[972], line_114[970], line_113[968], line_112[966], line_111[964], line_110[962], line_109[960], line_108[958], line_107[956], line_106[954], line_105[952], line_104[950], line_103[948], line_102[946], line_101[944], line_100[942], line_99[940], line_98[938], line_97[936], line_96[934], line_95[932], line_94[930], line_93[928], line_92[926], line_91[924], line_90[922], line_89[920], line_88[918], line_87[916], line_86[914], line_85[912], line_84[910], line_83[908], line_82[906], line_81[904], line_80[902], line_79[900], line_78[898], line_77[896], line_76[894], line_75[892], line_74[890], line_73[888], line_72[886], line_71[884], line_70[882], line_69[880], line_68[878], line_67[876], line_66[874], line_65[872], line_64[870], line_63[868], line_62[866], line_61[864], line_60[862], line_59[860], line_58[858], line_57[856], line_56[854], line_55[852], line_54[850], line_53[848], line_52[846], line_51[844], line_50[842], line_49[840], line_48[838], line_47[836], line_46[834], line_45[832], line_44[830], line_43[828], line_42[826], line_41[824], line_40[822], line_39[820], line_38[818], line_37[816], line_36[814], line_35[812], line_34[810], line_33[808], line_32[806], line_31[804], line_30[802], line_29[800], line_28[798], line_27[796], line_26[794], line_25[792], line_24[790], line_23[788], line_22[786], line_21[784], line_20[782], line_19[780], line_18[778], line_17[776], line_16[774], line_15[772], line_14[770], line_13[768], line_12[766], line_11[764], line_10[762], line_9[760], line_8[758], line_7[756], line_6[754], line_5[752], line_4[750], line_3[748], line_2[746], line_1[744] };
assign col_999 = {line_128[999], line_127[997], line_126[995], line_125[993], line_124[991], line_123[989], line_122[987], line_121[985], line_120[983], line_119[981], line_118[979], line_117[977], line_116[975], line_115[973], line_114[971], line_113[969], line_112[967], line_111[965], line_110[963], line_109[961], line_108[959], line_107[957], line_106[955], line_105[953], line_104[951], line_103[949], line_102[947], line_101[945], line_100[943], line_99[941], line_98[939], line_97[937], line_96[935], line_95[933], line_94[931], line_93[929], line_92[927], line_91[925], line_90[923], line_89[921], line_88[919], line_87[917], line_86[915], line_85[913], line_84[911], line_83[909], line_82[907], line_81[905], line_80[903], line_79[901], line_78[899], line_77[897], line_76[895], line_75[893], line_74[891], line_73[889], line_72[887], line_71[885], line_70[883], line_69[881], line_68[879], line_67[877], line_66[875], line_65[873], line_64[871], line_63[869], line_62[867], line_61[865], line_60[863], line_59[861], line_58[859], line_57[857], line_56[855], line_55[853], line_54[851], line_53[849], line_52[847], line_51[845], line_50[843], line_49[841], line_48[839], line_47[837], line_46[835], line_45[833], line_44[831], line_43[829], line_42[827], line_41[825], line_40[823], line_39[821], line_38[819], line_37[817], line_36[815], line_35[813], line_34[811], line_33[809], line_32[807], line_31[805], line_30[803], line_29[801], line_28[799], line_27[797], line_26[795], line_25[793], line_24[791], line_23[789], line_22[787], line_21[785], line_20[783], line_19[781], line_18[779], line_17[777], line_16[775], line_15[773], line_14[771], line_13[769], line_12[767], line_11[765], line_10[763], line_9[761], line_8[759], line_7[757], line_6[755], line_5[753], line_4[751], line_3[749], line_2[747], line_1[745] };
assign col_1000 = {line_128[1000], line_127[998], line_126[996], line_125[994], line_124[992], line_123[990], line_122[988], line_121[986], line_120[984], line_119[982], line_118[980], line_117[978], line_116[976], line_115[974], line_114[972], line_113[970], line_112[968], line_111[966], line_110[964], line_109[962], line_108[960], line_107[958], line_106[956], line_105[954], line_104[952], line_103[950], line_102[948], line_101[946], line_100[944], line_99[942], line_98[940], line_97[938], line_96[936], line_95[934], line_94[932], line_93[930], line_92[928], line_91[926], line_90[924], line_89[922], line_88[920], line_87[918], line_86[916], line_85[914], line_84[912], line_83[910], line_82[908], line_81[906], line_80[904], line_79[902], line_78[900], line_77[898], line_76[896], line_75[894], line_74[892], line_73[890], line_72[888], line_71[886], line_70[884], line_69[882], line_68[880], line_67[878], line_66[876], line_65[874], line_64[872], line_63[870], line_62[868], line_61[866], line_60[864], line_59[862], line_58[860], line_57[858], line_56[856], line_55[854], line_54[852], line_53[850], line_52[848], line_51[846], line_50[844], line_49[842], line_48[840], line_47[838], line_46[836], line_45[834], line_44[832], line_43[830], line_42[828], line_41[826], line_40[824], line_39[822], line_38[820], line_37[818], line_36[816], line_35[814], line_34[812], line_33[810], line_32[808], line_31[806], line_30[804], line_29[802], line_28[800], line_27[798], line_26[796], line_25[794], line_24[792], line_23[790], line_22[788], line_21[786], line_20[784], line_19[782], line_18[780], line_17[778], line_16[776], line_15[774], line_14[772], line_13[770], line_12[768], line_11[766], line_10[764], line_9[762], line_8[760], line_7[758], line_6[756], line_5[754], line_4[752], line_3[750], line_2[748], line_1[746] };
assign col_1001 = {line_128[1001], line_127[999], line_126[997], line_125[995], line_124[993], line_123[991], line_122[989], line_121[987], line_120[985], line_119[983], line_118[981], line_117[979], line_116[977], line_115[975], line_114[973], line_113[971], line_112[969], line_111[967], line_110[965], line_109[963], line_108[961], line_107[959], line_106[957], line_105[955], line_104[953], line_103[951], line_102[949], line_101[947], line_100[945], line_99[943], line_98[941], line_97[939], line_96[937], line_95[935], line_94[933], line_93[931], line_92[929], line_91[927], line_90[925], line_89[923], line_88[921], line_87[919], line_86[917], line_85[915], line_84[913], line_83[911], line_82[909], line_81[907], line_80[905], line_79[903], line_78[901], line_77[899], line_76[897], line_75[895], line_74[893], line_73[891], line_72[889], line_71[887], line_70[885], line_69[883], line_68[881], line_67[879], line_66[877], line_65[875], line_64[873], line_63[871], line_62[869], line_61[867], line_60[865], line_59[863], line_58[861], line_57[859], line_56[857], line_55[855], line_54[853], line_53[851], line_52[849], line_51[847], line_50[845], line_49[843], line_48[841], line_47[839], line_46[837], line_45[835], line_44[833], line_43[831], line_42[829], line_41[827], line_40[825], line_39[823], line_38[821], line_37[819], line_36[817], line_35[815], line_34[813], line_33[811], line_32[809], line_31[807], line_30[805], line_29[803], line_28[801], line_27[799], line_26[797], line_25[795], line_24[793], line_23[791], line_22[789], line_21[787], line_20[785], line_19[783], line_18[781], line_17[779], line_16[777], line_15[775], line_14[773], line_13[771], line_12[769], line_11[767], line_10[765], line_9[763], line_8[761], line_7[759], line_6[757], line_5[755], line_4[753], line_3[751], line_2[749], line_1[747] };
assign col_1002 = {line_128[1002], line_127[1000], line_126[998], line_125[996], line_124[994], line_123[992], line_122[990], line_121[988], line_120[986], line_119[984], line_118[982], line_117[980], line_116[978], line_115[976], line_114[974], line_113[972], line_112[970], line_111[968], line_110[966], line_109[964], line_108[962], line_107[960], line_106[958], line_105[956], line_104[954], line_103[952], line_102[950], line_101[948], line_100[946], line_99[944], line_98[942], line_97[940], line_96[938], line_95[936], line_94[934], line_93[932], line_92[930], line_91[928], line_90[926], line_89[924], line_88[922], line_87[920], line_86[918], line_85[916], line_84[914], line_83[912], line_82[910], line_81[908], line_80[906], line_79[904], line_78[902], line_77[900], line_76[898], line_75[896], line_74[894], line_73[892], line_72[890], line_71[888], line_70[886], line_69[884], line_68[882], line_67[880], line_66[878], line_65[876], line_64[874], line_63[872], line_62[870], line_61[868], line_60[866], line_59[864], line_58[862], line_57[860], line_56[858], line_55[856], line_54[854], line_53[852], line_52[850], line_51[848], line_50[846], line_49[844], line_48[842], line_47[840], line_46[838], line_45[836], line_44[834], line_43[832], line_42[830], line_41[828], line_40[826], line_39[824], line_38[822], line_37[820], line_36[818], line_35[816], line_34[814], line_33[812], line_32[810], line_31[808], line_30[806], line_29[804], line_28[802], line_27[800], line_26[798], line_25[796], line_24[794], line_23[792], line_22[790], line_21[788], line_20[786], line_19[784], line_18[782], line_17[780], line_16[778], line_15[776], line_14[774], line_13[772], line_12[770], line_11[768], line_10[766], line_9[764], line_8[762], line_7[760], line_6[758], line_5[756], line_4[754], line_3[752], line_2[750], line_1[748] };
assign col_1003 = {line_128[1003], line_127[1001], line_126[999], line_125[997], line_124[995], line_123[993], line_122[991], line_121[989], line_120[987], line_119[985], line_118[983], line_117[981], line_116[979], line_115[977], line_114[975], line_113[973], line_112[971], line_111[969], line_110[967], line_109[965], line_108[963], line_107[961], line_106[959], line_105[957], line_104[955], line_103[953], line_102[951], line_101[949], line_100[947], line_99[945], line_98[943], line_97[941], line_96[939], line_95[937], line_94[935], line_93[933], line_92[931], line_91[929], line_90[927], line_89[925], line_88[923], line_87[921], line_86[919], line_85[917], line_84[915], line_83[913], line_82[911], line_81[909], line_80[907], line_79[905], line_78[903], line_77[901], line_76[899], line_75[897], line_74[895], line_73[893], line_72[891], line_71[889], line_70[887], line_69[885], line_68[883], line_67[881], line_66[879], line_65[877], line_64[875], line_63[873], line_62[871], line_61[869], line_60[867], line_59[865], line_58[863], line_57[861], line_56[859], line_55[857], line_54[855], line_53[853], line_52[851], line_51[849], line_50[847], line_49[845], line_48[843], line_47[841], line_46[839], line_45[837], line_44[835], line_43[833], line_42[831], line_41[829], line_40[827], line_39[825], line_38[823], line_37[821], line_36[819], line_35[817], line_34[815], line_33[813], line_32[811], line_31[809], line_30[807], line_29[805], line_28[803], line_27[801], line_26[799], line_25[797], line_24[795], line_23[793], line_22[791], line_21[789], line_20[787], line_19[785], line_18[783], line_17[781], line_16[779], line_15[777], line_14[775], line_13[773], line_12[771], line_11[769], line_10[767], line_9[765], line_8[763], line_7[761], line_6[759], line_5[757], line_4[755], line_3[753], line_2[751], line_1[749] };
assign col_1004 = {line_128[1004], line_127[1002], line_126[1000], line_125[998], line_124[996], line_123[994], line_122[992], line_121[990], line_120[988], line_119[986], line_118[984], line_117[982], line_116[980], line_115[978], line_114[976], line_113[974], line_112[972], line_111[970], line_110[968], line_109[966], line_108[964], line_107[962], line_106[960], line_105[958], line_104[956], line_103[954], line_102[952], line_101[950], line_100[948], line_99[946], line_98[944], line_97[942], line_96[940], line_95[938], line_94[936], line_93[934], line_92[932], line_91[930], line_90[928], line_89[926], line_88[924], line_87[922], line_86[920], line_85[918], line_84[916], line_83[914], line_82[912], line_81[910], line_80[908], line_79[906], line_78[904], line_77[902], line_76[900], line_75[898], line_74[896], line_73[894], line_72[892], line_71[890], line_70[888], line_69[886], line_68[884], line_67[882], line_66[880], line_65[878], line_64[876], line_63[874], line_62[872], line_61[870], line_60[868], line_59[866], line_58[864], line_57[862], line_56[860], line_55[858], line_54[856], line_53[854], line_52[852], line_51[850], line_50[848], line_49[846], line_48[844], line_47[842], line_46[840], line_45[838], line_44[836], line_43[834], line_42[832], line_41[830], line_40[828], line_39[826], line_38[824], line_37[822], line_36[820], line_35[818], line_34[816], line_33[814], line_32[812], line_31[810], line_30[808], line_29[806], line_28[804], line_27[802], line_26[800], line_25[798], line_24[796], line_23[794], line_22[792], line_21[790], line_20[788], line_19[786], line_18[784], line_17[782], line_16[780], line_15[778], line_14[776], line_13[774], line_12[772], line_11[770], line_10[768], line_9[766], line_8[764], line_7[762], line_6[760], line_5[758], line_4[756], line_3[754], line_2[752], line_1[750] };
assign col_1005 = {line_128[1005], line_127[1003], line_126[1001], line_125[999], line_124[997], line_123[995], line_122[993], line_121[991], line_120[989], line_119[987], line_118[985], line_117[983], line_116[981], line_115[979], line_114[977], line_113[975], line_112[973], line_111[971], line_110[969], line_109[967], line_108[965], line_107[963], line_106[961], line_105[959], line_104[957], line_103[955], line_102[953], line_101[951], line_100[949], line_99[947], line_98[945], line_97[943], line_96[941], line_95[939], line_94[937], line_93[935], line_92[933], line_91[931], line_90[929], line_89[927], line_88[925], line_87[923], line_86[921], line_85[919], line_84[917], line_83[915], line_82[913], line_81[911], line_80[909], line_79[907], line_78[905], line_77[903], line_76[901], line_75[899], line_74[897], line_73[895], line_72[893], line_71[891], line_70[889], line_69[887], line_68[885], line_67[883], line_66[881], line_65[879], line_64[877], line_63[875], line_62[873], line_61[871], line_60[869], line_59[867], line_58[865], line_57[863], line_56[861], line_55[859], line_54[857], line_53[855], line_52[853], line_51[851], line_50[849], line_49[847], line_48[845], line_47[843], line_46[841], line_45[839], line_44[837], line_43[835], line_42[833], line_41[831], line_40[829], line_39[827], line_38[825], line_37[823], line_36[821], line_35[819], line_34[817], line_33[815], line_32[813], line_31[811], line_30[809], line_29[807], line_28[805], line_27[803], line_26[801], line_25[799], line_24[797], line_23[795], line_22[793], line_21[791], line_20[789], line_19[787], line_18[785], line_17[783], line_16[781], line_15[779], line_14[777], line_13[775], line_12[773], line_11[771], line_10[769], line_9[767], line_8[765], line_7[763], line_6[761], line_5[759], line_4[757], line_3[755], line_2[753], line_1[751] };
assign col_1006 = {line_128[1006], line_127[1004], line_126[1002], line_125[1000], line_124[998], line_123[996], line_122[994], line_121[992], line_120[990], line_119[988], line_118[986], line_117[984], line_116[982], line_115[980], line_114[978], line_113[976], line_112[974], line_111[972], line_110[970], line_109[968], line_108[966], line_107[964], line_106[962], line_105[960], line_104[958], line_103[956], line_102[954], line_101[952], line_100[950], line_99[948], line_98[946], line_97[944], line_96[942], line_95[940], line_94[938], line_93[936], line_92[934], line_91[932], line_90[930], line_89[928], line_88[926], line_87[924], line_86[922], line_85[920], line_84[918], line_83[916], line_82[914], line_81[912], line_80[910], line_79[908], line_78[906], line_77[904], line_76[902], line_75[900], line_74[898], line_73[896], line_72[894], line_71[892], line_70[890], line_69[888], line_68[886], line_67[884], line_66[882], line_65[880], line_64[878], line_63[876], line_62[874], line_61[872], line_60[870], line_59[868], line_58[866], line_57[864], line_56[862], line_55[860], line_54[858], line_53[856], line_52[854], line_51[852], line_50[850], line_49[848], line_48[846], line_47[844], line_46[842], line_45[840], line_44[838], line_43[836], line_42[834], line_41[832], line_40[830], line_39[828], line_38[826], line_37[824], line_36[822], line_35[820], line_34[818], line_33[816], line_32[814], line_31[812], line_30[810], line_29[808], line_28[806], line_27[804], line_26[802], line_25[800], line_24[798], line_23[796], line_22[794], line_21[792], line_20[790], line_19[788], line_18[786], line_17[784], line_16[782], line_15[780], line_14[778], line_13[776], line_12[774], line_11[772], line_10[770], line_9[768], line_8[766], line_7[764], line_6[762], line_5[760], line_4[758], line_3[756], line_2[754], line_1[752] };
assign col_1007 = {line_128[1007], line_127[1005], line_126[1003], line_125[1001], line_124[999], line_123[997], line_122[995], line_121[993], line_120[991], line_119[989], line_118[987], line_117[985], line_116[983], line_115[981], line_114[979], line_113[977], line_112[975], line_111[973], line_110[971], line_109[969], line_108[967], line_107[965], line_106[963], line_105[961], line_104[959], line_103[957], line_102[955], line_101[953], line_100[951], line_99[949], line_98[947], line_97[945], line_96[943], line_95[941], line_94[939], line_93[937], line_92[935], line_91[933], line_90[931], line_89[929], line_88[927], line_87[925], line_86[923], line_85[921], line_84[919], line_83[917], line_82[915], line_81[913], line_80[911], line_79[909], line_78[907], line_77[905], line_76[903], line_75[901], line_74[899], line_73[897], line_72[895], line_71[893], line_70[891], line_69[889], line_68[887], line_67[885], line_66[883], line_65[881], line_64[879], line_63[877], line_62[875], line_61[873], line_60[871], line_59[869], line_58[867], line_57[865], line_56[863], line_55[861], line_54[859], line_53[857], line_52[855], line_51[853], line_50[851], line_49[849], line_48[847], line_47[845], line_46[843], line_45[841], line_44[839], line_43[837], line_42[835], line_41[833], line_40[831], line_39[829], line_38[827], line_37[825], line_36[823], line_35[821], line_34[819], line_33[817], line_32[815], line_31[813], line_30[811], line_29[809], line_28[807], line_27[805], line_26[803], line_25[801], line_24[799], line_23[797], line_22[795], line_21[793], line_20[791], line_19[789], line_18[787], line_17[785], line_16[783], line_15[781], line_14[779], line_13[777], line_12[775], line_11[773], line_10[771], line_9[769], line_8[767], line_7[765], line_6[763], line_5[761], line_4[759], line_3[757], line_2[755], line_1[753] };
assign col_1008 = {line_128[1008], line_127[1006], line_126[1004], line_125[1002], line_124[1000], line_123[998], line_122[996], line_121[994], line_120[992], line_119[990], line_118[988], line_117[986], line_116[984], line_115[982], line_114[980], line_113[978], line_112[976], line_111[974], line_110[972], line_109[970], line_108[968], line_107[966], line_106[964], line_105[962], line_104[960], line_103[958], line_102[956], line_101[954], line_100[952], line_99[950], line_98[948], line_97[946], line_96[944], line_95[942], line_94[940], line_93[938], line_92[936], line_91[934], line_90[932], line_89[930], line_88[928], line_87[926], line_86[924], line_85[922], line_84[920], line_83[918], line_82[916], line_81[914], line_80[912], line_79[910], line_78[908], line_77[906], line_76[904], line_75[902], line_74[900], line_73[898], line_72[896], line_71[894], line_70[892], line_69[890], line_68[888], line_67[886], line_66[884], line_65[882], line_64[880], line_63[878], line_62[876], line_61[874], line_60[872], line_59[870], line_58[868], line_57[866], line_56[864], line_55[862], line_54[860], line_53[858], line_52[856], line_51[854], line_50[852], line_49[850], line_48[848], line_47[846], line_46[844], line_45[842], line_44[840], line_43[838], line_42[836], line_41[834], line_40[832], line_39[830], line_38[828], line_37[826], line_36[824], line_35[822], line_34[820], line_33[818], line_32[816], line_31[814], line_30[812], line_29[810], line_28[808], line_27[806], line_26[804], line_25[802], line_24[800], line_23[798], line_22[796], line_21[794], line_20[792], line_19[790], line_18[788], line_17[786], line_16[784], line_15[782], line_14[780], line_13[778], line_12[776], line_11[774], line_10[772], line_9[770], line_8[768], line_7[766], line_6[764], line_5[762], line_4[760], line_3[758], line_2[756], line_1[754] };
assign col_1009 = {line_128[1009], line_127[1007], line_126[1005], line_125[1003], line_124[1001], line_123[999], line_122[997], line_121[995], line_120[993], line_119[991], line_118[989], line_117[987], line_116[985], line_115[983], line_114[981], line_113[979], line_112[977], line_111[975], line_110[973], line_109[971], line_108[969], line_107[967], line_106[965], line_105[963], line_104[961], line_103[959], line_102[957], line_101[955], line_100[953], line_99[951], line_98[949], line_97[947], line_96[945], line_95[943], line_94[941], line_93[939], line_92[937], line_91[935], line_90[933], line_89[931], line_88[929], line_87[927], line_86[925], line_85[923], line_84[921], line_83[919], line_82[917], line_81[915], line_80[913], line_79[911], line_78[909], line_77[907], line_76[905], line_75[903], line_74[901], line_73[899], line_72[897], line_71[895], line_70[893], line_69[891], line_68[889], line_67[887], line_66[885], line_65[883], line_64[881], line_63[879], line_62[877], line_61[875], line_60[873], line_59[871], line_58[869], line_57[867], line_56[865], line_55[863], line_54[861], line_53[859], line_52[857], line_51[855], line_50[853], line_49[851], line_48[849], line_47[847], line_46[845], line_45[843], line_44[841], line_43[839], line_42[837], line_41[835], line_40[833], line_39[831], line_38[829], line_37[827], line_36[825], line_35[823], line_34[821], line_33[819], line_32[817], line_31[815], line_30[813], line_29[811], line_28[809], line_27[807], line_26[805], line_25[803], line_24[801], line_23[799], line_22[797], line_21[795], line_20[793], line_19[791], line_18[789], line_17[787], line_16[785], line_15[783], line_14[781], line_13[779], line_12[777], line_11[775], line_10[773], line_9[771], line_8[769], line_7[767], line_6[765], line_5[763], line_4[761], line_3[759], line_2[757], line_1[755] };
assign col_1010 = {line_128[1010], line_127[1008], line_126[1006], line_125[1004], line_124[1002], line_123[1000], line_122[998], line_121[996], line_120[994], line_119[992], line_118[990], line_117[988], line_116[986], line_115[984], line_114[982], line_113[980], line_112[978], line_111[976], line_110[974], line_109[972], line_108[970], line_107[968], line_106[966], line_105[964], line_104[962], line_103[960], line_102[958], line_101[956], line_100[954], line_99[952], line_98[950], line_97[948], line_96[946], line_95[944], line_94[942], line_93[940], line_92[938], line_91[936], line_90[934], line_89[932], line_88[930], line_87[928], line_86[926], line_85[924], line_84[922], line_83[920], line_82[918], line_81[916], line_80[914], line_79[912], line_78[910], line_77[908], line_76[906], line_75[904], line_74[902], line_73[900], line_72[898], line_71[896], line_70[894], line_69[892], line_68[890], line_67[888], line_66[886], line_65[884], line_64[882], line_63[880], line_62[878], line_61[876], line_60[874], line_59[872], line_58[870], line_57[868], line_56[866], line_55[864], line_54[862], line_53[860], line_52[858], line_51[856], line_50[854], line_49[852], line_48[850], line_47[848], line_46[846], line_45[844], line_44[842], line_43[840], line_42[838], line_41[836], line_40[834], line_39[832], line_38[830], line_37[828], line_36[826], line_35[824], line_34[822], line_33[820], line_32[818], line_31[816], line_30[814], line_29[812], line_28[810], line_27[808], line_26[806], line_25[804], line_24[802], line_23[800], line_22[798], line_21[796], line_20[794], line_19[792], line_18[790], line_17[788], line_16[786], line_15[784], line_14[782], line_13[780], line_12[778], line_11[776], line_10[774], line_9[772], line_8[770], line_7[768], line_6[766], line_5[764], line_4[762], line_3[760], line_2[758], line_1[756] };
assign col_1011 = {line_128[1011], line_127[1009], line_126[1007], line_125[1005], line_124[1003], line_123[1001], line_122[999], line_121[997], line_120[995], line_119[993], line_118[991], line_117[989], line_116[987], line_115[985], line_114[983], line_113[981], line_112[979], line_111[977], line_110[975], line_109[973], line_108[971], line_107[969], line_106[967], line_105[965], line_104[963], line_103[961], line_102[959], line_101[957], line_100[955], line_99[953], line_98[951], line_97[949], line_96[947], line_95[945], line_94[943], line_93[941], line_92[939], line_91[937], line_90[935], line_89[933], line_88[931], line_87[929], line_86[927], line_85[925], line_84[923], line_83[921], line_82[919], line_81[917], line_80[915], line_79[913], line_78[911], line_77[909], line_76[907], line_75[905], line_74[903], line_73[901], line_72[899], line_71[897], line_70[895], line_69[893], line_68[891], line_67[889], line_66[887], line_65[885], line_64[883], line_63[881], line_62[879], line_61[877], line_60[875], line_59[873], line_58[871], line_57[869], line_56[867], line_55[865], line_54[863], line_53[861], line_52[859], line_51[857], line_50[855], line_49[853], line_48[851], line_47[849], line_46[847], line_45[845], line_44[843], line_43[841], line_42[839], line_41[837], line_40[835], line_39[833], line_38[831], line_37[829], line_36[827], line_35[825], line_34[823], line_33[821], line_32[819], line_31[817], line_30[815], line_29[813], line_28[811], line_27[809], line_26[807], line_25[805], line_24[803], line_23[801], line_22[799], line_21[797], line_20[795], line_19[793], line_18[791], line_17[789], line_16[787], line_15[785], line_14[783], line_13[781], line_12[779], line_11[777], line_10[775], line_9[773], line_8[771], line_7[769], line_6[767], line_5[765], line_4[763], line_3[761], line_2[759], line_1[757] };
assign col_1012 = {line_128[1012], line_127[1010], line_126[1008], line_125[1006], line_124[1004], line_123[1002], line_122[1000], line_121[998], line_120[996], line_119[994], line_118[992], line_117[990], line_116[988], line_115[986], line_114[984], line_113[982], line_112[980], line_111[978], line_110[976], line_109[974], line_108[972], line_107[970], line_106[968], line_105[966], line_104[964], line_103[962], line_102[960], line_101[958], line_100[956], line_99[954], line_98[952], line_97[950], line_96[948], line_95[946], line_94[944], line_93[942], line_92[940], line_91[938], line_90[936], line_89[934], line_88[932], line_87[930], line_86[928], line_85[926], line_84[924], line_83[922], line_82[920], line_81[918], line_80[916], line_79[914], line_78[912], line_77[910], line_76[908], line_75[906], line_74[904], line_73[902], line_72[900], line_71[898], line_70[896], line_69[894], line_68[892], line_67[890], line_66[888], line_65[886], line_64[884], line_63[882], line_62[880], line_61[878], line_60[876], line_59[874], line_58[872], line_57[870], line_56[868], line_55[866], line_54[864], line_53[862], line_52[860], line_51[858], line_50[856], line_49[854], line_48[852], line_47[850], line_46[848], line_45[846], line_44[844], line_43[842], line_42[840], line_41[838], line_40[836], line_39[834], line_38[832], line_37[830], line_36[828], line_35[826], line_34[824], line_33[822], line_32[820], line_31[818], line_30[816], line_29[814], line_28[812], line_27[810], line_26[808], line_25[806], line_24[804], line_23[802], line_22[800], line_21[798], line_20[796], line_19[794], line_18[792], line_17[790], line_16[788], line_15[786], line_14[784], line_13[782], line_12[780], line_11[778], line_10[776], line_9[774], line_8[772], line_7[770], line_6[768], line_5[766], line_4[764], line_3[762], line_2[760], line_1[758] };
assign col_1013 = {line_128[1013], line_127[1011], line_126[1009], line_125[1007], line_124[1005], line_123[1003], line_122[1001], line_121[999], line_120[997], line_119[995], line_118[993], line_117[991], line_116[989], line_115[987], line_114[985], line_113[983], line_112[981], line_111[979], line_110[977], line_109[975], line_108[973], line_107[971], line_106[969], line_105[967], line_104[965], line_103[963], line_102[961], line_101[959], line_100[957], line_99[955], line_98[953], line_97[951], line_96[949], line_95[947], line_94[945], line_93[943], line_92[941], line_91[939], line_90[937], line_89[935], line_88[933], line_87[931], line_86[929], line_85[927], line_84[925], line_83[923], line_82[921], line_81[919], line_80[917], line_79[915], line_78[913], line_77[911], line_76[909], line_75[907], line_74[905], line_73[903], line_72[901], line_71[899], line_70[897], line_69[895], line_68[893], line_67[891], line_66[889], line_65[887], line_64[885], line_63[883], line_62[881], line_61[879], line_60[877], line_59[875], line_58[873], line_57[871], line_56[869], line_55[867], line_54[865], line_53[863], line_52[861], line_51[859], line_50[857], line_49[855], line_48[853], line_47[851], line_46[849], line_45[847], line_44[845], line_43[843], line_42[841], line_41[839], line_40[837], line_39[835], line_38[833], line_37[831], line_36[829], line_35[827], line_34[825], line_33[823], line_32[821], line_31[819], line_30[817], line_29[815], line_28[813], line_27[811], line_26[809], line_25[807], line_24[805], line_23[803], line_22[801], line_21[799], line_20[797], line_19[795], line_18[793], line_17[791], line_16[789], line_15[787], line_14[785], line_13[783], line_12[781], line_11[779], line_10[777], line_9[775], line_8[773], line_7[771], line_6[769], line_5[767], line_4[765], line_3[763], line_2[761], line_1[759] };
assign col_1014 = {line_128[1014], line_127[1012], line_126[1010], line_125[1008], line_124[1006], line_123[1004], line_122[1002], line_121[1000], line_120[998], line_119[996], line_118[994], line_117[992], line_116[990], line_115[988], line_114[986], line_113[984], line_112[982], line_111[980], line_110[978], line_109[976], line_108[974], line_107[972], line_106[970], line_105[968], line_104[966], line_103[964], line_102[962], line_101[960], line_100[958], line_99[956], line_98[954], line_97[952], line_96[950], line_95[948], line_94[946], line_93[944], line_92[942], line_91[940], line_90[938], line_89[936], line_88[934], line_87[932], line_86[930], line_85[928], line_84[926], line_83[924], line_82[922], line_81[920], line_80[918], line_79[916], line_78[914], line_77[912], line_76[910], line_75[908], line_74[906], line_73[904], line_72[902], line_71[900], line_70[898], line_69[896], line_68[894], line_67[892], line_66[890], line_65[888], line_64[886], line_63[884], line_62[882], line_61[880], line_60[878], line_59[876], line_58[874], line_57[872], line_56[870], line_55[868], line_54[866], line_53[864], line_52[862], line_51[860], line_50[858], line_49[856], line_48[854], line_47[852], line_46[850], line_45[848], line_44[846], line_43[844], line_42[842], line_41[840], line_40[838], line_39[836], line_38[834], line_37[832], line_36[830], line_35[828], line_34[826], line_33[824], line_32[822], line_31[820], line_30[818], line_29[816], line_28[814], line_27[812], line_26[810], line_25[808], line_24[806], line_23[804], line_22[802], line_21[800], line_20[798], line_19[796], line_18[794], line_17[792], line_16[790], line_15[788], line_14[786], line_13[784], line_12[782], line_11[780], line_10[778], line_9[776], line_8[774], line_7[772], line_6[770], line_5[768], line_4[766], line_3[764], line_2[762], line_1[760] };
assign col_1015 = {line_128[1015], line_127[1013], line_126[1011], line_125[1009], line_124[1007], line_123[1005], line_122[1003], line_121[1001], line_120[999], line_119[997], line_118[995], line_117[993], line_116[991], line_115[989], line_114[987], line_113[985], line_112[983], line_111[981], line_110[979], line_109[977], line_108[975], line_107[973], line_106[971], line_105[969], line_104[967], line_103[965], line_102[963], line_101[961], line_100[959], line_99[957], line_98[955], line_97[953], line_96[951], line_95[949], line_94[947], line_93[945], line_92[943], line_91[941], line_90[939], line_89[937], line_88[935], line_87[933], line_86[931], line_85[929], line_84[927], line_83[925], line_82[923], line_81[921], line_80[919], line_79[917], line_78[915], line_77[913], line_76[911], line_75[909], line_74[907], line_73[905], line_72[903], line_71[901], line_70[899], line_69[897], line_68[895], line_67[893], line_66[891], line_65[889], line_64[887], line_63[885], line_62[883], line_61[881], line_60[879], line_59[877], line_58[875], line_57[873], line_56[871], line_55[869], line_54[867], line_53[865], line_52[863], line_51[861], line_50[859], line_49[857], line_48[855], line_47[853], line_46[851], line_45[849], line_44[847], line_43[845], line_42[843], line_41[841], line_40[839], line_39[837], line_38[835], line_37[833], line_36[831], line_35[829], line_34[827], line_33[825], line_32[823], line_31[821], line_30[819], line_29[817], line_28[815], line_27[813], line_26[811], line_25[809], line_24[807], line_23[805], line_22[803], line_21[801], line_20[799], line_19[797], line_18[795], line_17[793], line_16[791], line_15[789], line_14[787], line_13[785], line_12[783], line_11[781], line_10[779], line_9[777], line_8[775], line_7[773], line_6[771], line_5[769], line_4[767], line_3[765], line_2[763], line_1[761] };
assign col_1016 = {line_128[1016], line_127[1014], line_126[1012], line_125[1010], line_124[1008], line_123[1006], line_122[1004], line_121[1002], line_120[1000], line_119[998], line_118[996], line_117[994], line_116[992], line_115[990], line_114[988], line_113[986], line_112[984], line_111[982], line_110[980], line_109[978], line_108[976], line_107[974], line_106[972], line_105[970], line_104[968], line_103[966], line_102[964], line_101[962], line_100[960], line_99[958], line_98[956], line_97[954], line_96[952], line_95[950], line_94[948], line_93[946], line_92[944], line_91[942], line_90[940], line_89[938], line_88[936], line_87[934], line_86[932], line_85[930], line_84[928], line_83[926], line_82[924], line_81[922], line_80[920], line_79[918], line_78[916], line_77[914], line_76[912], line_75[910], line_74[908], line_73[906], line_72[904], line_71[902], line_70[900], line_69[898], line_68[896], line_67[894], line_66[892], line_65[890], line_64[888], line_63[886], line_62[884], line_61[882], line_60[880], line_59[878], line_58[876], line_57[874], line_56[872], line_55[870], line_54[868], line_53[866], line_52[864], line_51[862], line_50[860], line_49[858], line_48[856], line_47[854], line_46[852], line_45[850], line_44[848], line_43[846], line_42[844], line_41[842], line_40[840], line_39[838], line_38[836], line_37[834], line_36[832], line_35[830], line_34[828], line_33[826], line_32[824], line_31[822], line_30[820], line_29[818], line_28[816], line_27[814], line_26[812], line_25[810], line_24[808], line_23[806], line_22[804], line_21[802], line_20[800], line_19[798], line_18[796], line_17[794], line_16[792], line_15[790], line_14[788], line_13[786], line_12[784], line_11[782], line_10[780], line_9[778], line_8[776], line_7[774], line_6[772], line_5[770], line_4[768], line_3[766], line_2[764], line_1[762] };
assign col_1017 = {line_128[1017], line_127[1015], line_126[1013], line_125[1011], line_124[1009], line_123[1007], line_122[1005], line_121[1003], line_120[1001], line_119[999], line_118[997], line_117[995], line_116[993], line_115[991], line_114[989], line_113[987], line_112[985], line_111[983], line_110[981], line_109[979], line_108[977], line_107[975], line_106[973], line_105[971], line_104[969], line_103[967], line_102[965], line_101[963], line_100[961], line_99[959], line_98[957], line_97[955], line_96[953], line_95[951], line_94[949], line_93[947], line_92[945], line_91[943], line_90[941], line_89[939], line_88[937], line_87[935], line_86[933], line_85[931], line_84[929], line_83[927], line_82[925], line_81[923], line_80[921], line_79[919], line_78[917], line_77[915], line_76[913], line_75[911], line_74[909], line_73[907], line_72[905], line_71[903], line_70[901], line_69[899], line_68[897], line_67[895], line_66[893], line_65[891], line_64[889], line_63[887], line_62[885], line_61[883], line_60[881], line_59[879], line_58[877], line_57[875], line_56[873], line_55[871], line_54[869], line_53[867], line_52[865], line_51[863], line_50[861], line_49[859], line_48[857], line_47[855], line_46[853], line_45[851], line_44[849], line_43[847], line_42[845], line_41[843], line_40[841], line_39[839], line_38[837], line_37[835], line_36[833], line_35[831], line_34[829], line_33[827], line_32[825], line_31[823], line_30[821], line_29[819], line_28[817], line_27[815], line_26[813], line_25[811], line_24[809], line_23[807], line_22[805], line_21[803], line_20[801], line_19[799], line_18[797], line_17[795], line_16[793], line_15[791], line_14[789], line_13[787], line_12[785], line_11[783], line_10[781], line_9[779], line_8[777], line_7[775], line_6[773], line_5[771], line_4[769], line_3[767], line_2[765], line_1[763] };
assign col_1018 = {line_128[1018], line_127[1016], line_126[1014], line_125[1012], line_124[1010], line_123[1008], line_122[1006], line_121[1004], line_120[1002], line_119[1000], line_118[998], line_117[996], line_116[994], line_115[992], line_114[990], line_113[988], line_112[986], line_111[984], line_110[982], line_109[980], line_108[978], line_107[976], line_106[974], line_105[972], line_104[970], line_103[968], line_102[966], line_101[964], line_100[962], line_99[960], line_98[958], line_97[956], line_96[954], line_95[952], line_94[950], line_93[948], line_92[946], line_91[944], line_90[942], line_89[940], line_88[938], line_87[936], line_86[934], line_85[932], line_84[930], line_83[928], line_82[926], line_81[924], line_80[922], line_79[920], line_78[918], line_77[916], line_76[914], line_75[912], line_74[910], line_73[908], line_72[906], line_71[904], line_70[902], line_69[900], line_68[898], line_67[896], line_66[894], line_65[892], line_64[890], line_63[888], line_62[886], line_61[884], line_60[882], line_59[880], line_58[878], line_57[876], line_56[874], line_55[872], line_54[870], line_53[868], line_52[866], line_51[864], line_50[862], line_49[860], line_48[858], line_47[856], line_46[854], line_45[852], line_44[850], line_43[848], line_42[846], line_41[844], line_40[842], line_39[840], line_38[838], line_37[836], line_36[834], line_35[832], line_34[830], line_33[828], line_32[826], line_31[824], line_30[822], line_29[820], line_28[818], line_27[816], line_26[814], line_25[812], line_24[810], line_23[808], line_22[806], line_21[804], line_20[802], line_19[800], line_18[798], line_17[796], line_16[794], line_15[792], line_14[790], line_13[788], line_12[786], line_11[784], line_10[782], line_9[780], line_8[778], line_7[776], line_6[774], line_5[772], line_4[770], line_3[768], line_2[766], line_1[764] };
assign col_1019 = {line_128[1019], line_127[1017], line_126[1015], line_125[1013], line_124[1011], line_123[1009], line_122[1007], line_121[1005], line_120[1003], line_119[1001], line_118[999], line_117[997], line_116[995], line_115[993], line_114[991], line_113[989], line_112[987], line_111[985], line_110[983], line_109[981], line_108[979], line_107[977], line_106[975], line_105[973], line_104[971], line_103[969], line_102[967], line_101[965], line_100[963], line_99[961], line_98[959], line_97[957], line_96[955], line_95[953], line_94[951], line_93[949], line_92[947], line_91[945], line_90[943], line_89[941], line_88[939], line_87[937], line_86[935], line_85[933], line_84[931], line_83[929], line_82[927], line_81[925], line_80[923], line_79[921], line_78[919], line_77[917], line_76[915], line_75[913], line_74[911], line_73[909], line_72[907], line_71[905], line_70[903], line_69[901], line_68[899], line_67[897], line_66[895], line_65[893], line_64[891], line_63[889], line_62[887], line_61[885], line_60[883], line_59[881], line_58[879], line_57[877], line_56[875], line_55[873], line_54[871], line_53[869], line_52[867], line_51[865], line_50[863], line_49[861], line_48[859], line_47[857], line_46[855], line_45[853], line_44[851], line_43[849], line_42[847], line_41[845], line_40[843], line_39[841], line_38[839], line_37[837], line_36[835], line_35[833], line_34[831], line_33[829], line_32[827], line_31[825], line_30[823], line_29[821], line_28[819], line_27[817], line_26[815], line_25[813], line_24[811], line_23[809], line_22[807], line_21[805], line_20[803], line_19[801], line_18[799], line_17[797], line_16[795], line_15[793], line_14[791], line_13[789], line_12[787], line_11[785], line_10[783], line_9[781], line_8[779], line_7[777], line_6[775], line_5[773], line_4[771], line_3[769], line_2[767], line_1[765] };
assign col_1020 = {line_128[1020], line_127[1018], line_126[1016], line_125[1014], line_124[1012], line_123[1010], line_122[1008], line_121[1006], line_120[1004], line_119[1002], line_118[1000], line_117[998], line_116[996], line_115[994], line_114[992], line_113[990], line_112[988], line_111[986], line_110[984], line_109[982], line_108[980], line_107[978], line_106[976], line_105[974], line_104[972], line_103[970], line_102[968], line_101[966], line_100[964], line_99[962], line_98[960], line_97[958], line_96[956], line_95[954], line_94[952], line_93[950], line_92[948], line_91[946], line_90[944], line_89[942], line_88[940], line_87[938], line_86[936], line_85[934], line_84[932], line_83[930], line_82[928], line_81[926], line_80[924], line_79[922], line_78[920], line_77[918], line_76[916], line_75[914], line_74[912], line_73[910], line_72[908], line_71[906], line_70[904], line_69[902], line_68[900], line_67[898], line_66[896], line_65[894], line_64[892], line_63[890], line_62[888], line_61[886], line_60[884], line_59[882], line_58[880], line_57[878], line_56[876], line_55[874], line_54[872], line_53[870], line_52[868], line_51[866], line_50[864], line_49[862], line_48[860], line_47[858], line_46[856], line_45[854], line_44[852], line_43[850], line_42[848], line_41[846], line_40[844], line_39[842], line_38[840], line_37[838], line_36[836], line_35[834], line_34[832], line_33[830], line_32[828], line_31[826], line_30[824], line_29[822], line_28[820], line_27[818], line_26[816], line_25[814], line_24[812], line_23[810], line_22[808], line_21[806], line_20[804], line_19[802], line_18[800], line_17[798], line_16[796], line_15[794], line_14[792], line_13[790], line_12[788], line_11[786], line_10[784], line_9[782], line_8[780], line_7[778], line_6[776], line_5[774], line_4[772], line_3[770], line_2[768], line_1[766] };
assign col_1021 = {line_128[1021], line_127[1019], line_126[1017], line_125[1015], line_124[1013], line_123[1011], line_122[1009], line_121[1007], line_120[1005], line_119[1003], line_118[1001], line_117[999], line_116[997], line_115[995], line_114[993], line_113[991], line_112[989], line_111[987], line_110[985], line_109[983], line_108[981], line_107[979], line_106[977], line_105[975], line_104[973], line_103[971], line_102[969], line_101[967], line_100[965], line_99[963], line_98[961], line_97[959], line_96[957], line_95[955], line_94[953], line_93[951], line_92[949], line_91[947], line_90[945], line_89[943], line_88[941], line_87[939], line_86[937], line_85[935], line_84[933], line_83[931], line_82[929], line_81[927], line_80[925], line_79[923], line_78[921], line_77[919], line_76[917], line_75[915], line_74[913], line_73[911], line_72[909], line_71[907], line_70[905], line_69[903], line_68[901], line_67[899], line_66[897], line_65[895], line_64[893], line_63[891], line_62[889], line_61[887], line_60[885], line_59[883], line_58[881], line_57[879], line_56[877], line_55[875], line_54[873], line_53[871], line_52[869], line_51[867], line_50[865], line_49[863], line_48[861], line_47[859], line_46[857], line_45[855], line_44[853], line_43[851], line_42[849], line_41[847], line_40[845], line_39[843], line_38[841], line_37[839], line_36[837], line_35[835], line_34[833], line_33[831], line_32[829], line_31[827], line_30[825], line_29[823], line_28[821], line_27[819], line_26[817], line_25[815], line_24[813], line_23[811], line_22[809], line_21[807], line_20[805], line_19[803], line_18[801], line_17[799], line_16[797], line_15[795], line_14[793], line_13[791], line_12[789], line_11[787], line_10[785], line_9[783], line_8[781], line_7[779], line_6[777], line_5[775], line_4[773], line_3[771], line_2[769], line_1[767] };
assign col_1022 = {line_128[1022], line_127[1020], line_126[1018], line_125[1016], line_124[1014], line_123[1012], line_122[1010], line_121[1008], line_120[1006], line_119[1004], line_118[1002], line_117[1000], line_116[998], line_115[996], line_114[994], line_113[992], line_112[990], line_111[988], line_110[986], line_109[984], line_108[982], line_107[980], line_106[978], line_105[976], line_104[974], line_103[972], line_102[970], line_101[968], line_100[966], line_99[964], line_98[962], line_97[960], line_96[958], line_95[956], line_94[954], line_93[952], line_92[950], line_91[948], line_90[946], line_89[944], line_88[942], line_87[940], line_86[938], line_85[936], line_84[934], line_83[932], line_82[930], line_81[928], line_80[926], line_79[924], line_78[922], line_77[920], line_76[918], line_75[916], line_74[914], line_73[912], line_72[910], line_71[908], line_70[906], line_69[904], line_68[902], line_67[900], line_66[898], line_65[896], line_64[894], line_63[892], line_62[890], line_61[888], line_60[886], line_59[884], line_58[882], line_57[880], line_56[878], line_55[876], line_54[874], line_53[872], line_52[870], line_51[868], line_50[866], line_49[864], line_48[862], line_47[860], line_46[858], line_45[856], line_44[854], line_43[852], line_42[850], line_41[848], line_40[846], line_39[844], line_38[842], line_37[840], line_36[838], line_35[836], line_34[834], line_33[832], line_32[830], line_31[828], line_30[826], line_29[824], line_28[822], line_27[820], line_26[818], line_25[816], line_24[814], line_23[812], line_22[810], line_21[808], line_20[806], line_19[804], line_18[802], line_17[800], line_16[798], line_15[796], line_14[794], line_13[792], line_12[790], line_11[788], line_10[786], line_9[784], line_8[782], line_7[780], line_6[778], line_5[776], line_4[774], line_3[772], line_2[770], line_1[768] };
assign col_1023 = {line_128[1023], line_127[1021], line_126[1019], line_125[1017], line_124[1015], line_123[1013], line_122[1011], line_121[1009], line_120[1007], line_119[1005], line_118[1003], line_117[1001], line_116[999], line_115[997], line_114[995], line_113[993], line_112[991], line_111[989], line_110[987], line_109[985], line_108[983], line_107[981], line_106[979], line_105[977], line_104[975], line_103[973], line_102[971], line_101[969], line_100[967], line_99[965], line_98[963], line_97[961], line_96[959], line_95[957], line_94[955], line_93[953], line_92[951], line_91[949], line_90[947], line_89[945], line_88[943], line_87[941], line_86[939], line_85[937], line_84[935], line_83[933], line_82[931], line_81[929], line_80[927], line_79[925], line_78[923], line_77[921], line_76[919], line_75[917], line_74[915], line_73[913], line_72[911], line_71[909], line_70[907], line_69[905], line_68[903], line_67[901], line_66[899], line_65[897], line_64[895], line_63[893], line_62[891], line_61[889], line_60[887], line_59[885], line_58[883], line_57[881], line_56[879], line_55[877], line_54[875], line_53[873], line_52[871], line_51[869], line_50[867], line_49[865], line_48[863], line_47[861], line_46[859], line_45[857], line_44[855], line_43[853], line_42[851], line_41[849], line_40[847], line_39[845], line_38[843], line_37[841], line_36[839], line_35[837], line_34[835], line_33[833], line_32[831], line_31[829], line_30[827], line_29[825], line_28[823], line_27[821], line_26[819], line_25[817], line_24[815], line_23[813], line_22[811], line_21[809], line_20[807], line_19[805], line_18[803], line_17[801], line_16[799], line_15[797], line_14[795], line_13[793], line_12[791], line_11[789], line_10[787], line_9[785], line_8[783], line_7[781], line_6[779], line_5[777], line_4[775], line_3[773], line_2[771], line_1[769] };
assign col_1024 = {line_128[1024], line_127[1022], line_126[1020], line_125[1018], line_124[1016], line_123[1014], line_122[1012], line_121[1010], line_120[1008], line_119[1006], line_118[1004], line_117[1002], line_116[1000], line_115[998], line_114[996], line_113[994], line_112[992], line_111[990], line_110[988], line_109[986], line_108[984], line_107[982], line_106[980], line_105[978], line_104[976], line_103[974], line_102[972], line_101[970], line_100[968], line_99[966], line_98[964], line_97[962], line_96[960], line_95[958], line_94[956], line_93[954], line_92[952], line_91[950], line_90[948], line_89[946], line_88[944], line_87[942], line_86[940], line_85[938], line_84[936], line_83[934], line_82[932], line_81[930], line_80[928], line_79[926], line_78[924], line_77[922], line_76[920], line_75[918], line_74[916], line_73[914], line_72[912], line_71[910], line_70[908], line_69[906], line_68[904], line_67[902], line_66[900], line_65[898], line_64[896], line_63[894], line_62[892], line_61[890], line_60[888], line_59[886], line_58[884], line_57[882], line_56[880], line_55[878], line_54[876], line_53[874], line_52[872], line_51[870], line_50[868], line_49[866], line_48[864], line_47[862], line_46[860], line_45[858], line_44[856], line_43[854], line_42[852], line_41[850], line_40[848], line_39[846], line_38[844], line_37[842], line_36[840], line_35[838], line_34[836], line_33[834], line_32[832], line_31[830], line_30[828], line_29[826], line_28[824], line_27[822], line_26[820], line_25[818], line_24[816], line_23[814], line_22[812], line_21[810], line_20[808], line_19[806], line_18[804], line_17[802], line_16[800], line_15[798], line_14[796], line_13[794], line_12[792], line_11[790], line_10[788], line_9[786], line_8[784], line_7[782], line_6[780], line_5[778], line_4[776], line_3[774], line_2[772], line_1[770] };
assign col_1025 = {line_128[1025], line_127[1023], line_126[1021], line_125[1019], line_124[1017], line_123[1015], line_122[1013], line_121[1011], line_120[1009], line_119[1007], line_118[1005], line_117[1003], line_116[1001], line_115[999], line_114[997], line_113[995], line_112[993], line_111[991], line_110[989], line_109[987], line_108[985], line_107[983], line_106[981], line_105[979], line_104[977], line_103[975], line_102[973], line_101[971], line_100[969], line_99[967], line_98[965], line_97[963], line_96[961], line_95[959], line_94[957], line_93[955], line_92[953], line_91[951], line_90[949], line_89[947], line_88[945], line_87[943], line_86[941], line_85[939], line_84[937], line_83[935], line_82[933], line_81[931], line_80[929], line_79[927], line_78[925], line_77[923], line_76[921], line_75[919], line_74[917], line_73[915], line_72[913], line_71[911], line_70[909], line_69[907], line_68[905], line_67[903], line_66[901], line_65[899], line_64[897], line_63[895], line_62[893], line_61[891], line_60[889], line_59[887], line_58[885], line_57[883], line_56[881], line_55[879], line_54[877], line_53[875], line_52[873], line_51[871], line_50[869], line_49[867], line_48[865], line_47[863], line_46[861], line_45[859], line_44[857], line_43[855], line_42[853], line_41[851], line_40[849], line_39[847], line_38[845], line_37[843], line_36[841], line_35[839], line_34[837], line_33[835], line_32[833], line_31[831], line_30[829], line_29[827], line_28[825], line_27[823], line_26[821], line_25[819], line_24[817], line_23[815], line_22[813], line_21[811], line_20[809], line_19[807], line_18[805], line_17[803], line_16[801], line_15[799], line_14[797], line_13[795], line_12[793], line_11[791], line_10[789], line_9[787], line_8[785], line_7[783], line_6[781], line_5[779], line_4[777], line_3[775], line_2[773], line_1[771] };

assign col_1026 = {line_127[1024], line_126[1022], line_125[1020], line_124[1018], line_123[1016], line_122[1014], line_121[1012], line_120[1010], line_119[1008], line_118[1006], line_117[1004], line_116[1002], line_115[1000], line_114[998], line_113[996], line_112[994], line_111[992], line_110[990], line_109[988], line_108[986], line_107[984], line_106[982], line_105[980], line_104[978], line_103[976], line_102[974], line_101[972], line_100[970], line_99[968], line_98[966], line_97[964], line_96[962], line_95[960], line_94[958], line_93[956], line_92[954], line_91[952], line_90[950], line_89[948], line_88[946], line_87[944], line_86[942], line_85[940], line_84[938], line_83[936], line_82[934], line_81[932], line_80[930], line_79[928], line_78[926], line_77[924], line_76[922], line_75[920], line_74[918], line_73[916], line_72[914], line_71[912], line_70[910], line_69[908], line_68[906], line_67[904], line_66[902], line_65[900], line_64[898], line_63[896], line_62[894], line_61[892], line_60[890], line_59[888], line_58[886], line_57[884], line_56[882], line_55[880], line_54[878], line_53[876], line_52[874], line_51[872], line_50[870], line_49[868], line_48[866], line_47[864], line_46[862], line_45[860], line_44[858], line_43[856], line_42[854], line_41[852], line_40[850], line_39[848], line_38[846], line_37[844], line_36[842], line_35[840], line_34[838], line_33[836], line_32[834], line_31[832], line_30[830], line_29[828], line_28[826], line_27[824], line_26[822], line_25[820], line_24[818], line_23[816], line_22[814], line_21[812], line_20[810], line_19[808], line_18[806], line_17[804], line_16[802], line_15[800], line_14[798], line_13[796], line_12[794], line_11[792], line_10[790], line_9[788], line_8[786], line_7[784], line_6[782], line_5[780], line_4[778], line_3[776], line_2[774], line_1[772], 1'b0};
assign col_1027 = {line_127[1025], line_126[1023], line_125[1021], line_124[1019], line_123[1017], line_122[1015], line_121[1013], line_120[1011], line_119[1009], line_118[1007], line_117[1005], line_116[1003], line_115[1001], line_114[999], line_113[997], line_112[995], line_111[993], line_110[991], line_109[989], line_108[987], line_107[985], line_106[983], line_105[981], line_104[979], line_103[977], line_102[975], line_101[973], line_100[971], line_99[969], line_98[967], line_97[965], line_96[963], line_95[961], line_94[959], line_93[957], line_92[955], line_91[953], line_90[951], line_89[949], line_88[947], line_87[945], line_86[943], line_85[941], line_84[939], line_83[937], line_82[935], line_81[933], line_80[931], line_79[929], line_78[927], line_77[925], line_76[923], line_75[921], line_74[919], line_73[917], line_72[915], line_71[913], line_70[911], line_69[909], line_68[907], line_67[905], line_66[903], line_65[901], line_64[899], line_63[897], line_62[895], line_61[893], line_60[891], line_59[889], line_58[887], line_57[885], line_56[883], line_55[881], line_54[879], line_53[877], line_52[875], line_51[873], line_50[871], line_49[869], line_48[867], line_47[865], line_46[863], line_45[861], line_44[859], line_43[857], line_42[855], line_41[853], line_40[851], line_39[849], line_38[847], line_37[845], line_36[843], line_35[841], line_34[839], line_33[837], line_32[835], line_31[833], line_30[831], line_29[829], line_28[827], line_27[825], line_26[823], line_25[821], line_24[819], line_23[817], line_22[815], line_21[813], line_20[811], line_19[809], line_18[807], line_17[805], line_16[803], line_15[801], line_14[799], line_13[797], line_12[795], line_11[793], line_10[791], line_9[789], line_8[787], line_7[785], line_6[783], line_5[781], line_4[779], line_3[777], line_2[775], line_1[773], 1'b0};
assign col_1028 = {line_126[1024], line_125[1022], line_124[1020], line_123[1018], line_122[1016], line_121[1014], line_120[1012], line_119[1010], line_118[1008], line_117[1006], line_116[1004], line_115[1002], line_114[1000], line_113[998], line_112[996], line_111[994], line_110[992], line_109[990], line_108[988], line_107[986], line_106[984], line_105[982], line_104[980], line_103[978], line_102[976], line_101[974], line_100[972], line_99[970], line_98[968], line_97[966], line_96[964], line_95[962], line_94[960], line_93[958], line_92[956], line_91[954], line_90[952], line_89[950], line_88[948], line_87[946], line_86[944], line_85[942], line_84[940], line_83[938], line_82[936], line_81[934], line_80[932], line_79[930], line_78[928], line_77[926], line_76[924], line_75[922], line_74[920], line_73[918], line_72[916], line_71[914], line_70[912], line_69[910], line_68[908], line_67[906], line_66[904], line_65[902], line_64[900], line_63[898], line_62[896], line_61[894], line_60[892], line_59[890], line_58[888], line_57[886], line_56[884], line_55[882], line_54[880], line_53[878], line_52[876], line_51[874], line_50[872], line_49[870], line_48[868], line_47[866], line_46[864], line_45[862], line_44[860], line_43[858], line_42[856], line_41[854], line_40[852], line_39[850], line_38[848], line_37[846], line_36[844], line_35[842], line_34[840], line_33[838], line_32[836], line_31[834], line_30[832], line_29[830], line_28[828], line_27[826], line_26[824], line_25[822], line_24[820], line_23[818], line_22[816], line_21[814], line_20[812], line_19[810], line_18[808], line_17[806], line_16[804], line_15[802], line_14[800], line_13[798], line_12[796], line_11[794], line_10[792], line_9[790], line_8[788], line_7[786], line_6[784], line_5[782], line_4[780], line_3[778], line_2[776], line_1[774], 2'b0};
assign col_1029 = {line_126[1025], line_125[1023], line_124[1021], line_123[1019], line_122[1017], line_121[1015], line_120[1013], line_119[1011], line_118[1009], line_117[1007], line_116[1005], line_115[1003], line_114[1001], line_113[999], line_112[997], line_111[995], line_110[993], line_109[991], line_108[989], line_107[987], line_106[985], line_105[983], line_104[981], line_103[979], line_102[977], line_101[975], line_100[973], line_99[971], line_98[969], line_97[967], line_96[965], line_95[963], line_94[961], line_93[959], line_92[957], line_91[955], line_90[953], line_89[951], line_88[949], line_87[947], line_86[945], line_85[943], line_84[941], line_83[939], line_82[937], line_81[935], line_80[933], line_79[931], line_78[929], line_77[927], line_76[925], line_75[923], line_74[921], line_73[919], line_72[917], line_71[915], line_70[913], line_69[911], line_68[909], line_67[907], line_66[905], line_65[903], line_64[901], line_63[899], line_62[897], line_61[895], line_60[893], line_59[891], line_58[889], line_57[887], line_56[885], line_55[883], line_54[881], line_53[879], line_52[877], line_51[875], line_50[873], line_49[871], line_48[869], line_47[867], line_46[865], line_45[863], line_44[861], line_43[859], line_42[857], line_41[855], line_40[853], line_39[851], line_38[849], line_37[847], line_36[845], line_35[843], line_34[841], line_33[839], line_32[837], line_31[835], line_30[833], line_29[831], line_28[829], line_27[827], line_26[825], line_25[823], line_24[821], line_23[819], line_22[817], line_21[815], line_20[813], line_19[811], line_18[809], line_17[807], line_16[805], line_15[803], line_14[801], line_13[799], line_12[797], line_11[795], line_10[793], line_9[791], line_8[789], line_7[787], line_6[785], line_5[783], line_4[781], line_3[779], line_2[777], line_1[775], 2'b0};
assign col_1030 = {line_125[1024], line_124[1022], line_123[1020], line_122[1018], line_121[1016], line_120[1014], line_119[1012], line_118[1010], line_117[1008], line_116[1006], line_115[1004], line_114[1002], line_113[1000], line_112[998], line_111[996], line_110[994], line_109[992], line_108[990], line_107[988], line_106[986], line_105[984], line_104[982], line_103[980], line_102[978], line_101[976], line_100[974], line_99[972], line_98[970], line_97[968], line_96[966], line_95[964], line_94[962], line_93[960], line_92[958], line_91[956], line_90[954], line_89[952], line_88[950], line_87[948], line_86[946], line_85[944], line_84[942], line_83[940], line_82[938], line_81[936], line_80[934], line_79[932], line_78[930], line_77[928], line_76[926], line_75[924], line_74[922], line_73[920], line_72[918], line_71[916], line_70[914], line_69[912], line_68[910], line_67[908], line_66[906], line_65[904], line_64[902], line_63[900], line_62[898], line_61[896], line_60[894], line_59[892], line_58[890], line_57[888], line_56[886], line_55[884], line_54[882], line_53[880], line_52[878], line_51[876], line_50[874], line_49[872], line_48[870], line_47[868], line_46[866], line_45[864], line_44[862], line_43[860], line_42[858], line_41[856], line_40[854], line_39[852], line_38[850], line_37[848], line_36[846], line_35[844], line_34[842], line_33[840], line_32[838], line_31[836], line_30[834], line_29[832], line_28[830], line_27[828], line_26[826], line_25[824], line_24[822], line_23[820], line_22[818], line_21[816], line_20[814], line_19[812], line_18[810], line_17[808], line_16[806], line_15[804], line_14[802], line_13[800], line_12[798], line_11[796], line_10[794], line_9[792], line_8[790], line_7[788], line_6[786], line_5[784], line_4[782], line_3[780], line_2[778], line_1[776], 3'b0};
assign col_1031 = {line_125[1025], line_124[1023], line_123[1021], line_122[1019], line_121[1017], line_120[1015], line_119[1013], line_118[1011], line_117[1009], line_116[1007], line_115[1005], line_114[1003], line_113[1001], line_112[999], line_111[997], line_110[995], line_109[993], line_108[991], line_107[989], line_106[987], line_105[985], line_104[983], line_103[981], line_102[979], line_101[977], line_100[975], line_99[973], line_98[971], line_97[969], line_96[967], line_95[965], line_94[963], line_93[961], line_92[959], line_91[957], line_90[955], line_89[953], line_88[951], line_87[949], line_86[947], line_85[945], line_84[943], line_83[941], line_82[939], line_81[937], line_80[935], line_79[933], line_78[931], line_77[929], line_76[927], line_75[925], line_74[923], line_73[921], line_72[919], line_71[917], line_70[915], line_69[913], line_68[911], line_67[909], line_66[907], line_65[905], line_64[903], line_63[901], line_62[899], line_61[897], line_60[895], line_59[893], line_58[891], line_57[889], line_56[887], line_55[885], line_54[883], line_53[881], line_52[879], line_51[877], line_50[875], line_49[873], line_48[871], line_47[869], line_46[867], line_45[865], line_44[863], line_43[861], line_42[859], line_41[857], line_40[855], line_39[853], line_38[851], line_37[849], line_36[847], line_35[845], line_34[843], line_33[841], line_32[839], line_31[837], line_30[835], line_29[833], line_28[831], line_27[829], line_26[827], line_25[825], line_24[823], line_23[821], line_22[819], line_21[817], line_20[815], line_19[813], line_18[811], line_17[809], line_16[807], line_15[805], line_14[803], line_13[801], line_12[799], line_11[797], line_10[795], line_9[793], line_8[791], line_7[789], line_6[787], line_5[785], line_4[783], line_3[781], line_2[779], line_1[777], 3'b0};
assign col_1032 = {line_124[1024], line_123[1022], line_122[1020], line_121[1018], line_120[1016], line_119[1014], line_118[1012], line_117[1010], line_116[1008], line_115[1006], line_114[1004], line_113[1002], line_112[1000], line_111[998], line_110[996], line_109[994], line_108[992], line_107[990], line_106[988], line_105[986], line_104[984], line_103[982], line_102[980], line_101[978], line_100[976], line_99[974], line_98[972], line_97[970], line_96[968], line_95[966], line_94[964], line_93[962], line_92[960], line_91[958], line_90[956], line_89[954], line_88[952], line_87[950], line_86[948], line_85[946], line_84[944], line_83[942], line_82[940], line_81[938], line_80[936], line_79[934], line_78[932], line_77[930], line_76[928], line_75[926], line_74[924], line_73[922], line_72[920], line_71[918], line_70[916], line_69[914], line_68[912], line_67[910], line_66[908], line_65[906], line_64[904], line_63[902], line_62[900], line_61[898], line_60[896], line_59[894], line_58[892], line_57[890], line_56[888], line_55[886], line_54[884], line_53[882], line_52[880], line_51[878], line_50[876], line_49[874], line_48[872], line_47[870], line_46[868], line_45[866], line_44[864], line_43[862], line_42[860], line_41[858], line_40[856], line_39[854], line_38[852], line_37[850], line_36[848], line_35[846], line_34[844], line_33[842], line_32[840], line_31[838], line_30[836], line_29[834], line_28[832], line_27[830], line_26[828], line_25[826], line_24[824], line_23[822], line_22[820], line_21[818], line_20[816], line_19[814], line_18[812], line_17[810], line_16[808], line_15[806], line_14[804], line_13[802], line_12[800], line_11[798], line_10[796], line_9[794], line_8[792], line_7[790], line_6[788], line_5[786], line_4[784], line_3[782], line_2[780], line_1[778], 4'b0};
assign col_1033 = {line_124[1025], line_123[1023], line_122[1021], line_121[1019], line_120[1017], line_119[1015], line_118[1013], line_117[1011], line_116[1009], line_115[1007], line_114[1005], line_113[1003], line_112[1001], line_111[999], line_110[997], line_109[995], line_108[993], line_107[991], line_106[989], line_105[987], line_104[985], line_103[983], line_102[981], line_101[979], line_100[977], line_99[975], line_98[973], line_97[971], line_96[969], line_95[967], line_94[965], line_93[963], line_92[961], line_91[959], line_90[957], line_89[955], line_88[953], line_87[951], line_86[949], line_85[947], line_84[945], line_83[943], line_82[941], line_81[939], line_80[937], line_79[935], line_78[933], line_77[931], line_76[929], line_75[927], line_74[925], line_73[923], line_72[921], line_71[919], line_70[917], line_69[915], line_68[913], line_67[911], line_66[909], line_65[907], line_64[905], line_63[903], line_62[901], line_61[899], line_60[897], line_59[895], line_58[893], line_57[891], line_56[889], line_55[887], line_54[885], line_53[883], line_52[881], line_51[879], line_50[877], line_49[875], line_48[873], line_47[871], line_46[869], line_45[867], line_44[865], line_43[863], line_42[861], line_41[859], line_40[857], line_39[855], line_38[853], line_37[851], line_36[849], line_35[847], line_34[845], line_33[843], line_32[841], line_31[839], line_30[837], line_29[835], line_28[833], line_27[831], line_26[829], line_25[827], line_24[825], line_23[823], line_22[821], line_21[819], line_20[817], line_19[815], line_18[813], line_17[811], line_16[809], line_15[807], line_14[805], line_13[803], line_12[801], line_11[799], line_10[797], line_9[795], line_8[793], line_7[791], line_6[789], line_5[787], line_4[785], line_3[783], line_2[781], line_1[779], 4'b0};
assign col_1034 = {line_123[1024], line_122[1022], line_121[1020], line_120[1018], line_119[1016], line_118[1014], line_117[1012], line_116[1010], line_115[1008], line_114[1006], line_113[1004], line_112[1002], line_111[1000], line_110[998], line_109[996], line_108[994], line_107[992], line_106[990], line_105[988], line_104[986], line_103[984], line_102[982], line_101[980], line_100[978], line_99[976], line_98[974], line_97[972], line_96[970], line_95[968], line_94[966], line_93[964], line_92[962], line_91[960], line_90[958], line_89[956], line_88[954], line_87[952], line_86[950], line_85[948], line_84[946], line_83[944], line_82[942], line_81[940], line_80[938], line_79[936], line_78[934], line_77[932], line_76[930], line_75[928], line_74[926], line_73[924], line_72[922], line_71[920], line_70[918], line_69[916], line_68[914], line_67[912], line_66[910], line_65[908], line_64[906], line_63[904], line_62[902], line_61[900], line_60[898], line_59[896], line_58[894], line_57[892], line_56[890], line_55[888], line_54[886], line_53[884], line_52[882], line_51[880], line_50[878], line_49[876], line_48[874], line_47[872], line_46[870], line_45[868], line_44[866], line_43[864], line_42[862], line_41[860], line_40[858], line_39[856], line_38[854], line_37[852], line_36[850], line_35[848], line_34[846], line_33[844], line_32[842], line_31[840], line_30[838], line_29[836], line_28[834], line_27[832], line_26[830], line_25[828], line_24[826], line_23[824], line_22[822], line_21[820], line_20[818], line_19[816], line_18[814], line_17[812], line_16[810], line_15[808], line_14[806], line_13[804], line_12[802], line_11[800], line_10[798], line_9[796], line_8[794], line_7[792], line_6[790], line_5[788], line_4[786], line_3[784], line_2[782], line_1[780], 5'b0};
assign col_1035 = {line_123[1025], line_122[1023], line_121[1021], line_120[1019], line_119[1017], line_118[1015], line_117[1013], line_116[1011], line_115[1009], line_114[1007], line_113[1005], line_112[1003], line_111[1001], line_110[999], line_109[997], line_108[995], line_107[993], line_106[991], line_105[989], line_104[987], line_103[985], line_102[983], line_101[981], line_100[979], line_99[977], line_98[975], line_97[973], line_96[971], line_95[969], line_94[967], line_93[965], line_92[963], line_91[961], line_90[959], line_89[957], line_88[955], line_87[953], line_86[951], line_85[949], line_84[947], line_83[945], line_82[943], line_81[941], line_80[939], line_79[937], line_78[935], line_77[933], line_76[931], line_75[929], line_74[927], line_73[925], line_72[923], line_71[921], line_70[919], line_69[917], line_68[915], line_67[913], line_66[911], line_65[909], line_64[907], line_63[905], line_62[903], line_61[901], line_60[899], line_59[897], line_58[895], line_57[893], line_56[891], line_55[889], line_54[887], line_53[885], line_52[883], line_51[881], line_50[879], line_49[877], line_48[875], line_47[873], line_46[871], line_45[869], line_44[867], line_43[865], line_42[863], line_41[861], line_40[859], line_39[857], line_38[855], line_37[853], line_36[851], line_35[849], line_34[847], line_33[845], line_32[843], line_31[841], line_30[839], line_29[837], line_28[835], line_27[833], line_26[831], line_25[829], line_24[827], line_23[825], line_22[823], line_21[821], line_20[819], line_19[817], line_18[815], line_17[813], line_16[811], line_15[809], line_14[807], line_13[805], line_12[803], line_11[801], line_10[799], line_9[797], line_8[795], line_7[793], line_6[791], line_5[789], line_4[787], line_3[785], line_2[783], line_1[781], 5'b0};
assign col_1036 = {line_122[1024], line_121[1022], line_120[1020], line_119[1018], line_118[1016], line_117[1014], line_116[1012], line_115[1010], line_114[1008], line_113[1006], line_112[1004], line_111[1002], line_110[1000], line_109[998], line_108[996], line_107[994], line_106[992], line_105[990], line_104[988], line_103[986], line_102[984], line_101[982], line_100[980], line_99[978], line_98[976], line_97[974], line_96[972], line_95[970], line_94[968], line_93[966], line_92[964], line_91[962], line_90[960], line_89[958], line_88[956], line_87[954], line_86[952], line_85[950], line_84[948], line_83[946], line_82[944], line_81[942], line_80[940], line_79[938], line_78[936], line_77[934], line_76[932], line_75[930], line_74[928], line_73[926], line_72[924], line_71[922], line_70[920], line_69[918], line_68[916], line_67[914], line_66[912], line_65[910], line_64[908], line_63[906], line_62[904], line_61[902], line_60[900], line_59[898], line_58[896], line_57[894], line_56[892], line_55[890], line_54[888], line_53[886], line_52[884], line_51[882], line_50[880], line_49[878], line_48[876], line_47[874], line_46[872], line_45[870], line_44[868], line_43[866], line_42[864], line_41[862], line_40[860], line_39[858], line_38[856], line_37[854], line_36[852], line_35[850], line_34[848], line_33[846], line_32[844], line_31[842], line_30[840], line_29[838], line_28[836], line_27[834], line_26[832], line_25[830], line_24[828], line_23[826], line_22[824], line_21[822], line_20[820], line_19[818], line_18[816], line_17[814], line_16[812], line_15[810], line_14[808], line_13[806], line_12[804], line_11[802], line_10[800], line_9[798], line_8[796], line_7[794], line_6[792], line_5[790], line_4[788], line_3[786], line_2[784], line_1[782], 6'b0};
assign col_1037 = {line_122[1025], line_121[1023], line_120[1021], line_119[1019], line_118[1017], line_117[1015], line_116[1013], line_115[1011], line_114[1009], line_113[1007], line_112[1005], line_111[1003], line_110[1001], line_109[999], line_108[997], line_107[995], line_106[993], line_105[991], line_104[989], line_103[987], line_102[985], line_101[983], line_100[981], line_99[979], line_98[977], line_97[975], line_96[973], line_95[971], line_94[969], line_93[967], line_92[965], line_91[963], line_90[961], line_89[959], line_88[957], line_87[955], line_86[953], line_85[951], line_84[949], line_83[947], line_82[945], line_81[943], line_80[941], line_79[939], line_78[937], line_77[935], line_76[933], line_75[931], line_74[929], line_73[927], line_72[925], line_71[923], line_70[921], line_69[919], line_68[917], line_67[915], line_66[913], line_65[911], line_64[909], line_63[907], line_62[905], line_61[903], line_60[901], line_59[899], line_58[897], line_57[895], line_56[893], line_55[891], line_54[889], line_53[887], line_52[885], line_51[883], line_50[881], line_49[879], line_48[877], line_47[875], line_46[873], line_45[871], line_44[869], line_43[867], line_42[865], line_41[863], line_40[861], line_39[859], line_38[857], line_37[855], line_36[853], line_35[851], line_34[849], line_33[847], line_32[845], line_31[843], line_30[841], line_29[839], line_28[837], line_27[835], line_26[833], line_25[831], line_24[829], line_23[827], line_22[825], line_21[823], line_20[821], line_19[819], line_18[817], line_17[815], line_16[813], line_15[811], line_14[809], line_13[807], line_12[805], line_11[803], line_10[801], line_9[799], line_8[797], line_7[795], line_6[793], line_5[791], line_4[789], line_3[787], line_2[785], line_1[783], 6'b0};
assign col_1038 = {line_121[1024], line_120[1022], line_119[1020], line_118[1018], line_117[1016], line_116[1014], line_115[1012], line_114[1010], line_113[1008], line_112[1006], line_111[1004], line_110[1002], line_109[1000], line_108[998], line_107[996], line_106[994], line_105[992], line_104[990], line_103[988], line_102[986], line_101[984], line_100[982], line_99[980], line_98[978], line_97[976], line_96[974], line_95[972], line_94[970], line_93[968], line_92[966], line_91[964], line_90[962], line_89[960], line_88[958], line_87[956], line_86[954], line_85[952], line_84[950], line_83[948], line_82[946], line_81[944], line_80[942], line_79[940], line_78[938], line_77[936], line_76[934], line_75[932], line_74[930], line_73[928], line_72[926], line_71[924], line_70[922], line_69[920], line_68[918], line_67[916], line_66[914], line_65[912], line_64[910], line_63[908], line_62[906], line_61[904], line_60[902], line_59[900], line_58[898], line_57[896], line_56[894], line_55[892], line_54[890], line_53[888], line_52[886], line_51[884], line_50[882], line_49[880], line_48[878], line_47[876], line_46[874], line_45[872], line_44[870], line_43[868], line_42[866], line_41[864], line_40[862], line_39[860], line_38[858], line_37[856], line_36[854], line_35[852], line_34[850], line_33[848], line_32[846], line_31[844], line_30[842], line_29[840], line_28[838], line_27[836], line_26[834], line_25[832], line_24[830], line_23[828], line_22[826], line_21[824], line_20[822], line_19[820], line_18[818], line_17[816], line_16[814], line_15[812], line_14[810], line_13[808], line_12[806], line_11[804], line_10[802], line_9[800], line_8[798], line_7[796], line_6[794], line_5[792], line_4[790], line_3[788], line_2[786], line_1[784], 7'b0};
assign col_1039 = {line_121[1025], line_120[1023], line_119[1021], line_118[1019], line_117[1017], line_116[1015], line_115[1013], line_114[1011], line_113[1009], line_112[1007], line_111[1005], line_110[1003], line_109[1001], line_108[999], line_107[997], line_106[995], line_105[993], line_104[991], line_103[989], line_102[987], line_101[985], line_100[983], line_99[981], line_98[979], line_97[977], line_96[975], line_95[973], line_94[971], line_93[969], line_92[967], line_91[965], line_90[963], line_89[961], line_88[959], line_87[957], line_86[955], line_85[953], line_84[951], line_83[949], line_82[947], line_81[945], line_80[943], line_79[941], line_78[939], line_77[937], line_76[935], line_75[933], line_74[931], line_73[929], line_72[927], line_71[925], line_70[923], line_69[921], line_68[919], line_67[917], line_66[915], line_65[913], line_64[911], line_63[909], line_62[907], line_61[905], line_60[903], line_59[901], line_58[899], line_57[897], line_56[895], line_55[893], line_54[891], line_53[889], line_52[887], line_51[885], line_50[883], line_49[881], line_48[879], line_47[877], line_46[875], line_45[873], line_44[871], line_43[869], line_42[867], line_41[865], line_40[863], line_39[861], line_38[859], line_37[857], line_36[855], line_35[853], line_34[851], line_33[849], line_32[847], line_31[845], line_30[843], line_29[841], line_28[839], line_27[837], line_26[835], line_25[833], line_24[831], line_23[829], line_22[827], line_21[825], line_20[823], line_19[821], line_18[819], line_17[817], line_16[815], line_15[813], line_14[811], line_13[809], line_12[807], line_11[805], line_10[803], line_9[801], line_8[799], line_7[797], line_6[795], line_5[793], line_4[791], line_3[789], line_2[787], line_1[785], 7'b0};
assign col_1040 = {line_120[1024], line_119[1022], line_118[1020], line_117[1018], line_116[1016], line_115[1014], line_114[1012], line_113[1010], line_112[1008], line_111[1006], line_110[1004], line_109[1002], line_108[1000], line_107[998], line_106[996], line_105[994], line_104[992], line_103[990], line_102[988], line_101[986], line_100[984], line_99[982], line_98[980], line_97[978], line_96[976], line_95[974], line_94[972], line_93[970], line_92[968], line_91[966], line_90[964], line_89[962], line_88[960], line_87[958], line_86[956], line_85[954], line_84[952], line_83[950], line_82[948], line_81[946], line_80[944], line_79[942], line_78[940], line_77[938], line_76[936], line_75[934], line_74[932], line_73[930], line_72[928], line_71[926], line_70[924], line_69[922], line_68[920], line_67[918], line_66[916], line_65[914], line_64[912], line_63[910], line_62[908], line_61[906], line_60[904], line_59[902], line_58[900], line_57[898], line_56[896], line_55[894], line_54[892], line_53[890], line_52[888], line_51[886], line_50[884], line_49[882], line_48[880], line_47[878], line_46[876], line_45[874], line_44[872], line_43[870], line_42[868], line_41[866], line_40[864], line_39[862], line_38[860], line_37[858], line_36[856], line_35[854], line_34[852], line_33[850], line_32[848], line_31[846], line_30[844], line_29[842], line_28[840], line_27[838], line_26[836], line_25[834], line_24[832], line_23[830], line_22[828], line_21[826], line_20[824], line_19[822], line_18[820], line_17[818], line_16[816], line_15[814], line_14[812], line_13[810], line_12[808], line_11[806], line_10[804], line_9[802], line_8[800], line_7[798], line_6[796], line_5[794], line_4[792], line_3[790], line_2[788], line_1[786], 8'b0};
assign col_1041 = {line_120[1025], line_119[1023], line_118[1021], line_117[1019], line_116[1017], line_115[1015], line_114[1013], line_113[1011], line_112[1009], line_111[1007], line_110[1005], line_109[1003], line_108[1001], line_107[999], line_106[997], line_105[995], line_104[993], line_103[991], line_102[989], line_101[987], line_100[985], line_99[983], line_98[981], line_97[979], line_96[977], line_95[975], line_94[973], line_93[971], line_92[969], line_91[967], line_90[965], line_89[963], line_88[961], line_87[959], line_86[957], line_85[955], line_84[953], line_83[951], line_82[949], line_81[947], line_80[945], line_79[943], line_78[941], line_77[939], line_76[937], line_75[935], line_74[933], line_73[931], line_72[929], line_71[927], line_70[925], line_69[923], line_68[921], line_67[919], line_66[917], line_65[915], line_64[913], line_63[911], line_62[909], line_61[907], line_60[905], line_59[903], line_58[901], line_57[899], line_56[897], line_55[895], line_54[893], line_53[891], line_52[889], line_51[887], line_50[885], line_49[883], line_48[881], line_47[879], line_46[877], line_45[875], line_44[873], line_43[871], line_42[869], line_41[867], line_40[865], line_39[863], line_38[861], line_37[859], line_36[857], line_35[855], line_34[853], line_33[851], line_32[849], line_31[847], line_30[845], line_29[843], line_28[841], line_27[839], line_26[837], line_25[835], line_24[833], line_23[831], line_22[829], line_21[827], line_20[825], line_19[823], line_18[821], line_17[819], line_16[817], line_15[815], line_14[813], line_13[811], line_12[809], line_11[807], line_10[805], line_9[803], line_8[801], line_7[799], line_6[797], line_5[795], line_4[793], line_3[791], line_2[789], line_1[787], 8'b0};
assign col_1042 = {line_119[1024], line_118[1022], line_117[1020], line_116[1018], line_115[1016], line_114[1014], line_113[1012], line_112[1010], line_111[1008], line_110[1006], line_109[1004], line_108[1002], line_107[1000], line_106[998], line_105[996], line_104[994], line_103[992], line_102[990], line_101[988], line_100[986], line_99[984], line_98[982], line_97[980], line_96[978], line_95[976], line_94[974], line_93[972], line_92[970], line_91[968], line_90[966], line_89[964], line_88[962], line_87[960], line_86[958], line_85[956], line_84[954], line_83[952], line_82[950], line_81[948], line_80[946], line_79[944], line_78[942], line_77[940], line_76[938], line_75[936], line_74[934], line_73[932], line_72[930], line_71[928], line_70[926], line_69[924], line_68[922], line_67[920], line_66[918], line_65[916], line_64[914], line_63[912], line_62[910], line_61[908], line_60[906], line_59[904], line_58[902], line_57[900], line_56[898], line_55[896], line_54[894], line_53[892], line_52[890], line_51[888], line_50[886], line_49[884], line_48[882], line_47[880], line_46[878], line_45[876], line_44[874], line_43[872], line_42[870], line_41[868], line_40[866], line_39[864], line_38[862], line_37[860], line_36[858], line_35[856], line_34[854], line_33[852], line_32[850], line_31[848], line_30[846], line_29[844], line_28[842], line_27[840], line_26[838], line_25[836], line_24[834], line_23[832], line_22[830], line_21[828], line_20[826], line_19[824], line_18[822], line_17[820], line_16[818], line_15[816], line_14[814], line_13[812], line_12[810], line_11[808], line_10[806], line_9[804], line_8[802], line_7[800], line_6[798], line_5[796], line_4[794], line_3[792], line_2[790], line_1[788], 9'b0};
assign col_1043 = {line_119[1025], line_118[1023], line_117[1021], line_116[1019], line_115[1017], line_114[1015], line_113[1013], line_112[1011], line_111[1009], line_110[1007], line_109[1005], line_108[1003], line_107[1001], line_106[999], line_105[997], line_104[995], line_103[993], line_102[991], line_101[989], line_100[987], line_99[985], line_98[983], line_97[981], line_96[979], line_95[977], line_94[975], line_93[973], line_92[971], line_91[969], line_90[967], line_89[965], line_88[963], line_87[961], line_86[959], line_85[957], line_84[955], line_83[953], line_82[951], line_81[949], line_80[947], line_79[945], line_78[943], line_77[941], line_76[939], line_75[937], line_74[935], line_73[933], line_72[931], line_71[929], line_70[927], line_69[925], line_68[923], line_67[921], line_66[919], line_65[917], line_64[915], line_63[913], line_62[911], line_61[909], line_60[907], line_59[905], line_58[903], line_57[901], line_56[899], line_55[897], line_54[895], line_53[893], line_52[891], line_51[889], line_50[887], line_49[885], line_48[883], line_47[881], line_46[879], line_45[877], line_44[875], line_43[873], line_42[871], line_41[869], line_40[867], line_39[865], line_38[863], line_37[861], line_36[859], line_35[857], line_34[855], line_33[853], line_32[851], line_31[849], line_30[847], line_29[845], line_28[843], line_27[841], line_26[839], line_25[837], line_24[835], line_23[833], line_22[831], line_21[829], line_20[827], line_19[825], line_18[823], line_17[821], line_16[819], line_15[817], line_14[815], line_13[813], line_12[811], line_11[809], line_10[807], line_9[805], line_8[803], line_7[801], line_6[799], line_5[797], line_4[795], line_3[793], line_2[791], line_1[789], 9'b0};
assign col_1044 = {line_118[1024], line_117[1022], line_116[1020], line_115[1018], line_114[1016], line_113[1014], line_112[1012], line_111[1010], line_110[1008], line_109[1006], line_108[1004], line_107[1002], line_106[1000], line_105[998], line_104[996], line_103[994], line_102[992], line_101[990], line_100[988], line_99[986], line_98[984], line_97[982], line_96[980], line_95[978], line_94[976], line_93[974], line_92[972], line_91[970], line_90[968], line_89[966], line_88[964], line_87[962], line_86[960], line_85[958], line_84[956], line_83[954], line_82[952], line_81[950], line_80[948], line_79[946], line_78[944], line_77[942], line_76[940], line_75[938], line_74[936], line_73[934], line_72[932], line_71[930], line_70[928], line_69[926], line_68[924], line_67[922], line_66[920], line_65[918], line_64[916], line_63[914], line_62[912], line_61[910], line_60[908], line_59[906], line_58[904], line_57[902], line_56[900], line_55[898], line_54[896], line_53[894], line_52[892], line_51[890], line_50[888], line_49[886], line_48[884], line_47[882], line_46[880], line_45[878], line_44[876], line_43[874], line_42[872], line_41[870], line_40[868], line_39[866], line_38[864], line_37[862], line_36[860], line_35[858], line_34[856], line_33[854], line_32[852], line_31[850], line_30[848], line_29[846], line_28[844], line_27[842], line_26[840], line_25[838], line_24[836], line_23[834], line_22[832], line_21[830], line_20[828], line_19[826], line_18[824], line_17[822], line_16[820], line_15[818], line_14[816], line_13[814], line_12[812], line_11[810], line_10[808], line_9[806], line_8[804], line_7[802], line_6[800], line_5[798], line_4[796], line_3[794], line_2[792], line_1[790], 10'b0};
assign col_1045 = {line_118[1025], line_117[1023], line_116[1021], line_115[1019], line_114[1017], line_113[1015], line_112[1013], line_111[1011], line_110[1009], line_109[1007], line_108[1005], line_107[1003], line_106[1001], line_105[999], line_104[997], line_103[995], line_102[993], line_101[991], line_100[989], line_99[987], line_98[985], line_97[983], line_96[981], line_95[979], line_94[977], line_93[975], line_92[973], line_91[971], line_90[969], line_89[967], line_88[965], line_87[963], line_86[961], line_85[959], line_84[957], line_83[955], line_82[953], line_81[951], line_80[949], line_79[947], line_78[945], line_77[943], line_76[941], line_75[939], line_74[937], line_73[935], line_72[933], line_71[931], line_70[929], line_69[927], line_68[925], line_67[923], line_66[921], line_65[919], line_64[917], line_63[915], line_62[913], line_61[911], line_60[909], line_59[907], line_58[905], line_57[903], line_56[901], line_55[899], line_54[897], line_53[895], line_52[893], line_51[891], line_50[889], line_49[887], line_48[885], line_47[883], line_46[881], line_45[879], line_44[877], line_43[875], line_42[873], line_41[871], line_40[869], line_39[867], line_38[865], line_37[863], line_36[861], line_35[859], line_34[857], line_33[855], line_32[853], line_31[851], line_30[849], line_29[847], line_28[845], line_27[843], line_26[841], line_25[839], line_24[837], line_23[835], line_22[833], line_21[831], line_20[829], line_19[827], line_18[825], line_17[823], line_16[821], line_15[819], line_14[817], line_13[815], line_12[813], line_11[811], line_10[809], line_9[807], line_8[805], line_7[803], line_6[801], line_5[799], line_4[797], line_3[795], line_2[793], line_1[791], 10'b0};
assign col_1046 = {line_117[1024], line_116[1022], line_115[1020], line_114[1018], line_113[1016], line_112[1014], line_111[1012], line_110[1010], line_109[1008], line_108[1006], line_107[1004], line_106[1002], line_105[1000], line_104[998], line_103[996], line_102[994], line_101[992], line_100[990], line_99[988], line_98[986], line_97[984], line_96[982], line_95[980], line_94[978], line_93[976], line_92[974], line_91[972], line_90[970], line_89[968], line_88[966], line_87[964], line_86[962], line_85[960], line_84[958], line_83[956], line_82[954], line_81[952], line_80[950], line_79[948], line_78[946], line_77[944], line_76[942], line_75[940], line_74[938], line_73[936], line_72[934], line_71[932], line_70[930], line_69[928], line_68[926], line_67[924], line_66[922], line_65[920], line_64[918], line_63[916], line_62[914], line_61[912], line_60[910], line_59[908], line_58[906], line_57[904], line_56[902], line_55[900], line_54[898], line_53[896], line_52[894], line_51[892], line_50[890], line_49[888], line_48[886], line_47[884], line_46[882], line_45[880], line_44[878], line_43[876], line_42[874], line_41[872], line_40[870], line_39[868], line_38[866], line_37[864], line_36[862], line_35[860], line_34[858], line_33[856], line_32[854], line_31[852], line_30[850], line_29[848], line_28[846], line_27[844], line_26[842], line_25[840], line_24[838], line_23[836], line_22[834], line_21[832], line_20[830], line_19[828], line_18[826], line_17[824], line_16[822], line_15[820], line_14[818], line_13[816], line_12[814], line_11[812], line_10[810], line_9[808], line_8[806], line_7[804], line_6[802], line_5[800], line_4[798], line_3[796], line_2[794], line_1[792], 11'b0};
assign col_1047 = {line_117[1025], line_116[1023], line_115[1021], line_114[1019], line_113[1017], line_112[1015], line_111[1013], line_110[1011], line_109[1009], line_108[1007], line_107[1005], line_106[1003], line_105[1001], line_104[999], line_103[997], line_102[995], line_101[993], line_100[991], line_99[989], line_98[987], line_97[985], line_96[983], line_95[981], line_94[979], line_93[977], line_92[975], line_91[973], line_90[971], line_89[969], line_88[967], line_87[965], line_86[963], line_85[961], line_84[959], line_83[957], line_82[955], line_81[953], line_80[951], line_79[949], line_78[947], line_77[945], line_76[943], line_75[941], line_74[939], line_73[937], line_72[935], line_71[933], line_70[931], line_69[929], line_68[927], line_67[925], line_66[923], line_65[921], line_64[919], line_63[917], line_62[915], line_61[913], line_60[911], line_59[909], line_58[907], line_57[905], line_56[903], line_55[901], line_54[899], line_53[897], line_52[895], line_51[893], line_50[891], line_49[889], line_48[887], line_47[885], line_46[883], line_45[881], line_44[879], line_43[877], line_42[875], line_41[873], line_40[871], line_39[869], line_38[867], line_37[865], line_36[863], line_35[861], line_34[859], line_33[857], line_32[855], line_31[853], line_30[851], line_29[849], line_28[847], line_27[845], line_26[843], line_25[841], line_24[839], line_23[837], line_22[835], line_21[833], line_20[831], line_19[829], line_18[827], line_17[825], line_16[823], line_15[821], line_14[819], line_13[817], line_12[815], line_11[813], line_10[811], line_9[809], line_8[807], line_7[805], line_6[803], line_5[801], line_4[799], line_3[797], line_2[795], line_1[793], 11'b0};
assign col_1048 = {line_116[1024], line_115[1022], line_114[1020], line_113[1018], line_112[1016], line_111[1014], line_110[1012], line_109[1010], line_108[1008], line_107[1006], line_106[1004], line_105[1002], line_104[1000], line_103[998], line_102[996], line_101[994], line_100[992], line_99[990], line_98[988], line_97[986], line_96[984], line_95[982], line_94[980], line_93[978], line_92[976], line_91[974], line_90[972], line_89[970], line_88[968], line_87[966], line_86[964], line_85[962], line_84[960], line_83[958], line_82[956], line_81[954], line_80[952], line_79[950], line_78[948], line_77[946], line_76[944], line_75[942], line_74[940], line_73[938], line_72[936], line_71[934], line_70[932], line_69[930], line_68[928], line_67[926], line_66[924], line_65[922], line_64[920], line_63[918], line_62[916], line_61[914], line_60[912], line_59[910], line_58[908], line_57[906], line_56[904], line_55[902], line_54[900], line_53[898], line_52[896], line_51[894], line_50[892], line_49[890], line_48[888], line_47[886], line_46[884], line_45[882], line_44[880], line_43[878], line_42[876], line_41[874], line_40[872], line_39[870], line_38[868], line_37[866], line_36[864], line_35[862], line_34[860], line_33[858], line_32[856], line_31[854], line_30[852], line_29[850], line_28[848], line_27[846], line_26[844], line_25[842], line_24[840], line_23[838], line_22[836], line_21[834], line_20[832], line_19[830], line_18[828], line_17[826], line_16[824], line_15[822], line_14[820], line_13[818], line_12[816], line_11[814], line_10[812], line_9[810], line_8[808], line_7[806], line_6[804], line_5[802], line_4[800], line_3[798], line_2[796], line_1[794], 12'b0};
assign col_1049 = {line_116[1025], line_115[1023], line_114[1021], line_113[1019], line_112[1017], line_111[1015], line_110[1013], line_109[1011], line_108[1009], line_107[1007], line_106[1005], line_105[1003], line_104[1001], line_103[999], line_102[997], line_101[995], line_100[993], line_99[991], line_98[989], line_97[987], line_96[985], line_95[983], line_94[981], line_93[979], line_92[977], line_91[975], line_90[973], line_89[971], line_88[969], line_87[967], line_86[965], line_85[963], line_84[961], line_83[959], line_82[957], line_81[955], line_80[953], line_79[951], line_78[949], line_77[947], line_76[945], line_75[943], line_74[941], line_73[939], line_72[937], line_71[935], line_70[933], line_69[931], line_68[929], line_67[927], line_66[925], line_65[923], line_64[921], line_63[919], line_62[917], line_61[915], line_60[913], line_59[911], line_58[909], line_57[907], line_56[905], line_55[903], line_54[901], line_53[899], line_52[897], line_51[895], line_50[893], line_49[891], line_48[889], line_47[887], line_46[885], line_45[883], line_44[881], line_43[879], line_42[877], line_41[875], line_40[873], line_39[871], line_38[869], line_37[867], line_36[865], line_35[863], line_34[861], line_33[859], line_32[857], line_31[855], line_30[853], line_29[851], line_28[849], line_27[847], line_26[845], line_25[843], line_24[841], line_23[839], line_22[837], line_21[835], line_20[833], line_19[831], line_18[829], line_17[827], line_16[825], line_15[823], line_14[821], line_13[819], line_12[817], line_11[815], line_10[813], line_9[811], line_8[809], line_7[807], line_6[805], line_5[803], line_4[801], line_3[799], line_2[797], line_1[795], 12'b0};
assign col_1050 = {line_115[1024], line_114[1022], line_113[1020], line_112[1018], line_111[1016], line_110[1014], line_109[1012], line_108[1010], line_107[1008], line_106[1006], line_105[1004], line_104[1002], line_103[1000], line_102[998], line_101[996], line_100[994], line_99[992], line_98[990], line_97[988], line_96[986], line_95[984], line_94[982], line_93[980], line_92[978], line_91[976], line_90[974], line_89[972], line_88[970], line_87[968], line_86[966], line_85[964], line_84[962], line_83[960], line_82[958], line_81[956], line_80[954], line_79[952], line_78[950], line_77[948], line_76[946], line_75[944], line_74[942], line_73[940], line_72[938], line_71[936], line_70[934], line_69[932], line_68[930], line_67[928], line_66[926], line_65[924], line_64[922], line_63[920], line_62[918], line_61[916], line_60[914], line_59[912], line_58[910], line_57[908], line_56[906], line_55[904], line_54[902], line_53[900], line_52[898], line_51[896], line_50[894], line_49[892], line_48[890], line_47[888], line_46[886], line_45[884], line_44[882], line_43[880], line_42[878], line_41[876], line_40[874], line_39[872], line_38[870], line_37[868], line_36[866], line_35[864], line_34[862], line_33[860], line_32[858], line_31[856], line_30[854], line_29[852], line_28[850], line_27[848], line_26[846], line_25[844], line_24[842], line_23[840], line_22[838], line_21[836], line_20[834], line_19[832], line_18[830], line_17[828], line_16[826], line_15[824], line_14[822], line_13[820], line_12[818], line_11[816], line_10[814], line_9[812], line_8[810], line_7[808], line_6[806], line_5[804], line_4[802], line_3[800], line_2[798], line_1[796], 13'b0};
assign col_1051 = {line_115[1025], line_114[1023], line_113[1021], line_112[1019], line_111[1017], line_110[1015], line_109[1013], line_108[1011], line_107[1009], line_106[1007], line_105[1005], line_104[1003], line_103[1001], line_102[999], line_101[997], line_100[995], line_99[993], line_98[991], line_97[989], line_96[987], line_95[985], line_94[983], line_93[981], line_92[979], line_91[977], line_90[975], line_89[973], line_88[971], line_87[969], line_86[967], line_85[965], line_84[963], line_83[961], line_82[959], line_81[957], line_80[955], line_79[953], line_78[951], line_77[949], line_76[947], line_75[945], line_74[943], line_73[941], line_72[939], line_71[937], line_70[935], line_69[933], line_68[931], line_67[929], line_66[927], line_65[925], line_64[923], line_63[921], line_62[919], line_61[917], line_60[915], line_59[913], line_58[911], line_57[909], line_56[907], line_55[905], line_54[903], line_53[901], line_52[899], line_51[897], line_50[895], line_49[893], line_48[891], line_47[889], line_46[887], line_45[885], line_44[883], line_43[881], line_42[879], line_41[877], line_40[875], line_39[873], line_38[871], line_37[869], line_36[867], line_35[865], line_34[863], line_33[861], line_32[859], line_31[857], line_30[855], line_29[853], line_28[851], line_27[849], line_26[847], line_25[845], line_24[843], line_23[841], line_22[839], line_21[837], line_20[835], line_19[833], line_18[831], line_17[829], line_16[827], line_15[825], line_14[823], line_13[821], line_12[819], line_11[817], line_10[815], line_9[813], line_8[811], line_7[809], line_6[807], line_5[805], line_4[803], line_3[801], line_2[799], line_1[797], 13'b0};
assign col_1052 = {line_114[1024], line_113[1022], line_112[1020], line_111[1018], line_110[1016], line_109[1014], line_108[1012], line_107[1010], line_106[1008], line_105[1006], line_104[1004], line_103[1002], line_102[1000], line_101[998], line_100[996], line_99[994], line_98[992], line_97[990], line_96[988], line_95[986], line_94[984], line_93[982], line_92[980], line_91[978], line_90[976], line_89[974], line_88[972], line_87[970], line_86[968], line_85[966], line_84[964], line_83[962], line_82[960], line_81[958], line_80[956], line_79[954], line_78[952], line_77[950], line_76[948], line_75[946], line_74[944], line_73[942], line_72[940], line_71[938], line_70[936], line_69[934], line_68[932], line_67[930], line_66[928], line_65[926], line_64[924], line_63[922], line_62[920], line_61[918], line_60[916], line_59[914], line_58[912], line_57[910], line_56[908], line_55[906], line_54[904], line_53[902], line_52[900], line_51[898], line_50[896], line_49[894], line_48[892], line_47[890], line_46[888], line_45[886], line_44[884], line_43[882], line_42[880], line_41[878], line_40[876], line_39[874], line_38[872], line_37[870], line_36[868], line_35[866], line_34[864], line_33[862], line_32[860], line_31[858], line_30[856], line_29[854], line_28[852], line_27[850], line_26[848], line_25[846], line_24[844], line_23[842], line_22[840], line_21[838], line_20[836], line_19[834], line_18[832], line_17[830], line_16[828], line_15[826], line_14[824], line_13[822], line_12[820], line_11[818], line_10[816], line_9[814], line_8[812], line_7[810], line_6[808], line_5[806], line_4[804], line_3[802], line_2[800], line_1[798], 14'b0};
assign col_1053 = {line_114[1025], line_113[1023], line_112[1021], line_111[1019], line_110[1017], line_109[1015], line_108[1013], line_107[1011], line_106[1009], line_105[1007], line_104[1005], line_103[1003], line_102[1001], line_101[999], line_100[997], line_99[995], line_98[993], line_97[991], line_96[989], line_95[987], line_94[985], line_93[983], line_92[981], line_91[979], line_90[977], line_89[975], line_88[973], line_87[971], line_86[969], line_85[967], line_84[965], line_83[963], line_82[961], line_81[959], line_80[957], line_79[955], line_78[953], line_77[951], line_76[949], line_75[947], line_74[945], line_73[943], line_72[941], line_71[939], line_70[937], line_69[935], line_68[933], line_67[931], line_66[929], line_65[927], line_64[925], line_63[923], line_62[921], line_61[919], line_60[917], line_59[915], line_58[913], line_57[911], line_56[909], line_55[907], line_54[905], line_53[903], line_52[901], line_51[899], line_50[897], line_49[895], line_48[893], line_47[891], line_46[889], line_45[887], line_44[885], line_43[883], line_42[881], line_41[879], line_40[877], line_39[875], line_38[873], line_37[871], line_36[869], line_35[867], line_34[865], line_33[863], line_32[861], line_31[859], line_30[857], line_29[855], line_28[853], line_27[851], line_26[849], line_25[847], line_24[845], line_23[843], line_22[841], line_21[839], line_20[837], line_19[835], line_18[833], line_17[831], line_16[829], line_15[827], line_14[825], line_13[823], line_12[821], line_11[819], line_10[817], line_9[815], line_8[813], line_7[811], line_6[809], line_5[807], line_4[805], line_3[803], line_2[801], line_1[799], 14'b0};
assign col_1054 = {line_113[1024], line_112[1022], line_111[1020], line_110[1018], line_109[1016], line_108[1014], line_107[1012], line_106[1010], line_105[1008], line_104[1006], line_103[1004], line_102[1002], line_101[1000], line_100[998], line_99[996], line_98[994], line_97[992], line_96[990], line_95[988], line_94[986], line_93[984], line_92[982], line_91[980], line_90[978], line_89[976], line_88[974], line_87[972], line_86[970], line_85[968], line_84[966], line_83[964], line_82[962], line_81[960], line_80[958], line_79[956], line_78[954], line_77[952], line_76[950], line_75[948], line_74[946], line_73[944], line_72[942], line_71[940], line_70[938], line_69[936], line_68[934], line_67[932], line_66[930], line_65[928], line_64[926], line_63[924], line_62[922], line_61[920], line_60[918], line_59[916], line_58[914], line_57[912], line_56[910], line_55[908], line_54[906], line_53[904], line_52[902], line_51[900], line_50[898], line_49[896], line_48[894], line_47[892], line_46[890], line_45[888], line_44[886], line_43[884], line_42[882], line_41[880], line_40[878], line_39[876], line_38[874], line_37[872], line_36[870], line_35[868], line_34[866], line_33[864], line_32[862], line_31[860], line_30[858], line_29[856], line_28[854], line_27[852], line_26[850], line_25[848], line_24[846], line_23[844], line_22[842], line_21[840], line_20[838], line_19[836], line_18[834], line_17[832], line_16[830], line_15[828], line_14[826], line_13[824], line_12[822], line_11[820], line_10[818], line_9[816], line_8[814], line_7[812], line_6[810], line_5[808], line_4[806], line_3[804], line_2[802], line_1[800], 15'b0};
assign col_1055 = {line_113[1025], line_112[1023], line_111[1021], line_110[1019], line_109[1017], line_108[1015], line_107[1013], line_106[1011], line_105[1009], line_104[1007], line_103[1005], line_102[1003], line_101[1001], line_100[999], line_99[997], line_98[995], line_97[993], line_96[991], line_95[989], line_94[987], line_93[985], line_92[983], line_91[981], line_90[979], line_89[977], line_88[975], line_87[973], line_86[971], line_85[969], line_84[967], line_83[965], line_82[963], line_81[961], line_80[959], line_79[957], line_78[955], line_77[953], line_76[951], line_75[949], line_74[947], line_73[945], line_72[943], line_71[941], line_70[939], line_69[937], line_68[935], line_67[933], line_66[931], line_65[929], line_64[927], line_63[925], line_62[923], line_61[921], line_60[919], line_59[917], line_58[915], line_57[913], line_56[911], line_55[909], line_54[907], line_53[905], line_52[903], line_51[901], line_50[899], line_49[897], line_48[895], line_47[893], line_46[891], line_45[889], line_44[887], line_43[885], line_42[883], line_41[881], line_40[879], line_39[877], line_38[875], line_37[873], line_36[871], line_35[869], line_34[867], line_33[865], line_32[863], line_31[861], line_30[859], line_29[857], line_28[855], line_27[853], line_26[851], line_25[849], line_24[847], line_23[845], line_22[843], line_21[841], line_20[839], line_19[837], line_18[835], line_17[833], line_16[831], line_15[829], line_14[827], line_13[825], line_12[823], line_11[821], line_10[819], line_9[817], line_8[815], line_7[813], line_6[811], line_5[809], line_4[807], line_3[805], line_2[803], line_1[801], 15'b0};
assign col_1056 = {line_112[1024], line_111[1022], line_110[1020], line_109[1018], line_108[1016], line_107[1014], line_106[1012], line_105[1010], line_104[1008], line_103[1006], line_102[1004], line_101[1002], line_100[1000], line_99[998], line_98[996], line_97[994], line_96[992], line_95[990], line_94[988], line_93[986], line_92[984], line_91[982], line_90[980], line_89[978], line_88[976], line_87[974], line_86[972], line_85[970], line_84[968], line_83[966], line_82[964], line_81[962], line_80[960], line_79[958], line_78[956], line_77[954], line_76[952], line_75[950], line_74[948], line_73[946], line_72[944], line_71[942], line_70[940], line_69[938], line_68[936], line_67[934], line_66[932], line_65[930], line_64[928], line_63[926], line_62[924], line_61[922], line_60[920], line_59[918], line_58[916], line_57[914], line_56[912], line_55[910], line_54[908], line_53[906], line_52[904], line_51[902], line_50[900], line_49[898], line_48[896], line_47[894], line_46[892], line_45[890], line_44[888], line_43[886], line_42[884], line_41[882], line_40[880], line_39[878], line_38[876], line_37[874], line_36[872], line_35[870], line_34[868], line_33[866], line_32[864], line_31[862], line_30[860], line_29[858], line_28[856], line_27[854], line_26[852], line_25[850], line_24[848], line_23[846], line_22[844], line_21[842], line_20[840], line_19[838], line_18[836], line_17[834], line_16[832], line_15[830], line_14[828], line_13[826], line_12[824], line_11[822], line_10[820], line_9[818], line_8[816], line_7[814], line_6[812], line_5[810], line_4[808], line_3[806], line_2[804], line_1[802], 16'b0};
assign col_1057 = {line_112[1025], line_111[1023], line_110[1021], line_109[1019], line_108[1017], line_107[1015], line_106[1013], line_105[1011], line_104[1009], line_103[1007], line_102[1005], line_101[1003], line_100[1001], line_99[999], line_98[997], line_97[995], line_96[993], line_95[991], line_94[989], line_93[987], line_92[985], line_91[983], line_90[981], line_89[979], line_88[977], line_87[975], line_86[973], line_85[971], line_84[969], line_83[967], line_82[965], line_81[963], line_80[961], line_79[959], line_78[957], line_77[955], line_76[953], line_75[951], line_74[949], line_73[947], line_72[945], line_71[943], line_70[941], line_69[939], line_68[937], line_67[935], line_66[933], line_65[931], line_64[929], line_63[927], line_62[925], line_61[923], line_60[921], line_59[919], line_58[917], line_57[915], line_56[913], line_55[911], line_54[909], line_53[907], line_52[905], line_51[903], line_50[901], line_49[899], line_48[897], line_47[895], line_46[893], line_45[891], line_44[889], line_43[887], line_42[885], line_41[883], line_40[881], line_39[879], line_38[877], line_37[875], line_36[873], line_35[871], line_34[869], line_33[867], line_32[865], line_31[863], line_30[861], line_29[859], line_28[857], line_27[855], line_26[853], line_25[851], line_24[849], line_23[847], line_22[845], line_21[843], line_20[841], line_19[839], line_18[837], line_17[835], line_16[833], line_15[831], line_14[829], line_13[827], line_12[825], line_11[823], line_10[821], line_9[819], line_8[817], line_7[815], line_6[813], line_5[811], line_4[809], line_3[807], line_2[805], line_1[803], 16'b0};
assign col_1058 = {line_111[1024], line_110[1022], line_109[1020], line_108[1018], line_107[1016], line_106[1014], line_105[1012], line_104[1010], line_103[1008], line_102[1006], line_101[1004], line_100[1002], line_99[1000], line_98[998], line_97[996], line_96[994], line_95[992], line_94[990], line_93[988], line_92[986], line_91[984], line_90[982], line_89[980], line_88[978], line_87[976], line_86[974], line_85[972], line_84[970], line_83[968], line_82[966], line_81[964], line_80[962], line_79[960], line_78[958], line_77[956], line_76[954], line_75[952], line_74[950], line_73[948], line_72[946], line_71[944], line_70[942], line_69[940], line_68[938], line_67[936], line_66[934], line_65[932], line_64[930], line_63[928], line_62[926], line_61[924], line_60[922], line_59[920], line_58[918], line_57[916], line_56[914], line_55[912], line_54[910], line_53[908], line_52[906], line_51[904], line_50[902], line_49[900], line_48[898], line_47[896], line_46[894], line_45[892], line_44[890], line_43[888], line_42[886], line_41[884], line_40[882], line_39[880], line_38[878], line_37[876], line_36[874], line_35[872], line_34[870], line_33[868], line_32[866], line_31[864], line_30[862], line_29[860], line_28[858], line_27[856], line_26[854], line_25[852], line_24[850], line_23[848], line_22[846], line_21[844], line_20[842], line_19[840], line_18[838], line_17[836], line_16[834], line_15[832], line_14[830], line_13[828], line_12[826], line_11[824], line_10[822], line_9[820], line_8[818], line_7[816], line_6[814], line_5[812], line_4[810], line_3[808], line_2[806], line_1[804], 17'b0};
assign col_1059 = {line_111[1025], line_110[1023], line_109[1021], line_108[1019], line_107[1017], line_106[1015], line_105[1013], line_104[1011], line_103[1009], line_102[1007], line_101[1005], line_100[1003], line_99[1001], line_98[999], line_97[997], line_96[995], line_95[993], line_94[991], line_93[989], line_92[987], line_91[985], line_90[983], line_89[981], line_88[979], line_87[977], line_86[975], line_85[973], line_84[971], line_83[969], line_82[967], line_81[965], line_80[963], line_79[961], line_78[959], line_77[957], line_76[955], line_75[953], line_74[951], line_73[949], line_72[947], line_71[945], line_70[943], line_69[941], line_68[939], line_67[937], line_66[935], line_65[933], line_64[931], line_63[929], line_62[927], line_61[925], line_60[923], line_59[921], line_58[919], line_57[917], line_56[915], line_55[913], line_54[911], line_53[909], line_52[907], line_51[905], line_50[903], line_49[901], line_48[899], line_47[897], line_46[895], line_45[893], line_44[891], line_43[889], line_42[887], line_41[885], line_40[883], line_39[881], line_38[879], line_37[877], line_36[875], line_35[873], line_34[871], line_33[869], line_32[867], line_31[865], line_30[863], line_29[861], line_28[859], line_27[857], line_26[855], line_25[853], line_24[851], line_23[849], line_22[847], line_21[845], line_20[843], line_19[841], line_18[839], line_17[837], line_16[835], line_15[833], line_14[831], line_13[829], line_12[827], line_11[825], line_10[823], line_9[821], line_8[819], line_7[817], line_6[815], line_5[813], line_4[811], line_3[809], line_2[807], line_1[805], 17'b0};
assign col_1060 = {line_110[1024], line_109[1022], line_108[1020], line_107[1018], line_106[1016], line_105[1014], line_104[1012], line_103[1010], line_102[1008], line_101[1006], line_100[1004], line_99[1002], line_98[1000], line_97[998], line_96[996], line_95[994], line_94[992], line_93[990], line_92[988], line_91[986], line_90[984], line_89[982], line_88[980], line_87[978], line_86[976], line_85[974], line_84[972], line_83[970], line_82[968], line_81[966], line_80[964], line_79[962], line_78[960], line_77[958], line_76[956], line_75[954], line_74[952], line_73[950], line_72[948], line_71[946], line_70[944], line_69[942], line_68[940], line_67[938], line_66[936], line_65[934], line_64[932], line_63[930], line_62[928], line_61[926], line_60[924], line_59[922], line_58[920], line_57[918], line_56[916], line_55[914], line_54[912], line_53[910], line_52[908], line_51[906], line_50[904], line_49[902], line_48[900], line_47[898], line_46[896], line_45[894], line_44[892], line_43[890], line_42[888], line_41[886], line_40[884], line_39[882], line_38[880], line_37[878], line_36[876], line_35[874], line_34[872], line_33[870], line_32[868], line_31[866], line_30[864], line_29[862], line_28[860], line_27[858], line_26[856], line_25[854], line_24[852], line_23[850], line_22[848], line_21[846], line_20[844], line_19[842], line_18[840], line_17[838], line_16[836], line_15[834], line_14[832], line_13[830], line_12[828], line_11[826], line_10[824], line_9[822], line_8[820], line_7[818], line_6[816], line_5[814], line_4[812], line_3[810], line_2[808], line_1[806], 18'b0};
assign col_1061 = {line_110[1025], line_109[1023], line_108[1021], line_107[1019], line_106[1017], line_105[1015], line_104[1013], line_103[1011], line_102[1009], line_101[1007], line_100[1005], line_99[1003], line_98[1001], line_97[999], line_96[997], line_95[995], line_94[993], line_93[991], line_92[989], line_91[987], line_90[985], line_89[983], line_88[981], line_87[979], line_86[977], line_85[975], line_84[973], line_83[971], line_82[969], line_81[967], line_80[965], line_79[963], line_78[961], line_77[959], line_76[957], line_75[955], line_74[953], line_73[951], line_72[949], line_71[947], line_70[945], line_69[943], line_68[941], line_67[939], line_66[937], line_65[935], line_64[933], line_63[931], line_62[929], line_61[927], line_60[925], line_59[923], line_58[921], line_57[919], line_56[917], line_55[915], line_54[913], line_53[911], line_52[909], line_51[907], line_50[905], line_49[903], line_48[901], line_47[899], line_46[897], line_45[895], line_44[893], line_43[891], line_42[889], line_41[887], line_40[885], line_39[883], line_38[881], line_37[879], line_36[877], line_35[875], line_34[873], line_33[871], line_32[869], line_31[867], line_30[865], line_29[863], line_28[861], line_27[859], line_26[857], line_25[855], line_24[853], line_23[851], line_22[849], line_21[847], line_20[845], line_19[843], line_18[841], line_17[839], line_16[837], line_15[835], line_14[833], line_13[831], line_12[829], line_11[827], line_10[825], line_9[823], line_8[821], line_7[819], line_6[817], line_5[815], line_4[813], line_3[811], line_2[809], line_1[807], 18'b0};
assign col_1062 = {line_109[1024], line_108[1022], line_107[1020], line_106[1018], line_105[1016], line_104[1014], line_103[1012], line_102[1010], line_101[1008], line_100[1006], line_99[1004], line_98[1002], line_97[1000], line_96[998], line_95[996], line_94[994], line_93[992], line_92[990], line_91[988], line_90[986], line_89[984], line_88[982], line_87[980], line_86[978], line_85[976], line_84[974], line_83[972], line_82[970], line_81[968], line_80[966], line_79[964], line_78[962], line_77[960], line_76[958], line_75[956], line_74[954], line_73[952], line_72[950], line_71[948], line_70[946], line_69[944], line_68[942], line_67[940], line_66[938], line_65[936], line_64[934], line_63[932], line_62[930], line_61[928], line_60[926], line_59[924], line_58[922], line_57[920], line_56[918], line_55[916], line_54[914], line_53[912], line_52[910], line_51[908], line_50[906], line_49[904], line_48[902], line_47[900], line_46[898], line_45[896], line_44[894], line_43[892], line_42[890], line_41[888], line_40[886], line_39[884], line_38[882], line_37[880], line_36[878], line_35[876], line_34[874], line_33[872], line_32[870], line_31[868], line_30[866], line_29[864], line_28[862], line_27[860], line_26[858], line_25[856], line_24[854], line_23[852], line_22[850], line_21[848], line_20[846], line_19[844], line_18[842], line_17[840], line_16[838], line_15[836], line_14[834], line_13[832], line_12[830], line_11[828], line_10[826], line_9[824], line_8[822], line_7[820], line_6[818], line_5[816], line_4[814], line_3[812], line_2[810], line_1[808], 19'b0};
assign col_1063 = {line_109[1025], line_108[1023], line_107[1021], line_106[1019], line_105[1017], line_104[1015], line_103[1013], line_102[1011], line_101[1009], line_100[1007], line_99[1005], line_98[1003], line_97[1001], line_96[999], line_95[997], line_94[995], line_93[993], line_92[991], line_91[989], line_90[987], line_89[985], line_88[983], line_87[981], line_86[979], line_85[977], line_84[975], line_83[973], line_82[971], line_81[969], line_80[967], line_79[965], line_78[963], line_77[961], line_76[959], line_75[957], line_74[955], line_73[953], line_72[951], line_71[949], line_70[947], line_69[945], line_68[943], line_67[941], line_66[939], line_65[937], line_64[935], line_63[933], line_62[931], line_61[929], line_60[927], line_59[925], line_58[923], line_57[921], line_56[919], line_55[917], line_54[915], line_53[913], line_52[911], line_51[909], line_50[907], line_49[905], line_48[903], line_47[901], line_46[899], line_45[897], line_44[895], line_43[893], line_42[891], line_41[889], line_40[887], line_39[885], line_38[883], line_37[881], line_36[879], line_35[877], line_34[875], line_33[873], line_32[871], line_31[869], line_30[867], line_29[865], line_28[863], line_27[861], line_26[859], line_25[857], line_24[855], line_23[853], line_22[851], line_21[849], line_20[847], line_19[845], line_18[843], line_17[841], line_16[839], line_15[837], line_14[835], line_13[833], line_12[831], line_11[829], line_10[827], line_9[825], line_8[823], line_7[821], line_6[819], line_5[817], line_4[815], line_3[813], line_2[811], line_1[809], 19'b0};
assign col_1064 = {line_108[1024], line_107[1022], line_106[1020], line_105[1018], line_104[1016], line_103[1014], line_102[1012], line_101[1010], line_100[1008], line_99[1006], line_98[1004], line_97[1002], line_96[1000], line_95[998], line_94[996], line_93[994], line_92[992], line_91[990], line_90[988], line_89[986], line_88[984], line_87[982], line_86[980], line_85[978], line_84[976], line_83[974], line_82[972], line_81[970], line_80[968], line_79[966], line_78[964], line_77[962], line_76[960], line_75[958], line_74[956], line_73[954], line_72[952], line_71[950], line_70[948], line_69[946], line_68[944], line_67[942], line_66[940], line_65[938], line_64[936], line_63[934], line_62[932], line_61[930], line_60[928], line_59[926], line_58[924], line_57[922], line_56[920], line_55[918], line_54[916], line_53[914], line_52[912], line_51[910], line_50[908], line_49[906], line_48[904], line_47[902], line_46[900], line_45[898], line_44[896], line_43[894], line_42[892], line_41[890], line_40[888], line_39[886], line_38[884], line_37[882], line_36[880], line_35[878], line_34[876], line_33[874], line_32[872], line_31[870], line_30[868], line_29[866], line_28[864], line_27[862], line_26[860], line_25[858], line_24[856], line_23[854], line_22[852], line_21[850], line_20[848], line_19[846], line_18[844], line_17[842], line_16[840], line_15[838], line_14[836], line_13[834], line_12[832], line_11[830], line_10[828], line_9[826], line_8[824], line_7[822], line_6[820], line_5[818], line_4[816], line_3[814], line_2[812], line_1[810], 20'b0};
assign col_1065 = {line_108[1025], line_107[1023], line_106[1021], line_105[1019], line_104[1017], line_103[1015], line_102[1013], line_101[1011], line_100[1009], line_99[1007], line_98[1005], line_97[1003], line_96[1001], line_95[999], line_94[997], line_93[995], line_92[993], line_91[991], line_90[989], line_89[987], line_88[985], line_87[983], line_86[981], line_85[979], line_84[977], line_83[975], line_82[973], line_81[971], line_80[969], line_79[967], line_78[965], line_77[963], line_76[961], line_75[959], line_74[957], line_73[955], line_72[953], line_71[951], line_70[949], line_69[947], line_68[945], line_67[943], line_66[941], line_65[939], line_64[937], line_63[935], line_62[933], line_61[931], line_60[929], line_59[927], line_58[925], line_57[923], line_56[921], line_55[919], line_54[917], line_53[915], line_52[913], line_51[911], line_50[909], line_49[907], line_48[905], line_47[903], line_46[901], line_45[899], line_44[897], line_43[895], line_42[893], line_41[891], line_40[889], line_39[887], line_38[885], line_37[883], line_36[881], line_35[879], line_34[877], line_33[875], line_32[873], line_31[871], line_30[869], line_29[867], line_28[865], line_27[863], line_26[861], line_25[859], line_24[857], line_23[855], line_22[853], line_21[851], line_20[849], line_19[847], line_18[845], line_17[843], line_16[841], line_15[839], line_14[837], line_13[835], line_12[833], line_11[831], line_10[829], line_9[827], line_8[825], line_7[823], line_6[821], line_5[819], line_4[817], line_3[815], line_2[813], line_1[811], 20'b0};
assign col_1066 = {line_107[1024], line_106[1022], line_105[1020], line_104[1018], line_103[1016], line_102[1014], line_101[1012], line_100[1010], line_99[1008], line_98[1006], line_97[1004], line_96[1002], line_95[1000], line_94[998], line_93[996], line_92[994], line_91[992], line_90[990], line_89[988], line_88[986], line_87[984], line_86[982], line_85[980], line_84[978], line_83[976], line_82[974], line_81[972], line_80[970], line_79[968], line_78[966], line_77[964], line_76[962], line_75[960], line_74[958], line_73[956], line_72[954], line_71[952], line_70[950], line_69[948], line_68[946], line_67[944], line_66[942], line_65[940], line_64[938], line_63[936], line_62[934], line_61[932], line_60[930], line_59[928], line_58[926], line_57[924], line_56[922], line_55[920], line_54[918], line_53[916], line_52[914], line_51[912], line_50[910], line_49[908], line_48[906], line_47[904], line_46[902], line_45[900], line_44[898], line_43[896], line_42[894], line_41[892], line_40[890], line_39[888], line_38[886], line_37[884], line_36[882], line_35[880], line_34[878], line_33[876], line_32[874], line_31[872], line_30[870], line_29[868], line_28[866], line_27[864], line_26[862], line_25[860], line_24[858], line_23[856], line_22[854], line_21[852], line_20[850], line_19[848], line_18[846], line_17[844], line_16[842], line_15[840], line_14[838], line_13[836], line_12[834], line_11[832], line_10[830], line_9[828], line_8[826], line_7[824], line_6[822], line_5[820], line_4[818], line_3[816], line_2[814], line_1[812], 21'b0};
assign col_1067 = {line_107[1025], line_106[1023], line_105[1021], line_104[1019], line_103[1017], line_102[1015], line_101[1013], line_100[1011], line_99[1009], line_98[1007], line_97[1005], line_96[1003], line_95[1001], line_94[999], line_93[997], line_92[995], line_91[993], line_90[991], line_89[989], line_88[987], line_87[985], line_86[983], line_85[981], line_84[979], line_83[977], line_82[975], line_81[973], line_80[971], line_79[969], line_78[967], line_77[965], line_76[963], line_75[961], line_74[959], line_73[957], line_72[955], line_71[953], line_70[951], line_69[949], line_68[947], line_67[945], line_66[943], line_65[941], line_64[939], line_63[937], line_62[935], line_61[933], line_60[931], line_59[929], line_58[927], line_57[925], line_56[923], line_55[921], line_54[919], line_53[917], line_52[915], line_51[913], line_50[911], line_49[909], line_48[907], line_47[905], line_46[903], line_45[901], line_44[899], line_43[897], line_42[895], line_41[893], line_40[891], line_39[889], line_38[887], line_37[885], line_36[883], line_35[881], line_34[879], line_33[877], line_32[875], line_31[873], line_30[871], line_29[869], line_28[867], line_27[865], line_26[863], line_25[861], line_24[859], line_23[857], line_22[855], line_21[853], line_20[851], line_19[849], line_18[847], line_17[845], line_16[843], line_15[841], line_14[839], line_13[837], line_12[835], line_11[833], line_10[831], line_9[829], line_8[827], line_7[825], line_6[823], line_5[821], line_4[819], line_3[817], line_2[815], line_1[813], 21'b0};
assign col_1068 = {line_106[1024], line_105[1022], line_104[1020], line_103[1018], line_102[1016], line_101[1014], line_100[1012], line_99[1010], line_98[1008], line_97[1006], line_96[1004], line_95[1002], line_94[1000], line_93[998], line_92[996], line_91[994], line_90[992], line_89[990], line_88[988], line_87[986], line_86[984], line_85[982], line_84[980], line_83[978], line_82[976], line_81[974], line_80[972], line_79[970], line_78[968], line_77[966], line_76[964], line_75[962], line_74[960], line_73[958], line_72[956], line_71[954], line_70[952], line_69[950], line_68[948], line_67[946], line_66[944], line_65[942], line_64[940], line_63[938], line_62[936], line_61[934], line_60[932], line_59[930], line_58[928], line_57[926], line_56[924], line_55[922], line_54[920], line_53[918], line_52[916], line_51[914], line_50[912], line_49[910], line_48[908], line_47[906], line_46[904], line_45[902], line_44[900], line_43[898], line_42[896], line_41[894], line_40[892], line_39[890], line_38[888], line_37[886], line_36[884], line_35[882], line_34[880], line_33[878], line_32[876], line_31[874], line_30[872], line_29[870], line_28[868], line_27[866], line_26[864], line_25[862], line_24[860], line_23[858], line_22[856], line_21[854], line_20[852], line_19[850], line_18[848], line_17[846], line_16[844], line_15[842], line_14[840], line_13[838], line_12[836], line_11[834], line_10[832], line_9[830], line_8[828], line_7[826], line_6[824], line_5[822], line_4[820], line_3[818], line_2[816], line_1[814], 22'b0};
assign col_1069 = {line_106[1025], line_105[1023], line_104[1021], line_103[1019], line_102[1017], line_101[1015], line_100[1013], line_99[1011], line_98[1009], line_97[1007], line_96[1005], line_95[1003], line_94[1001], line_93[999], line_92[997], line_91[995], line_90[993], line_89[991], line_88[989], line_87[987], line_86[985], line_85[983], line_84[981], line_83[979], line_82[977], line_81[975], line_80[973], line_79[971], line_78[969], line_77[967], line_76[965], line_75[963], line_74[961], line_73[959], line_72[957], line_71[955], line_70[953], line_69[951], line_68[949], line_67[947], line_66[945], line_65[943], line_64[941], line_63[939], line_62[937], line_61[935], line_60[933], line_59[931], line_58[929], line_57[927], line_56[925], line_55[923], line_54[921], line_53[919], line_52[917], line_51[915], line_50[913], line_49[911], line_48[909], line_47[907], line_46[905], line_45[903], line_44[901], line_43[899], line_42[897], line_41[895], line_40[893], line_39[891], line_38[889], line_37[887], line_36[885], line_35[883], line_34[881], line_33[879], line_32[877], line_31[875], line_30[873], line_29[871], line_28[869], line_27[867], line_26[865], line_25[863], line_24[861], line_23[859], line_22[857], line_21[855], line_20[853], line_19[851], line_18[849], line_17[847], line_16[845], line_15[843], line_14[841], line_13[839], line_12[837], line_11[835], line_10[833], line_9[831], line_8[829], line_7[827], line_6[825], line_5[823], line_4[821], line_3[819], line_2[817], line_1[815], 22'b0};
assign col_1070 = {line_105[1024], line_104[1022], line_103[1020], line_102[1018], line_101[1016], line_100[1014], line_99[1012], line_98[1010], line_97[1008], line_96[1006], line_95[1004], line_94[1002], line_93[1000], line_92[998], line_91[996], line_90[994], line_89[992], line_88[990], line_87[988], line_86[986], line_85[984], line_84[982], line_83[980], line_82[978], line_81[976], line_80[974], line_79[972], line_78[970], line_77[968], line_76[966], line_75[964], line_74[962], line_73[960], line_72[958], line_71[956], line_70[954], line_69[952], line_68[950], line_67[948], line_66[946], line_65[944], line_64[942], line_63[940], line_62[938], line_61[936], line_60[934], line_59[932], line_58[930], line_57[928], line_56[926], line_55[924], line_54[922], line_53[920], line_52[918], line_51[916], line_50[914], line_49[912], line_48[910], line_47[908], line_46[906], line_45[904], line_44[902], line_43[900], line_42[898], line_41[896], line_40[894], line_39[892], line_38[890], line_37[888], line_36[886], line_35[884], line_34[882], line_33[880], line_32[878], line_31[876], line_30[874], line_29[872], line_28[870], line_27[868], line_26[866], line_25[864], line_24[862], line_23[860], line_22[858], line_21[856], line_20[854], line_19[852], line_18[850], line_17[848], line_16[846], line_15[844], line_14[842], line_13[840], line_12[838], line_11[836], line_10[834], line_9[832], line_8[830], line_7[828], line_6[826], line_5[824], line_4[822], line_3[820], line_2[818], line_1[816], 23'b0};
assign col_1071 = {line_105[1025], line_104[1023], line_103[1021], line_102[1019], line_101[1017], line_100[1015], line_99[1013], line_98[1011], line_97[1009], line_96[1007], line_95[1005], line_94[1003], line_93[1001], line_92[999], line_91[997], line_90[995], line_89[993], line_88[991], line_87[989], line_86[987], line_85[985], line_84[983], line_83[981], line_82[979], line_81[977], line_80[975], line_79[973], line_78[971], line_77[969], line_76[967], line_75[965], line_74[963], line_73[961], line_72[959], line_71[957], line_70[955], line_69[953], line_68[951], line_67[949], line_66[947], line_65[945], line_64[943], line_63[941], line_62[939], line_61[937], line_60[935], line_59[933], line_58[931], line_57[929], line_56[927], line_55[925], line_54[923], line_53[921], line_52[919], line_51[917], line_50[915], line_49[913], line_48[911], line_47[909], line_46[907], line_45[905], line_44[903], line_43[901], line_42[899], line_41[897], line_40[895], line_39[893], line_38[891], line_37[889], line_36[887], line_35[885], line_34[883], line_33[881], line_32[879], line_31[877], line_30[875], line_29[873], line_28[871], line_27[869], line_26[867], line_25[865], line_24[863], line_23[861], line_22[859], line_21[857], line_20[855], line_19[853], line_18[851], line_17[849], line_16[847], line_15[845], line_14[843], line_13[841], line_12[839], line_11[837], line_10[835], line_9[833], line_8[831], line_7[829], line_6[827], line_5[825], line_4[823], line_3[821], line_2[819], line_1[817], 23'b0};
assign col_1072 = {line_104[1024], line_103[1022], line_102[1020], line_101[1018], line_100[1016], line_99[1014], line_98[1012], line_97[1010], line_96[1008], line_95[1006], line_94[1004], line_93[1002], line_92[1000], line_91[998], line_90[996], line_89[994], line_88[992], line_87[990], line_86[988], line_85[986], line_84[984], line_83[982], line_82[980], line_81[978], line_80[976], line_79[974], line_78[972], line_77[970], line_76[968], line_75[966], line_74[964], line_73[962], line_72[960], line_71[958], line_70[956], line_69[954], line_68[952], line_67[950], line_66[948], line_65[946], line_64[944], line_63[942], line_62[940], line_61[938], line_60[936], line_59[934], line_58[932], line_57[930], line_56[928], line_55[926], line_54[924], line_53[922], line_52[920], line_51[918], line_50[916], line_49[914], line_48[912], line_47[910], line_46[908], line_45[906], line_44[904], line_43[902], line_42[900], line_41[898], line_40[896], line_39[894], line_38[892], line_37[890], line_36[888], line_35[886], line_34[884], line_33[882], line_32[880], line_31[878], line_30[876], line_29[874], line_28[872], line_27[870], line_26[868], line_25[866], line_24[864], line_23[862], line_22[860], line_21[858], line_20[856], line_19[854], line_18[852], line_17[850], line_16[848], line_15[846], line_14[844], line_13[842], line_12[840], line_11[838], line_10[836], line_9[834], line_8[832], line_7[830], line_6[828], line_5[826], line_4[824], line_3[822], line_2[820], line_1[818], 24'b0};
assign col_1073 = {line_104[1025], line_103[1023], line_102[1021], line_101[1019], line_100[1017], line_99[1015], line_98[1013], line_97[1011], line_96[1009], line_95[1007], line_94[1005], line_93[1003], line_92[1001], line_91[999], line_90[997], line_89[995], line_88[993], line_87[991], line_86[989], line_85[987], line_84[985], line_83[983], line_82[981], line_81[979], line_80[977], line_79[975], line_78[973], line_77[971], line_76[969], line_75[967], line_74[965], line_73[963], line_72[961], line_71[959], line_70[957], line_69[955], line_68[953], line_67[951], line_66[949], line_65[947], line_64[945], line_63[943], line_62[941], line_61[939], line_60[937], line_59[935], line_58[933], line_57[931], line_56[929], line_55[927], line_54[925], line_53[923], line_52[921], line_51[919], line_50[917], line_49[915], line_48[913], line_47[911], line_46[909], line_45[907], line_44[905], line_43[903], line_42[901], line_41[899], line_40[897], line_39[895], line_38[893], line_37[891], line_36[889], line_35[887], line_34[885], line_33[883], line_32[881], line_31[879], line_30[877], line_29[875], line_28[873], line_27[871], line_26[869], line_25[867], line_24[865], line_23[863], line_22[861], line_21[859], line_20[857], line_19[855], line_18[853], line_17[851], line_16[849], line_15[847], line_14[845], line_13[843], line_12[841], line_11[839], line_10[837], line_9[835], line_8[833], line_7[831], line_6[829], line_5[827], line_4[825], line_3[823], line_2[821], line_1[819], 24'b0};
assign col_1074 = {line_103[1024], line_102[1022], line_101[1020], line_100[1018], line_99[1016], line_98[1014], line_97[1012], line_96[1010], line_95[1008], line_94[1006], line_93[1004], line_92[1002], line_91[1000], line_90[998], line_89[996], line_88[994], line_87[992], line_86[990], line_85[988], line_84[986], line_83[984], line_82[982], line_81[980], line_80[978], line_79[976], line_78[974], line_77[972], line_76[970], line_75[968], line_74[966], line_73[964], line_72[962], line_71[960], line_70[958], line_69[956], line_68[954], line_67[952], line_66[950], line_65[948], line_64[946], line_63[944], line_62[942], line_61[940], line_60[938], line_59[936], line_58[934], line_57[932], line_56[930], line_55[928], line_54[926], line_53[924], line_52[922], line_51[920], line_50[918], line_49[916], line_48[914], line_47[912], line_46[910], line_45[908], line_44[906], line_43[904], line_42[902], line_41[900], line_40[898], line_39[896], line_38[894], line_37[892], line_36[890], line_35[888], line_34[886], line_33[884], line_32[882], line_31[880], line_30[878], line_29[876], line_28[874], line_27[872], line_26[870], line_25[868], line_24[866], line_23[864], line_22[862], line_21[860], line_20[858], line_19[856], line_18[854], line_17[852], line_16[850], line_15[848], line_14[846], line_13[844], line_12[842], line_11[840], line_10[838], line_9[836], line_8[834], line_7[832], line_6[830], line_5[828], line_4[826], line_3[824], line_2[822], line_1[820], 25'b0};
assign col_1075 = {line_103[1025], line_102[1023], line_101[1021], line_100[1019], line_99[1017], line_98[1015], line_97[1013], line_96[1011], line_95[1009], line_94[1007], line_93[1005], line_92[1003], line_91[1001], line_90[999], line_89[997], line_88[995], line_87[993], line_86[991], line_85[989], line_84[987], line_83[985], line_82[983], line_81[981], line_80[979], line_79[977], line_78[975], line_77[973], line_76[971], line_75[969], line_74[967], line_73[965], line_72[963], line_71[961], line_70[959], line_69[957], line_68[955], line_67[953], line_66[951], line_65[949], line_64[947], line_63[945], line_62[943], line_61[941], line_60[939], line_59[937], line_58[935], line_57[933], line_56[931], line_55[929], line_54[927], line_53[925], line_52[923], line_51[921], line_50[919], line_49[917], line_48[915], line_47[913], line_46[911], line_45[909], line_44[907], line_43[905], line_42[903], line_41[901], line_40[899], line_39[897], line_38[895], line_37[893], line_36[891], line_35[889], line_34[887], line_33[885], line_32[883], line_31[881], line_30[879], line_29[877], line_28[875], line_27[873], line_26[871], line_25[869], line_24[867], line_23[865], line_22[863], line_21[861], line_20[859], line_19[857], line_18[855], line_17[853], line_16[851], line_15[849], line_14[847], line_13[845], line_12[843], line_11[841], line_10[839], line_9[837], line_8[835], line_7[833], line_6[831], line_5[829], line_4[827], line_3[825], line_2[823], line_1[821], 25'b0};
assign col_1076 = {line_102[1024], line_101[1022], line_100[1020], line_99[1018], line_98[1016], line_97[1014], line_96[1012], line_95[1010], line_94[1008], line_93[1006], line_92[1004], line_91[1002], line_90[1000], line_89[998], line_88[996], line_87[994], line_86[992], line_85[990], line_84[988], line_83[986], line_82[984], line_81[982], line_80[980], line_79[978], line_78[976], line_77[974], line_76[972], line_75[970], line_74[968], line_73[966], line_72[964], line_71[962], line_70[960], line_69[958], line_68[956], line_67[954], line_66[952], line_65[950], line_64[948], line_63[946], line_62[944], line_61[942], line_60[940], line_59[938], line_58[936], line_57[934], line_56[932], line_55[930], line_54[928], line_53[926], line_52[924], line_51[922], line_50[920], line_49[918], line_48[916], line_47[914], line_46[912], line_45[910], line_44[908], line_43[906], line_42[904], line_41[902], line_40[900], line_39[898], line_38[896], line_37[894], line_36[892], line_35[890], line_34[888], line_33[886], line_32[884], line_31[882], line_30[880], line_29[878], line_28[876], line_27[874], line_26[872], line_25[870], line_24[868], line_23[866], line_22[864], line_21[862], line_20[860], line_19[858], line_18[856], line_17[854], line_16[852], line_15[850], line_14[848], line_13[846], line_12[844], line_11[842], line_10[840], line_9[838], line_8[836], line_7[834], line_6[832], line_5[830], line_4[828], line_3[826], line_2[824], line_1[822], 26'b0};
assign col_1077 = {line_102[1025], line_101[1023], line_100[1021], line_99[1019], line_98[1017], line_97[1015], line_96[1013], line_95[1011], line_94[1009], line_93[1007], line_92[1005], line_91[1003], line_90[1001], line_89[999], line_88[997], line_87[995], line_86[993], line_85[991], line_84[989], line_83[987], line_82[985], line_81[983], line_80[981], line_79[979], line_78[977], line_77[975], line_76[973], line_75[971], line_74[969], line_73[967], line_72[965], line_71[963], line_70[961], line_69[959], line_68[957], line_67[955], line_66[953], line_65[951], line_64[949], line_63[947], line_62[945], line_61[943], line_60[941], line_59[939], line_58[937], line_57[935], line_56[933], line_55[931], line_54[929], line_53[927], line_52[925], line_51[923], line_50[921], line_49[919], line_48[917], line_47[915], line_46[913], line_45[911], line_44[909], line_43[907], line_42[905], line_41[903], line_40[901], line_39[899], line_38[897], line_37[895], line_36[893], line_35[891], line_34[889], line_33[887], line_32[885], line_31[883], line_30[881], line_29[879], line_28[877], line_27[875], line_26[873], line_25[871], line_24[869], line_23[867], line_22[865], line_21[863], line_20[861], line_19[859], line_18[857], line_17[855], line_16[853], line_15[851], line_14[849], line_13[847], line_12[845], line_11[843], line_10[841], line_9[839], line_8[837], line_7[835], line_6[833], line_5[831], line_4[829], line_3[827], line_2[825], line_1[823], 26'b0};
assign col_1078 = {line_101[1024], line_100[1022], line_99[1020], line_98[1018], line_97[1016], line_96[1014], line_95[1012], line_94[1010], line_93[1008], line_92[1006], line_91[1004], line_90[1002], line_89[1000], line_88[998], line_87[996], line_86[994], line_85[992], line_84[990], line_83[988], line_82[986], line_81[984], line_80[982], line_79[980], line_78[978], line_77[976], line_76[974], line_75[972], line_74[970], line_73[968], line_72[966], line_71[964], line_70[962], line_69[960], line_68[958], line_67[956], line_66[954], line_65[952], line_64[950], line_63[948], line_62[946], line_61[944], line_60[942], line_59[940], line_58[938], line_57[936], line_56[934], line_55[932], line_54[930], line_53[928], line_52[926], line_51[924], line_50[922], line_49[920], line_48[918], line_47[916], line_46[914], line_45[912], line_44[910], line_43[908], line_42[906], line_41[904], line_40[902], line_39[900], line_38[898], line_37[896], line_36[894], line_35[892], line_34[890], line_33[888], line_32[886], line_31[884], line_30[882], line_29[880], line_28[878], line_27[876], line_26[874], line_25[872], line_24[870], line_23[868], line_22[866], line_21[864], line_20[862], line_19[860], line_18[858], line_17[856], line_16[854], line_15[852], line_14[850], line_13[848], line_12[846], line_11[844], line_10[842], line_9[840], line_8[838], line_7[836], line_6[834], line_5[832], line_4[830], line_3[828], line_2[826], line_1[824], 27'b0};
assign col_1079 = {line_101[1025], line_100[1023], line_99[1021], line_98[1019], line_97[1017], line_96[1015], line_95[1013], line_94[1011], line_93[1009], line_92[1007], line_91[1005], line_90[1003], line_89[1001], line_88[999], line_87[997], line_86[995], line_85[993], line_84[991], line_83[989], line_82[987], line_81[985], line_80[983], line_79[981], line_78[979], line_77[977], line_76[975], line_75[973], line_74[971], line_73[969], line_72[967], line_71[965], line_70[963], line_69[961], line_68[959], line_67[957], line_66[955], line_65[953], line_64[951], line_63[949], line_62[947], line_61[945], line_60[943], line_59[941], line_58[939], line_57[937], line_56[935], line_55[933], line_54[931], line_53[929], line_52[927], line_51[925], line_50[923], line_49[921], line_48[919], line_47[917], line_46[915], line_45[913], line_44[911], line_43[909], line_42[907], line_41[905], line_40[903], line_39[901], line_38[899], line_37[897], line_36[895], line_35[893], line_34[891], line_33[889], line_32[887], line_31[885], line_30[883], line_29[881], line_28[879], line_27[877], line_26[875], line_25[873], line_24[871], line_23[869], line_22[867], line_21[865], line_20[863], line_19[861], line_18[859], line_17[857], line_16[855], line_15[853], line_14[851], line_13[849], line_12[847], line_11[845], line_10[843], line_9[841], line_8[839], line_7[837], line_6[835], line_5[833], line_4[831], line_3[829], line_2[827], line_1[825], 27'b0};
assign col_1080 = {line_100[1024], line_99[1022], line_98[1020], line_97[1018], line_96[1016], line_95[1014], line_94[1012], line_93[1010], line_92[1008], line_91[1006], line_90[1004], line_89[1002], line_88[1000], line_87[998], line_86[996], line_85[994], line_84[992], line_83[990], line_82[988], line_81[986], line_80[984], line_79[982], line_78[980], line_77[978], line_76[976], line_75[974], line_74[972], line_73[970], line_72[968], line_71[966], line_70[964], line_69[962], line_68[960], line_67[958], line_66[956], line_65[954], line_64[952], line_63[950], line_62[948], line_61[946], line_60[944], line_59[942], line_58[940], line_57[938], line_56[936], line_55[934], line_54[932], line_53[930], line_52[928], line_51[926], line_50[924], line_49[922], line_48[920], line_47[918], line_46[916], line_45[914], line_44[912], line_43[910], line_42[908], line_41[906], line_40[904], line_39[902], line_38[900], line_37[898], line_36[896], line_35[894], line_34[892], line_33[890], line_32[888], line_31[886], line_30[884], line_29[882], line_28[880], line_27[878], line_26[876], line_25[874], line_24[872], line_23[870], line_22[868], line_21[866], line_20[864], line_19[862], line_18[860], line_17[858], line_16[856], line_15[854], line_14[852], line_13[850], line_12[848], line_11[846], line_10[844], line_9[842], line_8[840], line_7[838], line_6[836], line_5[834], line_4[832], line_3[830], line_2[828], line_1[826], 28'b0};
assign col_1081 = {line_100[1025], line_99[1023], line_98[1021], line_97[1019], line_96[1017], line_95[1015], line_94[1013], line_93[1011], line_92[1009], line_91[1007], line_90[1005], line_89[1003], line_88[1001], line_87[999], line_86[997], line_85[995], line_84[993], line_83[991], line_82[989], line_81[987], line_80[985], line_79[983], line_78[981], line_77[979], line_76[977], line_75[975], line_74[973], line_73[971], line_72[969], line_71[967], line_70[965], line_69[963], line_68[961], line_67[959], line_66[957], line_65[955], line_64[953], line_63[951], line_62[949], line_61[947], line_60[945], line_59[943], line_58[941], line_57[939], line_56[937], line_55[935], line_54[933], line_53[931], line_52[929], line_51[927], line_50[925], line_49[923], line_48[921], line_47[919], line_46[917], line_45[915], line_44[913], line_43[911], line_42[909], line_41[907], line_40[905], line_39[903], line_38[901], line_37[899], line_36[897], line_35[895], line_34[893], line_33[891], line_32[889], line_31[887], line_30[885], line_29[883], line_28[881], line_27[879], line_26[877], line_25[875], line_24[873], line_23[871], line_22[869], line_21[867], line_20[865], line_19[863], line_18[861], line_17[859], line_16[857], line_15[855], line_14[853], line_13[851], line_12[849], line_11[847], line_10[845], line_9[843], line_8[841], line_7[839], line_6[837], line_5[835], line_4[833], line_3[831], line_2[829], line_1[827], 28'b0};
assign col_1082 = {line_99[1024], line_98[1022], line_97[1020], line_96[1018], line_95[1016], line_94[1014], line_93[1012], line_92[1010], line_91[1008], line_90[1006], line_89[1004], line_88[1002], line_87[1000], line_86[998], line_85[996], line_84[994], line_83[992], line_82[990], line_81[988], line_80[986], line_79[984], line_78[982], line_77[980], line_76[978], line_75[976], line_74[974], line_73[972], line_72[970], line_71[968], line_70[966], line_69[964], line_68[962], line_67[960], line_66[958], line_65[956], line_64[954], line_63[952], line_62[950], line_61[948], line_60[946], line_59[944], line_58[942], line_57[940], line_56[938], line_55[936], line_54[934], line_53[932], line_52[930], line_51[928], line_50[926], line_49[924], line_48[922], line_47[920], line_46[918], line_45[916], line_44[914], line_43[912], line_42[910], line_41[908], line_40[906], line_39[904], line_38[902], line_37[900], line_36[898], line_35[896], line_34[894], line_33[892], line_32[890], line_31[888], line_30[886], line_29[884], line_28[882], line_27[880], line_26[878], line_25[876], line_24[874], line_23[872], line_22[870], line_21[868], line_20[866], line_19[864], line_18[862], line_17[860], line_16[858], line_15[856], line_14[854], line_13[852], line_12[850], line_11[848], line_10[846], line_9[844], line_8[842], line_7[840], line_6[838], line_5[836], line_4[834], line_3[832], line_2[830], line_1[828], 29'b0};
assign col_1083 = {line_99[1025], line_98[1023], line_97[1021], line_96[1019], line_95[1017], line_94[1015], line_93[1013], line_92[1011], line_91[1009], line_90[1007], line_89[1005], line_88[1003], line_87[1001], line_86[999], line_85[997], line_84[995], line_83[993], line_82[991], line_81[989], line_80[987], line_79[985], line_78[983], line_77[981], line_76[979], line_75[977], line_74[975], line_73[973], line_72[971], line_71[969], line_70[967], line_69[965], line_68[963], line_67[961], line_66[959], line_65[957], line_64[955], line_63[953], line_62[951], line_61[949], line_60[947], line_59[945], line_58[943], line_57[941], line_56[939], line_55[937], line_54[935], line_53[933], line_52[931], line_51[929], line_50[927], line_49[925], line_48[923], line_47[921], line_46[919], line_45[917], line_44[915], line_43[913], line_42[911], line_41[909], line_40[907], line_39[905], line_38[903], line_37[901], line_36[899], line_35[897], line_34[895], line_33[893], line_32[891], line_31[889], line_30[887], line_29[885], line_28[883], line_27[881], line_26[879], line_25[877], line_24[875], line_23[873], line_22[871], line_21[869], line_20[867], line_19[865], line_18[863], line_17[861], line_16[859], line_15[857], line_14[855], line_13[853], line_12[851], line_11[849], line_10[847], line_9[845], line_8[843], line_7[841], line_6[839], line_5[837], line_4[835], line_3[833], line_2[831], line_1[829], 29'b0};
assign col_1084 = {line_98[1024], line_97[1022], line_96[1020], line_95[1018], line_94[1016], line_93[1014], line_92[1012], line_91[1010], line_90[1008], line_89[1006], line_88[1004], line_87[1002], line_86[1000], line_85[998], line_84[996], line_83[994], line_82[992], line_81[990], line_80[988], line_79[986], line_78[984], line_77[982], line_76[980], line_75[978], line_74[976], line_73[974], line_72[972], line_71[970], line_70[968], line_69[966], line_68[964], line_67[962], line_66[960], line_65[958], line_64[956], line_63[954], line_62[952], line_61[950], line_60[948], line_59[946], line_58[944], line_57[942], line_56[940], line_55[938], line_54[936], line_53[934], line_52[932], line_51[930], line_50[928], line_49[926], line_48[924], line_47[922], line_46[920], line_45[918], line_44[916], line_43[914], line_42[912], line_41[910], line_40[908], line_39[906], line_38[904], line_37[902], line_36[900], line_35[898], line_34[896], line_33[894], line_32[892], line_31[890], line_30[888], line_29[886], line_28[884], line_27[882], line_26[880], line_25[878], line_24[876], line_23[874], line_22[872], line_21[870], line_20[868], line_19[866], line_18[864], line_17[862], line_16[860], line_15[858], line_14[856], line_13[854], line_12[852], line_11[850], line_10[848], line_9[846], line_8[844], line_7[842], line_6[840], line_5[838], line_4[836], line_3[834], line_2[832], line_1[830], 30'b0};
assign col_1085 = {line_98[1025], line_97[1023], line_96[1021], line_95[1019], line_94[1017], line_93[1015], line_92[1013], line_91[1011], line_90[1009], line_89[1007], line_88[1005], line_87[1003], line_86[1001], line_85[999], line_84[997], line_83[995], line_82[993], line_81[991], line_80[989], line_79[987], line_78[985], line_77[983], line_76[981], line_75[979], line_74[977], line_73[975], line_72[973], line_71[971], line_70[969], line_69[967], line_68[965], line_67[963], line_66[961], line_65[959], line_64[957], line_63[955], line_62[953], line_61[951], line_60[949], line_59[947], line_58[945], line_57[943], line_56[941], line_55[939], line_54[937], line_53[935], line_52[933], line_51[931], line_50[929], line_49[927], line_48[925], line_47[923], line_46[921], line_45[919], line_44[917], line_43[915], line_42[913], line_41[911], line_40[909], line_39[907], line_38[905], line_37[903], line_36[901], line_35[899], line_34[897], line_33[895], line_32[893], line_31[891], line_30[889], line_29[887], line_28[885], line_27[883], line_26[881], line_25[879], line_24[877], line_23[875], line_22[873], line_21[871], line_20[869], line_19[867], line_18[865], line_17[863], line_16[861], line_15[859], line_14[857], line_13[855], line_12[853], line_11[851], line_10[849], line_9[847], line_8[845], line_7[843], line_6[841], line_5[839], line_4[837], line_3[835], line_2[833], line_1[831], 30'b0};
assign col_1086 = {line_97[1024], line_96[1022], line_95[1020], line_94[1018], line_93[1016], line_92[1014], line_91[1012], line_90[1010], line_89[1008], line_88[1006], line_87[1004], line_86[1002], line_85[1000], line_84[998], line_83[996], line_82[994], line_81[992], line_80[990], line_79[988], line_78[986], line_77[984], line_76[982], line_75[980], line_74[978], line_73[976], line_72[974], line_71[972], line_70[970], line_69[968], line_68[966], line_67[964], line_66[962], line_65[960], line_64[958], line_63[956], line_62[954], line_61[952], line_60[950], line_59[948], line_58[946], line_57[944], line_56[942], line_55[940], line_54[938], line_53[936], line_52[934], line_51[932], line_50[930], line_49[928], line_48[926], line_47[924], line_46[922], line_45[920], line_44[918], line_43[916], line_42[914], line_41[912], line_40[910], line_39[908], line_38[906], line_37[904], line_36[902], line_35[900], line_34[898], line_33[896], line_32[894], line_31[892], line_30[890], line_29[888], line_28[886], line_27[884], line_26[882], line_25[880], line_24[878], line_23[876], line_22[874], line_21[872], line_20[870], line_19[868], line_18[866], line_17[864], line_16[862], line_15[860], line_14[858], line_13[856], line_12[854], line_11[852], line_10[850], line_9[848], line_8[846], line_7[844], line_6[842], line_5[840], line_4[838], line_3[836], line_2[834], line_1[832], 31'b0};
assign col_1087 = {line_97[1025], line_96[1023], line_95[1021], line_94[1019], line_93[1017], line_92[1015], line_91[1013], line_90[1011], line_89[1009], line_88[1007], line_87[1005], line_86[1003], line_85[1001], line_84[999], line_83[997], line_82[995], line_81[993], line_80[991], line_79[989], line_78[987], line_77[985], line_76[983], line_75[981], line_74[979], line_73[977], line_72[975], line_71[973], line_70[971], line_69[969], line_68[967], line_67[965], line_66[963], line_65[961], line_64[959], line_63[957], line_62[955], line_61[953], line_60[951], line_59[949], line_58[947], line_57[945], line_56[943], line_55[941], line_54[939], line_53[937], line_52[935], line_51[933], line_50[931], line_49[929], line_48[927], line_47[925], line_46[923], line_45[921], line_44[919], line_43[917], line_42[915], line_41[913], line_40[911], line_39[909], line_38[907], line_37[905], line_36[903], line_35[901], line_34[899], line_33[897], line_32[895], line_31[893], line_30[891], line_29[889], line_28[887], line_27[885], line_26[883], line_25[881], line_24[879], line_23[877], line_22[875], line_21[873], line_20[871], line_19[869], line_18[867], line_17[865], line_16[863], line_15[861], line_14[859], line_13[857], line_12[855], line_11[853], line_10[851], line_9[849], line_8[847], line_7[845], line_6[843], line_5[841], line_4[839], line_3[837], line_2[835], line_1[833], 31'b0};
assign col_1088 = {line_96[1024], line_95[1022], line_94[1020], line_93[1018], line_92[1016], line_91[1014], line_90[1012], line_89[1010], line_88[1008], line_87[1006], line_86[1004], line_85[1002], line_84[1000], line_83[998], line_82[996], line_81[994], line_80[992], line_79[990], line_78[988], line_77[986], line_76[984], line_75[982], line_74[980], line_73[978], line_72[976], line_71[974], line_70[972], line_69[970], line_68[968], line_67[966], line_66[964], line_65[962], line_64[960], line_63[958], line_62[956], line_61[954], line_60[952], line_59[950], line_58[948], line_57[946], line_56[944], line_55[942], line_54[940], line_53[938], line_52[936], line_51[934], line_50[932], line_49[930], line_48[928], line_47[926], line_46[924], line_45[922], line_44[920], line_43[918], line_42[916], line_41[914], line_40[912], line_39[910], line_38[908], line_37[906], line_36[904], line_35[902], line_34[900], line_33[898], line_32[896], line_31[894], line_30[892], line_29[890], line_28[888], line_27[886], line_26[884], line_25[882], line_24[880], line_23[878], line_22[876], line_21[874], line_20[872], line_19[870], line_18[868], line_17[866], line_16[864], line_15[862], line_14[860], line_13[858], line_12[856], line_11[854], line_10[852], line_9[850], line_8[848], line_7[846], line_6[844], line_5[842], line_4[840], line_3[838], line_2[836], line_1[834], 32'b0};
assign col_1089 = {line_96[1025], line_95[1023], line_94[1021], line_93[1019], line_92[1017], line_91[1015], line_90[1013], line_89[1011], line_88[1009], line_87[1007], line_86[1005], line_85[1003], line_84[1001], line_83[999], line_82[997], line_81[995], line_80[993], line_79[991], line_78[989], line_77[987], line_76[985], line_75[983], line_74[981], line_73[979], line_72[977], line_71[975], line_70[973], line_69[971], line_68[969], line_67[967], line_66[965], line_65[963], line_64[961], line_63[959], line_62[957], line_61[955], line_60[953], line_59[951], line_58[949], line_57[947], line_56[945], line_55[943], line_54[941], line_53[939], line_52[937], line_51[935], line_50[933], line_49[931], line_48[929], line_47[927], line_46[925], line_45[923], line_44[921], line_43[919], line_42[917], line_41[915], line_40[913], line_39[911], line_38[909], line_37[907], line_36[905], line_35[903], line_34[901], line_33[899], line_32[897], line_31[895], line_30[893], line_29[891], line_28[889], line_27[887], line_26[885], line_25[883], line_24[881], line_23[879], line_22[877], line_21[875], line_20[873], line_19[871], line_18[869], line_17[867], line_16[865], line_15[863], line_14[861], line_13[859], line_12[857], line_11[855], line_10[853], line_9[851], line_8[849], line_7[847], line_6[845], line_5[843], line_4[841], line_3[839], line_2[837], line_1[835], 32'b0};
assign col_1090 = {line_95[1024], line_94[1022], line_93[1020], line_92[1018], line_91[1016], line_90[1014], line_89[1012], line_88[1010], line_87[1008], line_86[1006], line_85[1004], line_84[1002], line_83[1000], line_82[998], line_81[996], line_80[994], line_79[992], line_78[990], line_77[988], line_76[986], line_75[984], line_74[982], line_73[980], line_72[978], line_71[976], line_70[974], line_69[972], line_68[970], line_67[968], line_66[966], line_65[964], line_64[962], line_63[960], line_62[958], line_61[956], line_60[954], line_59[952], line_58[950], line_57[948], line_56[946], line_55[944], line_54[942], line_53[940], line_52[938], line_51[936], line_50[934], line_49[932], line_48[930], line_47[928], line_46[926], line_45[924], line_44[922], line_43[920], line_42[918], line_41[916], line_40[914], line_39[912], line_38[910], line_37[908], line_36[906], line_35[904], line_34[902], line_33[900], line_32[898], line_31[896], line_30[894], line_29[892], line_28[890], line_27[888], line_26[886], line_25[884], line_24[882], line_23[880], line_22[878], line_21[876], line_20[874], line_19[872], line_18[870], line_17[868], line_16[866], line_15[864], line_14[862], line_13[860], line_12[858], line_11[856], line_10[854], line_9[852], line_8[850], line_7[848], line_6[846], line_5[844], line_4[842], line_3[840], line_2[838], line_1[836], 33'b0};
assign col_1091 = {line_95[1025], line_94[1023], line_93[1021], line_92[1019], line_91[1017], line_90[1015], line_89[1013], line_88[1011], line_87[1009], line_86[1007], line_85[1005], line_84[1003], line_83[1001], line_82[999], line_81[997], line_80[995], line_79[993], line_78[991], line_77[989], line_76[987], line_75[985], line_74[983], line_73[981], line_72[979], line_71[977], line_70[975], line_69[973], line_68[971], line_67[969], line_66[967], line_65[965], line_64[963], line_63[961], line_62[959], line_61[957], line_60[955], line_59[953], line_58[951], line_57[949], line_56[947], line_55[945], line_54[943], line_53[941], line_52[939], line_51[937], line_50[935], line_49[933], line_48[931], line_47[929], line_46[927], line_45[925], line_44[923], line_43[921], line_42[919], line_41[917], line_40[915], line_39[913], line_38[911], line_37[909], line_36[907], line_35[905], line_34[903], line_33[901], line_32[899], line_31[897], line_30[895], line_29[893], line_28[891], line_27[889], line_26[887], line_25[885], line_24[883], line_23[881], line_22[879], line_21[877], line_20[875], line_19[873], line_18[871], line_17[869], line_16[867], line_15[865], line_14[863], line_13[861], line_12[859], line_11[857], line_10[855], line_9[853], line_8[851], line_7[849], line_6[847], line_5[845], line_4[843], line_3[841], line_2[839], line_1[837], 33'b0};
assign col_1092 = {line_94[1024], line_93[1022], line_92[1020], line_91[1018], line_90[1016], line_89[1014], line_88[1012], line_87[1010], line_86[1008], line_85[1006], line_84[1004], line_83[1002], line_82[1000], line_81[998], line_80[996], line_79[994], line_78[992], line_77[990], line_76[988], line_75[986], line_74[984], line_73[982], line_72[980], line_71[978], line_70[976], line_69[974], line_68[972], line_67[970], line_66[968], line_65[966], line_64[964], line_63[962], line_62[960], line_61[958], line_60[956], line_59[954], line_58[952], line_57[950], line_56[948], line_55[946], line_54[944], line_53[942], line_52[940], line_51[938], line_50[936], line_49[934], line_48[932], line_47[930], line_46[928], line_45[926], line_44[924], line_43[922], line_42[920], line_41[918], line_40[916], line_39[914], line_38[912], line_37[910], line_36[908], line_35[906], line_34[904], line_33[902], line_32[900], line_31[898], line_30[896], line_29[894], line_28[892], line_27[890], line_26[888], line_25[886], line_24[884], line_23[882], line_22[880], line_21[878], line_20[876], line_19[874], line_18[872], line_17[870], line_16[868], line_15[866], line_14[864], line_13[862], line_12[860], line_11[858], line_10[856], line_9[854], line_8[852], line_7[850], line_6[848], line_5[846], line_4[844], line_3[842], line_2[840], line_1[838], 34'b0};
assign col_1093 = {line_94[1025], line_93[1023], line_92[1021], line_91[1019], line_90[1017], line_89[1015], line_88[1013], line_87[1011], line_86[1009], line_85[1007], line_84[1005], line_83[1003], line_82[1001], line_81[999], line_80[997], line_79[995], line_78[993], line_77[991], line_76[989], line_75[987], line_74[985], line_73[983], line_72[981], line_71[979], line_70[977], line_69[975], line_68[973], line_67[971], line_66[969], line_65[967], line_64[965], line_63[963], line_62[961], line_61[959], line_60[957], line_59[955], line_58[953], line_57[951], line_56[949], line_55[947], line_54[945], line_53[943], line_52[941], line_51[939], line_50[937], line_49[935], line_48[933], line_47[931], line_46[929], line_45[927], line_44[925], line_43[923], line_42[921], line_41[919], line_40[917], line_39[915], line_38[913], line_37[911], line_36[909], line_35[907], line_34[905], line_33[903], line_32[901], line_31[899], line_30[897], line_29[895], line_28[893], line_27[891], line_26[889], line_25[887], line_24[885], line_23[883], line_22[881], line_21[879], line_20[877], line_19[875], line_18[873], line_17[871], line_16[869], line_15[867], line_14[865], line_13[863], line_12[861], line_11[859], line_10[857], line_9[855], line_8[853], line_7[851], line_6[849], line_5[847], line_4[845], line_3[843], line_2[841], line_1[839], 34'b0};
assign col_1094 = {line_93[1024], line_92[1022], line_91[1020], line_90[1018], line_89[1016], line_88[1014], line_87[1012], line_86[1010], line_85[1008], line_84[1006], line_83[1004], line_82[1002], line_81[1000], line_80[998], line_79[996], line_78[994], line_77[992], line_76[990], line_75[988], line_74[986], line_73[984], line_72[982], line_71[980], line_70[978], line_69[976], line_68[974], line_67[972], line_66[970], line_65[968], line_64[966], line_63[964], line_62[962], line_61[960], line_60[958], line_59[956], line_58[954], line_57[952], line_56[950], line_55[948], line_54[946], line_53[944], line_52[942], line_51[940], line_50[938], line_49[936], line_48[934], line_47[932], line_46[930], line_45[928], line_44[926], line_43[924], line_42[922], line_41[920], line_40[918], line_39[916], line_38[914], line_37[912], line_36[910], line_35[908], line_34[906], line_33[904], line_32[902], line_31[900], line_30[898], line_29[896], line_28[894], line_27[892], line_26[890], line_25[888], line_24[886], line_23[884], line_22[882], line_21[880], line_20[878], line_19[876], line_18[874], line_17[872], line_16[870], line_15[868], line_14[866], line_13[864], line_12[862], line_11[860], line_10[858], line_9[856], line_8[854], line_7[852], line_6[850], line_5[848], line_4[846], line_3[844], line_2[842], line_1[840], 35'b0};
assign col_1095 = {line_93[1025], line_92[1023], line_91[1021], line_90[1019], line_89[1017], line_88[1015], line_87[1013], line_86[1011], line_85[1009], line_84[1007], line_83[1005], line_82[1003], line_81[1001], line_80[999], line_79[997], line_78[995], line_77[993], line_76[991], line_75[989], line_74[987], line_73[985], line_72[983], line_71[981], line_70[979], line_69[977], line_68[975], line_67[973], line_66[971], line_65[969], line_64[967], line_63[965], line_62[963], line_61[961], line_60[959], line_59[957], line_58[955], line_57[953], line_56[951], line_55[949], line_54[947], line_53[945], line_52[943], line_51[941], line_50[939], line_49[937], line_48[935], line_47[933], line_46[931], line_45[929], line_44[927], line_43[925], line_42[923], line_41[921], line_40[919], line_39[917], line_38[915], line_37[913], line_36[911], line_35[909], line_34[907], line_33[905], line_32[903], line_31[901], line_30[899], line_29[897], line_28[895], line_27[893], line_26[891], line_25[889], line_24[887], line_23[885], line_22[883], line_21[881], line_20[879], line_19[877], line_18[875], line_17[873], line_16[871], line_15[869], line_14[867], line_13[865], line_12[863], line_11[861], line_10[859], line_9[857], line_8[855], line_7[853], line_6[851], line_5[849], line_4[847], line_3[845], line_2[843], line_1[841], 35'b0};
assign col_1096 = {line_92[1024], line_91[1022], line_90[1020], line_89[1018], line_88[1016], line_87[1014], line_86[1012], line_85[1010], line_84[1008], line_83[1006], line_82[1004], line_81[1002], line_80[1000], line_79[998], line_78[996], line_77[994], line_76[992], line_75[990], line_74[988], line_73[986], line_72[984], line_71[982], line_70[980], line_69[978], line_68[976], line_67[974], line_66[972], line_65[970], line_64[968], line_63[966], line_62[964], line_61[962], line_60[960], line_59[958], line_58[956], line_57[954], line_56[952], line_55[950], line_54[948], line_53[946], line_52[944], line_51[942], line_50[940], line_49[938], line_48[936], line_47[934], line_46[932], line_45[930], line_44[928], line_43[926], line_42[924], line_41[922], line_40[920], line_39[918], line_38[916], line_37[914], line_36[912], line_35[910], line_34[908], line_33[906], line_32[904], line_31[902], line_30[900], line_29[898], line_28[896], line_27[894], line_26[892], line_25[890], line_24[888], line_23[886], line_22[884], line_21[882], line_20[880], line_19[878], line_18[876], line_17[874], line_16[872], line_15[870], line_14[868], line_13[866], line_12[864], line_11[862], line_10[860], line_9[858], line_8[856], line_7[854], line_6[852], line_5[850], line_4[848], line_3[846], line_2[844], line_1[842], 36'b0};
assign col_1097 = {line_92[1025], line_91[1023], line_90[1021], line_89[1019], line_88[1017], line_87[1015], line_86[1013], line_85[1011], line_84[1009], line_83[1007], line_82[1005], line_81[1003], line_80[1001], line_79[999], line_78[997], line_77[995], line_76[993], line_75[991], line_74[989], line_73[987], line_72[985], line_71[983], line_70[981], line_69[979], line_68[977], line_67[975], line_66[973], line_65[971], line_64[969], line_63[967], line_62[965], line_61[963], line_60[961], line_59[959], line_58[957], line_57[955], line_56[953], line_55[951], line_54[949], line_53[947], line_52[945], line_51[943], line_50[941], line_49[939], line_48[937], line_47[935], line_46[933], line_45[931], line_44[929], line_43[927], line_42[925], line_41[923], line_40[921], line_39[919], line_38[917], line_37[915], line_36[913], line_35[911], line_34[909], line_33[907], line_32[905], line_31[903], line_30[901], line_29[899], line_28[897], line_27[895], line_26[893], line_25[891], line_24[889], line_23[887], line_22[885], line_21[883], line_20[881], line_19[879], line_18[877], line_17[875], line_16[873], line_15[871], line_14[869], line_13[867], line_12[865], line_11[863], line_10[861], line_9[859], line_8[857], line_7[855], line_6[853], line_5[851], line_4[849], line_3[847], line_2[845], line_1[843], 36'b0};
assign col_1098 = {line_91[1024], line_90[1022], line_89[1020], line_88[1018], line_87[1016], line_86[1014], line_85[1012], line_84[1010], line_83[1008], line_82[1006], line_81[1004], line_80[1002], line_79[1000], line_78[998], line_77[996], line_76[994], line_75[992], line_74[990], line_73[988], line_72[986], line_71[984], line_70[982], line_69[980], line_68[978], line_67[976], line_66[974], line_65[972], line_64[970], line_63[968], line_62[966], line_61[964], line_60[962], line_59[960], line_58[958], line_57[956], line_56[954], line_55[952], line_54[950], line_53[948], line_52[946], line_51[944], line_50[942], line_49[940], line_48[938], line_47[936], line_46[934], line_45[932], line_44[930], line_43[928], line_42[926], line_41[924], line_40[922], line_39[920], line_38[918], line_37[916], line_36[914], line_35[912], line_34[910], line_33[908], line_32[906], line_31[904], line_30[902], line_29[900], line_28[898], line_27[896], line_26[894], line_25[892], line_24[890], line_23[888], line_22[886], line_21[884], line_20[882], line_19[880], line_18[878], line_17[876], line_16[874], line_15[872], line_14[870], line_13[868], line_12[866], line_11[864], line_10[862], line_9[860], line_8[858], line_7[856], line_6[854], line_5[852], line_4[850], line_3[848], line_2[846], line_1[844], 37'b0};
assign col_1099 = {line_91[1025], line_90[1023], line_89[1021], line_88[1019], line_87[1017], line_86[1015], line_85[1013], line_84[1011], line_83[1009], line_82[1007], line_81[1005], line_80[1003], line_79[1001], line_78[999], line_77[997], line_76[995], line_75[993], line_74[991], line_73[989], line_72[987], line_71[985], line_70[983], line_69[981], line_68[979], line_67[977], line_66[975], line_65[973], line_64[971], line_63[969], line_62[967], line_61[965], line_60[963], line_59[961], line_58[959], line_57[957], line_56[955], line_55[953], line_54[951], line_53[949], line_52[947], line_51[945], line_50[943], line_49[941], line_48[939], line_47[937], line_46[935], line_45[933], line_44[931], line_43[929], line_42[927], line_41[925], line_40[923], line_39[921], line_38[919], line_37[917], line_36[915], line_35[913], line_34[911], line_33[909], line_32[907], line_31[905], line_30[903], line_29[901], line_28[899], line_27[897], line_26[895], line_25[893], line_24[891], line_23[889], line_22[887], line_21[885], line_20[883], line_19[881], line_18[879], line_17[877], line_16[875], line_15[873], line_14[871], line_13[869], line_12[867], line_11[865], line_10[863], line_9[861], line_8[859], line_7[857], line_6[855], line_5[853], line_4[851], line_3[849], line_2[847], line_1[845], 37'b0};
assign col_1100 = {line_90[1024], line_89[1022], line_88[1020], line_87[1018], line_86[1016], line_85[1014], line_84[1012], line_83[1010], line_82[1008], line_81[1006], line_80[1004], line_79[1002], line_78[1000], line_77[998], line_76[996], line_75[994], line_74[992], line_73[990], line_72[988], line_71[986], line_70[984], line_69[982], line_68[980], line_67[978], line_66[976], line_65[974], line_64[972], line_63[970], line_62[968], line_61[966], line_60[964], line_59[962], line_58[960], line_57[958], line_56[956], line_55[954], line_54[952], line_53[950], line_52[948], line_51[946], line_50[944], line_49[942], line_48[940], line_47[938], line_46[936], line_45[934], line_44[932], line_43[930], line_42[928], line_41[926], line_40[924], line_39[922], line_38[920], line_37[918], line_36[916], line_35[914], line_34[912], line_33[910], line_32[908], line_31[906], line_30[904], line_29[902], line_28[900], line_27[898], line_26[896], line_25[894], line_24[892], line_23[890], line_22[888], line_21[886], line_20[884], line_19[882], line_18[880], line_17[878], line_16[876], line_15[874], line_14[872], line_13[870], line_12[868], line_11[866], line_10[864], line_9[862], line_8[860], line_7[858], line_6[856], line_5[854], line_4[852], line_3[850], line_2[848], line_1[846], 38'b0};
assign col_1101 = {line_90[1025], line_89[1023], line_88[1021], line_87[1019], line_86[1017], line_85[1015], line_84[1013], line_83[1011], line_82[1009], line_81[1007], line_80[1005], line_79[1003], line_78[1001], line_77[999], line_76[997], line_75[995], line_74[993], line_73[991], line_72[989], line_71[987], line_70[985], line_69[983], line_68[981], line_67[979], line_66[977], line_65[975], line_64[973], line_63[971], line_62[969], line_61[967], line_60[965], line_59[963], line_58[961], line_57[959], line_56[957], line_55[955], line_54[953], line_53[951], line_52[949], line_51[947], line_50[945], line_49[943], line_48[941], line_47[939], line_46[937], line_45[935], line_44[933], line_43[931], line_42[929], line_41[927], line_40[925], line_39[923], line_38[921], line_37[919], line_36[917], line_35[915], line_34[913], line_33[911], line_32[909], line_31[907], line_30[905], line_29[903], line_28[901], line_27[899], line_26[897], line_25[895], line_24[893], line_23[891], line_22[889], line_21[887], line_20[885], line_19[883], line_18[881], line_17[879], line_16[877], line_15[875], line_14[873], line_13[871], line_12[869], line_11[867], line_10[865], line_9[863], line_8[861], line_7[859], line_6[857], line_5[855], line_4[853], line_3[851], line_2[849], line_1[847], 38'b0};
assign col_1102 = {line_89[1024], line_88[1022], line_87[1020], line_86[1018], line_85[1016], line_84[1014], line_83[1012], line_82[1010], line_81[1008], line_80[1006], line_79[1004], line_78[1002], line_77[1000], line_76[998], line_75[996], line_74[994], line_73[992], line_72[990], line_71[988], line_70[986], line_69[984], line_68[982], line_67[980], line_66[978], line_65[976], line_64[974], line_63[972], line_62[970], line_61[968], line_60[966], line_59[964], line_58[962], line_57[960], line_56[958], line_55[956], line_54[954], line_53[952], line_52[950], line_51[948], line_50[946], line_49[944], line_48[942], line_47[940], line_46[938], line_45[936], line_44[934], line_43[932], line_42[930], line_41[928], line_40[926], line_39[924], line_38[922], line_37[920], line_36[918], line_35[916], line_34[914], line_33[912], line_32[910], line_31[908], line_30[906], line_29[904], line_28[902], line_27[900], line_26[898], line_25[896], line_24[894], line_23[892], line_22[890], line_21[888], line_20[886], line_19[884], line_18[882], line_17[880], line_16[878], line_15[876], line_14[874], line_13[872], line_12[870], line_11[868], line_10[866], line_9[864], line_8[862], line_7[860], line_6[858], line_5[856], line_4[854], line_3[852], line_2[850], line_1[848], 39'b0};
assign col_1103 = {line_89[1025], line_88[1023], line_87[1021], line_86[1019], line_85[1017], line_84[1015], line_83[1013], line_82[1011], line_81[1009], line_80[1007], line_79[1005], line_78[1003], line_77[1001], line_76[999], line_75[997], line_74[995], line_73[993], line_72[991], line_71[989], line_70[987], line_69[985], line_68[983], line_67[981], line_66[979], line_65[977], line_64[975], line_63[973], line_62[971], line_61[969], line_60[967], line_59[965], line_58[963], line_57[961], line_56[959], line_55[957], line_54[955], line_53[953], line_52[951], line_51[949], line_50[947], line_49[945], line_48[943], line_47[941], line_46[939], line_45[937], line_44[935], line_43[933], line_42[931], line_41[929], line_40[927], line_39[925], line_38[923], line_37[921], line_36[919], line_35[917], line_34[915], line_33[913], line_32[911], line_31[909], line_30[907], line_29[905], line_28[903], line_27[901], line_26[899], line_25[897], line_24[895], line_23[893], line_22[891], line_21[889], line_20[887], line_19[885], line_18[883], line_17[881], line_16[879], line_15[877], line_14[875], line_13[873], line_12[871], line_11[869], line_10[867], line_9[865], line_8[863], line_7[861], line_6[859], line_5[857], line_4[855], line_3[853], line_2[851], line_1[849], 39'b0};
assign col_1104 = {line_88[1024], line_87[1022], line_86[1020], line_85[1018], line_84[1016], line_83[1014], line_82[1012], line_81[1010], line_80[1008], line_79[1006], line_78[1004], line_77[1002], line_76[1000], line_75[998], line_74[996], line_73[994], line_72[992], line_71[990], line_70[988], line_69[986], line_68[984], line_67[982], line_66[980], line_65[978], line_64[976], line_63[974], line_62[972], line_61[970], line_60[968], line_59[966], line_58[964], line_57[962], line_56[960], line_55[958], line_54[956], line_53[954], line_52[952], line_51[950], line_50[948], line_49[946], line_48[944], line_47[942], line_46[940], line_45[938], line_44[936], line_43[934], line_42[932], line_41[930], line_40[928], line_39[926], line_38[924], line_37[922], line_36[920], line_35[918], line_34[916], line_33[914], line_32[912], line_31[910], line_30[908], line_29[906], line_28[904], line_27[902], line_26[900], line_25[898], line_24[896], line_23[894], line_22[892], line_21[890], line_20[888], line_19[886], line_18[884], line_17[882], line_16[880], line_15[878], line_14[876], line_13[874], line_12[872], line_11[870], line_10[868], line_9[866], line_8[864], line_7[862], line_6[860], line_5[858], line_4[856], line_3[854], line_2[852], line_1[850], 40'b0};
assign col_1105 = {line_88[1025], line_87[1023], line_86[1021], line_85[1019], line_84[1017], line_83[1015], line_82[1013], line_81[1011], line_80[1009], line_79[1007], line_78[1005], line_77[1003], line_76[1001], line_75[999], line_74[997], line_73[995], line_72[993], line_71[991], line_70[989], line_69[987], line_68[985], line_67[983], line_66[981], line_65[979], line_64[977], line_63[975], line_62[973], line_61[971], line_60[969], line_59[967], line_58[965], line_57[963], line_56[961], line_55[959], line_54[957], line_53[955], line_52[953], line_51[951], line_50[949], line_49[947], line_48[945], line_47[943], line_46[941], line_45[939], line_44[937], line_43[935], line_42[933], line_41[931], line_40[929], line_39[927], line_38[925], line_37[923], line_36[921], line_35[919], line_34[917], line_33[915], line_32[913], line_31[911], line_30[909], line_29[907], line_28[905], line_27[903], line_26[901], line_25[899], line_24[897], line_23[895], line_22[893], line_21[891], line_20[889], line_19[887], line_18[885], line_17[883], line_16[881], line_15[879], line_14[877], line_13[875], line_12[873], line_11[871], line_10[869], line_9[867], line_8[865], line_7[863], line_6[861], line_5[859], line_4[857], line_3[855], line_2[853], line_1[851], 40'b0};
assign col_1106 = {line_87[1024], line_86[1022], line_85[1020], line_84[1018], line_83[1016], line_82[1014], line_81[1012], line_80[1010], line_79[1008], line_78[1006], line_77[1004], line_76[1002], line_75[1000], line_74[998], line_73[996], line_72[994], line_71[992], line_70[990], line_69[988], line_68[986], line_67[984], line_66[982], line_65[980], line_64[978], line_63[976], line_62[974], line_61[972], line_60[970], line_59[968], line_58[966], line_57[964], line_56[962], line_55[960], line_54[958], line_53[956], line_52[954], line_51[952], line_50[950], line_49[948], line_48[946], line_47[944], line_46[942], line_45[940], line_44[938], line_43[936], line_42[934], line_41[932], line_40[930], line_39[928], line_38[926], line_37[924], line_36[922], line_35[920], line_34[918], line_33[916], line_32[914], line_31[912], line_30[910], line_29[908], line_28[906], line_27[904], line_26[902], line_25[900], line_24[898], line_23[896], line_22[894], line_21[892], line_20[890], line_19[888], line_18[886], line_17[884], line_16[882], line_15[880], line_14[878], line_13[876], line_12[874], line_11[872], line_10[870], line_9[868], line_8[866], line_7[864], line_6[862], line_5[860], line_4[858], line_3[856], line_2[854], line_1[852], 41'b0};
assign col_1107 = {line_87[1025], line_86[1023], line_85[1021], line_84[1019], line_83[1017], line_82[1015], line_81[1013], line_80[1011], line_79[1009], line_78[1007], line_77[1005], line_76[1003], line_75[1001], line_74[999], line_73[997], line_72[995], line_71[993], line_70[991], line_69[989], line_68[987], line_67[985], line_66[983], line_65[981], line_64[979], line_63[977], line_62[975], line_61[973], line_60[971], line_59[969], line_58[967], line_57[965], line_56[963], line_55[961], line_54[959], line_53[957], line_52[955], line_51[953], line_50[951], line_49[949], line_48[947], line_47[945], line_46[943], line_45[941], line_44[939], line_43[937], line_42[935], line_41[933], line_40[931], line_39[929], line_38[927], line_37[925], line_36[923], line_35[921], line_34[919], line_33[917], line_32[915], line_31[913], line_30[911], line_29[909], line_28[907], line_27[905], line_26[903], line_25[901], line_24[899], line_23[897], line_22[895], line_21[893], line_20[891], line_19[889], line_18[887], line_17[885], line_16[883], line_15[881], line_14[879], line_13[877], line_12[875], line_11[873], line_10[871], line_9[869], line_8[867], line_7[865], line_6[863], line_5[861], line_4[859], line_3[857], line_2[855], line_1[853], 41'b0};
assign col_1108 = {line_86[1024], line_85[1022], line_84[1020], line_83[1018], line_82[1016], line_81[1014], line_80[1012], line_79[1010], line_78[1008], line_77[1006], line_76[1004], line_75[1002], line_74[1000], line_73[998], line_72[996], line_71[994], line_70[992], line_69[990], line_68[988], line_67[986], line_66[984], line_65[982], line_64[980], line_63[978], line_62[976], line_61[974], line_60[972], line_59[970], line_58[968], line_57[966], line_56[964], line_55[962], line_54[960], line_53[958], line_52[956], line_51[954], line_50[952], line_49[950], line_48[948], line_47[946], line_46[944], line_45[942], line_44[940], line_43[938], line_42[936], line_41[934], line_40[932], line_39[930], line_38[928], line_37[926], line_36[924], line_35[922], line_34[920], line_33[918], line_32[916], line_31[914], line_30[912], line_29[910], line_28[908], line_27[906], line_26[904], line_25[902], line_24[900], line_23[898], line_22[896], line_21[894], line_20[892], line_19[890], line_18[888], line_17[886], line_16[884], line_15[882], line_14[880], line_13[878], line_12[876], line_11[874], line_10[872], line_9[870], line_8[868], line_7[866], line_6[864], line_5[862], line_4[860], line_3[858], line_2[856], line_1[854], 42'b0};
assign col_1109 = {line_86[1025], line_85[1023], line_84[1021], line_83[1019], line_82[1017], line_81[1015], line_80[1013], line_79[1011], line_78[1009], line_77[1007], line_76[1005], line_75[1003], line_74[1001], line_73[999], line_72[997], line_71[995], line_70[993], line_69[991], line_68[989], line_67[987], line_66[985], line_65[983], line_64[981], line_63[979], line_62[977], line_61[975], line_60[973], line_59[971], line_58[969], line_57[967], line_56[965], line_55[963], line_54[961], line_53[959], line_52[957], line_51[955], line_50[953], line_49[951], line_48[949], line_47[947], line_46[945], line_45[943], line_44[941], line_43[939], line_42[937], line_41[935], line_40[933], line_39[931], line_38[929], line_37[927], line_36[925], line_35[923], line_34[921], line_33[919], line_32[917], line_31[915], line_30[913], line_29[911], line_28[909], line_27[907], line_26[905], line_25[903], line_24[901], line_23[899], line_22[897], line_21[895], line_20[893], line_19[891], line_18[889], line_17[887], line_16[885], line_15[883], line_14[881], line_13[879], line_12[877], line_11[875], line_10[873], line_9[871], line_8[869], line_7[867], line_6[865], line_5[863], line_4[861], line_3[859], line_2[857], line_1[855], 42'b0};
assign col_1110 = {line_85[1024], line_84[1022], line_83[1020], line_82[1018], line_81[1016], line_80[1014], line_79[1012], line_78[1010], line_77[1008], line_76[1006], line_75[1004], line_74[1002], line_73[1000], line_72[998], line_71[996], line_70[994], line_69[992], line_68[990], line_67[988], line_66[986], line_65[984], line_64[982], line_63[980], line_62[978], line_61[976], line_60[974], line_59[972], line_58[970], line_57[968], line_56[966], line_55[964], line_54[962], line_53[960], line_52[958], line_51[956], line_50[954], line_49[952], line_48[950], line_47[948], line_46[946], line_45[944], line_44[942], line_43[940], line_42[938], line_41[936], line_40[934], line_39[932], line_38[930], line_37[928], line_36[926], line_35[924], line_34[922], line_33[920], line_32[918], line_31[916], line_30[914], line_29[912], line_28[910], line_27[908], line_26[906], line_25[904], line_24[902], line_23[900], line_22[898], line_21[896], line_20[894], line_19[892], line_18[890], line_17[888], line_16[886], line_15[884], line_14[882], line_13[880], line_12[878], line_11[876], line_10[874], line_9[872], line_8[870], line_7[868], line_6[866], line_5[864], line_4[862], line_3[860], line_2[858], line_1[856], 43'b0};
assign col_1111 = {line_85[1025], line_84[1023], line_83[1021], line_82[1019], line_81[1017], line_80[1015], line_79[1013], line_78[1011], line_77[1009], line_76[1007], line_75[1005], line_74[1003], line_73[1001], line_72[999], line_71[997], line_70[995], line_69[993], line_68[991], line_67[989], line_66[987], line_65[985], line_64[983], line_63[981], line_62[979], line_61[977], line_60[975], line_59[973], line_58[971], line_57[969], line_56[967], line_55[965], line_54[963], line_53[961], line_52[959], line_51[957], line_50[955], line_49[953], line_48[951], line_47[949], line_46[947], line_45[945], line_44[943], line_43[941], line_42[939], line_41[937], line_40[935], line_39[933], line_38[931], line_37[929], line_36[927], line_35[925], line_34[923], line_33[921], line_32[919], line_31[917], line_30[915], line_29[913], line_28[911], line_27[909], line_26[907], line_25[905], line_24[903], line_23[901], line_22[899], line_21[897], line_20[895], line_19[893], line_18[891], line_17[889], line_16[887], line_15[885], line_14[883], line_13[881], line_12[879], line_11[877], line_10[875], line_9[873], line_8[871], line_7[869], line_6[867], line_5[865], line_4[863], line_3[861], line_2[859], line_1[857], 43'b0};
assign col_1112 = {line_84[1024], line_83[1022], line_82[1020], line_81[1018], line_80[1016], line_79[1014], line_78[1012], line_77[1010], line_76[1008], line_75[1006], line_74[1004], line_73[1002], line_72[1000], line_71[998], line_70[996], line_69[994], line_68[992], line_67[990], line_66[988], line_65[986], line_64[984], line_63[982], line_62[980], line_61[978], line_60[976], line_59[974], line_58[972], line_57[970], line_56[968], line_55[966], line_54[964], line_53[962], line_52[960], line_51[958], line_50[956], line_49[954], line_48[952], line_47[950], line_46[948], line_45[946], line_44[944], line_43[942], line_42[940], line_41[938], line_40[936], line_39[934], line_38[932], line_37[930], line_36[928], line_35[926], line_34[924], line_33[922], line_32[920], line_31[918], line_30[916], line_29[914], line_28[912], line_27[910], line_26[908], line_25[906], line_24[904], line_23[902], line_22[900], line_21[898], line_20[896], line_19[894], line_18[892], line_17[890], line_16[888], line_15[886], line_14[884], line_13[882], line_12[880], line_11[878], line_10[876], line_9[874], line_8[872], line_7[870], line_6[868], line_5[866], line_4[864], line_3[862], line_2[860], line_1[858], 44'b0};
assign col_1113 = {line_84[1025], line_83[1023], line_82[1021], line_81[1019], line_80[1017], line_79[1015], line_78[1013], line_77[1011], line_76[1009], line_75[1007], line_74[1005], line_73[1003], line_72[1001], line_71[999], line_70[997], line_69[995], line_68[993], line_67[991], line_66[989], line_65[987], line_64[985], line_63[983], line_62[981], line_61[979], line_60[977], line_59[975], line_58[973], line_57[971], line_56[969], line_55[967], line_54[965], line_53[963], line_52[961], line_51[959], line_50[957], line_49[955], line_48[953], line_47[951], line_46[949], line_45[947], line_44[945], line_43[943], line_42[941], line_41[939], line_40[937], line_39[935], line_38[933], line_37[931], line_36[929], line_35[927], line_34[925], line_33[923], line_32[921], line_31[919], line_30[917], line_29[915], line_28[913], line_27[911], line_26[909], line_25[907], line_24[905], line_23[903], line_22[901], line_21[899], line_20[897], line_19[895], line_18[893], line_17[891], line_16[889], line_15[887], line_14[885], line_13[883], line_12[881], line_11[879], line_10[877], line_9[875], line_8[873], line_7[871], line_6[869], line_5[867], line_4[865], line_3[863], line_2[861], line_1[859], 44'b0};
assign col_1114 = {line_83[1024], line_82[1022], line_81[1020], line_80[1018], line_79[1016], line_78[1014], line_77[1012], line_76[1010], line_75[1008], line_74[1006], line_73[1004], line_72[1002], line_71[1000], line_70[998], line_69[996], line_68[994], line_67[992], line_66[990], line_65[988], line_64[986], line_63[984], line_62[982], line_61[980], line_60[978], line_59[976], line_58[974], line_57[972], line_56[970], line_55[968], line_54[966], line_53[964], line_52[962], line_51[960], line_50[958], line_49[956], line_48[954], line_47[952], line_46[950], line_45[948], line_44[946], line_43[944], line_42[942], line_41[940], line_40[938], line_39[936], line_38[934], line_37[932], line_36[930], line_35[928], line_34[926], line_33[924], line_32[922], line_31[920], line_30[918], line_29[916], line_28[914], line_27[912], line_26[910], line_25[908], line_24[906], line_23[904], line_22[902], line_21[900], line_20[898], line_19[896], line_18[894], line_17[892], line_16[890], line_15[888], line_14[886], line_13[884], line_12[882], line_11[880], line_10[878], line_9[876], line_8[874], line_7[872], line_6[870], line_5[868], line_4[866], line_3[864], line_2[862], line_1[860], 45'b0};
assign col_1115 = {line_83[1025], line_82[1023], line_81[1021], line_80[1019], line_79[1017], line_78[1015], line_77[1013], line_76[1011], line_75[1009], line_74[1007], line_73[1005], line_72[1003], line_71[1001], line_70[999], line_69[997], line_68[995], line_67[993], line_66[991], line_65[989], line_64[987], line_63[985], line_62[983], line_61[981], line_60[979], line_59[977], line_58[975], line_57[973], line_56[971], line_55[969], line_54[967], line_53[965], line_52[963], line_51[961], line_50[959], line_49[957], line_48[955], line_47[953], line_46[951], line_45[949], line_44[947], line_43[945], line_42[943], line_41[941], line_40[939], line_39[937], line_38[935], line_37[933], line_36[931], line_35[929], line_34[927], line_33[925], line_32[923], line_31[921], line_30[919], line_29[917], line_28[915], line_27[913], line_26[911], line_25[909], line_24[907], line_23[905], line_22[903], line_21[901], line_20[899], line_19[897], line_18[895], line_17[893], line_16[891], line_15[889], line_14[887], line_13[885], line_12[883], line_11[881], line_10[879], line_9[877], line_8[875], line_7[873], line_6[871], line_5[869], line_4[867], line_3[865], line_2[863], line_1[861], 45'b0};
assign col_1116 = {line_82[1024], line_81[1022], line_80[1020], line_79[1018], line_78[1016], line_77[1014], line_76[1012], line_75[1010], line_74[1008], line_73[1006], line_72[1004], line_71[1002], line_70[1000], line_69[998], line_68[996], line_67[994], line_66[992], line_65[990], line_64[988], line_63[986], line_62[984], line_61[982], line_60[980], line_59[978], line_58[976], line_57[974], line_56[972], line_55[970], line_54[968], line_53[966], line_52[964], line_51[962], line_50[960], line_49[958], line_48[956], line_47[954], line_46[952], line_45[950], line_44[948], line_43[946], line_42[944], line_41[942], line_40[940], line_39[938], line_38[936], line_37[934], line_36[932], line_35[930], line_34[928], line_33[926], line_32[924], line_31[922], line_30[920], line_29[918], line_28[916], line_27[914], line_26[912], line_25[910], line_24[908], line_23[906], line_22[904], line_21[902], line_20[900], line_19[898], line_18[896], line_17[894], line_16[892], line_15[890], line_14[888], line_13[886], line_12[884], line_11[882], line_10[880], line_9[878], line_8[876], line_7[874], line_6[872], line_5[870], line_4[868], line_3[866], line_2[864], line_1[862], 46'b0};
assign col_1117 = {line_82[1025], line_81[1023], line_80[1021], line_79[1019], line_78[1017], line_77[1015], line_76[1013], line_75[1011], line_74[1009], line_73[1007], line_72[1005], line_71[1003], line_70[1001], line_69[999], line_68[997], line_67[995], line_66[993], line_65[991], line_64[989], line_63[987], line_62[985], line_61[983], line_60[981], line_59[979], line_58[977], line_57[975], line_56[973], line_55[971], line_54[969], line_53[967], line_52[965], line_51[963], line_50[961], line_49[959], line_48[957], line_47[955], line_46[953], line_45[951], line_44[949], line_43[947], line_42[945], line_41[943], line_40[941], line_39[939], line_38[937], line_37[935], line_36[933], line_35[931], line_34[929], line_33[927], line_32[925], line_31[923], line_30[921], line_29[919], line_28[917], line_27[915], line_26[913], line_25[911], line_24[909], line_23[907], line_22[905], line_21[903], line_20[901], line_19[899], line_18[897], line_17[895], line_16[893], line_15[891], line_14[889], line_13[887], line_12[885], line_11[883], line_10[881], line_9[879], line_8[877], line_7[875], line_6[873], line_5[871], line_4[869], line_3[867], line_2[865], line_1[863], 46'b0};
assign col_1118 = {line_81[1024], line_80[1022], line_79[1020], line_78[1018], line_77[1016], line_76[1014], line_75[1012], line_74[1010], line_73[1008], line_72[1006], line_71[1004], line_70[1002], line_69[1000], line_68[998], line_67[996], line_66[994], line_65[992], line_64[990], line_63[988], line_62[986], line_61[984], line_60[982], line_59[980], line_58[978], line_57[976], line_56[974], line_55[972], line_54[970], line_53[968], line_52[966], line_51[964], line_50[962], line_49[960], line_48[958], line_47[956], line_46[954], line_45[952], line_44[950], line_43[948], line_42[946], line_41[944], line_40[942], line_39[940], line_38[938], line_37[936], line_36[934], line_35[932], line_34[930], line_33[928], line_32[926], line_31[924], line_30[922], line_29[920], line_28[918], line_27[916], line_26[914], line_25[912], line_24[910], line_23[908], line_22[906], line_21[904], line_20[902], line_19[900], line_18[898], line_17[896], line_16[894], line_15[892], line_14[890], line_13[888], line_12[886], line_11[884], line_10[882], line_9[880], line_8[878], line_7[876], line_6[874], line_5[872], line_4[870], line_3[868], line_2[866], line_1[864], 47'b0};
assign col_1119 = {line_81[1025], line_80[1023], line_79[1021], line_78[1019], line_77[1017], line_76[1015], line_75[1013], line_74[1011], line_73[1009], line_72[1007], line_71[1005], line_70[1003], line_69[1001], line_68[999], line_67[997], line_66[995], line_65[993], line_64[991], line_63[989], line_62[987], line_61[985], line_60[983], line_59[981], line_58[979], line_57[977], line_56[975], line_55[973], line_54[971], line_53[969], line_52[967], line_51[965], line_50[963], line_49[961], line_48[959], line_47[957], line_46[955], line_45[953], line_44[951], line_43[949], line_42[947], line_41[945], line_40[943], line_39[941], line_38[939], line_37[937], line_36[935], line_35[933], line_34[931], line_33[929], line_32[927], line_31[925], line_30[923], line_29[921], line_28[919], line_27[917], line_26[915], line_25[913], line_24[911], line_23[909], line_22[907], line_21[905], line_20[903], line_19[901], line_18[899], line_17[897], line_16[895], line_15[893], line_14[891], line_13[889], line_12[887], line_11[885], line_10[883], line_9[881], line_8[879], line_7[877], line_6[875], line_5[873], line_4[871], line_3[869], line_2[867], line_1[865], 47'b0};
assign col_1120 = {line_80[1024], line_79[1022], line_78[1020], line_77[1018], line_76[1016], line_75[1014], line_74[1012], line_73[1010], line_72[1008], line_71[1006], line_70[1004], line_69[1002], line_68[1000], line_67[998], line_66[996], line_65[994], line_64[992], line_63[990], line_62[988], line_61[986], line_60[984], line_59[982], line_58[980], line_57[978], line_56[976], line_55[974], line_54[972], line_53[970], line_52[968], line_51[966], line_50[964], line_49[962], line_48[960], line_47[958], line_46[956], line_45[954], line_44[952], line_43[950], line_42[948], line_41[946], line_40[944], line_39[942], line_38[940], line_37[938], line_36[936], line_35[934], line_34[932], line_33[930], line_32[928], line_31[926], line_30[924], line_29[922], line_28[920], line_27[918], line_26[916], line_25[914], line_24[912], line_23[910], line_22[908], line_21[906], line_20[904], line_19[902], line_18[900], line_17[898], line_16[896], line_15[894], line_14[892], line_13[890], line_12[888], line_11[886], line_10[884], line_9[882], line_8[880], line_7[878], line_6[876], line_5[874], line_4[872], line_3[870], line_2[868], line_1[866], 48'b0};
assign col_1121 = {line_80[1025], line_79[1023], line_78[1021], line_77[1019], line_76[1017], line_75[1015], line_74[1013], line_73[1011], line_72[1009], line_71[1007], line_70[1005], line_69[1003], line_68[1001], line_67[999], line_66[997], line_65[995], line_64[993], line_63[991], line_62[989], line_61[987], line_60[985], line_59[983], line_58[981], line_57[979], line_56[977], line_55[975], line_54[973], line_53[971], line_52[969], line_51[967], line_50[965], line_49[963], line_48[961], line_47[959], line_46[957], line_45[955], line_44[953], line_43[951], line_42[949], line_41[947], line_40[945], line_39[943], line_38[941], line_37[939], line_36[937], line_35[935], line_34[933], line_33[931], line_32[929], line_31[927], line_30[925], line_29[923], line_28[921], line_27[919], line_26[917], line_25[915], line_24[913], line_23[911], line_22[909], line_21[907], line_20[905], line_19[903], line_18[901], line_17[899], line_16[897], line_15[895], line_14[893], line_13[891], line_12[889], line_11[887], line_10[885], line_9[883], line_8[881], line_7[879], line_6[877], line_5[875], line_4[873], line_3[871], line_2[869], line_1[867], 48'b0};
assign col_1122 = {line_79[1024], line_78[1022], line_77[1020], line_76[1018], line_75[1016], line_74[1014], line_73[1012], line_72[1010], line_71[1008], line_70[1006], line_69[1004], line_68[1002], line_67[1000], line_66[998], line_65[996], line_64[994], line_63[992], line_62[990], line_61[988], line_60[986], line_59[984], line_58[982], line_57[980], line_56[978], line_55[976], line_54[974], line_53[972], line_52[970], line_51[968], line_50[966], line_49[964], line_48[962], line_47[960], line_46[958], line_45[956], line_44[954], line_43[952], line_42[950], line_41[948], line_40[946], line_39[944], line_38[942], line_37[940], line_36[938], line_35[936], line_34[934], line_33[932], line_32[930], line_31[928], line_30[926], line_29[924], line_28[922], line_27[920], line_26[918], line_25[916], line_24[914], line_23[912], line_22[910], line_21[908], line_20[906], line_19[904], line_18[902], line_17[900], line_16[898], line_15[896], line_14[894], line_13[892], line_12[890], line_11[888], line_10[886], line_9[884], line_8[882], line_7[880], line_6[878], line_5[876], line_4[874], line_3[872], line_2[870], line_1[868], 49'b0};
assign col_1123 = {line_79[1025], line_78[1023], line_77[1021], line_76[1019], line_75[1017], line_74[1015], line_73[1013], line_72[1011], line_71[1009], line_70[1007], line_69[1005], line_68[1003], line_67[1001], line_66[999], line_65[997], line_64[995], line_63[993], line_62[991], line_61[989], line_60[987], line_59[985], line_58[983], line_57[981], line_56[979], line_55[977], line_54[975], line_53[973], line_52[971], line_51[969], line_50[967], line_49[965], line_48[963], line_47[961], line_46[959], line_45[957], line_44[955], line_43[953], line_42[951], line_41[949], line_40[947], line_39[945], line_38[943], line_37[941], line_36[939], line_35[937], line_34[935], line_33[933], line_32[931], line_31[929], line_30[927], line_29[925], line_28[923], line_27[921], line_26[919], line_25[917], line_24[915], line_23[913], line_22[911], line_21[909], line_20[907], line_19[905], line_18[903], line_17[901], line_16[899], line_15[897], line_14[895], line_13[893], line_12[891], line_11[889], line_10[887], line_9[885], line_8[883], line_7[881], line_6[879], line_5[877], line_4[875], line_3[873], line_2[871], line_1[869], 49'b0};
assign col_1124 = {line_78[1024], line_77[1022], line_76[1020], line_75[1018], line_74[1016], line_73[1014], line_72[1012], line_71[1010], line_70[1008], line_69[1006], line_68[1004], line_67[1002], line_66[1000], line_65[998], line_64[996], line_63[994], line_62[992], line_61[990], line_60[988], line_59[986], line_58[984], line_57[982], line_56[980], line_55[978], line_54[976], line_53[974], line_52[972], line_51[970], line_50[968], line_49[966], line_48[964], line_47[962], line_46[960], line_45[958], line_44[956], line_43[954], line_42[952], line_41[950], line_40[948], line_39[946], line_38[944], line_37[942], line_36[940], line_35[938], line_34[936], line_33[934], line_32[932], line_31[930], line_30[928], line_29[926], line_28[924], line_27[922], line_26[920], line_25[918], line_24[916], line_23[914], line_22[912], line_21[910], line_20[908], line_19[906], line_18[904], line_17[902], line_16[900], line_15[898], line_14[896], line_13[894], line_12[892], line_11[890], line_10[888], line_9[886], line_8[884], line_7[882], line_6[880], line_5[878], line_4[876], line_3[874], line_2[872], line_1[870], 50'b0};
assign col_1125 = {line_78[1025], line_77[1023], line_76[1021], line_75[1019], line_74[1017], line_73[1015], line_72[1013], line_71[1011], line_70[1009], line_69[1007], line_68[1005], line_67[1003], line_66[1001], line_65[999], line_64[997], line_63[995], line_62[993], line_61[991], line_60[989], line_59[987], line_58[985], line_57[983], line_56[981], line_55[979], line_54[977], line_53[975], line_52[973], line_51[971], line_50[969], line_49[967], line_48[965], line_47[963], line_46[961], line_45[959], line_44[957], line_43[955], line_42[953], line_41[951], line_40[949], line_39[947], line_38[945], line_37[943], line_36[941], line_35[939], line_34[937], line_33[935], line_32[933], line_31[931], line_30[929], line_29[927], line_28[925], line_27[923], line_26[921], line_25[919], line_24[917], line_23[915], line_22[913], line_21[911], line_20[909], line_19[907], line_18[905], line_17[903], line_16[901], line_15[899], line_14[897], line_13[895], line_12[893], line_11[891], line_10[889], line_9[887], line_8[885], line_7[883], line_6[881], line_5[879], line_4[877], line_3[875], line_2[873], line_1[871], 50'b0};
assign col_1126 = {line_77[1024], line_76[1022], line_75[1020], line_74[1018], line_73[1016], line_72[1014], line_71[1012], line_70[1010], line_69[1008], line_68[1006], line_67[1004], line_66[1002], line_65[1000], line_64[998], line_63[996], line_62[994], line_61[992], line_60[990], line_59[988], line_58[986], line_57[984], line_56[982], line_55[980], line_54[978], line_53[976], line_52[974], line_51[972], line_50[970], line_49[968], line_48[966], line_47[964], line_46[962], line_45[960], line_44[958], line_43[956], line_42[954], line_41[952], line_40[950], line_39[948], line_38[946], line_37[944], line_36[942], line_35[940], line_34[938], line_33[936], line_32[934], line_31[932], line_30[930], line_29[928], line_28[926], line_27[924], line_26[922], line_25[920], line_24[918], line_23[916], line_22[914], line_21[912], line_20[910], line_19[908], line_18[906], line_17[904], line_16[902], line_15[900], line_14[898], line_13[896], line_12[894], line_11[892], line_10[890], line_9[888], line_8[886], line_7[884], line_6[882], line_5[880], line_4[878], line_3[876], line_2[874], line_1[872], 51'b0};
assign col_1127 = {line_77[1025], line_76[1023], line_75[1021], line_74[1019], line_73[1017], line_72[1015], line_71[1013], line_70[1011], line_69[1009], line_68[1007], line_67[1005], line_66[1003], line_65[1001], line_64[999], line_63[997], line_62[995], line_61[993], line_60[991], line_59[989], line_58[987], line_57[985], line_56[983], line_55[981], line_54[979], line_53[977], line_52[975], line_51[973], line_50[971], line_49[969], line_48[967], line_47[965], line_46[963], line_45[961], line_44[959], line_43[957], line_42[955], line_41[953], line_40[951], line_39[949], line_38[947], line_37[945], line_36[943], line_35[941], line_34[939], line_33[937], line_32[935], line_31[933], line_30[931], line_29[929], line_28[927], line_27[925], line_26[923], line_25[921], line_24[919], line_23[917], line_22[915], line_21[913], line_20[911], line_19[909], line_18[907], line_17[905], line_16[903], line_15[901], line_14[899], line_13[897], line_12[895], line_11[893], line_10[891], line_9[889], line_8[887], line_7[885], line_6[883], line_5[881], line_4[879], line_3[877], line_2[875], line_1[873], 51'b0};
assign col_1128 = {line_76[1024], line_75[1022], line_74[1020], line_73[1018], line_72[1016], line_71[1014], line_70[1012], line_69[1010], line_68[1008], line_67[1006], line_66[1004], line_65[1002], line_64[1000], line_63[998], line_62[996], line_61[994], line_60[992], line_59[990], line_58[988], line_57[986], line_56[984], line_55[982], line_54[980], line_53[978], line_52[976], line_51[974], line_50[972], line_49[970], line_48[968], line_47[966], line_46[964], line_45[962], line_44[960], line_43[958], line_42[956], line_41[954], line_40[952], line_39[950], line_38[948], line_37[946], line_36[944], line_35[942], line_34[940], line_33[938], line_32[936], line_31[934], line_30[932], line_29[930], line_28[928], line_27[926], line_26[924], line_25[922], line_24[920], line_23[918], line_22[916], line_21[914], line_20[912], line_19[910], line_18[908], line_17[906], line_16[904], line_15[902], line_14[900], line_13[898], line_12[896], line_11[894], line_10[892], line_9[890], line_8[888], line_7[886], line_6[884], line_5[882], line_4[880], line_3[878], line_2[876], line_1[874], 52'b0};
assign col_1129 = {line_76[1025], line_75[1023], line_74[1021], line_73[1019], line_72[1017], line_71[1015], line_70[1013], line_69[1011], line_68[1009], line_67[1007], line_66[1005], line_65[1003], line_64[1001], line_63[999], line_62[997], line_61[995], line_60[993], line_59[991], line_58[989], line_57[987], line_56[985], line_55[983], line_54[981], line_53[979], line_52[977], line_51[975], line_50[973], line_49[971], line_48[969], line_47[967], line_46[965], line_45[963], line_44[961], line_43[959], line_42[957], line_41[955], line_40[953], line_39[951], line_38[949], line_37[947], line_36[945], line_35[943], line_34[941], line_33[939], line_32[937], line_31[935], line_30[933], line_29[931], line_28[929], line_27[927], line_26[925], line_25[923], line_24[921], line_23[919], line_22[917], line_21[915], line_20[913], line_19[911], line_18[909], line_17[907], line_16[905], line_15[903], line_14[901], line_13[899], line_12[897], line_11[895], line_10[893], line_9[891], line_8[889], line_7[887], line_6[885], line_5[883], line_4[881], line_3[879], line_2[877], line_1[875], 52'b0};
assign col_1130 = {line_75[1024], line_74[1022], line_73[1020], line_72[1018], line_71[1016], line_70[1014], line_69[1012], line_68[1010], line_67[1008], line_66[1006], line_65[1004], line_64[1002], line_63[1000], line_62[998], line_61[996], line_60[994], line_59[992], line_58[990], line_57[988], line_56[986], line_55[984], line_54[982], line_53[980], line_52[978], line_51[976], line_50[974], line_49[972], line_48[970], line_47[968], line_46[966], line_45[964], line_44[962], line_43[960], line_42[958], line_41[956], line_40[954], line_39[952], line_38[950], line_37[948], line_36[946], line_35[944], line_34[942], line_33[940], line_32[938], line_31[936], line_30[934], line_29[932], line_28[930], line_27[928], line_26[926], line_25[924], line_24[922], line_23[920], line_22[918], line_21[916], line_20[914], line_19[912], line_18[910], line_17[908], line_16[906], line_15[904], line_14[902], line_13[900], line_12[898], line_11[896], line_10[894], line_9[892], line_8[890], line_7[888], line_6[886], line_5[884], line_4[882], line_3[880], line_2[878], line_1[876], 53'b0};
assign col_1131 = {line_75[1025], line_74[1023], line_73[1021], line_72[1019], line_71[1017], line_70[1015], line_69[1013], line_68[1011], line_67[1009], line_66[1007], line_65[1005], line_64[1003], line_63[1001], line_62[999], line_61[997], line_60[995], line_59[993], line_58[991], line_57[989], line_56[987], line_55[985], line_54[983], line_53[981], line_52[979], line_51[977], line_50[975], line_49[973], line_48[971], line_47[969], line_46[967], line_45[965], line_44[963], line_43[961], line_42[959], line_41[957], line_40[955], line_39[953], line_38[951], line_37[949], line_36[947], line_35[945], line_34[943], line_33[941], line_32[939], line_31[937], line_30[935], line_29[933], line_28[931], line_27[929], line_26[927], line_25[925], line_24[923], line_23[921], line_22[919], line_21[917], line_20[915], line_19[913], line_18[911], line_17[909], line_16[907], line_15[905], line_14[903], line_13[901], line_12[899], line_11[897], line_10[895], line_9[893], line_8[891], line_7[889], line_6[887], line_5[885], line_4[883], line_3[881], line_2[879], line_1[877], 53'b0};
assign col_1132 = {line_74[1024], line_73[1022], line_72[1020], line_71[1018], line_70[1016], line_69[1014], line_68[1012], line_67[1010], line_66[1008], line_65[1006], line_64[1004], line_63[1002], line_62[1000], line_61[998], line_60[996], line_59[994], line_58[992], line_57[990], line_56[988], line_55[986], line_54[984], line_53[982], line_52[980], line_51[978], line_50[976], line_49[974], line_48[972], line_47[970], line_46[968], line_45[966], line_44[964], line_43[962], line_42[960], line_41[958], line_40[956], line_39[954], line_38[952], line_37[950], line_36[948], line_35[946], line_34[944], line_33[942], line_32[940], line_31[938], line_30[936], line_29[934], line_28[932], line_27[930], line_26[928], line_25[926], line_24[924], line_23[922], line_22[920], line_21[918], line_20[916], line_19[914], line_18[912], line_17[910], line_16[908], line_15[906], line_14[904], line_13[902], line_12[900], line_11[898], line_10[896], line_9[894], line_8[892], line_7[890], line_6[888], line_5[886], line_4[884], line_3[882], line_2[880], line_1[878], 54'b0};
assign col_1133 = {line_74[1025], line_73[1023], line_72[1021], line_71[1019], line_70[1017], line_69[1015], line_68[1013], line_67[1011], line_66[1009], line_65[1007], line_64[1005], line_63[1003], line_62[1001], line_61[999], line_60[997], line_59[995], line_58[993], line_57[991], line_56[989], line_55[987], line_54[985], line_53[983], line_52[981], line_51[979], line_50[977], line_49[975], line_48[973], line_47[971], line_46[969], line_45[967], line_44[965], line_43[963], line_42[961], line_41[959], line_40[957], line_39[955], line_38[953], line_37[951], line_36[949], line_35[947], line_34[945], line_33[943], line_32[941], line_31[939], line_30[937], line_29[935], line_28[933], line_27[931], line_26[929], line_25[927], line_24[925], line_23[923], line_22[921], line_21[919], line_20[917], line_19[915], line_18[913], line_17[911], line_16[909], line_15[907], line_14[905], line_13[903], line_12[901], line_11[899], line_10[897], line_9[895], line_8[893], line_7[891], line_6[889], line_5[887], line_4[885], line_3[883], line_2[881], line_1[879], 54'b0};
assign col_1134 = {line_73[1024], line_72[1022], line_71[1020], line_70[1018], line_69[1016], line_68[1014], line_67[1012], line_66[1010], line_65[1008], line_64[1006], line_63[1004], line_62[1002], line_61[1000], line_60[998], line_59[996], line_58[994], line_57[992], line_56[990], line_55[988], line_54[986], line_53[984], line_52[982], line_51[980], line_50[978], line_49[976], line_48[974], line_47[972], line_46[970], line_45[968], line_44[966], line_43[964], line_42[962], line_41[960], line_40[958], line_39[956], line_38[954], line_37[952], line_36[950], line_35[948], line_34[946], line_33[944], line_32[942], line_31[940], line_30[938], line_29[936], line_28[934], line_27[932], line_26[930], line_25[928], line_24[926], line_23[924], line_22[922], line_21[920], line_20[918], line_19[916], line_18[914], line_17[912], line_16[910], line_15[908], line_14[906], line_13[904], line_12[902], line_11[900], line_10[898], line_9[896], line_8[894], line_7[892], line_6[890], line_5[888], line_4[886], line_3[884], line_2[882], line_1[880], 55'b0};
assign col_1135 = {line_73[1025], line_72[1023], line_71[1021], line_70[1019], line_69[1017], line_68[1015], line_67[1013], line_66[1011], line_65[1009], line_64[1007], line_63[1005], line_62[1003], line_61[1001], line_60[999], line_59[997], line_58[995], line_57[993], line_56[991], line_55[989], line_54[987], line_53[985], line_52[983], line_51[981], line_50[979], line_49[977], line_48[975], line_47[973], line_46[971], line_45[969], line_44[967], line_43[965], line_42[963], line_41[961], line_40[959], line_39[957], line_38[955], line_37[953], line_36[951], line_35[949], line_34[947], line_33[945], line_32[943], line_31[941], line_30[939], line_29[937], line_28[935], line_27[933], line_26[931], line_25[929], line_24[927], line_23[925], line_22[923], line_21[921], line_20[919], line_19[917], line_18[915], line_17[913], line_16[911], line_15[909], line_14[907], line_13[905], line_12[903], line_11[901], line_10[899], line_9[897], line_8[895], line_7[893], line_6[891], line_5[889], line_4[887], line_3[885], line_2[883], line_1[881], 55'b0};
assign col_1136 = {line_72[1024], line_71[1022], line_70[1020], line_69[1018], line_68[1016], line_67[1014], line_66[1012], line_65[1010], line_64[1008], line_63[1006], line_62[1004], line_61[1002], line_60[1000], line_59[998], line_58[996], line_57[994], line_56[992], line_55[990], line_54[988], line_53[986], line_52[984], line_51[982], line_50[980], line_49[978], line_48[976], line_47[974], line_46[972], line_45[970], line_44[968], line_43[966], line_42[964], line_41[962], line_40[960], line_39[958], line_38[956], line_37[954], line_36[952], line_35[950], line_34[948], line_33[946], line_32[944], line_31[942], line_30[940], line_29[938], line_28[936], line_27[934], line_26[932], line_25[930], line_24[928], line_23[926], line_22[924], line_21[922], line_20[920], line_19[918], line_18[916], line_17[914], line_16[912], line_15[910], line_14[908], line_13[906], line_12[904], line_11[902], line_10[900], line_9[898], line_8[896], line_7[894], line_6[892], line_5[890], line_4[888], line_3[886], line_2[884], line_1[882], 56'b0};
assign col_1137 = {line_72[1025], line_71[1023], line_70[1021], line_69[1019], line_68[1017], line_67[1015], line_66[1013], line_65[1011], line_64[1009], line_63[1007], line_62[1005], line_61[1003], line_60[1001], line_59[999], line_58[997], line_57[995], line_56[993], line_55[991], line_54[989], line_53[987], line_52[985], line_51[983], line_50[981], line_49[979], line_48[977], line_47[975], line_46[973], line_45[971], line_44[969], line_43[967], line_42[965], line_41[963], line_40[961], line_39[959], line_38[957], line_37[955], line_36[953], line_35[951], line_34[949], line_33[947], line_32[945], line_31[943], line_30[941], line_29[939], line_28[937], line_27[935], line_26[933], line_25[931], line_24[929], line_23[927], line_22[925], line_21[923], line_20[921], line_19[919], line_18[917], line_17[915], line_16[913], line_15[911], line_14[909], line_13[907], line_12[905], line_11[903], line_10[901], line_9[899], line_8[897], line_7[895], line_6[893], line_5[891], line_4[889], line_3[887], line_2[885], line_1[883], 56'b0};
assign col_1138 = {line_71[1024], line_70[1022], line_69[1020], line_68[1018], line_67[1016], line_66[1014], line_65[1012], line_64[1010], line_63[1008], line_62[1006], line_61[1004], line_60[1002], line_59[1000], line_58[998], line_57[996], line_56[994], line_55[992], line_54[990], line_53[988], line_52[986], line_51[984], line_50[982], line_49[980], line_48[978], line_47[976], line_46[974], line_45[972], line_44[970], line_43[968], line_42[966], line_41[964], line_40[962], line_39[960], line_38[958], line_37[956], line_36[954], line_35[952], line_34[950], line_33[948], line_32[946], line_31[944], line_30[942], line_29[940], line_28[938], line_27[936], line_26[934], line_25[932], line_24[930], line_23[928], line_22[926], line_21[924], line_20[922], line_19[920], line_18[918], line_17[916], line_16[914], line_15[912], line_14[910], line_13[908], line_12[906], line_11[904], line_10[902], line_9[900], line_8[898], line_7[896], line_6[894], line_5[892], line_4[890], line_3[888], line_2[886], line_1[884], 57'b0};
assign col_1139 = {line_71[1025], line_70[1023], line_69[1021], line_68[1019], line_67[1017], line_66[1015], line_65[1013], line_64[1011], line_63[1009], line_62[1007], line_61[1005], line_60[1003], line_59[1001], line_58[999], line_57[997], line_56[995], line_55[993], line_54[991], line_53[989], line_52[987], line_51[985], line_50[983], line_49[981], line_48[979], line_47[977], line_46[975], line_45[973], line_44[971], line_43[969], line_42[967], line_41[965], line_40[963], line_39[961], line_38[959], line_37[957], line_36[955], line_35[953], line_34[951], line_33[949], line_32[947], line_31[945], line_30[943], line_29[941], line_28[939], line_27[937], line_26[935], line_25[933], line_24[931], line_23[929], line_22[927], line_21[925], line_20[923], line_19[921], line_18[919], line_17[917], line_16[915], line_15[913], line_14[911], line_13[909], line_12[907], line_11[905], line_10[903], line_9[901], line_8[899], line_7[897], line_6[895], line_5[893], line_4[891], line_3[889], line_2[887], line_1[885], 57'b0};
assign col_1140 = {line_70[1024], line_69[1022], line_68[1020], line_67[1018], line_66[1016], line_65[1014], line_64[1012], line_63[1010], line_62[1008], line_61[1006], line_60[1004], line_59[1002], line_58[1000], line_57[998], line_56[996], line_55[994], line_54[992], line_53[990], line_52[988], line_51[986], line_50[984], line_49[982], line_48[980], line_47[978], line_46[976], line_45[974], line_44[972], line_43[970], line_42[968], line_41[966], line_40[964], line_39[962], line_38[960], line_37[958], line_36[956], line_35[954], line_34[952], line_33[950], line_32[948], line_31[946], line_30[944], line_29[942], line_28[940], line_27[938], line_26[936], line_25[934], line_24[932], line_23[930], line_22[928], line_21[926], line_20[924], line_19[922], line_18[920], line_17[918], line_16[916], line_15[914], line_14[912], line_13[910], line_12[908], line_11[906], line_10[904], line_9[902], line_8[900], line_7[898], line_6[896], line_5[894], line_4[892], line_3[890], line_2[888], line_1[886], 58'b0};
assign col_1141 = {line_70[1025], line_69[1023], line_68[1021], line_67[1019], line_66[1017], line_65[1015], line_64[1013], line_63[1011], line_62[1009], line_61[1007], line_60[1005], line_59[1003], line_58[1001], line_57[999], line_56[997], line_55[995], line_54[993], line_53[991], line_52[989], line_51[987], line_50[985], line_49[983], line_48[981], line_47[979], line_46[977], line_45[975], line_44[973], line_43[971], line_42[969], line_41[967], line_40[965], line_39[963], line_38[961], line_37[959], line_36[957], line_35[955], line_34[953], line_33[951], line_32[949], line_31[947], line_30[945], line_29[943], line_28[941], line_27[939], line_26[937], line_25[935], line_24[933], line_23[931], line_22[929], line_21[927], line_20[925], line_19[923], line_18[921], line_17[919], line_16[917], line_15[915], line_14[913], line_13[911], line_12[909], line_11[907], line_10[905], line_9[903], line_8[901], line_7[899], line_6[897], line_5[895], line_4[893], line_3[891], line_2[889], line_1[887], 58'b0};
assign col_1142 = {line_69[1024], line_68[1022], line_67[1020], line_66[1018], line_65[1016], line_64[1014], line_63[1012], line_62[1010], line_61[1008], line_60[1006], line_59[1004], line_58[1002], line_57[1000], line_56[998], line_55[996], line_54[994], line_53[992], line_52[990], line_51[988], line_50[986], line_49[984], line_48[982], line_47[980], line_46[978], line_45[976], line_44[974], line_43[972], line_42[970], line_41[968], line_40[966], line_39[964], line_38[962], line_37[960], line_36[958], line_35[956], line_34[954], line_33[952], line_32[950], line_31[948], line_30[946], line_29[944], line_28[942], line_27[940], line_26[938], line_25[936], line_24[934], line_23[932], line_22[930], line_21[928], line_20[926], line_19[924], line_18[922], line_17[920], line_16[918], line_15[916], line_14[914], line_13[912], line_12[910], line_11[908], line_10[906], line_9[904], line_8[902], line_7[900], line_6[898], line_5[896], line_4[894], line_3[892], line_2[890], line_1[888], 59'b0};
assign col_1143 = {line_69[1025], line_68[1023], line_67[1021], line_66[1019], line_65[1017], line_64[1015], line_63[1013], line_62[1011], line_61[1009], line_60[1007], line_59[1005], line_58[1003], line_57[1001], line_56[999], line_55[997], line_54[995], line_53[993], line_52[991], line_51[989], line_50[987], line_49[985], line_48[983], line_47[981], line_46[979], line_45[977], line_44[975], line_43[973], line_42[971], line_41[969], line_40[967], line_39[965], line_38[963], line_37[961], line_36[959], line_35[957], line_34[955], line_33[953], line_32[951], line_31[949], line_30[947], line_29[945], line_28[943], line_27[941], line_26[939], line_25[937], line_24[935], line_23[933], line_22[931], line_21[929], line_20[927], line_19[925], line_18[923], line_17[921], line_16[919], line_15[917], line_14[915], line_13[913], line_12[911], line_11[909], line_10[907], line_9[905], line_8[903], line_7[901], line_6[899], line_5[897], line_4[895], line_3[893], line_2[891], line_1[889], 59'b0};
assign col_1144 = {line_68[1024], line_67[1022], line_66[1020], line_65[1018], line_64[1016], line_63[1014], line_62[1012], line_61[1010], line_60[1008], line_59[1006], line_58[1004], line_57[1002], line_56[1000], line_55[998], line_54[996], line_53[994], line_52[992], line_51[990], line_50[988], line_49[986], line_48[984], line_47[982], line_46[980], line_45[978], line_44[976], line_43[974], line_42[972], line_41[970], line_40[968], line_39[966], line_38[964], line_37[962], line_36[960], line_35[958], line_34[956], line_33[954], line_32[952], line_31[950], line_30[948], line_29[946], line_28[944], line_27[942], line_26[940], line_25[938], line_24[936], line_23[934], line_22[932], line_21[930], line_20[928], line_19[926], line_18[924], line_17[922], line_16[920], line_15[918], line_14[916], line_13[914], line_12[912], line_11[910], line_10[908], line_9[906], line_8[904], line_7[902], line_6[900], line_5[898], line_4[896], line_3[894], line_2[892], line_1[890], 60'b0};
assign col_1145 = {line_68[1025], line_67[1023], line_66[1021], line_65[1019], line_64[1017], line_63[1015], line_62[1013], line_61[1011], line_60[1009], line_59[1007], line_58[1005], line_57[1003], line_56[1001], line_55[999], line_54[997], line_53[995], line_52[993], line_51[991], line_50[989], line_49[987], line_48[985], line_47[983], line_46[981], line_45[979], line_44[977], line_43[975], line_42[973], line_41[971], line_40[969], line_39[967], line_38[965], line_37[963], line_36[961], line_35[959], line_34[957], line_33[955], line_32[953], line_31[951], line_30[949], line_29[947], line_28[945], line_27[943], line_26[941], line_25[939], line_24[937], line_23[935], line_22[933], line_21[931], line_20[929], line_19[927], line_18[925], line_17[923], line_16[921], line_15[919], line_14[917], line_13[915], line_12[913], line_11[911], line_10[909], line_9[907], line_8[905], line_7[903], line_6[901], line_5[899], line_4[897], line_3[895], line_2[893], line_1[891], 60'b0};
assign col_1146 = {line_67[1024], line_66[1022], line_65[1020], line_64[1018], line_63[1016], line_62[1014], line_61[1012], line_60[1010], line_59[1008], line_58[1006], line_57[1004], line_56[1002], line_55[1000], line_54[998], line_53[996], line_52[994], line_51[992], line_50[990], line_49[988], line_48[986], line_47[984], line_46[982], line_45[980], line_44[978], line_43[976], line_42[974], line_41[972], line_40[970], line_39[968], line_38[966], line_37[964], line_36[962], line_35[960], line_34[958], line_33[956], line_32[954], line_31[952], line_30[950], line_29[948], line_28[946], line_27[944], line_26[942], line_25[940], line_24[938], line_23[936], line_22[934], line_21[932], line_20[930], line_19[928], line_18[926], line_17[924], line_16[922], line_15[920], line_14[918], line_13[916], line_12[914], line_11[912], line_10[910], line_9[908], line_8[906], line_7[904], line_6[902], line_5[900], line_4[898], line_3[896], line_2[894], line_1[892], 61'b0};
assign col_1147 = {line_67[1025], line_66[1023], line_65[1021], line_64[1019], line_63[1017], line_62[1015], line_61[1013], line_60[1011], line_59[1009], line_58[1007], line_57[1005], line_56[1003], line_55[1001], line_54[999], line_53[997], line_52[995], line_51[993], line_50[991], line_49[989], line_48[987], line_47[985], line_46[983], line_45[981], line_44[979], line_43[977], line_42[975], line_41[973], line_40[971], line_39[969], line_38[967], line_37[965], line_36[963], line_35[961], line_34[959], line_33[957], line_32[955], line_31[953], line_30[951], line_29[949], line_28[947], line_27[945], line_26[943], line_25[941], line_24[939], line_23[937], line_22[935], line_21[933], line_20[931], line_19[929], line_18[927], line_17[925], line_16[923], line_15[921], line_14[919], line_13[917], line_12[915], line_11[913], line_10[911], line_9[909], line_8[907], line_7[905], line_6[903], line_5[901], line_4[899], line_3[897], line_2[895], line_1[893], 61'b0};
assign col_1148 = {line_66[1024], line_65[1022], line_64[1020], line_63[1018], line_62[1016], line_61[1014], line_60[1012], line_59[1010], line_58[1008], line_57[1006], line_56[1004], line_55[1002], line_54[1000], line_53[998], line_52[996], line_51[994], line_50[992], line_49[990], line_48[988], line_47[986], line_46[984], line_45[982], line_44[980], line_43[978], line_42[976], line_41[974], line_40[972], line_39[970], line_38[968], line_37[966], line_36[964], line_35[962], line_34[960], line_33[958], line_32[956], line_31[954], line_30[952], line_29[950], line_28[948], line_27[946], line_26[944], line_25[942], line_24[940], line_23[938], line_22[936], line_21[934], line_20[932], line_19[930], line_18[928], line_17[926], line_16[924], line_15[922], line_14[920], line_13[918], line_12[916], line_11[914], line_10[912], line_9[910], line_8[908], line_7[906], line_6[904], line_5[902], line_4[900], line_3[898], line_2[896], line_1[894], 62'b0};
assign col_1149 = {line_66[1025], line_65[1023], line_64[1021], line_63[1019], line_62[1017], line_61[1015], line_60[1013], line_59[1011], line_58[1009], line_57[1007], line_56[1005], line_55[1003], line_54[1001], line_53[999], line_52[997], line_51[995], line_50[993], line_49[991], line_48[989], line_47[987], line_46[985], line_45[983], line_44[981], line_43[979], line_42[977], line_41[975], line_40[973], line_39[971], line_38[969], line_37[967], line_36[965], line_35[963], line_34[961], line_33[959], line_32[957], line_31[955], line_30[953], line_29[951], line_28[949], line_27[947], line_26[945], line_25[943], line_24[941], line_23[939], line_22[937], line_21[935], line_20[933], line_19[931], line_18[929], line_17[927], line_16[925], line_15[923], line_14[921], line_13[919], line_12[917], line_11[915], line_10[913], line_9[911], line_8[909], line_7[907], line_6[905], line_5[903], line_4[901], line_3[899], line_2[897], line_1[895], 62'b0};
assign col_1150 = {line_65[1024], line_64[1022], line_63[1020], line_62[1018], line_61[1016], line_60[1014], line_59[1012], line_58[1010], line_57[1008], line_56[1006], line_55[1004], line_54[1002], line_53[1000], line_52[998], line_51[996], line_50[994], line_49[992], line_48[990], line_47[988], line_46[986], line_45[984], line_44[982], line_43[980], line_42[978], line_41[976], line_40[974], line_39[972], line_38[970], line_37[968], line_36[966], line_35[964], line_34[962], line_33[960], line_32[958], line_31[956], line_30[954], line_29[952], line_28[950], line_27[948], line_26[946], line_25[944], line_24[942], line_23[940], line_22[938], line_21[936], line_20[934], line_19[932], line_18[930], line_17[928], line_16[926], line_15[924], line_14[922], line_13[920], line_12[918], line_11[916], line_10[914], line_9[912], line_8[910], line_7[908], line_6[906], line_5[904], line_4[902], line_3[900], line_2[898], line_1[896], 63'b0};
assign col_1151 = {line_65[1025], line_64[1023], line_63[1021], line_62[1019], line_61[1017], line_60[1015], line_59[1013], line_58[1011], line_57[1009], line_56[1007], line_55[1005], line_54[1003], line_53[1001], line_52[999], line_51[997], line_50[995], line_49[993], line_48[991], line_47[989], line_46[987], line_45[985], line_44[983], line_43[981], line_42[979], line_41[977], line_40[975], line_39[973], line_38[971], line_37[969], line_36[967], line_35[965], line_34[963], line_33[961], line_32[959], line_31[957], line_30[955], line_29[953], line_28[951], line_27[949], line_26[947], line_25[945], line_24[943], line_23[941], line_22[939], line_21[937], line_20[935], line_19[933], line_18[931], line_17[929], line_16[927], line_15[925], line_14[923], line_13[921], line_12[919], line_11[917], line_10[915], line_9[913], line_8[911], line_7[909], line_6[907], line_5[905], line_4[903], line_3[901], line_2[899], line_1[897], 63'b0};
assign col_1152 = {line_64[1024], line_63[1022], line_62[1020], line_61[1018], line_60[1016], line_59[1014], line_58[1012], line_57[1010], line_56[1008], line_55[1006], line_54[1004], line_53[1002], line_52[1000], line_51[998], line_50[996], line_49[994], line_48[992], line_47[990], line_46[988], line_45[986], line_44[984], line_43[982], line_42[980], line_41[978], line_40[976], line_39[974], line_38[972], line_37[970], line_36[968], line_35[966], line_34[964], line_33[962], line_32[960], line_31[958], line_30[956], line_29[954], line_28[952], line_27[950], line_26[948], line_25[946], line_24[944], line_23[942], line_22[940], line_21[938], line_20[936], line_19[934], line_18[932], line_17[930], line_16[928], line_15[926], line_14[924], line_13[922], line_12[920], line_11[918], line_10[916], line_9[914], line_8[912], line_7[910], line_6[908], line_5[906], line_4[904], line_3[902], line_2[900], line_1[898], 64'b0};
assign col_1153 = {line_64[1025], line_63[1023], line_62[1021], line_61[1019], line_60[1017], line_59[1015], line_58[1013], line_57[1011], line_56[1009], line_55[1007], line_54[1005], line_53[1003], line_52[1001], line_51[999], line_50[997], line_49[995], line_48[993], line_47[991], line_46[989], line_45[987], line_44[985], line_43[983], line_42[981], line_41[979], line_40[977], line_39[975], line_38[973], line_37[971], line_36[969], line_35[967], line_34[965], line_33[963], line_32[961], line_31[959], line_30[957], line_29[955], line_28[953], line_27[951], line_26[949], line_25[947], line_24[945], line_23[943], line_22[941], line_21[939], line_20[937], line_19[935], line_18[933], line_17[931], line_16[929], line_15[927], line_14[925], line_13[923], line_12[921], line_11[919], line_10[917], line_9[915], line_8[913], line_7[911], line_6[909], line_5[907], line_4[905], line_3[903], line_2[901], line_1[899], 64'b0};
assign col_1154 = {line_63[1024], line_62[1022], line_61[1020], line_60[1018], line_59[1016], line_58[1014], line_57[1012], line_56[1010], line_55[1008], line_54[1006], line_53[1004], line_52[1002], line_51[1000], line_50[998], line_49[996], line_48[994], line_47[992], line_46[990], line_45[988], line_44[986], line_43[984], line_42[982], line_41[980], line_40[978], line_39[976], line_38[974], line_37[972], line_36[970], line_35[968], line_34[966], line_33[964], line_32[962], line_31[960], line_30[958], line_29[956], line_28[954], line_27[952], line_26[950], line_25[948], line_24[946], line_23[944], line_22[942], line_21[940], line_20[938], line_19[936], line_18[934], line_17[932], line_16[930], line_15[928], line_14[926], line_13[924], line_12[922], line_11[920], line_10[918], line_9[916], line_8[914], line_7[912], line_6[910], line_5[908], line_4[906], line_3[904], line_2[902], line_1[900], 65'b0};
assign col_1155 = {line_63[1025], line_62[1023], line_61[1021], line_60[1019], line_59[1017], line_58[1015], line_57[1013], line_56[1011], line_55[1009], line_54[1007], line_53[1005], line_52[1003], line_51[1001], line_50[999], line_49[997], line_48[995], line_47[993], line_46[991], line_45[989], line_44[987], line_43[985], line_42[983], line_41[981], line_40[979], line_39[977], line_38[975], line_37[973], line_36[971], line_35[969], line_34[967], line_33[965], line_32[963], line_31[961], line_30[959], line_29[957], line_28[955], line_27[953], line_26[951], line_25[949], line_24[947], line_23[945], line_22[943], line_21[941], line_20[939], line_19[937], line_18[935], line_17[933], line_16[931], line_15[929], line_14[927], line_13[925], line_12[923], line_11[921], line_10[919], line_9[917], line_8[915], line_7[913], line_6[911], line_5[909], line_4[907], line_3[905], line_2[903], line_1[901], 65'b0};
assign col_1156 = {line_62[1024], line_61[1022], line_60[1020], line_59[1018], line_58[1016], line_57[1014], line_56[1012], line_55[1010], line_54[1008], line_53[1006], line_52[1004], line_51[1002], line_50[1000], line_49[998], line_48[996], line_47[994], line_46[992], line_45[990], line_44[988], line_43[986], line_42[984], line_41[982], line_40[980], line_39[978], line_38[976], line_37[974], line_36[972], line_35[970], line_34[968], line_33[966], line_32[964], line_31[962], line_30[960], line_29[958], line_28[956], line_27[954], line_26[952], line_25[950], line_24[948], line_23[946], line_22[944], line_21[942], line_20[940], line_19[938], line_18[936], line_17[934], line_16[932], line_15[930], line_14[928], line_13[926], line_12[924], line_11[922], line_10[920], line_9[918], line_8[916], line_7[914], line_6[912], line_5[910], line_4[908], line_3[906], line_2[904], line_1[902], 66'b0};
assign col_1157 = {line_62[1025], line_61[1023], line_60[1021], line_59[1019], line_58[1017], line_57[1015], line_56[1013], line_55[1011], line_54[1009], line_53[1007], line_52[1005], line_51[1003], line_50[1001], line_49[999], line_48[997], line_47[995], line_46[993], line_45[991], line_44[989], line_43[987], line_42[985], line_41[983], line_40[981], line_39[979], line_38[977], line_37[975], line_36[973], line_35[971], line_34[969], line_33[967], line_32[965], line_31[963], line_30[961], line_29[959], line_28[957], line_27[955], line_26[953], line_25[951], line_24[949], line_23[947], line_22[945], line_21[943], line_20[941], line_19[939], line_18[937], line_17[935], line_16[933], line_15[931], line_14[929], line_13[927], line_12[925], line_11[923], line_10[921], line_9[919], line_8[917], line_7[915], line_6[913], line_5[911], line_4[909], line_3[907], line_2[905], line_1[903], 66'b0};
assign col_1158 = {line_61[1024], line_60[1022], line_59[1020], line_58[1018], line_57[1016], line_56[1014], line_55[1012], line_54[1010], line_53[1008], line_52[1006], line_51[1004], line_50[1002], line_49[1000], line_48[998], line_47[996], line_46[994], line_45[992], line_44[990], line_43[988], line_42[986], line_41[984], line_40[982], line_39[980], line_38[978], line_37[976], line_36[974], line_35[972], line_34[970], line_33[968], line_32[966], line_31[964], line_30[962], line_29[960], line_28[958], line_27[956], line_26[954], line_25[952], line_24[950], line_23[948], line_22[946], line_21[944], line_20[942], line_19[940], line_18[938], line_17[936], line_16[934], line_15[932], line_14[930], line_13[928], line_12[926], line_11[924], line_10[922], line_9[920], line_8[918], line_7[916], line_6[914], line_5[912], line_4[910], line_3[908], line_2[906], line_1[904], 67'b0};
assign col_1159 = {line_61[1025], line_60[1023], line_59[1021], line_58[1019], line_57[1017], line_56[1015], line_55[1013], line_54[1011], line_53[1009], line_52[1007], line_51[1005], line_50[1003], line_49[1001], line_48[999], line_47[997], line_46[995], line_45[993], line_44[991], line_43[989], line_42[987], line_41[985], line_40[983], line_39[981], line_38[979], line_37[977], line_36[975], line_35[973], line_34[971], line_33[969], line_32[967], line_31[965], line_30[963], line_29[961], line_28[959], line_27[957], line_26[955], line_25[953], line_24[951], line_23[949], line_22[947], line_21[945], line_20[943], line_19[941], line_18[939], line_17[937], line_16[935], line_15[933], line_14[931], line_13[929], line_12[927], line_11[925], line_10[923], line_9[921], line_8[919], line_7[917], line_6[915], line_5[913], line_4[911], line_3[909], line_2[907], line_1[905], 67'b0};
assign col_1160 = {line_60[1024], line_59[1022], line_58[1020], line_57[1018], line_56[1016], line_55[1014], line_54[1012], line_53[1010], line_52[1008], line_51[1006], line_50[1004], line_49[1002], line_48[1000], line_47[998], line_46[996], line_45[994], line_44[992], line_43[990], line_42[988], line_41[986], line_40[984], line_39[982], line_38[980], line_37[978], line_36[976], line_35[974], line_34[972], line_33[970], line_32[968], line_31[966], line_30[964], line_29[962], line_28[960], line_27[958], line_26[956], line_25[954], line_24[952], line_23[950], line_22[948], line_21[946], line_20[944], line_19[942], line_18[940], line_17[938], line_16[936], line_15[934], line_14[932], line_13[930], line_12[928], line_11[926], line_10[924], line_9[922], line_8[920], line_7[918], line_6[916], line_5[914], line_4[912], line_3[910], line_2[908], line_1[906], 68'b0};
assign col_1161 = {line_60[1025], line_59[1023], line_58[1021], line_57[1019], line_56[1017], line_55[1015], line_54[1013], line_53[1011], line_52[1009], line_51[1007], line_50[1005], line_49[1003], line_48[1001], line_47[999], line_46[997], line_45[995], line_44[993], line_43[991], line_42[989], line_41[987], line_40[985], line_39[983], line_38[981], line_37[979], line_36[977], line_35[975], line_34[973], line_33[971], line_32[969], line_31[967], line_30[965], line_29[963], line_28[961], line_27[959], line_26[957], line_25[955], line_24[953], line_23[951], line_22[949], line_21[947], line_20[945], line_19[943], line_18[941], line_17[939], line_16[937], line_15[935], line_14[933], line_13[931], line_12[929], line_11[927], line_10[925], line_9[923], line_8[921], line_7[919], line_6[917], line_5[915], line_4[913], line_3[911], line_2[909], line_1[907], 68'b0};
assign col_1162 = {line_59[1024], line_58[1022], line_57[1020], line_56[1018], line_55[1016], line_54[1014], line_53[1012], line_52[1010], line_51[1008], line_50[1006], line_49[1004], line_48[1002], line_47[1000], line_46[998], line_45[996], line_44[994], line_43[992], line_42[990], line_41[988], line_40[986], line_39[984], line_38[982], line_37[980], line_36[978], line_35[976], line_34[974], line_33[972], line_32[970], line_31[968], line_30[966], line_29[964], line_28[962], line_27[960], line_26[958], line_25[956], line_24[954], line_23[952], line_22[950], line_21[948], line_20[946], line_19[944], line_18[942], line_17[940], line_16[938], line_15[936], line_14[934], line_13[932], line_12[930], line_11[928], line_10[926], line_9[924], line_8[922], line_7[920], line_6[918], line_5[916], line_4[914], line_3[912], line_2[910], line_1[908], 69'b0};
assign col_1163 = {line_59[1025], line_58[1023], line_57[1021], line_56[1019], line_55[1017], line_54[1015], line_53[1013], line_52[1011], line_51[1009], line_50[1007], line_49[1005], line_48[1003], line_47[1001], line_46[999], line_45[997], line_44[995], line_43[993], line_42[991], line_41[989], line_40[987], line_39[985], line_38[983], line_37[981], line_36[979], line_35[977], line_34[975], line_33[973], line_32[971], line_31[969], line_30[967], line_29[965], line_28[963], line_27[961], line_26[959], line_25[957], line_24[955], line_23[953], line_22[951], line_21[949], line_20[947], line_19[945], line_18[943], line_17[941], line_16[939], line_15[937], line_14[935], line_13[933], line_12[931], line_11[929], line_10[927], line_9[925], line_8[923], line_7[921], line_6[919], line_5[917], line_4[915], line_3[913], line_2[911], line_1[909], 69'b0};
assign col_1164 = {line_58[1024], line_57[1022], line_56[1020], line_55[1018], line_54[1016], line_53[1014], line_52[1012], line_51[1010], line_50[1008], line_49[1006], line_48[1004], line_47[1002], line_46[1000], line_45[998], line_44[996], line_43[994], line_42[992], line_41[990], line_40[988], line_39[986], line_38[984], line_37[982], line_36[980], line_35[978], line_34[976], line_33[974], line_32[972], line_31[970], line_30[968], line_29[966], line_28[964], line_27[962], line_26[960], line_25[958], line_24[956], line_23[954], line_22[952], line_21[950], line_20[948], line_19[946], line_18[944], line_17[942], line_16[940], line_15[938], line_14[936], line_13[934], line_12[932], line_11[930], line_10[928], line_9[926], line_8[924], line_7[922], line_6[920], line_5[918], line_4[916], line_3[914], line_2[912], line_1[910], 70'b0};
assign col_1165 = {line_58[1025], line_57[1023], line_56[1021], line_55[1019], line_54[1017], line_53[1015], line_52[1013], line_51[1011], line_50[1009], line_49[1007], line_48[1005], line_47[1003], line_46[1001], line_45[999], line_44[997], line_43[995], line_42[993], line_41[991], line_40[989], line_39[987], line_38[985], line_37[983], line_36[981], line_35[979], line_34[977], line_33[975], line_32[973], line_31[971], line_30[969], line_29[967], line_28[965], line_27[963], line_26[961], line_25[959], line_24[957], line_23[955], line_22[953], line_21[951], line_20[949], line_19[947], line_18[945], line_17[943], line_16[941], line_15[939], line_14[937], line_13[935], line_12[933], line_11[931], line_10[929], line_9[927], line_8[925], line_7[923], line_6[921], line_5[919], line_4[917], line_3[915], line_2[913], line_1[911], 70'b0};
assign col_1166 = {line_57[1024], line_56[1022], line_55[1020], line_54[1018], line_53[1016], line_52[1014], line_51[1012], line_50[1010], line_49[1008], line_48[1006], line_47[1004], line_46[1002], line_45[1000], line_44[998], line_43[996], line_42[994], line_41[992], line_40[990], line_39[988], line_38[986], line_37[984], line_36[982], line_35[980], line_34[978], line_33[976], line_32[974], line_31[972], line_30[970], line_29[968], line_28[966], line_27[964], line_26[962], line_25[960], line_24[958], line_23[956], line_22[954], line_21[952], line_20[950], line_19[948], line_18[946], line_17[944], line_16[942], line_15[940], line_14[938], line_13[936], line_12[934], line_11[932], line_10[930], line_9[928], line_8[926], line_7[924], line_6[922], line_5[920], line_4[918], line_3[916], line_2[914], line_1[912], 71'b0};
assign col_1167 = {line_57[1025], line_56[1023], line_55[1021], line_54[1019], line_53[1017], line_52[1015], line_51[1013], line_50[1011], line_49[1009], line_48[1007], line_47[1005], line_46[1003], line_45[1001], line_44[999], line_43[997], line_42[995], line_41[993], line_40[991], line_39[989], line_38[987], line_37[985], line_36[983], line_35[981], line_34[979], line_33[977], line_32[975], line_31[973], line_30[971], line_29[969], line_28[967], line_27[965], line_26[963], line_25[961], line_24[959], line_23[957], line_22[955], line_21[953], line_20[951], line_19[949], line_18[947], line_17[945], line_16[943], line_15[941], line_14[939], line_13[937], line_12[935], line_11[933], line_10[931], line_9[929], line_8[927], line_7[925], line_6[923], line_5[921], line_4[919], line_3[917], line_2[915], line_1[913], 71'b0};
assign col_1168 = {line_56[1024], line_55[1022], line_54[1020], line_53[1018], line_52[1016], line_51[1014], line_50[1012], line_49[1010], line_48[1008], line_47[1006], line_46[1004], line_45[1002], line_44[1000], line_43[998], line_42[996], line_41[994], line_40[992], line_39[990], line_38[988], line_37[986], line_36[984], line_35[982], line_34[980], line_33[978], line_32[976], line_31[974], line_30[972], line_29[970], line_28[968], line_27[966], line_26[964], line_25[962], line_24[960], line_23[958], line_22[956], line_21[954], line_20[952], line_19[950], line_18[948], line_17[946], line_16[944], line_15[942], line_14[940], line_13[938], line_12[936], line_11[934], line_10[932], line_9[930], line_8[928], line_7[926], line_6[924], line_5[922], line_4[920], line_3[918], line_2[916], line_1[914], 72'b0};
assign col_1169 = {line_56[1025], line_55[1023], line_54[1021], line_53[1019], line_52[1017], line_51[1015], line_50[1013], line_49[1011], line_48[1009], line_47[1007], line_46[1005], line_45[1003], line_44[1001], line_43[999], line_42[997], line_41[995], line_40[993], line_39[991], line_38[989], line_37[987], line_36[985], line_35[983], line_34[981], line_33[979], line_32[977], line_31[975], line_30[973], line_29[971], line_28[969], line_27[967], line_26[965], line_25[963], line_24[961], line_23[959], line_22[957], line_21[955], line_20[953], line_19[951], line_18[949], line_17[947], line_16[945], line_15[943], line_14[941], line_13[939], line_12[937], line_11[935], line_10[933], line_9[931], line_8[929], line_7[927], line_6[925], line_5[923], line_4[921], line_3[919], line_2[917], line_1[915], 72'b0};
assign col_1170 = {line_55[1024], line_54[1022], line_53[1020], line_52[1018], line_51[1016], line_50[1014], line_49[1012], line_48[1010], line_47[1008], line_46[1006], line_45[1004], line_44[1002], line_43[1000], line_42[998], line_41[996], line_40[994], line_39[992], line_38[990], line_37[988], line_36[986], line_35[984], line_34[982], line_33[980], line_32[978], line_31[976], line_30[974], line_29[972], line_28[970], line_27[968], line_26[966], line_25[964], line_24[962], line_23[960], line_22[958], line_21[956], line_20[954], line_19[952], line_18[950], line_17[948], line_16[946], line_15[944], line_14[942], line_13[940], line_12[938], line_11[936], line_10[934], line_9[932], line_8[930], line_7[928], line_6[926], line_5[924], line_4[922], line_3[920], line_2[918], line_1[916], 73'b0};
assign col_1171 = {line_55[1025], line_54[1023], line_53[1021], line_52[1019], line_51[1017], line_50[1015], line_49[1013], line_48[1011], line_47[1009], line_46[1007], line_45[1005], line_44[1003], line_43[1001], line_42[999], line_41[997], line_40[995], line_39[993], line_38[991], line_37[989], line_36[987], line_35[985], line_34[983], line_33[981], line_32[979], line_31[977], line_30[975], line_29[973], line_28[971], line_27[969], line_26[967], line_25[965], line_24[963], line_23[961], line_22[959], line_21[957], line_20[955], line_19[953], line_18[951], line_17[949], line_16[947], line_15[945], line_14[943], line_13[941], line_12[939], line_11[937], line_10[935], line_9[933], line_8[931], line_7[929], line_6[927], line_5[925], line_4[923], line_3[921], line_2[919], line_1[917], 73'b0};
assign col_1172 = {line_54[1024], line_53[1022], line_52[1020], line_51[1018], line_50[1016], line_49[1014], line_48[1012], line_47[1010], line_46[1008], line_45[1006], line_44[1004], line_43[1002], line_42[1000], line_41[998], line_40[996], line_39[994], line_38[992], line_37[990], line_36[988], line_35[986], line_34[984], line_33[982], line_32[980], line_31[978], line_30[976], line_29[974], line_28[972], line_27[970], line_26[968], line_25[966], line_24[964], line_23[962], line_22[960], line_21[958], line_20[956], line_19[954], line_18[952], line_17[950], line_16[948], line_15[946], line_14[944], line_13[942], line_12[940], line_11[938], line_10[936], line_9[934], line_8[932], line_7[930], line_6[928], line_5[926], line_4[924], line_3[922], line_2[920], line_1[918], 74'b0};
assign col_1173 = {line_54[1025], line_53[1023], line_52[1021], line_51[1019], line_50[1017], line_49[1015], line_48[1013], line_47[1011], line_46[1009], line_45[1007], line_44[1005], line_43[1003], line_42[1001], line_41[999], line_40[997], line_39[995], line_38[993], line_37[991], line_36[989], line_35[987], line_34[985], line_33[983], line_32[981], line_31[979], line_30[977], line_29[975], line_28[973], line_27[971], line_26[969], line_25[967], line_24[965], line_23[963], line_22[961], line_21[959], line_20[957], line_19[955], line_18[953], line_17[951], line_16[949], line_15[947], line_14[945], line_13[943], line_12[941], line_11[939], line_10[937], line_9[935], line_8[933], line_7[931], line_6[929], line_5[927], line_4[925], line_3[923], line_2[921], line_1[919], 74'b0};
assign col_1174 = {line_53[1024], line_52[1022], line_51[1020], line_50[1018], line_49[1016], line_48[1014], line_47[1012], line_46[1010], line_45[1008], line_44[1006], line_43[1004], line_42[1002], line_41[1000], line_40[998], line_39[996], line_38[994], line_37[992], line_36[990], line_35[988], line_34[986], line_33[984], line_32[982], line_31[980], line_30[978], line_29[976], line_28[974], line_27[972], line_26[970], line_25[968], line_24[966], line_23[964], line_22[962], line_21[960], line_20[958], line_19[956], line_18[954], line_17[952], line_16[950], line_15[948], line_14[946], line_13[944], line_12[942], line_11[940], line_10[938], line_9[936], line_8[934], line_7[932], line_6[930], line_5[928], line_4[926], line_3[924], line_2[922], line_1[920], 75'b0};
assign col_1175 = {line_53[1025], line_52[1023], line_51[1021], line_50[1019], line_49[1017], line_48[1015], line_47[1013], line_46[1011], line_45[1009], line_44[1007], line_43[1005], line_42[1003], line_41[1001], line_40[999], line_39[997], line_38[995], line_37[993], line_36[991], line_35[989], line_34[987], line_33[985], line_32[983], line_31[981], line_30[979], line_29[977], line_28[975], line_27[973], line_26[971], line_25[969], line_24[967], line_23[965], line_22[963], line_21[961], line_20[959], line_19[957], line_18[955], line_17[953], line_16[951], line_15[949], line_14[947], line_13[945], line_12[943], line_11[941], line_10[939], line_9[937], line_8[935], line_7[933], line_6[931], line_5[929], line_4[927], line_3[925], line_2[923], line_1[921], 75'b0};
assign col_1176 = {line_52[1024], line_51[1022], line_50[1020], line_49[1018], line_48[1016], line_47[1014], line_46[1012], line_45[1010], line_44[1008], line_43[1006], line_42[1004], line_41[1002], line_40[1000], line_39[998], line_38[996], line_37[994], line_36[992], line_35[990], line_34[988], line_33[986], line_32[984], line_31[982], line_30[980], line_29[978], line_28[976], line_27[974], line_26[972], line_25[970], line_24[968], line_23[966], line_22[964], line_21[962], line_20[960], line_19[958], line_18[956], line_17[954], line_16[952], line_15[950], line_14[948], line_13[946], line_12[944], line_11[942], line_10[940], line_9[938], line_8[936], line_7[934], line_6[932], line_5[930], line_4[928], line_3[926], line_2[924], line_1[922], 76'b0};
assign col_1177 = {line_52[1025], line_51[1023], line_50[1021], line_49[1019], line_48[1017], line_47[1015], line_46[1013], line_45[1011], line_44[1009], line_43[1007], line_42[1005], line_41[1003], line_40[1001], line_39[999], line_38[997], line_37[995], line_36[993], line_35[991], line_34[989], line_33[987], line_32[985], line_31[983], line_30[981], line_29[979], line_28[977], line_27[975], line_26[973], line_25[971], line_24[969], line_23[967], line_22[965], line_21[963], line_20[961], line_19[959], line_18[957], line_17[955], line_16[953], line_15[951], line_14[949], line_13[947], line_12[945], line_11[943], line_10[941], line_9[939], line_8[937], line_7[935], line_6[933], line_5[931], line_4[929], line_3[927], line_2[925], line_1[923], 76'b0};
assign col_1178 = {line_51[1024], line_50[1022], line_49[1020], line_48[1018], line_47[1016], line_46[1014], line_45[1012], line_44[1010], line_43[1008], line_42[1006], line_41[1004], line_40[1002], line_39[1000], line_38[998], line_37[996], line_36[994], line_35[992], line_34[990], line_33[988], line_32[986], line_31[984], line_30[982], line_29[980], line_28[978], line_27[976], line_26[974], line_25[972], line_24[970], line_23[968], line_22[966], line_21[964], line_20[962], line_19[960], line_18[958], line_17[956], line_16[954], line_15[952], line_14[950], line_13[948], line_12[946], line_11[944], line_10[942], line_9[940], line_8[938], line_7[936], line_6[934], line_5[932], line_4[930], line_3[928], line_2[926], line_1[924], 77'b0};
assign col_1179 = {line_51[1025], line_50[1023], line_49[1021], line_48[1019], line_47[1017], line_46[1015], line_45[1013], line_44[1011], line_43[1009], line_42[1007], line_41[1005], line_40[1003], line_39[1001], line_38[999], line_37[997], line_36[995], line_35[993], line_34[991], line_33[989], line_32[987], line_31[985], line_30[983], line_29[981], line_28[979], line_27[977], line_26[975], line_25[973], line_24[971], line_23[969], line_22[967], line_21[965], line_20[963], line_19[961], line_18[959], line_17[957], line_16[955], line_15[953], line_14[951], line_13[949], line_12[947], line_11[945], line_10[943], line_9[941], line_8[939], line_7[937], line_6[935], line_5[933], line_4[931], line_3[929], line_2[927], line_1[925], 77'b0};
assign col_1180 = {line_50[1024], line_49[1022], line_48[1020], line_47[1018], line_46[1016], line_45[1014], line_44[1012], line_43[1010], line_42[1008], line_41[1006], line_40[1004], line_39[1002], line_38[1000], line_37[998], line_36[996], line_35[994], line_34[992], line_33[990], line_32[988], line_31[986], line_30[984], line_29[982], line_28[980], line_27[978], line_26[976], line_25[974], line_24[972], line_23[970], line_22[968], line_21[966], line_20[964], line_19[962], line_18[960], line_17[958], line_16[956], line_15[954], line_14[952], line_13[950], line_12[948], line_11[946], line_10[944], line_9[942], line_8[940], line_7[938], line_6[936], line_5[934], line_4[932], line_3[930], line_2[928], line_1[926], 78'b0};
assign col_1181 = {line_50[1025], line_49[1023], line_48[1021], line_47[1019], line_46[1017], line_45[1015], line_44[1013], line_43[1011], line_42[1009], line_41[1007], line_40[1005], line_39[1003], line_38[1001], line_37[999], line_36[997], line_35[995], line_34[993], line_33[991], line_32[989], line_31[987], line_30[985], line_29[983], line_28[981], line_27[979], line_26[977], line_25[975], line_24[973], line_23[971], line_22[969], line_21[967], line_20[965], line_19[963], line_18[961], line_17[959], line_16[957], line_15[955], line_14[953], line_13[951], line_12[949], line_11[947], line_10[945], line_9[943], line_8[941], line_7[939], line_6[937], line_5[935], line_4[933], line_3[931], line_2[929], line_1[927], 78'b0};
assign col_1182 = {line_49[1024], line_48[1022], line_47[1020], line_46[1018], line_45[1016], line_44[1014], line_43[1012], line_42[1010], line_41[1008], line_40[1006], line_39[1004], line_38[1002], line_37[1000], line_36[998], line_35[996], line_34[994], line_33[992], line_32[990], line_31[988], line_30[986], line_29[984], line_28[982], line_27[980], line_26[978], line_25[976], line_24[974], line_23[972], line_22[970], line_21[968], line_20[966], line_19[964], line_18[962], line_17[960], line_16[958], line_15[956], line_14[954], line_13[952], line_12[950], line_11[948], line_10[946], line_9[944], line_8[942], line_7[940], line_6[938], line_5[936], line_4[934], line_3[932], line_2[930], line_1[928], 79'b0};
assign col_1183 = {line_49[1025], line_48[1023], line_47[1021], line_46[1019], line_45[1017], line_44[1015], line_43[1013], line_42[1011], line_41[1009], line_40[1007], line_39[1005], line_38[1003], line_37[1001], line_36[999], line_35[997], line_34[995], line_33[993], line_32[991], line_31[989], line_30[987], line_29[985], line_28[983], line_27[981], line_26[979], line_25[977], line_24[975], line_23[973], line_22[971], line_21[969], line_20[967], line_19[965], line_18[963], line_17[961], line_16[959], line_15[957], line_14[955], line_13[953], line_12[951], line_11[949], line_10[947], line_9[945], line_8[943], line_7[941], line_6[939], line_5[937], line_4[935], line_3[933], line_2[931], line_1[929], 79'b0};
assign col_1184 = {line_48[1024], line_47[1022], line_46[1020], line_45[1018], line_44[1016], line_43[1014], line_42[1012], line_41[1010], line_40[1008], line_39[1006], line_38[1004], line_37[1002], line_36[1000], line_35[998], line_34[996], line_33[994], line_32[992], line_31[990], line_30[988], line_29[986], line_28[984], line_27[982], line_26[980], line_25[978], line_24[976], line_23[974], line_22[972], line_21[970], line_20[968], line_19[966], line_18[964], line_17[962], line_16[960], line_15[958], line_14[956], line_13[954], line_12[952], line_11[950], line_10[948], line_9[946], line_8[944], line_7[942], line_6[940], line_5[938], line_4[936], line_3[934], line_2[932], line_1[930], 80'b0};
assign col_1185 = {line_48[1025], line_47[1023], line_46[1021], line_45[1019], line_44[1017], line_43[1015], line_42[1013], line_41[1011], line_40[1009], line_39[1007], line_38[1005], line_37[1003], line_36[1001], line_35[999], line_34[997], line_33[995], line_32[993], line_31[991], line_30[989], line_29[987], line_28[985], line_27[983], line_26[981], line_25[979], line_24[977], line_23[975], line_22[973], line_21[971], line_20[969], line_19[967], line_18[965], line_17[963], line_16[961], line_15[959], line_14[957], line_13[955], line_12[953], line_11[951], line_10[949], line_9[947], line_8[945], line_7[943], line_6[941], line_5[939], line_4[937], line_3[935], line_2[933], line_1[931], 80'b0};
assign col_1186 = {line_47[1024], line_46[1022], line_45[1020], line_44[1018], line_43[1016], line_42[1014], line_41[1012], line_40[1010], line_39[1008], line_38[1006], line_37[1004], line_36[1002], line_35[1000], line_34[998], line_33[996], line_32[994], line_31[992], line_30[990], line_29[988], line_28[986], line_27[984], line_26[982], line_25[980], line_24[978], line_23[976], line_22[974], line_21[972], line_20[970], line_19[968], line_18[966], line_17[964], line_16[962], line_15[960], line_14[958], line_13[956], line_12[954], line_11[952], line_10[950], line_9[948], line_8[946], line_7[944], line_6[942], line_5[940], line_4[938], line_3[936], line_2[934], line_1[932], 81'b0};
assign col_1187 = {line_47[1025], line_46[1023], line_45[1021], line_44[1019], line_43[1017], line_42[1015], line_41[1013], line_40[1011], line_39[1009], line_38[1007], line_37[1005], line_36[1003], line_35[1001], line_34[999], line_33[997], line_32[995], line_31[993], line_30[991], line_29[989], line_28[987], line_27[985], line_26[983], line_25[981], line_24[979], line_23[977], line_22[975], line_21[973], line_20[971], line_19[969], line_18[967], line_17[965], line_16[963], line_15[961], line_14[959], line_13[957], line_12[955], line_11[953], line_10[951], line_9[949], line_8[947], line_7[945], line_6[943], line_5[941], line_4[939], line_3[937], line_2[935], line_1[933], 81'b0};
assign col_1188 = {line_46[1024], line_45[1022], line_44[1020], line_43[1018], line_42[1016], line_41[1014], line_40[1012], line_39[1010], line_38[1008], line_37[1006], line_36[1004], line_35[1002], line_34[1000], line_33[998], line_32[996], line_31[994], line_30[992], line_29[990], line_28[988], line_27[986], line_26[984], line_25[982], line_24[980], line_23[978], line_22[976], line_21[974], line_20[972], line_19[970], line_18[968], line_17[966], line_16[964], line_15[962], line_14[960], line_13[958], line_12[956], line_11[954], line_10[952], line_9[950], line_8[948], line_7[946], line_6[944], line_5[942], line_4[940], line_3[938], line_2[936], line_1[934], 82'b0};
assign col_1189 = {line_46[1025], line_45[1023], line_44[1021], line_43[1019], line_42[1017], line_41[1015], line_40[1013], line_39[1011], line_38[1009], line_37[1007], line_36[1005], line_35[1003], line_34[1001], line_33[999], line_32[997], line_31[995], line_30[993], line_29[991], line_28[989], line_27[987], line_26[985], line_25[983], line_24[981], line_23[979], line_22[977], line_21[975], line_20[973], line_19[971], line_18[969], line_17[967], line_16[965], line_15[963], line_14[961], line_13[959], line_12[957], line_11[955], line_10[953], line_9[951], line_8[949], line_7[947], line_6[945], line_5[943], line_4[941], line_3[939], line_2[937], line_1[935], 82'b0};
assign col_1190 = {line_45[1024], line_44[1022], line_43[1020], line_42[1018], line_41[1016], line_40[1014], line_39[1012], line_38[1010], line_37[1008], line_36[1006], line_35[1004], line_34[1002], line_33[1000], line_32[998], line_31[996], line_30[994], line_29[992], line_28[990], line_27[988], line_26[986], line_25[984], line_24[982], line_23[980], line_22[978], line_21[976], line_20[974], line_19[972], line_18[970], line_17[968], line_16[966], line_15[964], line_14[962], line_13[960], line_12[958], line_11[956], line_10[954], line_9[952], line_8[950], line_7[948], line_6[946], line_5[944], line_4[942], line_3[940], line_2[938], line_1[936], 83'b0};
assign col_1191 = {line_45[1025], line_44[1023], line_43[1021], line_42[1019], line_41[1017], line_40[1015], line_39[1013], line_38[1011], line_37[1009], line_36[1007], line_35[1005], line_34[1003], line_33[1001], line_32[999], line_31[997], line_30[995], line_29[993], line_28[991], line_27[989], line_26[987], line_25[985], line_24[983], line_23[981], line_22[979], line_21[977], line_20[975], line_19[973], line_18[971], line_17[969], line_16[967], line_15[965], line_14[963], line_13[961], line_12[959], line_11[957], line_10[955], line_9[953], line_8[951], line_7[949], line_6[947], line_5[945], line_4[943], line_3[941], line_2[939], line_1[937], 83'b0};
assign col_1192 = {line_44[1024], line_43[1022], line_42[1020], line_41[1018], line_40[1016], line_39[1014], line_38[1012], line_37[1010], line_36[1008], line_35[1006], line_34[1004], line_33[1002], line_32[1000], line_31[998], line_30[996], line_29[994], line_28[992], line_27[990], line_26[988], line_25[986], line_24[984], line_23[982], line_22[980], line_21[978], line_20[976], line_19[974], line_18[972], line_17[970], line_16[968], line_15[966], line_14[964], line_13[962], line_12[960], line_11[958], line_10[956], line_9[954], line_8[952], line_7[950], line_6[948], line_5[946], line_4[944], line_3[942], line_2[940], line_1[938], 84'b0};
assign col_1193 = {line_44[1025], line_43[1023], line_42[1021], line_41[1019], line_40[1017], line_39[1015], line_38[1013], line_37[1011], line_36[1009], line_35[1007], line_34[1005], line_33[1003], line_32[1001], line_31[999], line_30[997], line_29[995], line_28[993], line_27[991], line_26[989], line_25[987], line_24[985], line_23[983], line_22[981], line_21[979], line_20[977], line_19[975], line_18[973], line_17[971], line_16[969], line_15[967], line_14[965], line_13[963], line_12[961], line_11[959], line_10[957], line_9[955], line_8[953], line_7[951], line_6[949], line_5[947], line_4[945], line_3[943], line_2[941], line_1[939], 84'b0};
assign col_1194 = {line_43[1024], line_42[1022], line_41[1020], line_40[1018], line_39[1016], line_38[1014], line_37[1012], line_36[1010], line_35[1008], line_34[1006], line_33[1004], line_32[1002], line_31[1000], line_30[998], line_29[996], line_28[994], line_27[992], line_26[990], line_25[988], line_24[986], line_23[984], line_22[982], line_21[980], line_20[978], line_19[976], line_18[974], line_17[972], line_16[970], line_15[968], line_14[966], line_13[964], line_12[962], line_11[960], line_10[958], line_9[956], line_8[954], line_7[952], line_6[950], line_5[948], line_4[946], line_3[944], line_2[942], line_1[940], 85'b0};
assign col_1195 = {line_43[1025], line_42[1023], line_41[1021], line_40[1019], line_39[1017], line_38[1015], line_37[1013], line_36[1011], line_35[1009], line_34[1007], line_33[1005], line_32[1003], line_31[1001], line_30[999], line_29[997], line_28[995], line_27[993], line_26[991], line_25[989], line_24[987], line_23[985], line_22[983], line_21[981], line_20[979], line_19[977], line_18[975], line_17[973], line_16[971], line_15[969], line_14[967], line_13[965], line_12[963], line_11[961], line_10[959], line_9[957], line_8[955], line_7[953], line_6[951], line_5[949], line_4[947], line_3[945], line_2[943], line_1[941], 85'b0};
assign col_1196 = {line_42[1024], line_41[1022], line_40[1020], line_39[1018], line_38[1016], line_37[1014], line_36[1012], line_35[1010], line_34[1008], line_33[1006], line_32[1004], line_31[1002], line_30[1000], line_29[998], line_28[996], line_27[994], line_26[992], line_25[990], line_24[988], line_23[986], line_22[984], line_21[982], line_20[980], line_19[978], line_18[976], line_17[974], line_16[972], line_15[970], line_14[968], line_13[966], line_12[964], line_11[962], line_10[960], line_9[958], line_8[956], line_7[954], line_6[952], line_5[950], line_4[948], line_3[946], line_2[944], line_1[942], 86'b0};
assign col_1197 = {line_42[1025], line_41[1023], line_40[1021], line_39[1019], line_38[1017], line_37[1015], line_36[1013], line_35[1011], line_34[1009], line_33[1007], line_32[1005], line_31[1003], line_30[1001], line_29[999], line_28[997], line_27[995], line_26[993], line_25[991], line_24[989], line_23[987], line_22[985], line_21[983], line_20[981], line_19[979], line_18[977], line_17[975], line_16[973], line_15[971], line_14[969], line_13[967], line_12[965], line_11[963], line_10[961], line_9[959], line_8[957], line_7[955], line_6[953], line_5[951], line_4[949], line_3[947], line_2[945], line_1[943], 86'b0};
assign col_1198 = {line_41[1024], line_40[1022], line_39[1020], line_38[1018], line_37[1016], line_36[1014], line_35[1012], line_34[1010], line_33[1008], line_32[1006], line_31[1004], line_30[1002], line_29[1000], line_28[998], line_27[996], line_26[994], line_25[992], line_24[990], line_23[988], line_22[986], line_21[984], line_20[982], line_19[980], line_18[978], line_17[976], line_16[974], line_15[972], line_14[970], line_13[968], line_12[966], line_11[964], line_10[962], line_9[960], line_8[958], line_7[956], line_6[954], line_5[952], line_4[950], line_3[948], line_2[946], line_1[944], 87'b0};
assign col_1199 = {line_41[1025], line_40[1023], line_39[1021], line_38[1019], line_37[1017], line_36[1015], line_35[1013], line_34[1011], line_33[1009], line_32[1007], line_31[1005], line_30[1003], line_29[1001], line_28[999], line_27[997], line_26[995], line_25[993], line_24[991], line_23[989], line_22[987], line_21[985], line_20[983], line_19[981], line_18[979], line_17[977], line_16[975], line_15[973], line_14[971], line_13[969], line_12[967], line_11[965], line_10[963], line_9[961], line_8[959], line_7[957], line_6[955], line_5[953], line_4[951], line_3[949], line_2[947], line_1[945], 87'b0};
assign col_1200 = {line_40[1024], line_39[1022], line_38[1020], line_37[1018], line_36[1016], line_35[1014], line_34[1012], line_33[1010], line_32[1008], line_31[1006], line_30[1004], line_29[1002], line_28[1000], line_27[998], line_26[996], line_25[994], line_24[992], line_23[990], line_22[988], line_21[986], line_20[984], line_19[982], line_18[980], line_17[978], line_16[976], line_15[974], line_14[972], line_13[970], line_12[968], line_11[966], line_10[964], line_9[962], line_8[960], line_7[958], line_6[956], line_5[954], line_4[952], line_3[950], line_2[948], line_1[946], 88'b0};
assign col_1201 = {line_40[1025], line_39[1023], line_38[1021], line_37[1019], line_36[1017], line_35[1015], line_34[1013], line_33[1011], line_32[1009], line_31[1007], line_30[1005], line_29[1003], line_28[1001], line_27[999], line_26[997], line_25[995], line_24[993], line_23[991], line_22[989], line_21[987], line_20[985], line_19[983], line_18[981], line_17[979], line_16[977], line_15[975], line_14[973], line_13[971], line_12[969], line_11[967], line_10[965], line_9[963], line_8[961], line_7[959], line_6[957], line_5[955], line_4[953], line_3[951], line_2[949], line_1[947], 88'b0};
assign col_1202 = {line_39[1024], line_38[1022], line_37[1020], line_36[1018], line_35[1016], line_34[1014], line_33[1012], line_32[1010], line_31[1008], line_30[1006], line_29[1004], line_28[1002], line_27[1000], line_26[998], line_25[996], line_24[994], line_23[992], line_22[990], line_21[988], line_20[986], line_19[984], line_18[982], line_17[980], line_16[978], line_15[976], line_14[974], line_13[972], line_12[970], line_11[968], line_10[966], line_9[964], line_8[962], line_7[960], line_6[958], line_5[956], line_4[954], line_3[952], line_2[950], line_1[948], 89'b0};
assign col_1203 = {line_39[1025], line_38[1023], line_37[1021], line_36[1019], line_35[1017], line_34[1015], line_33[1013], line_32[1011], line_31[1009], line_30[1007], line_29[1005], line_28[1003], line_27[1001], line_26[999], line_25[997], line_24[995], line_23[993], line_22[991], line_21[989], line_20[987], line_19[985], line_18[983], line_17[981], line_16[979], line_15[977], line_14[975], line_13[973], line_12[971], line_11[969], line_10[967], line_9[965], line_8[963], line_7[961], line_6[959], line_5[957], line_4[955], line_3[953], line_2[951], line_1[949], 89'b0};
assign col_1204 = {line_38[1024], line_37[1022], line_36[1020], line_35[1018], line_34[1016], line_33[1014], line_32[1012], line_31[1010], line_30[1008], line_29[1006], line_28[1004], line_27[1002], line_26[1000], line_25[998], line_24[996], line_23[994], line_22[992], line_21[990], line_20[988], line_19[986], line_18[984], line_17[982], line_16[980], line_15[978], line_14[976], line_13[974], line_12[972], line_11[970], line_10[968], line_9[966], line_8[964], line_7[962], line_6[960], line_5[958], line_4[956], line_3[954], line_2[952], line_1[950], 90'b0};
assign col_1205 = {line_38[1025], line_37[1023], line_36[1021], line_35[1019], line_34[1017], line_33[1015], line_32[1013], line_31[1011], line_30[1009], line_29[1007], line_28[1005], line_27[1003], line_26[1001], line_25[999], line_24[997], line_23[995], line_22[993], line_21[991], line_20[989], line_19[987], line_18[985], line_17[983], line_16[981], line_15[979], line_14[977], line_13[975], line_12[973], line_11[971], line_10[969], line_9[967], line_8[965], line_7[963], line_6[961], line_5[959], line_4[957], line_3[955], line_2[953], line_1[951], 90'b0};
assign col_1206 = {line_37[1024], line_36[1022], line_35[1020], line_34[1018], line_33[1016], line_32[1014], line_31[1012], line_30[1010], line_29[1008], line_28[1006], line_27[1004], line_26[1002], line_25[1000], line_24[998], line_23[996], line_22[994], line_21[992], line_20[990], line_19[988], line_18[986], line_17[984], line_16[982], line_15[980], line_14[978], line_13[976], line_12[974], line_11[972], line_10[970], line_9[968], line_8[966], line_7[964], line_6[962], line_5[960], line_4[958], line_3[956], line_2[954], line_1[952], 91'b0};
assign col_1207 = {line_37[1025], line_36[1023], line_35[1021], line_34[1019], line_33[1017], line_32[1015], line_31[1013], line_30[1011], line_29[1009], line_28[1007], line_27[1005], line_26[1003], line_25[1001], line_24[999], line_23[997], line_22[995], line_21[993], line_20[991], line_19[989], line_18[987], line_17[985], line_16[983], line_15[981], line_14[979], line_13[977], line_12[975], line_11[973], line_10[971], line_9[969], line_8[967], line_7[965], line_6[963], line_5[961], line_4[959], line_3[957], line_2[955], line_1[953], 91'b0};
assign col_1208 = {line_36[1024], line_35[1022], line_34[1020], line_33[1018], line_32[1016], line_31[1014], line_30[1012], line_29[1010], line_28[1008], line_27[1006], line_26[1004], line_25[1002], line_24[1000], line_23[998], line_22[996], line_21[994], line_20[992], line_19[990], line_18[988], line_17[986], line_16[984], line_15[982], line_14[980], line_13[978], line_12[976], line_11[974], line_10[972], line_9[970], line_8[968], line_7[966], line_6[964], line_5[962], line_4[960], line_3[958], line_2[956], line_1[954], 92'b0};
assign col_1209 = {line_36[1025], line_35[1023], line_34[1021], line_33[1019], line_32[1017], line_31[1015], line_30[1013], line_29[1011], line_28[1009], line_27[1007], line_26[1005], line_25[1003], line_24[1001], line_23[999], line_22[997], line_21[995], line_20[993], line_19[991], line_18[989], line_17[987], line_16[985], line_15[983], line_14[981], line_13[979], line_12[977], line_11[975], line_10[973], line_9[971], line_8[969], line_7[967], line_6[965], line_5[963], line_4[961], line_3[959], line_2[957], line_1[955], 92'b0};
assign col_1210 = {line_35[1024], line_34[1022], line_33[1020], line_32[1018], line_31[1016], line_30[1014], line_29[1012], line_28[1010], line_27[1008], line_26[1006], line_25[1004], line_24[1002], line_23[1000], line_22[998], line_21[996], line_20[994], line_19[992], line_18[990], line_17[988], line_16[986], line_15[984], line_14[982], line_13[980], line_12[978], line_11[976], line_10[974], line_9[972], line_8[970], line_7[968], line_6[966], line_5[964], line_4[962], line_3[960], line_2[958], line_1[956], 93'b0};
assign col_1211 = {line_35[1025], line_34[1023], line_33[1021], line_32[1019], line_31[1017], line_30[1015], line_29[1013], line_28[1011], line_27[1009], line_26[1007], line_25[1005], line_24[1003], line_23[1001], line_22[999], line_21[997], line_20[995], line_19[993], line_18[991], line_17[989], line_16[987], line_15[985], line_14[983], line_13[981], line_12[979], line_11[977], line_10[975], line_9[973], line_8[971], line_7[969], line_6[967], line_5[965], line_4[963], line_3[961], line_2[959], line_1[957], 93'b0};
assign col_1212 = {line_34[1024], line_33[1022], line_32[1020], line_31[1018], line_30[1016], line_29[1014], line_28[1012], line_27[1010], line_26[1008], line_25[1006], line_24[1004], line_23[1002], line_22[1000], line_21[998], line_20[996], line_19[994], line_18[992], line_17[990], line_16[988], line_15[986], line_14[984], line_13[982], line_12[980], line_11[978], line_10[976], line_9[974], line_8[972], line_7[970], line_6[968], line_5[966], line_4[964], line_3[962], line_2[960], line_1[958], 94'b0};
assign col_1213 = {line_34[1025], line_33[1023], line_32[1021], line_31[1019], line_30[1017], line_29[1015], line_28[1013], line_27[1011], line_26[1009], line_25[1007], line_24[1005], line_23[1003], line_22[1001], line_21[999], line_20[997], line_19[995], line_18[993], line_17[991], line_16[989], line_15[987], line_14[985], line_13[983], line_12[981], line_11[979], line_10[977], line_9[975], line_8[973], line_7[971], line_6[969], line_5[967], line_4[965], line_3[963], line_2[961], line_1[959], 94'b0};
assign col_1214 = {line_33[1024], line_32[1022], line_31[1020], line_30[1018], line_29[1016], line_28[1014], line_27[1012], line_26[1010], line_25[1008], line_24[1006], line_23[1004], line_22[1002], line_21[1000], line_20[998], line_19[996], line_18[994], line_17[992], line_16[990], line_15[988], line_14[986], line_13[984], line_12[982], line_11[980], line_10[978], line_9[976], line_8[974], line_7[972], line_6[970], line_5[968], line_4[966], line_3[964], line_2[962], line_1[960], 95'b0};
assign col_1215 = {line_33[1025], line_32[1023], line_31[1021], line_30[1019], line_29[1017], line_28[1015], line_27[1013], line_26[1011], line_25[1009], line_24[1007], line_23[1005], line_22[1003], line_21[1001], line_20[999], line_19[997], line_18[995], line_17[993], line_16[991], line_15[989], line_14[987], line_13[985], line_12[983], line_11[981], line_10[979], line_9[977], line_8[975], line_7[973], line_6[971], line_5[969], line_4[967], line_3[965], line_2[963], line_1[961], 95'b0};
assign col_1216 = {line_32[1024], line_31[1022], line_30[1020], line_29[1018], line_28[1016], line_27[1014], line_26[1012], line_25[1010], line_24[1008], line_23[1006], line_22[1004], line_21[1002], line_20[1000], line_19[998], line_18[996], line_17[994], line_16[992], line_15[990], line_14[988], line_13[986], line_12[984], line_11[982], line_10[980], line_9[978], line_8[976], line_7[974], line_6[972], line_5[970], line_4[968], line_3[966], line_2[964], line_1[962], 96'b0};
assign col_1217 = {line_32[1025], line_31[1023], line_30[1021], line_29[1019], line_28[1017], line_27[1015], line_26[1013], line_25[1011], line_24[1009], line_23[1007], line_22[1005], line_21[1003], line_20[1001], line_19[999], line_18[997], line_17[995], line_16[993], line_15[991], line_14[989], line_13[987], line_12[985], line_11[983], line_10[981], line_9[979], line_8[977], line_7[975], line_6[973], line_5[971], line_4[969], line_3[967], line_2[965], line_1[963], 96'b0};
assign col_1218 = {line_31[1024], line_30[1022], line_29[1020], line_28[1018], line_27[1016], line_26[1014], line_25[1012], line_24[1010], line_23[1008], line_22[1006], line_21[1004], line_20[1002], line_19[1000], line_18[998], line_17[996], line_16[994], line_15[992], line_14[990], line_13[988], line_12[986], line_11[984], line_10[982], line_9[980], line_8[978], line_7[976], line_6[974], line_5[972], line_4[970], line_3[968], line_2[966], line_1[964], 97'b0};
assign col_1219 = {line_31[1025], line_30[1023], line_29[1021], line_28[1019], line_27[1017], line_26[1015], line_25[1013], line_24[1011], line_23[1009], line_22[1007], line_21[1005], line_20[1003], line_19[1001], line_18[999], line_17[997], line_16[995], line_15[993], line_14[991], line_13[989], line_12[987], line_11[985], line_10[983], line_9[981], line_8[979], line_7[977], line_6[975], line_5[973], line_4[971], line_3[969], line_2[967], line_1[965], 97'b0};
assign col_1220 = {line_30[1024], line_29[1022], line_28[1020], line_27[1018], line_26[1016], line_25[1014], line_24[1012], line_23[1010], line_22[1008], line_21[1006], line_20[1004], line_19[1002], line_18[1000], line_17[998], line_16[996], line_15[994], line_14[992], line_13[990], line_12[988], line_11[986], line_10[984], line_9[982], line_8[980], line_7[978], line_6[976], line_5[974], line_4[972], line_3[970], line_2[968], line_1[966], 98'b0};
assign col_1221 = {line_30[1025], line_29[1023], line_28[1021], line_27[1019], line_26[1017], line_25[1015], line_24[1013], line_23[1011], line_22[1009], line_21[1007], line_20[1005], line_19[1003], line_18[1001], line_17[999], line_16[997], line_15[995], line_14[993], line_13[991], line_12[989], line_11[987], line_10[985], line_9[983], line_8[981], line_7[979], line_6[977], line_5[975], line_4[973], line_3[971], line_2[969], line_1[967], 98'b0};
assign col_1222 = {line_29[1024], line_28[1022], line_27[1020], line_26[1018], line_25[1016], line_24[1014], line_23[1012], line_22[1010], line_21[1008], line_20[1006], line_19[1004], line_18[1002], line_17[1000], line_16[998], line_15[996], line_14[994], line_13[992], line_12[990], line_11[988], line_10[986], line_9[984], line_8[982], line_7[980], line_6[978], line_5[976], line_4[974], line_3[972], line_2[970], line_1[968], 99'b0};
assign col_1223 = {line_29[1025], line_28[1023], line_27[1021], line_26[1019], line_25[1017], line_24[1015], line_23[1013], line_22[1011], line_21[1009], line_20[1007], line_19[1005], line_18[1003], line_17[1001], line_16[999], line_15[997], line_14[995], line_13[993], line_12[991], line_11[989], line_10[987], line_9[985], line_8[983], line_7[981], line_6[979], line_5[977], line_4[975], line_3[973], line_2[971], line_1[969], 99'b0};
assign col_1224 = {line_28[1024], line_27[1022], line_26[1020], line_25[1018], line_24[1016], line_23[1014], line_22[1012], line_21[1010], line_20[1008], line_19[1006], line_18[1004], line_17[1002], line_16[1000], line_15[998], line_14[996], line_13[994], line_12[992], line_11[990], line_10[988], line_9[986], line_8[984], line_7[982], line_6[980], line_5[978], line_4[976], line_3[974], line_2[972], line_1[970], 100'b0};
assign col_1225 = {line_28[1025], line_27[1023], line_26[1021], line_25[1019], line_24[1017], line_23[1015], line_22[1013], line_21[1011], line_20[1009], line_19[1007], line_18[1005], line_17[1003], line_16[1001], line_15[999], line_14[997], line_13[995], line_12[993], line_11[991], line_10[989], line_9[987], line_8[985], line_7[983], line_6[981], line_5[979], line_4[977], line_3[975], line_2[973], line_1[971], 100'b0};
assign col_1226 = {line_27[1024], line_26[1022], line_25[1020], line_24[1018], line_23[1016], line_22[1014], line_21[1012], line_20[1010], line_19[1008], line_18[1006], line_17[1004], line_16[1002], line_15[1000], line_14[998], line_13[996], line_12[994], line_11[992], line_10[990], line_9[988], line_8[986], line_7[984], line_6[982], line_5[980], line_4[978], line_3[976], line_2[974], line_1[972], 101'b0};
assign col_1227 = {line_27[1025], line_26[1023], line_25[1021], line_24[1019], line_23[1017], line_22[1015], line_21[1013], line_20[1011], line_19[1009], line_18[1007], line_17[1005], line_16[1003], line_15[1001], line_14[999], line_13[997], line_12[995], line_11[993], line_10[991], line_9[989], line_8[987], line_7[985], line_6[983], line_5[981], line_4[979], line_3[977], line_2[975], line_1[973], 101'b0};
assign col_1228 = {line_26[1024], line_25[1022], line_24[1020], line_23[1018], line_22[1016], line_21[1014], line_20[1012], line_19[1010], line_18[1008], line_17[1006], line_16[1004], line_15[1002], line_14[1000], line_13[998], line_12[996], line_11[994], line_10[992], line_9[990], line_8[988], line_7[986], line_6[984], line_5[982], line_4[980], line_3[978], line_2[976], line_1[974], 102'b0};
assign col_1229 = {line_26[1025], line_25[1023], line_24[1021], line_23[1019], line_22[1017], line_21[1015], line_20[1013], line_19[1011], line_18[1009], line_17[1007], line_16[1005], line_15[1003], line_14[1001], line_13[999], line_12[997], line_11[995], line_10[993], line_9[991], line_8[989], line_7[987], line_6[985], line_5[983], line_4[981], line_3[979], line_2[977], line_1[975], 102'b0};
assign col_1230 = {line_25[1024], line_24[1022], line_23[1020], line_22[1018], line_21[1016], line_20[1014], line_19[1012], line_18[1010], line_17[1008], line_16[1006], line_15[1004], line_14[1002], line_13[1000], line_12[998], line_11[996], line_10[994], line_9[992], line_8[990], line_7[988], line_6[986], line_5[984], line_4[982], line_3[980], line_2[978], line_1[976], 103'b0};
assign col_1231 = {line_25[1025], line_24[1023], line_23[1021], line_22[1019], line_21[1017], line_20[1015], line_19[1013], line_18[1011], line_17[1009], line_16[1007], line_15[1005], line_14[1003], line_13[1001], line_12[999], line_11[997], line_10[995], line_9[993], line_8[991], line_7[989], line_6[987], line_5[985], line_4[983], line_3[981], line_2[979], line_1[977], 103'b0};
assign col_1232 = {line_24[1024], line_23[1022], line_22[1020], line_21[1018], line_20[1016], line_19[1014], line_18[1012], line_17[1010], line_16[1008], line_15[1006], line_14[1004], line_13[1002], line_12[1000], line_11[998], line_10[996], line_9[994], line_8[992], line_7[990], line_6[988], line_5[986], line_4[984], line_3[982], line_2[980], line_1[978], 104'b0};
assign col_1233 = {line_24[1025], line_23[1023], line_22[1021], line_21[1019], line_20[1017], line_19[1015], line_18[1013], line_17[1011], line_16[1009], line_15[1007], line_14[1005], line_13[1003], line_12[1001], line_11[999], line_10[997], line_9[995], line_8[993], line_7[991], line_6[989], line_5[987], line_4[985], line_3[983], line_2[981], line_1[979], 104'b0};
assign col_1234 = {line_23[1024], line_22[1022], line_21[1020], line_20[1018], line_19[1016], line_18[1014], line_17[1012], line_16[1010], line_15[1008], line_14[1006], line_13[1004], line_12[1002], line_11[1000], line_10[998], line_9[996], line_8[994], line_7[992], line_6[990], line_5[988], line_4[986], line_3[984], line_2[982], line_1[980], 105'b0};
assign col_1235 = {line_23[1025], line_22[1023], line_21[1021], line_20[1019], line_19[1017], line_18[1015], line_17[1013], line_16[1011], line_15[1009], line_14[1007], line_13[1005], line_12[1003], line_11[1001], line_10[999], line_9[997], line_8[995], line_7[993], line_6[991], line_5[989], line_4[987], line_3[985], line_2[983], line_1[981], 105'b0};
assign col_1236 = {line_22[1024], line_21[1022], line_20[1020], line_19[1018], line_18[1016], line_17[1014], line_16[1012], line_15[1010], line_14[1008], line_13[1006], line_12[1004], line_11[1002], line_10[1000], line_9[998], line_8[996], line_7[994], line_6[992], line_5[990], line_4[988], line_3[986], line_2[984], line_1[982], 106'b0};
assign col_1237 = {line_22[1025], line_21[1023], line_20[1021], line_19[1019], line_18[1017], line_17[1015], line_16[1013], line_15[1011], line_14[1009], line_13[1007], line_12[1005], line_11[1003], line_10[1001], line_9[999], line_8[997], line_7[995], line_6[993], line_5[991], line_4[989], line_3[987], line_2[985], line_1[983], 106'b0};
assign col_1238 = {line_21[1024], line_20[1022], line_19[1020], line_18[1018], line_17[1016], line_16[1014], line_15[1012], line_14[1010], line_13[1008], line_12[1006], line_11[1004], line_10[1002], line_9[1000], line_8[998], line_7[996], line_6[994], line_5[992], line_4[990], line_3[988], line_2[986], line_1[984], 107'b0};
assign col_1239 = {line_21[1025], line_20[1023], line_19[1021], line_18[1019], line_17[1017], line_16[1015], line_15[1013], line_14[1011], line_13[1009], line_12[1007], line_11[1005], line_10[1003], line_9[1001], line_8[999], line_7[997], line_6[995], line_5[993], line_4[991], line_3[989], line_2[987], line_1[985], 107'b0};
assign col_1240 = {line_20[1024], line_19[1022], line_18[1020], line_17[1018], line_16[1016], line_15[1014], line_14[1012], line_13[1010], line_12[1008], line_11[1006], line_10[1004], line_9[1002], line_8[1000], line_7[998], line_6[996], line_5[994], line_4[992], line_3[990], line_2[988], line_1[986], 108'b0};
assign col_1241 = {line_20[1025], line_19[1023], line_18[1021], line_17[1019], line_16[1017], line_15[1015], line_14[1013], line_13[1011], line_12[1009], line_11[1007], line_10[1005], line_9[1003], line_8[1001], line_7[999], line_6[997], line_5[995], line_4[993], line_3[991], line_2[989], line_1[987], 108'b0};
assign col_1242 = {line_19[1024], line_18[1022], line_17[1020], line_16[1018], line_15[1016], line_14[1014], line_13[1012], line_12[1010], line_11[1008], line_10[1006], line_9[1004], line_8[1002], line_7[1000], line_6[998], line_5[996], line_4[994], line_3[992], line_2[990], line_1[988], 109'b0};
assign col_1243 = {line_19[1025], line_18[1023], line_17[1021], line_16[1019], line_15[1017], line_14[1015], line_13[1013], line_12[1011], line_11[1009], line_10[1007], line_9[1005], line_8[1003], line_7[1001], line_6[999], line_5[997], line_4[995], line_3[993], line_2[991], line_1[989], 109'b0};
assign col_1244 = {line_18[1024], line_17[1022], line_16[1020], line_15[1018], line_14[1016], line_13[1014], line_12[1012], line_11[1010], line_10[1008], line_9[1006], line_8[1004], line_7[1002], line_6[1000], line_5[998], line_4[996], line_3[994], line_2[992], line_1[990], 110'b0};
assign col_1245 = {line_18[1025], line_17[1023], line_16[1021], line_15[1019], line_14[1017], line_13[1015], line_12[1013], line_11[1011], line_10[1009], line_9[1007], line_8[1005], line_7[1003], line_6[1001], line_5[999], line_4[997], line_3[995], line_2[993], line_1[991], 110'b0};
assign col_1246 = {line_17[1024], line_16[1022], line_15[1020], line_14[1018], line_13[1016], line_12[1014], line_11[1012], line_10[1010], line_9[1008], line_8[1006], line_7[1004], line_6[1002], line_5[1000], line_4[998], line_3[996], line_2[994], line_1[992], 111'b0};
assign col_1247 = {line_17[1025], line_16[1023], line_15[1021], line_14[1019], line_13[1017], line_12[1015], line_11[1013], line_10[1011], line_9[1009], line_8[1007], line_7[1005], line_6[1003], line_5[1001], line_4[999], line_3[997], line_2[995], line_1[993], 111'b0};
assign col_1248 = {line_16[1024], line_15[1022], line_14[1020], line_13[1018], line_12[1016], line_11[1014], line_10[1012], line_9[1010], line_8[1008], line_7[1006], line_6[1004], line_5[1002], line_4[1000], line_3[998], line_2[996], line_1[994], 112'b0};
assign col_1249 = {line_16[1025], line_15[1023], line_14[1021], line_13[1019], line_12[1017], line_11[1015], line_10[1013], line_9[1011], line_8[1009], line_7[1007], line_6[1005], line_5[1003], line_4[1001], line_3[999], line_2[997], line_1[995], 112'b0};
assign col_1250 = {line_15[1024], line_14[1022], line_13[1020], line_12[1018], line_11[1016], line_10[1014], line_9[1012], line_8[1010], line_7[1008], line_6[1006], line_5[1004], line_4[1002], line_3[1000], line_2[998], line_1[996], 113'b0};
assign col_1251 = {line_15[1025], line_14[1023], line_13[1021], line_12[1019], line_11[1017], line_10[1015], line_9[1013], line_8[1011], line_7[1009], line_6[1007], line_5[1005], line_4[1003], line_3[1001], line_2[999], line_1[997], 113'b0};
assign col_1252 = {line_14[1024], line_13[1022], line_12[1020], line_11[1018], line_10[1016], line_9[1014], line_8[1012], line_7[1010], line_6[1008], line_5[1006], line_4[1004], line_3[1002], line_2[1000], line_1[998], 114'b0};
assign col_1253 = {line_14[1025], line_13[1023], line_12[1021], line_11[1019], line_10[1017], line_9[1015], line_8[1013], line_7[1011], line_6[1009], line_5[1007], line_4[1005], line_3[1003], line_2[1001], line_1[999], 114'b0};
assign col_1254 = {line_13[1024], line_12[1022], line_11[1020], line_10[1018], line_9[1016], line_8[1014], line_7[1012], line_6[1010], line_5[1008], line_4[1006], line_3[1004], line_2[1002], line_1[1000], 115'b0};
assign col_1255 = {line_13[1025], line_12[1023], line_11[1021], line_10[1019], line_9[1017], line_8[1015], line_7[1013], line_6[1011], line_5[1009], line_4[1007], line_3[1005], line_2[1003], line_1[1001], 115'b0};
assign col_1256 = {line_12[1024], line_11[1022], line_10[1020], line_9[1018], line_8[1016], line_7[1014], line_6[1012], line_5[1010], line_4[1008], line_3[1006], line_2[1004], line_1[1002], 116'b0};
assign col_1257 = {line_12[1025], line_11[1023], line_10[1021], line_9[1019], line_8[1017], line_7[1015], line_6[1013], line_5[1011], line_4[1009], line_3[1007], line_2[1005], line_1[1003], 116'b0};
assign col_1258 = {line_11[1024], line_10[1022], line_9[1020], line_8[1018], line_7[1016], line_6[1014], line_5[1012], line_4[1010], line_3[1008], line_2[1006], line_1[1004], 117'b0};
assign col_1259 = {line_11[1025], line_10[1023], line_9[1021], line_8[1019], line_7[1017], line_6[1015], line_5[1013], line_4[1011], line_3[1009], line_2[1007], line_1[1005], 117'b0};
assign col_1260 = {line_10[1024], line_9[1022], line_8[1020], line_7[1018], line_6[1016], line_5[1014], line_4[1012], line_3[1010], line_2[1008], line_1[1006], 118'b0};
assign col_1261 = {line_10[1025], line_9[1023], line_8[1021], line_7[1019], line_6[1017], line_5[1015], line_4[1013], line_3[1011], line_2[1009], line_1[1007], 118'b0};
assign col_1262 = {line_9[1024], line_8[1022], line_7[1020], line_6[1018], line_5[1016], line_4[1014], line_3[1012], line_2[1010], line_1[1008], 119'b0};
assign col_1263 = {line_9[1025], line_8[1023], line_7[1021], line_6[1019], line_5[1017], line_4[1015], line_3[1013], line_2[1011], line_1[1009], 119'b0};
assign col_1264 = {line_8[1024], line_7[1022], line_6[1020], line_5[1018], line_4[1016], line_3[1014], line_2[1012], line_1[1010], 120'b0};
assign col_1265 = {line_8[1025], line_7[1023], line_6[1021], line_5[1019], line_4[1017], line_3[1015], line_2[1013], line_1[1011], 120'b0};
assign col_1266 = {line_7[1024], line_6[1022], line_5[1020], line_4[1018], line_3[1016], line_2[1014], line_1[1012], 121'b0};
assign col_1267 = {line_7[1025], line_6[1023], line_5[1021], line_4[1019], line_3[1017], line_2[1015], line_1[1013], 121'b0};
assign col_1268 = {line_6[1024], line_5[1022], line_4[1020], line_3[1018], line_2[1016], line_1[1014], 122'b0};
assign col_1269 = {line_6[1025], line_5[1023], line_4[1021], line_3[1019], line_2[1017], line_1[1015], 122'b0};
assign col_1270 = {line_5[1024], line_4[1022], line_3[1020], line_2[1018], line_1[1016], 123'b0};
assign col_1271 = {line_5[1025], line_4[1023], line_3[1021], line_2[1019], line_1[1017], 123'b0};
assign col_1272 = {line_4[1024], line_3[1022], line_2[1020], line_1[1018], 124'b0};
assign col_1273 = {line_4[1025], line_3[1023], line_2[1021], line_1[1019], 124'b0};
assign col_1274 = {line_3[1024], line_2[1022], line_1[1020], 125'b0};
assign col_1275 = {line_3[1025], line_2[1023], line_1[1021], 125'b0};
assign col_1276 = {line_2[1024], line_1[1022], 126'b0};
assign col_1277 = {line_2[1025], line_1[1023], 126'b0};
assign col_1278 = {line_1[1024], 127'b0};
assign col_1279 = {line_1[1025], 127'b0};

endmodule

module xpb_5_630
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h997c2b7f61d8ca35fedabd1772e665c0e43b3ed01d7aba6f0f005ab29e1a525758864987b795652ec0936754373c2ba16254acaad6e546bb6a1677303e720030e9281ae4bde97f17d59770f83d242e1e9db29880101394b0181464bdc56254b781af0f3b0872fef7ffff0fb0235c1b9740d9dbffbde40cc9bcd97bdbbe171b34;
    5'b00010 : xpb = 1024'h824b11a901c35fa332b00257d572843057007a6f657dd466a023fc0f8931f7a6adc41596a5044bcee1c88f618b1a4678608f316f8b17bd2b238daf0242118bb05e01011acc4200ea9894df4de16c980c4760376793a0fc4f7a9c3780d09a06dcd4568c4c601d0562793e38814ee8110532d9d91d2b7cbc6333437cb2f34bcffd;
    5'b00011 : xpb = 1024'h6b19f7d2a1adf5106685479837fea29fc9c5b60ead80ee5e31479d6c74499cf60301e1a59273326f02fdb76edef8614f5ec9b6343f4a339add04e6d445b1172fd2d9e750da9a82bd5b924da385b501f9f10dd64f172e63eedd240a43dbd1b90226fe095db7c70bccf27d61527a74067324d9d63a99156bfca9ad7d8a288084c6;
    5'b00100 : xpb = 1024'h53e8ddfc41988a7d9a5a8cd89a8ac10f3c8af1adf5840855c26b3ec95f614245583fadb47fe2190f2432df7c32d67c265d043af8f37caa0a967c1ea64950a2af47b2cd86e8f304901e8fbbf929fd6be79abb75369abbcb8e3fabdd06e7096b2779a5866f0f7112376bbc8a23a5fffbe116d9d35806ae1b9620177e615db5398f;
    5'b00101 : xpb = 1024'h3cb7c425e1831feace2fd218fd16df7eaf502d4d3d87224d538ee0264a78e794ad7d79c36d50ffaf4568078986b496fd5b3ebfbda7af207a4ff356784cf02e2ebc8bb3bcf74b8662e18d2a4ece45d5d54469141e1e49332da233afc9f2411d4ccc4d0380671b18a1e4fbb2f4d18bf14f08d9d0757446cb2f96817f3892e9ee58;
    5'b00110 : xpb = 1024'h2586aa4f816db558020517595fa2fdee221568ec858a3c44e4b2818335908ce402bb45d25abfe64f669d2f96da92b1d4597944825be196ea096a8e4a508fb9ae316499f305a40835a48a98a4728e3fc2ee16b305a1d69acd04bb828cfd78cf721ef48091bec51f0c5e3adbc5fd17e6bcfad9cd92e1df7ac90ceb800fc81ea321;
    5'b00111 : xpb = 1024'he55907921584ac535da5c99c22f1c5d94daa48bcd8d563c75d622e020a8323357f911e1482eccef87d257a42e70ccab57b3c94710140d59c2e1c61c542f452da63d802913fc8a08678806fa16d6a9b097c451ed2564026c6743555008b08197719bfda3166f2576d77a049728a3dc2aecd9cab04f782a62835580e6fd5357ea;
    5'b01000 : xpb = 1024'ha7d1bbf8833114fb34b519b13515821e7915e35beb0810ab84d67d92bec2848ab07f5b68ffc4321e4865bef865acf84cba0875f1e6f954152cf83d4c92a1455e8f659b0dd1e609203d1f77f253fad7cf3576ea6d3577971c7f57ba0dce12d64ef34b0cde1ee2246ed77914474bfff7c22db3a6b00d5c372c402efcc2bb6a731e;
    5'b01001 : xpb = 1024'h90a0a222231baa68688a5ef197a1a08debdb1efb330b2aa315fa1eefa9da29da05bd2777ed3318be699ae705b98b1323b842fab69b2bca84e66f751e9640d0de043e8143e03e8af3001ce647f84341bcdf248954b904febbe1df8cd0d94a887445f289ef768c2ad950b83d18778bed301fb3a3cd7af4e6c5b698fd99f09f27e7;
    5'b01010 : xpb = 1024'h796f884bc3063fd59c5fa431fa2dbefd5ea05a9a7b0e449aa71dc04c94f1cf295afaf386daa1ff5e8ad00f130d692dfab67d7f7b4f5e40f49fe6acf099e05c5d79176779ee970cc5c31a549d9c8babaa88d2283c3c92665b44675f93e4823a99989a0700ce363143c9f765e9a317e29e11b3a0eae88d965f2d02fe7125d3dcb0;
    5'b01011 : xpb = 1024'h623e6e7562f0d542d034e9725cb9dd6cd1659639c3115e92384161a980097478b038bf95c810e5feac053720614748d1b4b804400390b764595de4c29d7fe7dcedf04daffcef8e988617c2f340d41598327fc723c01fcdfaa6ef3256efb9ecbeeb41841225e037ae43368ebacea3d80c03b39e08562645f8a36cff485b089179;
    5'b01100 : xpb = 1024'h4b0d549f02db6ab0040a2eb2bf45fbdc442ad1d90b147889c96503066b2119c805768ba4b57fcc9ecd3a5f2db52563a8b2f28904b7c32dd412d51c94a11f735c62c933e60b48106b49153148e51c7f85dc2d660b43ad359a09770519faf19ee43de901237d8a3e18bc75b78bfa2fcd79f5b39b25c3bef59219d7001f903d4642;
    5'b01101 : xpb = 1024'h33dc3ac8a2c6001d37df73f321d21a4bb6f00d78531792815a88a4635638bf175ab457b3a2eeb33eee6f873b09037e7fb12d0dc96bf5a443cc4c5466a4befedbd7a21a1c19a0923e0c129f9e8964e97385db04f2c73a9d396bfed7dd0629510990907e34d534448335b4e05d25bbc2e7e7b398433157a52b904100f6c571fb0b;
    5'b01110 : xpb = 1024'h1cab20f242b0958a6bb4b933845e38bb29b549179b1aac78ebac45c041506466aff223c2905d99df0fa4af485ce19956af67928e20281ab385c38c38a85e8a5b4c7b005227f91410cf100df42dad53612f88a3da4ac804d8ce86aaa01161032ee337fb462cde4aedaef4092e5147b855d9b395609ef054c506ab01cdfaa6afd4;
    5'b01111 : xpb = 1024'h57a071be29b2af79f89fe73e6ea572a9c7a84b6e31dc6707ccfe71d2c6809b6052fefd17dcc807f30d9d755b0bfb42dada21752d45a91233f3ac40aabfe15dac153e688365195e3920d7c49d1f5bd4ed93642c1ce556c78310e7d631c98b55435df785784885158283331ff7cd3adc3cbb3927e0c89045e7d1502a52fdb649d;
    5'b10000 : xpb = 1024'h9ef6329b4473f52d9e64bb8b59d0bceb80b5c387009880df8bd041cfca825c0d5db639593561e5adf16d3ea9e7fbdfcf0ff6c3fdab3fd7dea9513b3aea70160baa7c016cf43b14fb67a4ed420f19eb6d76e8db41de6901284922e220e1fb0a0bb78e87928cfb5050283241afa02fc95b0c8d6e7dca6d112839ee7e80edf27fd1;
    5'b10001 : xpb = 1024'h87c518c4e45e8a9ad23a00cbbc5cdb5af37aff26489b9ad71cf3e32cb59a015cb2f4056822d0cc4e12a266b73bd9faa60e3148c25f724e4e62c8730cee0fa18b1f54e7a3029396ce2aa25b97b362555b20967a2961f668c7abaab4e3ed32bc310a3604a3e4a556baa1716a80cbbbbec8fe8d6b9b3805c0c1b0587f582327349a;
    5'b10010 : xpb = 1024'h7093feee84492008060f460c1ee8f9ca66403ac5909eb4ceae178489a0b1a6ac0831d177103fb2ee33d78ec48fb8157d0c6bcd8713a4c4be1c3faadef1af2d0a942dcdd910ec18a0ed9fc9ed57aabf48ca441910e583d0670e3287a6f86a6e565cdd81b53c4f5d251ab09351f747b436f08d68b8a59e705b26c2802f585be963;
    5'b10011 : xpb = 1024'h5962e5182433b57539e48b4c81751839d9057664d8a1cec63f3b25e68bc94bfb5d6f9d85fdae998e550cb6d1e39630540aa6524bc7d73b2dd5b6e2b0f54eb88a0906b40f1f449a73b09d3842fbf3293673f1b7f86911380670ba5a6a03a2207baf84fec693f9638f93efbc2322d3a9a4e28d65d613371ff49d2c81068d909e2c;
    5'b10100 : xpb = 1024'h4231cb41c41e4ae26db9d08ce40136a94bcab20420a4e8bdd05ec74376e0f14ab2ad6994eb1d802e7641dedf37744b2b08e0d7107c09b19d8f2e1a82f8ee44097ddf9a452d9d1c46739aa698a03b93241d9f56dfec9e9fa5d3422d2d0ed9d2a1022c7bd7eba369fa0d2ee4f44e5f9f12d48d62f380cfcf8e139681ddc2c552f5;
    5'b10101 : xpb = 1024'h2b00b16b6408e04fa18f15cd468d5518be8feda368a802b5618268a061f8969a07eb35a3d88c66ce977706ec8b526602071b5bd5303c280d48a55254fc8dcf88f2b8807b3bf59e19369814ee4483fd11c74cf5c7702c074535c9fff01a1184c654d3f8e9434d7064866e0dc579eb9480c68d6010ee687f278a0082b4f7fa07be;
    5'b10110 : xpb = 1024'h13cf979503f375bcd5645b0da919738831552942b0ab1cacf2a609fd4d103be95d2901b2c5fb4d6eb8ac2ef9df3080d90555e099e46e9e7d021c8a27002d5b08679166b14a4e1febf9958343e8cc66ff70fa94aef3b96ee49851d2b3254936eba77b75fa9af776ceffad3696a57789eeb88d5d2e5c012ec1006a838c2d2ebc87;
    5'b10111 : xpb = 1024'had4bc31465cc3ff2d43f18251bffd94915906812ce25d71c01a664afeb2a8e40b5af4b3a7d90b29d793f964e166cac7a67aa8d44bb53e5386c3301573e9f5b3950b9819608379f03cf2cf43c25f0951e0ead2d2f03cd0394b0663770eaab8ba3292a8535a36a75c6ffac4646c8d3a585f967392e19e53b8abd43ff67eb45d7bb;
    5'b11000 : xpb = 1024'h961aa93e05b6d56008145d657e8bf7b88855a3b21628f11392ca060cd64233900aed17496aff993d9a74be5b6a4ac75165e512096f865ba825aa3929423ee6b8c59267cc169020d6922a6291ca38ff0bb85acc16875a6b3412ee0a33f5e33dc87bd20246fb147c3178eb6f17f45f9af3eb67364b877deb2433ae003f207a8c84;
    5'b11001 : xpb = 1024'h7ee98f67a5a16acd3be9a2a5e1181627fb1adf515e2c0b0b23eda769c159d8df602ae358586e7fddbba9e668be28e228641f96ce23b8d217df2170fb45de72383a6b4e0224e8a2a95527d0e76e8168f962086afe0ae7d2d37575dcf7011aefedce797f5852be829bf22a97e91feb9061dd673368f5169abdaa18011655af414d;
    5'b11010 : xpb = 1024'h67b87591458c003a6fbee7e643a434976de01af0a62f2502b51148c6ac717e2eb568af6745dd667ddcdf0e761206fcff625a1b92d7eb48879898a8cd497dfdb7af4434383341247c18253f3d12c9d2e70bb609e58e753a72d7fdafba0c52a2132120fc69aa6889066b69c0ba4b7785cfcf67308662af4a57208201ed8ae3f616;
    5'b11011 : xpb = 1024'h50875bbae57695a7a3942d26a6305306e0a5568fee323efa4634ea239789237e0aa67b76334c4d1dfe14368365e517d66094a0578c1dbef7520fe09f4d1d8937241d1a6e4199a64edb22ad92b7123cd4b563a8cd1202a2123a85827d178a543873c8797b02128f70e4a8e98b77037b3dc1672da3d047f9f096ec02c4c018aadf;
    5'b11100 : xpb = 1024'h395641e485612b14d769726708bc7176536a922f363558f1d7588b8082a0c8cd5fe4478520bb33be1f495e90b9c332ad5ecf251c405035670b87187150bd14b698f600a44ff228219e201be85b5aa6c25f1147b4959009b19d0d554022c2065dc66ff68c59bc95db5de8125ca28f70abb3672ac13de0a98a0d56039bf54d5fa8;
    5'b11101 : xpb = 1024'h2225280e254bc0820b3eb7a76b488fe5c62fcdce7e3872e9687c2cdd6db86e1cb52213940e2a1a5e407e869e0da14d845d09a9e0f482abd6c4fe5043545ca0360dcee6da5e4aa9f4611d8a3dffa310b008bee69c191d7150ff9528032df9b8831917739db1669c45d7273b2dce1b6619a56727deab79592383c004732a821471;
    5'b11110 : xpb = 1024'haf40e37c53655ef3f13fce7cdd4ae5538f5096dc63b8ce0f99fce3a58d0136c0a5fdfa2fb9900fe61b3aeab617f685b5b442ea5a8b522467e75881557fc2bb582a7cd106ca32bc7241af893a3eb7a9db26c85839caad8f0621cfac639316aa86bbef0af0910a2b0506663fef9a75b87976724fc191208bcfa2a054a5fb6c93a;
    5'b11111 : xpb = 1024'ha47039b7270f20253deeb9ff40bb14161d30483de3b6475008a028ecf6ea65c362e6292ab32e662d224715ff98bb93fcbd98db507f9a6901e88bff45966e2be66bcfe7f52a8caadef9b2698be10fa8bc501f1e03acbe6da07a315f83fe93bf5fed6dffea1183a1a8506573af1d03771ed84100fbd6f61586b70381261dcde46e;
    endcase
end

endmodule

module compressor_array_16_2_1033
(
    input  [15:0] col_in_0,
    input  [15:0] col_in_1,
    input  [15:0] col_in_2,
    input  [15:0] col_in_3,
    input  [15:0] col_in_4,
    input  [15:0] col_in_5,
    input  [15:0] col_in_6,
    input  [15:0] col_in_7,
    input  [15:0] col_in_8,
    input  [15:0] col_in_9,
    input  [15:0] col_in_10,
    input  [15:0] col_in_11,
    input  [15:0] col_in_12,
    input  [15:0] col_in_13,
    input  [15:0] col_in_14,
    input  [15:0] col_in_15,
    input  [15:0] col_in_16,
    input  [15:0] col_in_17,
    input  [15:0] col_in_18,
    input  [15:0] col_in_19,
    input  [15:0] col_in_20,
    input  [15:0] col_in_21,
    input  [15:0] col_in_22,
    input  [15:0] col_in_23,
    input  [15:0] col_in_24,
    input  [15:0] col_in_25,
    input  [15:0] col_in_26,
    input  [15:0] col_in_27,
    input  [15:0] col_in_28,
    input  [15:0] col_in_29,
    input  [15:0] col_in_30,
    input  [15:0] col_in_31,
    input  [15:0] col_in_32,
    input  [15:0] col_in_33,
    input  [15:0] col_in_34,
    input  [15:0] col_in_35,
    input  [15:0] col_in_36,
    input  [15:0] col_in_37,
    input  [15:0] col_in_38,
    input  [15:0] col_in_39,
    input  [15:0] col_in_40,
    input  [15:0] col_in_41,
    input  [15:0] col_in_42,
    input  [15:0] col_in_43,
    input  [15:0] col_in_44,
    input  [15:0] col_in_45,
    input  [15:0] col_in_46,
    input  [15:0] col_in_47,
    input  [15:0] col_in_48,
    input  [15:0] col_in_49,
    input  [15:0] col_in_50,
    input  [15:0] col_in_51,
    input  [15:0] col_in_52,
    input  [15:0] col_in_53,
    input  [15:0] col_in_54,
    input  [15:0] col_in_55,
    input  [15:0] col_in_56,
    input  [15:0] col_in_57,
    input  [15:0] col_in_58,
    input  [15:0] col_in_59,
    input  [15:0] col_in_60,
    input  [15:0] col_in_61,
    input  [15:0] col_in_62,
    input  [15:0] col_in_63,
    input  [15:0] col_in_64,
    input  [15:0] col_in_65,
    input  [15:0] col_in_66,
    input  [15:0] col_in_67,
    input  [15:0] col_in_68,
    input  [15:0] col_in_69,
    input  [15:0] col_in_70,
    input  [15:0] col_in_71,
    input  [15:0] col_in_72,
    input  [15:0] col_in_73,
    input  [15:0] col_in_74,
    input  [15:0] col_in_75,
    input  [15:0] col_in_76,
    input  [15:0] col_in_77,
    input  [15:0] col_in_78,
    input  [15:0] col_in_79,
    input  [15:0] col_in_80,
    input  [15:0] col_in_81,
    input  [15:0] col_in_82,
    input  [15:0] col_in_83,
    input  [15:0] col_in_84,
    input  [15:0] col_in_85,
    input  [15:0] col_in_86,
    input  [15:0] col_in_87,
    input  [15:0] col_in_88,
    input  [15:0] col_in_89,
    input  [15:0] col_in_90,
    input  [15:0] col_in_91,
    input  [15:0] col_in_92,
    input  [15:0] col_in_93,
    input  [15:0] col_in_94,
    input  [15:0] col_in_95,
    input  [15:0] col_in_96,
    input  [15:0] col_in_97,
    input  [15:0] col_in_98,
    input  [15:0] col_in_99,
    input  [15:0] col_in_100,
    input  [15:0] col_in_101,
    input  [15:0] col_in_102,
    input  [15:0] col_in_103,
    input  [15:0] col_in_104,
    input  [15:0] col_in_105,
    input  [15:0] col_in_106,
    input  [15:0] col_in_107,
    input  [15:0] col_in_108,
    input  [15:0] col_in_109,
    input  [15:0] col_in_110,
    input  [15:0] col_in_111,
    input  [15:0] col_in_112,
    input  [15:0] col_in_113,
    input  [15:0] col_in_114,
    input  [15:0] col_in_115,
    input  [15:0] col_in_116,
    input  [15:0] col_in_117,
    input  [15:0] col_in_118,
    input  [15:0] col_in_119,
    input  [15:0] col_in_120,
    input  [15:0] col_in_121,
    input  [15:0] col_in_122,
    input  [15:0] col_in_123,
    input  [15:0] col_in_124,
    input  [15:0] col_in_125,
    input  [15:0] col_in_126,
    input  [15:0] col_in_127,
    input  [15:0] col_in_128,
    input  [15:0] col_in_129,
    input  [15:0] col_in_130,
    input  [15:0] col_in_131,
    input  [15:0] col_in_132,
    input  [15:0] col_in_133,
    input  [15:0] col_in_134,
    input  [15:0] col_in_135,
    input  [15:0] col_in_136,
    input  [15:0] col_in_137,
    input  [15:0] col_in_138,
    input  [15:0] col_in_139,
    input  [15:0] col_in_140,
    input  [15:0] col_in_141,
    input  [15:0] col_in_142,
    input  [15:0] col_in_143,
    input  [15:0] col_in_144,
    input  [15:0] col_in_145,
    input  [15:0] col_in_146,
    input  [15:0] col_in_147,
    input  [15:0] col_in_148,
    input  [15:0] col_in_149,
    input  [15:0] col_in_150,
    input  [15:0] col_in_151,
    input  [15:0] col_in_152,
    input  [15:0] col_in_153,
    input  [15:0] col_in_154,
    input  [15:0] col_in_155,
    input  [15:0] col_in_156,
    input  [15:0] col_in_157,
    input  [15:0] col_in_158,
    input  [15:0] col_in_159,
    input  [15:0] col_in_160,
    input  [15:0] col_in_161,
    input  [15:0] col_in_162,
    input  [15:0] col_in_163,
    input  [15:0] col_in_164,
    input  [15:0] col_in_165,
    input  [15:0] col_in_166,
    input  [15:0] col_in_167,
    input  [15:0] col_in_168,
    input  [15:0] col_in_169,
    input  [15:0] col_in_170,
    input  [15:0] col_in_171,
    input  [15:0] col_in_172,
    input  [15:0] col_in_173,
    input  [15:0] col_in_174,
    input  [15:0] col_in_175,
    input  [15:0] col_in_176,
    input  [15:0] col_in_177,
    input  [15:0] col_in_178,
    input  [15:0] col_in_179,
    input  [15:0] col_in_180,
    input  [15:0] col_in_181,
    input  [15:0] col_in_182,
    input  [15:0] col_in_183,
    input  [15:0] col_in_184,
    input  [15:0] col_in_185,
    input  [15:0] col_in_186,
    input  [15:0] col_in_187,
    input  [15:0] col_in_188,
    input  [15:0] col_in_189,
    input  [15:0] col_in_190,
    input  [15:0] col_in_191,
    input  [15:0] col_in_192,
    input  [15:0] col_in_193,
    input  [15:0] col_in_194,
    input  [15:0] col_in_195,
    input  [15:0] col_in_196,
    input  [15:0] col_in_197,
    input  [15:0] col_in_198,
    input  [15:0] col_in_199,
    input  [15:0] col_in_200,
    input  [15:0] col_in_201,
    input  [15:0] col_in_202,
    input  [15:0] col_in_203,
    input  [15:0] col_in_204,
    input  [15:0] col_in_205,
    input  [15:0] col_in_206,
    input  [15:0] col_in_207,
    input  [15:0] col_in_208,
    input  [15:0] col_in_209,
    input  [15:0] col_in_210,
    input  [15:0] col_in_211,
    input  [15:0] col_in_212,
    input  [15:0] col_in_213,
    input  [15:0] col_in_214,
    input  [15:0] col_in_215,
    input  [15:0] col_in_216,
    input  [15:0] col_in_217,
    input  [15:0] col_in_218,
    input  [15:0] col_in_219,
    input  [15:0] col_in_220,
    input  [15:0] col_in_221,
    input  [15:0] col_in_222,
    input  [15:0] col_in_223,
    input  [15:0] col_in_224,
    input  [15:0] col_in_225,
    input  [15:0] col_in_226,
    input  [15:0] col_in_227,
    input  [15:0] col_in_228,
    input  [15:0] col_in_229,
    input  [15:0] col_in_230,
    input  [15:0] col_in_231,
    input  [15:0] col_in_232,
    input  [15:0] col_in_233,
    input  [15:0] col_in_234,
    input  [15:0] col_in_235,
    input  [15:0] col_in_236,
    input  [15:0] col_in_237,
    input  [15:0] col_in_238,
    input  [15:0] col_in_239,
    input  [15:0] col_in_240,
    input  [15:0] col_in_241,
    input  [15:0] col_in_242,
    input  [15:0] col_in_243,
    input  [15:0] col_in_244,
    input  [15:0] col_in_245,
    input  [15:0] col_in_246,
    input  [15:0] col_in_247,
    input  [15:0] col_in_248,
    input  [15:0] col_in_249,
    input  [15:0] col_in_250,
    input  [15:0] col_in_251,
    input  [15:0] col_in_252,
    input  [15:0] col_in_253,
    input  [15:0] col_in_254,
    input  [15:0] col_in_255,
    input  [15:0] col_in_256,
    input  [15:0] col_in_257,
    input  [15:0] col_in_258,
    input  [15:0] col_in_259,
    input  [15:0] col_in_260,
    input  [15:0] col_in_261,
    input  [15:0] col_in_262,
    input  [15:0] col_in_263,
    input  [15:0] col_in_264,
    input  [15:0] col_in_265,
    input  [15:0] col_in_266,
    input  [15:0] col_in_267,
    input  [15:0] col_in_268,
    input  [15:0] col_in_269,
    input  [15:0] col_in_270,
    input  [15:0] col_in_271,
    input  [15:0] col_in_272,
    input  [15:0] col_in_273,
    input  [15:0] col_in_274,
    input  [15:0] col_in_275,
    input  [15:0] col_in_276,
    input  [15:0] col_in_277,
    input  [15:0] col_in_278,
    input  [15:0] col_in_279,
    input  [15:0] col_in_280,
    input  [15:0] col_in_281,
    input  [15:0] col_in_282,
    input  [15:0] col_in_283,
    input  [15:0] col_in_284,
    input  [15:0] col_in_285,
    input  [15:0] col_in_286,
    input  [15:0] col_in_287,
    input  [15:0] col_in_288,
    input  [15:0] col_in_289,
    input  [15:0] col_in_290,
    input  [15:0] col_in_291,
    input  [15:0] col_in_292,
    input  [15:0] col_in_293,
    input  [15:0] col_in_294,
    input  [15:0] col_in_295,
    input  [15:0] col_in_296,
    input  [15:0] col_in_297,
    input  [15:0] col_in_298,
    input  [15:0] col_in_299,
    input  [15:0] col_in_300,
    input  [15:0] col_in_301,
    input  [15:0] col_in_302,
    input  [15:0] col_in_303,
    input  [15:0] col_in_304,
    input  [15:0] col_in_305,
    input  [15:0] col_in_306,
    input  [15:0] col_in_307,
    input  [15:0] col_in_308,
    input  [15:0] col_in_309,
    input  [15:0] col_in_310,
    input  [15:0] col_in_311,
    input  [15:0] col_in_312,
    input  [15:0] col_in_313,
    input  [15:0] col_in_314,
    input  [15:0] col_in_315,
    input  [15:0] col_in_316,
    input  [15:0] col_in_317,
    input  [15:0] col_in_318,
    input  [15:0] col_in_319,
    input  [15:0] col_in_320,
    input  [15:0] col_in_321,
    input  [15:0] col_in_322,
    input  [15:0] col_in_323,
    input  [15:0] col_in_324,
    input  [15:0] col_in_325,
    input  [15:0] col_in_326,
    input  [15:0] col_in_327,
    input  [15:0] col_in_328,
    input  [15:0] col_in_329,
    input  [15:0] col_in_330,
    input  [15:0] col_in_331,
    input  [15:0] col_in_332,
    input  [15:0] col_in_333,
    input  [15:0] col_in_334,
    input  [15:0] col_in_335,
    input  [15:0] col_in_336,
    input  [15:0] col_in_337,
    input  [15:0] col_in_338,
    input  [15:0] col_in_339,
    input  [15:0] col_in_340,
    input  [15:0] col_in_341,
    input  [15:0] col_in_342,
    input  [15:0] col_in_343,
    input  [15:0] col_in_344,
    input  [15:0] col_in_345,
    input  [15:0] col_in_346,
    input  [15:0] col_in_347,
    input  [15:0] col_in_348,
    input  [15:0] col_in_349,
    input  [15:0] col_in_350,
    input  [15:0] col_in_351,
    input  [15:0] col_in_352,
    input  [15:0] col_in_353,
    input  [15:0] col_in_354,
    input  [15:0] col_in_355,
    input  [15:0] col_in_356,
    input  [15:0] col_in_357,
    input  [15:0] col_in_358,
    input  [15:0] col_in_359,
    input  [15:0] col_in_360,
    input  [15:0] col_in_361,
    input  [15:0] col_in_362,
    input  [15:0] col_in_363,
    input  [15:0] col_in_364,
    input  [15:0] col_in_365,
    input  [15:0] col_in_366,
    input  [15:0] col_in_367,
    input  [15:0] col_in_368,
    input  [15:0] col_in_369,
    input  [15:0] col_in_370,
    input  [15:0] col_in_371,
    input  [15:0] col_in_372,
    input  [15:0] col_in_373,
    input  [15:0] col_in_374,
    input  [15:0] col_in_375,
    input  [15:0] col_in_376,
    input  [15:0] col_in_377,
    input  [15:0] col_in_378,
    input  [15:0] col_in_379,
    input  [15:0] col_in_380,
    input  [15:0] col_in_381,
    input  [15:0] col_in_382,
    input  [15:0] col_in_383,
    input  [15:0] col_in_384,
    input  [15:0] col_in_385,
    input  [15:0] col_in_386,
    input  [15:0] col_in_387,
    input  [15:0] col_in_388,
    input  [15:0] col_in_389,
    input  [15:0] col_in_390,
    input  [15:0] col_in_391,
    input  [15:0] col_in_392,
    input  [15:0] col_in_393,
    input  [15:0] col_in_394,
    input  [15:0] col_in_395,
    input  [15:0] col_in_396,
    input  [15:0] col_in_397,
    input  [15:0] col_in_398,
    input  [15:0] col_in_399,
    input  [15:0] col_in_400,
    input  [15:0] col_in_401,
    input  [15:0] col_in_402,
    input  [15:0] col_in_403,
    input  [15:0] col_in_404,
    input  [15:0] col_in_405,
    input  [15:0] col_in_406,
    input  [15:0] col_in_407,
    input  [15:0] col_in_408,
    input  [15:0] col_in_409,
    input  [15:0] col_in_410,
    input  [15:0] col_in_411,
    input  [15:0] col_in_412,
    input  [15:0] col_in_413,
    input  [15:0] col_in_414,
    input  [15:0] col_in_415,
    input  [15:0] col_in_416,
    input  [15:0] col_in_417,
    input  [15:0] col_in_418,
    input  [15:0] col_in_419,
    input  [15:0] col_in_420,
    input  [15:0] col_in_421,
    input  [15:0] col_in_422,
    input  [15:0] col_in_423,
    input  [15:0] col_in_424,
    input  [15:0] col_in_425,
    input  [15:0] col_in_426,
    input  [15:0] col_in_427,
    input  [15:0] col_in_428,
    input  [15:0] col_in_429,
    input  [15:0] col_in_430,
    input  [15:0] col_in_431,
    input  [15:0] col_in_432,
    input  [15:0] col_in_433,
    input  [15:0] col_in_434,
    input  [15:0] col_in_435,
    input  [15:0] col_in_436,
    input  [15:0] col_in_437,
    input  [15:0] col_in_438,
    input  [15:0] col_in_439,
    input  [15:0] col_in_440,
    input  [15:0] col_in_441,
    input  [15:0] col_in_442,
    input  [15:0] col_in_443,
    input  [15:0] col_in_444,
    input  [15:0] col_in_445,
    input  [15:0] col_in_446,
    input  [15:0] col_in_447,
    input  [15:0] col_in_448,
    input  [15:0] col_in_449,
    input  [15:0] col_in_450,
    input  [15:0] col_in_451,
    input  [15:0] col_in_452,
    input  [15:0] col_in_453,
    input  [15:0] col_in_454,
    input  [15:0] col_in_455,
    input  [15:0] col_in_456,
    input  [15:0] col_in_457,
    input  [15:0] col_in_458,
    input  [15:0] col_in_459,
    input  [15:0] col_in_460,
    input  [15:0] col_in_461,
    input  [15:0] col_in_462,
    input  [15:0] col_in_463,
    input  [15:0] col_in_464,
    input  [15:0] col_in_465,
    input  [15:0] col_in_466,
    input  [15:0] col_in_467,
    input  [15:0] col_in_468,
    input  [15:0] col_in_469,
    input  [15:0] col_in_470,
    input  [15:0] col_in_471,
    input  [15:0] col_in_472,
    input  [15:0] col_in_473,
    input  [15:0] col_in_474,
    input  [15:0] col_in_475,
    input  [15:0] col_in_476,
    input  [15:0] col_in_477,
    input  [15:0] col_in_478,
    input  [15:0] col_in_479,
    input  [15:0] col_in_480,
    input  [15:0] col_in_481,
    input  [15:0] col_in_482,
    input  [15:0] col_in_483,
    input  [15:0] col_in_484,
    input  [15:0] col_in_485,
    input  [15:0] col_in_486,
    input  [15:0] col_in_487,
    input  [15:0] col_in_488,
    input  [15:0] col_in_489,
    input  [15:0] col_in_490,
    input  [15:0] col_in_491,
    input  [15:0] col_in_492,
    input  [15:0] col_in_493,
    input  [15:0] col_in_494,
    input  [15:0] col_in_495,
    input  [15:0] col_in_496,
    input  [15:0] col_in_497,
    input  [15:0] col_in_498,
    input  [15:0] col_in_499,
    input  [15:0] col_in_500,
    input  [15:0] col_in_501,
    input  [15:0] col_in_502,
    input  [15:0] col_in_503,
    input  [15:0] col_in_504,
    input  [15:0] col_in_505,
    input  [15:0] col_in_506,
    input  [15:0] col_in_507,
    input  [15:0] col_in_508,
    input  [15:0] col_in_509,
    input  [15:0] col_in_510,
    input  [15:0] col_in_511,
    input  [15:0] col_in_512,
    input  [15:0] col_in_513,
    input  [15:0] col_in_514,
    input  [15:0] col_in_515,
    input  [15:0] col_in_516,
    input  [15:0] col_in_517,
    input  [15:0] col_in_518,
    input  [15:0] col_in_519,
    input  [15:0] col_in_520,
    input  [15:0] col_in_521,
    input  [15:0] col_in_522,
    input  [15:0] col_in_523,
    input  [15:0] col_in_524,
    input  [15:0] col_in_525,
    input  [15:0] col_in_526,
    input  [15:0] col_in_527,
    input  [15:0] col_in_528,
    input  [15:0] col_in_529,
    input  [15:0] col_in_530,
    input  [15:0] col_in_531,
    input  [15:0] col_in_532,
    input  [15:0] col_in_533,
    input  [15:0] col_in_534,
    input  [15:0] col_in_535,
    input  [15:0] col_in_536,
    input  [15:0] col_in_537,
    input  [15:0] col_in_538,
    input  [15:0] col_in_539,
    input  [15:0] col_in_540,
    input  [15:0] col_in_541,
    input  [15:0] col_in_542,
    input  [15:0] col_in_543,
    input  [15:0] col_in_544,
    input  [15:0] col_in_545,
    input  [15:0] col_in_546,
    input  [15:0] col_in_547,
    input  [15:0] col_in_548,
    input  [15:0] col_in_549,
    input  [15:0] col_in_550,
    input  [15:0] col_in_551,
    input  [15:0] col_in_552,
    input  [15:0] col_in_553,
    input  [15:0] col_in_554,
    input  [15:0] col_in_555,
    input  [15:0] col_in_556,
    input  [15:0] col_in_557,
    input  [15:0] col_in_558,
    input  [15:0] col_in_559,
    input  [15:0] col_in_560,
    input  [15:0] col_in_561,
    input  [15:0] col_in_562,
    input  [15:0] col_in_563,
    input  [15:0] col_in_564,
    input  [15:0] col_in_565,
    input  [15:0] col_in_566,
    input  [15:0] col_in_567,
    input  [15:0] col_in_568,
    input  [15:0] col_in_569,
    input  [15:0] col_in_570,
    input  [15:0] col_in_571,
    input  [15:0] col_in_572,
    input  [15:0] col_in_573,
    input  [15:0] col_in_574,
    input  [15:0] col_in_575,
    input  [15:0] col_in_576,
    input  [15:0] col_in_577,
    input  [15:0] col_in_578,
    input  [15:0] col_in_579,
    input  [15:0] col_in_580,
    input  [15:0] col_in_581,
    input  [15:0] col_in_582,
    input  [15:0] col_in_583,
    input  [15:0] col_in_584,
    input  [15:0] col_in_585,
    input  [15:0] col_in_586,
    input  [15:0] col_in_587,
    input  [15:0] col_in_588,
    input  [15:0] col_in_589,
    input  [15:0] col_in_590,
    input  [15:0] col_in_591,
    input  [15:0] col_in_592,
    input  [15:0] col_in_593,
    input  [15:0] col_in_594,
    input  [15:0] col_in_595,
    input  [15:0] col_in_596,
    input  [15:0] col_in_597,
    input  [15:0] col_in_598,
    input  [15:0] col_in_599,
    input  [15:0] col_in_600,
    input  [15:0] col_in_601,
    input  [15:0] col_in_602,
    input  [15:0] col_in_603,
    input  [15:0] col_in_604,
    input  [15:0] col_in_605,
    input  [15:0] col_in_606,
    input  [15:0] col_in_607,
    input  [15:0] col_in_608,
    input  [15:0] col_in_609,
    input  [15:0] col_in_610,
    input  [15:0] col_in_611,
    input  [15:0] col_in_612,
    input  [15:0] col_in_613,
    input  [15:0] col_in_614,
    input  [15:0] col_in_615,
    input  [15:0] col_in_616,
    input  [15:0] col_in_617,
    input  [15:0] col_in_618,
    input  [15:0] col_in_619,
    input  [15:0] col_in_620,
    input  [15:0] col_in_621,
    input  [15:0] col_in_622,
    input  [15:0] col_in_623,
    input  [15:0] col_in_624,
    input  [15:0] col_in_625,
    input  [15:0] col_in_626,
    input  [15:0] col_in_627,
    input  [15:0] col_in_628,
    input  [15:0] col_in_629,
    input  [15:0] col_in_630,
    input  [15:0] col_in_631,
    input  [15:0] col_in_632,
    input  [15:0] col_in_633,
    input  [15:0] col_in_634,
    input  [15:0] col_in_635,
    input  [15:0] col_in_636,
    input  [15:0] col_in_637,
    input  [15:0] col_in_638,
    input  [15:0] col_in_639,
    input  [15:0] col_in_640,
    input  [15:0] col_in_641,
    input  [15:0] col_in_642,
    input  [15:0] col_in_643,
    input  [15:0] col_in_644,
    input  [15:0] col_in_645,
    input  [15:0] col_in_646,
    input  [15:0] col_in_647,
    input  [15:0] col_in_648,
    input  [15:0] col_in_649,
    input  [15:0] col_in_650,
    input  [15:0] col_in_651,
    input  [15:0] col_in_652,
    input  [15:0] col_in_653,
    input  [15:0] col_in_654,
    input  [15:0] col_in_655,
    input  [15:0] col_in_656,
    input  [15:0] col_in_657,
    input  [15:0] col_in_658,
    input  [15:0] col_in_659,
    input  [15:0] col_in_660,
    input  [15:0] col_in_661,
    input  [15:0] col_in_662,
    input  [15:0] col_in_663,
    input  [15:0] col_in_664,
    input  [15:0] col_in_665,
    input  [15:0] col_in_666,
    input  [15:0] col_in_667,
    input  [15:0] col_in_668,
    input  [15:0] col_in_669,
    input  [15:0] col_in_670,
    input  [15:0] col_in_671,
    input  [15:0] col_in_672,
    input  [15:0] col_in_673,
    input  [15:0] col_in_674,
    input  [15:0] col_in_675,
    input  [15:0] col_in_676,
    input  [15:0] col_in_677,
    input  [15:0] col_in_678,
    input  [15:0] col_in_679,
    input  [15:0] col_in_680,
    input  [15:0] col_in_681,
    input  [15:0] col_in_682,
    input  [15:0] col_in_683,
    input  [15:0] col_in_684,
    input  [15:0] col_in_685,
    input  [15:0] col_in_686,
    input  [15:0] col_in_687,
    input  [15:0] col_in_688,
    input  [15:0] col_in_689,
    input  [15:0] col_in_690,
    input  [15:0] col_in_691,
    input  [15:0] col_in_692,
    input  [15:0] col_in_693,
    input  [15:0] col_in_694,
    input  [15:0] col_in_695,
    input  [15:0] col_in_696,
    input  [15:0] col_in_697,
    input  [15:0] col_in_698,
    input  [15:0] col_in_699,
    input  [15:0] col_in_700,
    input  [15:0] col_in_701,
    input  [15:0] col_in_702,
    input  [15:0] col_in_703,
    input  [15:0] col_in_704,
    input  [15:0] col_in_705,
    input  [15:0] col_in_706,
    input  [15:0] col_in_707,
    input  [15:0] col_in_708,
    input  [15:0] col_in_709,
    input  [15:0] col_in_710,
    input  [15:0] col_in_711,
    input  [15:0] col_in_712,
    input  [15:0] col_in_713,
    input  [15:0] col_in_714,
    input  [15:0] col_in_715,
    input  [15:0] col_in_716,
    input  [15:0] col_in_717,
    input  [15:0] col_in_718,
    input  [15:0] col_in_719,
    input  [15:0] col_in_720,
    input  [15:0] col_in_721,
    input  [15:0] col_in_722,
    input  [15:0] col_in_723,
    input  [15:0] col_in_724,
    input  [15:0] col_in_725,
    input  [15:0] col_in_726,
    input  [15:0] col_in_727,
    input  [15:0] col_in_728,
    input  [15:0] col_in_729,
    input  [15:0] col_in_730,
    input  [15:0] col_in_731,
    input  [15:0] col_in_732,
    input  [15:0] col_in_733,
    input  [15:0] col_in_734,
    input  [15:0] col_in_735,
    input  [15:0] col_in_736,
    input  [15:0] col_in_737,
    input  [15:0] col_in_738,
    input  [15:0] col_in_739,
    input  [15:0] col_in_740,
    input  [15:0] col_in_741,
    input  [15:0] col_in_742,
    input  [15:0] col_in_743,
    input  [15:0] col_in_744,
    input  [15:0] col_in_745,
    input  [15:0] col_in_746,
    input  [15:0] col_in_747,
    input  [15:0] col_in_748,
    input  [15:0] col_in_749,
    input  [15:0] col_in_750,
    input  [15:0] col_in_751,
    input  [15:0] col_in_752,
    input  [15:0] col_in_753,
    input  [15:0] col_in_754,
    input  [15:0] col_in_755,
    input  [15:0] col_in_756,
    input  [15:0] col_in_757,
    input  [15:0] col_in_758,
    input  [15:0] col_in_759,
    input  [15:0] col_in_760,
    input  [15:0] col_in_761,
    input  [15:0] col_in_762,
    input  [15:0] col_in_763,
    input  [15:0] col_in_764,
    input  [15:0] col_in_765,
    input  [15:0] col_in_766,
    input  [15:0] col_in_767,
    input  [15:0] col_in_768,
    input  [15:0] col_in_769,
    input  [15:0] col_in_770,
    input  [15:0] col_in_771,
    input  [15:0] col_in_772,
    input  [15:0] col_in_773,
    input  [15:0] col_in_774,
    input  [15:0] col_in_775,
    input  [15:0] col_in_776,
    input  [15:0] col_in_777,
    input  [15:0] col_in_778,
    input  [15:0] col_in_779,
    input  [15:0] col_in_780,
    input  [15:0] col_in_781,
    input  [15:0] col_in_782,
    input  [15:0] col_in_783,
    input  [15:0] col_in_784,
    input  [15:0] col_in_785,
    input  [15:0] col_in_786,
    input  [15:0] col_in_787,
    input  [15:0] col_in_788,
    input  [15:0] col_in_789,
    input  [15:0] col_in_790,
    input  [15:0] col_in_791,
    input  [15:0] col_in_792,
    input  [15:0] col_in_793,
    input  [15:0] col_in_794,
    input  [15:0] col_in_795,
    input  [15:0] col_in_796,
    input  [15:0] col_in_797,
    input  [15:0] col_in_798,
    input  [15:0] col_in_799,
    input  [15:0] col_in_800,
    input  [15:0] col_in_801,
    input  [15:0] col_in_802,
    input  [15:0] col_in_803,
    input  [15:0] col_in_804,
    input  [15:0] col_in_805,
    input  [15:0] col_in_806,
    input  [15:0] col_in_807,
    input  [15:0] col_in_808,
    input  [15:0] col_in_809,
    input  [15:0] col_in_810,
    input  [15:0] col_in_811,
    input  [15:0] col_in_812,
    input  [15:0] col_in_813,
    input  [15:0] col_in_814,
    input  [15:0] col_in_815,
    input  [15:0] col_in_816,
    input  [15:0] col_in_817,
    input  [15:0] col_in_818,
    input  [15:0] col_in_819,
    input  [15:0] col_in_820,
    input  [15:0] col_in_821,
    input  [15:0] col_in_822,
    input  [15:0] col_in_823,
    input  [15:0] col_in_824,
    input  [15:0] col_in_825,
    input  [15:0] col_in_826,
    input  [15:0] col_in_827,
    input  [15:0] col_in_828,
    input  [15:0] col_in_829,
    input  [15:0] col_in_830,
    input  [15:0] col_in_831,
    input  [15:0] col_in_832,
    input  [15:0] col_in_833,
    input  [15:0] col_in_834,
    input  [15:0] col_in_835,
    input  [15:0] col_in_836,
    input  [15:0] col_in_837,
    input  [15:0] col_in_838,
    input  [15:0] col_in_839,
    input  [15:0] col_in_840,
    input  [15:0] col_in_841,
    input  [15:0] col_in_842,
    input  [15:0] col_in_843,
    input  [15:0] col_in_844,
    input  [15:0] col_in_845,
    input  [15:0] col_in_846,
    input  [15:0] col_in_847,
    input  [15:0] col_in_848,
    input  [15:0] col_in_849,
    input  [15:0] col_in_850,
    input  [15:0] col_in_851,
    input  [15:0] col_in_852,
    input  [15:0] col_in_853,
    input  [15:0] col_in_854,
    input  [15:0] col_in_855,
    input  [15:0] col_in_856,
    input  [15:0] col_in_857,
    input  [15:0] col_in_858,
    input  [15:0] col_in_859,
    input  [15:0] col_in_860,
    input  [15:0] col_in_861,
    input  [15:0] col_in_862,
    input  [15:0] col_in_863,
    input  [15:0] col_in_864,
    input  [15:0] col_in_865,
    input  [15:0] col_in_866,
    input  [15:0] col_in_867,
    input  [15:0] col_in_868,
    input  [15:0] col_in_869,
    input  [15:0] col_in_870,
    input  [15:0] col_in_871,
    input  [15:0] col_in_872,
    input  [15:0] col_in_873,
    input  [15:0] col_in_874,
    input  [15:0] col_in_875,
    input  [15:0] col_in_876,
    input  [15:0] col_in_877,
    input  [15:0] col_in_878,
    input  [15:0] col_in_879,
    input  [15:0] col_in_880,
    input  [15:0] col_in_881,
    input  [15:0] col_in_882,
    input  [15:0] col_in_883,
    input  [15:0] col_in_884,
    input  [15:0] col_in_885,
    input  [15:0] col_in_886,
    input  [15:0] col_in_887,
    input  [15:0] col_in_888,
    input  [15:0] col_in_889,
    input  [15:0] col_in_890,
    input  [15:0] col_in_891,
    input  [15:0] col_in_892,
    input  [15:0] col_in_893,
    input  [15:0] col_in_894,
    input  [15:0] col_in_895,
    input  [15:0] col_in_896,
    input  [15:0] col_in_897,
    input  [15:0] col_in_898,
    input  [15:0] col_in_899,
    input  [15:0] col_in_900,
    input  [15:0] col_in_901,
    input  [15:0] col_in_902,
    input  [15:0] col_in_903,
    input  [15:0] col_in_904,
    input  [15:0] col_in_905,
    input  [15:0] col_in_906,
    input  [15:0] col_in_907,
    input  [15:0] col_in_908,
    input  [15:0] col_in_909,
    input  [15:0] col_in_910,
    input  [15:0] col_in_911,
    input  [15:0] col_in_912,
    input  [15:0] col_in_913,
    input  [15:0] col_in_914,
    input  [15:0] col_in_915,
    input  [15:0] col_in_916,
    input  [15:0] col_in_917,
    input  [15:0] col_in_918,
    input  [15:0] col_in_919,
    input  [15:0] col_in_920,
    input  [15:0] col_in_921,
    input  [15:0] col_in_922,
    input  [15:0] col_in_923,
    input  [15:0] col_in_924,
    input  [15:0] col_in_925,
    input  [15:0] col_in_926,
    input  [15:0] col_in_927,
    input  [15:0] col_in_928,
    input  [15:0] col_in_929,
    input  [15:0] col_in_930,
    input  [15:0] col_in_931,
    input  [15:0] col_in_932,
    input  [15:0] col_in_933,
    input  [15:0] col_in_934,
    input  [15:0] col_in_935,
    input  [15:0] col_in_936,
    input  [15:0] col_in_937,
    input  [15:0] col_in_938,
    input  [15:0] col_in_939,
    input  [15:0] col_in_940,
    input  [15:0] col_in_941,
    input  [15:0] col_in_942,
    input  [15:0] col_in_943,
    input  [15:0] col_in_944,
    input  [15:0] col_in_945,
    input  [15:0] col_in_946,
    input  [15:0] col_in_947,
    input  [15:0] col_in_948,
    input  [15:0] col_in_949,
    input  [15:0] col_in_950,
    input  [15:0] col_in_951,
    input  [15:0] col_in_952,
    input  [15:0] col_in_953,
    input  [15:0] col_in_954,
    input  [15:0] col_in_955,
    input  [15:0] col_in_956,
    input  [15:0] col_in_957,
    input  [15:0] col_in_958,
    input  [15:0] col_in_959,
    input  [15:0] col_in_960,
    input  [15:0] col_in_961,
    input  [15:0] col_in_962,
    input  [15:0] col_in_963,
    input  [15:0] col_in_964,
    input  [15:0] col_in_965,
    input  [15:0] col_in_966,
    input  [15:0] col_in_967,
    input  [15:0] col_in_968,
    input  [15:0] col_in_969,
    input  [15:0] col_in_970,
    input  [15:0] col_in_971,
    input  [15:0] col_in_972,
    input  [15:0] col_in_973,
    input  [15:0] col_in_974,
    input  [15:0] col_in_975,
    input  [15:0] col_in_976,
    input  [15:0] col_in_977,
    input  [15:0] col_in_978,
    input  [15:0] col_in_979,
    input  [15:0] col_in_980,
    input  [15:0] col_in_981,
    input  [15:0] col_in_982,
    input  [15:0] col_in_983,
    input  [15:0] col_in_984,
    input  [15:0] col_in_985,
    input  [15:0] col_in_986,
    input  [15:0] col_in_987,
    input  [15:0] col_in_988,
    input  [15:0] col_in_989,
    input  [15:0] col_in_990,
    input  [15:0] col_in_991,
    input  [15:0] col_in_992,
    input  [15:0] col_in_993,
    input  [15:0] col_in_994,
    input  [15:0] col_in_995,
    input  [15:0] col_in_996,
    input  [15:0] col_in_997,
    input  [15:0] col_in_998,
    input  [15:0] col_in_999,
    input  [15:0] col_in_1000,
    input  [15:0] col_in_1001,
    input  [15:0] col_in_1002,
    input  [15:0] col_in_1003,
    input  [15:0] col_in_1004,
    input  [15:0] col_in_1005,
    input  [15:0] col_in_1006,
    input  [15:0] col_in_1007,
    input  [15:0] col_in_1008,
    input  [15:0] col_in_1009,
    input  [15:0] col_in_1010,
    input  [15:0] col_in_1011,
    input  [15:0] col_in_1012,
    input  [15:0] col_in_1013,
    input  [15:0] col_in_1014,
    input  [15:0] col_in_1015,
    input  [15:0] col_in_1016,
    input  [15:0] col_in_1017,
    input  [15:0] col_in_1018,
    input  [15:0] col_in_1019,
    input  [15:0] col_in_1020,
    input  [15:0] col_in_1021,
    input  [15:0] col_in_1022,
    input  [15:0] col_in_1023,
    input  [15:0] col_in_1024,
    input  [15:0] col_in_1025,
    input  [15:0] col_in_1026,
    input  [15:0] col_in_1027,
    input  [15:0] col_in_1028,
    input  [15:0] col_in_1029,
    input  [15:0] col_in_1030,
    input  [15:0] col_in_1031,
    input  [15:0] col_in_1032,

    output [1:0] col_out_0,
    output [1:0] col_out_1,
    output [1:0] col_out_2,
    output [1:0] col_out_3,
    output [1:0] col_out_4,
    output [1:0] col_out_5,
    output [1:0] col_out_6,
    output [1:0] col_out_7,
    output [1:0] col_out_8,
    output [1:0] col_out_9,
    output [1:0] col_out_10,
    output [1:0] col_out_11,
    output [1:0] col_out_12,
    output [1:0] col_out_13,
    output [1:0] col_out_14,
    output [1:0] col_out_15,
    output [1:0] col_out_16,
    output [1:0] col_out_17,
    output [1:0] col_out_18,
    output [1:0] col_out_19,
    output [1:0] col_out_20,
    output [1:0] col_out_21,
    output [1:0] col_out_22,
    output [1:0] col_out_23,
    output [1:0] col_out_24,
    output [1:0] col_out_25,
    output [1:0] col_out_26,
    output [1:0] col_out_27,
    output [1:0] col_out_28,
    output [1:0] col_out_29,
    output [1:0] col_out_30,
    output [1:0] col_out_31,
    output [1:0] col_out_32,
    output [1:0] col_out_33,
    output [1:0] col_out_34,
    output [1:0] col_out_35,
    output [1:0] col_out_36,
    output [1:0] col_out_37,
    output [1:0] col_out_38,
    output [1:0] col_out_39,
    output [1:0] col_out_40,
    output [1:0] col_out_41,
    output [1:0] col_out_42,
    output [1:0] col_out_43,
    output [1:0] col_out_44,
    output [1:0] col_out_45,
    output [1:0] col_out_46,
    output [1:0] col_out_47,
    output [1:0] col_out_48,
    output [1:0] col_out_49,
    output [1:0] col_out_50,
    output [1:0] col_out_51,
    output [1:0] col_out_52,
    output [1:0] col_out_53,
    output [1:0] col_out_54,
    output [1:0] col_out_55,
    output [1:0] col_out_56,
    output [1:0] col_out_57,
    output [1:0] col_out_58,
    output [1:0] col_out_59,
    output [1:0] col_out_60,
    output [1:0] col_out_61,
    output [1:0] col_out_62,
    output [1:0] col_out_63,
    output [1:0] col_out_64,
    output [1:0] col_out_65,
    output [1:0] col_out_66,
    output [1:0] col_out_67,
    output [1:0] col_out_68,
    output [1:0] col_out_69,
    output [1:0] col_out_70,
    output [1:0] col_out_71,
    output [1:0] col_out_72,
    output [1:0] col_out_73,
    output [1:0] col_out_74,
    output [1:0] col_out_75,
    output [1:0] col_out_76,
    output [1:0] col_out_77,
    output [1:0] col_out_78,
    output [1:0] col_out_79,
    output [1:0] col_out_80,
    output [1:0] col_out_81,
    output [1:0] col_out_82,
    output [1:0] col_out_83,
    output [1:0] col_out_84,
    output [1:0] col_out_85,
    output [1:0] col_out_86,
    output [1:0] col_out_87,
    output [1:0] col_out_88,
    output [1:0] col_out_89,
    output [1:0] col_out_90,
    output [1:0] col_out_91,
    output [1:0] col_out_92,
    output [1:0] col_out_93,
    output [1:0] col_out_94,
    output [1:0] col_out_95,
    output [1:0] col_out_96,
    output [1:0] col_out_97,
    output [1:0] col_out_98,
    output [1:0] col_out_99,
    output [1:0] col_out_100,
    output [1:0] col_out_101,
    output [1:0] col_out_102,
    output [1:0] col_out_103,
    output [1:0] col_out_104,
    output [1:0] col_out_105,
    output [1:0] col_out_106,
    output [1:0] col_out_107,
    output [1:0] col_out_108,
    output [1:0] col_out_109,
    output [1:0] col_out_110,
    output [1:0] col_out_111,
    output [1:0] col_out_112,
    output [1:0] col_out_113,
    output [1:0] col_out_114,
    output [1:0] col_out_115,
    output [1:0] col_out_116,
    output [1:0] col_out_117,
    output [1:0] col_out_118,
    output [1:0] col_out_119,
    output [1:0] col_out_120,
    output [1:0] col_out_121,
    output [1:0] col_out_122,
    output [1:0] col_out_123,
    output [1:0] col_out_124,
    output [1:0] col_out_125,
    output [1:0] col_out_126,
    output [1:0] col_out_127,
    output [1:0] col_out_128,
    output [1:0] col_out_129,
    output [1:0] col_out_130,
    output [1:0] col_out_131,
    output [1:0] col_out_132,
    output [1:0] col_out_133,
    output [1:0] col_out_134,
    output [1:0] col_out_135,
    output [1:0] col_out_136,
    output [1:0] col_out_137,
    output [1:0] col_out_138,
    output [1:0] col_out_139,
    output [1:0] col_out_140,
    output [1:0] col_out_141,
    output [1:0] col_out_142,
    output [1:0] col_out_143,
    output [1:0] col_out_144,
    output [1:0] col_out_145,
    output [1:0] col_out_146,
    output [1:0] col_out_147,
    output [1:0] col_out_148,
    output [1:0] col_out_149,
    output [1:0] col_out_150,
    output [1:0] col_out_151,
    output [1:0] col_out_152,
    output [1:0] col_out_153,
    output [1:0] col_out_154,
    output [1:0] col_out_155,
    output [1:0] col_out_156,
    output [1:0] col_out_157,
    output [1:0] col_out_158,
    output [1:0] col_out_159,
    output [1:0] col_out_160,
    output [1:0] col_out_161,
    output [1:0] col_out_162,
    output [1:0] col_out_163,
    output [1:0] col_out_164,
    output [1:0] col_out_165,
    output [1:0] col_out_166,
    output [1:0] col_out_167,
    output [1:0] col_out_168,
    output [1:0] col_out_169,
    output [1:0] col_out_170,
    output [1:0] col_out_171,
    output [1:0] col_out_172,
    output [1:0] col_out_173,
    output [1:0] col_out_174,
    output [1:0] col_out_175,
    output [1:0] col_out_176,
    output [1:0] col_out_177,
    output [1:0] col_out_178,
    output [1:0] col_out_179,
    output [1:0] col_out_180,
    output [1:0] col_out_181,
    output [1:0] col_out_182,
    output [1:0] col_out_183,
    output [1:0] col_out_184,
    output [1:0] col_out_185,
    output [1:0] col_out_186,
    output [1:0] col_out_187,
    output [1:0] col_out_188,
    output [1:0] col_out_189,
    output [1:0] col_out_190,
    output [1:0] col_out_191,
    output [1:0] col_out_192,
    output [1:0] col_out_193,
    output [1:0] col_out_194,
    output [1:0] col_out_195,
    output [1:0] col_out_196,
    output [1:0] col_out_197,
    output [1:0] col_out_198,
    output [1:0] col_out_199,
    output [1:0] col_out_200,
    output [1:0] col_out_201,
    output [1:0] col_out_202,
    output [1:0] col_out_203,
    output [1:0] col_out_204,
    output [1:0] col_out_205,
    output [1:0] col_out_206,
    output [1:0] col_out_207,
    output [1:0] col_out_208,
    output [1:0] col_out_209,
    output [1:0] col_out_210,
    output [1:0] col_out_211,
    output [1:0] col_out_212,
    output [1:0] col_out_213,
    output [1:0] col_out_214,
    output [1:0] col_out_215,
    output [1:0] col_out_216,
    output [1:0] col_out_217,
    output [1:0] col_out_218,
    output [1:0] col_out_219,
    output [1:0] col_out_220,
    output [1:0] col_out_221,
    output [1:0] col_out_222,
    output [1:0] col_out_223,
    output [1:0] col_out_224,
    output [1:0] col_out_225,
    output [1:0] col_out_226,
    output [1:0] col_out_227,
    output [1:0] col_out_228,
    output [1:0] col_out_229,
    output [1:0] col_out_230,
    output [1:0] col_out_231,
    output [1:0] col_out_232,
    output [1:0] col_out_233,
    output [1:0] col_out_234,
    output [1:0] col_out_235,
    output [1:0] col_out_236,
    output [1:0] col_out_237,
    output [1:0] col_out_238,
    output [1:0] col_out_239,
    output [1:0] col_out_240,
    output [1:0] col_out_241,
    output [1:0] col_out_242,
    output [1:0] col_out_243,
    output [1:0] col_out_244,
    output [1:0] col_out_245,
    output [1:0] col_out_246,
    output [1:0] col_out_247,
    output [1:0] col_out_248,
    output [1:0] col_out_249,
    output [1:0] col_out_250,
    output [1:0] col_out_251,
    output [1:0] col_out_252,
    output [1:0] col_out_253,
    output [1:0] col_out_254,
    output [1:0] col_out_255,
    output [1:0] col_out_256,
    output [1:0] col_out_257,
    output [1:0] col_out_258,
    output [1:0] col_out_259,
    output [1:0] col_out_260,
    output [1:0] col_out_261,
    output [1:0] col_out_262,
    output [1:0] col_out_263,
    output [1:0] col_out_264,
    output [1:0] col_out_265,
    output [1:0] col_out_266,
    output [1:0] col_out_267,
    output [1:0] col_out_268,
    output [1:0] col_out_269,
    output [1:0] col_out_270,
    output [1:0] col_out_271,
    output [1:0] col_out_272,
    output [1:0] col_out_273,
    output [1:0] col_out_274,
    output [1:0] col_out_275,
    output [1:0] col_out_276,
    output [1:0] col_out_277,
    output [1:0] col_out_278,
    output [1:0] col_out_279,
    output [1:0] col_out_280,
    output [1:0] col_out_281,
    output [1:0] col_out_282,
    output [1:0] col_out_283,
    output [1:0] col_out_284,
    output [1:0] col_out_285,
    output [1:0] col_out_286,
    output [1:0] col_out_287,
    output [1:0] col_out_288,
    output [1:0] col_out_289,
    output [1:0] col_out_290,
    output [1:0] col_out_291,
    output [1:0] col_out_292,
    output [1:0] col_out_293,
    output [1:0] col_out_294,
    output [1:0] col_out_295,
    output [1:0] col_out_296,
    output [1:0] col_out_297,
    output [1:0] col_out_298,
    output [1:0] col_out_299,
    output [1:0] col_out_300,
    output [1:0] col_out_301,
    output [1:0] col_out_302,
    output [1:0] col_out_303,
    output [1:0] col_out_304,
    output [1:0] col_out_305,
    output [1:0] col_out_306,
    output [1:0] col_out_307,
    output [1:0] col_out_308,
    output [1:0] col_out_309,
    output [1:0] col_out_310,
    output [1:0] col_out_311,
    output [1:0] col_out_312,
    output [1:0] col_out_313,
    output [1:0] col_out_314,
    output [1:0] col_out_315,
    output [1:0] col_out_316,
    output [1:0] col_out_317,
    output [1:0] col_out_318,
    output [1:0] col_out_319,
    output [1:0] col_out_320,
    output [1:0] col_out_321,
    output [1:0] col_out_322,
    output [1:0] col_out_323,
    output [1:0] col_out_324,
    output [1:0] col_out_325,
    output [1:0] col_out_326,
    output [1:0] col_out_327,
    output [1:0] col_out_328,
    output [1:0] col_out_329,
    output [1:0] col_out_330,
    output [1:0] col_out_331,
    output [1:0] col_out_332,
    output [1:0] col_out_333,
    output [1:0] col_out_334,
    output [1:0] col_out_335,
    output [1:0] col_out_336,
    output [1:0] col_out_337,
    output [1:0] col_out_338,
    output [1:0] col_out_339,
    output [1:0] col_out_340,
    output [1:0] col_out_341,
    output [1:0] col_out_342,
    output [1:0] col_out_343,
    output [1:0] col_out_344,
    output [1:0] col_out_345,
    output [1:0] col_out_346,
    output [1:0] col_out_347,
    output [1:0] col_out_348,
    output [1:0] col_out_349,
    output [1:0] col_out_350,
    output [1:0] col_out_351,
    output [1:0] col_out_352,
    output [1:0] col_out_353,
    output [1:0] col_out_354,
    output [1:0] col_out_355,
    output [1:0] col_out_356,
    output [1:0] col_out_357,
    output [1:0] col_out_358,
    output [1:0] col_out_359,
    output [1:0] col_out_360,
    output [1:0] col_out_361,
    output [1:0] col_out_362,
    output [1:0] col_out_363,
    output [1:0] col_out_364,
    output [1:0] col_out_365,
    output [1:0] col_out_366,
    output [1:0] col_out_367,
    output [1:0] col_out_368,
    output [1:0] col_out_369,
    output [1:0] col_out_370,
    output [1:0] col_out_371,
    output [1:0] col_out_372,
    output [1:0] col_out_373,
    output [1:0] col_out_374,
    output [1:0] col_out_375,
    output [1:0] col_out_376,
    output [1:0] col_out_377,
    output [1:0] col_out_378,
    output [1:0] col_out_379,
    output [1:0] col_out_380,
    output [1:0] col_out_381,
    output [1:0] col_out_382,
    output [1:0] col_out_383,
    output [1:0] col_out_384,
    output [1:0] col_out_385,
    output [1:0] col_out_386,
    output [1:0] col_out_387,
    output [1:0] col_out_388,
    output [1:0] col_out_389,
    output [1:0] col_out_390,
    output [1:0] col_out_391,
    output [1:0] col_out_392,
    output [1:0] col_out_393,
    output [1:0] col_out_394,
    output [1:0] col_out_395,
    output [1:0] col_out_396,
    output [1:0] col_out_397,
    output [1:0] col_out_398,
    output [1:0] col_out_399,
    output [1:0] col_out_400,
    output [1:0] col_out_401,
    output [1:0] col_out_402,
    output [1:0] col_out_403,
    output [1:0] col_out_404,
    output [1:0] col_out_405,
    output [1:0] col_out_406,
    output [1:0] col_out_407,
    output [1:0] col_out_408,
    output [1:0] col_out_409,
    output [1:0] col_out_410,
    output [1:0] col_out_411,
    output [1:0] col_out_412,
    output [1:0] col_out_413,
    output [1:0] col_out_414,
    output [1:0] col_out_415,
    output [1:0] col_out_416,
    output [1:0] col_out_417,
    output [1:0] col_out_418,
    output [1:0] col_out_419,
    output [1:0] col_out_420,
    output [1:0] col_out_421,
    output [1:0] col_out_422,
    output [1:0] col_out_423,
    output [1:0] col_out_424,
    output [1:0] col_out_425,
    output [1:0] col_out_426,
    output [1:0] col_out_427,
    output [1:0] col_out_428,
    output [1:0] col_out_429,
    output [1:0] col_out_430,
    output [1:0] col_out_431,
    output [1:0] col_out_432,
    output [1:0] col_out_433,
    output [1:0] col_out_434,
    output [1:0] col_out_435,
    output [1:0] col_out_436,
    output [1:0] col_out_437,
    output [1:0] col_out_438,
    output [1:0] col_out_439,
    output [1:0] col_out_440,
    output [1:0] col_out_441,
    output [1:0] col_out_442,
    output [1:0] col_out_443,
    output [1:0] col_out_444,
    output [1:0] col_out_445,
    output [1:0] col_out_446,
    output [1:0] col_out_447,
    output [1:0] col_out_448,
    output [1:0] col_out_449,
    output [1:0] col_out_450,
    output [1:0] col_out_451,
    output [1:0] col_out_452,
    output [1:0] col_out_453,
    output [1:0] col_out_454,
    output [1:0] col_out_455,
    output [1:0] col_out_456,
    output [1:0] col_out_457,
    output [1:0] col_out_458,
    output [1:0] col_out_459,
    output [1:0] col_out_460,
    output [1:0] col_out_461,
    output [1:0] col_out_462,
    output [1:0] col_out_463,
    output [1:0] col_out_464,
    output [1:0] col_out_465,
    output [1:0] col_out_466,
    output [1:0] col_out_467,
    output [1:0] col_out_468,
    output [1:0] col_out_469,
    output [1:0] col_out_470,
    output [1:0] col_out_471,
    output [1:0] col_out_472,
    output [1:0] col_out_473,
    output [1:0] col_out_474,
    output [1:0] col_out_475,
    output [1:0] col_out_476,
    output [1:0] col_out_477,
    output [1:0] col_out_478,
    output [1:0] col_out_479,
    output [1:0] col_out_480,
    output [1:0] col_out_481,
    output [1:0] col_out_482,
    output [1:0] col_out_483,
    output [1:0] col_out_484,
    output [1:0] col_out_485,
    output [1:0] col_out_486,
    output [1:0] col_out_487,
    output [1:0] col_out_488,
    output [1:0] col_out_489,
    output [1:0] col_out_490,
    output [1:0] col_out_491,
    output [1:0] col_out_492,
    output [1:0] col_out_493,
    output [1:0] col_out_494,
    output [1:0] col_out_495,
    output [1:0] col_out_496,
    output [1:0] col_out_497,
    output [1:0] col_out_498,
    output [1:0] col_out_499,
    output [1:0] col_out_500,
    output [1:0] col_out_501,
    output [1:0] col_out_502,
    output [1:0] col_out_503,
    output [1:0] col_out_504,
    output [1:0] col_out_505,
    output [1:0] col_out_506,
    output [1:0] col_out_507,
    output [1:0] col_out_508,
    output [1:0] col_out_509,
    output [1:0] col_out_510,
    output [1:0] col_out_511,
    output [1:0] col_out_512,
    output [1:0] col_out_513,
    output [1:0] col_out_514,
    output [1:0] col_out_515,
    output [1:0] col_out_516,
    output [1:0] col_out_517,
    output [1:0] col_out_518,
    output [1:0] col_out_519,
    output [1:0] col_out_520,
    output [1:0] col_out_521,
    output [1:0] col_out_522,
    output [1:0] col_out_523,
    output [1:0] col_out_524,
    output [1:0] col_out_525,
    output [1:0] col_out_526,
    output [1:0] col_out_527,
    output [1:0] col_out_528,
    output [1:0] col_out_529,
    output [1:0] col_out_530,
    output [1:0] col_out_531,
    output [1:0] col_out_532,
    output [1:0] col_out_533,
    output [1:0] col_out_534,
    output [1:0] col_out_535,
    output [1:0] col_out_536,
    output [1:0] col_out_537,
    output [1:0] col_out_538,
    output [1:0] col_out_539,
    output [1:0] col_out_540,
    output [1:0] col_out_541,
    output [1:0] col_out_542,
    output [1:0] col_out_543,
    output [1:0] col_out_544,
    output [1:0] col_out_545,
    output [1:0] col_out_546,
    output [1:0] col_out_547,
    output [1:0] col_out_548,
    output [1:0] col_out_549,
    output [1:0] col_out_550,
    output [1:0] col_out_551,
    output [1:0] col_out_552,
    output [1:0] col_out_553,
    output [1:0] col_out_554,
    output [1:0] col_out_555,
    output [1:0] col_out_556,
    output [1:0] col_out_557,
    output [1:0] col_out_558,
    output [1:0] col_out_559,
    output [1:0] col_out_560,
    output [1:0] col_out_561,
    output [1:0] col_out_562,
    output [1:0] col_out_563,
    output [1:0] col_out_564,
    output [1:0] col_out_565,
    output [1:0] col_out_566,
    output [1:0] col_out_567,
    output [1:0] col_out_568,
    output [1:0] col_out_569,
    output [1:0] col_out_570,
    output [1:0] col_out_571,
    output [1:0] col_out_572,
    output [1:0] col_out_573,
    output [1:0] col_out_574,
    output [1:0] col_out_575,
    output [1:0] col_out_576,
    output [1:0] col_out_577,
    output [1:0] col_out_578,
    output [1:0] col_out_579,
    output [1:0] col_out_580,
    output [1:0] col_out_581,
    output [1:0] col_out_582,
    output [1:0] col_out_583,
    output [1:0] col_out_584,
    output [1:0] col_out_585,
    output [1:0] col_out_586,
    output [1:0] col_out_587,
    output [1:0] col_out_588,
    output [1:0] col_out_589,
    output [1:0] col_out_590,
    output [1:0] col_out_591,
    output [1:0] col_out_592,
    output [1:0] col_out_593,
    output [1:0] col_out_594,
    output [1:0] col_out_595,
    output [1:0] col_out_596,
    output [1:0] col_out_597,
    output [1:0] col_out_598,
    output [1:0] col_out_599,
    output [1:0] col_out_600,
    output [1:0] col_out_601,
    output [1:0] col_out_602,
    output [1:0] col_out_603,
    output [1:0] col_out_604,
    output [1:0] col_out_605,
    output [1:0] col_out_606,
    output [1:0] col_out_607,
    output [1:0] col_out_608,
    output [1:0] col_out_609,
    output [1:0] col_out_610,
    output [1:0] col_out_611,
    output [1:0] col_out_612,
    output [1:0] col_out_613,
    output [1:0] col_out_614,
    output [1:0] col_out_615,
    output [1:0] col_out_616,
    output [1:0] col_out_617,
    output [1:0] col_out_618,
    output [1:0] col_out_619,
    output [1:0] col_out_620,
    output [1:0] col_out_621,
    output [1:0] col_out_622,
    output [1:0] col_out_623,
    output [1:0] col_out_624,
    output [1:0] col_out_625,
    output [1:0] col_out_626,
    output [1:0] col_out_627,
    output [1:0] col_out_628,
    output [1:0] col_out_629,
    output [1:0] col_out_630,
    output [1:0] col_out_631,
    output [1:0] col_out_632,
    output [1:0] col_out_633,
    output [1:0] col_out_634,
    output [1:0] col_out_635,
    output [1:0] col_out_636,
    output [1:0] col_out_637,
    output [1:0] col_out_638,
    output [1:0] col_out_639,
    output [1:0] col_out_640,
    output [1:0] col_out_641,
    output [1:0] col_out_642,
    output [1:0] col_out_643,
    output [1:0] col_out_644,
    output [1:0] col_out_645,
    output [1:0] col_out_646,
    output [1:0] col_out_647,
    output [1:0] col_out_648,
    output [1:0] col_out_649,
    output [1:0] col_out_650,
    output [1:0] col_out_651,
    output [1:0] col_out_652,
    output [1:0] col_out_653,
    output [1:0] col_out_654,
    output [1:0] col_out_655,
    output [1:0] col_out_656,
    output [1:0] col_out_657,
    output [1:0] col_out_658,
    output [1:0] col_out_659,
    output [1:0] col_out_660,
    output [1:0] col_out_661,
    output [1:0] col_out_662,
    output [1:0] col_out_663,
    output [1:0] col_out_664,
    output [1:0] col_out_665,
    output [1:0] col_out_666,
    output [1:0] col_out_667,
    output [1:0] col_out_668,
    output [1:0] col_out_669,
    output [1:0] col_out_670,
    output [1:0] col_out_671,
    output [1:0] col_out_672,
    output [1:0] col_out_673,
    output [1:0] col_out_674,
    output [1:0] col_out_675,
    output [1:0] col_out_676,
    output [1:0] col_out_677,
    output [1:0] col_out_678,
    output [1:0] col_out_679,
    output [1:0] col_out_680,
    output [1:0] col_out_681,
    output [1:0] col_out_682,
    output [1:0] col_out_683,
    output [1:0] col_out_684,
    output [1:0] col_out_685,
    output [1:0] col_out_686,
    output [1:0] col_out_687,
    output [1:0] col_out_688,
    output [1:0] col_out_689,
    output [1:0] col_out_690,
    output [1:0] col_out_691,
    output [1:0] col_out_692,
    output [1:0] col_out_693,
    output [1:0] col_out_694,
    output [1:0] col_out_695,
    output [1:0] col_out_696,
    output [1:0] col_out_697,
    output [1:0] col_out_698,
    output [1:0] col_out_699,
    output [1:0] col_out_700,
    output [1:0] col_out_701,
    output [1:0] col_out_702,
    output [1:0] col_out_703,
    output [1:0] col_out_704,
    output [1:0] col_out_705,
    output [1:0] col_out_706,
    output [1:0] col_out_707,
    output [1:0] col_out_708,
    output [1:0] col_out_709,
    output [1:0] col_out_710,
    output [1:0] col_out_711,
    output [1:0] col_out_712,
    output [1:0] col_out_713,
    output [1:0] col_out_714,
    output [1:0] col_out_715,
    output [1:0] col_out_716,
    output [1:0] col_out_717,
    output [1:0] col_out_718,
    output [1:0] col_out_719,
    output [1:0] col_out_720,
    output [1:0] col_out_721,
    output [1:0] col_out_722,
    output [1:0] col_out_723,
    output [1:0] col_out_724,
    output [1:0] col_out_725,
    output [1:0] col_out_726,
    output [1:0] col_out_727,
    output [1:0] col_out_728,
    output [1:0] col_out_729,
    output [1:0] col_out_730,
    output [1:0] col_out_731,
    output [1:0] col_out_732,
    output [1:0] col_out_733,
    output [1:0] col_out_734,
    output [1:0] col_out_735,
    output [1:0] col_out_736,
    output [1:0] col_out_737,
    output [1:0] col_out_738,
    output [1:0] col_out_739,
    output [1:0] col_out_740,
    output [1:0] col_out_741,
    output [1:0] col_out_742,
    output [1:0] col_out_743,
    output [1:0] col_out_744,
    output [1:0] col_out_745,
    output [1:0] col_out_746,
    output [1:0] col_out_747,
    output [1:0] col_out_748,
    output [1:0] col_out_749,
    output [1:0] col_out_750,
    output [1:0] col_out_751,
    output [1:0] col_out_752,
    output [1:0] col_out_753,
    output [1:0] col_out_754,
    output [1:0] col_out_755,
    output [1:0] col_out_756,
    output [1:0] col_out_757,
    output [1:0] col_out_758,
    output [1:0] col_out_759,
    output [1:0] col_out_760,
    output [1:0] col_out_761,
    output [1:0] col_out_762,
    output [1:0] col_out_763,
    output [1:0] col_out_764,
    output [1:0] col_out_765,
    output [1:0] col_out_766,
    output [1:0] col_out_767,
    output [1:0] col_out_768,
    output [1:0] col_out_769,
    output [1:0] col_out_770,
    output [1:0] col_out_771,
    output [1:0] col_out_772,
    output [1:0] col_out_773,
    output [1:0] col_out_774,
    output [1:0] col_out_775,
    output [1:0] col_out_776,
    output [1:0] col_out_777,
    output [1:0] col_out_778,
    output [1:0] col_out_779,
    output [1:0] col_out_780,
    output [1:0] col_out_781,
    output [1:0] col_out_782,
    output [1:0] col_out_783,
    output [1:0] col_out_784,
    output [1:0] col_out_785,
    output [1:0] col_out_786,
    output [1:0] col_out_787,
    output [1:0] col_out_788,
    output [1:0] col_out_789,
    output [1:0] col_out_790,
    output [1:0] col_out_791,
    output [1:0] col_out_792,
    output [1:0] col_out_793,
    output [1:0] col_out_794,
    output [1:0] col_out_795,
    output [1:0] col_out_796,
    output [1:0] col_out_797,
    output [1:0] col_out_798,
    output [1:0] col_out_799,
    output [1:0] col_out_800,
    output [1:0] col_out_801,
    output [1:0] col_out_802,
    output [1:0] col_out_803,
    output [1:0] col_out_804,
    output [1:0] col_out_805,
    output [1:0] col_out_806,
    output [1:0] col_out_807,
    output [1:0] col_out_808,
    output [1:0] col_out_809,
    output [1:0] col_out_810,
    output [1:0] col_out_811,
    output [1:0] col_out_812,
    output [1:0] col_out_813,
    output [1:0] col_out_814,
    output [1:0] col_out_815,
    output [1:0] col_out_816,
    output [1:0] col_out_817,
    output [1:0] col_out_818,
    output [1:0] col_out_819,
    output [1:0] col_out_820,
    output [1:0] col_out_821,
    output [1:0] col_out_822,
    output [1:0] col_out_823,
    output [1:0] col_out_824,
    output [1:0] col_out_825,
    output [1:0] col_out_826,
    output [1:0] col_out_827,
    output [1:0] col_out_828,
    output [1:0] col_out_829,
    output [1:0] col_out_830,
    output [1:0] col_out_831,
    output [1:0] col_out_832,
    output [1:0] col_out_833,
    output [1:0] col_out_834,
    output [1:0] col_out_835,
    output [1:0] col_out_836,
    output [1:0] col_out_837,
    output [1:0] col_out_838,
    output [1:0] col_out_839,
    output [1:0] col_out_840,
    output [1:0] col_out_841,
    output [1:0] col_out_842,
    output [1:0] col_out_843,
    output [1:0] col_out_844,
    output [1:0] col_out_845,
    output [1:0] col_out_846,
    output [1:0] col_out_847,
    output [1:0] col_out_848,
    output [1:0] col_out_849,
    output [1:0] col_out_850,
    output [1:0] col_out_851,
    output [1:0] col_out_852,
    output [1:0] col_out_853,
    output [1:0] col_out_854,
    output [1:0] col_out_855,
    output [1:0] col_out_856,
    output [1:0] col_out_857,
    output [1:0] col_out_858,
    output [1:0] col_out_859,
    output [1:0] col_out_860,
    output [1:0] col_out_861,
    output [1:0] col_out_862,
    output [1:0] col_out_863,
    output [1:0] col_out_864,
    output [1:0] col_out_865,
    output [1:0] col_out_866,
    output [1:0] col_out_867,
    output [1:0] col_out_868,
    output [1:0] col_out_869,
    output [1:0] col_out_870,
    output [1:0] col_out_871,
    output [1:0] col_out_872,
    output [1:0] col_out_873,
    output [1:0] col_out_874,
    output [1:0] col_out_875,
    output [1:0] col_out_876,
    output [1:0] col_out_877,
    output [1:0] col_out_878,
    output [1:0] col_out_879,
    output [1:0] col_out_880,
    output [1:0] col_out_881,
    output [1:0] col_out_882,
    output [1:0] col_out_883,
    output [1:0] col_out_884,
    output [1:0] col_out_885,
    output [1:0] col_out_886,
    output [1:0] col_out_887,
    output [1:0] col_out_888,
    output [1:0] col_out_889,
    output [1:0] col_out_890,
    output [1:0] col_out_891,
    output [1:0] col_out_892,
    output [1:0] col_out_893,
    output [1:0] col_out_894,
    output [1:0] col_out_895,
    output [1:0] col_out_896,
    output [1:0] col_out_897,
    output [1:0] col_out_898,
    output [1:0] col_out_899,
    output [1:0] col_out_900,
    output [1:0] col_out_901,
    output [1:0] col_out_902,
    output [1:0] col_out_903,
    output [1:0] col_out_904,
    output [1:0] col_out_905,
    output [1:0] col_out_906,
    output [1:0] col_out_907,
    output [1:0] col_out_908,
    output [1:0] col_out_909,
    output [1:0] col_out_910,
    output [1:0] col_out_911,
    output [1:0] col_out_912,
    output [1:0] col_out_913,
    output [1:0] col_out_914,
    output [1:0] col_out_915,
    output [1:0] col_out_916,
    output [1:0] col_out_917,
    output [1:0] col_out_918,
    output [1:0] col_out_919,
    output [1:0] col_out_920,
    output [1:0] col_out_921,
    output [1:0] col_out_922,
    output [1:0] col_out_923,
    output [1:0] col_out_924,
    output [1:0] col_out_925,
    output [1:0] col_out_926,
    output [1:0] col_out_927,
    output [1:0] col_out_928,
    output [1:0] col_out_929,
    output [1:0] col_out_930,
    output [1:0] col_out_931,
    output [1:0] col_out_932,
    output [1:0] col_out_933,
    output [1:0] col_out_934,
    output [1:0] col_out_935,
    output [1:0] col_out_936,
    output [1:0] col_out_937,
    output [1:0] col_out_938,
    output [1:0] col_out_939,
    output [1:0] col_out_940,
    output [1:0] col_out_941,
    output [1:0] col_out_942,
    output [1:0] col_out_943,
    output [1:0] col_out_944,
    output [1:0] col_out_945,
    output [1:0] col_out_946,
    output [1:0] col_out_947,
    output [1:0] col_out_948,
    output [1:0] col_out_949,
    output [1:0] col_out_950,
    output [1:0] col_out_951,
    output [1:0] col_out_952,
    output [1:0] col_out_953,
    output [1:0] col_out_954,
    output [1:0] col_out_955,
    output [1:0] col_out_956,
    output [1:0] col_out_957,
    output [1:0] col_out_958,
    output [1:0] col_out_959,
    output [1:0] col_out_960,
    output [1:0] col_out_961,
    output [1:0] col_out_962,
    output [1:0] col_out_963,
    output [1:0] col_out_964,
    output [1:0] col_out_965,
    output [1:0] col_out_966,
    output [1:0] col_out_967,
    output [1:0] col_out_968,
    output [1:0] col_out_969,
    output [1:0] col_out_970,
    output [1:0] col_out_971,
    output [1:0] col_out_972,
    output [1:0] col_out_973,
    output [1:0] col_out_974,
    output [1:0] col_out_975,
    output [1:0] col_out_976,
    output [1:0] col_out_977,
    output [1:0] col_out_978,
    output [1:0] col_out_979,
    output [1:0] col_out_980,
    output [1:0] col_out_981,
    output [1:0] col_out_982,
    output [1:0] col_out_983,
    output [1:0] col_out_984,
    output [1:0] col_out_985,
    output [1:0] col_out_986,
    output [1:0] col_out_987,
    output [1:0] col_out_988,
    output [1:0] col_out_989,
    output [1:0] col_out_990,
    output [1:0] col_out_991,
    output [1:0] col_out_992,
    output [1:0] col_out_993,
    output [1:0] col_out_994,
    output [1:0] col_out_995,
    output [1:0] col_out_996,
    output [1:0] col_out_997,
    output [1:0] col_out_998,
    output [1:0] col_out_999,
    output [1:0] col_out_1000,
    output [1:0] col_out_1001,
    output [1:0] col_out_1002,
    output [1:0] col_out_1003,
    output [1:0] col_out_1004,
    output [1:0] col_out_1005,
    output [1:0] col_out_1006,
    output [1:0] col_out_1007,
    output [1:0] col_out_1008,
    output [1:0] col_out_1009,
    output [1:0] col_out_1010,
    output [1:0] col_out_1011,
    output [1:0] col_out_1012,
    output [1:0] col_out_1013,
    output [1:0] col_out_1014,
    output [1:0] col_out_1015,
    output [1:0] col_out_1016,
    output [1:0] col_out_1017,
    output [1:0] col_out_1018,
    output [1:0] col_out_1019,
    output [1:0] col_out_1020,
    output [1:0] col_out_1021,
    output [1:0] col_out_1022,
    output [1:0] col_out_1023,
    output [1:0] col_out_1024,
    output [1:0] col_out_1025,
    output [1:0] col_out_1026,
    output [1:0] col_out_1027,
    output [1:0] col_out_1028,
    output [1:0] col_out_1029,
    output [1:0] col_out_1030,
    output [1:0] col_out_1031,
    output [1:0] col_out_1032
);

// compressor_array_16_12_1033 Outputs
wire  [11:0]  u0_col_out_0;
wire  [11:0]  u0_col_out_1;
wire  [11:0]  u0_col_out_2;
wire  [11:0]  u0_col_out_3;
wire  [11:0]  u0_col_out_4;
wire  [11:0]  u0_col_out_5;
wire  [11:0]  u0_col_out_6;
wire  [11:0]  u0_col_out_7;
wire  [11:0]  u0_col_out_8;
wire  [11:0]  u0_col_out_9;
wire  [11:0]  u0_col_out_10;
wire  [11:0]  u0_col_out_11;
wire  [11:0]  u0_col_out_12;
wire  [11:0]  u0_col_out_13;
wire  [11:0]  u0_col_out_14;
wire  [11:0]  u0_col_out_15;
wire  [11:0]  u0_col_out_16;
wire  [11:0]  u0_col_out_17;
wire  [11:0]  u0_col_out_18;
wire  [11:0]  u0_col_out_19;
wire  [11:0]  u0_col_out_20;
wire  [11:0]  u0_col_out_21;
wire  [11:0]  u0_col_out_22;
wire  [11:0]  u0_col_out_23;
wire  [11:0]  u0_col_out_24;
wire  [11:0]  u0_col_out_25;
wire  [11:0]  u0_col_out_26;
wire  [11:0]  u0_col_out_27;
wire  [11:0]  u0_col_out_28;
wire  [11:0]  u0_col_out_29;
wire  [11:0]  u0_col_out_30;
wire  [11:0]  u0_col_out_31;
wire  [11:0]  u0_col_out_32;
wire  [11:0]  u0_col_out_33;
wire  [11:0]  u0_col_out_34;
wire  [11:0]  u0_col_out_35;
wire  [11:0]  u0_col_out_36;
wire  [11:0]  u0_col_out_37;
wire  [11:0]  u0_col_out_38;
wire  [11:0]  u0_col_out_39;
wire  [11:0]  u0_col_out_40;
wire  [11:0]  u0_col_out_41;
wire  [11:0]  u0_col_out_42;
wire  [11:0]  u0_col_out_43;
wire  [11:0]  u0_col_out_44;
wire  [11:0]  u0_col_out_45;
wire  [11:0]  u0_col_out_46;
wire  [11:0]  u0_col_out_47;
wire  [11:0]  u0_col_out_48;
wire  [11:0]  u0_col_out_49;
wire  [11:0]  u0_col_out_50;
wire  [11:0]  u0_col_out_51;
wire  [11:0]  u0_col_out_52;
wire  [11:0]  u0_col_out_53;
wire  [11:0]  u0_col_out_54;
wire  [11:0]  u0_col_out_55;
wire  [11:0]  u0_col_out_56;
wire  [11:0]  u0_col_out_57;
wire  [11:0]  u0_col_out_58;
wire  [11:0]  u0_col_out_59;
wire  [11:0]  u0_col_out_60;
wire  [11:0]  u0_col_out_61;
wire  [11:0]  u0_col_out_62;
wire  [11:0]  u0_col_out_63;
wire  [11:0]  u0_col_out_64;
wire  [11:0]  u0_col_out_65;
wire  [11:0]  u0_col_out_66;
wire  [11:0]  u0_col_out_67;
wire  [11:0]  u0_col_out_68;
wire  [11:0]  u0_col_out_69;
wire  [11:0]  u0_col_out_70;
wire  [11:0]  u0_col_out_71;
wire  [11:0]  u0_col_out_72;
wire  [11:0]  u0_col_out_73;
wire  [11:0]  u0_col_out_74;
wire  [11:0]  u0_col_out_75;
wire  [11:0]  u0_col_out_76;
wire  [11:0]  u0_col_out_77;
wire  [11:0]  u0_col_out_78;
wire  [11:0]  u0_col_out_79;
wire  [11:0]  u0_col_out_80;
wire  [11:0]  u0_col_out_81;
wire  [11:0]  u0_col_out_82;
wire  [11:0]  u0_col_out_83;
wire  [11:0]  u0_col_out_84;
wire  [11:0]  u0_col_out_85;
wire  [11:0]  u0_col_out_86;
wire  [11:0]  u0_col_out_87;
wire  [11:0]  u0_col_out_88;
wire  [11:0]  u0_col_out_89;
wire  [11:0]  u0_col_out_90;
wire  [11:0]  u0_col_out_91;
wire  [11:0]  u0_col_out_92;
wire  [11:0]  u0_col_out_93;
wire  [11:0]  u0_col_out_94;
wire  [11:0]  u0_col_out_95;
wire  [11:0]  u0_col_out_96;
wire  [11:0]  u0_col_out_97;
wire  [11:0]  u0_col_out_98;
wire  [11:0]  u0_col_out_99;
wire  [11:0]  u0_col_out_100;
wire  [11:0]  u0_col_out_101;
wire  [11:0]  u0_col_out_102;
wire  [11:0]  u0_col_out_103;
wire  [11:0]  u0_col_out_104;
wire  [11:0]  u0_col_out_105;
wire  [11:0]  u0_col_out_106;
wire  [11:0]  u0_col_out_107;
wire  [11:0]  u0_col_out_108;
wire  [11:0]  u0_col_out_109;
wire  [11:0]  u0_col_out_110;
wire  [11:0]  u0_col_out_111;
wire  [11:0]  u0_col_out_112;
wire  [11:0]  u0_col_out_113;
wire  [11:0]  u0_col_out_114;
wire  [11:0]  u0_col_out_115;
wire  [11:0]  u0_col_out_116;
wire  [11:0]  u0_col_out_117;
wire  [11:0]  u0_col_out_118;
wire  [11:0]  u0_col_out_119;
wire  [11:0]  u0_col_out_120;
wire  [11:0]  u0_col_out_121;
wire  [11:0]  u0_col_out_122;
wire  [11:0]  u0_col_out_123;
wire  [11:0]  u0_col_out_124;
wire  [11:0]  u0_col_out_125;
wire  [11:0]  u0_col_out_126;
wire  [11:0]  u0_col_out_127;
wire  [11:0]  u0_col_out_128;
wire  [11:0]  u0_col_out_129;
wire  [11:0]  u0_col_out_130;
wire  [11:0]  u0_col_out_131;
wire  [11:0]  u0_col_out_132;
wire  [11:0]  u0_col_out_133;
wire  [11:0]  u0_col_out_134;
wire  [11:0]  u0_col_out_135;
wire  [11:0]  u0_col_out_136;
wire  [11:0]  u0_col_out_137;
wire  [11:0]  u0_col_out_138;
wire  [11:0]  u0_col_out_139;
wire  [11:0]  u0_col_out_140;
wire  [11:0]  u0_col_out_141;
wire  [11:0]  u0_col_out_142;
wire  [11:0]  u0_col_out_143;
wire  [11:0]  u0_col_out_144;
wire  [11:0]  u0_col_out_145;
wire  [11:0]  u0_col_out_146;
wire  [11:0]  u0_col_out_147;
wire  [11:0]  u0_col_out_148;
wire  [11:0]  u0_col_out_149;
wire  [11:0]  u0_col_out_150;
wire  [11:0]  u0_col_out_151;
wire  [11:0]  u0_col_out_152;
wire  [11:0]  u0_col_out_153;
wire  [11:0]  u0_col_out_154;
wire  [11:0]  u0_col_out_155;
wire  [11:0]  u0_col_out_156;
wire  [11:0]  u0_col_out_157;
wire  [11:0]  u0_col_out_158;
wire  [11:0]  u0_col_out_159;
wire  [11:0]  u0_col_out_160;
wire  [11:0]  u0_col_out_161;
wire  [11:0]  u0_col_out_162;
wire  [11:0]  u0_col_out_163;
wire  [11:0]  u0_col_out_164;
wire  [11:0]  u0_col_out_165;
wire  [11:0]  u0_col_out_166;
wire  [11:0]  u0_col_out_167;
wire  [11:0]  u0_col_out_168;
wire  [11:0]  u0_col_out_169;
wire  [11:0]  u0_col_out_170;
wire  [11:0]  u0_col_out_171;
wire  [11:0]  u0_col_out_172;
wire  [11:0]  u0_col_out_173;
wire  [11:0]  u0_col_out_174;
wire  [11:0]  u0_col_out_175;
wire  [11:0]  u0_col_out_176;
wire  [11:0]  u0_col_out_177;
wire  [11:0]  u0_col_out_178;
wire  [11:0]  u0_col_out_179;
wire  [11:0]  u0_col_out_180;
wire  [11:0]  u0_col_out_181;
wire  [11:0]  u0_col_out_182;
wire  [11:0]  u0_col_out_183;
wire  [11:0]  u0_col_out_184;
wire  [11:0]  u0_col_out_185;
wire  [11:0]  u0_col_out_186;
wire  [11:0]  u0_col_out_187;
wire  [11:0]  u0_col_out_188;
wire  [11:0]  u0_col_out_189;
wire  [11:0]  u0_col_out_190;
wire  [11:0]  u0_col_out_191;
wire  [11:0]  u0_col_out_192;
wire  [11:0]  u0_col_out_193;
wire  [11:0]  u0_col_out_194;
wire  [11:0]  u0_col_out_195;
wire  [11:0]  u0_col_out_196;
wire  [11:0]  u0_col_out_197;
wire  [11:0]  u0_col_out_198;
wire  [11:0]  u0_col_out_199;
wire  [11:0]  u0_col_out_200;
wire  [11:0]  u0_col_out_201;
wire  [11:0]  u0_col_out_202;
wire  [11:0]  u0_col_out_203;
wire  [11:0]  u0_col_out_204;
wire  [11:0]  u0_col_out_205;
wire  [11:0]  u0_col_out_206;
wire  [11:0]  u0_col_out_207;
wire  [11:0]  u0_col_out_208;
wire  [11:0]  u0_col_out_209;
wire  [11:0]  u0_col_out_210;
wire  [11:0]  u0_col_out_211;
wire  [11:0]  u0_col_out_212;
wire  [11:0]  u0_col_out_213;
wire  [11:0]  u0_col_out_214;
wire  [11:0]  u0_col_out_215;
wire  [11:0]  u0_col_out_216;
wire  [11:0]  u0_col_out_217;
wire  [11:0]  u0_col_out_218;
wire  [11:0]  u0_col_out_219;
wire  [11:0]  u0_col_out_220;
wire  [11:0]  u0_col_out_221;
wire  [11:0]  u0_col_out_222;
wire  [11:0]  u0_col_out_223;
wire  [11:0]  u0_col_out_224;
wire  [11:0]  u0_col_out_225;
wire  [11:0]  u0_col_out_226;
wire  [11:0]  u0_col_out_227;
wire  [11:0]  u0_col_out_228;
wire  [11:0]  u0_col_out_229;
wire  [11:0]  u0_col_out_230;
wire  [11:0]  u0_col_out_231;
wire  [11:0]  u0_col_out_232;
wire  [11:0]  u0_col_out_233;
wire  [11:0]  u0_col_out_234;
wire  [11:0]  u0_col_out_235;
wire  [11:0]  u0_col_out_236;
wire  [11:0]  u0_col_out_237;
wire  [11:0]  u0_col_out_238;
wire  [11:0]  u0_col_out_239;
wire  [11:0]  u0_col_out_240;
wire  [11:0]  u0_col_out_241;
wire  [11:0]  u0_col_out_242;
wire  [11:0]  u0_col_out_243;
wire  [11:0]  u0_col_out_244;
wire  [11:0]  u0_col_out_245;
wire  [11:0]  u0_col_out_246;
wire  [11:0]  u0_col_out_247;
wire  [11:0]  u0_col_out_248;
wire  [11:0]  u0_col_out_249;
wire  [11:0]  u0_col_out_250;
wire  [11:0]  u0_col_out_251;
wire  [11:0]  u0_col_out_252;
wire  [11:0]  u0_col_out_253;
wire  [11:0]  u0_col_out_254;
wire  [11:0]  u0_col_out_255;
wire  [11:0]  u0_col_out_256;
wire  [11:0]  u0_col_out_257;
wire  [11:0]  u0_col_out_258;
wire  [11:0]  u0_col_out_259;
wire  [11:0]  u0_col_out_260;
wire  [11:0]  u0_col_out_261;
wire  [11:0]  u0_col_out_262;
wire  [11:0]  u0_col_out_263;
wire  [11:0]  u0_col_out_264;
wire  [11:0]  u0_col_out_265;
wire  [11:0]  u0_col_out_266;
wire  [11:0]  u0_col_out_267;
wire  [11:0]  u0_col_out_268;
wire  [11:0]  u0_col_out_269;
wire  [11:0]  u0_col_out_270;
wire  [11:0]  u0_col_out_271;
wire  [11:0]  u0_col_out_272;
wire  [11:0]  u0_col_out_273;
wire  [11:0]  u0_col_out_274;
wire  [11:0]  u0_col_out_275;
wire  [11:0]  u0_col_out_276;
wire  [11:0]  u0_col_out_277;
wire  [11:0]  u0_col_out_278;
wire  [11:0]  u0_col_out_279;
wire  [11:0]  u0_col_out_280;
wire  [11:0]  u0_col_out_281;
wire  [11:0]  u0_col_out_282;
wire  [11:0]  u0_col_out_283;
wire  [11:0]  u0_col_out_284;
wire  [11:0]  u0_col_out_285;
wire  [11:0]  u0_col_out_286;
wire  [11:0]  u0_col_out_287;
wire  [11:0]  u0_col_out_288;
wire  [11:0]  u0_col_out_289;
wire  [11:0]  u0_col_out_290;
wire  [11:0]  u0_col_out_291;
wire  [11:0]  u0_col_out_292;
wire  [11:0]  u0_col_out_293;
wire  [11:0]  u0_col_out_294;
wire  [11:0]  u0_col_out_295;
wire  [11:0]  u0_col_out_296;
wire  [11:0]  u0_col_out_297;
wire  [11:0]  u0_col_out_298;
wire  [11:0]  u0_col_out_299;
wire  [11:0]  u0_col_out_300;
wire  [11:0]  u0_col_out_301;
wire  [11:0]  u0_col_out_302;
wire  [11:0]  u0_col_out_303;
wire  [11:0]  u0_col_out_304;
wire  [11:0]  u0_col_out_305;
wire  [11:0]  u0_col_out_306;
wire  [11:0]  u0_col_out_307;
wire  [11:0]  u0_col_out_308;
wire  [11:0]  u0_col_out_309;
wire  [11:0]  u0_col_out_310;
wire  [11:0]  u0_col_out_311;
wire  [11:0]  u0_col_out_312;
wire  [11:0]  u0_col_out_313;
wire  [11:0]  u0_col_out_314;
wire  [11:0]  u0_col_out_315;
wire  [11:0]  u0_col_out_316;
wire  [11:0]  u0_col_out_317;
wire  [11:0]  u0_col_out_318;
wire  [11:0]  u0_col_out_319;
wire  [11:0]  u0_col_out_320;
wire  [11:0]  u0_col_out_321;
wire  [11:0]  u0_col_out_322;
wire  [11:0]  u0_col_out_323;
wire  [11:0]  u0_col_out_324;
wire  [11:0]  u0_col_out_325;
wire  [11:0]  u0_col_out_326;
wire  [11:0]  u0_col_out_327;
wire  [11:0]  u0_col_out_328;
wire  [11:0]  u0_col_out_329;
wire  [11:0]  u0_col_out_330;
wire  [11:0]  u0_col_out_331;
wire  [11:0]  u0_col_out_332;
wire  [11:0]  u0_col_out_333;
wire  [11:0]  u0_col_out_334;
wire  [11:0]  u0_col_out_335;
wire  [11:0]  u0_col_out_336;
wire  [11:0]  u0_col_out_337;
wire  [11:0]  u0_col_out_338;
wire  [11:0]  u0_col_out_339;
wire  [11:0]  u0_col_out_340;
wire  [11:0]  u0_col_out_341;
wire  [11:0]  u0_col_out_342;
wire  [11:0]  u0_col_out_343;
wire  [11:0]  u0_col_out_344;
wire  [11:0]  u0_col_out_345;
wire  [11:0]  u0_col_out_346;
wire  [11:0]  u0_col_out_347;
wire  [11:0]  u0_col_out_348;
wire  [11:0]  u0_col_out_349;
wire  [11:0]  u0_col_out_350;
wire  [11:0]  u0_col_out_351;
wire  [11:0]  u0_col_out_352;
wire  [11:0]  u0_col_out_353;
wire  [11:0]  u0_col_out_354;
wire  [11:0]  u0_col_out_355;
wire  [11:0]  u0_col_out_356;
wire  [11:0]  u0_col_out_357;
wire  [11:0]  u0_col_out_358;
wire  [11:0]  u0_col_out_359;
wire  [11:0]  u0_col_out_360;
wire  [11:0]  u0_col_out_361;
wire  [11:0]  u0_col_out_362;
wire  [11:0]  u0_col_out_363;
wire  [11:0]  u0_col_out_364;
wire  [11:0]  u0_col_out_365;
wire  [11:0]  u0_col_out_366;
wire  [11:0]  u0_col_out_367;
wire  [11:0]  u0_col_out_368;
wire  [11:0]  u0_col_out_369;
wire  [11:0]  u0_col_out_370;
wire  [11:0]  u0_col_out_371;
wire  [11:0]  u0_col_out_372;
wire  [11:0]  u0_col_out_373;
wire  [11:0]  u0_col_out_374;
wire  [11:0]  u0_col_out_375;
wire  [11:0]  u0_col_out_376;
wire  [11:0]  u0_col_out_377;
wire  [11:0]  u0_col_out_378;
wire  [11:0]  u0_col_out_379;
wire  [11:0]  u0_col_out_380;
wire  [11:0]  u0_col_out_381;
wire  [11:0]  u0_col_out_382;
wire  [11:0]  u0_col_out_383;
wire  [11:0]  u0_col_out_384;
wire  [11:0]  u0_col_out_385;
wire  [11:0]  u0_col_out_386;
wire  [11:0]  u0_col_out_387;
wire  [11:0]  u0_col_out_388;
wire  [11:0]  u0_col_out_389;
wire  [11:0]  u0_col_out_390;
wire  [11:0]  u0_col_out_391;
wire  [11:0]  u0_col_out_392;
wire  [11:0]  u0_col_out_393;
wire  [11:0]  u0_col_out_394;
wire  [11:0]  u0_col_out_395;
wire  [11:0]  u0_col_out_396;
wire  [11:0]  u0_col_out_397;
wire  [11:0]  u0_col_out_398;
wire  [11:0]  u0_col_out_399;
wire  [11:0]  u0_col_out_400;
wire  [11:0]  u0_col_out_401;
wire  [11:0]  u0_col_out_402;
wire  [11:0]  u0_col_out_403;
wire  [11:0]  u0_col_out_404;
wire  [11:0]  u0_col_out_405;
wire  [11:0]  u0_col_out_406;
wire  [11:0]  u0_col_out_407;
wire  [11:0]  u0_col_out_408;
wire  [11:0]  u0_col_out_409;
wire  [11:0]  u0_col_out_410;
wire  [11:0]  u0_col_out_411;
wire  [11:0]  u0_col_out_412;
wire  [11:0]  u0_col_out_413;
wire  [11:0]  u0_col_out_414;
wire  [11:0]  u0_col_out_415;
wire  [11:0]  u0_col_out_416;
wire  [11:0]  u0_col_out_417;
wire  [11:0]  u0_col_out_418;
wire  [11:0]  u0_col_out_419;
wire  [11:0]  u0_col_out_420;
wire  [11:0]  u0_col_out_421;
wire  [11:0]  u0_col_out_422;
wire  [11:0]  u0_col_out_423;
wire  [11:0]  u0_col_out_424;
wire  [11:0]  u0_col_out_425;
wire  [11:0]  u0_col_out_426;
wire  [11:0]  u0_col_out_427;
wire  [11:0]  u0_col_out_428;
wire  [11:0]  u0_col_out_429;
wire  [11:0]  u0_col_out_430;
wire  [11:0]  u0_col_out_431;
wire  [11:0]  u0_col_out_432;
wire  [11:0]  u0_col_out_433;
wire  [11:0]  u0_col_out_434;
wire  [11:0]  u0_col_out_435;
wire  [11:0]  u0_col_out_436;
wire  [11:0]  u0_col_out_437;
wire  [11:0]  u0_col_out_438;
wire  [11:0]  u0_col_out_439;
wire  [11:0]  u0_col_out_440;
wire  [11:0]  u0_col_out_441;
wire  [11:0]  u0_col_out_442;
wire  [11:0]  u0_col_out_443;
wire  [11:0]  u0_col_out_444;
wire  [11:0]  u0_col_out_445;
wire  [11:0]  u0_col_out_446;
wire  [11:0]  u0_col_out_447;
wire  [11:0]  u0_col_out_448;
wire  [11:0]  u0_col_out_449;
wire  [11:0]  u0_col_out_450;
wire  [11:0]  u0_col_out_451;
wire  [11:0]  u0_col_out_452;
wire  [11:0]  u0_col_out_453;
wire  [11:0]  u0_col_out_454;
wire  [11:0]  u0_col_out_455;
wire  [11:0]  u0_col_out_456;
wire  [11:0]  u0_col_out_457;
wire  [11:0]  u0_col_out_458;
wire  [11:0]  u0_col_out_459;
wire  [11:0]  u0_col_out_460;
wire  [11:0]  u0_col_out_461;
wire  [11:0]  u0_col_out_462;
wire  [11:0]  u0_col_out_463;
wire  [11:0]  u0_col_out_464;
wire  [11:0]  u0_col_out_465;
wire  [11:0]  u0_col_out_466;
wire  [11:0]  u0_col_out_467;
wire  [11:0]  u0_col_out_468;
wire  [11:0]  u0_col_out_469;
wire  [11:0]  u0_col_out_470;
wire  [11:0]  u0_col_out_471;
wire  [11:0]  u0_col_out_472;
wire  [11:0]  u0_col_out_473;
wire  [11:0]  u0_col_out_474;
wire  [11:0]  u0_col_out_475;
wire  [11:0]  u0_col_out_476;
wire  [11:0]  u0_col_out_477;
wire  [11:0]  u0_col_out_478;
wire  [11:0]  u0_col_out_479;
wire  [11:0]  u0_col_out_480;
wire  [11:0]  u0_col_out_481;
wire  [11:0]  u0_col_out_482;
wire  [11:0]  u0_col_out_483;
wire  [11:0]  u0_col_out_484;
wire  [11:0]  u0_col_out_485;
wire  [11:0]  u0_col_out_486;
wire  [11:0]  u0_col_out_487;
wire  [11:0]  u0_col_out_488;
wire  [11:0]  u0_col_out_489;
wire  [11:0]  u0_col_out_490;
wire  [11:0]  u0_col_out_491;
wire  [11:0]  u0_col_out_492;
wire  [11:0]  u0_col_out_493;
wire  [11:0]  u0_col_out_494;
wire  [11:0]  u0_col_out_495;
wire  [11:0]  u0_col_out_496;
wire  [11:0]  u0_col_out_497;
wire  [11:0]  u0_col_out_498;
wire  [11:0]  u0_col_out_499;
wire  [11:0]  u0_col_out_500;
wire  [11:0]  u0_col_out_501;
wire  [11:0]  u0_col_out_502;
wire  [11:0]  u0_col_out_503;
wire  [11:0]  u0_col_out_504;
wire  [11:0]  u0_col_out_505;
wire  [11:0]  u0_col_out_506;
wire  [11:0]  u0_col_out_507;
wire  [11:0]  u0_col_out_508;
wire  [11:0]  u0_col_out_509;
wire  [11:0]  u0_col_out_510;
wire  [11:0]  u0_col_out_511;
wire  [11:0]  u0_col_out_512;
wire  [11:0]  u0_col_out_513;
wire  [11:0]  u0_col_out_514;
wire  [11:0]  u0_col_out_515;
wire  [11:0]  u0_col_out_516;
wire  [11:0]  u0_col_out_517;
wire  [11:0]  u0_col_out_518;
wire  [11:0]  u0_col_out_519;
wire  [11:0]  u0_col_out_520;
wire  [11:0]  u0_col_out_521;
wire  [11:0]  u0_col_out_522;
wire  [11:0]  u0_col_out_523;
wire  [11:0]  u0_col_out_524;
wire  [11:0]  u0_col_out_525;
wire  [11:0]  u0_col_out_526;
wire  [11:0]  u0_col_out_527;
wire  [11:0]  u0_col_out_528;
wire  [11:0]  u0_col_out_529;
wire  [11:0]  u0_col_out_530;
wire  [11:0]  u0_col_out_531;
wire  [11:0]  u0_col_out_532;
wire  [11:0]  u0_col_out_533;
wire  [11:0]  u0_col_out_534;
wire  [11:0]  u0_col_out_535;
wire  [11:0]  u0_col_out_536;
wire  [11:0]  u0_col_out_537;
wire  [11:0]  u0_col_out_538;
wire  [11:0]  u0_col_out_539;
wire  [11:0]  u0_col_out_540;
wire  [11:0]  u0_col_out_541;
wire  [11:0]  u0_col_out_542;
wire  [11:0]  u0_col_out_543;
wire  [11:0]  u0_col_out_544;
wire  [11:0]  u0_col_out_545;
wire  [11:0]  u0_col_out_546;
wire  [11:0]  u0_col_out_547;
wire  [11:0]  u0_col_out_548;
wire  [11:0]  u0_col_out_549;
wire  [11:0]  u0_col_out_550;
wire  [11:0]  u0_col_out_551;
wire  [11:0]  u0_col_out_552;
wire  [11:0]  u0_col_out_553;
wire  [11:0]  u0_col_out_554;
wire  [11:0]  u0_col_out_555;
wire  [11:0]  u0_col_out_556;
wire  [11:0]  u0_col_out_557;
wire  [11:0]  u0_col_out_558;
wire  [11:0]  u0_col_out_559;
wire  [11:0]  u0_col_out_560;
wire  [11:0]  u0_col_out_561;
wire  [11:0]  u0_col_out_562;
wire  [11:0]  u0_col_out_563;
wire  [11:0]  u0_col_out_564;
wire  [11:0]  u0_col_out_565;
wire  [11:0]  u0_col_out_566;
wire  [11:0]  u0_col_out_567;
wire  [11:0]  u0_col_out_568;
wire  [11:0]  u0_col_out_569;
wire  [11:0]  u0_col_out_570;
wire  [11:0]  u0_col_out_571;
wire  [11:0]  u0_col_out_572;
wire  [11:0]  u0_col_out_573;
wire  [11:0]  u0_col_out_574;
wire  [11:0]  u0_col_out_575;
wire  [11:0]  u0_col_out_576;
wire  [11:0]  u0_col_out_577;
wire  [11:0]  u0_col_out_578;
wire  [11:0]  u0_col_out_579;
wire  [11:0]  u0_col_out_580;
wire  [11:0]  u0_col_out_581;
wire  [11:0]  u0_col_out_582;
wire  [11:0]  u0_col_out_583;
wire  [11:0]  u0_col_out_584;
wire  [11:0]  u0_col_out_585;
wire  [11:0]  u0_col_out_586;
wire  [11:0]  u0_col_out_587;
wire  [11:0]  u0_col_out_588;
wire  [11:0]  u0_col_out_589;
wire  [11:0]  u0_col_out_590;
wire  [11:0]  u0_col_out_591;
wire  [11:0]  u0_col_out_592;
wire  [11:0]  u0_col_out_593;
wire  [11:0]  u0_col_out_594;
wire  [11:0]  u0_col_out_595;
wire  [11:0]  u0_col_out_596;
wire  [11:0]  u0_col_out_597;
wire  [11:0]  u0_col_out_598;
wire  [11:0]  u0_col_out_599;
wire  [11:0]  u0_col_out_600;
wire  [11:0]  u0_col_out_601;
wire  [11:0]  u0_col_out_602;
wire  [11:0]  u0_col_out_603;
wire  [11:0]  u0_col_out_604;
wire  [11:0]  u0_col_out_605;
wire  [11:0]  u0_col_out_606;
wire  [11:0]  u0_col_out_607;
wire  [11:0]  u0_col_out_608;
wire  [11:0]  u0_col_out_609;
wire  [11:0]  u0_col_out_610;
wire  [11:0]  u0_col_out_611;
wire  [11:0]  u0_col_out_612;
wire  [11:0]  u0_col_out_613;
wire  [11:0]  u0_col_out_614;
wire  [11:0]  u0_col_out_615;
wire  [11:0]  u0_col_out_616;
wire  [11:0]  u0_col_out_617;
wire  [11:0]  u0_col_out_618;
wire  [11:0]  u0_col_out_619;
wire  [11:0]  u0_col_out_620;
wire  [11:0]  u0_col_out_621;
wire  [11:0]  u0_col_out_622;
wire  [11:0]  u0_col_out_623;
wire  [11:0]  u0_col_out_624;
wire  [11:0]  u0_col_out_625;
wire  [11:0]  u0_col_out_626;
wire  [11:0]  u0_col_out_627;
wire  [11:0]  u0_col_out_628;
wire  [11:0]  u0_col_out_629;
wire  [11:0]  u0_col_out_630;
wire  [11:0]  u0_col_out_631;
wire  [11:0]  u0_col_out_632;
wire  [11:0]  u0_col_out_633;
wire  [11:0]  u0_col_out_634;
wire  [11:0]  u0_col_out_635;
wire  [11:0]  u0_col_out_636;
wire  [11:0]  u0_col_out_637;
wire  [11:0]  u0_col_out_638;
wire  [11:0]  u0_col_out_639;
wire  [11:0]  u0_col_out_640;
wire  [11:0]  u0_col_out_641;
wire  [11:0]  u0_col_out_642;
wire  [11:0]  u0_col_out_643;
wire  [11:0]  u0_col_out_644;
wire  [11:0]  u0_col_out_645;
wire  [11:0]  u0_col_out_646;
wire  [11:0]  u0_col_out_647;
wire  [11:0]  u0_col_out_648;
wire  [11:0]  u0_col_out_649;
wire  [11:0]  u0_col_out_650;
wire  [11:0]  u0_col_out_651;
wire  [11:0]  u0_col_out_652;
wire  [11:0]  u0_col_out_653;
wire  [11:0]  u0_col_out_654;
wire  [11:0]  u0_col_out_655;
wire  [11:0]  u0_col_out_656;
wire  [11:0]  u0_col_out_657;
wire  [11:0]  u0_col_out_658;
wire  [11:0]  u0_col_out_659;
wire  [11:0]  u0_col_out_660;
wire  [11:0]  u0_col_out_661;
wire  [11:0]  u0_col_out_662;
wire  [11:0]  u0_col_out_663;
wire  [11:0]  u0_col_out_664;
wire  [11:0]  u0_col_out_665;
wire  [11:0]  u0_col_out_666;
wire  [11:0]  u0_col_out_667;
wire  [11:0]  u0_col_out_668;
wire  [11:0]  u0_col_out_669;
wire  [11:0]  u0_col_out_670;
wire  [11:0]  u0_col_out_671;
wire  [11:0]  u0_col_out_672;
wire  [11:0]  u0_col_out_673;
wire  [11:0]  u0_col_out_674;
wire  [11:0]  u0_col_out_675;
wire  [11:0]  u0_col_out_676;
wire  [11:0]  u0_col_out_677;
wire  [11:0]  u0_col_out_678;
wire  [11:0]  u0_col_out_679;
wire  [11:0]  u0_col_out_680;
wire  [11:0]  u0_col_out_681;
wire  [11:0]  u0_col_out_682;
wire  [11:0]  u0_col_out_683;
wire  [11:0]  u0_col_out_684;
wire  [11:0]  u0_col_out_685;
wire  [11:0]  u0_col_out_686;
wire  [11:0]  u0_col_out_687;
wire  [11:0]  u0_col_out_688;
wire  [11:0]  u0_col_out_689;
wire  [11:0]  u0_col_out_690;
wire  [11:0]  u0_col_out_691;
wire  [11:0]  u0_col_out_692;
wire  [11:0]  u0_col_out_693;
wire  [11:0]  u0_col_out_694;
wire  [11:0]  u0_col_out_695;
wire  [11:0]  u0_col_out_696;
wire  [11:0]  u0_col_out_697;
wire  [11:0]  u0_col_out_698;
wire  [11:0]  u0_col_out_699;
wire  [11:0]  u0_col_out_700;
wire  [11:0]  u0_col_out_701;
wire  [11:0]  u0_col_out_702;
wire  [11:0]  u0_col_out_703;
wire  [11:0]  u0_col_out_704;
wire  [11:0]  u0_col_out_705;
wire  [11:0]  u0_col_out_706;
wire  [11:0]  u0_col_out_707;
wire  [11:0]  u0_col_out_708;
wire  [11:0]  u0_col_out_709;
wire  [11:0]  u0_col_out_710;
wire  [11:0]  u0_col_out_711;
wire  [11:0]  u0_col_out_712;
wire  [11:0]  u0_col_out_713;
wire  [11:0]  u0_col_out_714;
wire  [11:0]  u0_col_out_715;
wire  [11:0]  u0_col_out_716;
wire  [11:0]  u0_col_out_717;
wire  [11:0]  u0_col_out_718;
wire  [11:0]  u0_col_out_719;
wire  [11:0]  u0_col_out_720;
wire  [11:0]  u0_col_out_721;
wire  [11:0]  u0_col_out_722;
wire  [11:0]  u0_col_out_723;
wire  [11:0]  u0_col_out_724;
wire  [11:0]  u0_col_out_725;
wire  [11:0]  u0_col_out_726;
wire  [11:0]  u0_col_out_727;
wire  [11:0]  u0_col_out_728;
wire  [11:0]  u0_col_out_729;
wire  [11:0]  u0_col_out_730;
wire  [11:0]  u0_col_out_731;
wire  [11:0]  u0_col_out_732;
wire  [11:0]  u0_col_out_733;
wire  [11:0]  u0_col_out_734;
wire  [11:0]  u0_col_out_735;
wire  [11:0]  u0_col_out_736;
wire  [11:0]  u0_col_out_737;
wire  [11:0]  u0_col_out_738;
wire  [11:0]  u0_col_out_739;
wire  [11:0]  u0_col_out_740;
wire  [11:0]  u0_col_out_741;
wire  [11:0]  u0_col_out_742;
wire  [11:0]  u0_col_out_743;
wire  [11:0]  u0_col_out_744;
wire  [11:0]  u0_col_out_745;
wire  [11:0]  u0_col_out_746;
wire  [11:0]  u0_col_out_747;
wire  [11:0]  u0_col_out_748;
wire  [11:0]  u0_col_out_749;
wire  [11:0]  u0_col_out_750;
wire  [11:0]  u0_col_out_751;
wire  [11:0]  u0_col_out_752;
wire  [11:0]  u0_col_out_753;
wire  [11:0]  u0_col_out_754;
wire  [11:0]  u0_col_out_755;
wire  [11:0]  u0_col_out_756;
wire  [11:0]  u0_col_out_757;
wire  [11:0]  u0_col_out_758;
wire  [11:0]  u0_col_out_759;
wire  [11:0]  u0_col_out_760;
wire  [11:0]  u0_col_out_761;
wire  [11:0]  u0_col_out_762;
wire  [11:0]  u0_col_out_763;
wire  [11:0]  u0_col_out_764;
wire  [11:0]  u0_col_out_765;
wire  [11:0]  u0_col_out_766;
wire  [11:0]  u0_col_out_767;
wire  [11:0]  u0_col_out_768;
wire  [11:0]  u0_col_out_769;
wire  [11:0]  u0_col_out_770;
wire  [11:0]  u0_col_out_771;
wire  [11:0]  u0_col_out_772;
wire  [11:0]  u0_col_out_773;
wire  [11:0]  u0_col_out_774;
wire  [11:0]  u0_col_out_775;
wire  [11:0]  u0_col_out_776;
wire  [11:0]  u0_col_out_777;
wire  [11:0]  u0_col_out_778;
wire  [11:0]  u0_col_out_779;
wire  [11:0]  u0_col_out_780;
wire  [11:0]  u0_col_out_781;
wire  [11:0]  u0_col_out_782;
wire  [11:0]  u0_col_out_783;
wire  [11:0]  u0_col_out_784;
wire  [11:0]  u0_col_out_785;
wire  [11:0]  u0_col_out_786;
wire  [11:0]  u0_col_out_787;
wire  [11:0]  u0_col_out_788;
wire  [11:0]  u0_col_out_789;
wire  [11:0]  u0_col_out_790;
wire  [11:0]  u0_col_out_791;
wire  [11:0]  u0_col_out_792;
wire  [11:0]  u0_col_out_793;
wire  [11:0]  u0_col_out_794;
wire  [11:0]  u0_col_out_795;
wire  [11:0]  u0_col_out_796;
wire  [11:0]  u0_col_out_797;
wire  [11:0]  u0_col_out_798;
wire  [11:0]  u0_col_out_799;
wire  [11:0]  u0_col_out_800;
wire  [11:0]  u0_col_out_801;
wire  [11:0]  u0_col_out_802;
wire  [11:0]  u0_col_out_803;
wire  [11:0]  u0_col_out_804;
wire  [11:0]  u0_col_out_805;
wire  [11:0]  u0_col_out_806;
wire  [11:0]  u0_col_out_807;
wire  [11:0]  u0_col_out_808;
wire  [11:0]  u0_col_out_809;
wire  [11:0]  u0_col_out_810;
wire  [11:0]  u0_col_out_811;
wire  [11:0]  u0_col_out_812;
wire  [11:0]  u0_col_out_813;
wire  [11:0]  u0_col_out_814;
wire  [11:0]  u0_col_out_815;
wire  [11:0]  u0_col_out_816;
wire  [11:0]  u0_col_out_817;
wire  [11:0]  u0_col_out_818;
wire  [11:0]  u0_col_out_819;
wire  [11:0]  u0_col_out_820;
wire  [11:0]  u0_col_out_821;
wire  [11:0]  u0_col_out_822;
wire  [11:0]  u0_col_out_823;
wire  [11:0]  u0_col_out_824;
wire  [11:0]  u0_col_out_825;
wire  [11:0]  u0_col_out_826;
wire  [11:0]  u0_col_out_827;
wire  [11:0]  u0_col_out_828;
wire  [11:0]  u0_col_out_829;
wire  [11:0]  u0_col_out_830;
wire  [11:0]  u0_col_out_831;
wire  [11:0]  u0_col_out_832;
wire  [11:0]  u0_col_out_833;
wire  [11:0]  u0_col_out_834;
wire  [11:0]  u0_col_out_835;
wire  [11:0]  u0_col_out_836;
wire  [11:0]  u0_col_out_837;
wire  [11:0]  u0_col_out_838;
wire  [11:0]  u0_col_out_839;
wire  [11:0]  u0_col_out_840;
wire  [11:0]  u0_col_out_841;
wire  [11:0]  u0_col_out_842;
wire  [11:0]  u0_col_out_843;
wire  [11:0]  u0_col_out_844;
wire  [11:0]  u0_col_out_845;
wire  [11:0]  u0_col_out_846;
wire  [11:0]  u0_col_out_847;
wire  [11:0]  u0_col_out_848;
wire  [11:0]  u0_col_out_849;
wire  [11:0]  u0_col_out_850;
wire  [11:0]  u0_col_out_851;
wire  [11:0]  u0_col_out_852;
wire  [11:0]  u0_col_out_853;
wire  [11:0]  u0_col_out_854;
wire  [11:0]  u0_col_out_855;
wire  [11:0]  u0_col_out_856;
wire  [11:0]  u0_col_out_857;
wire  [11:0]  u0_col_out_858;
wire  [11:0]  u0_col_out_859;
wire  [11:0]  u0_col_out_860;
wire  [11:0]  u0_col_out_861;
wire  [11:0]  u0_col_out_862;
wire  [11:0]  u0_col_out_863;
wire  [11:0]  u0_col_out_864;
wire  [11:0]  u0_col_out_865;
wire  [11:0]  u0_col_out_866;
wire  [11:0]  u0_col_out_867;
wire  [11:0]  u0_col_out_868;
wire  [11:0]  u0_col_out_869;
wire  [11:0]  u0_col_out_870;
wire  [11:0]  u0_col_out_871;
wire  [11:0]  u0_col_out_872;
wire  [11:0]  u0_col_out_873;
wire  [11:0]  u0_col_out_874;
wire  [11:0]  u0_col_out_875;
wire  [11:0]  u0_col_out_876;
wire  [11:0]  u0_col_out_877;
wire  [11:0]  u0_col_out_878;
wire  [11:0]  u0_col_out_879;
wire  [11:0]  u0_col_out_880;
wire  [11:0]  u0_col_out_881;
wire  [11:0]  u0_col_out_882;
wire  [11:0]  u0_col_out_883;
wire  [11:0]  u0_col_out_884;
wire  [11:0]  u0_col_out_885;
wire  [11:0]  u0_col_out_886;
wire  [11:0]  u0_col_out_887;
wire  [11:0]  u0_col_out_888;
wire  [11:0]  u0_col_out_889;
wire  [11:0]  u0_col_out_890;
wire  [11:0]  u0_col_out_891;
wire  [11:0]  u0_col_out_892;
wire  [11:0]  u0_col_out_893;
wire  [11:0]  u0_col_out_894;
wire  [11:0]  u0_col_out_895;
wire  [11:0]  u0_col_out_896;
wire  [11:0]  u0_col_out_897;
wire  [11:0]  u0_col_out_898;
wire  [11:0]  u0_col_out_899;
wire  [11:0]  u0_col_out_900;
wire  [11:0]  u0_col_out_901;
wire  [11:0]  u0_col_out_902;
wire  [11:0]  u0_col_out_903;
wire  [11:0]  u0_col_out_904;
wire  [11:0]  u0_col_out_905;
wire  [11:0]  u0_col_out_906;
wire  [11:0]  u0_col_out_907;
wire  [11:0]  u0_col_out_908;
wire  [11:0]  u0_col_out_909;
wire  [11:0]  u0_col_out_910;
wire  [11:0]  u0_col_out_911;
wire  [11:0]  u0_col_out_912;
wire  [11:0]  u0_col_out_913;
wire  [11:0]  u0_col_out_914;
wire  [11:0]  u0_col_out_915;
wire  [11:0]  u0_col_out_916;
wire  [11:0]  u0_col_out_917;
wire  [11:0]  u0_col_out_918;
wire  [11:0]  u0_col_out_919;
wire  [11:0]  u0_col_out_920;
wire  [11:0]  u0_col_out_921;
wire  [11:0]  u0_col_out_922;
wire  [11:0]  u0_col_out_923;
wire  [11:0]  u0_col_out_924;
wire  [11:0]  u0_col_out_925;
wire  [11:0]  u0_col_out_926;
wire  [11:0]  u0_col_out_927;
wire  [11:0]  u0_col_out_928;
wire  [11:0]  u0_col_out_929;
wire  [11:0]  u0_col_out_930;
wire  [11:0]  u0_col_out_931;
wire  [11:0]  u0_col_out_932;
wire  [11:0]  u0_col_out_933;
wire  [11:0]  u0_col_out_934;
wire  [11:0]  u0_col_out_935;
wire  [11:0]  u0_col_out_936;
wire  [11:0]  u0_col_out_937;
wire  [11:0]  u0_col_out_938;
wire  [11:0]  u0_col_out_939;
wire  [11:0]  u0_col_out_940;
wire  [11:0]  u0_col_out_941;
wire  [11:0]  u0_col_out_942;
wire  [11:0]  u0_col_out_943;
wire  [11:0]  u0_col_out_944;
wire  [11:0]  u0_col_out_945;
wire  [11:0]  u0_col_out_946;
wire  [11:0]  u0_col_out_947;
wire  [11:0]  u0_col_out_948;
wire  [11:0]  u0_col_out_949;
wire  [11:0]  u0_col_out_950;
wire  [11:0]  u0_col_out_951;
wire  [11:0]  u0_col_out_952;
wire  [11:0]  u0_col_out_953;
wire  [11:0]  u0_col_out_954;
wire  [11:0]  u0_col_out_955;
wire  [11:0]  u0_col_out_956;
wire  [11:0]  u0_col_out_957;
wire  [11:0]  u0_col_out_958;
wire  [11:0]  u0_col_out_959;
wire  [11:0]  u0_col_out_960;
wire  [11:0]  u0_col_out_961;
wire  [11:0]  u0_col_out_962;
wire  [11:0]  u0_col_out_963;
wire  [11:0]  u0_col_out_964;
wire  [11:0]  u0_col_out_965;
wire  [11:0]  u0_col_out_966;
wire  [11:0]  u0_col_out_967;
wire  [11:0]  u0_col_out_968;
wire  [11:0]  u0_col_out_969;
wire  [11:0]  u0_col_out_970;
wire  [11:0]  u0_col_out_971;
wire  [11:0]  u0_col_out_972;
wire  [11:0]  u0_col_out_973;
wire  [11:0]  u0_col_out_974;
wire  [11:0]  u0_col_out_975;
wire  [11:0]  u0_col_out_976;
wire  [11:0]  u0_col_out_977;
wire  [11:0]  u0_col_out_978;
wire  [11:0]  u0_col_out_979;
wire  [11:0]  u0_col_out_980;
wire  [11:0]  u0_col_out_981;
wire  [11:0]  u0_col_out_982;
wire  [11:0]  u0_col_out_983;
wire  [11:0]  u0_col_out_984;
wire  [11:0]  u0_col_out_985;
wire  [11:0]  u0_col_out_986;
wire  [11:0]  u0_col_out_987;
wire  [11:0]  u0_col_out_988;
wire  [11:0]  u0_col_out_989;
wire  [11:0]  u0_col_out_990;
wire  [11:0]  u0_col_out_991;
wire  [11:0]  u0_col_out_992;
wire  [11:0]  u0_col_out_993;
wire  [11:0]  u0_col_out_994;
wire  [11:0]  u0_col_out_995;
wire  [11:0]  u0_col_out_996;
wire  [11:0]  u0_col_out_997;
wire  [11:0]  u0_col_out_998;
wire  [11:0]  u0_col_out_999;
wire  [11:0]  u0_col_out_1000;
wire  [11:0]  u0_col_out_1001;
wire  [11:0]  u0_col_out_1002;
wire  [11:0]  u0_col_out_1003;
wire  [11:0]  u0_col_out_1004;
wire  [11:0]  u0_col_out_1005;
wire  [11:0]  u0_col_out_1006;
wire  [11:0]  u0_col_out_1007;
wire  [11:0]  u0_col_out_1008;
wire  [11:0]  u0_col_out_1009;
wire  [11:0]  u0_col_out_1010;
wire  [11:0]  u0_col_out_1011;
wire  [11:0]  u0_col_out_1012;
wire  [11:0]  u0_col_out_1013;
wire  [11:0]  u0_col_out_1014;
wire  [11:0]  u0_col_out_1015;
wire  [11:0]  u0_col_out_1016;
wire  [11:0]  u0_col_out_1017;
wire  [11:0]  u0_col_out_1018;
wire  [11:0]  u0_col_out_1019;
wire  [11:0]  u0_col_out_1020;
wire  [11:0]  u0_col_out_1021;
wire  [11:0]  u0_col_out_1022;
wire  [11:0]  u0_col_out_1023;
wire  [11:0]  u0_col_out_1024;
wire  [11:0]  u0_col_out_1025;
wire  [11:0]  u0_col_out_1026;
wire  [11:0]  u0_col_out_1027;
wire  [11:0]  u0_col_out_1028;
wire  [11:0]  u0_col_out_1029;
wire  [11:0]  u0_col_out_1030;
wire  [11:0]  u0_col_out_1031;
wire  [11:0]  u0_col_out_1032;
wire  [11:0]  u0_col_out_1033;

compressor_array_16_12_1033  u0_compressor_array_16_12_1033 (
    .col_in_0                ( col_in_0       ),
    .col_in_1                ( col_in_1       ),
    .col_in_2                ( col_in_2       ),
    .col_in_3                ( col_in_3       ),
    .col_in_4                ( col_in_4       ),
    .col_in_5                ( col_in_5       ),
    .col_in_6                ( col_in_6       ),
    .col_in_7                ( col_in_7       ),
    .col_in_8                ( col_in_8       ),
    .col_in_9                ( col_in_9       ),
    .col_in_10               ( col_in_10      ),
    .col_in_11               ( col_in_11      ),
    .col_in_12               ( col_in_12      ),
    .col_in_13               ( col_in_13      ),
    .col_in_14               ( col_in_14      ),
    .col_in_15               ( col_in_15      ),
    .col_in_16               ( col_in_16      ),
    .col_in_17               ( col_in_17      ),
    .col_in_18               ( col_in_18      ),
    .col_in_19               ( col_in_19      ),
    .col_in_20               ( col_in_20      ),
    .col_in_21               ( col_in_21      ),
    .col_in_22               ( col_in_22      ),
    .col_in_23               ( col_in_23      ),
    .col_in_24               ( col_in_24      ),
    .col_in_25               ( col_in_25      ),
    .col_in_26               ( col_in_26      ),
    .col_in_27               ( col_in_27      ),
    .col_in_28               ( col_in_28      ),
    .col_in_29               ( col_in_29      ),
    .col_in_30               ( col_in_30      ),
    .col_in_31               ( col_in_31      ),
    .col_in_32               ( col_in_32      ),
    .col_in_33               ( col_in_33      ),
    .col_in_34               ( col_in_34      ),
    .col_in_35               ( col_in_35      ),
    .col_in_36               ( col_in_36      ),
    .col_in_37               ( col_in_37      ),
    .col_in_38               ( col_in_38      ),
    .col_in_39               ( col_in_39      ),
    .col_in_40               ( col_in_40      ),
    .col_in_41               ( col_in_41      ),
    .col_in_42               ( col_in_42      ),
    .col_in_43               ( col_in_43      ),
    .col_in_44               ( col_in_44      ),
    .col_in_45               ( col_in_45      ),
    .col_in_46               ( col_in_46      ),
    .col_in_47               ( col_in_47      ),
    .col_in_48               ( col_in_48      ),
    .col_in_49               ( col_in_49      ),
    .col_in_50               ( col_in_50      ),
    .col_in_51               ( col_in_51      ),
    .col_in_52               ( col_in_52      ),
    .col_in_53               ( col_in_53      ),
    .col_in_54               ( col_in_54      ),
    .col_in_55               ( col_in_55      ),
    .col_in_56               ( col_in_56      ),
    .col_in_57               ( col_in_57      ),
    .col_in_58               ( col_in_58      ),
    .col_in_59               ( col_in_59      ),
    .col_in_60               ( col_in_60      ),
    .col_in_61               ( col_in_61      ),
    .col_in_62               ( col_in_62      ),
    .col_in_63               ( col_in_63      ),
    .col_in_64               ( col_in_64      ),
    .col_in_65               ( col_in_65      ),
    .col_in_66               ( col_in_66      ),
    .col_in_67               ( col_in_67      ),
    .col_in_68               ( col_in_68      ),
    .col_in_69               ( col_in_69      ),
    .col_in_70               ( col_in_70      ),
    .col_in_71               ( col_in_71      ),
    .col_in_72               ( col_in_72      ),
    .col_in_73               ( col_in_73      ),
    .col_in_74               ( col_in_74      ),
    .col_in_75               ( col_in_75      ),
    .col_in_76               ( col_in_76      ),
    .col_in_77               ( col_in_77      ),
    .col_in_78               ( col_in_78      ),
    .col_in_79               ( col_in_79      ),
    .col_in_80               ( col_in_80      ),
    .col_in_81               ( col_in_81      ),
    .col_in_82               ( col_in_82      ),
    .col_in_83               ( col_in_83      ),
    .col_in_84               ( col_in_84      ),
    .col_in_85               ( col_in_85      ),
    .col_in_86               ( col_in_86      ),
    .col_in_87               ( col_in_87      ),
    .col_in_88               ( col_in_88      ),
    .col_in_89               ( col_in_89      ),
    .col_in_90               ( col_in_90      ),
    .col_in_91               ( col_in_91      ),
    .col_in_92               ( col_in_92      ),
    .col_in_93               ( col_in_93      ),
    .col_in_94               ( col_in_94      ),
    .col_in_95               ( col_in_95      ),
    .col_in_96               ( col_in_96      ),
    .col_in_97               ( col_in_97      ),
    .col_in_98               ( col_in_98      ),
    .col_in_99               ( col_in_99      ),
    .col_in_100              ( col_in_100     ),
    .col_in_101              ( col_in_101     ),
    .col_in_102              ( col_in_102     ),
    .col_in_103              ( col_in_103     ),
    .col_in_104              ( col_in_104     ),
    .col_in_105              ( col_in_105     ),
    .col_in_106              ( col_in_106     ),
    .col_in_107              ( col_in_107     ),
    .col_in_108              ( col_in_108     ),
    .col_in_109              ( col_in_109     ),
    .col_in_110              ( col_in_110     ),
    .col_in_111              ( col_in_111     ),
    .col_in_112              ( col_in_112     ),
    .col_in_113              ( col_in_113     ),
    .col_in_114              ( col_in_114     ),
    .col_in_115              ( col_in_115     ),
    .col_in_116              ( col_in_116     ),
    .col_in_117              ( col_in_117     ),
    .col_in_118              ( col_in_118     ),
    .col_in_119              ( col_in_119     ),
    .col_in_120              ( col_in_120     ),
    .col_in_121              ( col_in_121     ),
    .col_in_122              ( col_in_122     ),
    .col_in_123              ( col_in_123     ),
    .col_in_124              ( col_in_124     ),
    .col_in_125              ( col_in_125     ),
    .col_in_126              ( col_in_126     ),
    .col_in_127              ( col_in_127     ),
    .col_in_128              ( col_in_128     ),
    .col_in_129              ( col_in_129     ),
    .col_in_130              ( col_in_130     ),
    .col_in_131              ( col_in_131     ),
    .col_in_132              ( col_in_132     ),
    .col_in_133              ( col_in_133     ),
    .col_in_134              ( col_in_134     ),
    .col_in_135              ( col_in_135     ),
    .col_in_136              ( col_in_136     ),
    .col_in_137              ( col_in_137     ),
    .col_in_138              ( col_in_138     ),
    .col_in_139              ( col_in_139     ),
    .col_in_140              ( col_in_140     ),
    .col_in_141              ( col_in_141     ),
    .col_in_142              ( col_in_142     ),
    .col_in_143              ( col_in_143     ),
    .col_in_144              ( col_in_144     ),
    .col_in_145              ( col_in_145     ),
    .col_in_146              ( col_in_146     ),
    .col_in_147              ( col_in_147     ),
    .col_in_148              ( col_in_148     ),
    .col_in_149              ( col_in_149     ),
    .col_in_150              ( col_in_150     ),
    .col_in_151              ( col_in_151     ),
    .col_in_152              ( col_in_152     ),
    .col_in_153              ( col_in_153     ),
    .col_in_154              ( col_in_154     ),
    .col_in_155              ( col_in_155     ),
    .col_in_156              ( col_in_156     ),
    .col_in_157              ( col_in_157     ),
    .col_in_158              ( col_in_158     ),
    .col_in_159              ( col_in_159     ),
    .col_in_160              ( col_in_160     ),
    .col_in_161              ( col_in_161     ),
    .col_in_162              ( col_in_162     ),
    .col_in_163              ( col_in_163     ),
    .col_in_164              ( col_in_164     ),
    .col_in_165              ( col_in_165     ),
    .col_in_166              ( col_in_166     ),
    .col_in_167              ( col_in_167     ),
    .col_in_168              ( col_in_168     ),
    .col_in_169              ( col_in_169     ),
    .col_in_170              ( col_in_170     ),
    .col_in_171              ( col_in_171     ),
    .col_in_172              ( col_in_172     ),
    .col_in_173              ( col_in_173     ),
    .col_in_174              ( col_in_174     ),
    .col_in_175              ( col_in_175     ),
    .col_in_176              ( col_in_176     ),
    .col_in_177              ( col_in_177     ),
    .col_in_178              ( col_in_178     ),
    .col_in_179              ( col_in_179     ),
    .col_in_180              ( col_in_180     ),
    .col_in_181              ( col_in_181     ),
    .col_in_182              ( col_in_182     ),
    .col_in_183              ( col_in_183     ),
    .col_in_184              ( col_in_184     ),
    .col_in_185              ( col_in_185     ),
    .col_in_186              ( col_in_186     ),
    .col_in_187              ( col_in_187     ),
    .col_in_188              ( col_in_188     ),
    .col_in_189              ( col_in_189     ),
    .col_in_190              ( col_in_190     ),
    .col_in_191              ( col_in_191     ),
    .col_in_192              ( col_in_192     ),
    .col_in_193              ( col_in_193     ),
    .col_in_194              ( col_in_194     ),
    .col_in_195              ( col_in_195     ),
    .col_in_196              ( col_in_196     ),
    .col_in_197              ( col_in_197     ),
    .col_in_198              ( col_in_198     ),
    .col_in_199              ( col_in_199     ),
    .col_in_200              ( col_in_200     ),
    .col_in_201              ( col_in_201     ),
    .col_in_202              ( col_in_202     ),
    .col_in_203              ( col_in_203     ),
    .col_in_204              ( col_in_204     ),
    .col_in_205              ( col_in_205     ),
    .col_in_206              ( col_in_206     ),
    .col_in_207              ( col_in_207     ),
    .col_in_208              ( col_in_208     ),
    .col_in_209              ( col_in_209     ),
    .col_in_210              ( col_in_210     ),
    .col_in_211              ( col_in_211     ),
    .col_in_212              ( col_in_212     ),
    .col_in_213              ( col_in_213     ),
    .col_in_214              ( col_in_214     ),
    .col_in_215              ( col_in_215     ),
    .col_in_216              ( col_in_216     ),
    .col_in_217              ( col_in_217     ),
    .col_in_218              ( col_in_218     ),
    .col_in_219              ( col_in_219     ),
    .col_in_220              ( col_in_220     ),
    .col_in_221              ( col_in_221     ),
    .col_in_222              ( col_in_222     ),
    .col_in_223              ( col_in_223     ),
    .col_in_224              ( col_in_224     ),
    .col_in_225              ( col_in_225     ),
    .col_in_226              ( col_in_226     ),
    .col_in_227              ( col_in_227     ),
    .col_in_228              ( col_in_228     ),
    .col_in_229              ( col_in_229     ),
    .col_in_230              ( col_in_230     ),
    .col_in_231              ( col_in_231     ),
    .col_in_232              ( col_in_232     ),
    .col_in_233              ( col_in_233     ),
    .col_in_234              ( col_in_234     ),
    .col_in_235              ( col_in_235     ),
    .col_in_236              ( col_in_236     ),
    .col_in_237              ( col_in_237     ),
    .col_in_238              ( col_in_238     ),
    .col_in_239              ( col_in_239     ),
    .col_in_240              ( col_in_240     ),
    .col_in_241              ( col_in_241     ),
    .col_in_242              ( col_in_242     ),
    .col_in_243              ( col_in_243     ),
    .col_in_244              ( col_in_244     ),
    .col_in_245              ( col_in_245     ),
    .col_in_246              ( col_in_246     ),
    .col_in_247              ( col_in_247     ),
    .col_in_248              ( col_in_248     ),
    .col_in_249              ( col_in_249     ),
    .col_in_250              ( col_in_250     ),
    .col_in_251              ( col_in_251     ),
    .col_in_252              ( col_in_252     ),
    .col_in_253              ( col_in_253     ),
    .col_in_254              ( col_in_254     ),
    .col_in_255              ( col_in_255     ),
    .col_in_256              ( col_in_256     ),
    .col_in_257              ( col_in_257     ),
    .col_in_258              ( col_in_258     ),
    .col_in_259              ( col_in_259     ),
    .col_in_260              ( col_in_260     ),
    .col_in_261              ( col_in_261     ),
    .col_in_262              ( col_in_262     ),
    .col_in_263              ( col_in_263     ),
    .col_in_264              ( col_in_264     ),
    .col_in_265              ( col_in_265     ),
    .col_in_266              ( col_in_266     ),
    .col_in_267              ( col_in_267     ),
    .col_in_268              ( col_in_268     ),
    .col_in_269              ( col_in_269     ),
    .col_in_270              ( col_in_270     ),
    .col_in_271              ( col_in_271     ),
    .col_in_272              ( col_in_272     ),
    .col_in_273              ( col_in_273     ),
    .col_in_274              ( col_in_274     ),
    .col_in_275              ( col_in_275     ),
    .col_in_276              ( col_in_276     ),
    .col_in_277              ( col_in_277     ),
    .col_in_278              ( col_in_278     ),
    .col_in_279              ( col_in_279     ),
    .col_in_280              ( col_in_280     ),
    .col_in_281              ( col_in_281     ),
    .col_in_282              ( col_in_282     ),
    .col_in_283              ( col_in_283     ),
    .col_in_284              ( col_in_284     ),
    .col_in_285              ( col_in_285     ),
    .col_in_286              ( col_in_286     ),
    .col_in_287              ( col_in_287     ),
    .col_in_288              ( col_in_288     ),
    .col_in_289              ( col_in_289     ),
    .col_in_290              ( col_in_290     ),
    .col_in_291              ( col_in_291     ),
    .col_in_292              ( col_in_292     ),
    .col_in_293              ( col_in_293     ),
    .col_in_294              ( col_in_294     ),
    .col_in_295              ( col_in_295     ),
    .col_in_296              ( col_in_296     ),
    .col_in_297              ( col_in_297     ),
    .col_in_298              ( col_in_298     ),
    .col_in_299              ( col_in_299     ),
    .col_in_300              ( col_in_300     ),
    .col_in_301              ( col_in_301     ),
    .col_in_302              ( col_in_302     ),
    .col_in_303              ( col_in_303     ),
    .col_in_304              ( col_in_304     ),
    .col_in_305              ( col_in_305     ),
    .col_in_306              ( col_in_306     ),
    .col_in_307              ( col_in_307     ),
    .col_in_308              ( col_in_308     ),
    .col_in_309              ( col_in_309     ),
    .col_in_310              ( col_in_310     ),
    .col_in_311              ( col_in_311     ),
    .col_in_312              ( col_in_312     ),
    .col_in_313              ( col_in_313     ),
    .col_in_314              ( col_in_314     ),
    .col_in_315              ( col_in_315     ),
    .col_in_316              ( col_in_316     ),
    .col_in_317              ( col_in_317     ),
    .col_in_318              ( col_in_318     ),
    .col_in_319              ( col_in_319     ),
    .col_in_320              ( col_in_320     ),
    .col_in_321              ( col_in_321     ),
    .col_in_322              ( col_in_322     ),
    .col_in_323              ( col_in_323     ),
    .col_in_324              ( col_in_324     ),
    .col_in_325              ( col_in_325     ),
    .col_in_326              ( col_in_326     ),
    .col_in_327              ( col_in_327     ),
    .col_in_328              ( col_in_328     ),
    .col_in_329              ( col_in_329     ),
    .col_in_330              ( col_in_330     ),
    .col_in_331              ( col_in_331     ),
    .col_in_332              ( col_in_332     ),
    .col_in_333              ( col_in_333     ),
    .col_in_334              ( col_in_334     ),
    .col_in_335              ( col_in_335     ),
    .col_in_336              ( col_in_336     ),
    .col_in_337              ( col_in_337     ),
    .col_in_338              ( col_in_338     ),
    .col_in_339              ( col_in_339     ),
    .col_in_340              ( col_in_340     ),
    .col_in_341              ( col_in_341     ),
    .col_in_342              ( col_in_342     ),
    .col_in_343              ( col_in_343     ),
    .col_in_344              ( col_in_344     ),
    .col_in_345              ( col_in_345     ),
    .col_in_346              ( col_in_346     ),
    .col_in_347              ( col_in_347     ),
    .col_in_348              ( col_in_348     ),
    .col_in_349              ( col_in_349     ),
    .col_in_350              ( col_in_350     ),
    .col_in_351              ( col_in_351     ),
    .col_in_352              ( col_in_352     ),
    .col_in_353              ( col_in_353     ),
    .col_in_354              ( col_in_354     ),
    .col_in_355              ( col_in_355     ),
    .col_in_356              ( col_in_356     ),
    .col_in_357              ( col_in_357     ),
    .col_in_358              ( col_in_358     ),
    .col_in_359              ( col_in_359     ),
    .col_in_360              ( col_in_360     ),
    .col_in_361              ( col_in_361     ),
    .col_in_362              ( col_in_362     ),
    .col_in_363              ( col_in_363     ),
    .col_in_364              ( col_in_364     ),
    .col_in_365              ( col_in_365     ),
    .col_in_366              ( col_in_366     ),
    .col_in_367              ( col_in_367     ),
    .col_in_368              ( col_in_368     ),
    .col_in_369              ( col_in_369     ),
    .col_in_370              ( col_in_370     ),
    .col_in_371              ( col_in_371     ),
    .col_in_372              ( col_in_372     ),
    .col_in_373              ( col_in_373     ),
    .col_in_374              ( col_in_374     ),
    .col_in_375              ( col_in_375     ),
    .col_in_376              ( col_in_376     ),
    .col_in_377              ( col_in_377     ),
    .col_in_378              ( col_in_378     ),
    .col_in_379              ( col_in_379     ),
    .col_in_380              ( col_in_380     ),
    .col_in_381              ( col_in_381     ),
    .col_in_382              ( col_in_382     ),
    .col_in_383              ( col_in_383     ),
    .col_in_384              ( col_in_384     ),
    .col_in_385              ( col_in_385     ),
    .col_in_386              ( col_in_386     ),
    .col_in_387              ( col_in_387     ),
    .col_in_388              ( col_in_388     ),
    .col_in_389              ( col_in_389     ),
    .col_in_390              ( col_in_390     ),
    .col_in_391              ( col_in_391     ),
    .col_in_392              ( col_in_392     ),
    .col_in_393              ( col_in_393     ),
    .col_in_394              ( col_in_394     ),
    .col_in_395              ( col_in_395     ),
    .col_in_396              ( col_in_396     ),
    .col_in_397              ( col_in_397     ),
    .col_in_398              ( col_in_398     ),
    .col_in_399              ( col_in_399     ),
    .col_in_400              ( col_in_400     ),
    .col_in_401              ( col_in_401     ),
    .col_in_402              ( col_in_402     ),
    .col_in_403              ( col_in_403     ),
    .col_in_404              ( col_in_404     ),
    .col_in_405              ( col_in_405     ),
    .col_in_406              ( col_in_406     ),
    .col_in_407              ( col_in_407     ),
    .col_in_408              ( col_in_408     ),
    .col_in_409              ( col_in_409     ),
    .col_in_410              ( col_in_410     ),
    .col_in_411              ( col_in_411     ),
    .col_in_412              ( col_in_412     ),
    .col_in_413              ( col_in_413     ),
    .col_in_414              ( col_in_414     ),
    .col_in_415              ( col_in_415     ),
    .col_in_416              ( col_in_416     ),
    .col_in_417              ( col_in_417     ),
    .col_in_418              ( col_in_418     ),
    .col_in_419              ( col_in_419     ),
    .col_in_420              ( col_in_420     ),
    .col_in_421              ( col_in_421     ),
    .col_in_422              ( col_in_422     ),
    .col_in_423              ( col_in_423     ),
    .col_in_424              ( col_in_424     ),
    .col_in_425              ( col_in_425     ),
    .col_in_426              ( col_in_426     ),
    .col_in_427              ( col_in_427     ),
    .col_in_428              ( col_in_428     ),
    .col_in_429              ( col_in_429     ),
    .col_in_430              ( col_in_430     ),
    .col_in_431              ( col_in_431     ),
    .col_in_432              ( col_in_432     ),
    .col_in_433              ( col_in_433     ),
    .col_in_434              ( col_in_434     ),
    .col_in_435              ( col_in_435     ),
    .col_in_436              ( col_in_436     ),
    .col_in_437              ( col_in_437     ),
    .col_in_438              ( col_in_438     ),
    .col_in_439              ( col_in_439     ),
    .col_in_440              ( col_in_440     ),
    .col_in_441              ( col_in_441     ),
    .col_in_442              ( col_in_442     ),
    .col_in_443              ( col_in_443     ),
    .col_in_444              ( col_in_444     ),
    .col_in_445              ( col_in_445     ),
    .col_in_446              ( col_in_446     ),
    .col_in_447              ( col_in_447     ),
    .col_in_448              ( col_in_448     ),
    .col_in_449              ( col_in_449     ),
    .col_in_450              ( col_in_450     ),
    .col_in_451              ( col_in_451     ),
    .col_in_452              ( col_in_452     ),
    .col_in_453              ( col_in_453     ),
    .col_in_454              ( col_in_454     ),
    .col_in_455              ( col_in_455     ),
    .col_in_456              ( col_in_456     ),
    .col_in_457              ( col_in_457     ),
    .col_in_458              ( col_in_458     ),
    .col_in_459              ( col_in_459     ),
    .col_in_460              ( col_in_460     ),
    .col_in_461              ( col_in_461     ),
    .col_in_462              ( col_in_462     ),
    .col_in_463              ( col_in_463     ),
    .col_in_464              ( col_in_464     ),
    .col_in_465              ( col_in_465     ),
    .col_in_466              ( col_in_466     ),
    .col_in_467              ( col_in_467     ),
    .col_in_468              ( col_in_468     ),
    .col_in_469              ( col_in_469     ),
    .col_in_470              ( col_in_470     ),
    .col_in_471              ( col_in_471     ),
    .col_in_472              ( col_in_472     ),
    .col_in_473              ( col_in_473     ),
    .col_in_474              ( col_in_474     ),
    .col_in_475              ( col_in_475     ),
    .col_in_476              ( col_in_476     ),
    .col_in_477              ( col_in_477     ),
    .col_in_478              ( col_in_478     ),
    .col_in_479              ( col_in_479     ),
    .col_in_480              ( col_in_480     ),
    .col_in_481              ( col_in_481     ),
    .col_in_482              ( col_in_482     ),
    .col_in_483              ( col_in_483     ),
    .col_in_484              ( col_in_484     ),
    .col_in_485              ( col_in_485     ),
    .col_in_486              ( col_in_486     ),
    .col_in_487              ( col_in_487     ),
    .col_in_488              ( col_in_488     ),
    .col_in_489              ( col_in_489     ),
    .col_in_490              ( col_in_490     ),
    .col_in_491              ( col_in_491     ),
    .col_in_492              ( col_in_492     ),
    .col_in_493              ( col_in_493     ),
    .col_in_494              ( col_in_494     ),
    .col_in_495              ( col_in_495     ),
    .col_in_496              ( col_in_496     ),
    .col_in_497              ( col_in_497     ),
    .col_in_498              ( col_in_498     ),
    .col_in_499              ( col_in_499     ),
    .col_in_500              ( col_in_500     ),
    .col_in_501              ( col_in_501     ),
    .col_in_502              ( col_in_502     ),
    .col_in_503              ( col_in_503     ),
    .col_in_504              ( col_in_504     ),
    .col_in_505              ( col_in_505     ),
    .col_in_506              ( col_in_506     ),
    .col_in_507              ( col_in_507     ),
    .col_in_508              ( col_in_508     ),
    .col_in_509              ( col_in_509     ),
    .col_in_510              ( col_in_510     ),
    .col_in_511              ( col_in_511     ),
    .col_in_512              ( col_in_512     ),
    .col_in_513              ( col_in_513     ),
    .col_in_514              ( col_in_514     ),
    .col_in_515              ( col_in_515     ),
    .col_in_516              ( col_in_516     ),
    .col_in_517              ( col_in_517     ),
    .col_in_518              ( col_in_518     ),
    .col_in_519              ( col_in_519     ),
    .col_in_520              ( col_in_520     ),
    .col_in_521              ( col_in_521     ),
    .col_in_522              ( col_in_522     ),
    .col_in_523              ( col_in_523     ),
    .col_in_524              ( col_in_524     ),
    .col_in_525              ( col_in_525     ),
    .col_in_526              ( col_in_526     ),
    .col_in_527              ( col_in_527     ),
    .col_in_528              ( col_in_528     ),
    .col_in_529              ( col_in_529     ),
    .col_in_530              ( col_in_530     ),
    .col_in_531              ( col_in_531     ),
    .col_in_532              ( col_in_532     ),
    .col_in_533              ( col_in_533     ),
    .col_in_534              ( col_in_534     ),
    .col_in_535              ( col_in_535     ),
    .col_in_536              ( col_in_536     ),
    .col_in_537              ( col_in_537     ),
    .col_in_538              ( col_in_538     ),
    .col_in_539              ( col_in_539     ),
    .col_in_540              ( col_in_540     ),
    .col_in_541              ( col_in_541     ),
    .col_in_542              ( col_in_542     ),
    .col_in_543              ( col_in_543     ),
    .col_in_544              ( col_in_544     ),
    .col_in_545              ( col_in_545     ),
    .col_in_546              ( col_in_546     ),
    .col_in_547              ( col_in_547     ),
    .col_in_548              ( col_in_548     ),
    .col_in_549              ( col_in_549     ),
    .col_in_550              ( col_in_550     ),
    .col_in_551              ( col_in_551     ),
    .col_in_552              ( col_in_552     ),
    .col_in_553              ( col_in_553     ),
    .col_in_554              ( col_in_554     ),
    .col_in_555              ( col_in_555     ),
    .col_in_556              ( col_in_556     ),
    .col_in_557              ( col_in_557     ),
    .col_in_558              ( col_in_558     ),
    .col_in_559              ( col_in_559     ),
    .col_in_560              ( col_in_560     ),
    .col_in_561              ( col_in_561     ),
    .col_in_562              ( col_in_562     ),
    .col_in_563              ( col_in_563     ),
    .col_in_564              ( col_in_564     ),
    .col_in_565              ( col_in_565     ),
    .col_in_566              ( col_in_566     ),
    .col_in_567              ( col_in_567     ),
    .col_in_568              ( col_in_568     ),
    .col_in_569              ( col_in_569     ),
    .col_in_570              ( col_in_570     ),
    .col_in_571              ( col_in_571     ),
    .col_in_572              ( col_in_572     ),
    .col_in_573              ( col_in_573     ),
    .col_in_574              ( col_in_574     ),
    .col_in_575              ( col_in_575     ),
    .col_in_576              ( col_in_576     ),
    .col_in_577              ( col_in_577     ),
    .col_in_578              ( col_in_578     ),
    .col_in_579              ( col_in_579     ),
    .col_in_580              ( col_in_580     ),
    .col_in_581              ( col_in_581     ),
    .col_in_582              ( col_in_582     ),
    .col_in_583              ( col_in_583     ),
    .col_in_584              ( col_in_584     ),
    .col_in_585              ( col_in_585     ),
    .col_in_586              ( col_in_586     ),
    .col_in_587              ( col_in_587     ),
    .col_in_588              ( col_in_588     ),
    .col_in_589              ( col_in_589     ),
    .col_in_590              ( col_in_590     ),
    .col_in_591              ( col_in_591     ),
    .col_in_592              ( col_in_592     ),
    .col_in_593              ( col_in_593     ),
    .col_in_594              ( col_in_594     ),
    .col_in_595              ( col_in_595     ),
    .col_in_596              ( col_in_596     ),
    .col_in_597              ( col_in_597     ),
    .col_in_598              ( col_in_598     ),
    .col_in_599              ( col_in_599     ),
    .col_in_600              ( col_in_600     ),
    .col_in_601              ( col_in_601     ),
    .col_in_602              ( col_in_602     ),
    .col_in_603              ( col_in_603     ),
    .col_in_604              ( col_in_604     ),
    .col_in_605              ( col_in_605     ),
    .col_in_606              ( col_in_606     ),
    .col_in_607              ( col_in_607     ),
    .col_in_608              ( col_in_608     ),
    .col_in_609              ( col_in_609     ),
    .col_in_610              ( col_in_610     ),
    .col_in_611              ( col_in_611     ),
    .col_in_612              ( col_in_612     ),
    .col_in_613              ( col_in_613     ),
    .col_in_614              ( col_in_614     ),
    .col_in_615              ( col_in_615     ),
    .col_in_616              ( col_in_616     ),
    .col_in_617              ( col_in_617     ),
    .col_in_618              ( col_in_618     ),
    .col_in_619              ( col_in_619     ),
    .col_in_620              ( col_in_620     ),
    .col_in_621              ( col_in_621     ),
    .col_in_622              ( col_in_622     ),
    .col_in_623              ( col_in_623     ),
    .col_in_624              ( col_in_624     ),
    .col_in_625              ( col_in_625     ),
    .col_in_626              ( col_in_626     ),
    .col_in_627              ( col_in_627     ),
    .col_in_628              ( col_in_628     ),
    .col_in_629              ( col_in_629     ),
    .col_in_630              ( col_in_630     ),
    .col_in_631              ( col_in_631     ),
    .col_in_632              ( col_in_632     ),
    .col_in_633              ( col_in_633     ),
    .col_in_634              ( col_in_634     ),
    .col_in_635              ( col_in_635     ),
    .col_in_636              ( col_in_636     ),
    .col_in_637              ( col_in_637     ),
    .col_in_638              ( col_in_638     ),
    .col_in_639              ( col_in_639     ),
    .col_in_640              ( col_in_640     ),
    .col_in_641              ( col_in_641     ),
    .col_in_642              ( col_in_642     ),
    .col_in_643              ( col_in_643     ),
    .col_in_644              ( col_in_644     ),
    .col_in_645              ( col_in_645     ),
    .col_in_646              ( col_in_646     ),
    .col_in_647              ( col_in_647     ),
    .col_in_648              ( col_in_648     ),
    .col_in_649              ( col_in_649     ),
    .col_in_650              ( col_in_650     ),
    .col_in_651              ( col_in_651     ),
    .col_in_652              ( col_in_652     ),
    .col_in_653              ( col_in_653     ),
    .col_in_654              ( col_in_654     ),
    .col_in_655              ( col_in_655     ),
    .col_in_656              ( col_in_656     ),
    .col_in_657              ( col_in_657     ),
    .col_in_658              ( col_in_658     ),
    .col_in_659              ( col_in_659     ),
    .col_in_660              ( col_in_660     ),
    .col_in_661              ( col_in_661     ),
    .col_in_662              ( col_in_662     ),
    .col_in_663              ( col_in_663     ),
    .col_in_664              ( col_in_664     ),
    .col_in_665              ( col_in_665     ),
    .col_in_666              ( col_in_666     ),
    .col_in_667              ( col_in_667     ),
    .col_in_668              ( col_in_668     ),
    .col_in_669              ( col_in_669     ),
    .col_in_670              ( col_in_670     ),
    .col_in_671              ( col_in_671     ),
    .col_in_672              ( col_in_672     ),
    .col_in_673              ( col_in_673     ),
    .col_in_674              ( col_in_674     ),
    .col_in_675              ( col_in_675     ),
    .col_in_676              ( col_in_676     ),
    .col_in_677              ( col_in_677     ),
    .col_in_678              ( col_in_678     ),
    .col_in_679              ( col_in_679     ),
    .col_in_680              ( col_in_680     ),
    .col_in_681              ( col_in_681     ),
    .col_in_682              ( col_in_682     ),
    .col_in_683              ( col_in_683     ),
    .col_in_684              ( col_in_684     ),
    .col_in_685              ( col_in_685     ),
    .col_in_686              ( col_in_686     ),
    .col_in_687              ( col_in_687     ),
    .col_in_688              ( col_in_688     ),
    .col_in_689              ( col_in_689     ),
    .col_in_690              ( col_in_690     ),
    .col_in_691              ( col_in_691     ),
    .col_in_692              ( col_in_692     ),
    .col_in_693              ( col_in_693     ),
    .col_in_694              ( col_in_694     ),
    .col_in_695              ( col_in_695     ),
    .col_in_696              ( col_in_696     ),
    .col_in_697              ( col_in_697     ),
    .col_in_698              ( col_in_698     ),
    .col_in_699              ( col_in_699     ),
    .col_in_700              ( col_in_700     ),
    .col_in_701              ( col_in_701     ),
    .col_in_702              ( col_in_702     ),
    .col_in_703              ( col_in_703     ),
    .col_in_704              ( col_in_704     ),
    .col_in_705              ( col_in_705     ),
    .col_in_706              ( col_in_706     ),
    .col_in_707              ( col_in_707     ),
    .col_in_708              ( col_in_708     ),
    .col_in_709              ( col_in_709     ),
    .col_in_710              ( col_in_710     ),
    .col_in_711              ( col_in_711     ),
    .col_in_712              ( col_in_712     ),
    .col_in_713              ( col_in_713     ),
    .col_in_714              ( col_in_714     ),
    .col_in_715              ( col_in_715     ),
    .col_in_716              ( col_in_716     ),
    .col_in_717              ( col_in_717     ),
    .col_in_718              ( col_in_718     ),
    .col_in_719              ( col_in_719     ),
    .col_in_720              ( col_in_720     ),
    .col_in_721              ( col_in_721     ),
    .col_in_722              ( col_in_722     ),
    .col_in_723              ( col_in_723     ),
    .col_in_724              ( col_in_724     ),
    .col_in_725              ( col_in_725     ),
    .col_in_726              ( col_in_726     ),
    .col_in_727              ( col_in_727     ),
    .col_in_728              ( col_in_728     ),
    .col_in_729              ( col_in_729     ),
    .col_in_730              ( col_in_730     ),
    .col_in_731              ( col_in_731     ),
    .col_in_732              ( col_in_732     ),
    .col_in_733              ( col_in_733     ),
    .col_in_734              ( col_in_734     ),
    .col_in_735              ( col_in_735     ),
    .col_in_736              ( col_in_736     ),
    .col_in_737              ( col_in_737     ),
    .col_in_738              ( col_in_738     ),
    .col_in_739              ( col_in_739     ),
    .col_in_740              ( col_in_740     ),
    .col_in_741              ( col_in_741     ),
    .col_in_742              ( col_in_742     ),
    .col_in_743              ( col_in_743     ),
    .col_in_744              ( col_in_744     ),
    .col_in_745              ( col_in_745     ),
    .col_in_746              ( col_in_746     ),
    .col_in_747              ( col_in_747     ),
    .col_in_748              ( col_in_748     ),
    .col_in_749              ( col_in_749     ),
    .col_in_750              ( col_in_750     ),
    .col_in_751              ( col_in_751     ),
    .col_in_752              ( col_in_752     ),
    .col_in_753              ( col_in_753     ),
    .col_in_754              ( col_in_754     ),
    .col_in_755              ( col_in_755     ),
    .col_in_756              ( col_in_756     ),
    .col_in_757              ( col_in_757     ),
    .col_in_758              ( col_in_758     ),
    .col_in_759              ( col_in_759     ),
    .col_in_760              ( col_in_760     ),
    .col_in_761              ( col_in_761     ),
    .col_in_762              ( col_in_762     ),
    .col_in_763              ( col_in_763     ),
    .col_in_764              ( col_in_764     ),
    .col_in_765              ( col_in_765     ),
    .col_in_766              ( col_in_766     ),
    .col_in_767              ( col_in_767     ),
    .col_in_768              ( col_in_768     ),
    .col_in_769              ( col_in_769     ),
    .col_in_770              ( col_in_770     ),
    .col_in_771              ( col_in_771     ),
    .col_in_772              ( col_in_772     ),
    .col_in_773              ( col_in_773     ),
    .col_in_774              ( col_in_774     ),
    .col_in_775              ( col_in_775     ),
    .col_in_776              ( col_in_776     ),
    .col_in_777              ( col_in_777     ),
    .col_in_778              ( col_in_778     ),
    .col_in_779              ( col_in_779     ),
    .col_in_780              ( col_in_780     ),
    .col_in_781              ( col_in_781     ),
    .col_in_782              ( col_in_782     ),
    .col_in_783              ( col_in_783     ),
    .col_in_784              ( col_in_784     ),
    .col_in_785              ( col_in_785     ),
    .col_in_786              ( col_in_786     ),
    .col_in_787              ( col_in_787     ),
    .col_in_788              ( col_in_788     ),
    .col_in_789              ( col_in_789     ),
    .col_in_790              ( col_in_790     ),
    .col_in_791              ( col_in_791     ),
    .col_in_792              ( col_in_792     ),
    .col_in_793              ( col_in_793     ),
    .col_in_794              ( col_in_794     ),
    .col_in_795              ( col_in_795     ),
    .col_in_796              ( col_in_796     ),
    .col_in_797              ( col_in_797     ),
    .col_in_798              ( col_in_798     ),
    .col_in_799              ( col_in_799     ),
    .col_in_800              ( col_in_800     ),
    .col_in_801              ( col_in_801     ),
    .col_in_802              ( col_in_802     ),
    .col_in_803              ( col_in_803     ),
    .col_in_804              ( col_in_804     ),
    .col_in_805              ( col_in_805     ),
    .col_in_806              ( col_in_806     ),
    .col_in_807              ( col_in_807     ),
    .col_in_808              ( col_in_808     ),
    .col_in_809              ( col_in_809     ),
    .col_in_810              ( col_in_810     ),
    .col_in_811              ( col_in_811     ),
    .col_in_812              ( col_in_812     ),
    .col_in_813              ( col_in_813     ),
    .col_in_814              ( col_in_814     ),
    .col_in_815              ( col_in_815     ),
    .col_in_816              ( col_in_816     ),
    .col_in_817              ( col_in_817     ),
    .col_in_818              ( col_in_818     ),
    .col_in_819              ( col_in_819     ),
    .col_in_820              ( col_in_820     ),
    .col_in_821              ( col_in_821     ),
    .col_in_822              ( col_in_822     ),
    .col_in_823              ( col_in_823     ),
    .col_in_824              ( col_in_824     ),
    .col_in_825              ( col_in_825     ),
    .col_in_826              ( col_in_826     ),
    .col_in_827              ( col_in_827     ),
    .col_in_828              ( col_in_828     ),
    .col_in_829              ( col_in_829     ),
    .col_in_830              ( col_in_830     ),
    .col_in_831              ( col_in_831     ),
    .col_in_832              ( col_in_832     ),
    .col_in_833              ( col_in_833     ),
    .col_in_834              ( col_in_834     ),
    .col_in_835              ( col_in_835     ),
    .col_in_836              ( col_in_836     ),
    .col_in_837              ( col_in_837     ),
    .col_in_838              ( col_in_838     ),
    .col_in_839              ( col_in_839     ),
    .col_in_840              ( col_in_840     ),
    .col_in_841              ( col_in_841     ),
    .col_in_842              ( col_in_842     ),
    .col_in_843              ( col_in_843     ),
    .col_in_844              ( col_in_844     ),
    .col_in_845              ( col_in_845     ),
    .col_in_846              ( col_in_846     ),
    .col_in_847              ( col_in_847     ),
    .col_in_848              ( col_in_848     ),
    .col_in_849              ( col_in_849     ),
    .col_in_850              ( col_in_850     ),
    .col_in_851              ( col_in_851     ),
    .col_in_852              ( col_in_852     ),
    .col_in_853              ( col_in_853     ),
    .col_in_854              ( col_in_854     ),
    .col_in_855              ( col_in_855     ),
    .col_in_856              ( col_in_856     ),
    .col_in_857              ( col_in_857     ),
    .col_in_858              ( col_in_858     ),
    .col_in_859              ( col_in_859     ),
    .col_in_860              ( col_in_860     ),
    .col_in_861              ( col_in_861     ),
    .col_in_862              ( col_in_862     ),
    .col_in_863              ( col_in_863     ),
    .col_in_864              ( col_in_864     ),
    .col_in_865              ( col_in_865     ),
    .col_in_866              ( col_in_866     ),
    .col_in_867              ( col_in_867     ),
    .col_in_868              ( col_in_868     ),
    .col_in_869              ( col_in_869     ),
    .col_in_870              ( col_in_870     ),
    .col_in_871              ( col_in_871     ),
    .col_in_872              ( col_in_872     ),
    .col_in_873              ( col_in_873     ),
    .col_in_874              ( col_in_874     ),
    .col_in_875              ( col_in_875     ),
    .col_in_876              ( col_in_876     ),
    .col_in_877              ( col_in_877     ),
    .col_in_878              ( col_in_878     ),
    .col_in_879              ( col_in_879     ),
    .col_in_880              ( col_in_880     ),
    .col_in_881              ( col_in_881     ),
    .col_in_882              ( col_in_882     ),
    .col_in_883              ( col_in_883     ),
    .col_in_884              ( col_in_884     ),
    .col_in_885              ( col_in_885     ),
    .col_in_886              ( col_in_886     ),
    .col_in_887              ( col_in_887     ),
    .col_in_888              ( col_in_888     ),
    .col_in_889              ( col_in_889     ),
    .col_in_890              ( col_in_890     ),
    .col_in_891              ( col_in_891     ),
    .col_in_892              ( col_in_892     ),
    .col_in_893              ( col_in_893     ),
    .col_in_894              ( col_in_894     ),
    .col_in_895              ( col_in_895     ),
    .col_in_896              ( col_in_896     ),
    .col_in_897              ( col_in_897     ),
    .col_in_898              ( col_in_898     ),
    .col_in_899              ( col_in_899     ),
    .col_in_900              ( col_in_900     ),
    .col_in_901              ( col_in_901     ),
    .col_in_902              ( col_in_902     ),
    .col_in_903              ( col_in_903     ),
    .col_in_904              ( col_in_904     ),
    .col_in_905              ( col_in_905     ),
    .col_in_906              ( col_in_906     ),
    .col_in_907              ( col_in_907     ),
    .col_in_908              ( col_in_908     ),
    .col_in_909              ( col_in_909     ),
    .col_in_910              ( col_in_910     ),
    .col_in_911              ( col_in_911     ),
    .col_in_912              ( col_in_912     ),
    .col_in_913              ( col_in_913     ),
    .col_in_914              ( col_in_914     ),
    .col_in_915              ( col_in_915     ),
    .col_in_916              ( col_in_916     ),
    .col_in_917              ( col_in_917     ),
    .col_in_918              ( col_in_918     ),
    .col_in_919              ( col_in_919     ),
    .col_in_920              ( col_in_920     ),
    .col_in_921              ( col_in_921     ),
    .col_in_922              ( col_in_922     ),
    .col_in_923              ( col_in_923     ),
    .col_in_924              ( col_in_924     ),
    .col_in_925              ( col_in_925     ),
    .col_in_926              ( col_in_926     ),
    .col_in_927              ( col_in_927     ),
    .col_in_928              ( col_in_928     ),
    .col_in_929              ( col_in_929     ),
    .col_in_930              ( col_in_930     ),
    .col_in_931              ( col_in_931     ),
    .col_in_932              ( col_in_932     ),
    .col_in_933              ( col_in_933     ),
    .col_in_934              ( col_in_934     ),
    .col_in_935              ( col_in_935     ),
    .col_in_936              ( col_in_936     ),
    .col_in_937              ( col_in_937     ),
    .col_in_938              ( col_in_938     ),
    .col_in_939              ( col_in_939     ),
    .col_in_940              ( col_in_940     ),
    .col_in_941              ( col_in_941     ),
    .col_in_942              ( col_in_942     ),
    .col_in_943              ( col_in_943     ),
    .col_in_944              ( col_in_944     ),
    .col_in_945              ( col_in_945     ),
    .col_in_946              ( col_in_946     ),
    .col_in_947              ( col_in_947     ),
    .col_in_948              ( col_in_948     ),
    .col_in_949              ( col_in_949     ),
    .col_in_950              ( col_in_950     ),
    .col_in_951              ( col_in_951     ),
    .col_in_952              ( col_in_952     ),
    .col_in_953              ( col_in_953     ),
    .col_in_954              ( col_in_954     ),
    .col_in_955              ( col_in_955     ),
    .col_in_956              ( col_in_956     ),
    .col_in_957              ( col_in_957     ),
    .col_in_958              ( col_in_958     ),
    .col_in_959              ( col_in_959     ),
    .col_in_960              ( col_in_960     ),
    .col_in_961              ( col_in_961     ),
    .col_in_962              ( col_in_962     ),
    .col_in_963              ( col_in_963     ),
    .col_in_964              ( col_in_964     ),
    .col_in_965              ( col_in_965     ),
    .col_in_966              ( col_in_966     ),
    .col_in_967              ( col_in_967     ),
    .col_in_968              ( col_in_968     ),
    .col_in_969              ( col_in_969     ),
    .col_in_970              ( col_in_970     ),
    .col_in_971              ( col_in_971     ),
    .col_in_972              ( col_in_972     ),
    .col_in_973              ( col_in_973     ),
    .col_in_974              ( col_in_974     ),
    .col_in_975              ( col_in_975     ),
    .col_in_976              ( col_in_976     ),
    .col_in_977              ( col_in_977     ),
    .col_in_978              ( col_in_978     ),
    .col_in_979              ( col_in_979     ),
    .col_in_980              ( col_in_980     ),
    .col_in_981              ( col_in_981     ),
    .col_in_982              ( col_in_982     ),
    .col_in_983              ( col_in_983     ),
    .col_in_984              ( col_in_984     ),
    .col_in_985              ( col_in_985     ),
    .col_in_986              ( col_in_986     ),
    .col_in_987              ( col_in_987     ),
    .col_in_988              ( col_in_988     ),
    .col_in_989              ( col_in_989     ),
    .col_in_990              ( col_in_990     ),
    .col_in_991              ( col_in_991     ),
    .col_in_992              ( col_in_992     ),
    .col_in_993              ( col_in_993     ),
    .col_in_994              ( col_in_994     ),
    .col_in_995              ( col_in_995     ),
    .col_in_996              ( col_in_996     ),
    .col_in_997              ( col_in_997     ),
    .col_in_998              ( col_in_998     ),
    .col_in_999              ( col_in_999     ),
    .col_in_1000             ( col_in_1000    ),
    .col_in_1001             ( col_in_1001    ),
    .col_in_1002             ( col_in_1002    ),
    .col_in_1003             ( col_in_1003    ),
    .col_in_1004             ( col_in_1004    ),
    .col_in_1005             ( col_in_1005    ),
    .col_in_1006             ( col_in_1006    ),
    .col_in_1007             ( col_in_1007    ),
    .col_in_1008             ( col_in_1008    ),
    .col_in_1009             ( col_in_1009    ),
    .col_in_1010             ( col_in_1010    ),
    .col_in_1011             ( col_in_1011    ),
    .col_in_1012             ( col_in_1012    ),
    .col_in_1013             ( col_in_1013    ),
    .col_in_1014             ( col_in_1014    ),
    .col_in_1015             ( col_in_1015    ),
    .col_in_1016             ( col_in_1016    ),
    .col_in_1017             ( col_in_1017    ),
    .col_in_1018             ( col_in_1018    ),
    .col_in_1019             ( col_in_1019    ),
    .col_in_1020             ( col_in_1020    ),
    .col_in_1021             ( col_in_1021    ),
    .col_in_1022             ( col_in_1022    ),
    .col_in_1023             ( col_in_1023    ),
    .col_in_1024             ( col_in_1024    ),
    .col_in_1025             ( col_in_1025    ),
    .col_in_1026             ( col_in_1026    ),
    .col_in_1027             ( col_in_1027    ),
    .col_in_1028             ( col_in_1028    ),
    .col_in_1029             ( col_in_1029    ),
    .col_in_1030             ( col_in_1030    ),
    .col_in_1031             ( col_in_1031    ),
    .col_in_1032             ( col_in_1032    ),

    .col_out_0               ( u0_col_out_0      ),
    .col_out_1               ( u0_col_out_1      ),
    .col_out_2               ( u0_col_out_2      ),
    .col_out_3               ( u0_col_out_3      ),
    .col_out_4               ( u0_col_out_4      ),
    .col_out_5               ( u0_col_out_5      ),
    .col_out_6               ( u0_col_out_6      ),
    .col_out_7               ( u0_col_out_7      ),
    .col_out_8               ( u0_col_out_8      ),
    .col_out_9               ( u0_col_out_9      ),
    .col_out_10              ( u0_col_out_10     ),
    .col_out_11              ( u0_col_out_11     ),
    .col_out_12              ( u0_col_out_12     ),
    .col_out_13              ( u0_col_out_13     ),
    .col_out_14              ( u0_col_out_14     ),
    .col_out_15              ( u0_col_out_15     ),
    .col_out_16              ( u0_col_out_16     ),
    .col_out_17              ( u0_col_out_17     ),
    .col_out_18              ( u0_col_out_18     ),
    .col_out_19              ( u0_col_out_19     ),
    .col_out_20              ( u0_col_out_20     ),
    .col_out_21              ( u0_col_out_21     ),
    .col_out_22              ( u0_col_out_22     ),
    .col_out_23              ( u0_col_out_23     ),
    .col_out_24              ( u0_col_out_24     ),
    .col_out_25              ( u0_col_out_25     ),
    .col_out_26              ( u0_col_out_26     ),
    .col_out_27              ( u0_col_out_27     ),
    .col_out_28              ( u0_col_out_28     ),
    .col_out_29              ( u0_col_out_29     ),
    .col_out_30              ( u0_col_out_30     ),
    .col_out_31              ( u0_col_out_31     ),
    .col_out_32              ( u0_col_out_32     ),
    .col_out_33              ( u0_col_out_33     ),
    .col_out_34              ( u0_col_out_34     ),
    .col_out_35              ( u0_col_out_35     ),
    .col_out_36              ( u0_col_out_36     ),
    .col_out_37              ( u0_col_out_37     ),
    .col_out_38              ( u0_col_out_38     ),
    .col_out_39              ( u0_col_out_39     ),
    .col_out_40              ( u0_col_out_40     ),
    .col_out_41              ( u0_col_out_41     ),
    .col_out_42              ( u0_col_out_42     ),
    .col_out_43              ( u0_col_out_43     ),
    .col_out_44              ( u0_col_out_44     ),
    .col_out_45              ( u0_col_out_45     ),
    .col_out_46              ( u0_col_out_46     ),
    .col_out_47              ( u0_col_out_47     ),
    .col_out_48              ( u0_col_out_48     ),
    .col_out_49              ( u0_col_out_49     ),
    .col_out_50              ( u0_col_out_50     ),
    .col_out_51              ( u0_col_out_51     ),
    .col_out_52              ( u0_col_out_52     ),
    .col_out_53              ( u0_col_out_53     ),
    .col_out_54              ( u0_col_out_54     ),
    .col_out_55              ( u0_col_out_55     ),
    .col_out_56              ( u0_col_out_56     ),
    .col_out_57              ( u0_col_out_57     ),
    .col_out_58              ( u0_col_out_58     ),
    .col_out_59              ( u0_col_out_59     ),
    .col_out_60              ( u0_col_out_60     ),
    .col_out_61              ( u0_col_out_61     ),
    .col_out_62              ( u0_col_out_62     ),
    .col_out_63              ( u0_col_out_63     ),
    .col_out_64              ( u0_col_out_64     ),
    .col_out_65              ( u0_col_out_65     ),
    .col_out_66              ( u0_col_out_66     ),
    .col_out_67              ( u0_col_out_67     ),
    .col_out_68              ( u0_col_out_68     ),
    .col_out_69              ( u0_col_out_69     ),
    .col_out_70              ( u0_col_out_70     ),
    .col_out_71              ( u0_col_out_71     ),
    .col_out_72              ( u0_col_out_72     ),
    .col_out_73              ( u0_col_out_73     ),
    .col_out_74              ( u0_col_out_74     ),
    .col_out_75              ( u0_col_out_75     ),
    .col_out_76              ( u0_col_out_76     ),
    .col_out_77              ( u0_col_out_77     ),
    .col_out_78              ( u0_col_out_78     ),
    .col_out_79              ( u0_col_out_79     ),
    .col_out_80              ( u0_col_out_80     ),
    .col_out_81              ( u0_col_out_81     ),
    .col_out_82              ( u0_col_out_82     ),
    .col_out_83              ( u0_col_out_83     ),
    .col_out_84              ( u0_col_out_84     ),
    .col_out_85              ( u0_col_out_85     ),
    .col_out_86              ( u0_col_out_86     ),
    .col_out_87              ( u0_col_out_87     ),
    .col_out_88              ( u0_col_out_88     ),
    .col_out_89              ( u0_col_out_89     ),
    .col_out_90              ( u0_col_out_90     ),
    .col_out_91              ( u0_col_out_91     ),
    .col_out_92              ( u0_col_out_92     ),
    .col_out_93              ( u0_col_out_93     ),
    .col_out_94              ( u0_col_out_94     ),
    .col_out_95              ( u0_col_out_95     ),
    .col_out_96              ( u0_col_out_96     ),
    .col_out_97              ( u0_col_out_97     ),
    .col_out_98              ( u0_col_out_98     ),
    .col_out_99              ( u0_col_out_99     ),
    .col_out_100             ( u0_col_out_100    ),
    .col_out_101             ( u0_col_out_101    ),
    .col_out_102             ( u0_col_out_102    ),
    .col_out_103             ( u0_col_out_103    ),
    .col_out_104             ( u0_col_out_104    ),
    .col_out_105             ( u0_col_out_105    ),
    .col_out_106             ( u0_col_out_106    ),
    .col_out_107             ( u0_col_out_107    ),
    .col_out_108             ( u0_col_out_108    ),
    .col_out_109             ( u0_col_out_109    ),
    .col_out_110             ( u0_col_out_110    ),
    .col_out_111             ( u0_col_out_111    ),
    .col_out_112             ( u0_col_out_112    ),
    .col_out_113             ( u0_col_out_113    ),
    .col_out_114             ( u0_col_out_114    ),
    .col_out_115             ( u0_col_out_115    ),
    .col_out_116             ( u0_col_out_116    ),
    .col_out_117             ( u0_col_out_117    ),
    .col_out_118             ( u0_col_out_118    ),
    .col_out_119             ( u0_col_out_119    ),
    .col_out_120             ( u0_col_out_120    ),
    .col_out_121             ( u0_col_out_121    ),
    .col_out_122             ( u0_col_out_122    ),
    .col_out_123             ( u0_col_out_123    ),
    .col_out_124             ( u0_col_out_124    ),
    .col_out_125             ( u0_col_out_125    ),
    .col_out_126             ( u0_col_out_126    ),
    .col_out_127             ( u0_col_out_127    ),
    .col_out_128             ( u0_col_out_128    ),
    .col_out_129             ( u0_col_out_129    ),
    .col_out_130             ( u0_col_out_130    ),
    .col_out_131             ( u0_col_out_131    ),
    .col_out_132             ( u0_col_out_132    ),
    .col_out_133             ( u0_col_out_133    ),
    .col_out_134             ( u0_col_out_134    ),
    .col_out_135             ( u0_col_out_135    ),
    .col_out_136             ( u0_col_out_136    ),
    .col_out_137             ( u0_col_out_137    ),
    .col_out_138             ( u0_col_out_138    ),
    .col_out_139             ( u0_col_out_139    ),
    .col_out_140             ( u0_col_out_140    ),
    .col_out_141             ( u0_col_out_141    ),
    .col_out_142             ( u0_col_out_142    ),
    .col_out_143             ( u0_col_out_143    ),
    .col_out_144             ( u0_col_out_144    ),
    .col_out_145             ( u0_col_out_145    ),
    .col_out_146             ( u0_col_out_146    ),
    .col_out_147             ( u0_col_out_147    ),
    .col_out_148             ( u0_col_out_148    ),
    .col_out_149             ( u0_col_out_149    ),
    .col_out_150             ( u0_col_out_150    ),
    .col_out_151             ( u0_col_out_151    ),
    .col_out_152             ( u0_col_out_152    ),
    .col_out_153             ( u0_col_out_153    ),
    .col_out_154             ( u0_col_out_154    ),
    .col_out_155             ( u0_col_out_155    ),
    .col_out_156             ( u0_col_out_156    ),
    .col_out_157             ( u0_col_out_157    ),
    .col_out_158             ( u0_col_out_158    ),
    .col_out_159             ( u0_col_out_159    ),
    .col_out_160             ( u0_col_out_160    ),
    .col_out_161             ( u0_col_out_161    ),
    .col_out_162             ( u0_col_out_162    ),
    .col_out_163             ( u0_col_out_163    ),
    .col_out_164             ( u0_col_out_164    ),
    .col_out_165             ( u0_col_out_165    ),
    .col_out_166             ( u0_col_out_166    ),
    .col_out_167             ( u0_col_out_167    ),
    .col_out_168             ( u0_col_out_168    ),
    .col_out_169             ( u0_col_out_169    ),
    .col_out_170             ( u0_col_out_170    ),
    .col_out_171             ( u0_col_out_171    ),
    .col_out_172             ( u0_col_out_172    ),
    .col_out_173             ( u0_col_out_173    ),
    .col_out_174             ( u0_col_out_174    ),
    .col_out_175             ( u0_col_out_175    ),
    .col_out_176             ( u0_col_out_176    ),
    .col_out_177             ( u0_col_out_177    ),
    .col_out_178             ( u0_col_out_178    ),
    .col_out_179             ( u0_col_out_179    ),
    .col_out_180             ( u0_col_out_180    ),
    .col_out_181             ( u0_col_out_181    ),
    .col_out_182             ( u0_col_out_182    ),
    .col_out_183             ( u0_col_out_183    ),
    .col_out_184             ( u0_col_out_184    ),
    .col_out_185             ( u0_col_out_185    ),
    .col_out_186             ( u0_col_out_186    ),
    .col_out_187             ( u0_col_out_187    ),
    .col_out_188             ( u0_col_out_188    ),
    .col_out_189             ( u0_col_out_189    ),
    .col_out_190             ( u0_col_out_190    ),
    .col_out_191             ( u0_col_out_191    ),
    .col_out_192             ( u0_col_out_192    ),
    .col_out_193             ( u0_col_out_193    ),
    .col_out_194             ( u0_col_out_194    ),
    .col_out_195             ( u0_col_out_195    ),
    .col_out_196             ( u0_col_out_196    ),
    .col_out_197             ( u0_col_out_197    ),
    .col_out_198             ( u0_col_out_198    ),
    .col_out_199             ( u0_col_out_199    ),
    .col_out_200             ( u0_col_out_200    ),
    .col_out_201             ( u0_col_out_201    ),
    .col_out_202             ( u0_col_out_202    ),
    .col_out_203             ( u0_col_out_203    ),
    .col_out_204             ( u0_col_out_204    ),
    .col_out_205             ( u0_col_out_205    ),
    .col_out_206             ( u0_col_out_206    ),
    .col_out_207             ( u0_col_out_207    ),
    .col_out_208             ( u0_col_out_208    ),
    .col_out_209             ( u0_col_out_209    ),
    .col_out_210             ( u0_col_out_210    ),
    .col_out_211             ( u0_col_out_211    ),
    .col_out_212             ( u0_col_out_212    ),
    .col_out_213             ( u0_col_out_213    ),
    .col_out_214             ( u0_col_out_214    ),
    .col_out_215             ( u0_col_out_215    ),
    .col_out_216             ( u0_col_out_216    ),
    .col_out_217             ( u0_col_out_217    ),
    .col_out_218             ( u0_col_out_218    ),
    .col_out_219             ( u0_col_out_219    ),
    .col_out_220             ( u0_col_out_220    ),
    .col_out_221             ( u0_col_out_221    ),
    .col_out_222             ( u0_col_out_222    ),
    .col_out_223             ( u0_col_out_223    ),
    .col_out_224             ( u0_col_out_224    ),
    .col_out_225             ( u0_col_out_225    ),
    .col_out_226             ( u0_col_out_226    ),
    .col_out_227             ( u0_col_out_227    ),
    .col_out_228             ( u0_col_out_228    ),
    .col_out_229             ( u0_col_out_229    ),
    .col_out_230             ( u0_col_out_230    ),
    .col_out_231             ( u0_col_out_231    ),
    .col_out_232             ( u0_col_out_232    ),
    .col_out_233             ( u0_col_out_233    ),
    .col_out_234             ( u0_col_out_234    ),
    .col_out_235             ( u0_col_out_235    ),
    .col_out_236             ( u0_col_out_236    ),
    .col_out_237             ( u0_col_out_237    ),
    .col_out_238             ( u0_col_out_238    ),
    .col_out_239             ( u0_col_out_239    ),
    .col_out_240             ( u0_col_out_240    ),
    .col_out_241             ( u0_col_out_241    ),
    .col_out_242             ( u0_col_out_242    ),
    .col_out_243             ( u0_col_out_243    ),
    .col_out_244             ( u0_col_out_244    ),
    .col_out_245             ( u0_col_out_245    ),
    .col_out_246             ( u0_col_out_246    ),
    .col_out_247             ( u0_col_out_247    ),
    .col_out_248             ( u0_col_out_248    ),
    .col_out_249             ( u0_col_out_249    ),
    .col_out_250             ( u0_col_out_250    ),
    .col_out_251             ( u0_col_out_251    ),
    .col_out_252             ( u0_col_out_252    ),
    .col_out_253             ( u0_col_out_253    ),
    .col_out_254             ( u0_col_out_254    ),
    .col_out_255             ( u0_col_out_255    ),
    .col_out_256             ( u0_col_out_256    ),
    .col_out_257             ( u0_col_out_257    ),
    .col_out_258             ( u0_col_out_258    ),
    .col_out_259             ( u0_col_out_259    ),
    .col_out_260             ( u0_col_out_260    ),
    .col_out_261             ( u0_col_out_261    ),
    .col_out_262             ( u0_col_out_262    ),
    .col_out_263             ( u0_col_out_263    ),
    .col_out_264             ( u0_col_out_264    ),
    .col_out_265             ( u0_col_out_265    ),
    .col_out_266             ( u0_col_out_266    ),
    .col_out_267             ( u0_col_out_267    ),
    .col_out_268             ( u0_col_out_268    ),
    .col_out_269             ( u0_col_out_269    ),
    .col_out_270             ( u0_col_out_270    ),
    .col_out_271             ( u0_col_out_271    ),
    .col_out_272             ( u0_col_out_272    ),
    .col_out_273             ( u0_col_out_273    ),
    .col_out_274             ( u0_col_out_274    ),
    .col_out_275             ( u0_col_out_275    ),
    .col_out_276             ( u0_col_out_276    ),
    .col_out_277             ( u0_col_out_277    ),
    .col_out_278             ( u0_col_out_278    ),
    .col_out_279             ( u0_col_out_279    ),
    .col_out_280             ( u0_col_out_280    ),
    .col_out_281             ( u0_col_out_281    ),
    .col_out_282             ( u0_col_out_282    ),
    .col_out_283             ( u0_col_out_283    ),
    .col_out_284             ( u0_col_out_284    ),
    .col_out_285             ( u0_col_out_285    ),
    .col_out_286             ( u0_col_out_286    ),
    .col_out_287             ( u0_col_out_287    ),
    .col_out_288             ( u0_col_out_288    ),
    .col_out_289             ( u0_col_out_289    ),
    .col_out_290             ( u0_col_out_290    ),
    .col_out_291             ( u0_col_out_291    ),
    .col_out_292             ( u0_col_out_292    ),
    .col_out_293             ( u0_col_out_293    ),
    .col_out_294             ( u0_col_out_294    ),
    .col_out_295             ( u0_col_out_295    ),
    .col_out_296             ( u0_col_out_296    ),
    .col_out_297             ( u0_col_out_297    ),
    .col_out_298             ( u0_col_out_298    ),
    .col_out_299             ( u0_col_out_299    ),
    .col_out_300             ( u0_col_out_300    ),
    .col_out_301             ( u0_col_out_301    ),
    .col_out_302             ( u0_col_out_302    ),
    .col_out_303             ( u0_col_out_303    ),
    .col_out_304             ( u0_col_out_304    ),
    .col_out_305             ( u0_col_out_305    ),
    .col_out_306             ( u0_col_out_306    ),
    .col_out_307             ( u0_col_out_307    ),
    .col_out_308             ( u0_col_out_308    ),
    .col_out_309             ( u0_col_out_309    ),
    .col_out_310             ( u0_col_out_310    ),
    .col_out_311             ( u0_col_out_311    ),
    .col_out_312             ( u0_col_out_312    ),
    .col_out_313             ( u0_col_out_313    ),
    .col_out_314             ( u0_col_out_314    ),
    .col_out_315             ( u0_col_out_315    ),
    .col_out_316             ( u0_col_out_316    ),
    .col_out_317             ( u0_col_out_317    ),
    .col_out_318             ( u0_col_out_318    ),
    .col_out_319             ( u0_col_out_319    ),
    .col_out_320             ( u0_col_out_320    ),
    .col_out_321             ( u0_col_out_321    ),
    .col_out_322             ( u0_col_out_322    ),
    .col_out_323             ( u0_col_out_323    ),
    .col_out_324             ( u0_col_out_324    ),
    .col_out_325             ( u0_col_out_325    ),
    .col_out_326             ( u0_col_out_326    ),
    .col_out_327             ( u0_col_out_327    ),
    .col_out_328             ( u0_col_out_328    ),
    .col_out_329             ( u0_col_out_329    ),
    .col_out_330             ( u0_col_out_330    ),
    .col_out_331             ( u0_col_out_331    ),
    .col_out_332             ( u0_col_out_332    ),
    .col_out_333             ( u0_col_out_333    ),
    .col_out_334             ( u0_col_out_334    ),
    .col_out_335             ( u0_col_out_335    ),
    .col_out_336             ( u0_col_out_336    ),
    .col_out_337             ( u0_col_out_337    ),
    .col_out_338             ( u0_col_out_338    ),
    .col_out_339             ( u0_col_out_339    ),
    .col_out_340             ( u0_col_out_340    ),
    .col_out_341             ( u0_col_out_341    ),
    .col_out_342             ( u0_col_out_342    ),
    .col_out_343             ( u0_col_out_343    ),
    .col_out_344             ( u0_col_out_344    ),
    .col_out_345             ( u0_col_out_345    ),
    .col_out_346             ( u0_col_out_346    ),
    .col_out_347             ( u0_col_out_347    ),
    .col_out_348             ( u0_col_out_348    ),
    .col_out_349             ( u0_col_out_349    ),
    .col_out_350             ( u0_col_out_350    ),
    .col_out_351             ( u0_col_out_351    ),
    .col_out_352             ( u0_col_out_352    ),
    .col_out_353             ( u0_col_out_353    ),
    .col_out_354             ( u0_col_out_354    ),
    .col_out_355             ( u0_col_out_355    ),
    .col_out_356             ( u0_col_out_356    ),
    .col_out_357             ( u0_col_out_357    ),
    .col_out_358             ( u0_col_out_358    ),
    .col_out_359             ( u0_col_out_359    ),
    .col_out_360             ( u0_col_out_360    ),
    .col_out_361             ( u0_col_out_361    ),
    .col_out_362             ( u0_col_out_362    ),
    .col_out_363             ( u0_col_out_363    ),
    .col_out_364             ( u0_col_out_364    ),
    .col_out_365             ( u0_col_out_365    ),
    .col_out_366             ( u0_col_out_366    ),
    .col_out_367             ( u0_col_out_367    ),
    .col_out_368             ( u0_col_out_368    ),
    .col_out_369             ( u0_col_out_369    ),
    .col_out_370             ( u0_col_out_370    ),
    .col_out_371             ( u0_col_out_371    ),
    .col_out_372             ( u0_col_out_372    ),
    .col_out_373             ( u0_col_out_373    ),
    .col_out_374             ( u0_col_out_374    ),
    .col_out_375             ( u0_col_out_375    ),
    .col_out_376             ( u0_col_out_376    ),
    .col_out_377             ( u0_col_out_377    ),
    .col_out_378             ( u0_col_out_378    ),
    .col_out_379             ( u0_col_out_379    ),
    .col_out_380             ( u0_col_out_380    ),
    .col_out_381             ( u0_col_out_381    ),
    .col_out_382             ( u0_col_out_382    ),
    .col_out_383             ( u0_col_out_383    ),
    .col_out_384             ( u0_col_out_384    ),
    .col_out_385             ( u0_col_out_385    ),
    .col_out_386             ( u0_col_out_386    ),
    .col_out_387             ( u0_col_out_387    ),
    .col_out_388             ( u0_col_out_388    ),
    .col_out_389             ( u0_col_out_389    ),
    .col_out_390             ( u0_col_out_390    ),
    .col_out_391             ( u0_col_out_391    ),
    .col_out_392             ( u0_col_out_392    ),
    .col_out_393             ( u0_col_out_393    ),
    .col_out_394             ( u0_col_out_394    ),
    .col_out_395             ( u0_col_out_395    ),
    .col_out_396             ( u0_col_out_396    ),
    .col_out_397             ( u0_col_out_397    ),
    .col_out_398             ( u0_col_out_398    ),
    .col_out_399             ( u0_col_out_399    ),
    .col_out_400             ( u0_col_out_400    ),
    .col_out_401             ( u0_col_out_401    ),
    .col_out_402             ( u0_col_out_402    ),
    .col_out_403             ( u0_col_out_403    ),
    .col_out_404             ( u0_col_out_404    ),
    .col_out_405             ( u0_col_out_405    ),
    .col_out_406             ( u0_col_out_406    ),
    .col_out_407             ( u0_col_out_407    ),
    .col_out_408             ( u0_col_out_408    ),
    .col_out_409             ( u0_col_out_409    ),
    .col_out_410             ( u0_col_out_410    ),
    .col_out_411             ( u0_col_out_411    ),
    .col_out_412             ( u0_col_out_412    ),
    .col_out_413             ( u0_col_out_413    ),
    .col_out_414             ( u0_col_out_414    ),
    .col_out_415             ( u0_col_out_415    ),
    .col_out_416             ( u0_col_out_416    ),
    .col_out_417             ( u0_col_out_417    ),
    .col_out_418             ( u0_col_out_418    ),
    .col_out_419             ( u0_col_out_419    ),
    .col_out_420             ( u0_col_out_420    ),
    .col_out_421             ( u0_col_out_421    ),
    .col_out_422             ( u0_col_out_422    ),
    .col_out_423             ( u0_col_out_423    ),
    .col_out_424             ( u0_col_out_424    ),
    .col_out_425             ( u0_col_out_425    ),
    .col_out_426             ( u0_col_out_426    ),
    .col_out_427             ( u0_col_out_427    ),
    .col_out_428             ( u0_col_out_428    ),
    .col_out_429             ( u0_col_out_429    ),
    .col_out_430             ( u0_col_out_430    ),
    .col_out_431             ( u0_col_out_431    ),
    .col_out_432             ( u0_col_out_432    ),
    .col_out_433             ( u0_col_out_433    ),
    .col_out_434             ( u0_col_out_434    ),
    .col_out_435             ( u0_col_out_435    ),
    .col_out_436             ( u0_col_out_436    ),
    .col_out_437             ( u0_col_out_437    ),
    .col_out_438             ( u0_col_out_438    ),
    .col_out_439             ( u0_col_out_439    ),
    .col_out_440             ( u0_col_out_440    ),
    .col_out_441             ( u0_col_out_441    ),
    .col_out_442             ( u0_col_out_442    ),
    .col_out_443             ( u0_col_out_443    ),
    .col_out_444             ( u0_col_out_444    ),
    .col_out_445             ( u0_col_out_445    ),
    .col_out_446             ( u0_col_out_446    ),
    .col_out_447             ( u0_col_out_447    ),
    .col_out_448             ( u0_col_out_448    ),
    .col_out_449             ( u0_col_out_449    ),
    .col_out_450             ( u0_col_out_450    ),
    .col_out_451             ( u0_col_out_451    ),
    .col_out_452             ( u0_col_out_452    ),
    .col_out_453             ( u0_col_out_453    ),
    .col_out_454             ( u0_col_out_454    ),
    .col_out_455             ( u0_col_out_455    ),
    .col_out_456             ( u0_col_out_456    ),
    .col_out_457             ( u0_col_out_457    ),
    .col_out_458             ( u0_col_out_458    ),
    .col_out_459             ( u0_col_out_459    ),
    .col_out_460             ( u0_col_out_460    ),
    .col_out_461             ( u0_col_out_461    ),
    .col_out_462             ( u0_col_out_462    ),
    .col_out_463             ( u0_col_out_463    ),
    .col_out_464             ( u0_col_out_464    ),
    .col_out_465             ( u0_col_out_465    ),
    .col_out_466             ( u0_col_out_466    ),
    .col_out_467             ( u0_col_out_467    ),
    .col_out_468             ( u0_col_out_468    ),
    .col_out_469             ( u0_col_out_469    ),
    .col_out_470             ( u0_col_out_470    ),
    .col_out_471             ( u0_col_out_471    ),
    .col_out_472             ( u0_col_out_472    ),
    .col_out_473             ( u0_col_out_473    ),
    .col_out_474             ( u0_col_out_474    ),
    .col_out_475             ( u0_col_out_475    ),
    .col_out_476             ( u0_col_out_476    ),
    .col_out_477             ( u0_col_out_477    ),
    .col_out_478             ( u0_col_out_478    ),
    .col_out_479             ( u0_col_out_479    ),
    .col_out_480             ( u0_col_out_480    ),
    .col_out_481             ( u0_col_out_481    ),
    .col_out_482             ( u0_col_out_482    ),
    .col_out_483             ( u0_col_out_483    ),
    .col_out_484             ( u0_col_out_484    ),
    .col_out_485             ( u0_col_out_485    ),
    .col_out_486             ( u0_col_out_486    ),
    .col_out_487             ( u0_col_out_487    ),
    .col_out_488             ( u0_col_out_488    ),
    .col_out_489             ( u0_col_out_489    ),
    .col_out_490             ( u0_col_out_490    ),
    .col_out_491             ( u0_col_out_491    ),
    .col_out_492             ( u0_col_out_492    ),
    .col_out_493             ( u0_col_out_493    ),
    .col_out_494             ( u0_col_out_494    ),
    .col_out_495             ( u0_col_out_495    ),
    .col_out_496             ( u0_col_out_496    ),
    .col_out_497             ( u0_col_out_497    ),
    .col_out_498             ( u0_col_out_498    ),
    .col_out_499             ( u0_col_out_499    ),
    .col_out_500             ( u0_col_out_500    ),
    .col_out_501             ( u0_col_out_501    ),
    .col_out_502             ( u0_col_out_502    ),
    .col_out_503             ( u0_col_out_503    ),
    .col_out_504             ( u0_col_out_504    ),
    .col_out_505             ( u0_col_out_505    ),
    .col_out_506             ( u0_col_out_506    ),
    .col_out_507             ( u0_col_out_507    ),
    .col_out_508             ( u0_col_out_508    ),
    .col_out_509             ( u0_col_out_509    ),
    .col_out_510             ( u0_col_out_510    ),
    .col_out_511             ( u0_col_out_511    ),
    .col_out_512             ( u0_col_out_512    ),
    .col_out_513             ( u0_col_out_513    ),
    .col_out_514             ( u0_col_out_514    ),
    .col_out_515             ( u0_col_out_515    ),
    .col_out_516             ( u0_col_out_516    ),
    .col_out_517             ( u0_col_out_517    ),
    .col_out_518             ( u0_col_out_518    ),
    .col_out_519             ( u0_col_out_519    ),
    .col_out_520             ( u0_col_out_520    ),
    .col_out_521             ( u0_col_out_521    ),
    .col_out_522             ( u0_col_out_522    ),
    .col_out_523             ( u0_col_out_523    ),
    .col_out_524             ( u0_col_out_524    ),
    .col_out_525             ( u0_col_out_525    ),
    .col_out_526             ( u0_col_out_526    ),
    .col_out_527             ( u0_col_out_527    ),
    .col_out_528             ( u0_col_out_528    ),
    .col_out_529             ( u0_col_out_529    ),
    .col_out_530             ( u0_col_out_530    ),
    .col_out_531             ( u0_col_out_531    ),
    .col_out_532             ( u0_col_out_532    ),
    .col_out_533             ( u0_col_out_533    ),
    .col_out_534             ( u0_col_out_534    ),
    .col_out_535             ( u0_col_out_535    ),
    .col_out_536             ( u0_col_out_536    ),
    .col_out_537             ( u0_col_out_537    ),
    .col_out_538             ( u0_col_out_538    ),
    .col_out_539             ( u0_col_out_539    ),
    .col_out_540             ( u0_col_out_540    ),
    .col_out_541             ( u0_col_out_541    ),
    .col_out_542             ( u0_col_out_542    ),
    .col_out_543             ( u0_col_out_543    ),
    .col_out_544             ( u0_col_out_544    ),
    .col_out_545             ( u0_col_out_545    ),
    .col_out_546             ( u0_col_out_546    ),
    .col_out_547             ( u0_col_out_547    ),
    .col_out_548             ( u0_col_out_548    ),
    .col_out_549             ( u0_col_out_549    ),
    .col_out_550             ( u0_col_out_550    ),
    .col_out_551             ( u0_col_out_551    ),
    .col_out_552             ( u0_col_out_552    ),
    .col_out_553             ( u0_col_out_553    ),
    .col_out_554             ( u0_col_out_554    ),
    .col_out_555             ( u0_col_out_555    ),
    .col_out_556             ( u0_col_out_556    ),
    .col_out_557             ( u0_col_out_557    ),
    .col_out_558             ( u0_col_out_558    ),
    .col_out_559             ( u0_col_out_559    ),
    .col_out_560             ( u0_col_out_560    ),
    .col_out_561             ( u0_col_out_561    ),
    .col_out_562             ( u0_col_out_562    ),
    .col_out_563             ( u0_col_out_563    ),
    .col_out_564             ( u0_col_out_564    ),
    .col_out_565             ( u0_col_out_565    ),
    .col_out_566             ( u0_col_out_566    ),
    .col_out_567             ( u0_col_out_567    ),
    .col_out_568             ( u0_col_out_568    ),
    .col_out_569             ( u0_col_out_569    ),
    .col_out_570             ( u0_col_out_570    ),
    .col_out_571             ( u0_col_out_571    ),
    .col_out_572             ( u0_col_out_572    ),
    .col_out_573             ( u0_col_out_573    ),
    .col_out_574             ( u0_col_out_574    ),
    .col_out_575             ( u0_col_out_575    ),
    .col_out_576             ( u0_col_out_576    ),
    .col_out_577             ( u0_col_out_577    ),
    .col_out_578             ( u0_col_out_578    ),
    .col_out_579             ( u0_col_out_579    ),
    .col_out_580             ( u0_col_out_580    ),
    .col_out_581             ( u0_col_out_581    ),
    .col_out_582             ( u0_col_out_582    ),
    .col_out_583             ( u0_col_out_583    ),
    .col_out_584             ( u0_col_out_584    ),
    .col_out_585             ( u0_col_out_585    ),
    .col_out_586             ( u0_col_out_586    ),
    .col_out_587             ( u0_col_out_587    ),
    .col_out_588             ( u0_col_out_588    ),
    .col_out_589             ( u0_col_out_589    ),
    .col_out_590             ( u0_col_out_590    ),
    .col_out_591             ( u0_col_out_591    ),
    .col_out_592             ( u0_col_out_592    ),
    .col_out_593             ( u0_col_out_593    ),
    .col_out_594             ( u0_col_out_594    ),
    .col_out_595             ( u0_col_out_595    ),
    .col_out_596             ( u0_col_out_596    ),
    .col_out_597             ( u0_col_out_597    ),
    .col_out_598             ( u0_col_out_598    ),
    .col_out_599             ( u0_col_out_599    ),
    .col_out_600             ( u0_col_out_600    ),
    .col_out_601             ( u0_col_out_601    ),
    .col_out_602             ( u0_col_out_602    ),
    .col_out_603             ( u0_col_out_603    ),
    .col_out_604             ( u0_col_out_604    ),
    .col_out_605             ( u0_col_out_605    ),
    .col_out_606             ( u0_col_out_606    ),
    .col_out_607             ( u0_col_out_607    ),
    .col_out_608             ( u0_col_out_608    ),
    .col_out_609             ( u0_col_out_609    ),
    .col_out_610             ( u0_col_out_610    ),
    .col_out_611             ( u0_col_out_611    ),
    .col_out_612             ( u0_col_out_612    ),
    .col_out_613             ( u0_col_out_613    ),
    .col_out_614             ( u0_col_out_614    ),
    .col_out_615             ( u0_col_out_615    ),
    .col_out_616             ( u0_col_out_616    ),
    .col_out_617             ( u0_col_out_617    ),
    .col_out_618             ( u0_col_out_618    ),
    .col_out_619             ( u0_col_out_619    ),
    .col_out_620             ( u0_col_out_620    ),
    .col_out_621             ( u0_col_out_621    ),
    .col_out_622             ( u0_col_out_622    ),
    .col_out_623             ( u0_col_out_623    ),
    .col_out_624             ( u0_col_out_624    ),
    .col_out_625             ( u0_col_out_625    ),
    .col_out_626             ( u0_col_out_626    ),
    .col_out_627             ( u0_col_out_627    ),
    .col_out_628             ( u0_col_out_628    ),
    .col_out_629             ( u0_col_out_629    ),
    .col_out_630             ( u0_col_out_630    ),
    .col_out_631             ( u0_col_out_631    ),
    .col_out_632             ( u0_col_out_632    ),
    .col_out_633             ( u0_col_out_633    ),
    .col_out_634             ( u0_col_out_634    ),
    .col_out_635             ( u0_col_out_635    ),
    .col_out_636             ( u0_col_out_636    ),
    .col_out_637             ( u0_col_out_637    ),
    .col_out_638             ( u0_col_out_638    ),
    .col_out_639             ( u0_col_out_639    ),
    .col_out_640             ( u0_col_out_640    ),
    .col_out_641             ( u0_col_out_641    ),
    .col_out_642             ( u0_col_out_642    ),
    .col_out_643             ( u0_col_out_643    ),
    .col_out_644             ( u0_col_out_644    ),
    .col_out_645             ( u0_col_out_645    ),
    .col_out_646             ( u0_col_out_646    ),
    .col_out_647             ( u0_col_out_647    ),
    .col_out_648             ( u0_col_out_648    ),
    .col_out_649             ( u0_col_out_649    ),
    .col_out_650             ( u0_col_out_650    ),
    .col_out_651             ( u0_col_out_651    ),
    .col_out_652             ( u0_col_out_652    ),
    .col_out_653             ( u0_col_out_653    ),
    .col_out_654             ( u0_col_out_654    ),
    .col_out_655             ( u0_col_out_655    ),
    .col_out_656             ( u0_col_out_656    ),
    .col_out_657             ( u0_col_out_657    ),
    .col_out_658             ( u0_col_out_658    ),
    .col_out_659             ( u0_col_out_659    ),
    .col_out_660             ( u0_col_out_660    ),
    .col_out_661             ( u0_col_out_661    ),
    .col_out_662             ( u0_col_out_662    ),
    .col_out_663             ( u0_col_out_663    ),
    .col_out_664             ( u0_col_out_664    ),
    .col_out_665             ( u0_col_out_665    ),
    .col_out_666             ( u0_col_out_666    ),
    .col_out_667             ( u0_col_out_667    ),
    .col_out_668             ( u0_col_out_668    ),
    .col_out_669             ( u0_col_out_669    ),
    .col_out_670             ( u0_col_out_670    ),
    .col_out_671             ( u0_col_out_671    ),
    .col_out_672             ( u0_col_out_672    ),
    .col_out_673             ( u0_col_out_673    ),
    .col_out_674             ( u0_col_out_674    ),
    .col_out_675             ( u0_col_out_675    ),
    .col_out_676             ( u0_col_out_676    ),
    .col_out_677             ( u0_col_out_677    ),
    .col_out_678             ( u0_col_out_678    ),
    .col_out_679             ( u0_col_out_679    ),
    .col_out_680             ( u0_col_out_680    ),
    .col_out_681             ( u0_col_out_681    ),
    .col_out_682             ( u0_col_out_682    ),
    .col_out_683             ( u0_col_out_683    ),
    .col_out_684             ( u0_col_out_684    ),
    .col_out_685             ( u0_col_out_685    ),
    .col_out_686             ( u0_col_out_686    ),
    .col_out_687             ( u0_col_out_687    ),
    .col_out_688             ( u0_col_out_688    ),
    .col_out_689             ( u0_col_out_689    ),
    .col_out_690             ( u0_col_out_690    ),
    .col_out_691             ( u0_col_out_691    ),
    .col_out_692             ( u0_col_out_692    ),
    .col_out_693             ( u0_col_out_693    ),
    .col_out_694             ( u0_col_out_694    ),
    .col_out_695             ( u0_col_out_695    ),
    .col_out_696             ( u0_col_out_696    ),
    .col_out_697             ( u0_col_out_697    ),
    .col_out_698             ( u0_col_out_698    ),
    .col_out_699             ( u0_col_out_699    ),
    .col_out_700             ( u0_col_out_700    ),
    .col_out_701             ( u0_col_out_701    ),
    .col_out_702             ( u0_col_out_702    ),
    .col_out_703             ( u0_col_out_703    ),
    .col_out_704             ( u0_col_out_704    ),
    .col_out_705             ( u0_col_out_705    ),
    .col_out_706             ( u0_col_out_706    ),
    .col_out_707             ( u0_col_out_707    ),
    .col_out_708             ( u0_col_out_708    ),
    .col_out_709             ( u0_col_out_709    ),
    .col_out_710             ( u0_col_out_710    ),
    .col_out_711             ( u0_col_out_711    ),
    .col_out_712             ( u0_col_out_712    ),
    .col_out_713             ( u0_col_out_713    ),
    .col_out_714             ( u0_col_out_714    ),
    .col_out_715             ( u0_col_out_715    ),
    .col_out_716             ( u0_col_out_716    ),
    .col_out_717             ( u0_col_out_717    ),
    .col_out_718             ( u0_col_out_718    ),
    .col_out_719             ( u0_col_out_719    ),
    .col_out_720             ( u0_col_out_720    ),
    .col_out_721             ( u0_col_out_721    ),
    .col_out_722             ( u0_col_out_722    ),
    .col_out_723             ( u0_col_out_723    ),
    .col_out_724             ( u0_col_out_724    ),
    .col_out_725             ( u0_col_out_725    ),
    .col_out_726             ( u0_col_out_726    ),
    .col_out_727             ( u0_col_out_727    ),
    .col_out_728             ( u0_col_out_728    ),
    .col_out_729             ( u0_col_out_729    ),
    .col_out_730             ( u0_col_out_730    ),
    .col_out_731             ( u0_col_out_731    ),
    .col_out_732             ( u0_col_out_732    ),
    .col_out_733             ( u0_col_out_733    ),
    .col_out_734             ( u0_col_out_734    ),
    .col_out_735             ( u0_col_out_735    ),
    .col_out_736             ( u0_col_out_736    ),
    .col_out_737             ( u0_col_out_737    ),
    .col_out_738             ( u0_col_out_738    ),
    .col_out_739             ( u0_col_out_739    ),
    .col_out_740             ( u0_col_out_740    ),
    .col_out_741             ( u0_col_out_741    ),
    .col_out_742             ( u0_col_out_742    ),
    .col_out_743             ( u0_col_out_743    ),
    .col_out_744             ( u0_col_out_744    ),
    .col_out_745             ( u0_col_out_745    ),
    .col_out_746             ( u0_col_out_746    ),
    .col_out_747             ( u0_col_out_747    ),
    .col_out_748             ( u0_col_out_748    ),
    .col_out_749             ( u0_col_out_749    ),
    .col_out_750             ( u0_col_out_750    ),
    .col_out_751             ( u0_col_out_751    ),
    .col_out_752             ( u0_col_out_752    ),
    .col_out_753             ( u0_col_out_753    ),
    .col_out_754             ( u0_col_out_754    ),
    .col_out_755             ( u0_col_out_755    ),
    .col_out_756             ( u0_col_out_756    ),
    .col_out_757             ( u0_col_out_757    ),
    .col_out_758             ( u0_col_out_758    ),
    .col_out_759             ( u0_col_out_759    ),
    .col_out_760             ( u0_col_out_760    ),
    .col_out_761             ( u0_col_out_761    ),
    .col_out_762             ( u0_col_out_762    ),
    .col_out_763             ( u0_col_out_763    ),
    .col_out_764             ( u0_col_out_764    ),
    .col_out_765             ( u0_col_out_765    ),
    .col_out_766             ( u0_col_out_766    ),
    .col_out_767             ( u0_col_out_767    ),
    .col_out_768             ( u0_col_out_768    ),
    .col_out_769             ( u0_col_out_769    ),
    .col_out_770             ( u0_col_out_770    ),
    .col_out_771             ( u0_col_out_771    ),
    .col_out_772             ( u0_col_out_772    ),
    .col_out_773             ( u0_col_out_773    ),
    .col_out_774             ( u0_col_out_774    ),
    .col_out_775             ( u0_col_out_775    ),
    .col_out_776             ( u0_col_out_776    ),
    .col_out_777             ( u0_col_out_777    ),
    .col_out_778             ( u0_col_out_778    ),
    .col_out_779             ( u0_col_out_779    ),
    .col_out_780             ( u0_col_out_780    ),
    .col_out_781             ( u0_col_out_781    ),
    .col_out_782             ( u0_col_out_782    ),
    .col_out_783             ( u0_col_out_783    ),
    .col_out_784             ( u0_col_out_784    ),
    .col_out_785             ( u0_col_out_785    ),
    .col_out_786             ( u0_col_out_786    ),
    .col_out_787             ( u0_col_out_787    ),
    .col_out_788             ( u0_col_out_788    ),
    .col_out_789             ( u0_col_out_789    ),
    .col_out_790             ( u0_col_out_790    ),
    .col_out_791             ( u0_col_out_791    ),
    .col_out_792             ( u0_col_out_792    ),
    .col_out_793             ( u0_col_out_793    ),
    .col_out_794             ( u0_col_out_794    ),
    .col_out_795             ( u0_col_out_795    ),
    .col_out_796             ( u0_col_out_796    ),
    .col_out_797             ( u0_col_out_797    ),
    .col_out_798             ( u0_col_out_798    ),
    .col_out_799             ( u0_col_out_799    ),
    .col_out_800             ( u0_col_out_800    ),
    .col_out_801             ( u0_col_out_801    ),
    .col_out_802             ( u0_col_out_802    ),
    .col_out_803             ( u0_col_out_803    ),
    .col_out_804             ( u0_col_out_804    ),
    .col_out_805             ( u0_col_out_805    ),
    .col_out_806             ( u0_col_out_806    ),
    .col_out_807             ( u0_col_out_807    ),
    .col_out_808             ( u0_col_out_808    ),
    .col_out_809             ( u0_col_out_809    ),
    .col_out_810             ( u0_col_out_810    ),
    .col_out_811             ( u0_col_out_811    ),
    .col_out_812             ( u0_col_out_812    ),
    .col_out_813             ( u0_col_out_813    ),
    .col_out_814             ( u0_col_out_814    ),
    .col_out_815             ( u0_col_out_815    ),
    .col_out_816             ( u0_col_out_816    ),
    .col_out_817             ( u0_col_out_817    ),
    .col_out_818             ( u0_col_out_818    ),
    .col_out_819             ( u0_col_out_819    ),
    .col_out_820             ( u0_col_out_820    ),
    .col_out_821             ( u0_col_out_821    ),
    .col_out_822             ( u0_col_out_822    ),
    .col_out_823             ( u0_col_out_823    ),
    .col_out_824             ( u0_col_out_824    ),
    .col_out_825             ( u0_col_out_825    ),
    .col_out_826             ( u0_col_out_826    ),
    .col_out_827             ( u0_col_out_827    ),
    .col_out_828             ( u0_col_out_828    ),
    .col_out_829             ( u0_col_out_829    ),
    .col_out_830             ( u0_col_out_830    ),
    .col_out_831             ( u0_col_out_831    ),
    .col_out_832             ( u0_col_out_832    ),
    .col_out_833             ( u0_col_out_833    ),
    .col_out_834             ( u0_col_out_834    ),
    .col_out_835             ( u0_col_out_835    ),
    .col_out_836             ( u0_col_out_836    ),
    .col_out_837             ( u0_col_out_837    ),
    .col_out_838             ( u0_col_out_838    ),
    .col_out_839             ( u0_col_out_839    ),
    .col_out_840             ( u0_col_out_840    ),
    .col_out_841             ( u0_col_out_841    ),
    .col_out_842             ( u0_col_out_842    ),
    .col_out_843             ( u0_col_out_843    ),
    .col_out_844             ( u0_col_out_844    ),
    .col_out_845             ( u0_col_out_845    ),
    .col_out_846             ( u0_col_out_846    ),
    .col_out_847             ( u0_col_out_847    ),
    .col_out_848             ( u0_col_out_848    ),
    .col_out_849             ( u0_col_out_849    ),
    .col_out_850             ( u0_col_out_850    ),
    .col_out_851             ( u0_col_out_851    ),
    .col_out_852             ( u0_col_out_852    ),
    .col_out_853             ( u0_col_out_853    ),
    .col_out_854             ( u0_col_out_854    ),
    .col_out_855             ( u0_col_out_855    ),
    .col_out_856             ( u0_col_out_856    ),
    .col_out_857             ( u0_col_out_857    ),
    .col_out_858             ( u0_col_out_858    ),
    .col_out_859             ( u0_col_out_859    ),
    .col_out_860             ( u0_col_out_860    ),
    .col_out_861             ( u0_col_out_861    ),
    .col_out_862             ( u0_col_out_862    ),
    .col_out_863             ( u0_col_out_863    ),
    .col_out_864             ( u0_col_out_864    ),
    .col_out_865             ( u0_col_out_865    ),
    .col_out_866             ( u0_col_out_866    ),
    .col_out_867             ( u0_col_out_867    ),
    .col_out_868             ( u0_col_out_868    ),
    .col_out_869             ( u0_col_out_869    ),
    .col_out_870             ( u0_col_out_870    ),
    .col_out_871             ( u0_col_out_871    ),
    .col_out_872             ( u0_col_out_872    ),
    .col_out_873             ( u0_col_out_873    ),
    .col_out_874             ( u0_col_out_874    ),
    .col_out_875             ( u0_col_out_875    ),
    .col_out_876             ( u0_col_out_876    ),
    .col_out_877             ( u0_col_out_877    ),
    .col_out_878             ( u0_col_out_878    ),
    .col_out_879             ( u0_col_out_879    ),
    .col_out_880             ( u0_col_out_880    ),
    .col_out_881             ( u0_col_out_881    ),
    .col_out_882             ( u0_col_out_882    ),
    .col_out_883             ( u0_col_out_883    ),
    .col_out_884             ( u0_col_out_884    ),
    .col_out_885             ( u0_col_out_885    ),
    .col_out_886             ( u0_col_out_886    ),
    .col_out_887             ( u0_col_out_887    ),
    .col_out_888             ( u0_col_out_888    ),
    .col_out_889             ( u0_col_out_889    ),
    .col_out_890             ( u0_col_out_890    ),
    .col_out_891             ( u0_col_out_891    ),
    .col_out_892             ( u0_col_out_892    ),
    .col_out_893             ( u0_col_out_893    ),
    .col_out_894             ( u0_col_out_894    ),
    .col_out_895             ( u0_col_out_895    ),
    .col_out_896             ( u0_col_out_896    ),
    .col_out_897             ( u0_col_out_897    ),
    .col_out_898             ( u0_col_out_898    ),
    .col_out_899             ( u0_col_out_899    ),
    .col_out_900             ( u0_col_out_900    ),
    .col_out_901             ( u0_col_out_901    ),
    .col_out_902             ( u0_col_out_902    ),
    .col_out_903             ( u0_col_out_903    ),
    .col_out_904             ( u0_col_out_904    ),
    .col_out_905             ( u0_col_out_905    ),
    .col_out_906             ( u0_col_out_906    ),
    .col_out_907             ( u0_col_out_907    ),
    .col_out_908             ( u0_col_out_908    ),
    .col_out_909             ( u0_col_out_909    ),
    .col_out_910             ( u0_col_out_910    ),
    .col_out_911             ( u0_col_out_911    ),
    .col_out_912             ( u0_col_out_912    ),
    .col_out_913             ( u0_col_out_913    ),
    .col_out_914             ( u0_col_out_914    ),
    .col_out_915             ( u0_col_out_915    ),
    .col_out_916             ( u0_col_out_916    ),
    .col_out_917             ( u0_col_out_917    ),
    .col_out_918             ( u0_col_out_918    ),
    .col_out_919             ( u0_col_out_919    ),
    .col_out_920             ( u0_col_out_920    ),
    .col_out_921             ( u0_col_out_921    ),
    .col_out_922             ( u0_col_out_922    ),
    .col_out_923             ( u0_col_out_923    ),
    .col_out_924             ( u0_col_out_924    ),
    .col_out_925             ( u0_col_out_925    ),
    .col_out_926             ( u0_col_out_926    ),
    .col_out_927             ( u0_col_out_927    ),
    .col_out_928             ( u0_col_out_928    ),
    .col_out_929             ( u0_col_out_929    ),
    .col_out_930             ( u0_col_out_930    ),
    .col_out_931             ( u0_col_out_931    ),
    .col_out_932             ( u0_col_out_932    ),
    .col_out_933             ( u0_col_out_933    ),
    .col_out_934             ( u0_col_out_934    ),
    .col_out_935             ( u0_col_out_935    ),
    .col_out_936             ( u0_col_out_936    ),
    .col_out_937             ( u0_col_out_937    ),
    .col_out_938             ( u0_col_out_938    ),
    .col_out_939             ( u0_col_out_939    ),
    .col_out_940             ( u0_col_out_940    ),
    .col_out_941             ( u0_col_out_941    ),
    .col_out_942             ( u0_col_out_942    ),
    .col_out_943             ( u0_col_out_943    ),
    .col_out_944             ( u0_col_out_944    ),
    .col_out_945             ( u0_col_out_945    ),
    .col_out_946             ( u0_col_out_946    ),
    .col_out_947             ( u0_col_out_947    ),
    .col_out_948             ( u0_col_out_948    ),
    .col_out_949             ( u0_col_out_949    ),
    .col_out_950             ( u0_col_out_950    ),
    .col_out_951             ( u0_col_out_951    ),
    .col_out_952             ( u0_col_out_952    ),
    .col_out_953             ( u0_col_out_953    ),
    .col_out_954             ( u0_col_out_954    ),
    .col_out_955             ( u0_col_out_955    ),
    .col_out_956             ( u0_col_out_956    ),
    .col_out_957             ( u0_col_out_957    ),
    .col_out_958             ( u0_col_out_958    ),
    .col_out_959             ( u0_col_out_959    ),
    .col_out_960             ( u0_col_out_960    ),
    .col_out_961             ( u0_col_out_961    ),
    .col_out_962             ( u0_col_out_962    ),
    .col_out_963             ( u0_col_out_963    ),
    .col_out_964             ( u0_col_out_964    ),
    .col_out_965             ( u0_col_out_965    ),
    .col_out_966             ( u0_col_out_966    ),
    .col_out_967             ( u0_col_out_967    ),
    .col_out_968             ( u0_col_out_968    ),
    .col_out_969             ( u0_col_out_969    ),
    .col_out_970             ( u0_col_out_970    ),
    .col_out_971             ( u0_col_out_971    ),
    .col_out_972             ( u0_col_out_972    ),
    .col_out_973             ( u0_col_out_973    ),
    .col_out_974             ( u0_col_out_974    ),
    .col_out_975             ( u0_col_out_975    ),
    .col_out_976             ( u0_col_out_976    ),
    .col_out_977             ( u0_col_out_977    ),
    .col_out_978             ( u0_col_out_978    ),
    .col_out_979             ( u0_col_out_979    ),
    .col_out_980             ( u0_col_out_980    ),
    .col_out_981             ( u0_col_out_981    ),
    .col_out_982             ( u0_col_out_982    ),
    .col_out_983             ( u0_col_out_983    ),
    .col_out_984             ( u0_col_out_984    ),
    .col_out_985             ( u0_col_out_985    ),
    .col_out_986             ( u0_col_out_986    ),
    .col_out_987             ( u0_col_out_987    ),
    .col_out_988             ( u0_col_out_988    ),
    .col_out_989             ( u0_col_out_989    ),
    .col_out_990             ( u0_col_out_990    ),
    .col_out_991             ( u0_col_out_991    ),
    .col_out_992             ( u0_col_out_992    ),
    .col_out_993             ( u0_col_out_993    ),
    .col_out_994             ( u0_col_out_994    ),
    .col_out_995             ( u0_col_out_995    ),
    .col_out_996             ( u0_col_out_996    ),
    .col_out_997             ( u0_col_out_997    ),
    .col_out_998             ( u0_col_out_998    ),
    .col_out_999             ( u0_col_out_999    ),
    .col_out_1000            ( u0_col_out_1000   ),
    .col_out_1001            ( u0_col_out_1001   ),
    .col_out_1002            ( u0_col_out_1002   ),
    .col_out_1003            ( u0_col_out_1003   ),
    .col_out_1004            ( u0_col_out_1004   ),
    .col_out_1005            ( u0_col_out_1005   ),
    .col_out_1006            ( u0_col_out_1006   ),
    .col_out_1007            ( u0_col_out_1007   ),
    .col_out_1008            ( u0_col_out_1008   ),
    .col_out_1009            ( u0_col_out_1009   ),
    .col_out_1010            ( u0_col_out_1010   ),
    .col_out_1011            ( u0_col_out_1011   ),
    .col_out_1012            ( u0_col_out_1012   ),
    .col_out_1013            ( u0_col_out_1013   ),
    .col_out_1014            ( u0_col_out_1014   ),
    .col_out_1015            ( u0_col_out_1015   ),
    .col_out_1016            ( u0_col_out_1016   ),
    .col_out_1017            ( u0_col_out_1017   ),
    .col_out_1018            ( u0_col_out_1018   ),
    .col_out_1019            ( u0_col_out_1019   ),
    .col_out_1020            ( u0_col_out_1020   ),
    .col_out_1021            ( u0_col_out_1021   ),
    .col_out_1022            ( u0_col_out_1022   ),
    .col_out_1023            ( u0_col_out_1023   ),
    .col_out_1024            ( u0_col_out_1024   ),
    .col_out_1025            ( u0_col_out_1025   ),
    .col_out_1026            ( u0_col_out_1026   ),
    .col_out_1027            ( u0_col_out_1027   ),
    .col_out_1028            ( u0_col_out_1028   ),
    .col_out_1029            ( u0_col_out_1029   ),
    .col_out_1030            ( u0_col_out_1030   ),
    .col_out_1031            ( u0_col_out_1031   ),
    .col_out_1032            ( u0_col_out_1032   ),
    .col_out_1033            ( u0_col_out_1033   )
);
















// compressor_array_12_8_1033 Outputs
wire  [7:0]  u1_col_out_0;
wire  [7:0]  u1_col_out_1;
wire  [7:0]  u1_col_out_2;
wire  [7:0]  u1_col_out_3;
wire  [7:0]  u1_col_out_4;
wire  [7:0]  u1_col_out_5;
wire  [7:0]  u1_col_out_6;
wire  [7:0]  u1_col_out_7;
wire  [7:0]  u1_col_out_8;
wire  [7:0]  u1_col_out_9;
wire  [7:0]  u1_col_out_10;
wire  [7:0]  u1_col_out_11;
wire  [7:0]  u1_col_out_12;
wire  [7:0]  u1_col_out_13;
wire  [7:0]  u1_col_out_14;
wire  [7:0]  u1_col_out_15;
wire  [7:0]  u1_col_out_16;
wire  [7:0]  u1_col_out_17;
wire  [7:0]  u1_col_out_18;
wire  [7:0]  u1_col_out_19;
wire  [7:0]  u1_col_out_20;
wire  [7:0]  u1_col_out_21;
wire  [7:0]  u1_col_out_22;
wire  [7:0]  u1_col_out_23;
wire  [7:0]  u1_col_out_24;
wire  [7:0]  u1_col_out_25;
wire  [7:0]  u1_col_out_26;
wire  [7:0]  u1_col_out_27;
wire  [7:0]  u1_col_out_28;
wire  [7:0]  u1_col_out_29;
wire  [7:0]  u1_col_out_30;
wire  [7:0]  u1_col_out_31;
wire  [7:0]  u1_col_out_32;
wire  [7:0]  u1_col_out_33;
wire  [7:0]  u1_col_out_34;
wire  [7:0]  u1_col_out_35;
wire  [7:0]  u1_col_out_36;
wire  [7:0]  u1_col_out_37;
wire  [7:0]  u1_col_out_38;
wire  [7:0]  u1_col_out_39;
wire  [7:0]  u1_col_out_40;
wire  [7:0]  u1_col_out_41;
wire  [7:0]  u1_col_out_42;
wire  [7:0]  u1_col_out_43;
wire  [7:0]  u1_col_out_44;
wire  [7:0]  u1_col_out_45;
wire  [7:0]  u1_col_out_46;
wire  [7:0]  u1_col_out_47;
wire  [7:0]  u1_col_out_48;
wire  [7:0]  u1_col_out_49;
wire  [7:0]  u1_col_out_50;
wire  [7:0]  u1_col_out_51;
wire  [7:0]  u1_col_out_52;
wire  [7:0]  u1_col_out_53;
wire  [7:0]  u1_col_out_54;
wire  [7:0]  u1_col_out_55;
wire  [7:0]  u1_col_out_56;
wire  [7:0]  u1_col_out_57;
wire  [7:0]  u1_col_out_58;
wire  [7:0]  u1_col_out_59;
wire  [7:0]  u1_col_out_60;
wire  [7:0]  u1_col_out_61;
wire  [7:0]  u1_col_out_62;
wire  [7:0]  u1_col_out_63;
wire  [7:0]  u1_col_out_64;
wire  [7:0]  u1_col_out_65;
wire  [7:0]  u1_col_out_66;
wire  [7:0]  u1_col_out_67;
wire  [7:0]  u1_col_out_68;
wire  [7:0]  u1_col_out_69;
wire  [7:0]  u1_col_out_70;
wire  [7:0]  u1_col_out_71;
wire  [7:0]  u1_col_out_72;
wire  [7:0]  u1_col_out_73;
wire  [7:0]  u1_col_out_74;
wire  [7:0]  u1_col_out_75;
wire  [7:0]  u1_col_out_76;
wire  [7:0]  u1_col_out_77;
wire  [7:0]  u1_col_out_78;
wire  [7:0]  u1_col_out_79;
wire  [7:0]  u1_col_out_80;
wire  [7:0]  u1_col_out_81;
wire  [7:0]  u1_col_out_82;
wire  [7:0]  u1_col_out_83;
wire  [7:0]  u1_col_out_84;
wire  [7:0]  u1_col_out_85;
wire  [7:0]  u1_col_out_86;
wire  [7:0]  u1_col_out_87;
wire  [7:0]  u1_col_out_88;
wire  [7:0]  u1_col_out_89;
wire  [7:0]  u1_col_out_90;
wire  [7:0]  u1_col_out_91;
wire  [7:0]  u1_col_out_92;
wire  [7:0]  u1_col_out_93;
wire  [7:0]  u1_col_out_94;
wire  [7:0]  u1_col_out_95;
wire  [7:0]  u1_col_out_96;
wire  [7:0]  u1_col_out_97;
wire  [7:0]  u1_col_out_98;
wire  [7:0]  u1_col_out_99;
wire  [7:0]  u1_col_out_100;
wire  [7:0]  u1_col_out_101;
wire  [7:0]  u1_col_out_102;
wire  [7:0]  u1_col_out_103;
wire  [7:0]  u1_col_out_104;
wire  [7:0]  u1_col_out_105;
wire  [7:0]  u1_col_out_106;
wire  [7:0]  u1_col_out_107;
wire  [7:0]  u1_col_out_108;
wire  [7:0]  u1_col_out_109;
wire  [7:0]  u1_col_out_110;
wire  [7:0]  u1_col_out_111;
wire  [7:0]  u1_col_out_112;
wire  [7:0]  u1_col_out_113;
wire  [7:0]  u1_col_out_114;
wire  [7:0]  u1_col_out_115;
wire  [7:0]  u1_col_out_116;
wire  [7:0]  u1_col_out_117;
wire  [7:0]  u1_col_out_118;
wire  [7:0]  u1_col_out_119;
wire  [7:0]  u1_col_out_120;
wire  [7:0]  u1_col_out_121;
wire  [7:0]  u1_col_out_122;
wire  [7:0]  u1_col_out_123;
wire  [7:0]  u1_col_out_124;
wire  [7:0]  u1_col_out_125;
wire  [7:0]  u1_col_out_126;
wire  [7:0]  u1_col_out_127;
wire  [7:0]  u1_col_out_128;
wire  [7:0]  u1_col_out_129;
wire  [7:0]  u1_col_out_130;
wire  [7:0]  u1_col_out_131;
wire  [7:0]  u1_col_out_132;
wire  [7:0]  u1_col_out_133;
wire  [7:0]  u1_col_out_134;
wire  [7:0]  u1_col_out_135;
wire  [7:0]  u1_col_out_136;
wire  [7:0]  u1_col_out_137;
wire  [7:0]  u1_col_out_138;
wire  [7:0]  u1_col_out_139;
wire  [7:0]  u1_col_out_140;
wire  [7:0]  u1_col_out_141;
wire  [7:0]  u1_col_out_142;
wire  [7:0]  u1_col_out_143;
wire  [7:0]  u1_col_out_144;
wire  [7:0]  u1_col_out_145;
wire  [7:0]  u1_col_out_146;
wire  [7:0]  u1_col_out_147;
wire  [7:0]  u1_col_out_148;
wire  [7:0]  u1_col_out_149;
wire  [7:0]  u1_col_out_150;
wire  [7:0]  u1_col_out_151;
wire  [7:0]  u1_col_out_152;
wire  [7:0]  u1_col_out_153;
wire  [7:0]  u1_col_out_154;
wire  [7:0]  u1_col_out_155;
wire  [7:0]  u1_col_out_156;
wire  [7:0]  u1_col_out_157;
wire  [7:0]  u1_col_out_158;
wire  [7:0]  u1_col_out_159;
wire  [7:0]  u1_col_out_160;
wire  [7:0]  u1_col_out_161;
wire  [7:0]  u1_col_out_162;
wire  [7:0]  u1_col_out_163;
wire  [7:0]  u1_col_out_164;
wire  [7:0]  u1_col_out_165;
wire  [7:0]  u1_col_out_166;
wire  [7:0]  u1_col_out_167;
wire  [7:0]  u1_col_out_168;
wire  [7:0]  u1_col_out_169;
wire  [7:0]  u1_col_out_170;
wire  [7:0]  u1_col_out_171;
wire  [7:0]  u1_col_out_172;
wire  [7:0]  u1_col_out_173;
wire  [7:0]  u1_col_out_174;
wire  [7:0]  u1_col_out_175;
wire  [7:0]  u1_col_out_176;
wire  [7:0]  u1_col_out_177;
wire  [7:0]  u1_col_out_178;
wire  [7:0]  u1_col_out_179;
wire  [7:0]  u1_col_out_180;
wire  [7:0]  u1_col_out_181;
wire  [7:0]  u1_col_out_182;
wire  [7:0]  u1_col_out_183;
wire  [7:0]  u1_col_out_184;
wire  [7:0]  u1_col_out_185;
wire  [7:0]  u1_col_out_186;
wire  [7:0]  u1_col_out_187;
wire  [7:0]  u1_col_out_188;
wire  [7:0]  u1_col_out_189;
wire  [7:0]  u1_col_out_190;
wire  [7:0]  u1_col_out_191;
wire  [7:0]  u1_col_out_192;
wire  [7:0]  u1_col_out_193;
wire  [7:0]  u1_col_out_194;
wire  [7:0]  u1_col_out_195;
wire  [7:0]  u1_col_out_196;
wire  [7:0]  u1_col_out_197;
wire  [7:0]  u1_col_out_198;
wire  [7:0]  u1_col_out_199;
wire  [7:0]  u1_col_out_200;
wire  [7:0]  u1_col_out_201;
wire  [7:0]  u1_col_out_202;
wire  [7:0]  u1_col_out_203;
wire  [7:0]  u1_col_out_204;
wire  [7:0]  u1_col_out_205;
wire  [7:0]  u1_col_out_206;
wire  [7:0]  u1_col_out_207;
wire  [7:0]  u1_col_out_208;
wire  [7:0]  u1_col_out_209;
wire  [7:0]  u1_col_out_210;
wire  [7:0]  u1_col_out_211;
wire  [7:0]  u1_col_out_212;
wire  [7:0]  u1_col_out_213;
wire  [7:0]  u1_col_out_214;
wire  [7:0]  u1_col_out_215;
wire  [7:0]  u1_col_out_216;
wire  [7:0]  u1_col_out_217;
wire  [7:0]  u1_col_out_218;
wire  [7:0]  u1_col_out_219;
wire  [7:0]  u1_col_out_220;
wire  [7:0]  u1_col_out_221;
wire  [7:0]  u1_col_out_222;
wire  [7:0]  u1_col_out_223;
wire  [7:0]  u1_col_out_224;
wire  [7:0]  u1_col_out_225;
wire  [7:0]  u1_col_out_226;
wire  [7:0]  u1_col_out_227;
wire  [7:0]  u1_col_out_228;
wire  [7:0]  u1_col_out_229;
wire  [7:0]  u1_col_out_230;
wire  [7:0]  u1_col_out_231;
wire  [7:0]  u1_col_out_232;
wire  [7:0]  u1_col_out_233;
wire  [7:0]  u1_col_out_234;
wire  [7:0]  u1_col_out_235;
wire  [7:0]  u1_col_out_236;
wire  [7:0]  u1_col_out_237;
wire  [7:0]  u1_col_out_238;
wire  [7:0]  u1_col_out_239;
wire  [7:0]  u1_col_out_240;
wire  [7:0]  u1_col_out_241;
wire  [7:0]  u1_col_out_242;
wire  [7:0]  u1_col_out_243;
wire  [7:0]  u1_col_out_244;
wire  [7:0]  u1_col_out_245;
wire  [7:0]  u1_col_out_246;
wire  [7:0]  u1_col_out_247;
wire  [7:0]  u1_col_out_248;
wire  [7:0]  u1_col_out_249;
wire  [7:0]  u1_col_out_250;
wire  [7:0]  u1_col_out_251;
wire  [7:0]  u1_col_out_252;
wire  [7:0]  u1_col_out_253;
wire  [7:0]  u1_col_out_254;
wire  [7:0]  u1_col_out_255;
wire  [7:0]  u1_col_out_256;
wire  [7:0]  u1_col_out_257;
wire  [7:0]  u1_col_out_258;
wire  [7:0]  u1_col_out_259;
wire  [7:0]  u1_col_out_260;
wire  [7:0]  u1_col_out_261;
wire  [7:0]  u1_col_out_262;
wire  [7:0]  u1_col_out_263;
wire  [7:0]  u1_col_out_264;
wire  [7:0]  u1_col_out_265;
wire  [7:0]  u1_col_out_266;
wire  [7:0]  u1_col_out_267;
wire  [7:0]  u1_col_out_268;
wire  [7:0]  u1_col_out_269;
wire  [7:0]  u1_col_out_270;
wire  [7:0]  u1_col_out_271;
wire  [7:0]  u1_col_out_272;
wire  [7:0]  u1_col_out_273;
wire  [7:0]  u1_col_out_274;
wire  [7:0]  u1_col_out_275;
wire  [7:0]  u1_col_out_276;
wire  [7:0]  u1_col_out_277;
wire  [7:0]  u1_col_out_278;
wire  [7:0]  u1_col_out_279;
wire  [7:0]  u1_col_out_280;
wire  [7:0]  u1_col_out_281;
wire  [7:0]  u1_col_out_282;
wire  [7:0]  u1_col_out_283;
wire  [7:0]  u1_col_out_284;
wire  [7:0]  u1_col_out_285;
wire  [7:0]  u1_col_out_286;
wire  [7:0]  u1_col_out_287;
wire  [7:0]  u1_col_out_288;
wire  [7:0]  u1_col_out_289;
wire  [7:0]  u1_col_out_290;
wire  [7:0]  u1_col_out_291;
wire  [7:0]  u1_col_out_292;
wire  [7:0]  u1_col_out_293;
wire  [7:0]  u1_col_out_294;
wire  [7:0]  u1_col_out_295;
wire  [7:0]  u1_col_out_296;
wire  [7:0]  u1_col_out_297;
wire  [7:0]  u1_col_out_298;
wire  [7:0]  u1_col_out_299;
wire  [7:0]  u1_col_out_300;
wire  [7:0]  u1_col_out_301;
wire  [7:0]  u1_col_out_302;
wire  [7:0]  u1_col_out_303;
wire  [7:0]  u1_col_out_304;
wire  [7:0]  u1_col_out_305;
wire  [7:0]  u1_col_out_306;
wire  [7:0]  u1_col_out_307;
wire  [7:0]  u1_col_out_308;
wire  [7:0]  u1_col_out_309;
wire  [7:0]  u1_col_out_310;
wire  [7:0]  u1_col_out_311;
wire  [7:0]  u1_col_out_312;
wire  [7:0]  u1_col_out_313;
wire  [7:0]  u1_col_out_314;
wire  [7:0]  u1_col_out_315;
wire  [7:0]  u1_col_out_316;
wire  [7:0]  u1_col_out_317;
wire  [7:0]  u1_col_out_318;
wire  [7:0]  u1_col_out_319;
wire  [7:0]  u1_col_out_320;
wire  [7:0]  u1_col_out_321;
wire  [7:0]  u1_col_out_322;
wire  [7:0]  u1_col_out_323;
wire  [7:0]  u1_col_out_324;
wire  [7:0]  u1_col_out_325;
wire  [7:0]  u1_col_out_326;
wire  [7:0]  u1_col_out_327;
wire  [7:0]  u1_col_out_328;
wire  [7:0]  u1_col_out_329;
wire  [7:0]  u1_col_out_330;
wire  [7:0]  u1_col_out_331;
wire  [7:0]  u1_col_out_332;
wire  [7:0]  u1_col_out_333;
wire  [7:0]  u1_col_out_334;
wire  [7:0]  u1_col_out_335;
wire  [7:0]  u1_col_out_336;
wire  [7:0]  u1_col_out_337;
wire  [7:0]  u1_col_out_338;
wire  [7:0]  u1_col_out_339;
wire  [7:0]  u1_col_out_340;
wire  [7:0]  u1_col_out_341;
wire  [7:0]  u1_col_out_342;
wire  [7:0]  u1_col_out_343;
wire  [7:0]  u1_col_out_344;
wire  [7:0]  u1_col_out_345;
wire  [7:0]  u1_col_out_346;
wire  [7:0]  u1_col_out_347;
wire  [7:0]  u1_col_out_348;
wire  [7:0]  u1_col_out_349;
wire  [7:0]  u1_col_out_350;
wire  [7:0]  u1_col_out_351;
wire  [7:0]  u1_col_out_352;
wire  [7:0]  u1_col_out_353;
wire  [7:0]  u1_col_out_354;
wire  [7:0]  u1_col_out_355;
wire  [7:0]  u1_col_out_356;
wire  [7:0]  u1_col_out_357;
wire  [7:0]  u1_col_out_358;
wire  [7:0]  u1_col_out_359;
wire  [7:0]  u1_col_out_360;
wire  [7:0]  u1_col_out_361;
wire  [7:0]  u1_col_out_362;
wire  [7:0]  u1_col_out_363;
wire  [7:0]  u1_col_out_364;
wire  [7:0]  u1_col_out_365;
wire  [7:0]  u1_col_out_366;
wire  [7:0]  u1_col_out_367;
wire  [7:0]  u1_col_out_368;
wire  [7:0]  u1_col_out_369;
wire  [7:0]  u1_col_out_370;
wire  [7:0]  u1_col_out_371;
wire  [7:0]  u1_col_out_372;
wire  [7:0]  u1_col_out_373;
wire  [7:0]  u1_col_out_374;
wire  [7:0]  u1_col_out_375;
wire  [7:0]  u1_col_out_376;
wire  [7:0]  u1_col_out_377;
wire  [7:0]  u1_col_out_378;
wire  [7:0]  u1_col_out_379;
wire  [7:0]  u1_col_out_380;
wire  [7:0]  u1_col_out_381;
wire  [7:0]  u1_col_out_382;
wire  [7:0]  u1_col_out_383;
wire  [7:0]  u1_col_out_384;
wire  [7:0]  u1_col_out_385;
wire  [7:0]  u1_col_out_386;
wire  [7:0]  u1_col_out_387;
wire  [7:0]  u1_col_out_388;
wire  [7:0]  u1_col_out_389;
wire  [7:0]  u1_col_out_390;
wire  [7:0]  u1_col_out_391;
wire  [7:0]  u1_col_out_392;
wire  [7:0]  u1_col_out_393;
wire  [7:0]  u1_col_out_394;
wire  [7:0]  u1_col_out_395;
wire  [7:0]  u1_col_out_396;
wire  [7:0]  u1_col_out_397;
wire  [7:0]  u1_col_out_398;
wire  [7:0]  u1_col_out_399;
wire  [7:0]  u1_col_out_400;
wire  [7:0]  u1_col_out_401;
wire  [7:0]  u1_col_out_402;
wire  [7:0]  u1_col_out_403;
wire  [7:0]  u1_col_out_404;
wire  [7:0]  u1_col_out_405;
wire  [7:0]  u1_col_out_406;
wire  [7:0]  u1_col_out_407;
wire  [7:0]  u1_col_out_408;
wire  [7:0]  u1_col_out_409;
wire  [7:0]  u1_col_out_410;
wire  [7:0]  u1_col_out_411;
wire  [7:0]  u1_col_out_412;
wire  [7:0]  u1_col_out_413;
wire  [7:0]  u1_col_out_414;
wire  [7:0]  u1_col_out_415;
wire  [7:0]  u1_col_out_416;
wire  [7:0]  u1_col_out_417;
wire  [7:0]  u1_col_out_418;
wire  [7:0]  u1_col_out_419;
wire  [7:0]  u1_col_out_420;
wire  [7:0]  u1_col_out_421;
wire  [7:0]  u1_col_out_422;
wire  [7:0]  u1_col_out_423;
wire  [7:0]  u1_col_out_424;
wire  [7:0]  u1_col_out_425;
wire  [7:0]  u1_col_out_426;
wire  [7:0]  u1_col_out_427;
wire  [7:0]  u1_col_out_428;
wire  [7:0]  u1_col_out_429;
wire  [7:0]  u1_col_out_430;
wire  [7:0]  u1_col_out_431;
wire  [7:0]  u1_col_out_432;
wire  [7:0]  u1_col_out_433;
wire  [7:0]  u1_col_out_434;
wire  [7:0]  u1_col_out_435;
wire  [7:0]  u1_col_out_436;
wire  [7:0]  u1_col_out_437;
wire  [7:0]  u1_col_out_438;
wire  [7:0]  u1_col_out_439;
wire  [7:0]  u1_col_out_440;
wire  [7:0]  u1_col_out_441;
wire  [7:0]  u1_col_out_442;
wire  [7:0]  u1_col_out_443;
wire  [7:0]  u1_col_out_444;
wire  [7:0]  u1_col_out_445;
wire  [7:0]  u1_col_out_446;
wire  [7:0]  u1_col_out_447;
wire  [7:0]  u1_col_out_448;
wire  [7:0]  u1_col_out_449;
wire  [7:0]  u1_col_out_450;
wire  [7:0]  u1_col_out_451;
wire  [7:0]  u1_col_out_452;
wire  [7:0]  u1_col_out_453;
wire  [7:0]  u1_col_out_454;
wire  [7:0]  u1_col_out_455;
wire  [7:0]  u1_col_out_456;
wire  [7:0]  u1_col_out_457;
wire  [7:0]  u1_col_out_458;
wire  [7:0]  u1_col_out_459;
wire  [7:0]  u1_col_out_460;
wire  [7:0]  u1_col_out_461;
wire  [7:0]  u1_col_out_462;
wire  [7:0]  u1_col_out_463;
wire  [7:0]  u1_col_out_464;
wire  [7:0]  u1_col_out_465;
wire  [7:0]  u1_col_out_466;
wire  [7:0]  u1_col_out_467;
wire  [7:0]  u1_col_out_468;
wire  [7:0]  u1_col_out_469;
wire  [7:0]  u1_col_out_470;
wire  [7:0]  u1_col_out_471;
wire  [7:0]  u1_col_out_472;
wire  [7:0]  u1_col_out_473;
wire  [7:0]  u1_col_out_474;
wire  [7:0]  u1_col_out_475;
wire  [7:0]  u1_col_out_476;
wire  [7:0]  u1_col_out_477;
wire  [7:0]  u1_col_out_478;
wire  [7:0]  u1_col_out_479;
wire  [7:0]  u1_col_out_480;
wire  [7:0]  u1_col_out_481;
wire  [7:0]  u1_col_out_482;
wire  [7:0]  u1_col_out_483;
wire  [7:0]  u1_col_out_484;
wire  [7:0]  u1_col_out_485;
wire  [7:0]  u1_col_out_486;
wire  [7:0]  u1_col_out_487;
wire  [7:0]  u1_col_out_488;
wire  [7:0]  u1_col_out_489;
wire  [7:0]  u1_col_out_490;
wire  [7:0]  u1_col_out_491;
wire  [7:0]  u1_col_out_492;
wire  [7:0]  u1_col_out_493;
wire  [7:0]  u1_col_out_494;
wire  [7:0]  u1_col_out_495;
wire  [7:0]  u1_col_out_496;
wire  [7:0]  u1_col_out_497;
wire  [7:0]  u1_col_out_498;
wire  [7:0]  u1_col_out_499;
wire  [7:0]  u1_col_out_500;
wire  [7:0]  u1_col_out_501;
wire  [7:0]  u1_col_out_502;
wire  [7:0]  u1_col_out_503;
wire  [7:0]  u1_col_out_504;
wire  [7:0]  u1_col_out_505;
wire  [7:0]  u1_col_out_506;
wire  [7:0]  u1_col_out_507;
wire  [7:0]  u1_col_out_508;
wire  [7:0]  u1_col_out_509;
wire  [7:0]  u1_col_out_510;
wire  [7:0]  u1_col_out_511;
wire  [7:0]  u1_col_out_512;
wire  [7:0]  u1_col_out_513;
wire  [7:0]  u1_col_out_514;
wire  [7:0]  u1_col_out_515;
wire  [7:0]  u1_col_out_516;
wire  [7:0]  u1_col_out_517;
wire  [7:0]  u1_col_out_518;
wire  [7:0]  u1_col_out_519;
wire  [7:0]  u1_col_out_520;
wire  [7:0]  u1_col_out_521;
wire  [7:0]  u1_col_out_522;
wire  [7:0]  u1_col_out_523;
wire  [7:0]  u1_col_out_524;
wire  [7:0]  u1_col_out_525;
wire  [7:0]  u1_col_out_526;
wire  [7:0]  u1_col_out_527;
wire  [7:0]  u1_col_out_528;
wire  [7:0]  u1_col_out_529;
wire  [7:0]  u1_col_out_530;
wire  [7:0]  u1_col_out_531;
wire  [7:0]  u1_col_out_532;
wire  [7:0]  u1_col_out_533;
wire  [7:0]  u1_col_out_534;
wire  [7:0]  u1_col_out_535;
wire  [7:0]  u1_col_out_536;
wire  [7:0]  u1_col_out_537;
wire  [7:0]  u1_col_out_538;
wire  [7:0]  u1_col_out_539;
wire  [7:0]  u1_col_out_540;
wire  [7:0]  u1_col_out_541;
wire  [7:0]  u1_col_out_542;
wire  [7:0]  u1_col_out_543;
wire  [7:0]  u1_col_out_544;
wire  [7:0]  u1_col_out_545;
wire  [7:0]  u1_col_out_546;
wire  [7:0]  u1_col_out_547;
wire  [7:0]  u1_col_out_548;
wire  [7:0]  u1_col_out_549;
wire  [7:0]  u1_col_out_550;
wire  [7:0]  u1_col_out_551;
wire  [7:0]  u1_col_out_552;
wire  [7:0]  u1_col_out_553;
wire  [7:0]  u1_col_out_554;
wire  [7:0]  u1_col_out_555;
wire  [7:0]  u1_col_out_556;
wire  [7:0]  u1_col_out_557;
wire  [7:0]  u1_col_out_558;
wire  [7:0]  u1_col_out_559;
wire  [7:0]  u1_col_out_560;
wire  [7:0]  u1_col_out_561;
wire  [7:0]  u1_col_out_562;
wire  [7:0]  u1_col_out_563;
wire  [7:0]  u1_col_out_564;
wire  [7:0]  u1_col_out_565;
wire  [7:0]  u1_col_out_566;
wire  [7:0]  u1_col_out_567;
wire  [7:0]  u1_col_out_568;
wire  [7:0]  u1_col_out_569;
wire  [7:0]  u1_col_out_570;
wire  [7:0]  u1_col_out_571;
wire  [7:0]  u1_col_out_572;
wire  [7:0]  u1_col_out_573;
wire  [7:0]  u1_col_out_574;
wire  [7:0]  u1_col_out_575;
wire  [7:0]  u1_col_out_576;
wire  [7:0]  u1_col_out_577;
wire  [7:0]  u1_col_out_578;
wire  [7:0]  u1_col_out_579;
wire  [7:0]  u1_col_out_580;
wire  [7:0]  u1_col_out_581;
wire  [7:0]  u1_col_out_582;
wire  [7:0]  u1_col_out_583;
wire  [7:0]  u1_col_out_584;
wire  [7:0]  u1_col_out_585;
wire  [7:0]  u1_col_out_586;
wire  [7:0]  u1_col_out_587;
wire  [7:0]  u1_col_out_588;
wire  [7:0]  u1_col_out_589;
wire  [7:0]  u1_col_out_590;
wire  [7:0]  u1_col_out_591;
wire  [7:0]  u1_col_out_592;
wire  [7:0]  u1_col_out_593;
wire  [7:0]  u1_col_out_594;
wire  [7:0]  u1_col_out_595;
wire  [7:0]  u1_col_out_596;
wire  [7:0]  u1_col_out_597;
wire  [7:0]  u1_col_out_598;
wire  [7:0]  u1_col_out_599;
wire  [7:0]  u1_col_out_600;
wire  [7:0]  u1_col_out_601;
wire  [7:0]  u1_col_out_602;
wire  [7:0]  u1_col_out_603;
wire  [7:0]  u1_col_out_604;
wire  [7:0]  u1_col_out_605;
wire  [7:0]  u1_col_out_606;
wire  [7:0]  u1_col_out_607;
wire  [7:0]  u1_col_out_608;
wire  [7:0]  u1_col_out_609;
wire  [7:0]  u1_col_out_610;
wire  [7:0]  u1_col_out_611;
wire  [7:0]  u1_col_out_612;
wire  [7:0]  u1_col_out_613;
wire  [7:0]  u1_col_out_614;
wire  [7:0]  u1_col_out_615;
wire  [7:0]  u1_col_out_616;
wire  [7:0]  u1_col_out_617;
wire  [7:0]  u1_col_out_618;
wire  [7:0]  u1_col_out_619;
wire  [7:0]  u1_col_out_620;
wire  [7:0]  u1_col_out_621;
wire  [7:0]  u1_col_out_622;
wire  [7:0]  u1_col_out_623;
wire  [7:0]  u1_col_out_624;
wire  [7:0]  u1_col_out_625;
wire  [7:0]  u1_col_out_626;
wire  [7:0]  u1_col_out_627;
wire  [7:0]  u1_col_out_628;
wire  [7:0]  u1_col_out_629;
wire  [7:0]  u1_col_out_630;
wire  [7:0]  u1_col_out_631;
wire  [7:0]  u1_col_out_632;
wire  [7:0]  u1_col_out_633;
wire  [7:0]  u1_col_out_634;
wire  [7:0]  u1_col_out_635;
wire  [7:0]  u1_col_out_636;
wire  [7:0]  u1_col_out_637;
wire  [7:0]  u1_col_out_638;
wire  [7:0]  u1_col_out_639;
wire  [7:0]  u1_col_out_640;
wire  [7:0]  u1_col_out_641;
wire  [7:0]  u1_col_out_642;
wire  [7:0]  u1_col_out_643;
wire  [7:0]  u1_col_out_644;
wire  [7:0]  u1_col_out_645;
wire  [7:0]  u1_col_out_646;
wire  [7:0]  u1_col_out_647;
wire  [7:0]  u1_col_out_648;
wire  [7:0]  u1_col_out_649;
wire  [7:0]  u1_col_out_650;
wire  [7:0]  u1_col_out_651;
wire  [7:0]  u1_col_out_652;
wire  [7:0]  u1_col_out_653;
wire  [7:0]  u1_col_out_654;
wire  [7:0]  u1_col_out_655;
wire  [7:0]  u1_col_out_656;
wire  [7:0]  u1_col_out_657;
wire  [7:0]  u1_col_out_658;
wire  [7:0]  u1_col_out_659;
wire  [7:0]  u1_col_out_660;
wire  [7:0]  u1_col_out_661;
wire  [7:0]  u1_col_out_662;
wire  [7:0]  u1_col_out_663;
wire  [7:0]  u1_col_out_664;
wire  [7:0]  u1_col_out_665;
wire  [7:0]  u1_col_out_666;
wire  [7:0]  u1_col_out_667;
wire  [7:0]  u1_col_out_668;
wire  [7:0]  u1_col_out_669;
wire  [7:0]  u1_col_out_670;
wire  [7:0]  u1_col_out_671;
wire  [7:0]  u1_col_out_672;
wire  [7:0]  u1_col_out_673;
wire  [7:0]  u1_col_out_674;
wire  [7:0]  u1_col_out_675;
wire  [7:0]  u1_col_out_676;
wire  [7:0]  u1_col_out_677;
wire  [7:0]  u1_col_out_678;
wire  [7:0]  u1_col_out_679;
wire  [7:0]  u1_col_out_680;
wire  [7:0]  u1_col_out_681;
wire  [7:0]  u1_col_out_682;
wire  [7:0]  u1_col_out_683;
wire  [7:0]  u1_col_out_684;
wire  [7:0]  u1_col_out_685;
wire  [7:0]  u1_col_out_686;
wire  [7:0]  u1_col_out_687;
wire  [7:0]  u1_col_out_688;
wire  [7:0]  u1_col_out_689;
wire  [7:0]  u1_col_out_690;
wire  [7:0]  u1_col_out_691;
wire  [7:0]  u1_col_out_692;
wire  [7:0]  u1_col_out_693;
wire  [7:0]  u1_col_out_694;
wire  [7:0]  u1_col_out_695;
wire  [7:0]  u1_col_out_696;
wire  [7:0]  u1_col_out_697;
wire  [7:0]  u1_col_out_698;
wire  [7:0]  u1_col_out_699;
wire  [7:0]  u1_col_out_700;
wire  [7:0]  u1_col_out_701;
wire  [7:0]  u1_col_out_702;
wire  [7:0]  u1_col_out_703;
wire  [7:0]  u1_col_out_704;
wire  [7:0]  u1_col_out_705;
wire  [7:0]  u1_col_out_706;
wire  [7:0]  u1_col_out_707;
wire  [7:0]  u1_col_out_708;
wire  [7:0]  u1_col_out_709;
wire  [7:0]  u1_col_out_710;
wire  [7:0]  u1_col_out_711;
wire  [7:0]  u1_col_out_712;
wire  [7:0]  u1_col_out_713;
wire  [7:0]  u1_col_out_714;
wire  [7:0]  u1_col_out_715;
wire  [7:0]  u1_col_out_716;
wire  [7:0]  u1_col_out_717;
wire  [7:0]  u1_col_out_718;
wire  [7:0]  u1_col_out_719;
wire  [7:0]  u1_col_out_720;
wire  [7:0]  u1_col_out_721;
wire  [7:0]  u1_col_out_722;
wire  [7:0]  u1_col_out_723;
wire  [7:0]  u1_col_out_724;
wire  [7:0]  u1_col_out_725;
wire  [7:0]  u1_col_out_726;
wire  [7:0]  u1_col_out_727;
wire  [7:0]  u1_col_out_728;
wire  [7:0]  u1_col_out_729;
wire  [7:0]  u1_col_out_730;
wire  [7:0]  u1_col_out_731;
wire  [7:0]  u1_col_out_732;
wire  [7:0]  u1_col_out_733;
wire  [7:0]  u1_col_out_734;
wire  [7:0]  u1_col_out_735;
wire  [7:0]  u1_col_out_736;
wire  [7:0]  u1_col_out_737;
wire  [7:0]  u1_col_out_738;
wire  [7:0]  u1_col_out_739;
wire  [7:0]  u1_col_out_740;
wire  [7:0]  u1_col_out_741;
wire  [7:0]  u1_col_out_742;
wire  [7:0]  u1_col_out_743;
wire  [7:0]  u1_col_out_744;
wire  [7:0]  u1_col_out_745;
wire  [7:0]  u1_col_out_746;
wire  [7:0]  u1_col_out_747;
wire  [7:0]  u1_col_out_748;
wire  [7:0]  u1_col_out_749;
wire  [7:0]  u1_col_out_750;
wire  [7:0]  u1_col_out_751;
wire  [7:0]  u1_col_out_752;
wire  [7:0]  u1_col_out_753;
wire  [7:0]  u1_col_out_754;
wire  [7:0]  u1_col_out_755;
wire  [7:0]  u1_col_out_756;
wire  [7:0]  u1_col_out_757;
wire  [7:0]  u1_col_out_758;
wire  [7:0]  u1_col_out_759;
wire  [7:0]  u1_col_out_760;
wire  [7:0]  u1_col_out_761;
wire  [7:0]  u1_col_out_762;
wire  [7:0]  u1_col_out_763;
wire  [7:0]  u1_col_out_764;
wire  [7:0]  u1_col_out_765;
wire  [7:0]  u1_col_out_766;
wire  [7:0]  u1_col_out_767;
wire  [7:0]  u1_col_out_768;
wire  [7:0]  u1_col_out_769;
wire  [7:0]  u1_col_out_770;
wire  [7:0]  u1_col_out_771;
wire  [7:0]  u1_col_out_772;
wire  [7:0]  u1_col_out_773;
wire  [7:0]  u1_col_out_774;
wire  [7:0]  u1_col_out_775;
wire  [7:0]  u1_col_out_776;
wire  [7:0]  u1_col_out_777;
wire  [7:0]  u1_col_out_778;
wire  [7:0]  u1_col_out_779;
wire  [7:0]  u1_col_out_780;
wire  [7:0]  u1_col_out_781;
wire  [7:0]  u1_col_out_782;
wire  [7:0]  u1_col_out_783;
wire  [7:0]  u1_col_out_784;
wire  [7:0]  u1_col_out_785;
wire  [7:0]  u1_col_out_786;
wire  [7:0]  u1_col_out_787;
wire  [7:0]  u1_col_out_788;
wire  [7:0]  u1_col_out_789;
wire  [7:0]  u1_col_out_790;
wire  [7:0]  u1_col_out_791;
wire  [7:0]  u1_col_out_792;
wire  [7:0]  u1_col_out_793;
wire  [7:0]  u1_col_out_794;
wire  [7:0]  u1_col_out_795;
wire  [7:0]  u1_col_out_796;
wire  [7:0]  u1_col_out_797;
wire  [7:0]  u1_col_out_798;
wire  [7:0]  u1_col_out_799;
wire  [7:0]  u1_col_out_800;
wire  [7:0]  u1_col_out_801;
wire  [7:0]  u1_col_out_802;
wire  [7:0]  u1_col_out_803;
wire  [7:0]  u1_col_out_804;
wire  [7:0]  u1_col_out_805;
wire  [7:0]  u1_col_out_806;
wire  [7:0]  u1_col_out_807;
wire  [7:0]  u1_col_out_808;
wire  [7:0]  u1_col_out_809;
wire  [7:0]  u1_col_out_810;
wire  [7:0]  u1_col_out_811;
wire  [7:0]  u1_col_out_812;
wire  [7:0]  u1_col_out_813;
wire  [7:0]  u1_col_out_814;
wire  [7:0]  u1_col_out_815;
wire  [7:0]  u1_col_out_816;
wire  [7:0]  u1_col_out_817;
wire  [7:0]  u1_col_out_818;
wire  [7:0]  u1_col_out_819;
wire  [7:0]  u1_col_out_820;
wire  [7:0]  u1_col_out_821;
wire  [7:0]  u1_col_out_822;
wire  [7:0]  u1_col_out_823;
wire  [7:0]  u1_col_out_824;
wire  [7:0]  u1_col_out_825;
wire  [7:0]  u1_col_out_826;
wire  [7:0]  u1_col_out_827;
wire  [7:0]  u1_col_out_828;
wire  [7:0]  u1_col_out_829;
wire  [7:0]  u1_col_out_830;
wire  [7:0]  u1_col_out_831;
wire  [7:0]  u1_col_out_832;
wire  [7:0]  u1_col_out_833;
wire  [7:0]  u1_col_out_834;
wire  [7:0]  u1_col_out_835;
wire  [7:0]  u1_col_out_836;
wire  [7:0]  u1_col_out_837;
wire  [7:0]  u1_col_out_838;
wire  [7:0]  u1_col_out_839;
wire  [7:0]  u1_col_out_840;
wire  [7:0]  u1_col_out_841;
wire  [7:0]  u1_col_out_842;
wire  [7:0]  u1_col_out_843;
wire  [7:0]  u1_col_out_844;
wire  [7:0]  u1_col_out_845;
wire  [7:0]  u1_col_out_846;
wire  [7:0]  u1_col_out_847;
wire  [7:0]  u1_col_out_848;
wire  [7:0]  u1_col_out_849;
wire  [7:0]  u1_col_out_850;
wire  [7:0]  u1_col_out_851;
wire  [7:0]  u1_col_out_852;
wire  [7:0]  u1_col_out_853;
wire  [7:0]  u1_col_out_854;
wire  [7:0]  u1_col_out_855;
wire  [7:0]  u1_col_out_856;
wire  [7:0]  u1_col_out_857;
wire  [7:0]  u1_col_out_858;
wire  [7:0]  u1_col_out_859;
wire  [7:0]  u1_col_out_860;
wire  [7:0]  u1_col_out_861;
wire  [7:0]  u1_col_out_862;
wire  [7:0]  u1_col_out_863;
wire  [7:0]  u1_col_out_864;
wire  [7:0]  u1_col_out_865;
wire  [7:0]  u1_col_out_866;
wire  [7:0]  u1_col_out_867;
wire  [7:0]  u1_col_out_868;
wire  [7:0]  u1_col_out_869;
wire  [7:0]  u1_col_out_870;
wire  [7:0]  u1_col_out_871;
wire  [7:0]  u1_col_out_872;
wire  [7:0]  u1_col_out_873;
wire  [7:0]  u1_col_out_874;
wire  [7:0]  u1_col_out_875;
wire  [7:0]  u1_col_out_876;
wire  [7:0]  u1_col_out_877;
wire  [7:0]  u1_col_out_878;
wire  [7:0]  u1_col_out_879;
wire  [7:0]  u1_col_out_880;
wire  [7:0]  u1_col_out_881;
wire  [7:0]  u1_col_out_882;
wire  [7:0]  u1_col_out_883;
wire  [7:0]  u1_col_out_884;
wire  [7:0]  u1_col_out_885;
wire  [7:0]  u1_col_out_886;
wire  [7:0]  u1_col_out_887;
wire  [7:0]  u1_col_out_888;
wire  [7:0]  u1_col_out_889;
wire  [7:0]  u1_col_out_890;
wire  [7:0]  u1_col_out_891;
wire  [7:0]  u1_col_out_892;
wire  [7:0]  u1_col_out_893;
wire  [7:0]  u1_col_out_894;
wire  [7:0]  u1_col_out_895;
wire  [7:0]  u1_col_out_896;
wire  [7:0]  u1_col_out_897;
wire  [7:0]  u1_col_out_898;
wire  [7:0]  u1_col_out_899;
wire  [7:0]  u1_col_out_900;
wire  [7:0]  u1_col_out_901;
wire  [7:0]  u1_col_out_902;
wire  [7:0]  u1_col_out_903;
wire  [7:0]  u1_col_out_904;
wire  [7:0]  u1_col_out_905;
wire  [7:0]  u1_col_out_906;
wire  [7:0]  u1_col_out_907;
wire  [7:0]  u1_col_out_908;
wire  [7:0]  u1_col_out_909;
wire  [7:0]  u1_col_out_910;
wire  [7:0]  u1_col_out_911;
wire  [7:0]  u1_col_out_912;
wire  [7:0]  u1_col_out_913;
wire  [7:0]  u1_col_out_914;
wire  [7:0]  u1_col_out_915;
wire  [7:0]  u1_col_out_916;
wire  [7:0]  u1_col_out_917;
wire  [7:0]  u1_col_out_918;
wire  [7:0]  u1_col_out_919;
wire  [7:0]  u1_col_out_920;
wire  [7:0]  u1_col_out_921;
wire  [7:0]  u1_col_out_922;
wire  [7:0]  u1_col_out_923;
wire  [7:0]  u1_col_out_924;
wire  [7:0]  u1_col_out_925;
wire  [7:0]  u1_col_out_926;
wire  [7:0]  u1_col_out_927;
wire  [7:0]  u1_col_out_928;
wire  [7:0]  u1_col_out_929;
wire  [7:0]  u1_col_out_930;
wire  [7:0]  u1_col_out_931;
wire  [7:0]  u1_col_out_932;
wire  [7:0]  u1_col_out_933;
wire  [7:0]  u1_col_out_934;
wire  [7:0]  u1_col_out_935;
wire  [7:0]  u1_col_out_936;
wire  [7:0]  u1_col_out_937;
wire  [7:0]  u1_col_out_938;
wire  [7:0]  u1_col_out_939;
wire  [7:0]  u1_col_out_940;
wire  [7:0]  u1_col_out_941;
wire  [7:0]  u1_col_out_942;
wire  [7:0]  u1_col_out_943;
wire  [7:0]  u1_col_out_944;
wire  [7:0]  u1_col_out_945;
wire  [7:0]  u1_col_out_946;
wire  [7:0]  u1_col_out_947;
wire  [7:0]  u1_col_out_948;
wire  [7:0]  u1_col_out_949;
wire  [7:0]  u1_col_out_950;
wire  [7:0]  u1_col_out_951;
wire  [7:0]  u1_col_out_952;
wire  [7:0]  u1_col_out_953;
wire  [7:0]  u1_col_out_954;
wire  [7:0]  u1_col_out_955;
wire  [7:0]  u1_col_out_956;
wire  [7:0]  u1_col_out_957;
wire  [7:0]  u1_col_out_958;
wire  [7:0]  u1_col_out_959;
wire  [7:0]  u1_col_out_960;
wire  [7:0]  u1_col_out_961;
wire  [7:0]  u1_col_out_962;
wire  [7:0]  u1_col_out_963;
wire  [7:0]  u1_col_out_964;
wire  [7:0]  u1_col_out_965;
wire  [7:0]  u1_col_out_966;
wire  [7:0]  u1_col_out_967;
wire  [7:0]  u1_col_out_968;
wire  [7:0]  u1_col_out_969;
wire  [7:0]  u1_col_out_970;
wire  [7:0]  u1_col_out_971;
wire  [7:0]  u1_col_out_972;
wire  [7:0]  u1_col_out_973;
wire  [7:0]  u1_col_out_974;
wire  [7:0]  u1_col_out_975;
wire  [7:0]  u1_col_out_976;
wire  [7:0]  u1_col_out_977;
wire  [7:0]  u1_col_out_978;
wire  [7:0]  u1_col_out_979;
wire  [7:0]  u1_col_out_980;
wire  [7:0]  u1_col_out_981;
wire  [7:0]  u1_col_out_982;
wire  [7:0]  u1_col_out_983;
wire  [7:0]  u1_col_out_984;
wire  [7:0]  u1_col_out_985;
wire  [7:0]  u1_col_out_986;
wire  [7:0]  u1_col_out_987;
wire  [7:0]  u1_col_out_988;
wire  [7:0]  u1_col_out_989;
wire  [7:0]  u1_col_out_990;
wire  [7:0]  u1_col_out_991;
wire  [7:0]  u1_col_out_992;
wire  [7:0]  u1_col_out_993;
wire  [7:0]  u1_col_out_994;
wire  [7:0]  u1_col_out_995;
wire  [7:0]  u1_col_out_996;
wire  [7:0]  u1_col_out_997;
wire  [7:0]  u1_col_out_998;
wire  [7:0]  u1_col_out_999;
wire  [7:0]  u1_col_out_1000;
wire  [7:0]  u1_col_out_1001;
wire  [7:0]  u1_col_out_1002;
wire  [7:0]  u1_col_out_1003;
wire  [7:0]  u1_col_out_1004;
wire  [7:0]  u1_col_out_1005;
wire  [7:0]  u1_col_out_1006;
wire  [7:0]  u1_col_out_1007;
wire  [7:0]  u1_col_out_1008;
wire  [7:0]  u1_col_out_1009;
wire  [7:0]  u1_col_out_1010;
wire  [7:0]  u1_col_out_1011;
wire  [7:0]  u1_col_out_1012;
wire  [7:0]  u1_col_out_1013;
wire  [7:0]  u1_col_out_1014;
wire  [7:0]  u1_col_out_1015;
wire  [7:0]  u1_col_out_1016;
wire  [7:0]  u1_col_out_1017;
wire  [7:0]  u1_col_out_1018;
wire  [7:0]  u1_col_out_1019;
wire  [7:0]  u1_col_out_1020;
wire  [7:0]  u1_col_out_1021;
wire  [7:0]  u1_col_out_1022;
wire  [7:0]  u1_col_out_1023;
wire  [7:0]  u1_col_out_1024;
wire  [7:0]  u1_col_out_1025;
wire  [7:0]  u1_col_out_1026;
wire  [7:0]  u1_col_out_1027;
wire  [7:0]  u1_col_out_1028;
wire  [7:0]  u1_col_out_1029;
wire  [7:0]  u1_col_out_1030;
wire  [7:0]  u1_col_out_1031;
wire  [7:0]  u1_col_out_1032;
wire  [7:0]  u1_col_out_1033;

compressor_array_12_8_1033  u1_compressor_array_12_8_1033 (
    .col_in_0                ( u0_col_out_0       ),
    .col_in_1                ( u0_col_out_1       ),
    .col_in_2                ( u0_col_out_2       ),
    .col_in_3                ( u0_col_out_3       ),
    .col_in_4                ( u0_col_out_4       ),
    .col_in_5                ( u0_col_out_5       ),
    .col_in_6                ( u0_col_out_6       ),
    .col_in_7                ( u0_col_out_7       ),
    .col_in_8                ( u0_col_out_8       ),
    .col_in_9                ( u0_col_out_9       ),
    .col_in_10               ( u0_col_out_10      ),
    .col_in_11               ( u0_col_out_11      ),
    .col_in_12               ( u0_col_out_12      ),
    .col_in_13               ( u0_col_out_13      ),
    .col_in_14               ( u0_col_out_14      ),
    .col_in_15               ( u0_col_out_15      ),
    .col_in_16               ( u0_col_out_16      ),
    .col_in_17               ( u0_col_out_17      ),
    .col_in_18               ( u0_col_out_18      ),
    .col_in_19               ( u0_col_out_19      ),
    .col_in_20               ( u0_col_out_20      ),
    .col_in_21               ( u0_col_out_21      ),
    .col_in_22               ( u0_col_out_22      ),
    .col_in_23               ( u0_col_out_23      ),
    .col_in_24               ( u0_col_out_24      ),
    .col_in_25               ( u0_col_out_25      ),
    .col_in_26               ( u0_col_out_26      ),
    .col_in_27               ( u0_col_out_27      ),
    .col_in_28               ( u0_col_out_28      ),
    .col_in_29               ( u0_col_out_29      ),
    .col_in_30               ( u0_col_out_30      ),
    .col_in_31               ( u0_col_out_31      ),
    .col_in_32               ( u0_col_out_32      ),
    .col_in_33               ( u0_col_out_33      ),
    .col_in_34               ( u0_col_out_34      ),
    .col_in_35               ( u0_col_out_35      ),
    .col_in_36               ( u0_col_out_36      ),
    .col_in_37               ( u0_col_out_37      ),
    .col_in_38               ( u0_col_out_38      ),
    .col_in_39               ( u0_col_out_39      ),
    .col_in_40               ( u0_col_out_40      ),
    .col_in_41               ( u0_col_out_41      ),
    .col_in_42               ( u0_col_out_42      ),
    .col_in_43               ( u0_col_out_43      ),
    .col_in_44               ( u0_col_out_44      ),
    .col_in_45               ( u0_col_out_45      ),
    .col_in_46               ( u0_col_out_46      ),
    .col_in_47               ( u0_col_out_47      ),
    .col_in_48               ( u0_col_out_48      ),
    .col_in_49               ( u0_col_out_49      ),
    .col_in_50               ( u0_col_out_50      ),
    .col_in_51               ( u0_col_out_51      ),
    .col_in_52               ( u0_col_out_52      ),
    .col_in_53               ( u0_col_out_53      ),
    .col_in_54               ( u0_col_out_54      ),
    .col_in_55               ( u0_col_out_55      ),
    .col_in_56               ( u0_col_out_56      ),
    .col_in_57               ( u0_col_out_57      ),
    .col_in_58               ( u0_col_out_58      ),
    .col_in_59               ( u0_col_out_59      ),
    .col_in_60               ( u0_col_out_60      ),
    .col_in_61               ( u0_col_out_61      ),
    .col_in_62               ( u0_col_out_62      ),
    .col_in_63               ( u0_col_out_63      ),
    .col_in_64               ( u0_col_out_64      ),
    .col_in_65               ( u0_col_out_65      ),
    .col_in_66               ( u0_col_out_66      ),
    .col_in_67               ( u0_col_out_67      ),
    .col_in_68               ( u0_col_out_68      ),
    .col_in_69               ( u0_col_out_69      ),
    .col_in_70               ( u0_col_out_70      ),
    .col_in_71               ( u0_col_out_71      ),
    .col_in_72               ( u0_col_out_72      ),
    .col_in_73               ( u0_col_out_73      ),
    .col_in_74               ( u0_col_out_74      ),
    .col_in_75               ( u0_col_out_75      ),
    .col_in_76               ( u0_col_out_76      ),
    .col_in_77               ( u0_col_out_77      ),
    .col_in_78               ( u0_col_out_78      ),
    .col_in_79               ( u0_col_out_79      ),
    .col_in_80               ( u0_col_out_80      ),
    .col_in_81               ( u0_col_out_81      ),
    .col_in_82               ( u0_col_out_82      ),
    .col_in_83               ( u0_col_out_83      ),
    .col_in_84               ( u0_col_out_84      ),
    .col_in_85               ( u0_col_out_85      ),
    .col_in_86               ( u0_col_out_86      ),
    .col_in_87               ( u0_col_out_87      ),
    .col_in_88               ( u0_col_out_88      ),
    .col_in_89               ( u0_col_out_89      ),
    .col_in_90               ( u0_col_out_90      ),
    .col_in_91               ( u0_col_out_91      ),
    .col_in_92               ( u0_col_out_92      ),
    .col_in_93               ( u0_col_out_93      ),
    .col_in_94               ( u0_col_out_94      ),
    .col_in_95               ( u0_col_out_95      ),
    .col_in_96               ( u0_col_out_96      ),
    .col_in_97               ( u0_col_out_97      ),
    .col_in_98               ( u0_col_out_98      ),
    .col_in_99               ( u0_col_out_99      ),
    .col_in_100              ( u0_col_out_100     ),
    .col_in_101              ( u0_col_out_101     ),
    .col_in_102              ( u0_col_out_102     ),
    .col_in_103              ( u0_col_out_103     ),
    .col_in_104              ( u0_col_out_104     ),
    .col_in_105              ( u0_col_out_105     ),
    .col_in_106              ( u0_col_out_106     ),
    .col_in_107              ( u0_col_out_107     ),
    .col_in_108              ( u0_col_out_108     ),
    .col_in_109              ( u0_col_out_109     ),
    .col_in_110              ( u0_col_out_110     ),
    .col_in_111              ( u0_col_out_111     ),
    .col_in_112              ( u0_col_out_112     ),
    .col_in_113              ( u0_col_out_113     ),
    .col_in_114              ( u0_col_out_114     ),
    .col_in_115              ( u0_col_out_115     ),
    .col_in_116              ( u0_col_out_116     ),
    .col_in_117              ( u0_col_out_117     ),
    .col_in_118              ( u0_col_out_118     ),
    .col_in_119              ( u0_col_out_119     ),
    .col_in_120              ( u0_col_out_120     ),
    .col_in_121              ( u0_col_out_121     ),
    .col_in_122              ( u0_col_out_122     ),
    .col_in_123              ( u0_col_out_123     ),
    .col_in_124              ( u0_col_out_124     ),
    .col_in_125              ( u0_col_out_125     ),
    .col_in_126              ( u0_col_out_126     ),
    .col_in_127              ( u0_col_out_127     ),
    .col_in_128              ( u0_col_out_128     ),
    .col_in_129              ( u0_col_out_129     ),
    .col_in_130              ( u0_col_out_130     ),
    .col_in_131              ( u0_col_out_131     ),
    .col_in_132              ( u0_col_out_132     ),
    .col_in_133              ( u0_col_out_133     ),
    .col_in_134              ( u0_col_out_134     ),
    .col_in_135              ( u0_col_out_135     ),
    .col_in_136              ( u0_col_out_136     ),
    .col_in_137              ( u0_col_out_137     ),
    .col_in_138              ( u0_col_out_138     ),
    .col_in_139              ( u0_col_out_139     ),
    .col_in_140              ( u0_col_out_140     ),
    .col_in_141              ( u0_col_out_141     ),
    .col_in_142              ( u0_col_out_142     ),
    .col_in_143              ( u0_col_out_143     ),
    .col_in_144              ( u0_col_out_144     ),
    .col_in_145              ( u0_col_out_145     ),
    .col_in_146              ( u0_col_out_146     ),
    .col_in_147              ( u0_col_out_147     ),
    .col_in_148              ( u0_col_out_148     ),
    .col_in_149              ( u0_col_out_149     ),
    .col_in_150              ( u0_col_out_150     ),
    .col_in_151              ( u0_col_out_151     ),
    .col_in_152              ( u0_col_out_152     ),
    .col_in_153              ( u0_col_out_153     ),
    .col_in_154              ( u0_col_out_154     ),
    .col_in_155              ( u0_col_out_155     ),
    .col_in_156              ( u0_col_out_156     ),
    .col_in_157              ( u0_col_out_157     ),
    .col_in_158              ( u0_col_out_158     ),
    .col_in_159              ( u0_col_out_159     ),
    .col_in_160              ( u0_col_out_160     ),
    .col_in_161              ( u0_col_out_161     ),
    .col_in_162              ( u0_col_out_162     ),
    .col_in_163              ( u0_col_out_163     ),
    .col_in_164              ( u0_col_out_164     ),
    .col_in_165              ( u0_col_out_165     ),
    .col_in_166              ( u0_col_out_166     ),
    .col_in_167              ( u0_col_out_167     ),
    .col_in_168              ( u0_col_out_168     ),
    .col_in_169              ( u0_col_out_169     ),
    .col_in_170              ( u0_col_out_170     ),
    .col_in_171              ( u0_col_out_171     ),
    .col_in_172              ( u0_col_out_172     ),
    .col_in_173              ( u0_col_out_173     ),
    .col_in_174              ( u0_col_out_174     ),
    .col_in_175              ( u0_col_out_175     ),
    .col_in_176              ( u0_col_out_176     ),
    .col_in_177              ( u0_col_out_177     ),
    .col_in_178              ( u0_col_out_178     ),
    .col_in_179              ( u0_col_out_179     ),
    .col_in_180              ( u0_col_out_180     ),
    .col_in_181              ( u0_col_out_181     ),
    .col_in_182              ( u0_col_out_182     ),
    .col_in_183              ( u0_col_out_183     ),
    .col_in_184              ( u0_col_out_184     ),
    .col_in_185              ( u0_col_out_185     ),
    .col_in_186              ( u0_col_out_186     ),
    .col_in_187              ( u0_col_out_187     ),
    .col_in_188              ( u0_col_out_188     ),
    .col_in_189              ( u0_col_out_189     ),
    .col_in_190              ( u0_col_out_190     ),
    .col_in_191              ( u0_col_out_191     ),
    .col_in_192              ( u0_col_out_192     ),
    .col_in_193              ( u0_col_out_193     ),
    .col_in_194              ( u0_col_out_194     ),
    .col_in_195              ( u0_col_out_195     ),
    .col_in_196              ( u0_col_out_196     ),
    .col_in_197              ( u0_col_out_197     ),
    .col_in_198              ( u0_col_out_198     ),
    .col_in_199              ( u0_col_out_199     ),
    .col_in_200              ( u0_col_out_200     ),
    .col_in_201              ( u0_col_out_201     ),
    .col_in_202              ( u0_col_out_202     ),
    .col_in_203              ( u0_col_out_203     ),
    .col_in_204              ( u0_col_out_204     ),
    .col_in_205              ( u0_col_out_205     ),
    .col_in_206              ( u0_col_out_206     ),
    .col_in_207              ( u0_col_out_207     ),
    .col_in_208              ( u0_col_out_208     ),
    .col_in_209              ( u0_col_out_209     ),
    .col_in_210              ( u0_col_out_210     ),
    .col_in_211              ( u0_col_out_211     ),
    .col_in_212              ( u0_col_out_212     ),
    .col_in_213              ( u0_col_out_213     ),
    .col_in_214              ( u0_col_out_214     ),
    .col_in_215              ( u0_col_out_215     ),
    .col_in_216              ( u0_col_out_216     ),
    .col_in_217              ( u0_col_out_217     ),
    .col_in_218              ( u0_col_out_218     ),
    .col_in_219              ( u0_col_out_219     ),
    .col_in_220              ( u0_col_out_220     ),
    .col_in_221              ( u0_col_out_221     ),
    .col_in_222              ( u0_col_out_222     ),
    .col_in_223              ( u0_col_out_223     ),
    .col_in_224              ( u0_col_out_224     ),
    .col_in_225              ( u0_col_out_225     ),
    .col_in_226              ( u0_col_out_226     ),
    .col_in_227              ( u0_col_out_227     ),
    .col_in_228              ( u0_col_out_228     ),
    .col_in_229              ( u0_col_out_229     ),
    .col_in_230              ( u0_col_out_230     ),
    .col_in_231              ( u0_col_out_231     ),
    .col_in_232              ( u0_col_out_232     ),
    .col_in_233              ( u0_col_out_233     ),
    .col_in_234              ( u0_col_out_234     ),
    .col_in_235              ( u0_col_out_235     ),
    .col_in_236              ( u0_col_out_236     ),
    .col_in_237              ( u0_col_out_237     ),
    .col_in_238              ( u0_col_out_238     ),
    .col_in_239              ( u0_col_out_239     ),
    .col_in_240              ( u0_col_out_240     ),
    .col_in_241              ( u0_col_out_241     ),
    .col_in_242              ( u0_col_out_242     ),
    .col_in_243              ( u0_col_out_243     ),
    .col_in_244              ( u0_col_out_244     ),
    .col_in_245              ( u0_col_out_245     ),
    .col_in_246              ( u0_col_out_246     ),
    .col_in_247              ( u0_col_out_247     ),
    .col_in_248              ( u0_col_out_248     ),
    .col_in_249              ( u0_col_out_249     ),
    .col_in_250              ( u0_col_out_250     ),
    .col_in_251              ( u0_col_out_251     ),
    .col_in_252              ( u0_col_out_252     ),
    .col_in_253              ( u0_col_out_253     ),
    .col_in_254              ( u0_col_out_254     ),
    .col_in_255              ( u0_col_out_255     ),
    .col_in_256              ( u0_col_out_256     ),
    .col_in_257              ( u0_col_out_257     ),
    .col_in_258              ( u0_col_out_258     ),
    .col_in_259              ( u0_col_out_259     ),
    .col_in_260              ( u0_col_out_260     ),
    .col_in_261              ( u0_col_out_261     ),
    .col_in_262              ( u0_col_out_262     ),
    .col_in_263              ( u0_col_out_263     ),
    .col_in_264              ( u0_col_out_264     ),
    .col_in_265              ( u0_col_out_265     ),
    .col_in_266              ( u0_col_out_266     ),
    .col_in_267              ( u0_col_out_267     ),
    .col_in_268              ( u0_col_out_268     ),
    .col_in_269              ( u0_col_out_269     ),
    .col_in_270              ( u0_col_out_270     ),
    .col_in_271              ( u0_col_out_271     ),
    .col_in_272              ( u0_col_out_272     ),
    .col_in_273              ( u0_col_out_273     ),
    .col_in_274              ( u0_col_out_274     ),
    .col_in_275              ( u0_col_out_275     ),
    .col_in_276              ( u0_col_out_276     ),
    .col_in_277              ( u0_col_out_277     ),
    .col_in_278              ( u0_col_out_278     ),
    .col_in_279              ( u0_col_out_279     ),
    .col_in_280              ( u0_col_out_280     ),
    .col_in_281              ( u0_col_out_281     ),
    .col_in_282              ( u0_col_out_282     ),
    .col_in_283              ( u0_col_out_283     ),
    .col_in_284              ( u0_col_out_284     ),
    .col_in_285              ( u0_col_out_285     ),
    .col_in_286              ( u0_col_out_286     ),
    .col_in_287              ( u0_col_out_287     ),
    .col_in_288              ( u0_col_out_288     ),
    .col_in_289              ( u0_col_out_289     ),
    .col_in_290              ( u0_col_out_290     ),
    .col_in_291              ( u0_col_out_291     ),
    .col_in_292              ( u0_col_out_292     ),
    .col_in_293              ( u0_col_out_293     ),
    .col_in_294              ( u0_col_out_294     ),
    .col_in_295              ( u0_col_out_295     ),
    .col_in_296              ( u0_col_out_296     ),
    .col_in_297              ( u0_col_out_297     ),
    .col_in_298              ( u0_col_out_298     ),
    .col_in_299              ( u0_col_out_299     ),
    .col_in_300              ( u0_col_out_300     ),
    .col_in_301              ( u0_col_out_301     ),
    .col_in_302              ( u0_col_out_302     ),
    .col_in_303              ( u0_col_out_303     ),
    .col_in_304              ( u0_col_out_304     ),
    .col_in_305              ( u0_col_out_305     ),
    .col_in_306              ( u0_col_out_306     ),
    .col_in_307              ( u0_col_out_307     ),
    .col_in_308              ( u0_col_out_308     ),
    .col_in_309              ( u0_col_out_309     ),
    .col_in_310              ( u0_col_out_310     ),
    .col_in_311              ( u0_col_out_311     ),
    .col_in_312              ( u0_col_out_312     ),
    .col_in_313              ( u0_col_out_313     ),
    .col_in_314              ( u0_col_out_314     ),
    .col_in_315              ( u0_col_out_315     ),
    .col_in_316              ( u0_col_out_316     ),
    .col_in_317              ( u0_col_out_317     ),
    .col_in_318              ( u0_col_out_318     ),
    .col_in_319              ( u0_col_out_319     ),
    .col_in_320              ( u0_col_out_320     ),
    .col_in_321              ( u0_col_out_321     ),
    .col_in_322              ( u0_col_out_322     ),
    .col_in_323              ( u0_col_out_323     ),
    .col_in_324              ( u0_col_out_324     ),
    .col_in_325              ( u0_col_out_325     ),
    .col_in_326              ( u0_col_out_326     ),
    .col_in_327              ( u0_col_out_327     ),
    .col_in_328              ( u0_col_out_328     ),
    .col_in_329              ( u0_col_out_329     ),
    .col_in_330              ( u0_col_out_330     ),
    .col_in_331              ( u0_col_out_331     ),
    .col_in_332              ( u0_col_out_332     ),
    .col_in_333              ( u0_col_out_333     ),
    .col_in_334              ( u0_col_out_334     ),
    .col_in_335              ( u0_col_out_335     ),
    .col_in_336              ( u0_col_out_336     ),
    .col_in_337              ( u0_col_out_337     ),
    .col_in_338              ( u0_col_out_338     ),
    .col_in_339              ( u0_col_out_339     ),
    .col_in_340              ( u0_col_out_340     ),
    .col_in_341              ( u0_col_out_341     ),
    .col_in_342              ( u0_col_out_342     ),
    .col_in_343              ( u0_col_out_343     ),
    .col_in_344              ( u0_col_out_344     ),
    .col_in_345              ( u0_col_out_345     ),
    .col_in_346              ( u0_col_out_346     ),
    .col_in_347              ( u0_col_out_347     ),
    .col_in_348              ( u0_col_out_348     ),
    .col_in_349              ( u0_col_out_349     ),
    .col_in_350              ( u0_col_out_350     ),
    .col_in_351              ( u0_col_out_351     ),
    .col_in_352              ( u0_col_out_352     ),
    .col_in_353              ( u0_col_out_353     ),
    .col_in_354              ( u0_col_out_354     ),
    .col_in_355              ( u0_col_out_355     ),
    .col_in_356              ( u0_col_out_356     ),
    .col_in_357              ( u0_col_out_357     ),
    .col_in_358              ( u0_col_out_358     ),
    .col_in_359              ( u0_col_out_359     ),
    .col_in_360              ( u0_col_out_360     ),
    .col_in_361              ( u0_col_out_361     ),
    .col_in_362              ( u0_col_out_362     ),
    .col_in_363              ( u0_col_out_363     ),
    .col_in_364              ( u0_col_out_364     ),
    .col_in_365              ( u0_col_out_365     ),
    .col_in_366              ( u0_col_out_366     ),
    .col_in_367              ( u0_col_out_367     ),
    .col_in_368              ( u0_col_out_368     ),
    .col_in_369              ( u0_col_out_369     ),
    .col_in_370              ( u0_col_out_370     ),
    .col_in_371              ( u0_col_out_371     ),
    .col_in_372              ( u0_col_out_372     ),
    .col_in_373              ( u0_col_out_373     ),
    .col_in_374              ( u0_col_out_374     ),
    .col_in_375              ( u0_col_out_375     ),
    .col_in_376              ( u0_col_out_376     ),
    .col_in_377              ( u0_col_out_377     ),
    .col_in_378              ( u0_col_out_378     ),
    .col_in_379              ( u0_col_out_379     ),
    .col_in_380              ( u0_col_out_380     ),
    .col_in_381              ( u0_col_out_381     ),
    .col_in_382              ( u0_col_out_382     ),
    .col_in_383              ( u0_col_out_383     ),
    .col_in_384              ( u0_col_out_384     ),
    .col_in_385              ( u0_col_out_385     ),
    .col_in_386              ( u0_col_out_386     ),
    .col_in_387              ( u0_col_out_387     ),
    .col_in_388              ( u0_col_out_388     ),
    .col_in_389              ( u0_col_out_389     ),
    .col_in_390              ( u0_col_out_390     ),
    .col_in_391              ( u0_col_out_391     ),
    .col_in_392              ( u0_col_out_392     ),
    .col_in_393              ( u0_col_out_393     ),
    .col_in_394              ( u0_col_out_394     ),
    .col_in_395              ( u0_col_out_395     ),
    .col_in_396              ( u0_col_out_396     ),
    .col_in_397              ( u0_col_out_397     ),
    .col_in_398              ( u0_col_out_398     ),
    .col_in_399              ( u0_col_out_399     ),
    .col_in_400              ( u0_col_out_400     ),
    .col_in_401              ( u0_col_out_401     ),
    .col_in_402              ( u0_col_out_402     ),
    .col_in_403              ( u0_col_out_403     ),
    .col_in_404              ( u0_col_out_404     ),
    .col_in_405              ( u0_col_out_405     ),
    .col_in_406              ( u0_col_out_406     ),
    .col_in_407              ( u0_col_out_407     ),
    .col_in_408              ( u0_col_out_408     ),
    .col_in_409              ( u0_col_out_409     ),
    .col_in_410              ( u0_col_out_410     ),
    .col_in_411              ( u0_col_out_411     ),
    .col_in_412              ( u0_col_out_412     ),
    .col_in_413              ( u0_col_out_413     ),
    .col_in_414              ( u0_col_out_414     ),
    .col_in_415              ( u0_col_out_415     ),
    .col_in_416              ( u0_col_out_416     ),
    .col_in_417              ( u0_col_out_417     ),
    .col_in_418              ( u0_col_out_418     ),
    .col_in_419              ( u0_col_out_419     ),
    .col_in_420              ( u0_col_out_420     ),
    .col_in_421              ( u0_col_out_421     ),
    .col_in_422              ( u0_col_out_422     ),
    .col_in_423              ( u0_col_out_423     ),
    .col_in_424              ( u0_col_out_424     ),
    .col_in_425              ( u0_col_out_425     ),
    .col_in_426              ( u0_col_out_426     ),
    .col_in_427              ( u0_col_out_427     ),
    .col_in_428              ( u0_col_out_428     ),
    .col_in_429              ( u0_col_out_429     ),
    .col_in_430              ( u0_col_out_430     ),
    .col_in_431              ( u0_col_out_431     ),
    .col_in_432              ( u0_col_out_432     ),
    .col_in_433              ( u0_col_out_433     ),
    .col_in_434              ( u0_col_out_434     ),
    .col_in_435              ( u0_col_out_435     ),
    .col_in_436              ( u0_col_out_436     ),
    .col_in_437              ( u0_col_out_437     ),
    .col_in_438              ( u0_col_out_438     ),
    .col_in_439              ( u0_col_out_439     ),
    .col_in_440              ( u0_col_out_440     ),
    .col_in_441              ( u0_col_out_441     ),
    .col_in_442              ( u0_col_out_442     ),
    .col_in_443              ( u0_col_out_443     ),
    .col_in_444              ( u0_col_out_444     ),
    .col_in_445              ( u0_col_out_445     ),
    .col_in_446              ( u0_col_out_446     ),
    .col_in_447              ( u0_col_out_447     ),
    .col_in_448              ( u0_col_out_448     ),
    .col_in_449              ( u0_col_out_449     ),
    .col_in_450              ( u0_col_out_450     ),
    .col_in_451              ( u0_col_out_451     ),
    .col_in_452              ( u0_col_out_452     ),
    .col_in_453              ( u0_col_out_453     ),
    .col_in_454              ( u0_col_out_454     ),
    .col_in_455              ( u0_col_out_455     ),
    .col_in_456              ( u0_col_out_456     ),
    .col_in_457              ( u0_col_out_457     ),
    .col_in_458              ( u0_col_out_458     ),
    .col_in_459              ( u0_col_out_459     ),
    .col_in_460              ( u0_col_out_460     ),
    .col_in_461              ( u0_col_out_461     ),
    .col_in_462              ( u0_col_out_462     ),
    .col_in_463              ( u0_col_out_463     ),
    .col_in_464              ( u0_col_out_464     ),
    .col_in_465              ( u0_col_out_465     ),
    .col_in_466              ( u0_col_out_466     ),
    .col_in_467              ( u0_col_out_467     ),
    .col_in_468              ( u0_col_out_468     ),
    .col_in_469              ( u0_col_out_469     ),
    .col_in_470              ( u0_col_out_470     ),
    .col_in_471              ( u0_col_out_471     ),
    .col_in_472              ( u0_col_out_472     ),
    .col_in_473              ( u0_col_out_473     ),
    .col_in_474              ( u0_col_out_474     ),
    .col_in_475              ( u0_col_out_475     ),
    .col_in_476              ( u0_col_out_476     ),
    .col_in_477              ( u0_col_out_477     ),
    .col_in_478              ( u0_col_out_478     ),
    .col_in_479              ( u0_col_out_479     ),
    .col_in_480              ( u0_col_out_480     ),
    .col_in_481              ( u0_col_out_481     ),
    .col_in_482              ( u0_col_out_482     ),
    .col_in_483              ( u0_col_out_483     ),
    .col_in_484              ( u0_col_out_484     ),
    .col_in_485              ( u0_col_out_485     ),
    .col_in_486              ( u0_col_out_486     ),
    .col_in_487              ( u0_col_out_487     ),
    .col_in_488              ( u0_col_out_488     ),
    .col_in_489              ( u0_col_out_489     ),
    .col_in_490              ( u0_col_out_490     ),
    .col_in_491              ( u0_col_out_491     ),
    .col_in_492              ( u0_col_out_492     ),
    .col_in_493              ( u0_col_out_493     ),
    .col_in_494              ( u0_col_out_494     ),
    .col_in_495              ( u0_col_out_495     ),
    .col_in_496              ( u0_col_out_496     ),
    .col_in_497              ( u0_col_out_497     ),
    .col_in_498              ( u0_col_out_498     ),
    .col_in_499              ( u0_col_out_499     ),
    .col_in_500              ( u0_col_out_500     ),
    .col_in_501              ( u0_col_out_501     ),
    .col_in_502              ( u0_col_out_502     ),
    .col_in_503              ( u0_col_out_503     ),
    .col_in_504              ( u0_col_out_504     ),
    .col_in_505              ( u0_col_out_505     ),
    .col_in_506              ( u0_col_out_506     ),
    .col_in_507              ( u0_col_out_507     ),
    .col_in_508              ( u0_col_out_508     ),
    .col_in_509              ( u0_col_out_509     ),
    .col_in_510              ( u0_col_out_510     ),
    .col_in_511              ( u0_col_out_511     ),
    .col_in_512              ( u0_col_out_512     ),
    .col_in_513              ( u0_col_out_513     ),
    .col_in_514              ( u0_col_out_514     ),
    .col_in_515              ( u0_col_out_515     ),
    .col_in_516              ( u0_col_out_516     ),
    .col_in_517              ( u0_col_out_517     ),
    .col_in_518              ( u0_col_out_518     ),
    .col_in_519              ( u0_col_out_519     ),
    .col_in_520              ( u0_col_out_520     ),
    .col_in_521              ( u0_col_out_521     ),
    .col_in_522              ( u0_col_out_522     ),
    .col_in_523              ( u0_col_out_523     ),
    .col_in_524              ( u0_col_out_524     ),
    .col_in_525              ( u0_col_out_525     ),
    .col_in_526              ( u0_col_out_526     ),
    .col_in_527              ( u0_col_out_527     ),
    .col_in_528              ( u0_col_out_528     ),
    .col_in_529              ( u0_col_out_529     ),
    .col_in_530              ( u0_col_out_530     ),
    .col_in_531              ( u0_col_out_531     ),
    .col_in_532              ( u0_col_out_532     ),
    .col_in_533              ( u0_col_out_533     ),
    .col_in_534              ( u0_col_out_534     ),
    .col_in_535              ( u0_col_out_535     ),
    .col_in_536              ( u0_col_out_536     ),
    .col_in_537              ( u0_col_out_537     ),
    .col_in_538              ( u0_col_out_538     ),
    .col_in_539              ( u0_col_out_539     ),
    .col_in_540              ( u0_col_out_540     ),
    .col_in_541              ( u0_col_out_541     ),
    .col_in_542              ( u0_col_out_542     ),
    .col_in_543              ( u0_col_out_543     ),
    .col_in_544              ( u0_col_out_544     ),
    .col_in_545              ( u0_col_out_545     ),
    .col_in_546              ( u0_col_out_546     ),
    .col_in_547              ( u0_col_out_547     ),
    .col_in_548              ( u0_col_out_548     ),
    .col_in_549              ( u0_col_out_549     ),
    .col_in_550              ( u0_col_out_550     ),
    .col_in_551              ( u0_col_out_551     ),
    .col_in_552              ( u0_col_out_552     ),
    .col_in_553              ( u0_col_out_553     ),
    .col_in_554              ( u0_col_out_554     ),
    .col_in_555              ( u0_col_out_555     ),
    .col_in_556              ( u0_col_out_556     ),
    .col_in_557              ( u0_col_out_557     ),
    .col_in_558              ( u0_col_out_558     ),
    .col_in_559              ( u0_col_out_559     ),
    .col_in_560              ( u0_col_out_560     ),
    .col_in_561              ( u0_col_out_561     ),
    .col_in_562              ( u0_col_out_562     ),
    .col_in_563              ( u0_col_out_563     ),
    .col_in_564              ( u0_col_out_564     ),
    .col_in_565              ( u0_col_out_565     ),
    .col_in_566              ( u0_col_out_566     ),
    .col_in_567              ( u0_col_out_567     ),
    .col_in_568              ( u0_col_out_568     ),
    .col_in_569              ( u0_col_out_569     ),
    .col_in_570              ( u0_col_out_570     ),
    .col_in_571              ( u0_col_out_571     ),
    .col_in_572              ( u0_col_out_572     ),
    .col_in_573              ( u0_col_out_573     ),
    .col_in_574              ( u0_col_out_574     ),
    .col_in_575              ( u0_col_out_575     ),
    .col_in_576              ( u0_col_out_576     ),
    .col_in_577              ( u0_col_out_577     ),
    .col_in_578              ( u0_col_out_578     ),
    .col_in_579              ( u0_col_out_579     ),
    .col_in_580              ( u0_col_out_580     ),
    .col_in_581              ( u0_col_out_581     ),
    .col_in_582              ( u0_col_out_582     ),
    .col_in_583              ( u0_col_out_583     ),
    .col_in_584              ( u0_col_out_584     ),
    .col_in_585              ( u0_col_out_585     ),
    .col_in_586              ( u0_col_out_586     ),
    .col_in_587              ( u0_col_out_587     ),
    .col_in_588              ( u0_col_out_588     ),
    .col_in_589              ( u0_col_out_589     ),
    .col_in_590              ( u0_col_out_590     ),
    .col_in_591              ( u0_col_out_591     ),
    .col_in_592              ( u0_col_out_592     ),
    .col_in_593              ( u0_col_out_593     ),
    .col_in_594              ( u0_col_out_594     ),
    .col_in_595              ( u0_col_out_595     ),
    .col_in_596              ( u0_col_out_596     ),
    .col_in_597              ( u0_col_out_597     ),
    .col_in_598              ( u0_col_out_598     ),
    .col_in_599              ( u0_col_out_599     ),
    .col_in_600              ( u0_col_out_600     ),
    .col_in_601              ( u0_col_out_601     ),
    .col_in_602              ( u0_col_out_602     ),
    .col_in_603              ( u0_col_out_603     ),
    .col_in_604              ( u0_col_out_604     ),
    .col_in_605              ( u0_col_out_605     ),
    .col_in_606              ( u0_col_out_606     ),
    .col_in_607              ( u0_col_out_607     ),
    .col_in_608              ( u0_col_out_608     ),
    .col_in_609              ( u0_col_out_609     ),
    .col_in_610              ( u0_col_out_610     ),
    .col_in_611              ( u0_col_out_611     ),
    .col_in_612              ( u0_col_out_612     ),
    .col_in_613              ( u0_col_out_613     ),
    .col_in_614              ( u0_col_out_614     ),
    .col_in_615              ( u0_col_out_615     ),
    .col_in_616              ( u0_col_out_616     ),
    .col_in_617              ( u0_col_out_617     ),
    .col_in_618              ( u0_col_out_618     ),
    .col_in_619              ( u0_col_out_619     ),
    .col_in_620              ( u0_col_out_620     ),
    .col_in_621              ( u0_col_out_621     ),
    .col_in_622              ( u0_col_out_622     ),
    .col_in_623              ( u0_col_out_623     ),
    .col_in_624              ( u0_col_out_624     ),
    .col_in_625              ( u0_col_out_625     ),
    .col_in_626              ( u0_col_out_626     ),
    .col_in_627              ( u0_col_out_627     ),
    .col_in_628              ( u0_col_out_628     ),
    .col_in_629              ( u0_col_out_629     ),
    .col_in_630              ( u0_col_out_630     ),
    .col_in_631              ( u0_col_out_631     ),
    .col_in_632              ( u0_col_out_632     ),
    .col_in_633              ( u0_col_out_633     ),
    .col_in_634              ( u0_col_out_634     ),
    .col_in_635              ( u0_col_out_635     ),
    .col_in_636              ( u0_col_out_636     ),
    .col_in_637              ( u0_col_out_637     ),
    .col_in_638              ( u0_col_out_638     ),
    .col_in_639              ( u0_col_out_639     ),
    .col_in_640              ( u0_col_out_640     ),
    .col_in_641              ( u0_col_out_641     ),
    .col_in_642              ( u0_col_out_642     ),
    .col_in_643              ( u0_col_out_643     ),
    .col_in_644              ( u0_col_out_644     ),
    .col_in_645              ( u0_col_out_645     ),
    .col_in_646              ( u0_col_out_646     ),
    .col_in_647              ( u0_col_out_647     ),
    .col_in_648              ( u0_col_out_648     ),
    .col_in_649              ( u0_col_out_649     ),
    .col_in_650              ( u0_col_out_650     ),
    .col_in_651              ( u0_col_out_651     ),
    .col_in_652              ( u0_col_out_652     ),
    .col_in_653              ( u0_col_out_653     ),
    .col_in_654              ( u0_col_out_654     ),
    .col_in_655              ( u0_col_out_655     ),
    .col_in_656              ( u0_col_out_656     ),
    .col_in_657              ( u0_col_out_657     ),
    .col_in_658              ( u0_col_out_658     ),
    .col_in_659              ( u0_col_out_659     ),
    .col_in_660              ( u0_col_out_660     ),
    .col_in_661              ( u0_col_out_661     ),
    .col_in_662              ( u0_col_out_662     ),
    .col_in_663              ( u0_col_out_663     ),
    .col_in_664              ( u0_col_out_664     ),
    .col_in_665              ( u0_col_out_665     ),
    .col_in_666              ( u0_col_out_666     ),
    .col_in_667              ( u0_col_out_667     ),
    .col_in_668              ( u0_col_out_668     ),
    .col_in_669              ( u0_col_out_669     ),
    .col_in_670              ( u0_col_out_670     ),
    .col_in_671              ( u0_col_out_671     ),
    .col_in_672              ( u0_col_out_672     ),
    .col_in_673              ( u0_col_out_673     ),
    .col_in_674              ( u0_col_out_674     ),
    .col_in_675              ( u0_col_out_675     ),
    .col_in_676              ( u0_col_out_676     ),
    .col_in_677              ( u0_col_out_677     ),
    .col_in_678              ( u0_col_out_678     ),
    .col_in_679              ( u0_col_out_679     ),
    .col_in_680              ( u0_col_out_680     ),
    .col_in_681              ( u0_col_out_681     ),
    .col_in_682              ( u0_col_out_682     ),
    .col_in_683              ( u0_col_out_683     ),
    .col_in_684              ( u0_col_out_684     ),
    .col_in_685              ( u0_col_out_685     ),
    .col_in_686              ( u0_col_out_686     ),
    .col_in_687              ( u0_col_out_687     ),
    .col_in_688              ( u0_col_out_688     ),
    .col_in_689              ( u0_col_out_689     ),
    .col_in_690              ( u0_col_out_690     ),
    .col_in_691              ( u0_col_out_691     ),
    .col_in_692              ( u0_col_out_692     ),
    .col_in_693              ( u0_col_out_693     ),
    .col_in_694              ( u0_col_out_694     ),
    .col_in_695              ( u0_col_out_695     ),
    .col_in_696              ( u0_col_out_696     ),
    .col_in_697              ( u0_col_out_697     ),
    .col_in_698              ( u0_col_out_698     ),
    .col_in_699              ( u0_col_out_699     ),
    .col_in_700              ( u0_col_out_700     ),
    .col_in_701              ( u0_col_out_701     ),
    .col_in_702              ( u0_col_out_702     ),
    .col_in_703              ( u0_col_out_703     ),
    .col_in_704              ( u0_col_out_704     ),
    .col_in_705              ( u0_col_out_705     ),
    .col_in_706              ( u0_col_out_706     ),
    .col_in_707              ( u0_col_out_707     ),
    .col_in_708              ( u0_col_out_708     ),
    .col_in_709              ( u0_col_out_709     ),
    .col_in_710              ( u0_col_out_710     ),
    .col_in_711              ( u0_col_out_711     ),
    .col_in_712              ( u0_col_out_712     ),
    .col_in_713              ( u0_col_out_713     ),
    .col_in_714              ( u0_col_out_714     ),
    .col_in_715              ( u0_col_out_715     ),
    .col_in_716              ( u0_col_out_716     ),
    .col_in_717              ( u0_col_out_717     ),
    .col_in_718              ( u0_col_out_718     ),
    .col_in_719              ( u0_col_out_719     ),
    .col_in_720              ( u0_col_out_720     ),
    .col_in_721              ( u0_col_out_721     ),
    .col_in_722              ( u0_col_out_722     ),
    .col_in_723              ( u0_col_out_723     ),
    .col_in_724              ( u0_col_out_724     ),
    .col_in_725              ( u0_col_out_725     ),
    .col_in_726              ( u0_col_out_726     ),
    .col_in_727              ( u0_col_out_727     ),
    .col_in_728              ( u0_col_out_728     ),
    .col_in_729              ( u0_col_out_729     ),
    .col_in_730              ( u0_col_out_730     ),
    .col_in_731              ( u0_col_out_731     ),
    .col_in_732              ( u0_col_out_732     ),
    .col_in_733              ( u0_col_out_733     ),
    .col_in_734              ( u0_col_out_734     ),
    .col_in_735              ( u0_col_out_735     ),
    .col_in_736              ( u0_col_out_736     ),
    .col_in_737              ( u0_col_out_737     ),
    .col_in_738              ( u0_col_out_738     ),
    .col_in_739              ( u0_col_out_739     ),
    .col_in_740              ( u0_col_out_740     ),
    .col_in_741              ( u0_col_out_741     ),
    .col_in_742              ( u0_col_out_742     ),
    .col_in_743              ( u0_col_out_743     ),
    .col_in_744              ( u0_col_out_744     ),
    .col_in_745              ( u0_col_out_745     ),
    .col_in_746              ( u0_col_out_746     ),
    .col_in_747              ( u0_col_out_747     ),
    .col_in_748              ( u0_col_out_748     ),
    .col_in_749              ( u0_col_out_749     ),
    .col_in_750              ( u0_col_out_750     ),
    .col_in_751              ( u0_col_out_751     ),
    .col_in_752              ( u0_col_out_752     ),
    .col_in_753              ( u0_col_out_753     ),
    .col_in_754              ( u0_col_out_754     ),
    .col_in_755              ( u0_col_out_755     ),
    .col_in_756              ( u0_col_out_756     ),
    .col_in_757              ( u0_col_out_757     ),
    .col_in_758              ( u0_col_out_758     ),
    .col_in_759              ( u0_col_out_759     ),
    .col_in_760              ( u0_col_out_760     ),
    .col_in_761              ( u0_col_out_761     ),
    .col_in_762              ( u0_col_out_762     ),
    .col_in_763              ( u0_col_out_763     ),
    .col_in_764              ( u0_col_out_764     ),
    .col_in_765              ( u0_col_out_765     ),
    .col_in_766              ( u0_col_out_766     ),
    .col_in_767              ( u0_col_out_767     ),
    .col_in_768              ( u0_col_out_768     ),
    .col_in_769              ( u0_col_out_769     ),
    .col_in_770              ( u0_col_out_770     ),
    .col_in_771              ( u0_col_out_771     ),
    .col_in_772              ( u0_col_out_772     ),
    .col_in_773              ( u0_col_out_773     ),
    .col_in_774              ( u0_col_out_774     ),
    .col_in_775              ( u0_col_out_775     ),
    .col_in_776              ( u0_col_out_776     ),
    .col_in_777              ( u0_col_out_777     ),
    .col_in_778              ( u0_col_out_778     ),
    .col_in_779              ( u0_col_out_779     ),
    .col_in_780              ( u0_col_out_780     ),
    .col_in_781              ( u0_col_out_781     ),
    .col_in_782              ( u0_col_out_782     ),
    .col_in_783              ( u0_col_out_783     ),
    .col_in_784              ( u0_col_out_784     ),
    .col_in_785              ( u0_col_out_785     ),
    .col_in_786              ( u0_col_out_786     ),
    .col_in_787              ( u0_col_out_787     ),
    .col_in_788              ( u0_col_out_788     ),
    .col_in_789              ( u0_col_out_789     ),
    .col_in_790              ( u0_col_out_790     ),
    .col_in_791              ( u0_col_out_791     ),
    .col_in_792              ( u0_col_out_792     ),
    .col_in_793              ( u0_col_out_793     ),
    .col_in_794              ( u0_col_out_794     ),
    .col_in_795              ( u0_col_out_795     ),
    .col_in_796              ( u0_col_out_796     ),
    .col_in_797              ( u0_col_out_797     ),
    .col_in_798              ( u0_col_out_798     ),
    .col_in_799              ( u0_col_out_799     ),
    .col_in_800              ( u0_col_out_800     ),
    .col_in_801              ( u0_col_out_801     ),
    .col_in_802              ( u0_col_out_802     ),
    .col_in_803              ( u0_col_out_803     ),
    .col_in_804              ( u0_col_out_804     ),
    .col_in_805              ( u0_col_out_805     ),
    .col_in_806              ( u0_col_out_806     ),
    .col_in_807              ( u0_col_out_807     ),
    .col_in_808              ( u0_col_out_808     ),
    .col_in_809              ( u0_col_out_809     ),
    .col_in_810              ( u0_col_out_810     ),
    .col_in_811              ( u0_col_out_811     ),
    .col_in_812              ( u0_col_out_812     ),
    .col_in_813              ( u0_col_out_813     ),
    .col_in_814              ( u0_col_out_814     ),
    .col_in_815              ( u0_col_out_815     ),
    .col_in_816              ( u0_col_out_816     ),
    .col_in_817              ( u0_col_out_817     ),
    .col_in_818              ( u0_col_out_818     ),
    .col_in_819              ( u0_col_out_819     ),
    .col_in_820              ( u0_col_out_820     ),
    .col_in_821              ( u0_col_out_821     ),
    .col_in_822              ( u0_col_out_822     ),
    .col_in_823              ( u0_col_out_823     ),
    .col_in_824              ( u0_col_out_824     ),
    .col_in_825              ( u0_col_out_825     ),
    .col_in_826              ( u0_col_out_826     ),
    .col_in_827              ( u0_col_out_827     ),
    .col_in_828              ( u0_col_out_828     ),
    .col_in_829              ( u0_col_out_829     ),
    .col_in_830              ( u0_col_out_830     ),
    .col_in_831              ( u0_col_out_831     ),
    .col_in_832              ( u0_col_out_832     ),
    .col_in_833              ( u0_col_out_833     ),
    .col_in_834              ( u0_col_out_834     ),
    .col_in_835              ( u0_col_out_835     ),
    .col_in_836              ( u0_col_out_836     ),
    .col_in_837              ( u0_col_out_837     ),
    .col_in_838              ( u0_col_out_838     ),
    .col_in_839              ( u0_col_out_839     ),
    .col_in_840              ( u0_col_out_840     ),
    .col_in_841              ( u0_col_out_841     ),
    .col_in_842              ( u0_col_out_842     ),
    .col_in_843              ( u0_col_out_843     ),
    .col_in_844              ( u0_col_out_844     ),
    .col_in_845              ( u0_col_out_845     ),
    .col_in_846              ( u0_col_out_846     ),
    .col_in_847              ( u0_col_out_847     ),
    .col_in_848              ( u0_col_out_848     ),
    .col_in_849              ( u0_col_out_849     ),
    .col_in_850              ( u0_col_out_850     ),
    .col_in_851              ( u0_col_out_851     ),
    .col_in_852              ( u0_col_out_852     ),
    .col_in_853              ( u0_col_out_853     ),
    .col_in_854              ( u0_col_out_854     ),
    .col_in_855              ( u0_col_out_855     ),
    .col_in_856              ( u0_col_out_856     ),
    .col_in_857              ( u0_col_out_857     ),
    .col_in_858              ( u0_col_out_858     ),
    .col_in_859              ( u0_col_out_859     ),
    .col_in_860              ( u0_col_out_860     ),
    .col_in_861              ( u0_col_out_861     ),
    .col_in_862              ( u0_col_out_862     ),
    .col_in_863              ( u0_col_out_863     ),
    .col_in_864              ( u0_col_out_864     ),
    .col_in_865              ( u0_col_out_865     ),
    .col_in_866              ( u0_col_out_866     ),
    .col_in_867              ( u0_col_out_867     ),
    .col_in_868              ( u0_col_out_868     ),
    .col_in_869              ( u0_col_out_869     ),
    .col_in_870              ( u0_col_out_870     ),
    .col_in_871              ( u0_col_out_871     ),
    .col_in_872              ( u0_col_out_872     ),
    .col_in_873              ( u0_col_out_873     ),
    .col_in_874              ( u0_col_out_874     ),
    .col_in_875              ( u0_col_out_875     ),
    .col_in_876              ( u0_col_out_876     ),
    .col_in_877              ( u0_col_out_877     ),
    .col_in_878              ( u0_col_out_878     ),
    .col_in_879              ( u0_col_out_879     ),
    .col_in_880              ( u0_col_out_880     ),
    .col_in_881              ( u0_col_out_881     ),
    .col_in_882              ( u0_col_out_882     ),
    .col_in_883              ( u0_col_out_883     ),
    .col_in_884              ( u0_col_out_884     ),
    .col_in_885              ( u0_col_out_885     ),
    .col_in_886              ( u0_col_out_886     ),
    .col_in_887              ( u0_col_out_887     ),
    .col_in_888              ( u0_col_out_888     ),
    .col_in_889              ( u0_col_out_889     ),
    .col_in_890              ( u0_col_out_890     ),
    .col_in_891              ( u0_col_out_891     ),
    .col_in_892              ( u0_col_out_892     ),
    .col_in_893              ( u0_col_out_893     ),
    .col_in_894              ( u0_col_out_894     ),
    .col_in_895              ( u0_col_out_895     ),
    .col_in_896              ( u0_col_out_896     ),
    .col_in_897              ( u0_col_out_897     ),
    .col_in_898              ( u0_col_out_898     ),
    .col_in_899              ( u0_col_out_899     ),
    .col_in_900              ( u0_col_out_900     ),
    .col_in_901              ( u0_col_out_901     ),
    .col_in_902              ( u0_col_out_902     ),
    .col_in_903              ( u0_col_out_903     ),
    .col_in_904              ( u0_col_out_904     ),
    .col_in_905              ( u0_col_out_905     ),
    .col_in_906              ( u0_col_out_906     ),
    .col_in_907              ( u0_col_out_907     ),
    .col_in_908              ( u0_col_out_908     ),
    .col_in_909              ( u0_col_out_909     ),
    .col_in_910              ( u0_col_out_910     ),
    .col_in_911              ( u0_col_out_911     ),
    .col_in_912              ( u0_col_out_912     ),
    .col_in_913              ( u0_col_out_913     ),
    .col_in_914              ( u0_col_out_914     ),
    .col_in_915              ( u0_col_out_915     ),
    .col_in_916              ( u0_col_out_916     ),
    .col_in_917              ( u0_col_out_917     ),
    .col_in_918              ( u0_col_out_918     ),
    .col_in_919              ( u0_col_out_919     ),
    .col_in_920              ( u0_col_out_920     ),
    .col_in_921              ( u0_col_out_921     ),
    .col_in_922              ( u0_col_out_922     ),
    .col_in_923              ( u0_col_out_923     ),
    .col_in_924              ( u0_col_out_924     ),
    .col_in_925              ( u0_col_out_925     ),
    .col_in_926              ( u0_col_out_926     ),
    .col_in_927              ( u0_col_out_927     ),
    .col_in_928              ( u0_col_out_928     ),
    .col_in_929              ( u0_col_out_929     ),
    .col_in_930              ( u0_col_out_930     ),
    .col_in_931              ( u0_col_out_931     ),
    .col_in_932              ( u0_col_out_932     ),
    .col_in_933              ( u0_col_out_933     ),
    .col_in_934              ( u0_col_out_934     ),
    .col_in_935              ( u0_col_out_935     ),
    .col_in_936              ( u0_col_out_936     ),
    .col_in_937              ( u0_col_out_937     ),
    .col_in_938              ( u0_col_out_938     ),
    .col_in_939              ( u0_col_out_939     ),
    .col_in_940              ( u0_col_out_940     ),
    .col_in_941              ( u0_col_out_941     ),
    .col_in_942              ( u0_col_out_942     ),
    .col_in_943              ( u0_col_out_943     ),
    .col_in_944              ( u0_col_out_944     ),
    .col_in_945              ( u0_col_out_945     ),
    .col_in_946              ( u0_col_out_946     ),
    .col_in_947              ( u0_col_out_947     ),
    .col_in_948              ( u0_col_out_948     ),
    .col_in_949              ( u0_col_out_949     ),
    .col_in_950              ( u0_col_out_950     ),
    .col_in_951              ( u0_col_out_951     ),
    .col_in_952              ( u0_col_out_952     ),
    .col_in_953              ( u0_col_out_953     ),
    .col_in_954              ( u0_col_out_954     ),
    .col_in_955              ( u0_col_out_955     ),
    .col_in_956              ( u0_col_out_956     ),
    .col_in_957              ( u0_col_out_957     ),
    .col_in_958              ( u0_col_out_958     ),
    .col_in_959              ( u0_col_out_959     ),
    .col_in_960              ( u0_col_out_960     ),
    .col_in_961              ( u0_col_out_961     ),
    .col_in_962              ( u0_col_out_962     ),
    .col_in_963              ( u0_col_out_963     ),
    .col_in_964              ( u0_col_out_964     ),
    .col_in_965              ( u0_col_out_965     ),
    .col_in_966              ( u0_col_out_966     ),
    .col_in_967              ( u0_col_out_967     ),
    .col_in_968              ( u0_col_out_968     ),
    .col_in_969              ( u0_col_out_969     ),
    .col_in_970              ( u0_col_out_970     ),
    .col_in_971              ( u0_col_out_971     ),
    .col_in_972              ( u0_col_out_972     ),
    .col_in_973              ( u0_col_out_973     ),
    .col_in_974              ( u0_col_out_974     ),
    .col_in_975              ( u0_col_out_975     ),
    .col_in_976              ( u0_col_out_976     ),
    .col_in_977              ( u0_col_out_977     ),
    .col_in_978              ( u0_col_out_978     ),
    .col_in_979              ( u0_col_out_979     ),
    .col_in_980              ( u0_col_out_980     ),
    .col_in_981              ( u0_col_out_981     ),
    .col_in_982              ( u0_col_out_982     ),
    .col_in_983              ( u0_col_out_983     ),
    .col_in_984              ( u0_col_out_984     ),
    .col_in_985              ( u0_col_out_985     ),
    .col_in_986              ( u0_col_out_986     ),
    .col_in_987              ( u0_col_out_987     ),
    .col_in_988              ( u0_col_out_988     ),
    .col_in_989              ( u0_col_out_989     ),
    .col_in_990              ( u0_col_out_990     ),
    .col_in_991              ( u0_col_out_991     ),
    .col_in_992              ( u0_col_out_992     ),
    .col_in_993              ( u0_col_out_993     ),
    .col_in_994              ( u0_col_out_994     ),
    .col_in_995              ( u0_col_out_995     ),
    .col_in_996              ( u0_col_out_996     ),
    .col_in_997              ( u0_col_out_997     ),
    .col_in_998              ( u0_col_out_998     ),
    .col_in_999              ( u0_col_out_999     ),
    .col_in_1000             ( u0_col_out_1000    ),
    .col_in_1001             ( u0_col_out_1001    ),
    .col_in_1002             ( u0_col_out_1002    ),
    .col_in_1003             ( u0_col_out_1003    ),
    .col_in_1004             ( u0_col_out_1004    ),
    .col_in_1005             ( u0_col_out_1005    ),
    .col_in_1006             ( u0_col_out_1006    ),
    .col_in_1007             ( u0_col_out_1007    ),
    .col_in_1008             ( u0_col_out_1008    ),
    .col_in_1009             ( u0_col_out_1009    ),
    .col_in_1010             ( u0_col_out_1010    ),
    .col_in_1011             ( u0_col_out_1011    ),
    .col_in_1012             ( u0_col_out_1012    ),
    .col_in_1013             ( u0_col_out_1013    ),
    .col_in_1014             ( u0_col_out_1014    ),
    .col_in_1015             ( u0_col_out_1015    ),
    .col_in_1016             ( u0_col_out_1016    ),
    .col_in_1017             ( u0_col_out_1017    ),
    .col_in_1018             ( u0_col_out_1018    ),
    .col_in_1019             ( u0_col_out_1019    ),
    .col_in_1020             ( u0_col_out_1020    ),
    .col_in_1021             ( u0_col_out_1021    ),
    .col_in_1022             ( u0_col_out_1022    ),
    .col_in_1023             ( u0_col_out_1023    ),
    .col_in_1024             ( u0_col_out_1024    ),
    .col_in_1025             ( u0_col_out_1025    ),
    .col_in_1026             ( u0_col_out_1026    ),
    .col_in_1027             ( u0_col_out_1027    ),
    .col_in_1028             ( u0_col_out_1028    ),
    .col_in_1029             ( u0_col_out_1029    ),
    .col_in_1030             ( u0_col_out_1030    ),
    .col_in_1031             ( u0_col_out_1031    ),
    .col_in_1032             ( u0_col_out_1032    ),


    .col_out_0               ( u1_col_out_0      ),
    .col_out_1               ( u1_col_out_1      ),
    .col_out_2               ( u1_col_out_2      ),
    .col_out_3               ( u1_col_out_3      ),
    .col_out_4               ( u1_col_out_4      ),
    .col_out_5               ( u1_col_out_5      ),
    .col_out_6               ( u1_col_out_6      ),
    .col_out_7               ( u1_col_out_7      ),
    .col_out_8               ( u1_col_out_8      ),
    .col_out_9               ( u1_col_out_9      ),
    .col_out_10              ( u1_col_out_10     ),
    .col_out_11              ( u1_col_out_11     ),
    .col_out_12              ( u1_col_out_12     ),
    .col_out_13              ( u1_col_out_13     ),
    .col_out_14              ( u1_col_out_14     ),
    .col_out_15              ( u1_col_out_15     ),
    .col_out_16              ( u1_col_out_16     ),
    .col_out_17              ( u1_col_out_17     ),
    .col_out_18              ( u1_col_out_18     ),
    .col_out_19              ( u1_col_out_19     ),
    .col_out_20              ( u1_col_out_20     ),
    .col_out_21              ( u1_col_out_21     ),
    .col_out_22              ( u1_col_out_22     ),
    .col_out_23              ( u1_col_out_23     ),
    .col_out_24              ( u1_col_out_24     ),
    .col_out_25              ( u1_col_out_25     ),
    .col_out_26              ( u1_col_out_26     ),
    .col_out_27              ( u1_col_out_27     ),
    .col_out_28              ( u1_col_out_28     ),
    .col_out_29              ( u1_col_out_29     ),
    .col_out_30              ( u1_col_out_30     ),
    .col_out_31              ( u1_col_out_31     ),
    .col_out_32              ( u1_col_out_32     ),
    .col_out_33              ( u1_col_out_33     ),
    .col_out_34              ( u1_col_out_34     ),
    .col_out_35              ( u1_col_out_35     ),
    .col_out_36              ( u1_col_out_36     ),
    .col_out_37              ( u1_col_out_37     ),
    .col_out_38              ( u1_col_out_38     ),
    .col_out_39              ( u1_col_out_39     ),
    .col_out_40              ( u1_col_out_40     ),
    .col_out_41              ( u1_col_out_41     ),
    .col_out_42              ( u1_col_out_42     ),
    .col_out_43              ( u1_col_out_43     ),
    .col_out_44              ( u1_col_out_44     ),
    .col_out_45              ( u1_col_out_45     ),
    .col_out_46              ( u1_col_out_46     ),
    .col_out_47              ( u1_col_out_47     ),
    .col_out_48              ( u1_col_out_48     ),
    .col_out_49              ( u1_col_out_49     ),
    .col_out_50              ( u1_col_out_50     ),
    .col_out_51              ( u1_col_out_51     ),
    .col_out_52              ( u1_col_out_52     ),
    .col_out_53              ( u1_col_out_53     ),
    .col_out_54              ( u1_col_out_54     ),
    .col_out_55              ( u1_col_out_55     ),
    .col_out_56              ( u1_col_out_56     ),
    .col_out_57              ( u1_col_out_57     ),
    .col_out_58              ( u1_col_out_58     ),
    .col_out_59              ( u1_col_out_59     ),
    .col_out_60              ( u1_col_out_60     ),
    .col_out_61              ( u1_col_out_61     ),
    .col_out_62              ( u1_col_out_62     ),
    .col_out_63              ( u1_col_out_63     ),
    .col_out_64              ( u1_col_out_64     ),
    .col_out_65              ( u1_col_out_65     ),
    .col_out_66              ( u1_col_out_66     ),
    .col_out_67              ( u1_col_out_67     ),
    .col_out_68              ( u1_col_out_68     ),
    .col_out_69              ( u1_col_out_69     ),
    .col_out_70              ( u1_col_out_70     ),
    .col_out_71              ( u1_col_out_71     ),
    .col_out_72              ( u1_col_out_72     ),
    .col_out_73              ( u1_col_out_73     ),
    .col_out_74              ( u1_col_out_74     ),
    .col_out_75              ( u1_col_out_75     ),
    .col_out_76              ( u1_col_out_76     ),
    .col_out_77              ( u1_col_out_77     ),
    .col_out_78              ( u1_col_out_78     ),
    .col_out_79              ( u1_col_out_79     ),
    .col_out_80              ( u1_col_out_80     ),
    .col_out_81              ( u1_col_out_81     ),
    .col_out_82              ( u1_col_out_82     ),
    .col_out_83              ( u1_col_out_83     ),
    .col_out_84              ( u1_col_out_84     ),
    .col_out_85              ( u1_col_out_85     ),
    .col_out_86              ( u1_col_out_86     ),
    .col_out_87              ( u1_col_out_87     ),
    .col_out_88              ( u1_col_out_88     ),
    .col_out_89              ( u1_col_out_89     ),
    .col_out_90              ( u1_col_out_90     ),
    .col_out_91              ( u1_col_out_91     ),
    .col_out_92              ( u1_col_out_92     ),
    .col_out_93              ( u1_col_out_93     ),
    .col_out_94              ( u1_col_out_94     ),
    .col_out_95              ( u1_col_out_95     ),
    .col_out_96              ( u1_col_out_96     ),
    .col_out_97              ( u1_col_out_97     ),
    .col_out_98              ( u1_col_out_98     ),
    .col_out_99              ( u1_col_out_99     ),
    .col_out_100             ( u1_col_out_100    ),
    .col_out_101             ( u1_col_out_101    ),
    .col_out_102             ( u1_col_out_102    ),
    .col_out_103             ( u1_col_out_103    ),
    .col_out_104             ( u1_col_out_104    ),
    .col_out_105             ( u1_col_out_105    ),
    .col_out_106             ( u1_col_out_106    ),
    .col_out_107             ( u1_col_out_107    ),
    .col_out_108             ( u1_col_out_108    ),
    .col_out_109             ( u1_col_out_109    ),
    .col_out_110             ( u1_col_out_110    ),
    .col_out_111             ( u1_col_out_111    ),
    .col_out_112             ( u1_col_out_112    ),
    .col_out_113             ( u1_col_out_113    ),
    .col_out_114             ( u1_col_out_114    ),
    .col_out_115             ( u1_col_out_115    ),
    .col_out_116             ( u1_col_out_116    ),
    .col_out_117             ( u1_col_out_117    ),
    .col_out_118             ( u1_col_out_118    ),
    .col_out_119             ( u1_col_out_119    ),
    .col_out_120             ( u1_col_out_120    ),
    .col_out_121             ( u1_col_out_121    ),
    .col_out_122             ( u1_col_out_122    ),
    .col_out_123             ( u1_col_out_123    ),
    .col_out_124             ( u1_col_out_124    ),
    .col_out_125             ( u1_col_out_125    ),
    .col_out_126             ( u1_col_out_126    ),
    .col_out_127             ( u1_col_out_127    ),
    .col_out_128             ( u1_col_out_128    ),
    .col_out_129             ( u1_col_out_129    ),
    .col_out_130             ( u1_col_out_130    ),
    .col_out_131             ( u1_col_out_131    ),
    .col_out_132             ( u1_col_out_132    ),
    .col_out_133             ( u1_col_out_133    ),
    .col_out_134             ( u1_col_out_134    ),
    .col_out_135             ( u1_col_out_135    ),
    .col_out_136             ( u1_col_out_136    ),
    .col_out_137             ( u1_col_out_137    ),
    .col_out_138             ( u1_col_out_138    ),
    .col_out_139             ( u1_col_out_139    ),
    .col_out_140             ( u1_col_out_140    ),
    .col_out_141             ( u1_col_out_141    ),
    .col_out_142             ( u1_col_out_142    ),
    .col_out_143             ( u1_col_out_143    ),
    .col_out_144             ( u1_col_out_144    ),
    .col_out_145             ( u1_col_out_145    ),
    .col_out_146             ( u1_col_out_146    ),
    .col_out_147             ( u1_col_out_147    ),
    .col_out_148             ( u1_col_out_148    ),
    .col_out_149             ( u1_col_out_149    ),
    .col_out_150             ( u1_col_out_150    ),
    .col_out_151             ( u1_col_out_151    ),
    .col_out_152             ( u1_col_out_152    ),
    .col_out_153             ( u1_col_out_153    ),
    .col_out_154             ( u1_col_out_154    ),
    .col_out_155             ( u1_col_out_155    ),
    .col_out_156             ( u1_col_out_156    ),
    .col_out_157             ( u1_col_out_157    ),
    .col_out_158             ( u1_col_out_158    ),
    .col_out_159             ( u1_col_out_159    ),
    .col_out_160             ( u1_col_out_160    ),
    .col_out_161             ( u1_col_out_161    ),
    .col_out_162             ( u1_col_out_162    ),
    .col_out_163             ( u1_col_out_163    ),
    .col_out_164             ( u1_col_out_164    ),
    .col_out_165             ( u1_col_out_165    ),
    .col_out_166             ( u1_col_out_166    ),
    .col_out_167             ( u1_col_out_167    ),
    .col_out_168             ( u1_col_out_168    ),
    .col_out_169             ( u1_col_out_169    ),
    .col_out_170             ( u1_col_out_170    ),
    .col_out_171             ( u1_col_out_171    ),
    .col_out_172             ( u1_col_out_172    ),
    .col_out_173             ( u1_col_out_173    ),
    .col_out_174             ( u1_col_out_174    ),
    .col_out_175             ( u1_col_out_175    ),
    .col_out_176             ( u1_col_out_176    ),
    .col_out_177             ( u1_col_out_177    ),
    .col_out_178             ( u1_col_out_178    ),
    .col_out_179             ( u1_col_out_179    ),
    .col_out_180             ( u1_col_out_180    ),
    .col_out_181             ( u1_col_out_181    ),
    .col_out_182             ( u1_col_out_182    ),
    .col_out_183             ( u1_col_out_183    ),
    .col_out_184             ( u1_col_out_184    ),
    .col_out_185             ( u1_col_out_185    ),
    .col_out_186             ( u1_col_out_186    ),
    .col_out_187             ( u1_col_out_187    ),
    .col_out_188             ( u1_col_out_188    ),
    .col_out_189             ( u1_col_out_189    ),
    .col_out_190             ( u1_col_out_190    ),
    .col_out_191             ( u1_col_out_191    ),
    .col_out_192             ( u1_col_out_192    ),
    .col_out_193             ( u1_col_out_193    ),
    .col_out_194             ( u1_col_out_194    ),
    .col_out_195             ( u1_col_out_195    ),
    .col_out_196             ( u1_col_out_196    ),
    .col_out_197             ( u1_col_out_197    ),
    .col_out_198             ( u1_col_out_198    ),
    .col_out_199             ( u1_col_out_199    ),
    .col_out_200             ( u1_col_out_200    ),
    .col_out_201             ( u1_col_out_201    ),
    .col_out_202             ( u1_col_out_202    ),
    .col_out_203             ( u1_col_out_203    ),
    .col_out_204             ( u1_col_out_204    ),
    .col_out_205             ( u1_col_out_205    ),
    .col_out_206             ( u1_col_out_206    ),
    .col_out_207             ( u1_col_out_207    ),
    .col_out_208             ( u1_col_out_208    ),
    .col_out_209             ( u1_col_out_209    ),
    .col_out_210             ( u1_col_out_210    ),
    .col_out_211             ( u1_col_out_211    ),
    .col_out_212             ( u1_col_out_212    ),
    .col_out_213             ( u1_col_out_213    ),
    .col_out_214             ( u1_col_out_214    ),
    .col_out_215             ( u1_col_out_215    ),
    .col_out_216             ( u1_col_out_216    ),
    .col_out_217             ( u1_col_out_217    ),
    .col_out_218             ( u1_col_out_218    ),
    .col_out_219             ( u1_col_out_219    ),
    .col_out_220             ( u1_col_out_220    ),
    .col_out_221             ( u1_col_out_221    ),
    .col_out_222             ( u1_col_out_222    ),
    .col_out_223             ( u1_col_out_223    ),
    .col_out_224             ( u1_col_out_224    ),
    .col_out_225             ( u1_col_out_225    ),
    .col_out_226             ( u1_col_out_226    ),
    .col_out_227             ( u1_col_out_227    ),
    .col_out_228             ( u1_col_out_228    ),
    .col_out_229             ( u1_col_out_229    ),
    .col_out_230             ( u1_col_out_230    ),
    .col_out_231             ( u1_col_out_231    ),
    .col_out_232             ( u1_col_out_232    ),
    .col_out_233             ( u1_col_out_233    ),
    .col_out_234             ( u1_col_out_234    ),
    .col_out_235             ( u1_col_out_235    ),
    .col_out_236             ( u1_col_out_236    ),
    .col_out_237             ( u1_col_out_237    ),
    .col_out_238             ( u1_col_out_238    ),
    .col_out_239             ( u1_col_out_239    ),
    .col_out_240             ( u1_col_out_240    ),
    .col_out_241             ( u1_col_out_241    ),
    .col_out_242             ( u1_col_out_242    ),
    .col_out_243             ( u1_col_out_243    ),
    .col_out_244             ( u1_col_out_244    ),
    .col_out_245             ( u1_col_out_245    ),
    .col_out_246             ( u1_col_out_246    ),
    .col_out_247             ( u1_col_out_247    ),
    .col_out_248             ( u1_col_out_248    ),
    .col_out_249             ( u1_col_out_249    ),
    .col_out_250             ( u1_col_out_250    ),
    .col_out_251             ( u1_col_out_251    ),
    .col_out_252             ( u1_col_out_252    ),
    .col_out_253             ( u1_col_out_253    ),
    .col_out_254             ( u1_col_out_254    ),
    .col_out_255             ( u1_col_out_255    ),
    .col_out_256             ( u1_col_out_256    ),
    .col_out_257             ( u1_col_out_257    ),
    .col_out_258             ( u1_col_out_258    ),
    .col_out_259             ( u1_col_out_259    ),
    .col_out_260             ( u1_col_out_260    ),
    .col_out_261             ( u1_col_out_261    ),
    .col_out_262             ( u1_col_out_262    ),
    .col_out_263             ( u1_col_out_263    ),
    .col_out_264             ( u1_col_out_264    ),
    .col_out_265             ( u1_col_out_265    ),
    .col_out_266             ( u1_col_out_266    ),
    .col_out_267             ( u1_col_out_267    ),
    .col_out_268             ( u1_col_out_268    ),
    .col_out_269             ( u1_col_out_269    ),
    .col_out_270             ( u1_col_out_270    ),
    .col_out_271             ( u1_col_out_271    ),
    .col_out_272             ( u1_col_out_272    ),
    .col_out_273             ( u1_col_out_273    ),
    .col_out_274             ( u1_col_out_274    ),
    .col_out_275             ( u1_col_out_275    ),
    .col_out_276             ( u1_col_out_276    ),
    .col_out_277             ( u1_col_out_277    ),
    .col_out_278             ( u1_col_out_278    ),
    .col_out_279             ( u1_col_out_279    ),
    .col_out_280             ( u1_col_out_280    ),
    .col_out_281             ( u1_col_out_281    ),
    .col_out_282             ( u1_col_out_282    ),
    .col_out_283             ( u1_col_out_283    ),
    .col_out_284             ( u1_col_out_284    ),
    .col_out_285             ( u1_col_out_285    ),
    .col_out_286             ( u1_col_out_286    ),
    .col_out_287             ( u1_col_out_287    ),
    .col_out_288             ( u1_col_out_288    ),
    .col_out_289             ( u1_col_out_289    ),
    .col_out_290             ( u1_col_out_290    ),
    .col_out_291             ( u1_col_out_291    ),
    .col_out_292             ( u1_col_out_292    ),
    .col_out_293             ( u1_col_out_293    ),
    .col_out_294             ( u1_col_out_294    ),
    .col_out_295             ( u1_col_out_295    ),
    .col_out_296             ( u1_col_out_296    ),
    .col_out_297             ( u1_col_out_297    ),
    .col_out_298             ( u1_col_out_298    ),
    .col_out_299             ( u1_col_out_299    ),
    .col_out_300             ( u1_col_out_300    ),
    .col_out_301             ( u1_col_out_301    ),
    .col_out_302             ( u1_col_out_302    ),
    .col_out_303             ( u1_col_out_303    ),
    .col_out_304             ( u1_col_out_304    ),
    .col_out_305             ( u1_col_out_305    ),
    .col_out_306             ( u1_col_out_306    ),
    .col_out_307             ( u1_col_out_307    ),
    .col_out_308             ( u1_col_out_308    ),
    .col_out_309             ( u1_col_out_309    ),
    .col_out_310             ( u1_col_out_310    ),
    .col_out_311             ( u1_col_out_311    ),
    .col_out_312             ( u1_col_out_312    ),
    .col_out_313             ( u1_col_out_313    ),
    .col_out_314             ( u1_col_out_314    ),
    .col_out_315             ( u1_col_out_315    ),
    .col_out_316             ( u1_col_out_316    ),
    .col_out_317             ( u1_col_out_317    ),
    .col_out_318             ( u1_col_out_318    ),
    .col_out_319             ( u1_col_out_319    ),
    .col_out_320             ( u1_col_out_320    ),
    .col_out_321             ( u1_col_out_321    ),
    .col_out_322             ( u1_col_out_322    ),
    .col_out_323             ( u1_col_out_323    ),
    .col_out_324             ( u1_col_out_324    ),
    .col_out_325             ( u1_col_out_325    ),
    .col_out_326             ( u1_col_out_326    ),
    .col_out_327             ( u1_col_out_327    ),
    .col_out_328             ( u1_col_out_328    ),
    .col_out_329             ( u1_col_out_329    ),
    .col_out_330             ( u1_col_out_330    ),
    .col_out_331             ( u1_col_out_331    ),
    .col_out_332             ( u1_col_out_332    ),
    .col_out_333             ( u1_col_out_333    ),
    .col_out_334             ( u1_col_out_334    ),
    .col_out_335             ( u1_col_out_335    ),
    .col_out_336             ( u1_col_out_336    ),
    .col_out_337             ( u1_col_out_337    ),
    .col_out_338             ( u1_col_out_338    ),
    .col_out_339             ( u1_col_out_339    ),
    .col_out_340             ( u1_col_out_340    ),
    .col_out_341             ( u1_col_out_341    ),
    .col_out_342             ( u1_col_out_342    ),
    .col_out_343             ( u1_col_out_343    ),
    .col_out_344             ( u1_col_out_344    ),
    .col_out_345             ( u1_col_out_345    ),
    .col_out_346             ( u1_col_out_346    ),
    .col_out_347             ( u1_col_out_347    ),
    .col_out_348             ( u1_col_out_348    ),
    .col_out_349             ( u1_col_out_349    ),
    .col_out_350             ( u1_col_out_350    ),
    .col_out_351             ( u1_col_out_351    ),
    .col_out_352             ( u1_col_out_352    ),
    .col_out_353             ( u1_col_out_353    ),
    .col_out_354             ( u1_col_out_354    ),
    .col_out_355             ( u1_col_out_355    ),
    .col_out_356             ( u1_col_out_356    ),
    .col_out_357             ( u1_col_out_357    ),
    .col_out_358             ( u1_col_out_358    ),
    .col_out_359             ( u1_col_out_359    ),
    .col_out_360             ( u1_col_out_360    ),
    .col_out_361             ( u1_col_out_361    ),
    .col_out_362             ( u1_col_out_362    ),
    .col_out_363             ( u1_col_out_363    ),
    .col_out_364             ( u1_col_out_364    ),
    .col_out_365             ( u1_col_out_365    ),
    .col_out_366             ( u1_col_out_366    ),
    .col_out_367             ( u1_col_out_367    ),
    .col_out_368             ( u1_col_out_368    ),
    .col_out_369             ( u1_col_out_369    ),
    .col_out_370             ( u1_col_out_370    ),
    .col_out_371             ( u1_col_out_371    ),
    .col_out_372             ( u1_col_out_372    ),
    .col_out_373             ( u1_col_out_373    ),
    .col_out_374             ( u1_col_out_374    ),
    .col_out_375             ( u1_col_out_375    ),
    .col_out_376             ( u1_col_out_376    ),
    .col_out_377             ( u1_col_out_377    ),
    .col_out_378             ( u1_col_out_378    ),
    .col_out_379             ( u1_col_out_379    ),
    .col_out_380             ( u1_col_out_380    ),
    .col_out_381             ( u1_col_out_381    ),
    .col_out_382             ( u1_col_out_382    ),
    .col_out_383             ( u1_col_out_383    ),
    .col_out_384             ( u1_col_out_384    ),
    .col_out_385             ( u1_col_out_385    ),
    .col_out_386             ( u1_col_out_386    ),
    .col_out_387             ( u1_col_out_387    ),
    .col_out_388             ( u1_col_out_388    ),
    .col_out_389             ( u1_col_out_389    ),
    .col_out_390             ( u1_col_out_390    ),
    .col_out_391             ( u1_col_out_391    ),
    .col_out_392             ( u1_col_out_392    ),
    .col_out_393             ( u1_col_out_393    ),
    .col_out_394             ( u1_col_out_394    ),
    .col_out_395             ( u1_col_out_395    ),
    .col_out_396             ( u1_col_out_396    ),
    .col_out_397             ( u1_col_out_397    ),
    .col_out_398             ( u1_col_out_398    ),
    .col_out_399             ( u1_col_out_399    ),
    .col_out_400             ( u1_col_out_400    ),
    .col_out_401             ( u1_col_out_401    ),
    .col_out_402             ( u1_col_out_402    ),
    .col_out_403             ( u1_col_out_403    ),
    .col_out_404             ( u1_col_out_404    ),
    .col_out_405             ( u1_col_out_405    ),
    .col_out_406             ( u1_col_out_406    ),
    .col_out_407             ( u1_col_out_407    ),
    .col_out_408             ( u1_col_out_408    ),
    .col_out_409             ( u1_col_out_409    ),
    .col_out_410             ( u1_col_out_410    ),
    .col_out_411             ( u1_col_out_411    ),
    .col_out_412             ( u1_col_out_412    ),
    .col_out_413             ( u1_col_out_413    ),
    .col_out_414             ( u1_col_out_414    ),
    .col_out_415             ( u1_col_out_415    ),
    .col_out_416             ( u1_col_out_416    ),
    .col_out_417             ( u1_col_out_417    ),
    .col_out_418             ( u1_col_out_418    ),
    .col_out_419             ( u1_col_out_419    ),
    .col_out_420             ( u1_col_out_420    ),
    .col_out_421             ( u1_col_out_421    ),
    .col_out_422             ( u1_col_out_422    ),
    .col_out_423             ( u1_col_out_423    ),
    .col_out_424             ( u1_col_out_424    ),
    .col_out_425             ( u1_col_out_425    ),
    .col_out_426             ( u1_col_out_426    ),
    .col_out_427             ( u1_col_out_427    ),
    .col_out_428             ( u1_col_out_428    ),
    .col_out_429             ( u1_col_out_429    ),
    .col_out_430             ( u1_col_out_430    ),
    .col_out_431             ( u1_col_out_431    ),
    .col_out_432             ( u1_col_out_432    ),
    .col_out_433             ( u1_col_out_433    ),
    .col_out_434             ( u1_col_out_434    ),
    .col_out_435             ( u1_col_out_435    ),
    .col_out_436             ( u1_col_out_436    ),
    .col_out_437             ( u1_col_out_437    ),
    .col_out_438             ( u1_col_out_438    ),
    .col_out_439             ( u1_col_out_439    ),
    .col_out_440             ( u1_col_out_440    ),
    .col_out_441             ( u1_col_out_441    ),
    .col_out_442             ( u1_col_out_442    ),
    .col_out_443             ( u1_col_out_443    ),
    .col_out_444             ( u1_col_out_444    ),
    .col_out_445             ( u1_col_out_445    ),
    .col_out_446             ( u1_col_out_446    ),
    .col_out_447             ( u1_col_out_447    ),
    .col_out_448             ( u1_col_out_448    ),
    .col_out_449             ( u1_col_out_449    ),
    .col_out_450             ( u1_col_out_450    ),
    .col_out_451             ( u1_col_out_451    ),
    .col_out_452             ( u1_col_out_452    ),
    .col_out_453             ( u1_col_out_453    ),
    .col_out_454             ( u1_col_out_454    ),
    .col_out_455             ( u1_col_out_455    ),
    .col_out_456             ( u1_col_out_456    ),
    .col_out_457             ( u1_col_out_457    ),
    .col_out_458             ( u1_col_out_458    ),
    .col_out_459             ( u1_col_out_459    ),
    .col_out_460             ( u1_col_out_460    ),
    .col_out_461             ( u1_col_out_461    ),
    .col_out_462             ( u1_col_out_462    ),
    .col_out_463             ( u1_col_out_463    ),
    .col_out_464             ( u1_col_out_464    ),
    .col_out_465             ( u1_col_out_465    ),
    .col_out_466             ( u1_col_out_466    ),
    .col_out_467             ( u1_col_out_467    ),
    .col_out_468             ( u1_col_out_468    ),
    .col_out_469             ( u1_col_out_469    ),
    .col_out_470             ( u1_col_out_470    ),
    .col_out_471             ( u1_col_out_471    ),
    .col_out_472             ( u1_col_out_472    ),
    .col_out_473             ( u1_col_out_473    ),
    .col_out_474             ( u1_col_out_474    ),
    .col_out_475             ( u1_col_out_475    ),
    .col_out_476             ( u1_col_out_476    ),
    .col_out_477             ( u1_col_out_477    ),
    .col_out_478             ( u1_col_out_478    ),
    .col_out_479             ( u1_col_out_479    ),
    .col_out_480             ( u1_col_out_480    ),
    .col_out_481             ( u1_col_out_481    ),
    .col_out_482             ( u1_col_out_482    ),
    .col_out_483             ( u1_col_out_483    ),
    .col_out_484             ( u1_col_out_484    ),
    .col_out_485             ( u1_col_out_485    ),
    .col_out_486             ( u1_col_out_486    ),
    .col_out_487             ( u1_col_out_487    ),
    .col_out_488             ( u1_col_out_488    ),
    .col_out_489             ( u1_col_out_489    ),
    .col_out_490             ( u1_col_out_490    ),
    .col_out_491             ( u1_col_out_491    ),
    .col_out_492             ( u1_col_out_492    ),
    .col_out_493             ( u1_col_out_493    ),
    .col_out_494             ( u1_col_out_494    ),
    .col_out_495             ( u1_col_out_495    ),
    .col_out_496             ( u1_col_out_496    ),
    .col_out_497             ( u1_col_out_497    ),
    .col_out_498             ( u1_col_out_498    ),
    .col_out_499             ( u1_col_out_499    ),
    .col_out_500             ( u1_col_out_500    ),
    .col_out_501             ( u1_col_out_501    ),
    .col_out_502             ( u1_col_out_502    ),
    .col_out_503             ( u1_col_out_503    ),
    .col_out_504             ( u1_col_out_504    ),
    .col_out_505             ( u1_col_out_505    ),
    .col_out_506             ( u1_col_out_506    ),
    .col_out_507             ( u1_col_out_507    ),
    .col_out_508             ( u1_col_out_508    ),
    .col_out_509             ( u1_col_out_509    ),
    .col_out_510             ( u1_col_out_510    ),
    .col_out_511             ( u1_col_out_511    ),
    .col_out_512             ( u1_col_out_512    ),
    .col_out_513             ( u1_col_out_513    ),
    .col_out_514             ( u1_col_out_514    ),
    .col_out_515             ( u1_col_out_515    ),
    .col_out_516             ( u1_col_out_516    ),
    .col_out_517             ( u1_col_out_517    ),
    .col_out_518             ( u1_col_out_518    ),
    .col_out_519             ( u1_col_out_519    ),
    .col_out_520             ( u1_col_out_520    ),
    .col_out_521             ( u1_col_out_521    ),
    .col_out_522             ( u1_col_out_522    ),
    .col_out_523             ( u1_col_out_523    ),
    .col_out_524             ( u1_col_out_524    ),
    .col_out_525             ( u1_col_out_525    ),
    .col_out_526             ( u1_col_out_526    ),
    .col_out_527             ( u1_col_out_527    ),
    .col_out_528             ( u1_col_out_528    ),
    .col_out_529             ( u1_col_out_529    ),
    .col_out_530             ( u1_col_out_530    ),
    .col_out_531             ( u1_col_out_531    ),
    .col_out_532             ( u1_col_out_532    ),
    .col_out_533             ( u1_col_out_533    ),
    .col_out_534             ( u1_col_out_534    ),
    .col_out_535             ( u1_col_out_535    ),
    .col_out_536             ( u1_col_out_536    ),
    .col_out_537             ( u1_col_out_537    ),
    .col_out_538             ( u1_col_out_538    ),
    .col_out_539             ( u1_col_out_539    ),
    .col_out_540             ( u1_col_out_540    ),
    .col_out_541             ( u1_col_out_541    ),
    .col_out_542             ( u1_col_out_542    ),
    .col_out_543             ( u1_col_out_543    ),
    .col_out_544             ( u1_col_out_544    ),
    .col_out_545             ( u1_col_out_545    ),
    .col_out_546             ( u1_col_out_546    ),
    .col_out_547             ( u1_col_out_547    ),
    .col_out_548             ( u1_col_out_548    ),
    .col_out_549             ( u1_col_out_549    ),
    .col_out_550             ( u1_col_out_550    ),
    .col_out_551             ( u1_col_out_551    ),
    .col_out_552             ( u1_col_out_552    ),
    .col_out_553             ( u1_col_out_553    ),
    .col_out_554             ( u1_col_out_554    ),
    .col_out_555             ( u1_col_out_555    ),
    .col_out_556             ( u1_col_out_556    ),
    .col_out_557             ( u1_col_out_557    ),
    .col_out_558             ( u1_col_out_558    ),
    .col_out_559             ( u1_col_out_559    ),
    .col_out_560             ( u1_col_out_560    ),
    .col_out_561             ( u1_col_out_561    ),
    .col_out_562             ( u1_col_out_562    ),
    .col_out_563             ( u1_col_out_563    ),
    .col_out_564             ( u1_col_out_564    ),
    .col_out_565             ( u1_col_out_565    ),
    .col_out_566             ( u1_col_out_566    ),
    .col_out_567             ( u1_col_out_567    ),
    .col_out_568             ( u1_col_out_568    ),
    .col_out_569             ( u1_col_out_569    ),
    .col_out_570             ( u1_col_out_570    ),
    .col_out_571             ( u1_col_out_571    ),
    .col_out_572             ( u1_col_out_572    ),
    .col_out_573             ( u1_col_out_573    ),
    .col_out_574             ( u1_col_out_574    ),
    .col_out_575             ( u1_col_out_575    ),
    .col_out_576             ( u1_col_out_576    ),
    .col_out_577             ( u1_col_out_577    ),
    .col_out_578             ( u1_col_out_578    ),
    .col_out_579             ( u1_col_out_579    ),
    .col_out_580             ( u1_col_out_580    ),
    .col_out_581             ( u1_col_out_581    ),
    .col_out_582             ( u1_col_out_582    ),
    .col_out_583             ( u1_col_out_583    ),
    .col_out_584             ( u1_col_out_584    ),
    .col_out_585             ( u1_col_out_585    ),
    .col_out_586             ( u1_col_out_586    ),
    .col_out_587             ( u1_col_out_587    ),
    .col_out_588             ( u1_col_out_588    ),
    .col_out_589             ( u1_col_out_589    ),
    .col_out_590             ( u1_col_out_590    ),
    .col_out_591             ( u1_col_out_591    ),
    .col_out_592             ( u1_col_out_592    ),
    .col_out_593             ( u1_col_out_593    ),
    .col_out_594             ( u1_col_out_594    ),
    .col_out_595             ( u1_col_out_595    ),
    .col_out_596             ( u1_col_out_596    ),
    .col_out_597             ( u1_col_out_597    ),
    .col_out_598             ( u1_col_out_598    ),
    .col_out_599             ( u1_col_out_599    ),
    .col_out_600             ( u1_col_out_600    ),
    .col_out_601             ( u1_col_out_601    ),
    .col_out_602             ( u1_col_out_602    ),
    .col_out_603             ( u1_col_out_603    ),
    .col_out_604             ( u1_col_out_604    ),
    .col_out_605             ( u1_col_out_605    ),
    .col_out_606             ( u1_col_out_606    ),
    .col_out_607             ( u1_col_out_607    ),
    .col_out_608             ( u1_col_out_608    ),
    .col_out_609             ( u1_col_out_609    ),
    .col_out_610             ( u1_col_out_610    ),
    .col_out_611             ( u1_col_out_611    ),
    .col_out_612             ( u1_col_out_612    ),
    .col_out_613             ( u1_col_out_613    ),
    .col_out_614             ( u1_col_out_614    ),
    .col_out_615             ( u1_col_out_615    ),
    .col_out_616             ( u1_col_out_616    ),
    .col_out_617             ( u1_col_out_617    ),
    .col_out_618             ( u1_col_out_618    ),
    .col_out_619             ( u1_col_out_619    ),
    .col_out_620             ( u1_col_out_620    ),
    .col_out_621             ( u1_col_out_621    ),
    .col_out_622             ( u1_col_out_622    ),
    .col_out_623             ( u1_col_out_623    ),
    .col_out_624             ( u1_col_out_624    ),
    .col_out_625             ( u1_col_out_625    ),
    .col_out_626             ( u1_col_out_626    ),
    .col_out_627             ( u1_col_out_627    ),
    .col_out_628             ( u1_col_out_628    ),
    .col_out_629             ( u1_col_out_629    ),
    .col_out_630             ( u1_col_out_630    ),
    .col_out_631             ( u1_col_out_631    ),
    .col_out_632             ( u1_col_out_632    ),
    .col_out_633             ( u1_col_out_633    ),
    .col_out_634             ( u1_col_out_634    ),
    .col_out_635             ( u1_col_out_635    ),
    .col_out_636             ( u1_col_out_636    ),
    .col_out_637             ( u1_col_out_637    ),
    .col_out_638             ( u1_col_out_638    ),
    .col_out_639             ( u1_col_out_639    ),
    .col_out_640             ( u1_col_out_640    ),
    .col_out_641             ( u1_col_out_641    ),
    .col_out_642             ( u1_col_out_642    ),
    .col_out_643             ( u1_col_out_643    ),
    .col_out_644             ( u1_col_out_644    ),
    .col_out_645             ( u1_col_out_645    ),
    .col_out_646             ( u1_col_out_646    ),
    .col_out_647             ( u1_col_out_647    ),
    .col_out_648             ( u1_col_out_648    ),
    .col_out_649             ( u1_col_out_649    ),
    .col_out_650             ( u1_col_out_650    ),
    .col_out_651             ( u1_col_out_651    ),
    .col_out_652             ( u1_col_out_652    ),
    .col_out_653             ( u1_col_out_653    ),
    .col_out_654             ( u1_col_out_654    ),
    .col_out_655             ( u1_col_out_655    ),
    .col_out_656             ( u1_col_out_656    ),
    .col_out_657             ( u1_col_out_657    ),
    .col_out_658             ( u1_col_out_658    ),
    .col_out_659             ( u1_col_out_659    ),
    .col_out_660             ( u1_col_out_660    ),
    .col_out_661             ( u1_col_out_661    ),
    .col_out_662             ( u1_col_out_662    ),
    .col_out_663             ( u1_col_out_663    ),
    .col_out_664             ( u1_col_out_664    ),
    .col_out_665             ( u1_col_out_665    ),
    .col_out_666             ( u1_col_out_666    ),
    .col_out_667             ( u1_col_out_667    ),
    .col_out_668             ( u1_col_out_668    ),
    .col_out_669             ( u1_col_out_669    ),
    .col_out_670             ( u1_col_out_670    ),
    .col_out_671             ( u1_col_out_671    ),
    .col_out_672             ( u1_col_out_672    ),
    .col_out_673             ( u1_col_out_673    ),
    .col_out_674             ( u1_col_out_674    ),
    .col_out_675             ( u1_col_out_675    ),
    .col_out_676             ( u1_col_out_676    ),
    .col_out_677             ( u1_col_out_677    ),
    .col_out_678             ( u1_col_out_678    ),
    .col_out_679             ( u1_col_out_679    ),
    .col_out_680             ( u1_col_out_680    ),
    .col_out_681             ( u1_col_out_681    ),
    .col_out_682             ( u1_col_out_682    ),
    .col_out_683             ( u1_col_out_683    ),
    .col_out_684             ( u1_col_out_684    ),
    .col_out_685             ( u1_col_out_685    ),
    .col_out_686             ( u1_col_out_686    ),
    .col_out_687             ( u1_col_out_687    ),
    .col_out_688             ( u1_col_out_688    ),
    .col_out_689             ( u1_col_out_689    ),
    .col_out_690             ( u1_col_out_690    ),
    .col_out_691             ( u1_col_out_691    ),
    .col_out_692             ( u1_col_out_692    ),
    .col_out_693             ( u1_col_out_693    ),
    .col_out_694             ( u1_col_out_694    ),
    .col_out_695             ( u1_col_out_695    ),
    .col_out_696             ( u1_col_out_696    ),
    .col_out_697             ( u1_col_out_697    ),
    .col_out_698             ( u1_col_out_698    ),
    .col_out_699             ( u1_col_out_699    ),
    .col_out_700             ( u1_col_out_700    ),
    .col_out_701             ( u1_col_out_701    ),
    .col_out_702             ( u1_col_out_702    ),
    .col_out_703             ( u1_col_out_703    ),
    .col_out_704             ( u1_col_out_704    ),
    .col_out_705             ( u1_col_out_705    ),
    .col_out_706             ( u1_col_out_706    ),
    .col_out_707             ( u1_col_out_707    ),
    .col_out_708             ( u1_col_out_708    ),
    .col_out_709             ( u1_col_out_709    ),
    .col_out_710             ( u1_col_out_710    ),
    .col_out_711             ( u1_col_out_711    ),
    .col_out_712             ( u1_col_out_712    ),
    .col_out_713             ( u1_col_out_713    ),
    .col_out_714             ( u1_col_out_714    ),
    .col_out_715             ( u1_col_out_715    ),
    .col_out_716             ( u1_col_out_716    ),
    .col_out_717             ( u1_col_out_717    ),
    .col_out_718             ( u1_col_out_718    ),
    .col_out_719             ( u1_col_out_719    ),
    .col_out_720             ( u1_col_out_720    ),
    .col_out_721             ( u1_col_out_721    ),
    .col_out_722             ( u1_col_out_722    ),
    .col_out_723             ( u1_col_out_723    ),
    .col_out_724             ( u1_col_out_724    ),
    .col_out_725             ( u1_col_out_725    ),
    .col_out_726             ( u1_col_out_726    ),
    .col_out_727             ( u1_col_out_727    ),
    .col_out_728             ( u1_col_out_728    ),
    .col_out_729             ( u1_col_out_729    ),
    .col_out_730             ( u1_col_out_730    ),
    .col_out_731             ( u1_col_out_731    ),
    .col_out_732             ( u1_col_out_732    ),
    .col_out_733             ( u1_col_out_733    ),
    .col_out_734             ( u1_col_out_734    ),
    .col_out_735             ( u1_col_out_735    ),
    .col_out_736             ( u1_col_out_736    ),
    .col_out_737             ( u1_col_out_737    ),
    .col_out_738             ( u1_col_out_738    ),
    .col_out_739             ( u1_col_out_739    ),
    .col_out_740             ( u1_col_out_740    ),
    .col_out_741             ( u1_col_out_741    ),
    .col_out_742             ( u1_col_out_742    ),
    .col_out_743             ( u1_col_out_743    ),
    .col_out_744             ( u1_col_out_744    ),
    .col_out_745             ( u1_col_out_745    ),
    .col_out_746             ( u1_col_out_746    ),
    .col_out_747             ( u1_col_out_747    ),
    .col_out_748             ( u1_col_out_748    ),
    .col_out_749             ( u1_col_out_749    ),
    .col_out_750             ( u1_col_out_750    ),
    .col_out_751             ( u1_col_out_751    ),
    .col_out_752             ( u1_col_out_752    ),
    .col_out_753             ( u1_col_out_753    ),
    .col_out_754             ( u1_col_out_754    ),
    .col_out_755             ( u1_col_out_755    ),
    .col_out_756             ( u1_col_out_756    ),
    .col_out_757             ( u1_col_out_757    ),
    .col_out_758             ( u1_col_out_758    ),
    .col_out_759             ( u1_col_out_759    ),
    .col_out_760             ( u1_col_out_760    ),
    .col_out_761             ( u1_col_out_761    ),
    .col_out_762             ( u1_col_out_762    ),
    .col_out_763             ( u1_col_out_763    ),
    .col_out_764             ( u1_col_out_764    ),
    .col_out_765             ( u1_col_out_765    ),
    .col_out_766             ( u1_col_out_766    ),
    .col_out_767             ( u1_col_out_767    ),
    .col_out_768             ( u1_col_out_768    ),
    .col_out_769             ( u1_col_out_769    ),
    .col_out_770             ( u1_col_out_770    ),
    .col_out_771             ( u1_col_out_771    ),
    .col_out_772             ( u1_col_out_772    ),
    .col_out_773             ( u1_col_out_773    ),
    .col_out_774             ( u1_col_out_774    ),
    .col_out_775             ( u1_col_out_775    ),
    .col_out_776             ( u1_col_out_776    ),
    .col_out_777             ( u1_col_out_777    ),
    .col_out_778             ( u1_col_out_778    ),
    .col_out_779             ( u1_col_out_779    ),
    .col_out_780             ( u1_col_out_780    ),
    .col_out_781             ( u1_col_out_781    ),
    .col_out_782             ( u1_col_out_782    ),
    .col_out_783             ( u1_col_out_783    ),
    .col_out_784             ( u1_col_out_784    ),
    .col_out_785             ( u1_col_out_785    ),
    .col_out_786             ( u1_col_out_786    ),
    .col_out_787             ( u1_col_out_787    ),
    .col_out_788             ( u1_col_out_788    ),
    .col_out_789             ( u1_col_out_789    ),
    .col_out_790             ( u1_col_out_790    ),
    .col_out_791             ( u1_col_out_791    ),
    .col_out_792             ( u1_col_out_792    ),
    .col_out_793             ( u1_col_out_793    ),
    .col_out_794             ( u1_col_out_794    ),
    .col_out_795             ( u1_col_out_795    ),
    .col_out_796             ( u1_col_out_796    ),
    .col_out_797             ( u1_col_out_797    ),
    .col_out_798             ( u1_col_out_798    ),
    .col_out_799             ( u1_col_out_799    ),
    .col_out_800             ( u1_col_out_800    ),
    .col_out_801             ( u1_col_out_801    ),
    .col_out_802             ( u1_col_out_802    ),
    .col_out_803             ( u1_col_out_803    ),
    .col_out_804             ( u1_col_out_804    ),
    .col_out_805             ( u1_col_out_805    ),
    .col_out_806             ( u1_col_out_806    ),
    .col_out_807             ( u1_col_out_807    ),
    .col_out_808             ( u1_col_out_808    ),
    .col_out_809             ( u1_col_out_809    ),
    .col_out_810             ( u1_col_out_810    ),
    .col_out_811             ( u1_col_out_811    ),
    .col_out_812             ( u1_col_out_812    ),
    .col_out_813             ( u1_col_out_813    ),
    .col_out_814             ( u1_col_out_814    ),
    .col_out_815             ( u1_col_out_815    ),
    .col_out_816             ( u1_col_out_816    ),
    .col_out_817             ( u1_col_out_817    ),
    .col_out_818             ( u1_col_out_818    ),
    .col_out_819             ( u1_col_out_819    ),
    .col_out_820             ( u1_col_out_820    ),
    .col_out_821             ( u1_col_out_821    ),
    .col_out_822             ( u1_col_out_822    ),
    .col_out_823             ( u1_col_out_823    ),
    .col_out_824             ( u1_col_out_824    ),
    .col_out_825             ( u1_col_out_825    ),
    .col_out_826             ( u1_col_out_826    ),
    .col_out_827             ( u1_col_out_827    ),
    .col_out_828             ( u1_col_out_828    ),
    .col_out_829             ( u1_col_out_829    ),
    .col_out_830             ( u1_col_out_830    ),
    .col_out_831             ( u1_col_out_831    ),
    .col_out_832             ( u1_col_out_832    ),
    .col_out_833             ( u1_col_out_833    ),
    .col_out_834             ( u1_col_out_834    ),
    .col_out_835             ( u1_col_out_835    ),
    .col_out_836             ( u1_col_out_836    ),
    .col_out_837             ( u1_col_out_837    ),
    .col_out_838             ( u1_col_out_838    ),
    .col_out_839             ( u1_col_out_839    ),
    .col_out_840             ( u1_col_out_840    ),
    .col_out_841             ( u1_col_out_841    ),
    .col_out_842             ( u1_col_out_842    ),
    .col_out_843             ( u1_col_out_843    ),
    .col_out_844             ( u1_col_out_844    ),
    .col_out_845             ( u1_col_out_845    ),
    .col_out_846             ( u1_col_out_846    ),
    .col_out_847             ( u1_col_out_847    ),
    .col_out_848             ( u1_col_out_848    ),
    .col_out_849             ( u1_col_out_849    ),
    .col_out_850             ( u1_col_out_850    ),
    .col_out_851             ( u1_col_out_851    ),
    .col_out_852             ( u1_col_out_852    ),
    .col_out_853             ( u1_col_out_853    ),
    .col_out_854             ( u1_col_out_854    ),
    .col_out_855             ( u1_col_out_855    ),
    .col_out_856             ( u1_col_out_856    ),
    .col_out_857             ( u1_col_out_857    ),
    .col_out_858             ( u1_col_out_858    ),
    .col_out_859             ( u1_col_out_859    ),
    .col_out_860             ( u1_col_out_860    ),
    .col_out_861             ( u1_col_out_861    ),
    .col_out_862             ( u1_col_out_862    ),
    .col_out_863             ( u1_col_out_863    ),
    .col_out_864             ( u1_col_out_864    ),
    .col_out_865             ( u1_col_out_865    ),
    .col_out_866             ( u1_col_out_866    ),
    .col_out_867             ( u1_col_out_867    ),
    .col_out_868             ( u1_col_out_868    ),
    .col_out_869             ( u1_col_out_869    ),
    .col_out_870             ( u1_col_out_870    ),
    .col_out_871             ( u1_col_out_871    ),
    .col_out_872             ( u1_col_out_872    ),
    .col_out_873             ( u1_col_out_873    ),
    .col_out_874             ( u1_col_out_874    ),
    .col_out_875             ( u1_col_out_875    ),
    .col_out_876             ( u1_col_out_876    ),
    .col_out_877             ( u1_col_out_877    ),
    .col_out_878             ( u1_col_out_878    ),
    .col_out_879             ( u1_col_out_879    ),
    .col_out_880             ( u1_col_out_880    ),
    .col_out_881             ( u1_col_out_881    ),
    .col_out_882             ( u1_col_out_882    ),
    .col_out_883             ( u1_col_out_883    ),
    .col_out_884             ( u1_col_out_884    ),
    .col_out_885             ( u1_col_out_885    ),
    .col_out_886             ( u1_col_out_886    ),
    .col_out_887             ( u1_col_out_887    ),
    .col_out_888             ( u1_col_out_888    ),
    .col_out_889             ( u1_col_out_889    ),
    .col_out_890             ( u1_col_out_890    ),
    .col_out_891             ( u1_col_out_891    ),
    .col_out_892             ( u1_col_out_892    ),
    .col_out_893             ( u1_col_out_893    ),
    .col_out_894             ( u1_col_out_894    ),
    .col_out_895             ( u1_col_out_895    ),
    .col_out_896             ( u1_col_out_896    ),
    .col_out_897             ( u1_col_out_897    ),
    .col_out_898             ( u1_col_out_898    ),
    .col_out_899             ( u1_col_out_899    ),
    .col_out_900             ( u1_col_out_900    ),
    .col_out_901             ( u1_col_out_901    ),
    .col_out_902             ( u1_col_out_902    ),
    .col_out_903             ( u1_col_out_903    ),
    .col_out_904             ( u1_col_out_904    ),
    .col_out_905             ( u1_col_out_905    ),
    .col_out_906             ( u1_col_out_906    ),
    .col_out_907             ( u1_col_out_907    ),
    .col_out_908             ( u1_col_out_908    ),
    .col_out_909             ( u1_col_out_909    ),
    .col_out_910             ( u1_col_out_910    ),
    .col_out_911             ( u1_col_out_911    ),
    .col_out_912             ( u1_col_out_912    ),
    .col_out_913             ( u1_col_out_913    ),
    .col_out_914             ( u1_col_out_914    ),
    .col_out_915             ( u1_col_out_915    ),
    .col_out_916             ( u1_col_out_916    ),
    .col_out_917             ( u1_col_out_917    ),
    .col_out_918             ( u1_col_out_918    ),
    .col_out_919             ( u1_col_out_919    ),
    .col_out_920             ( u1_col_out_920    ),
    .col_out_921             ( u1_col_out_921    ),
    .col_out_922             ( u1_col_out_922    ),
    .col_out_923             ( u1_col_out_923    ),
    .col_out_924             ( u1_col_out_924    ),
    .col_out_925             ( u1_col_out_925    ),
    .col_out_926             ( u1_col_out_926    ),
    .col_out_927             ( u1_col_out_927    ),
    .col_out_928             ( u1_col_out_928    ),
    .col_out_929             ( u1_col_out_929    ),
    .col_out_930             ( u1_col_out_930    ),
    .col_out_931             ( u1_col_out_931    ),
    .col_out_932             ( u1_col_out_932    ),
    .col_out_933             ( u1_col_out_933    ),
    .col_out_934             ( u1_col_out_934    ),
    .col_out_935             ( u1_col_out_935    ),
    .col_out_936             ( u1_col_out_936    ),
    .col_out_937             ( u1_col_out_937    ),
    .col_out_938             ( u1_col_out_938    ),
    .col_out_939             ( u1_col_out_939    ),
    .col_out_940             ( u1_col_out_940    ),
    .col_out_941             ( u1_col_out_941    ),
    .col_out_942             ( u1_col_out_942    ),
    .col_out_943             ( u1_col_out_943    ),
    .col_out_944             ( u1_col_out_944    ),
    .col_out_945             ( u1_col_out_945    ),
    .col_out_946             ( u1_col_out_946    ),
    .col_out_947             ( u1_col_out_947    ),
    .col_out_948             ( u1_col_out_948    ),
    .col_out_949             ( u1_col_out_949    ),
    .col_out_950             ( u1_col_out_950    ),
    .col_out_951             ( u1_col_out_951    ),
    .col_out_952             ( u1_col_out_952    ),
    .col_out_953             ( u1_col_out_953    ),
    .col_out_954             ( u1_col_out_954    ),
    .col_out_955             ( u1_col_out_955    ),
    .col_out_956             ( u1_col_out_956    ),
    .col_out_957             ( u1_col_out_957    ),
    .col_out_958             ( u1_col_out_958    ),
    .col_out_959             ( u1_col_out_959    ),
    .col_out_960             ( u1_col_out_960    ),
    .col_out_961             ( u1_col_out_961    ),
    .col_out_962             ( u1_col_out_962    ),
    .col_out_963             ( u1_col_out_963    ),
    .col_out_964             ( u1_col_out_964    ),
    .col_out_965             ( u1_col_out_965    ),
    .col_out_966             ( u1_col_out_966    ),
    .col_out_967             ( u1_col_out_967    ),
    .col_out_968             ( u1_col_out_968    ),
    .col_out_969             ( u1_col_out_969    ),
    .col_out_970             ( u1_col_out_970    ),
    .col_out_971             ( u1_col_out_971    ),
    .col_out_972             ( u1_col_out_972    ),
    .col_out_973             ( u1_col_out_973    ),
    .col_out_974             ( u1_col_out_974    ),
    .col_out_975             ( u1_col_out_975    ),
    .col_out_976             ( u1_col_out_976    ),
    .col_out_977             ( u1_col_out_977    ),
    .col_out_978             ( u1_col_out_978    ),
    .col_out_979             ( u1_col_out_979    ),
    .col_out_980             ( u1_col_out_980    ),
    .col_out_981             ( u1_col_out_981    ),
    .col_out_982             ( u1_col_out_982    ),
    .col_out_983             ( u1_col_out_983    ),
    .col_out_984             ( u1_col_out_984    ),
    .col_out_985             ( u1_col_out_985    ),
    .col_out_986             ( u1_col_out_986    ),
    .col_out_987             ( u1_col_out_987    ),
    .col_out_988             ( u1_col_out_988    ),
    .col_out_989             ( u1_col_out_989    ),
    .col_out_990             ( u1_col_out_990    ),
    .col_out_991             ( u1_col_out_991    ),
    .col_out_992             ( u1_col_out_992    ),
    .col_out_993             ( u1_col_out_993    ),
    .col_out_994             ( u1_col_out_994    ),
    .col_out_995             ( u1_col_out_995    ),
    .col_out_996             ( u1_col_out_996    ),
    .col_out_997             ( u1_col_out_997    ),
    .col_out_998             ( u1_col_out_998    ),
    .col_out_999             ( u1_col_out_999    ),
    .col_out_1000            ( u1_col_out_1000   ),
    .col_out_1001            ( u1_col_out_1001   ),
    .col_out_1002            ( u1_col_out_1002   ),
    .col_out_1003            ( u1_col_out_1003   ),
    .col_out_1004            ( u1_col_out_1004   ),
    .col_out_1005            ( u1_col_out_1005   ),
    .col_out_1006            ( u1_col_out_1006   ),
    .col_out_1007            ( u1_col_out_1007   ),
    .col_out_1008            ( u1_col_out_1008   ),
    .col_out_1009            ( u1_col_out_1009   ),
    .col_out_1010            ( u1_col_out_1010   ),
    .col_out_1011            ( u1_col_out_1011   ),
    .col_out_1012            ( u1_col_out_1012   ),
    .col_out_1013            ( u1_col_out_1013   ),
    .col_out_1014            ( u1_col_out_1014   ),
    .col_out_1015            ( u1_col_out_1015   ),
    .col_out_1016            ( u1_col_out_1016   ),
    .col_out_1017            ( u1_col_out_1017   ),
    .col_out_1018            ( u1_col_out_1018   ),
    .col_out_1019            ( u1_col_out_1019   ),
    .col_out_1020            ( u1_col_out_1020   ),
    .col_out_1021            ( u1_col_out_1021   ),
    .col_out_1022            ( u1_col_out_1022   ),
    .col_out_1023            ( u1_col_out_1023   ),
    .col_out_1024            ( u1_col_out_1024   ),
    .col_out_1025            ( u1_col_out_1025   ),
    .col_out_1026            ( u1_col_out_1026   ),
    .col_out_1027            ( u1_col_out_1027   ),
    .col_out_1028            ( u1_col_out_1028   ),
    .col_out_1029            ( u1_col_out_1029   ),
    .col_out_1030            ( u1_col_out_1030   ),
    .col_out_1031            ( u1_col_out_1031   ),
    .col_out_1032            ( u1_col_out_1032   ),
    .col_out_1033            ( u1_col_out_1033   )
);


























// compressor_array_8_6_1033 Outputs
wire  [5:0]  u2_col_out_0;
wire  [5:0]  u2_col_out_1;
wire  [5:0]  u2_col_out_2;
wire  [5:0]  u2_col_out_3;
wire  [5:0]  u2_col_out_4;
wire  [5:0]  u2_col_out_5;
wire  [5:0]  u2_col_out_6;
wire  [5:0]  u2_col_out_7;
wire  [5:0]  u2_col_out_8;
wire  [5:0]  u2_col_out_9;
wire  [5:0]  u2_col_out_10;
wire  [5:0]  u2_col_out_11;
wire  [5:0]  u2_col_out_12;
wire  [5:0]  u2_col_out_13;
wire  [5:0]  u2_col_out_14;
wire  [5:0]  u2_col_out_15;
wire  [5:0]  u2_col_out_16;
wire  [5:0]  u2_col_out_17;
wire  [5:0]  u2_col_out_18;
wire  [5:0]  u2_col_out_19;
wire  [5:0]  u2_col_out_20;
wire  [5:0]  u2_col_out_21;
wire  [5:0]  u2_col_out_22;
wire  [5:0]  u2_col_out_23;
wire  [5:0]  u2_col_out_24;
wire  [5:0]  u2_col_out_25;
wire  [5:0]  u2_col_out_26;
wire  [5:0]  u2_col_out_27;
wire  [5:0]  u2_col_out_28;
wire  [5:0]  u2_col_out_29;
wire  [5:0]  u2_col_out_30;
wire  [5:0]  u2_col_out_31;
wire  [5:0]  u2_col_out_32;
wire  [5:0]  u2_col_out_33;
wire  [5:0]  u2_col_out_34;
wire  [5:0]  u2_col_out_35;
wire  [5:0]  u2_col_out_36;
wire  [5:0]  u2_col_out_37;
wire  [5:0]  u2_col_out_38;
wire  [5:0]  u2_col_out_39;
wire  [5:0]  u2_col_out_40;
wire  [5:0]  u2_col_out_41;
wire  [5:0]  u2_col_out_42;
wire  [5:0]  u2_col_out_43;
wire  [5:0]  u2_col_out_44;
wire  [5:0]  u2_col_out_45;
wire  [5:0]  u2_col_out_46;
wire  [5:0]  u2_col_out_47;
wire  [5:0]  u2_col_out_48;
wire  [5:0]  u2_col_out_49;
wire  [5:0]  u2_col_out_50;
wire  [5:0]  u2_col_out_51;
wire  [5:0]  u2_col_out_52;
wire  [5:0]  u2_col_out_53;
wire  [5:0]  u2_col_out_54;
wire  [5:0]  u2_col_out_55;
wire  [5:0]  u2_col_out_56;
wire  [5:0]  u2_col_out_57;
wire  [5:0]  u2_col_out_58;
wire  [5:0]  u2_col_out_59;
wire  [5:0]  u2_col_out_60;
wire  [5:0]  u2_col_out_61;
wire  [5:0]  u2_col_out_62;
wire  [5:0]  u2_col_out_63;
wire  [5:0]  u2_col_out_64;
wire  [5:0]  u2_col_out_65;
wire  [5:0]  u2_col_out_66;
wire  [5:0]  u2_col_out_67;
wire  [5:0]  u2_col_out_68;
wire  [5:0]  u2_col_out_69;
wire  [5:0]  u2_col_out_70;
wire  [5:0]  u2_col_out_71;
wire  [5:0]  u2_col_out_72;
wire  [5:0]  u2_col_out_73;
wire  [5:0]  u2_col_out_74;
wire  [5:0]  u2_col_out_75;
wire  [5:0]  u2_col_out_76;
wire  [5:0]  u2_col_out_77;
wire  [5:0]  u2_col_out_78;
wire  [5:0]  u2_col_out_79;
wire  [5:0]  u2_col_out_80;
wire  [5:0]  u2_col_out_81;
wire  [5:0]  u2_col_out_82;
wire  [5:0]  u2_col_out_83;
wire  [5:0]  u2_col_out_84;
wire  [5:0]  u2_col_out_85;
wire  [5:0]  u2_col_out_86;
wire  [5:0]  u2_col_out_87;
wire  [5:0]  u2_col_out_88;
wire  [5:0]  u2_col_out_89;
wire  [5:0]  u2_col_out_90;
wire  [5:0]  u2_col_out_91;
wire  [5:0]  u2_col_out_92;
wire  [5:0]  u2_col_out_93;
wire  [5:0]  u2_col_out_94;
wire  [5:0]  u2_col_out_95;
wire  [5:0]  u2_col_out_96;
wire  [5:0]  u2_col_out_97;
wire  [5:0]  u2_col_out_98;
wire  [5:0]  u2_col_out_99;
wire  [5:0]  u2_col_out_100;
wire  [5:0]  u2_col_out_101;
wire  [5:0]  u2_col_out_102;
wire  [5:0]  u2_col_out_103;
wire  [5:0]  u2_col_out_104;
wire  [5:0]  u2_col_out_105;
wire  [5:0]  u2_col_out_106;
wire  [5:0]  u2_col_out_107;
wire  [5:0]  u2_col_out_108;
wire  [5:0]  u2_col_out_109;
wire  [5:0]  u2_col_out_110;
wire  [5:0]  u2_col_out_111;
wire  [5:0]  u2_col_out_112;
wire  [5:0]  u2_col_out_113;
wire  [5:0]  u2_col_out_114;
wire  [5:0]  u2_col_out_115;
wire  [5:0]  u2_col_out_116;
wire  [5:0]  u2_col_out_117;
wire  [5:0]  u2_col_out_118;
wire  [5:0]  u2_col_out_119;
wire  [5:0]  u2_col_out_120;
wire  [5:0]  u2_col_out_121;
wire  [5:0]  u2_col_out_122;
wire  [5:0]  u2_col_out_123;
wire  [5:0]  u2_col_out_124;
wire  [5:0]  u2_col_out_125;
wire  [5:0]  u2_col_out_126;
wire  [5:0]  u2_col_out_127;
wire  [5:0]  u2_col_out_128;
wire  [5:0]  u2_col_out_129;
wire  [5:0]  u2_col_out_130;
wire  [5:0]  u2_col_out_131;
wire  [5:0]  u2_col_out_132;
wire  [5:0]  u2_col_out_133;
wire  [5:0]  u2_col_out_134;
wire  [5:0]  u2_col_out_135;
wire  [5:0]  u2_col_out_136;
wire  [5:0]  u2_col_out_137;
wire  [5:0]  u2_col_out_138;
wire  [5:0]  u2_col_out_139;
wire  [5:0]  u2_col_out_140;
wire  [5:0]  u2_col_out_141;
wire  [5:0]  u2_col_out_142;
wire  [5:0]  u2_col_out_143;
wire  [5:0]  u2_col_out_144;
wire  [5:0]  u2_col_out_145;
wire  [5:0]  u2_col_out_146;
wire  [5:0]  u2_col_out_147;
wire  [5:0]  u2_col_out_148;
wire  [5:0]  u2_col_out_149;
wire  [5:0]  u2_col_out_150;
wire  [5:0]  u2_col_out_151;
wire  [5:0]  u2_col_out_152;
wire  [5:0]  u2_col_out_153;
wire  [5:0]  u2_col_out_154;
wire  [5:0]  u2_col_out_155;
wire  [5:0]  u2_col_out_156;
wire  [5:0]  u2_col_out_157;
wire  [5:0]  u2_col_out_158;
wire  [5:0]  u2_col_out_159;
wire  [5:0]  u2_col_out_160;
wire  [5:0]  u2_col_out_161;
wire  [5:0]  u2_col_out_162;
wire  [5:0]  u2_col_out_163;
wire  [5:0]  u2_col_out_164;
wire  [5:0]  u2_col_out_165;
wire  [5:0]  u2_col_out_166;
wire  [5:0]  u2_col_out_167;
wire  [5:0]  u2_col_out_168;
wire  [5:0]  u2_col_out_169;
wire  [5:0]  u2_col_out_170;
wire  [5:0]  u2_col_out_171;
wire  [5:0]  u2_col_out_172;
wire  [5:0]  u2_col_out_173;
wire  [5:0]  u2_col_out_174;
wire  [5:0]  u2_col_out_175;
wire  [5:0]  u2_col_out_176;
wire  [5:0]  u2_col_out_177;
wire  [5:0]  u2_col_out_178;
wire  [5:0]  u2_col_out_179;
wire  [5:0]  u2_col_out_180;
wire  [5:0]  u2_col_out_181;
wire  [5:0]  u2_col_out_182;
wire  [5:0]  u2_col_out_183;
wire  [5:0]  u2_col_out_184;
wire  [5:0]  u2_col_out_185;
wire  [5:0]  u2_col_out_186;
wire  [5:0]  u2_col_out_187;
wire  [5:0]  u2_col_out_188;
wire  [5:0]  u2_col_out_189;
wire  [5:0]  u2_col_out_190;
wire  [5:0]  u2_col_out_191;
wire  [5:0]  u2_col_out_192;
wire  [5:0]  u2_col_out_193;
wire  [5:0]  u2_col_out_194;
wire  [5:0]  u2_col_out_195;
wire  [5:0]  u2_col_out_196;
wire  [5:0]  u2_col_out_197;
wire  [5:0]  u2_col_out_198;
wire  [5:0]  u2_col_out_199;
wire  [5:0]  u2_col_out_200;
wire  [5:0]  u2_col_out_201;
wire  [5:0]  u2_col_out_202;
wire  [5:0]  u2_col_out_203;
wire  [5:0]  u2_col_out_204;
wire  [5:0]  u2_col_out_205;
wire  [5:0]  u2_col_out_206;
wire  [5:0]  u2_col_out_207;
wire  [5:0]  u2_col_out_208;
wire  [5:0]  u2_col_out_209;
wire  [5:0]  u2_col_out_210;
wire  [5:0]  u2_col_out_211;
wire  [5:0]  u2_col_out_212;
wire  [5:0]  u2_col_out_213;
wire  [5:0]  u2_col_out_214;
wire  [5:0]  u2_col_out_215;
wire  [5:0]  u2_col_out_216;
wire  [5:0]  u2_col_out_217;
wire  [5:0]  u2_col_out_218;
wire  [5:0]  u2_col_out_219;
wire  [5:0]  u2_col_out_220;
wire  [5:0]  u2_col_out_221;
wire  [5:0]  u2_col_out_222;
wire  [5:0]  u2_col_out_223;
wire  [5:0]  u2_col_out_224;
wire  [5:0]  u2_col_out_225;
wire  [5:0]  u2_col_out_226;
wire  [5:0]  u2_col_out_227;
wire  [5:0]  u2_col_out_228;
wire  [5:0]  u2_col_out_229;
wire  [5:0]  u2_col_out_230;
wire  [5:0]  u2_col_out_231;
wire  [5:0]  u2_col_out_232;
wire  [5:0]  u2_col_out_233;
wire  [5:0]  u2_col_out_234;
wire  [5:0]  u2_col_out_235;
wire  [5:0]  u2_col_out_236;
wire  [5:0]  u2_col_out_237;
wire  [5:0]  u2_col_out_238;
wire  [5:0]  u2_col_out_239;
wire  [5:0]  u2_col_out_240;
wire  [5:0]  u2_col_out_241;
wire  [5:0]  u2_col_out_242;
wire  [5:0]  u2_col_out_243;
wire  [5:0]  u2_col_out_244;
wire  [5:0]  u2_col_out_245;
wire  [5:0]  u2_col_out_246;
wire  [5:0]  u2_col_out_247;
wire  [5:0]  u2_col_out_248;
wire  [5:0]  u2_col_out_249;
wire  [5:0]  u2_col_out_250;
wire  [5:0]  u2_col_out_251;
wire  [5:0]  u2_col_out_252;
wire  [5:0]  u2_col_out_253;
wire  [5:0]  u2_col_out_254;
wire  [5:0]  u2_col_out_255;
wire  [5:0]  u2_col_out_256;
wire  [5:0]  u2_col_out_257;
wire  [5:0]  u2_col_out_258;
wire  [5:0]  u2_col_out_259;
wire  [5:0]  u2_col_out_260;
wire  [5:0]  u2_col_out_261;
wire  [5:0]  u2_col_out_262;
wire  [5:0]  u2_col_out_263;
wire  [5:0]  u2_col_out_264;
wire  [5:0]  u2_col_out_265;
wire  [5:0]  u2_col_out_266;
wire  [5:0]  u2_col_out_267;
wire  [5:0]  u2_col_out_268;
wire  [5:0]  u2_col_out_269;
wire  [5:0]  u2_col_out_270;
wire  [5:0]  u2_col_out_271;
wire  [5:0]  u2_col_out_272;
wire  [5:0]  u2_col_out_273;
wire  [5:0]  u2_col_out_274;
wire  [5:0]  u2_col_out_275;
wire  [5:0]  u2_col_out_276;
wire  [5:0]  u2_col_out_277;
wire  [5:0]  u2_col_out_278;
wire  [5:0]  u2_col_out_279;
wire  [5:0]  u2_col_out_280;
wire  [5:0]  u2_col_out_281;
wire  [5:0]  u2_col_out_282;
wire  [5:0]  u2_col_out_283;
wire  [5:0]  u2_col_out_284;
wire  [5:0]  u2_col_out_285;
wire  [5:0]  u2_col_out_286;
wire  [5:0]  u2_col_out_287;
wire  [5:0]  u2_col_out_288;
wire  [5:0]  u2_col_out_289;
wire  [5:0]  u2_col_out_290;
wire  [5:0]  u2_col_out_291;
wire  [5:0]  u2_col_out_292;
wire  [5:0]  u2_col_out_293;
wire  [5:0]  u2_col_out_294;
wire  [5:0]  u2_col_out_295;
wire  [5:0]  u2_col_out_296;
wire  [5:0]  u2_col_out_297;
wire  [5:0]  u2_col_out_298;
wire  [5:0]  u2_col_out_299;
wire  [5:0]  u2_col_out_300;
wire  [5:0]  u2_col_out_301;
wire  [5:0]  u2_col_out_302;
wire  [5:0]  u2_col_out_303;
wire  [5:0]  u2_col_out_304;
wire  [5:0]  u2_col_out_305;
wire  [5:0]  u2_col_out_306;
wire  [5:0]  u2_col_out_307;
wire  [5:0]  u2_col_out_308;
wire  [5:0]  u2_col_out_309;
wire  [5:0]  u2_col_out_310;
wire  [5:0]  u2_col_out_311;
wire  [5:0]  u2_col_out_312;
wire  [5:0]  u2_col_out_313;
wire  [5:0]  u2_col_out_314;
wire  [5:0]  u2_col_out_315;
wire  [5:0]  u2_col_out_316;
wire  [5:0]  u2_col_out_317;
wire  [5:0]  u2_col_out_318;
wire  [5:0]  u2_col_out_319;
wire  [5:0]  u2_col_out_320;
wire  [5:0]  u2_col_out_321;
wire  [5:0]  u2_col_out_322;
wire  [5:0]  u2_col_out_323;
wire  [5:0]  u2_col_out_324;
wire  [5:0]  u2_col_out_325;
wire  [5:0]  u2_col_out_326;
wire  [5:0]  u2_col_out_327;
wire  [5:0]  u2_col_out_328;
wire  [5:0]  u2_col_out_329;
wire  [5:0]  u2_col_out_330;
wire  [5:0]  u2_col_out_331;
wire  [5:0]  u2_col_out_332;
wire  [5:0]  u2_col_out_333;
wire  [5:0]  u2_col_out_334;
wire  [5:0]  u2_col_out_335;
wire  [5:0]  u2_col_out_336;
wire  [5:0]  u2_col_out_337;
wire  [5:0]  u2_col_out_338;
wire  [5:0]  u2_col_out_339;
wire  [5:0]  u2_col_out_340;
wire  [5:0]  u2_col_out_341;
wire  [5:0]  u2_col_out_342;
wire  [5:0]  u2_col_out_343;
wire  [5:0]  u2_col_out_344;
wire  [5:0]  u2_col_out_345;
wire  [5:0]  u2_col_out_346;
wire  [5:0]  u2_col_out_347;
wire  [5:0]  u2_col_out_348;
wire  [5:0]  u2_col_out_349;
wire  [5:0]  u2_col_out_350;
wire  [5:0]  u2_col_out_351;
wire  [5:0]  u2_col_out_352;
wire  [5:0]  u2_col_out_353;
wire  [5:0]  u2_col_out_354;
wire  [5:0]  u2_col_out_355;
wire  [5:0]  u2_col_out_356;
wire  [5:0]  u2_col_out_357;
wire  [5:0]  u2_col_out_358;
wire  [5:0]  u2_col_out_359;
wire  [5:0]  u2_col_out_360;
wire  [5:0]  u2_col_out_361;
wire  [5:0]  u2_col_out_362;
wire  [5:0]  u2_col_out_363;
wire  [5:0]  u2_col_out_364;
wire  [5:0]  u2_col_out_365;
wire  [5:0]  u2_col_out_366;
wire  [5:0]  u2_col_out_367;
wire  [5:0]  u2_col_out_368;
wire  [5:0]  u2_col_out_369;
wire  [5:0]  u2_col_out_370;
wire  [5:0]  u2_col_out_371;
wire  [5:0]  u2_col_out_372;
wire  [5:0]  u2_col_out_373;
wire  [5:0]  u2_col_out_374;
wire  [5:0]  u2_col_out_375;
wire  [5:0]  u2_col_out_376;
wire  [5:0]  u2_col_out_377;
wire  [5:0]  u2_col_out_378;
wire  [5:0]  u2_col_out_379;
wire  [5:0]  u2_col_out_380;
wire  [5:0]  u2_col_out_381;
wire  [5:0]  u2_col_out_382;
wire  [5:0]  u2_col_out_383;
wire  [5:0]  u2_col_out_384;
wire  [5:0]  u2_col_out_385;
wire  [5:0]  u2_col_out_386;
wire  [5:0]  u2_col_out_387;
wire  [5:0]  u2_col_out_388;
wire  [5:0]  u2_col_out_389;
wire  [5:0]  u2_col_out_390;
wire  [5:0]  u2_col_out_391;
wire  [5:0]  u2_col_out_392;
wire  [5:0]  u2_col_out_393;
wire  [5:0]  u2_col_out_394;
wire  [5:0]  u2_col_out_395;
wire  [5:0]  u2_col_out_396;
wire  [5:0]  u2_col_out_397;
wire  [5:0]  u2_col_out_398;
wire  [5:0]  u2_col_out_399;
wire  [5:0]  u2_col_out_400;
wire  [5:0]  u2_col_out_401;
wire  [5:0]  u2_col_out_402;
wire  [5:0]  u2_col_out_403;
wire  [5:0]  u2_col_out_404;
wire  [5:0]  u2_col_out_405;
wire  [5:0]  u2_col_out_406;
wire  [5:0]  u2_col_out_407;
wire  [5:0]  u2_col_out_408;
wire  [5:0]  u2_col_out_409;
wire  [5:0]  u2_col_out_410;
wire  [5:0]  u2_col_out_411;
wire  [5:0]  u2_col_out_412;
wire  [5:0]  u2_col_out_413;
wire  [5:0]  u2_col_out_414;
wire  [5:0]  u2_col_out_415;
wire  [5:0]  u2_col_out_416;
wire  [5:0]  u2_col_out_417;
wire  [5:0]  u2_col_out_418;
wire  [5:0]  u2_col_out_419;
wire  [5:0]  u2_col_out_420;
wire  [5:0]  u2_col_out_421;
wire  [5:0]  u2_col_out_422;
wire  [5:0]  u2_col_out_423;
wire  [5:0]  u2_col_out_424;
wire  [5:0]  u2_col_out_425;
wire  [5:0]  u2_col_out_426;
wire  [5:0]  u2_col_out_427;
wire  [5:0]  u2_col_out_428;
wire  [5:0]  u2_col_out_429;
wire  [5:0]  u2_col_out_430;
wire  [5:0]  u2_col_out_431;
wire  [5:0]  u2_col_out_432;
wire  [5:0]  u2_col_out_433;
wire  [5:0]  u2_col_out_434;
wire  [5:0]  u2_col_out_435;
wire  [5:0]  u2_col_out_436;
wire  [5:0]  u2_col_out_437;
wire  [5:0]  u2_col_out_438;
wire  [5:0]  u2_col_out_439;
wire  [5:0]  u2_col_out_440;
wire  [5:0]  u2_col_out_441;
wire  [5:0]  u2_col_out_442;
wire  [5:0]  u2_col_out_443;
wire  [5:0]  u2_col_out_444;
wire  [5:0]  u2_col_out_445;
wire  [5:0]  u2_col_out_446;
wire  [5:0]  u2_col_out_447;
wire  [5:0]  u2_col_out_448;
wire  [5:0]  u2_col_out_449;
wire  [5:0]  u2_col_out_450;
wire  [5:0]  u2_col_out_451;
wire  [5:0]  u2_col_out_452;
wire  [5:0]  u2_col_out_453;
wire  [5:0]  u2_col_out_454;
wire  [5:0]  u2_col_out_455;
wire  [5:0]  u2_col_out_456;
wire  [5:0]  u2_col_out_457;
wire  [5:0]  u2_col_out_458;
wire  [5:0]  u2_col_out_459;
wire  [5:0]  u2_col_out_460;
wire  [5:0]  u2_col_out_461;
wire  [5:0]  u2_col_out_462;
wire  [5:0]  u2_col_out_463;
wire  [5:0]  u2_col_out_464;
wire  [5:0]  u2_col_out_465;
wire  [5:0]  u2_col_out_466;
wire  [5:0]  u2_col_out_467;
wire  [5:0]  u2_col_out_468;
wire  [5:0]  u2_col_out_469;
wire  [5:0]  u2_col_out_470;
wire  [5:0]  u2_col_out_471;
wire  [5:0]  u2_col_out_472;
wire  [5:0]  u2_col_out_473;
wire  [5:0]  u2_col_out_474;
wire  [5:0]  u2_col_out_475;
wire  [5:0]  u2_col_out_476;
wire  [5:0]  u2_col_out_477;
wire  [5:0]  u2_col_out_478;
wire  [5:0]  u2_col_out_479;
wire  [5:0]  u2_col_out_480;
wire  [5:0]  u2_col_out_481;
wire  [5:0]  u2_col_out_482;
wire  [5:0]  u2_col_out_483;
wire  [5:0]  u2_col_out_484;
wire  [5:0]  u2_col_out_485;
wire  [5:0]  u2_col_out_486;
wire  [5:0]  u2_col_out_487;
wire  [5:0]  u2_col_out_488;
wire  [5:0]  u2_col_out_489;
wire  [5:0]  u2_col_out_490;
wire  [5:0]  u2_col_out_491;
wire  [5:0]  u2_col_out_492;
wire  [5:0]  u2_col_out_493;
wire  [5:0]  u2_col_out_494;
wire  [5:0]  u2_col_out_495;
wire  [5:0]  u2_col_out_496;
wire  [5:0]  u2_col_out_497;
wire  [5:0]  u2_col_out_498;
wire  [5:0]  u2_col_out_499;
wire  [5:0]  u2_col_out_500;
wire  [5:0]  u2_col_out_501;
wire  [5:0]  u2_col_out_502;
wire  [5:0]  u2_col_out_503;
wire  [5:0]  u2_col_out_504;
wire  [5:0]  u2_col_out_505;
wire  [5:0]  u2_col_out_506;
wire  [5:0]  u2_col_out_507;
wire  [5:0]  u2_col_out_508;
wire  [5:0]  u2_col_out_509;
wire  [5:0]  u2_col_out_510;
wire  [5:0]  u2_col_out_511;
wire  [5:0]  u2_col_out_512;
wire  [5:0]  u2_col_out_513;
wire  [5:0]  u2_col_out_514;
wire  [5:0]  u2_col_out_515;
wire  [5:0]  u2_col_out_516;
wire  [5:0]  u2_col_out_517;
wire  [5:0]  u2_col_out_518;
wire  [5:0]  u2_col_out_519;
wire  [5:0]  u2_col_out_520;
wire  [5:0]  u2_col_out_521;
wire  [5:0]  u2_col_out_522;
wire  [5:0]  u2_col_out_523;
wire  [5:0]  u2_col_out_524;
wire  [5:0]  u2_col_out_525;
wire  [5:0]  u2_col_out_526;
wire  [5:0]  u2_col_out_527;
wire  [5:0]  u2_col_out_528;
wire  [5:0]  u2_col_out_529;
wire  [5:0]  u2_col_out_530;
wire  [5:0]  u2_col_out_531;
wire  [5:0]  u2_col_out_532;
wire  [5:0]  u2_col_out_533;
wire  [5:0]  u2_col_out_534;
wire  [5:0]  u2_col_out_535;
wire  [5:0]  u2_col_out_536;
wire  [5:0]  u2_col_out_537;
wire  [5:0]  u2_col_out_538;
wire  [5:0]  u2_col_out_539;
wire  [5:0]  u2_col_out_540;
wire  [5:0]  u2_col_out_541;
wire  [5:0]  u2_col_out_542;
wire  [5:0]  u2_col_out_543;
wire  [5:0]  u2_col_out_544;
wire  [5:0]  u2_col_out_545;
wire  [5:0]  u2_col_out_546;
wire  [5:0]  u2_col_out_547;
wire  [5:0]  u2_col_out_548;
wire  [5:0]  u2_col_out_549;
wire  [5:0]  u2_col_out_550;
wire  [5:0]  u2_col_out_551;
wire  [5:0]  u2_col_out_552;
wire  [5:0]  u2_col_out_553;
wire  [5:0]  u2_col_out_554;
wire  [5:0]  u2_col_out_555;
wire  [5:0]  u2_col_out_556;
wire  [5:0]  u2_col_out_557;
wire  [5:0]  u2_col_out_558;
wire  [5:0]  u2_col_out_559;
wire  [5:0]  u2_col_out_560;
wire  [5:0]  u2_col_out_561;
wire  [5:0]  u2_col_out_562;
wire  [5:0]  u2_col_out_563;
wire  [5:0]  u2_col_out_564;
wire  [5:0]  u2_col_out_565;
wire  [5:0]  u2_col_out_566;
wire  [5:0]  u2_col_out_567;
wire  [5:0]  u2_col_out_568;
wire  [5:0]  u2_col_out_569;
wire  [5:0]  u2_col_out_570;
wire  [5:0]  u2_col_out_571;
wire  [5:0]  u2_col_out_572;
wire  [5:0]  u2_col_out_573;
wire  [5:0]  u2_col_out_574;
wire  [5:0]  u2_col_out_575;
wire  [5:0]  u2_col_out_576;
wire  [5:0]  u2_col_out_577;
wire  [5:0]  u2_col_out_578;
wire  [5:0]  u2_col_out_579;
wire  [5:0]  u2_col_out_580;
wire  [5:0]  u2_col_out_581;
wire  [5:0]  u2_col_out_582;
wire  [5:0]  u2_col_out_583;
wire  [5:0]  u2_col_out_584;
wire  [5:0]  u2_col_out_585;
wire  [5:0]  u2_col_out_586;
wire  [5:0]  u2_col_out_587;
wire  [5:0]  u2_col_out_588;
wire  [5:0]  u2_col_out_589;
wire  [5:0]  u2_col_out_590;
wire  [5:0]  u2_col_out_591;
wire  [5:0]  u2_col_out_592;
wire  [5:0]  u2_col_out_593;
wire  [5:0]  u2_col_out_594;
wire  [5:0]  u2_col_out_595;
wire  [5:0]  u2_col_out_596;
wire  [5:0]  u2_col_out_597;
wire  [5:0]  u2_col_out_598;
wire  [5:0]  u2_col_out_599;
wire  [5:0]  u2_col_out_600;
wire  [5:0]  u2_col_out_601;
wire  [5:0]  u2_col_out_602;
wire  [5:0]  u2_col_out_603;
wire  [5:0]  u2_col_out_604;
wire  [5:0]  u2_col_out_605;
wire  [5:0]  u2_col_out_606;
wire  [5:0]  u2_col_out_607;
wire  [5:0]  u2_col_out_608;
wire  [5:0]  u2_col_out_609;
wire  [5:0]  u2_col_out_610;
wire  [5:0]  u2_col_out_611;
wire  [5:0]  u2_col_out_612;
wire  [5:0]  u2_col_out_613;
wire  [5:0]  u2_col_out_614;
wire  [5:0]  u2_col_out_615;
wire  [5:0]  u2_col_out_616;
wire  [5:0]  u2_col_out_617;
wire  [5:0]  u2_col_out_618;
wire  [5:0]  u2_col_out_619;
wire  [5:0]  u2_col_out_620;
wire  [5:0]  u2_col_out_621;
wire  [5:0]  u2_col_out_622;
wire  [5:0]  u2_col_out_623;
wire  [5:0]  u2_col_out_624;
wire  [5:0]  u2_col_out_625;
wire  [5:0]  u2_col_out_626;
wire  [5:0]  u2_col_out_627;
wire  [5:0]  u2_col_out_628;
wire  [5:0]  u2_col_out_629;
wire  [5:0]  u2_col_out_630;
wire  [5:0]  u2_col_out_631;
wire  [5:0]  u2_col_out_632;
wire  [5:0]  u2_col_out_633;
wire  [5:0]  u2_col_out_634;
wire  [5:0]  u2_col_out_635;
wire  [5:0]  u2_col_out_636;
wire  [5:0]  u2_col_out_637;
wire  [5:0]  u2_col_out_638;
wire  [5:0]  u2_col_out_639;
wire  [5:0]  u2_col_out_640;
wire  [5:0]  u2_col_out_641;
wire  [5:0]  u2_col_out_642;
wire  [5:0]  u2_col_out_643;
wire  [5:0]  u2_col_out_644;
wire  [5:0]  u2_col_out_645;
wire  [5:0]  u2_col_out_646;
wire  [5:0]  u2_col_out_647;
wire  [5:0]  u2_col_out_648;
wire  [5:0]  u2_col_out_649;
wire  [5:0]  u2_col_out_650;
wire  [5:0]  u2_col_out_651;
wire  [5:0]  u2_col_out_652;
wire  [5:0]  u2_col_out_653;
wire  [5:0]  u2_col_out_654;
wire  [5:0]  u2_col_out_655;
wire  [5:0]  u2_col_out_656;
wire  [5:0]  u2_col_out_657;
wire  [5:0]  u2_col_out_658;
wire  [5:0]  u2_col_out_659;
wire  [5:0]  u2_col_out_660;
wire  [5:0]  u2_col_out_661;
wire  [5:0]  u2_col_out_662;
wire  [5:0]  u2_col_out_663;
wire  [5:0]  u2_col_out_664;
wire  [5:0]  u2_col_out_665;
wire  [5:0]  u2_col_out_666;
wire  [5:0]  u2_col_out_667;
wire  [5:0]  u2_col_out_668;
wire  [5:0]  u2_col_out_669;
wire  [5:0]  u2_col_out_670;
wire  [5:0]  u2_col_out_671;
wire  [5:0]  u2_col_out_672;
wire  [5:0]  u2_col_out_673;
wire  [5:0]  u2_col_out_674;
wire  [5:0]  u2_col_out_675;
wire  [5:0]  u2_col_out_676;
wire  [5:0]  u2_col_out_677;
wire  [5:0]  u2_col_out_678;
wire  [5:0]  u2_col_out_679;
wire  [5:0]  u2_col_out_680;
wire  [5:0]  u2_col_out_681;
wire  [5:0]  u2_col_out_682;
wire  [5:0]  u2_col_out_683;
wire  [5:0]  u2_col_out_684;
wire  [5:0]  u2_col_out_685;
wire  [5:0]  u2_col_out_686;
wire  [5:0]  u2_col_out_687;
wire  [5:0]  u2_col_out_688;
wire  [5:0]  u2_col_out_689;
wire  [5:0]  u2_col_out_690;
wire  [5:0]  u2_col_out_691;
wire  [5:0]  u2_col_out_692;
wire  [5:0]  u2_col_out_693;
wire  [5:0]  u2_col_out_694;
wire  [5:0]  u2_col_out_695;
wire  [5:0]  u2_col_out_696;
wire  [5:0]  u2_col_out_697;
wire  [5:0]  u2_col_out_698;
wire  [5:0]  u2_col_out_699;
wire  [5:0]  u2_col_out_700;
wire  [5:0]  u2_col_out_701;
wire  [5:0]  u2_col_out_702;
wire  [5:0]  u2_col_out_703;
wire  [5:0]  u2_col_out_704;
wire  [5:0]  u2_col_out_705;
wire  [5:0]  u2_col_out_706;
wire  [5:0]  u2_col_out_707;
wire  [5:0]  u2_col_out_708;
wire  [5:0]  u2_col_out_709;
wire  [5:0]  u2_col_out_710;
wire  [5:0]  u2_col_out_711;
wire  [5:0]  u2_col_out_712;
wire  [5:0]  u2_col_out_713;
wire  [5:0]  u2_col_out_714;
wire  [5:0]  u2_col_out_715;
wire  [5:0]  u2_col_out_716;
wire  [5:0]  u2_col_out_717;
wire  [5:0]  u2_col_out_718;
wire  [5:0]  u2_col_out_719;
wire  [5:0]  u2_col_out_720;
wire  [5:0]  u2_col_out_721;
wire  [5:0]  u2_col_out_722;
wire  [5:0]  u2_col_out_723;
wire  [5:0]  u2_col_out_724;
wire  [5:0]  u2_col_out_725;
wire  [5:0]  u2_col_out_726;
wire  [5:0]  u2_col_out_727;
wire  [5:0]  u2_col_out_728;
wire  [5:0]  u2_col_out_729;
wire  [5:0]  u2_col_out_730;
wire  [5:0]  u2_col_out_731;
wire  [5:0]  u2_col_out_732;
wire  [5:0]  u2_col_out_733;
wire  [5:0]  u2_col_out_734;
wire  [5:0]  u2_col_out_735;
wire  [5:0]  u2_col_out_736;
wire  [5:0]  u2_col_out_737;
wire  [5:0]  u2_col_out_738;
wire  [5:0]  u2_col_out_739;
wire  [5:0]  u2_col_out_740;
wire  [5:0]  u2_col_out_741;
wire  [5:0]  u2_col_out_742;
wire  [5:0]  u2_col_out_743;
wire  [5:0]  u2_col_out_744;
wire  [5:0]  u2_col_out_745;
wire  [5:0]  u2_col_out_746;
wire  [5:0]  u2_col_out_747;
wire  [5:0]  u2_col_out_748;
wire  [5:0]  u2_col_out_749;
wire  [5:0]  u2_col_out_750;
wire  [5:0]  u2_col_out_751;
wire  [5:0]  u2_col_out_752;
wire  [5:0]  u2_col_out_753;
wire  [5:0]  u2_col_out_754;
wire  [5:0]  u2_col_out_755;
wire  [5:0]  u2_col_out_756;
wire  [5:0]  u2_col_out_757;
wire  [5:0]  u2_col_out_758;
wire  [5:0]  u2_col_out_759;
wire  [5:0]  u2_col_out_760;
wire  [5:0]  u2_col_out_761;
wire  [5:0]  u2_col_out_762;
wire  [5:0]  u2_col_out_763;
wire  [5:0]  u2_col_out_764;
wire  [5:0]  u2_col_out_765;
wire  [5:0]  u2_col_out_766;
wire  [5:0]  u2_col_out_767;
wire  [5:0]  u2_col_out_768;
wire  [5:0]  u2_col_out_769;
wire  [5:0]  u2_col_out_770;
wire  [5:0]  u2_col_out_771;
wire  [5:0]  u2_col_out_772;
wire  [5:0]  u2_col_out_773;
wire  [5:0]  u2_col_out_774;
wire  [5:0]  u2_col_out_775;
wire  [5:0]  u2_col_out_776;
wire  [5:0]  u2_col_out_777;
wire  [5:0]  u2_col_out_778;
wire  [5:0]  u2_col_out_779;
wire  [5:0]  u2_col_out_780;
wire  [5:0]  u2_col_out_781;
wire  [5:0]  u2_col_out_782;
wire  [5:0]  u2_col_out_783;
wire  [5:0]  u2_col_out_784;
wire  [5:0]  u2_col_out_785;
wire  [5:0]  u2_col_out_786;
wire  [5:0]  u2_col_out_787;
wire  [5:0]  u2_col_out_788;
wire  [5:0]  u2_col_out_789;
wire  [5:0]  u2_col_out_790;
wire  [5:0]  u2_col_out_791;
wire  [5:0]  u2_col_out_792;
wire  [5:0]  u2_col_out_793;
wire  [5:0]  u2_col_out_794;
wire  [5:0]  u2_col_out_795;
wire  [5:0]  u2_col_out_796;
wire  [5:0]  u2_col_out_797;
wire  [5:0]  u2_col_out_798;
wire  [5:0]  u2_col_out_799;
wire  [5:0]  u2_col_out_800;
wire  [5:0]  u2_col_out_801;
wire  [5:0]  u2_col_out_802;
wire  [5:0]  u2_col_out_803;
wire  [5:0]  u2_col_out_804;
wire  [5:0]  u2_col_out_805;
wire  [5:0]  u2_col_out_806;
wire  [5:0]  u2_col_out_807;
wire  [5:0]  u2_col_out_808;
wire  [5:0]  u2_col_out_809;
wire  [5:0]  u2_col_out_810;
wire  [5:0]  u2_col_out_811;
wire  [5:0]  u2_col_out_812;
wire  [5:0]  u2_col_out_813;
wire  [5:0]  u2_col_out_814;
wire  [5:0]  u2_col_out_815;
wire  [5:0]  u2_col_out_816;
wire  [5:0]  u2_col_out_817;
wire  [5:0]  u2_col_out_818;
wire  [5:0]  u2_col_out_819;
wire  [5:0]  u2_col_out_820;
wire  [5:0]  u2_col_out_821;
wire  [5:0]  u2_col_out_822;
wire  [5:0]  u2_col_out_823;
wire  [5:0]  u2_col_out_824;
wire  [5:0]  u2_col_out_825;
wire  [5:0]  u2_col_out_826;
wire  [5:0]  u2_col_out_827;
wire  [5:0]  u2_col_out_828;
wire  [5:0]  u2_col_out_829;
wire  [5:0]  u2_col_out_830;
wire  [5:0]  u2_col_out_831;
wire  [5:0]  u2_col_out_832;
wire  [5:0]  u2_col_out_833;
wire  [5:0]  u2_col_out_834;
wire  [5:0]  u2_col_out_835;
wire  [5:0]  u2_col_out_836;
wire  [5:0]  u2_col_out_837;
wire  [5:0]  u2_col_out_838;
wire  [5:0]  u2_col_out_839;
wire  [5:0]  u2_col_out_840;
wire  [5:0]  u2_col_out_841;
wire  [5:0]  u2_col_out_842;
wire  [5:0]  u2_col_out_843;
wire  [5:0]  u2_col_out_844;
wire  [5:0]  u2_col_out_845;
wire  [5:0]  u2_col_out_846;
wire  [5:0]  u2_col_out_847;
wire  [5:0]  u2_col_out_848;
wire  [5:0]  u2_col_out_849;
wire  [5:0]  u2_col_out_850;
wire  [5:0]  u2_col_out_851;
wire  [5:0]  u2_col_out_852;
wire  [5:0]  u2_col_out_853;
wire  [5:0]  u2_col_out_854;
wire  [5:0]  u2_col_out_855;
wire  [5:0]  u2_col_out_856;
wire  [5:0]  u2_col_out_857;
wire  [5:0]  u2_col_out_858;
wire  [5:0]  u2_col_out_859;
wire  [5:0]  u2_col_out_860;
wire  [5:0]  u2_col_out_861;
wire  [5:0]  u2_col_out_862;
wire  [5:0]  u2_col_out_863;
wire  [5:0]  u2_col_out_864;
wire  [5:0]  u2_col_out_865;
wire  [5:0]  u2_col_out_866;
wire  [5:0]  u2_col_out_867;
wire  [5:0]  u2_col_out_868;
wire  [5:0]  u2_col_out_869;
wire  [5:0]  u2_col_out_870;
wire  [5:0]  u2_col_out_871;
wire  [5:0]  u2_col_out_872;
wire  [5:0]  u2_col_out_873;
wire  [5:0]  u2_col_out_874;
wire  [5:0]  u2_col_out_875;
wire  [5:0]  u2_col_out_876;
wire  [5:0]  u2_col_out_877;
wire  [5:0]  u2_col_out_878;
wire  [5:0]  u2_col_out_879;
wire  [5:0]  u2_col_out_880;
wire  [5:0]  u2_col_out_881;
wire  [5:0]  u2_col_out_882;
wire  [5:0]  u2_col_out_883;
wire  [5:0]  u2_col_out_884;
wire  [5:0]  u2_col_out_885;
wire  [5:0]  u2_col_out_886;
wire  [5:0]  u2_col_out_887;
wire  [5:0]  u2_col_out_888;
wire  [5:0]  u2_col_out_889;
wire  [5:0]  u2_col_out_890;
wire  [5:0]  u2_col_out_891;
wire  [5:0]  u2_col_out_892;
wire  [5:0]  u2_col_out_893;
wire  [5:0]  u2_col_out_894;
wire  [5:0]  u2_col_out_895;
wire  [5:0]  u2_col_out_896;
wire  [5:0]  u2_col_out_897;
wire  [5:0]  u2_col_out_898;
wire  [5:0]  u2_col_out_899;
wire  [5:0]  u2_col_out_900;
wire  [5:0]  u2_col_out_901;
wire  [5:0]  u2_col_out_902;
wire  [5:0]  u2_col_out_903;
wire  [5:0]  u2_col_out_904;
wire  [5:0]  u2_col_out_905;
wire  [5:0]  u2_col_out_906;
wire  [5:0]  u2_col_out_907;
wire  [5:0]  u2_col_out_908;
wire  [5:0]  u2_col_out_909;
wire  [5:0]  u2_col_out_910;
wire  [5:0]  u2_col_out_911;
wire  [5:0]  u2_col_out_912;
wire  [5:0]  u2_col_out_913;
wire  [5:0]  u2_col_out_914;
wire  [5:0]  u2_col_out_915;
wire  [5:0]  u2_col_out_916;
wire  [5:0]  u2_col_out_917;
wire  [5:0]  u2_col_out_918;
wire  [5:0]  u2_col_out_919;
wire  [5:0]  u2_col_out_920;
wire  [5:0]  u2_col_out_921;
wire  [5:0]  u2_col_out_922;
wire  [5:0]  u2_col_out_923;
wire  [5:0]  u2_col_out_924;
wire  [5:0]  u2_col_out_925;
wire  [5:0]  u2_col_out_926;
wire  [5:0]  u2_col_out_927;
wire  [5:0]  u2_col_out_928;
wire  [5:0]  u2_col_out_929;
wire  [5:0]  u2_col_out_930;
wire  [5:0]  u2_col_out_931;
wire  [5:0]  u2_col_out_932;
wire  [5:0]  u2_col_out_933;
wire  [5:0]  u2_col_out_934;
wire  [5:0]  u2_col_out_935;
wire  [5:0]  u2_col_out_936;
wire  [5:0]  u2_col_out_937;
wire  [5:0]  u2_col_out_938;
wire  [5:0]  u2_col_out_939;
wire  [5:0]  u2_col_out_940;
wire  [5:0]  u2_col_out_941;
wire  [5:0]  u2_col_out_942;
wire  [5:0]  u2_col_out_943;
wire  [5:0]  u2_col_out_944;
wire  [5:0]  u2_col_out_945;
wire  [5:0]  u2_col_out_946;
wire  [5:0]  u2_col_out_947;
wire  [5:0]  u2_col_out_948;
wire  [5:0]  u2_col_out_949;
wire  [5:0]  u2_col_out_950;
wire  [5:0]  u2_col_out_951;
wire  [5:0]  u2_col_out_952;
wire  [5:0]  u2_col_out_953;
wire  [5:0]  u2_col_out_954;
wire  [5:0]  u2_col_out_955;
wire  [5:0]  u2_col_out_956;
wire  [5:0]  u2_col_out_957;
wire  [5:0]  u2_col_out_958;
wire  [5:0]  u2_col_out_959;
wire  [5:0]  u2_col_out_960;
wire  [5:0]  u2_col_out_961;
wire  [5:0]  u2_col_out_962;
wire  [5:0]  u2_col_out_963;
wire  [5:0]  u2_col_out_964;
wire  [5:0]  u2_col_out_965;
wire  [5:0]  u2_col_out_966;
wire  [5:0]  u2_col_out_967;
wire  [5:0]  u2_col_out_968;
wire  [5:0]  u2_col_out_969;
wire  [5:0]  u2_col_out_970;
wire  [5:0]  u2_col_out_971;
wire  [5:0]  u2_col_out_972;
wire  [5:0]  u2_col_out_973;
wire  [5:0]  u2_col_out_974;
wire  [5:0]  u2_col_out_975;
wire  [5:0]  u2_col_out_976;
wire  [5:0]  u2_col_out_977;
wire  [5:0]  u2_col_out_978;
wire  [5:0]  u2_col_out_979;
wire  [5:0]  u2_col_out_980;
wire  [5:0]  u2_col_out_981;
wire  [5:0]  u2_col_out_982;
wire  [5:0]  u2_col_out_983;
wire  [5:0]  u2_col_out_984;
wire  [5:0]  u2_col_out_985;
wire  [5:0]  u2_col_out_986;
wire  [5:0]  u2_col_out_987;
wire  [5:0]  u2_col_out_988;
wire  [5:0]  u2_col_out_989;
wire  [5:0]  u2_col_out_990;
wire  [5:0]  u2_col_out_991;
wire  [5:0]  u2_col_out_992;
wire  [5:0]  u2_col_out_993;
wire  [5:0]  u2_col_out_994;
wire  [5:0]  u2_col_out_995;
wire  [5:0]  u2_col_out_996;
wire  [5:0]  u2_col_out_997;
wire  [5:0]  u2_col_out_998;
wire  [5:0]  u2_col_out_999;
wire  [5:0]  u2_col_out_1000;
wire  [5:0]  u2_col_out_1001;
wire  [5:0]  u2_col_out_1002;
wire  [5:0]  u2_col_out_1003;
wire  [5:0]  u2_col_out_1004;
wire  [5:0]  u2_col_out_1005;
wire  [5:0]  u2_col_out_1006;
wire  [5:0]  u2_col_out_1007;
wire  [5:0]  u2_col_out_1008;
wire  [5:0]  u2_col_out_1009;
wire  [5:0]  u2_col_out_1010;
wire  [5:0]  u2_col_out_1011;
wire  [5:0]  u2_col_out_1012;
wire  [5:0]  u2_col_out_1013;
wire  [5:0]  u2_col_out_1014;
wire  [5:0]  u2_col_out_1015;
wire  [5:0]  u2_col_out_1016;
wire  [5:0]  u2_col_out_1017;
wire  [5:0]  u2_col_out_1018;
wire  [5:0]  u2_col_out_1019;
wire  [5:0]  u2_col_out_1020;
wire  [5:0]  u2_col_out_1021;
wire  [5:0]  u2_col_out_1022;
wire  [5:0]  u2_col_out_1023;
wire  [5:0]  u2_col_out_1024;
wire  [5:0]  u2_col_out_1025;
wire  [5:0]  u2_col_out_1026;
wire  [5:0]  u2_col_out_1027;
wire  [5:0]  u2_col_out_1028;
wire  [5:0]  u2_col_out_1029;
wire  [5:0]  u2_col_out_1030;
wire  [5:0]  u2_col_out_1031;
wire  [5:0]  u2_col_out_1032;
wire  [5:0]  u2_col_out_1033;

compressor_array_8_6_1033  u2_compressor_array_8_6_1033 (
    .col_in_0                ( u1_col_out_0       ),
    .col_in_1                ( u1_col_out_1       ),
    .col_in_2                ( u1_col_out_2       ),
    .col_in_3                ( u1_col_out_3       ),
    .col_in_4                ( u1_col_out_4       ),
    .col_in_5                ( u1_col_out_5       ),
    .col_in_6                ( u1_col_out_6       ),
    .col_in_7                ( u1_col_out_7       ),
    .col_in_8                ( u1_col_out_8       ),
    .col_in_9                ( u1_col_out_9       ),
    .col_in_10               ( u1_col_out_10      ),
    .col_in_11               ( u1_col_out_11      ),
    .col_in_12               ( u1_col_out_12      ),
    .col_in_13               ( u1_col_out_13      ),
    .col_in_14               ( u1_col_out_14      ),
    .col_in_15               ( u1_col_out_15      ),
    .col_in_16               ( u1_col_out_16      ),
    .col_in_17               ( u1_col_out_17      ),
    .col_in_18               ( u1_col_out_18      ),
    .col_in_19               ( u1_col_out_19      ),
    .col_in_20               ( u1_col_out_20      ),
    .col_in_21               ( u1_col_out_21      ),
    .col_in_22               ( u1_col_out_22      ),
    .col_in_23               ( u1_col_out_23      ),
    .col_in_24               ( u1_col_out_24      ),
    .col_in_25               ( u1_col_out_25      ),
    .col_in_26               ( u1_col_out_26      ),
    .col_in_27               ( u1_col_out_27      ),
    .col_in_28               ( u1_col_out_28      ),
    .col_in_29               ( u1_col_out_29      ),
    .col_in_30               ( u1_col_out_30      ),
    .col_in_31               ( u1_col_out_31      ),
    .col_in_32               ( u1_col_out_32      ),
    .col_in_33               ( u1_col_out_33      ),
    .col_in_34               ( u1_col_out_34      ),
    .col_in_35               ( u1_col_out_35      ),
    .col_in_36               ( u1_col_out_36      ),
    .col_in_37               ( u1_col_out_37      ),
    .col_in_38               ( u1_col_out_38      ),
    .col_in_39               ( u1_col_out_39      ),
    .col_in_40               ( u1_col_out_40      ),
    .col_in_41               ( u1_col_out_41      ),
    .col_in_42               ( u1_col_out_42      ),
    .col_in_43               ( u1_col_out_43      ),
    .col_in_44               ( u1_col_out_44      ),
    .col_in_45               ( u1_col_out_45      ),
    .col_in_46               ( u1_col_out_46      ),
    .col_in_47               ( u1_col_out_47      ),
    .col_in_48               ( u1_col_out_48      ),
    .col_in_49               ( u1_col_out_49      ),
    .col_in_50               ( u1_col_out_50      ),
    .col_in_51               ( u1_col_out_51      ),
    .col_in_52               ( u1_col_out_52      ),
    .col_in_53               ( u1_col_out_53      ),
    .col_in_54               ( u1_col_out_54      ),
    .col_in_55               ( u1_col_out_55      ),
    .col_in_56               ( u1_col_out_56      ),
    .col_in_57               ( u1_col_out_57      ),
    .col_in_58               ( u1_col_out_58      ),
    .col_in_59               ( u1_col_out_59      ),
    .col_in_60               ( u1_col_out_60      ),
    .col_in_61               ( u1_col_out_61      ),
    .col_in_62               ( u1_col_out_62      ),
    .col_in_63               ( u1_col_out_63      ),
    .col_in_64               ( u1_col_out_64      ),
    .col_in_65               ( u1_col_out_65      ),
    .col_in_66               ( u1_col_out_66      ),
    .col_in_67               ( u1_col_out_67      ),
    .col_in_68               ( u1_col_out_68      ),
    .col_in_69               ( u1_col_out_69      ),
    .col_in_70               ( u1_col_out_70      ),
    .col_in_71               ( u1_col_out_71      ),
    .col_in_72               ( u1_col_out_72      ),
    .col_in_73               ( u1_col_out_73      ),
    .col_in_74               ( u1_col_out_74      ),
    .col_in_75               ( u1_col_out_75      ),
    .col_in_76               ( u1_col_out_76      ),
    .col_in_77               ( u1_col_out_77      ),
    .col_in_78               ( u1_col_out_78      ),
    .col_in_79               ( u1_col_out_79      ),
    .col_in_80               ( u1_col_out_80      ),
    .col_in_81               ( u1_col_out_81      ),
    .col_in_82               ( u1_col_out_82      ),
    .col_in_83               ( u1_col_out_83      ),
    .col_in_84               ( u1_col_out_84      ),
    .col_in_85               ( u1_col_out_85      ),
    .col_in_86               ( u1_col_out_86      ),
    .col_in_87               ( u1_col_out_87      ),
    .col_in_88               ( u1_col_out_88      ),
    .col_in_89               ( u1_col_out_89      ),
    .col_in_90               ( u1_col_out_90      ),
    .col_in_91               ( u1_col_out_91      ),
    .col_in_92               ( u1_col_out_92      ),
    .col_in_93               ( u1_col_out_93      ),
    .col_in_94               ( u1_col_out_94      ),
    .col_in_95               ( u1_col_out_95      ),
    .col_in_96               ( u1_col_out_96      ),
    .col_in_97               ( u1_col_out_97      ),
    .col_in_98               ( u1_col_out_98      ),
    .col_in_99               ( u1_col_out_99      ),
    .col_in_100              ( u1_col_out_100     ),
    .col_in_101              ( u1_col_out_101     ),
    .col_in_102              ( u1_col_out_102     ),
    .col_in_103              ( u1_col_out_103     ),
    .col_in_104              ( u1_col_out_104     ),
    .col_in_105              ( u1_col_out_105     ),
    .col_in_106              ( u1_col_out_106     ),
    .col_in_107              ( u1_col_out_107     ),
    .col_in_108              ( u1_col_out_108     ),
    .col_in_109              ( u1_col_out_109     ),
    .col_in_110              ( u1_col_out_110     ),
    .col_in_111              ( u1_col_out_111     ),
    .col_in_112              ( u1_col_out_112     ),
    .col_in_113              ( u1_col_out_113     ),
    .col_in_114              ( u1_col_out_114     ),
    .col_in_115              ( u1_col_out_115     ),
    .col_in_116              ( u1_col_out_116     ),
    .col_in_117              ( u1_col_out_117     ),
    .col_in_118              ( u1_col_out_118     ),
    .col_in_119              ( u1_col_out_119     ),
    .col_in_120              ( u1_col_out_120     ),
    .col_in_121              ( u1_col_out_121     ),
    .col_in_122              ( u1_col_out_122     ),
    .col_in_123              ( u1_col_out_123     ),
    .col_in_124              ( u1_col_out_124     ),
    .col_in_125              ( u1_col_out_125     ),
    .col_in_126              ( u1_col_out_126     ),
    .col_in_127              ( u1_col_out_127     ),
    .col_in_128              ( u1_col_out_128     ),
    .col_in_129              ( u1_col_out_129     ),
    .col_in_130              ( u1_col_out_130     ),
    .col_in_131              ( u1_col_out_131     ),
    .col_in_132              ( u1_col_out_132     ),
    .col_in_133              ( u1_col_out_133     ),
    .col_in_134              ( u1_col_out_134     ),
    .col_in_135              ( u1_col_out_135     ),
    .col_in_136              ( u1_col_out_136     ),
    .col_in_137              ( u1_col_out_137     ),
    .col_in_138              ( u1_col_out_138     ),
    .col_in_139              ( u1_col_out_139     ),
    .col_in_140              ( u1_col_out_140     ),
    .col_in_141              ( u1_col_out_141     ),
    .col_in_142              ( u1_col_out_142     ),
    .col_in_143              ( u1_col_out_143     ),
    .col_in_144              ( u1_col_out_144     ),
    .col_in_145              ( u1_col_out_145     ),
    .col_in_146              ( u1_col_out_146     ),
    .col_in_147              ( u1_col_out_147     ),
    .col_in_148              ( u1_col_out_148     ),
    .col_in_149              ( u1_col_out_149     ),
    .col_in_150              ( u1_col_out_150     ),
    .col_in_151              ( u1_col_out_151     ),
    .col_in_152              ( u1_col_out_152     ),
    .col_in_153              ( u1_col_out_153     ),
    .col_in_154              ( u1_col_out_154     ),
    .col_in_155              ( u1_col_out_155     ),
    .col_in_156              ( u1_col_out_156     ),
    .col_in_157              ( u1_col_out_157     ),
    .col_in_158              ( u1_col_out_158     ),
    .col_in_159              ( u1_col_out_159     ),
    .col_in_160              ( u1_col_out_160     ),
    .col_in_161              ( u1_col_out_161     ),
    .col_in_162              ( u1_col_out_162     ),
    .col_in_163              ( u1_col_out_163     ),
    .col_in_164              ( u1_col_out_164     ),
    .col_in_165              ( u1_col_out_165     ),
    .col_in_166              ( u1_col_out_166     ),
    .col_in_167              ( u1_col_out_167     ),
    .col_in_168              ( u1_col_out_168     ),
    .col_in_169              ( u1_col_out_169     ),
    .col_in_170              ( u1_col_out_170     ),
    .col_in_171              ( u1_col_out_171     ),
    .col_in_172              ( u1_col_out_172     ),
    .col_in_173              ( u1_col_out_173     ),
    .col_in_174              ( u1_col_out_174     ),
    .col_in_175              ( u1_col_out_175     ),
    .col_in_176              ( u1_col_out_176     ),
    .col_in_177              ( u1_col_out_177     ),
    .col_in_178              ( u1_col_out_178     ),
    .col_in_179              ( u1_col_out_179     ),
    .col_in_180              ( u1_col_out_180     ),
    .col_in_181              ( u1_col_out_181     ),
    .col_in_182              ( u1_col_out_182     ),
    .col_in_183              ( u1_col_out_183     ),
    .col_in_184              ( u1_col_out_184     ),
    .col_in_185              ( u1_col_out_185     ),
    .col_in_186              ( u1_col_out_186     ),
    .col_in_187              ( u1_col_out_187     ),
    .col_in_188              ( u1_col_out_188     ),
    .col_in_189              ( u1_col_out_189     ),
    .col_in_190              ( u1_col_out_190     ),
    .col_in_191              ( u1_col_out_191     ),
    .col_in_192              ( u1_col_out_192     ),
    .col_in_193              ( u1_col_out_193     ),
    .col_in_194              ( u1_col_out_194     ),
    .col_in_195              ( u1_col_out_195     ),
    .col_in_196              ( u1_col_out_196     ),
    .col_in_197              ( u1_col_out_197     ),
    .col_in_198              ( u1_col_out_198     ),
    .col_in_199              ( u1_col_out_199     ),
    .col_in_200              ( u1_col_out_200     ),
    .col_in_201              ( u1_col_out_201     ),
    .col_in_202              ( u1_col_out_202     ),
    .col_in_203              ( u1_col_out_203     ),
    .col_in_204              ( u1_col_out_204     ),
    .col_in_205              ( u1_col_out_205     ),
    .col_in_206              ( u1_col_out_206     ),
    .col_in_207              ( u1_col_out_207     ),
    .col_in_208              ( u1_col_out_208     ),
    .col_in_209              ( u1_col_out_209     ),
    .col_in_210              ( u1_col_out_210     ),
    .col_in_211              ( u1_col_out_211     ),
    .col_in_212              ( u1_col_out_212     ),
    .col_in_213              ( u1_col_out_213     ),
    .col_in_214              ( u1_col_out_214     ),
    .col_in_215              ( u1_col_out_215     ),
    .col_in_216              ( u1_col_out_216     ),
    .col_in_217              ( u1_col_out_217     ),
    .col_in_218              ( u1_col_out_218     ),
    .col_in_219              ( u1_col_out_219     ),
    .col_in_220              ( u1_col_out_220     ),
    .col_in_221              ( u1_col_out_221     ),
    .col_in_222              ( u1_col_out_222     ),
    .col_in_223              ( u1_col_out_223     ),
    .col_in_224              ( u1_col_out_224     ),
    .col_in_225              ( u1_col_out_225     ),
    .col_in_226              ( u1_col_out_226     ),
    .col_in_227              ( u1_col_out_227     ),
    .col_in_228              ( u1_col_out_228     ),
    .col_in_229              ( u1_col_out_229     ),
    .col_in_230              ( u1_col_out_230     ),
    .col_in_231              ( u1_col_out_231     ),
    .col_in_232              ( u1_col_out_232     ),
    .col_in_233              ( u1_col_out_233     ),
    .col_in_234              ( u1_col_out_234     ),
    .col_in_235              ( u1_col_out_235     ),
    .col_in_236              ( u1_col_out_236     ),
    .col_in_237              ( u1_col_out_237     ),
    .col_in_238              ( u1_col_out_238     ),
    .col_in_239              ( u1_col_out_239     ),
    .col_in_240              ( u1_col_out_240     ),
    .col_in_241              ( u1_col_out_241     ),
    .col_in_242              ( u1_col_out_242     ),
    .col_in_243              ( u1_col_out_243     ),
    .col_in_244              ( u1_col_out_244     ),
    .col_in_245              ( u1_col_out_245     ),
    .col_in_246              ( u1_col_out_246     ),
    .col_in_247              ( u1_col_out_247     ),
    .col_in_248              ( u1_col_out_248     ),
    .col_in_249              ( u1_col_out_249     ),
    .col_in_250              ( u1_col_out_250     ),
    .col_in_251              ( u1_col_out_251     ),
    .col_in_252              ( u1_col_out_252     ),
    .col_in_253              ( u1_col_out_253     ),
    .col_in_254              ( u1_col_out_254     ),
    .col_in_255              ( u1_col_out_255     ),
    .col_in_256              ( u1_col_out_256     ),
    .col_in_257              ( u1_col_out_257     ),
    .col_in_258              ( u1_col_out_258     ),
    .col_in_259              ( u1_col_out_259     ),
    .col_in_260              ( u1_col_out_260     ),
    .col_in_261              ( u1_col_out_261     ),
    .col_in_262              ( u1_col_out_262     ),
    .col_in_263              ( u1_col_out_263     ),
    .col_in_264              ( u1_col_out_264     ),
    .col_in_265              ( u1_col_out_265     ),
    .col_in_266              ( u1_col_out_266     ),
    .col_in_267              ( u1_col_out_267     ),
    .col_in_268              ( u1_col_out_268     ),
    .col_in_269              ( u1_col_out_269     ),
    .col_in_270              ( u1_col_out_270     ),
    .col_in_271              ( u1_col_out_271     ),
    .col_in_272              ( u1_col_out_272     ),
    .col_in_273              ( u1_col_out_273     ),
    .col_in_274              ( u1_col_out_274     ),
    .col_in_275              ( u1_col_out_275     ),
    .col_in_276              ( u1_col_out_276     ),
    .col_in_277              ( u1_col_out_277     ),
    .col_in_278              ( u1_col_out_278     ),
    .col_in_279              ( u1_col_out_279     ),
    .col_in_280              ( u1_col_out_280     ),
    .col_in_281              ( u1_col_out_281     ),
    .col_in_282              ( u1_col_out_282     ),
    .col_in_283              ( u1_col_out_283     ),
    .col_in_284              ( u1_col_out_284     ),
    .col_in_285              ( u1_col_out_285     ),
    .col_in_286              ( u1_col_out_286     ),
    .col_in_287              ( u1_col_out_287     ),
    .col_in_288              ( u1_col_out_288     ),
    .col_in_289              ( u1_col_out_289     ),
    .col_in_290              ( u1_col_out_290     ),
    .col_in_291              ( u1_col_out_291     ),
    .col_in_292              ( u1_col_out_292     ),
    .col_in_293              ( u1_col_out_293     ),
    .col_in_294              ( u1_col_out_294     ),
    .col_in_295              ( u1_col_out_295     ),
    .col_in_296              ( u1_col_out_296     ),
    .col_in_297              ( u1_col_out_297     ),
    .col_in_298              ( u1_col_out_298     ),
    .col_in_299              ( u1_col_out_299     ),
    .col_in_300              ( u1_col_out_300     ),
    .col_in_301              ( u1_col_out_301     ),
    .col_in_302              ( u1_col_out_302     ),
    .col_in_303              ( u1_col_out_303     ),
    .col_in_304              ( u1_col_out_304     ),
    .col_in_305              ( u1_col_out_305     ),
    .col_in_306              ( u1_col_out_306     ),
    .col_in_307              ( u1_col_out_307     ),
    .col_in_308              ( u1_col_out_308     ),
    .col_in_309              ( u1_col_out_309     ),
    .col_in_310              ( u1_col_out_310     ),
    .col_in_311              ( u1_col_out_311     ),
    .col_in_312              ( u1_col_out_312     ),
    .col_in_313              ( u1_col_out_313     ),
    .col_in_314              ( u1_col_out_314     ),
    .col_in_315              ( u1_col_out_315     ),
    .col_in_316              ( u1_col_out_316     ),
    .col_in_317              ( u1_col_out_317     ),
    .col_in_318              ( u1_col_out_318     ),
    .col_in_319              ( u1_col_out_319     ),
    .col_in_320              ( u1_col_out_320     ),
    .col_in_321              ( u1_col_out_321     ),
    .col_in_322              ( u1_col_out_322     ),
    .col_in_323              ( u1_col_out_323     ),
    .col_in_324              ( u1_col_out_324     ),
    .col_in_325              ( u1_col_out_325     ),
    .col_in_326              ( u1_col_out_326     ),
    .col_in_327              ( u1_col_out_327     ),
    .col_in_328              ( u1_col_out_328     ),
    .col_in_329              ( u1_col_out_329     ),
    .col_in_330              ( u1_col_out_330     ),
    .col_in_331              ( u1_col_out_331     ),
    .col_in_332              ( u1_col_out_332     ),
    .col_in_333              ( u1_col_out_333     ),
    .col_in_334              ( u1_col_out_334     ),
    .col_in_335              ( u1_col_out_335     ),
    .col_in_336              ( u1_col_out_336     ),
    .col_in_337              ( u1_col_out_337     ),
    .col_in_338              ( u1_col_out_338     ),
    .col_in_339              ( u1_col_out_339     ),
    .col_in_340              ( u1_col_out_340     ),
    .col_in_341              ( u1_col_out_341     ),
    .col_in_342              ( u1_col_out_342     ),
    .col_in_343              ( u1_col_out_343     ),
    .col_in_344              ( u1_col_out_344     ),
    .col_in_345              ( u1_col_out_345     ),
    .col_in_346              ( u1_col_out_346     ),
    .col_in_347              ( u1_col_out_347     ),
    .col_in_348              ( u1_col_out_348     ),
    .col_in_349              ( u1_col_out_349     ),
    .col_in_350              ( u1_col_out_350     ),
    .col_in_351              ( u1_col_out_351     ),
    .col_in_352              ( u1_col_out_352     ),
    .col_in_353              ( u1_col_out_353     ),
    .col_in_354              ( u1_col_out_354     ),
    .col_in_355              ( u1_col_out_355     ),
    .col_in_356              ( u1_col_out_356     ),
    .col_in_357              ( u1_col_out_357     ),
    .col_in_358              ( u1_col_out_358     ),
    .col_in_359              ( u1_col_out_359     ),
    .col_in_360              ( u1_col_out_360     ),
    .col_in_361              ( u1_col_out_361     ),
    .col_in_362              ( u1_col_out_362     ),
    .col_in_363              ( u1_col_out_363     ),
    .col_in_364              ( u1_col_out_364     ),
    .col_in_365              ( u1_col_out_365     ),
    .col_in_366              ( u1_col_out_366     ),
    .col_in_367              ( u1_col_out_367     ),
    .col_in_368              ( u1_col_out_368     ),
    .col_in_369              ( u1_col_out_369     ),
    .col_in_370              ( u1_col_out_370     ),
    .col_in_371              ( u1_col_out_371     ),
    .col_in_372              ( u1_col_out_372     ),
    .col_in_373              ( u1_col_out_373     ),
    .col_in_374              ( u1_col_out_374     ),
    .col_in_375              ( u1_col_out_375     ),
    .col_in_376              ( u1_col_out_376     ),
    .col_in_377              ( u1_col_out_377     ),
    .col_in_378              ( u1_col_out_378     ),
    .col_in_379              ( u1_col_out_379     ),
    .col_in_380              ( u1_col_out_380     ),
    .col_in_381              ( u1_col_out_381     ),
    .col_in_382              ( u1_col_out_382     ),
    .col_in_383              ( u1_col_out_383     ),
    .col_in_384              ( u1_col_out_384     ),
    .col_in_385              ( u1_col_out_385     ),
    .col_in_386              ( u1_col_out_386     ),
    .col_in_387              ( u1_col_out_387     ),
    .col_in_388              ( u1_col_out_388     ),
    .col_in_389              ( u1_col_out_389     ),
    .col_in_390              ( u1_col_out_390     ),
    .col_in_391              ( u1_col_out_391     ),
    .col_in_392              ( u1_col_out_392     ),
    .col_in_393              ( u1_col_out_393     ),
    .col_in_394              ( u1_col_out_394     ),
    .col_in_395              ( u1_col_out_395     ),
    .col_in_396              ( u1_col_out_396     ),
    .col_in_397              ( u1_col_out_397     ),
    .col_in_398              ( u1_col_out_398     ),
    .col_in_399              ( u1_col_out_399     ),
    .col_in_400              ( u1_col_out_400     ),
    .col_in_401              ( u1_col_out_401     ),
    .col_in_402              ( u1_col_out_402     ),
    .col_in_403              ( u1_col_out_403     ),
    .col_in_404              ( u1_col_out_404     ),
    .col_in_405              ( u1_col_out_405     ),
    .col_in_406              ( u1_col_out_406     ),
    .col_in_407              ( u1_col_out_407     ),
    .col_in_408              ( u1_col_out_408     ),
    .col_in_409              ( u1_col_out_409     ),
    .col_in_410              ( u1_col_out_410     ),
    .col_in_411              ( u1_col_out_411     ),
    .col_in_412              ( u1_col_out_412     ),
    .col_in_413              ( u1_col_out_413     ),
    .col_in_414              ( u1_col_out_414     ),
    .col_in_415              ( u1_col_out_415     ),
    .col_in_416              ( u1_col_out_416     ),
    .col_in_417              ( u1_col_out_417     ),
    .col_in_418              ( u1_col_out_418     ),
    .col_in_419              ( u1_col_out_419     ),
    .col_in_420              ( u1_col_out_420     ),
    .col_in_421              ( u1_col_out_421     ),
    .col_in_422              ( u1_col_out_422     ),
    .col_in_423              ( u1_col_out_423     ),
    .col_in_424              ( u1_col_out_424     ),
    .col_in_425              ( u1_col_out_425     ),
    .col_in_426              ( u1_col_out_426     ),
    .col_in_427              ( u1_col_out_427     ),
    .col_in_428              ( u1_col_out_428     ),
    .col_in_429              ( u1_col_out_429     ),
    .col_in_430              ( u1_col_out_430     ),
    .col_in_431              ( u1_col_out_431     ),
    .col_in_432              ( u1_col_out_432     ),
    .col_in_433              ( u1_col_out_433     ),
    .col_in_434              ( u1_col_out_434     ),
    .col_in_435              ( u1_col_out_435     ),
    .col_in_436              ( u1_col_out_436     ),
    .col_in_437              ( u1_col_out_437     ),
    .col_in_438              ( u1_col_out_438     ),
    .col_in_439              ( u1_col_out_439     ),
    .col_in_440              ( u1_col_out_440     ),
    .col_in_441              ( u1_col_out_441     ),
    .col_in_442              ( u1_col_out_442     ),
    .col_in_443              ( u1_col_out_443     ),
    .col_in_444              ( u1_col_out_444     ),
    .col_in_445              ( u1_col_out_445     ),
    .col_in_446              ( u1_col_out_446     ),
    .col_in_447              ( u1_col_out_447     ),
    .col_in_448              ( u1_col_out_448     ),
    .col_in_449              ( u1_col_out_449     ),
    .col_in_450              ( u1_col_out_450     ),
    .col_in_451              ( u1_col_out_451     ),
    .col_in_452              ( u1_col_out_452     ),
    .col_in_453              ( u1_col_out_453     ),
    .col_in_454              ( u1_col_out_454     ),
    .col_in_455              ( u1_col_out_455     ),
    .col_in_456              ( u1_col_out_456     ),
    .col_in_457              ( u1_col_out_457     ),
    .col_in_458              ( u1_col_out_458     ),
    .col_in_459              ( u1_col_out_459     ),
    .col_in_460              ( u1_col_out_460     ),
    .col_in_461              ( u1_col_out_461     ),
    .col_in_462              ( u1_col_out_462     ),
    .col_in_463              ( u1_col_out_463     ),
    .col_in_464              ( u1_col_out_464     ),
    .col_in_465              ( u1_col_out_465     ),
    .col_in_466              ( u1_col_out_466     ),
    .col_in_467              ( u1_col_out_467     ),
    .col_in_468              ( u1_col_out_468     ),
    .col_in_469              ( u1_col_out_469     ),
    .col_in_470              ( u1_col_out_470     ),
    .col_in_471              ( u1_col_out_471     ),
    .col_in_472              ( u1_col_out_472     ),
    .col_in_473              ( u1_col_out_473     ),
    .col_in_474              ( u1_col_out_474     ),
    .col_in_475              ( u1_col_out_475     ),
    .col_in_476              ( u1_col_out_476     ),
    .col_in_477              ( u1_col_out_477     ),
    .col_in_478              ( u1_col_out_478     ),
    .col_in_479              ( u1_col_out_479     ),
    .col_in_480              ( u1_col_out_480     ),
    .col_in_481              ( u1_col_out_481     ),
    .col_in_482              ( u1_col_out_482     ),
    .col_in_483              ( u1_col_out_483     ),
    .col_in_484              ( u1_col_out_484     ),
    .col_in_485              ( u1_col_out_485     ),
    .col_in_486              ( u1_col_out_486     ),
    .col_in_487              ( u1_col_out_487     ),
    .col_in_488              ( u1_col_out_488     ),
    .col_in_489              ( u1_col_out_489     ),
    .col_in_490              ( u1_col_out_490     ),
    .col_in_491              ( u1_col_out_491     ),
    .col_in_492              ( u1_col_out_492     ),
    .col_in_493              ( u1_col_out_493     ),
    .col_in_494              ( u1_col_out_494     ),
    .col_in_495              ( u1_col_out_495     ),
    .col_in_496              ( u1_col_out_496     ),
    .col_in_497              ( u1_col_out_497     ),
    .col_in_498              ( u1_col_out_498     ),
    .col_in_499              ( u1_col_out_499     ),
    .col_in_500              ( u1_col_out_500     ),
    .col_in_501              ( u1_col_out_501     ),
    .col_in_502              ( u1_col_out_502     ),
    .col_in_503              ( u1_col_out_503     ),
    .col_in_504              ( u1_col_out_504     ),
    .col_in_505              ( u1_col_out_505     ),
    .col_in_506              ( u1_col_out_506     ),
    .col_in_507              ( u1_col_out_507     ),
    .col_in_508              ( u1_col_out_508     ),
    .col_in_509              ( u1_col_out_509     ),
    .col_in_510              ( u1_col_out_510     ),
    .col_in_511              ( u1_col_out_511     ),
    .col_in_512              ( u1_col_out_512     ),
    .col_in_513              ( u1_col_out_513     ),
    .col_in_514              ( u1_col_out_514     ),
    .col_in_515              ( u1_col_out_515     ),
    .col_in_516              ( u1_col_out_516     ),
    .col_in_517              ( u1_col_out_517     ),
    .col_in_518              ( u1_col_out_518     ),
    .col_in_519              ( u1_col_out_519     ),
    .col_in_520              ( u1_col_out_520     ),
    .col_in_521              ( u1_col_out_521     ),
    .col_in_522              ( u1_col_out_522     ),
    .col_in_523              ( u1_col_out_523     ),
    .col_in_524              ( u1_col_out_524     ),
    .col_in_525              ( u1_col_out_525     ),
    .col_in_526              ( u1_col_out_526     ),
    .col_in_527              ( u1_col_out_527     ),
    .col_in_528              ( u1_col_out_528     ),
    .col_in_529              ( u1_col_out_529     ),
    .col_in_530              ( u1_col_out_530     ),
    .col_in_531              ( u1_col_out_531     ),
    .col_in_532              ( u1_col_out_532     ),
    .col_in_533              ( u1_col_out_533     ),
    .col_in_534              ( u1_col_out_534     ),
    .col_in_535              ( u1_col_out_535     ),
    .col_in_536              ( u1_col_out_536     ),
    .col_in_537              ( u1_col_out_537     ),
    .col_in_538              ( u1_col_out_538     ),
    .col_in_539              ( u1_col_out_539     ),
    .col_in_540              ( u1_col_out_540     ),
    .col_in_541              ( u1_col_out_541     ),
    .col_in_542              ( u1_col_out_542     ),
    .col_in_543              ( u1_col_out_543     ),
    .col_in_544              ( u1_col_out_544     ),
    .col_in_545              ( u1_col_out_545     ),
    .col_in_546              ( u1_col_out_546     ),
    .col_in_547              ( u1_col_out_547     ),
    .col_in_548              ( u1_col_out_548     ),
    .col_in_549              ( u1_col_out_549     ),
    .col_in_550              ( u1_col_out_550     ),
    .col_in_551              ( u1_col_out_551     ),
    .col_in_552              ( u1_col_out_552     ),
    .col_in_553              ( u1_col_out_553     ),
    .col_in_554              ( u1_col_out_554     ),
    .col_in_555              ( u1_col_out_555     ),
    .col_in_556              ( u1_col_out_556     ),
    .col_in_557              ( u1_col_out_557     ),
    .col_in_558              ( u1_col_out_558     ),
    .col_in_559              ( u1_col_out_559     ),
    .col_in_560              ( u1_col_out_560     ),
    .col_in_561              ( u1_col_out_561     ),
    .col_in_562              ( u1_col_out_562     ),
    .col_in_563              ( u1_col_out_563     ),
    .col_in_564              ( u1_col_out_564     ),
    .col_in_565              ( u1_col_out_565     ),
    .col_in_566              ( u1_col_out_566     ),
    .col_in_567              ( u1_col_out_567     ),
    .col_in_568              ( u1_col_out_568     ),
    .col_in_569              ( u1_col_out_569     ),
    .col_in_570              ( u1_col_out_570     ),
    .col_in_571              ( u1_col_out_571     ),
    .col_in_572              ( u1_col_out_572     ),
    .col_in_573              ( u1_col_out_573     ),
    .col_in_574              ( u1_col_out_574     ),
    .col_in_575              ( u1_col_out_575     ),
    .col_in_576              ( u1_col_out_576     ),
    .col_in_577              ( u1_col_out_577     ),
    .col_in_578              ( u1_col_out_578     ),
    .col_in_579              ( u1_col_out_579     ),
    .col_in_580              ( u1_col_out_580     ),
    .col_in_581              ( u1_col_out_581     ),
    .col_in_582              ( u1_col_out_582     ),
    .col_in_583              ( u1_col_out_583     ),
    .col_in_584              ( u1_col_out_584     ),
    .col_in_585              ( u1_col_out_585     ),
    .col_in_586              ( u1_col_out_586     ),
    .col_in_587              ( u1_col_out_587     ),
    .col_in_588              ( u1_col_out_588     ),
    .col_in_589              ( u1_col_out_589     ),
    .col_in_590              ( u1_col_out_590     ),
    .col_in_591              ( u1_col_out_591     ),
    .col_in_592              ( u1_col_out_592     ),
    .col_in_593              ( u1_col_out_593     ),
    .col_in_594              ( u1_col_out_594     ),
    .col_in_595              ( u1_col_out_595     ),
    .col_in_596              ( u1_col_out_596     ),
    .col_in_597              ( u1_col_out_597     ),
    .col_in_598              ( u1_col_out_598     ),
    .col_in_599              ( u1_col_out_599     ),
    .col_in_600              ( u1_col_out_600     ),
    .col_in_601              ( u1_col_out_601     ),
    .col_in_602              ( u1_col_out_602     ),
    .col_in_603              ( u1_col_out_603     ),
    .col_in_604              ( u1_col_out_604     ),
    .col_in_605              ( u1_col_out_605     ),
    .col_in_606              ( u1_col_out_606     ),
    .col_in_607              ( u1_col_out_607     ),
    .col_in_608              ( u1_col_out_608     ),
    .col_in_609              ( u1_col_out_609     ),
    .col_in_610              ( u1_col_out_610     ),
    .col_in_611              ( u1_col_out_611     ),
    .col_in_612              ( u1_col_out_612     ),
    .col_in_613              ( u1_col_out_613     ),
    .col_in_614              ( u1_col_out_614     ),
    .col_in_615              ( u1_col_out_615     ),
    .col_in_616              ( u1_col_out_616     ),
    .col_in_617              ( u1_col_out_617     ),
    .col_in_618              ( u1_col_out_618     ),
    .col_in_619              ( u1_col_out_619     ),
    .col_in_620              ( u1_col_out_620     ),
    .col_in_621              ( u1_col_out_621     ),
    .col_in_622              ( u1_col_out_622     ),
    .col_in_623              ( u1_col_out_623     ),
    .col_in_624              ( u1_col_out_624     ),
    .col_in_625              ( u1_col_out_625     ),
    .col_in_626              ( u1_col_out_626     ),
    .col_in_627              ( u1_col_out_627     ),
    .col_in_628              ( u1_col_out_628     ),
    .col_in_629              ( u1_col_out_629     ),
    .col_in_630              ( u1_col_out_630     ),
    .col_in_631              ( u1_col_out_631     ),
    .col_in_632              ( u1_col_out_632     ),
    .col_in_633              ( u1_col_out_633     ),
    .col_in_634              ( u1_col_out_634     ),
    .col_in_635              ( u1_col_out_635     ),
    .col_in_636              ( u1_col_out_636     ),
    .col_in_637              ( u1_col_out_637     ),
    .col_in_638              ( u1_col_out_638     ),
    .col_in_639              ( u1_col_out_639     ),
    .col_in_640              ( u1_col_out_640     ),
    .col_in_641              ( u1_col_out_641     ),
    .col_in_642              ( u1_col_out_642     ),
    .col_in_643              ( u1_col_out_643     ),
    .col_in_644              ( u1_col_out_644     ),
    .col_in_645              ( u1_col_out_645     ),
    .col_in_646              ( u1_col_out_646     ),
    .col_in_647              ( u1_col_out_647     ),
    .col_in_648              ( u1_col_out_648     ),
    .col_in_649              ( u1_col_out_649     ),
    .col_in_650              ( u1_col_out_650     ),
    .col_in_651              ( u1_col_out_651     ),
    .col_in_652              ( u1_col_out_652     ),
    .col_in_653              ( u1_col_out_653     ),
    .col_in_654              ( u1_col_out_654     ),
    .col_in_655              ( u1_col_out_655     ),
    .col_in_656              ( u1_col_out_656     ),
    .col_in_657              ( u1_col_out_657     ),
    .col_in_658              ( u1_col_out_658     ),
    .col_in_659              ( u1_col_out_659     ),
    .col_in_660              ( u1_col_out_660     ),
    .col_in_661              ( u1_col_out_661     ),
    .col_in_662              ( u1_col_out_662     ),
    .col_in_663              ( u1_col_out_663     ),
    .col_in_664              ( u1_col_out_664     ),
    .col_in_665              ( u1_col_out_665     ),
    .col_in_666              ( u1_col_out_666     ),
    .col_in_667              ( u1_col_out_667     ),
    .col_in_668              ( u1_col_out_668     ),
    .col_in_669              ( u1_col_out_669     ),
    .col_in_670              ( u1_col_out_670     ),
    .col_in_671              ( u1_col_out_671     ),
    .col_in_672              ( u1_col_out_672     ),
    .col_in_673              ( u1_col_out_673     ),
    .col_in_674              ( u1_col_out_674     ),
    .col_in_675              ( u1_col_out_675     ),
    .col_in_676              ( u1_col_out_676     ),
    .col_in_677              ( u1_col_out_677     ),
    .col_in_678              ( u1_col_out_678     ),
    .col_in_679              ( u1_col_out_679     ),
    .col_in_680              ( u1_col_out_680     ),
    .col_in_681              ( u1_col_out_681     ),
    .col_in_682              ( u1_col_out_682     ),
    .col_in_683              ( u1_col_out_683     ),
    .col_in_684              ( u1_col_out_684     ),
    .col_in_685              ( u1_col_out_685     ),
    .col_in_686              ( u1_col_out_686     ),
    .col_in_687              ( u1_col_out_687     ),
    .col_in_688              ( u1_col_out_688     ),
    .col_in_689              ( u1_col_out_689     ),
    .col_in_690              ( u1_col_out_690     ),
    .col_in_691              ( u1_col_out_691     ),
    .col_in_692              ( u1_col_out_692     ),
    .col_in_693              ( u1_col_out_693     ),
    .col_in_694              ( u1_col_out_694     ),
    .col_in_695              ( u1_col_out_695     ),
    .col_in_696              ( u1_col_out_696     ),
    .col_in_697              ( u1_col_out_697     ),
    .col_in_698              ( u1_col_out_698     ),
    .col_in_699              ( u1_col_out_699     ),
    .col_in_700              ( u1_col_out_700     ),
    .col_in_701              ( u1_col_out_701     ),
    .col_in_702              ( u1_col_out_702     ),
    .col_in_703              ( u1_col_out_703     ),
    .col_in_704              ( u1_col_out_704     ),
    .col_in_705              ( u1_col_out_705     ),
    .col_in_706              ( u1_col_out_706     ),
    .col_in_707              ( u1_col_out_707     ),
    .col_in_708              ( u1_col_out_708     ),
    .col_in_709              ( u1_col_out_709     ),
    .col_in_710              ( u1_col_out_710     ),
    .col_in_711              ( u1_col_out_711     ),
    .col_in_712              ( u1_col_out_712     ),
    .col_in_713              ( u1_col_out_713     ),
    .col_in_714              ( u1_col_out_714     ),
    .col_in_715              ( u1_col_out_715     ),
    .col_in_716              ( u1_col_out_716     ),
    .col_in_717              ( u1_col_out_717     ),
    .col_in_718              ( u1_col_out_718     ),
    .col_in_719              ( u1_col_out_719     ),
    .col_in_720              ( u1_col_out_720     ),
    .col_in_721              ( u1_col_out_721     ),
    .col_in_722              ( u1_col_out_722     ),
    .col_in_723              ( u1_col_out_723     ),
    .col_in_724              ( u1_col_out_724     ),
    .col_in_725              ( u1_col_out_725     ),
    .col_in_726              ( u1_col_out_726     ),
    .col_in_727              ( u1_col_out_727     ),
    .col_in_728              ( u1_col_out_728     ),
    .col_in_729              ( u1_col_out_729     ),
    .col_in_730              ( u1_col_out_730     ),
    .col_in_731              ( u1_col_out_731     ),
    .col_in_732              ( u1_col_out_732     ),
    .col_in_733              ( u1_col_out_733     ),
    .col_in_734              ( u1_col_out_734     ),
    .col_in_735              ( u1_col_out_735     ),
    .col_in_736              ( u1_col_out_736     ),
    .col_in_737              ( u1_col_out_737     ),
    .col_in_738              ( u1_col_out_738     ),
    .col_in_739              ( u1_col_out_739     ),
    .col_in_740              ( u1_col_out_740     ),
    .col_in_741              ( u1_col_out_741     ),
    .col_in_742              ( u1_col_out_742     ),
    .col_in_743              ( u1_col_out_743     ),
    .col_in_744              ( u1_col_out_744     ),
    .col_in_745              ( u1_col_out_745     ),
    .col_in_746              ( u1_col_out_746     ),
    .col_in_747              ( u1_col_out_747     ),
    .col_in_748              ( u1_col_out_748     ),
    .col_in_749              ( u1_col_out_749     ),
    .col_in_750              ( u1_col_out_750     ),
    .col_in_751              ( u1_col_out_751     ),
    .col_in_752              ( u1_col_out_752     ),
    .col_in_753              ( u1_col_out_753     ),
    .col_in_754              ( u1_col_out_754     ),
    .col_in_755              ( u1_col_out_755     ),
    .col_in_756              ( u1_col_out_756     ),
    .col_in_757              ( u1_col_out_757     ),
    .col_in_758              ( u1_col_out_758     ),
    .col_in_759              ( u1_col_out_759     ),
    .col_in_760              ( u1_col_out_760     ),
    .col_in_761              ( u1_col_out_761     ),
    .col_in_762              ( u1_col_out_762     ),
    .col_in_763              ( u1_col_out_763     ),
    .col_in_764              ( u1_col_out_764     ),
    .col_in_765              ( u1_col_out_765     ),
    .col_in_766              ( u1_col_out_766     ),
    .col_in_767              ( u1_col_out_767     ),
    .col_in_768              ( u1_col_out_768     ),
    .col_in_769              ( u1_col_out_769     ),
    .col_in_770              ( u1_col_out_770     ),
    .col_in_771              ( u1_col_out_771     ),
    .col_in_772              ( u1_col_out_772     ),
    .col_in_773              ( u1_col_out_773     ),
    .col_in_774              ( u1_col_out_774     ),
    .col_in_775              ( u1_col_out_775     ),
    .col_in_776              ( u1_col_out_776     ),
    .col_in_777              ( u1_col_out_777     ),
    .col_in_778              ( u1_col_out_778     ),
    .col_in_779              ( u1_col_out_779     ),
    .col_in_780              ( u1_col_out_780     ),
    .col_in_781              ( u1_col_out_781     ),
    .col_in_782              ( u1_col_out_782     ),
    .col_in_783              ( u1_col_out_783     ),
    .col_in_784              ( u1_col_out_784     ),
    .col_in_785              ( u1_col_out_785     ),
    .col_in_786              ( u1_col_out_786     ),
    .col_in_787              ( u1_col_out_787     ),
    .col_in_788              ( u1_col_out_788     ),
    .col_in_789              ( u1_col_out_789     ),
    .col_in_790              ( u1_col_out_790     ),
    .col_in_791              ( u1_col_out_791     ),
    .col_in_792              ( u1_col_out_792     ),
    .col_in_793              ( u1_col_out_793     ),
    .col_in_794              ( u1_col_out_794     ),
    .col_in_795              ( u1_col_out_795     ),
    .col_in_796              ( u1_col_out_796     ),
    .col_in_797              ( u1_col_out_797     ),
    .col_in_798              ( u1_col_out_798     ),
    .col_in_799              ( u1_col_out_799     ),
    .col_in_800              ( u1_col_out_800     ),
    .col_in_801              ( u1_col_out_801     ),
    .col_in_802              ( u1_col_out_802     ),
    .col_in_803              ( u1_col_out_803     ),
    .col_in_804              ( u1_col_out_804     ),
    .col_in_805              ( u1_col_out_805     ),
    .col_in_806              ( u1_col_out_806     ),
    .col_in_807              ( u1_col_out_807     ),
    .col_in_808              ( u1_col_out_808     ),
    .col_in_809              ( u1_col_out_809     ),
    .col_in_810              ( u1_col_out_810     ),
    .col_in_811              ( u1_col_out_811     ),
    .col_in_812              ( u1_col_out_812     ),
    .col_in_813              ( u1_col_out_813     ),
    .col_in_814              ( u1_col_out_814     ),
    .col_in_815              ( u1_col_out_815     ),
    .col_in_816              ( u1_col_out_816     ),
    .col_in_817              ( u1_col_out_817     ),
    .col_in_818              ( u1_col_out_818     ),
    .col_in_819              ( u1_col_out_819     ),
    .col_in_820              ( u1_col_out_820     ),
    .col_in_821              ( u1_col_out_821     ),
    .col_in_822              ( u1_col_out_822     ),
    .col_in_823              ( u1_col_out_823     ),
    .col_in_824              ( u1_col_out_824     ),
    .col_in_825              ( u1_col_out_825     ),
    .col_in_826              ( u1_col_out_826     ),
    .col_in_827              ( u1_col_out_827     ),
    .col_in_828              ( u1_col_out_828     ),
    .col_in_829              ( u1_col_out_829     ),
    .col_in_830              ( u1_col_out_830     ),
    .col_in_831              ( u1_col_out_831     ),
    .col_in_832              ( u1_col_out_832     ),
    .col_in_833              ( u1_col_out_833     ),
    .col_in_834              ( u1_col_out_834     ),
    .col_in_835              ( u1_col_out_835     ),
    .col_in_836              ( u1_col_out_836     ),
    .col_in_837              ( u1_col_out_837     ),
    .col_in_838              ( u1_col_out_838     ),
    .col_in_839              ( u1_col_out_839     ),
    .col_in_840              ( u1_col_out_840     ),
    .col_in_841              ( u1_col_out_841     ),
    .col_in_842              ( u1_col_out_842     ),
    .col_in_843              ( u1_col_out_843     ),
    .col_in_844              ( u1_col_out_844     ),
    .col_in_845              ( u1_col_out_845     ),
    .col_in_846              ( u1_col_out_846     ),
    .col_in_847              ( u1_col_out_847     ),
    .col_in_848              ( u1_col_out_848     ),
    .col_in_849              ( u1_col_out_849     ),
    .col_in_850              ( u1_col_out_850     ),
    .col_in_851              ( u1_col_out_851     ),
    .col_in_852              ( u1_col_out_852     ),
    .col_in_853              ( u1_col_out_853     ),
    .col_in_854              ( u1_col_out_854     ),
    .col_in_855              ( u1_col_out_855     ),
    .col_in_856              ( u1_col_out_856     ),
    .col_in_857              ( u1_col_out_857     ),
    .col_in_858              ( u1_col_out_858     ),
    .col_in_859              ( u1_col_out_859     ),
    .col_in_860              ( u1_col_out_860     ),
    .col_in_861              ( u1_col_out_861     ),
    .col_in_862              ( u1_col_out_862     ),
    .col_in_863              ( u1_col_out_863     ),
    .col_in_864              ( u1_col_out_864     ),
    .col_in_865              ( u1_col_out_865     ),
    .col_in_866              ( u1_col_out_866     ),
    .col_in_867              ( u1_col_out_867     ),
    .col_in_868              ( u1_col_out_868     ),
    .col_in_869              ( u1_col_out_869     ),
    .col_in_870              ( u1_col_out_870     ),
    .col_in_871              ( u1_col_out_871     ),
    .col_in_872              ( u1_col_out_872     ),
    .col_in_873              ( u1_col_out_873     ),
    .col_in_874              ( u1_col_out_874     ),
    .col_in_875              ( u1_col_out_875     ),
    .col_in_876              ( u1_col_out_876     ),
    .col_in_877              ( u1_col_out_877     ),
    .col_in_878              ( u1_col_out_878     ),
    .col_in_879              ( u1_col_out_879     ),
    .col_in_880              ( u1_col_out_880     ),
    .col_in_881              ( u1_col_out_881     ),
    .col_in_882              ( u1_col_out_882     ),
    .col_in_883              ( u1_col_out_883     ),
    .col_in_884              ( u1_col_out_884     ),
    .col_in_885              ( u1_col_out_885     ),
    .col_in_886              ( u1_col_out_886     ),
    .col_in_887              ( u1_col_out_887     ),
    .col_in_888              ( u1_col_out_888     ),
    .col_in_889              ( u1_col_out_889     ),
    .col_in_890              ( u1_col_out_890     ),
    .col_in_891              ( u1_col_out_891     ),
    .col_in_892              ( u1_col_out_892     ),
    .col_in_893              ( u1_col_out_893     ),
    .col_in_894              ( u1_col_out_894     ),
    .col_in_895              ( u1_col_out_895     ),
    .col_in_896              ( u1_col_out_896     ),
    .col_in_897              ( u1_col_out_897     ),
    .col_in_898              ( u1_col_out_898     ),
    .col_in_899              ( u1_col_out_899     ),
    .col_in_900              ( u1_col_out_900     ),
    .col_in_901              ( u1_col_out_901     ),
    .col_in_902              ( u1_col_out_902     ),
    .col_in_903              ( u1_col_out_903     ),
    .col_in_904              ( u1_col_out_904     ),
    .col_in_905              ( u1_col_out_905     ),
    .col_in_906              ( u1_col_out_906     ),
    .col_in_907              ( u1_col_out_907     ),
    .col_in_908              ( u1_col_out_908     ),
    .col_in_909              ( u1_col_out_909     ),
    .col_in_910              ( u1_col_out_910     ),
    .col_in_911              ( u1_col_out_911     ),
    .col_in_912              ( u1_col_out_912     ),
    .col_in_913              ( u1_col_out_913     ),
    .col_in_914              ( u1_col_out_914     ),
    .col_in_915              ( u1_col_out_915     ),
    .col_in_916              ( u1_col_out_916     ),
    .col_in_917              ( u1_col_out_917     ),
    .col_in_918              ( u1_col_out_918     ),
    .col_in_919              ( u1_col_out_919     ),
    .col_in_920              ( u1_col_out_920     ),
    .col_in_921              ( u1_col_out_921     ),
    .col_in_922              ( u1_col_out_922     ),
    .col_in_923              ( u1_col_out_923     ),
    .col_in_924              ( u1_col_out_924     ),
    .col_in_925              ( u1_col_out_925     ),
    .col_in_926              ( u1_col_out_926     ),
    .col_in_927              ( u1_col_out_927     ),
    .col_in_928              ( u1_col_out_928     ),
    .col_in_929              ( u1_col_out_929     ),
    .col_in_930              ( u1_col_out_930     ),
    .col_in_931              ( u1_col_out_931     ),
    .col_in_932              ( u1_col_out_932     ),
    .col_in_933              ( u1_col_out_933     ),
    .col_in_934              ( u1_col_out_934     ),
    .col_in_935              ( u1_col_out_935     ),
    .col_in_936              ( u1_col_out_936     ),
    .col_in_937              ( u1_col_out_937     ),
    .col_in_938              ( u1_col_out_938     ),
    .col_in_939              ( u1_col_out_939     ),
    .col_in_940              ( u1_col_out_940     ),
    .col_in_941              ( u1_col_out_941     ),
    .col_in_942              ( u1_col_out_942     ),
    .col_in_943              ( u1_col_out_943     ),
    .col_in_944              ( u1_col_out_944     ),
    .col_in_945              ( u1_col_out_945     ),
    .col_in_946              ( u1_col_out_946     ),
    .col_in_947              ( u1_col_out_947     ),
    .col_in_948              ( u1_col_out_948     ),
    .col_in_949              ( u1_col_out_949     ),
    .col_in_950              ( u1_col_out_950     ),
    .col_in_951              ( u1_col_out_951     ),
    .col_in_952              ( u1_col_out_952     ),
    .col_in_953              ( u1_col_out_953     ),
    .col_in_954              ( u1_col_out_954     ),
    .col_in_955              ( u1_col_out_955     ),
    .col_in_956              ( u1_col_out_956     ),
    .col_in_957              ( u1_col_out_957     ),
    .col_in_958              ( u1_col_out_958     ),
    .col_in_959              ( u1_col_out_959     ),
    .col_in_960              ( u1_col_out_960     ),
    .col_in_961              ( u1_col_out_961     ),
    .col_in_962              ( u1_col_out_962     ),
    .col_in_963              ( u1_col_out_963     ),
    .col_in_964              ( u1_col_out_964     ),
    .col_in_965              ( u1_col_out_965     ),
    .col_in_966              ( u1_col_out_966     ),
    .col_in_967              ( u1_col_out_967     ),
    .col_in_968              ( u1_col_out_968     ),
    .col_in_969              ( u1_col_out_969     ),
    .col_in_970              ( u1_col_out_970     ),
    .col_in_971              ( u1_col_out_971     ),
    .col_in_972              ( u1_col_out_972     ),
    .col_in_973              ( u1_col_out_973     ),
    .col_in_974              ( u1_col_out_974     ),
    .col_in_975              ( u1_col_out_975     ),
    .col_in_976              ( u1_col_out_976     ),
    .col_in_977              ( u1_col_out_977     ),
    .col_in_978              ( u1_col_out_978     ),
    .col_in_979              ( u1_col_out_979     ),
    .col_in_980              ( u1_col_out_980     ),
    .col_in_981              ( u1_col_out_981     ),
    .col_in_982              ( u1_col_out_982     ),
    .col_in_983              ( u1_col_out_983     ),
    .col_in_984              ( u1_col_out_984     ),
    .col_in_985              ( u1_col_out_985     ),
    .col_in_986              ( u1_col_out_986     ),
    .col_in_987              ( u1_col_out_987     ),
    .col_in_988              ( u1_col_out_988     ),
    .col_in_989              ( u1_col_out_989     ),
    .col_in_990              ( u1_col_out_990     ),
    .col_in_991              ( u1_col_out_991     ),
    .col_in_992              ( u1_col_out_992     ),
    .col_in_993              ( u1_col_out_993     ),
    .col_in_994              ( u1_col_out_994     ),
    .col_in_995              ( u1_col_out_995     ),
    .col_in_996              ( u1_col_out_996     ),
    .col_in_997              ( u1_col_out_997     ),
    .col_in_998              ( u1_col_out_998     ),
    .col_in_999              ( u1_col_out_999     ),
    .col_in_1000             ( u1_col_out_1000    ),
    .col_in_1001             ( u1_col_out_1001    ),
    .col_in_1002             ( u1_col_out_1002    ),
    .col_in_1003             ( u1_col_out_1003    ),
    .col_in_1004             ( u1_col_out_1004    ),
    .col_in_1005             ( u1_col_out_1005    ),
    .col_in_1006             ( u1_col_out_1006    ),
    .col_in_1007             ( u1_col_out_1007    ),
    .col_in_1008             ( u1_col_out_1008    ),
    .col_in_1009             ( u1_col_out_1009    ),
    .col_in_1010             ( u1_col_out_1010    ),
    .col_in_1011             ( u1_col_out_1011    ),
    .col_in_1012             ( u1_col_out_1012    ),
    .col_in_1013             ( u1_col_out_1013    ),
    .col_in_1014             ( u1_col_out_1014    ),
    .col_in_1015             ( u1_col_out_1015    ),
    .col_in_1016             ( u1_col_out_1016    ),
    .col_in_1017             ( u1_col_out_1017    ),
    .col_in_1018             ( u1_col_out_1018    ),
    .col_in_1019             ( u1_col_out_1019    ),
    .col_in_1020             ( u1_col_out_1020    ),
    .col_in_1021             ( u1_col_out_1021    ),
    .col_in_1022             ( u1_col_out_1022    ),
    .col_in_1023             ( u1_col_out_1023    ),
    .col_in_1024             ( u1_col_out_1024    ),
    .col_in_1025             ( u1_col_out_1025    ),
    .col_in_1026             ( u1_col_out_1026    ),
    .col_in_1027             ( u1_col_out_1027    ),
    .col_in_1028             ( u1_col_out_1028    ),
    .col_in_1029             ( u1_col_out_1029    ),
    .col_in_1030             ( u1_col_out_1030    ),
    .col_in_1031             ( u1_col_out_1031    ),
    .col_in_1032             ( u1_col_out_1032    ),

    .col_out_0               ( u2_col_out_0      ),
    .col_out_1               ( u2_col_out_1      ),
    .col_out_2               ( u2_col_out_2      ),
    .col_out_3               ( u2_col_out_3      ),
    .col_out_4               ( u2_col_out_4      ),
    .col_out_5               ( u2_col_out_5      ),
    .col_out_6               ( u2_col_out_6      ),
    .col_out_7               ( u2_col_out_7      ),
    .col_out_8               ( u2_col_out_8      ),
    .col_out_9               ( u2_col_out_9      ),
    .col_out_10              ( u2_col_out_10     ),
    .col_out_11              ( u2_col_out_11     ),
    .col_out_12              ( u2_col_out_12     ),
    .col_out_13              ( u2_col_out_13     ),
    .col_out_14              ( u2_col_out_14     ),
    .col_out_15              ( u2_col_out_15     ),
    .col_out_16              ( u2_col_out_16     ),
    .col_out_17              ( u2_col_out_17     ),
    .col_out_18              ( u2_col_out_18     ),
    .col_out_19              ( u2_col_out_19     ),
    .col_out_20              ( u2_col_out_20     ),
    .col_out_21              ( u2_col_out_21     ),
    .col_out_22              ( u2_col_out_22     ),
    .col_out_23              ( u2_col_out_23     ),
    .col_out_24              ( u2_col_out_24     ),
    .col_out_25              ( u2_col_out_25     ),
    .col_out_26              ( u2_col_out_26     ),
    .col_out_27              ( u2_col_out_27     ),
    .col_out_28              ( u2_col_out_28     ),
    .col_out_29              ( u2_col_out_29     ),
    .col_out_30              ( u2_col_out_30     ),
    .col_out_31              ( u2_col_out_31     ),
    .col_out_32              ( u2_col_out_32     ),
    .col_out_33              ( u2_col_out_33     ),
    .col_out_34              ( u2_col_out_34     ),
    .col_out_35              ( u2_col_out_35     ),
    .col_out_36              ( u2_col_out_36     ),
    .col_out_37              ( u2_col_out_37     ),
    .col_out_38              ( u2_col_out_38     ),
    .col_out_39              ( u2_col_out_39     ),
    .col_out_40              ( u2_col_out_40     ),
    .col_out_41              ( u2_col_out_41     ),
    .col_out_42              ( u2_col_out_42     ),
    .col_out_43              ( u2_col_out_43     ),
    .col_out_44              ( u2_col_out_44     ),
    .col_out_45              ( u2_col_out_45     ),
    .col_out_46              ( u2_col_out_46     ),
    .col_out_47              ( u2_col_out_47     ),
    .col_out_48              ( u2_col_out_48     ),
    .col_out_49              ( u2_col_out_49     ),
    .col_out_50              ( u2_col_out_50     ),
    .col_out_51              ( u2_col_out_51     ),
    .col_out_52              ( u2_col_out_52     ),
    .col_out_53              ( u2_col_out_53     ),
    .col_out_54              ( u2_col_out_54     ),
    .col_out_55              ( u2_col_out_55     ),
    .col_out_56              ( u2_col_out_56     ),
    .col_out_57              ( u2_col_out_57     ),
    .col_out_58              ( u2_col_out_58     ),
    .col_out_59              ( u2_col_out_59     ),
    .col_out_60              ( u2_col_out_60     ),
    .col_out_61              ( u2_col_out_61     ),
    .col_out_62              ( u2_col_out_62     ),
    .col_out_63              ( u2_col_out_63     ),
    .col_out_64              ( u2_col_out_64     ),
    .col_out_65              ( u2_col_out_65     ),
    .col_out_66              ( u2_col_out_66     ),
    .col_out_67              ( u2_col_out_67     ),
    .col_out_68              ( u2_col_out_68     ),
    .col_out_69              ( u2_col_out_69     ),
    .col_out_70              ( u2_col_out_70     ),
    .col_out_71              ( u2_col_out_71     ),
    .col_out_72              ( u2_col_out_72     ),
    .col_out_73              ( u2_col_out_73     ),
    .col_out_74              ( u2_col_out_74     ),
    .col_out_75              ( u2_col_out_75     ),
    .col_out_76              ( u2_col_out_76     ),
    .col_out_77              ( u2_col_out_77     ),
    .col_out_78              ( u2_col_out_78     ),
    .col_out_79              ( u2_col_out_79     ),
    .col_out_80              ( u2_col_out_80     ),
    .col_out_81              ( u2_col_out_81     ),
    .col_out_82              ( u2_col_out_82     ),
    .col_out_83              ( u2_col_out_83     ),
    .col_out_84              ( u2_col_out_84     ),
    .col_out_85              ( u2_col_out_85     ),
    .col_out_86              ( u2_col_out_86     ),
    .col_out_87              ( u2_col_out_87     ),
    .col_out_88              ( u2_col_out_88     ),
    .col_out_89              ( u2_col_out_89     ),
    .col_out_90              ( u2_col_out_90     ),
    .col_out_91              ( u2_col_out_91     ),
    .col_out_92              ( u2_col_out_92     ),
    .col_out_93              ( u2_col_out_93     ),
    .col_out_94              ( u2_col_out_94     ),
    .col_out_95              ( u2_col_out_95     ),
    .col_out_96              ( u2_col_out_96     ),
    .col_out_97              ( u2_col_out_97     ),
    .col_out_98              ( u2_col_out_98     ),
    .col_out_99              ( u2_col_out_99     ),
    .col_out_100             ( u2_col_out_100    ),
    .col_out_101             ( u2_col_out_101    ),
    .col_out_102             ( u2_col_out_102    ),
    .col_out_103             ( u2_col_out_103    ),
    .col_out_104             ( u2_col_out_104    ),
    .col_out_105             ( u2_col_out_105    ),
    .col_out_106             ( u2_col_out_106    ),
    .col_out_107             ( u2_col_out_107    ),
    .col_out_108             ( u2_col_out_108    ),
    .col_out_109             ( u2_col_out_109    ),
    .col_out_110             ( u2_col_out_110    ),
    .col_out_111             ( u2_col_out_111    ),
    .col_out_112             ( u2_col_out_112    ),
    .col_out_113             ( u2_col_out_113    ),
    .col_out_114             ( u2_col_out_114    ),
    .col_out_115             ( u2_col_out_115    ),
    .col_out_116             ( u2_col_out_116    ),
    .col_out_117             ( u2_col_out_117    ),
    .col_out_118             ( u2_col_out_118    ),
    .col_out_119             ( u2_col_out_119    ),
    .col_out_120             ( u2_col_out_120    ),
    .col_out_121             ( u2_col_out_121    ),
    .col_out_122             ( u2_col_out_122    ),
    .col_out_123             ( u2_col_out_123    ),
    .col_out_124             ( u2_col_out_124    ),
    .col_out_125             ( u2_col_out_125    ),
    .col_out_126             ( u2_col_out_126    ),
    .col_out_127             ( u2_col_out_127    ),
    .col_out_128             ( u2_col_out_128    ),
    .col_out_129             ( u2_col_out_129    ),
    .col_out_130             ( u2_col_out_130    ),
    .col_out_131             ( u2_col_out_131    ),
    .col_out_132             ( u2_col_out_132    ),
    .col_out_133             ( u2_col_out_133    ),
    .col_out_134             ( u2_col_out_134    ),
    .col_out_135             ( u2_col_out_135    ),
    .col_out_136             ( u2_col_out_136    ),
    .col_out_137             ( u2_col_out_137    ),
    .col_out_138             ( u2_col_out_138    ),
    .col_out_139             ( u2_col_out_139    ),
    .col_out_140             ( u2_col_out_140    ),
    .col_out_141             ( u2_col_out_141    ),
    .col_out_142             ( u2_col_out_142    ),
    .col_out_143             ( u2_col_out_143    ),
    .col_out_144             ( u2_col_out_144    ),
    .col_out_145             ( u2_col_out_145    ),
    .col_out_146             ( u2_col_out_146    ),
    .col_out_147             ( u2_col_out_147    ),
    .col_out_148             ( u2_col_out_148    ),
    .col_out_149             ( u2_col_out_149    ),
    .col_out_150             ( u2_col_out_150    ),
    .col_out_151             ( u2_col_out_151    ),
    .col_out_152             ( u2_col_out_152    ),
    .col_out_153             ( u2_col_out_153    ),
    .col_out_154             ( u2_col_out_154    ),
    .col_out_155             ( u2_col_out_155    ),
    .col_out_156             ( u2_col_out_156    ),
    .col_out_157             ( u2_col_out_157    ),
    .col_out_158             ( u2_col_out_158    ),
    .col_out_159             ( u2_col_out_159    ),
    .col_out_160             ( u2_col_out_160    ),
    .col_out_161             ( u2_col_out_161    ),
    .col_out_162             ( u2_col_out_162    ),
    .col_out_163             ( u2_col_out_163    ),
    .col_out_164             ( u2_col_out_164    ),
    .col_out_165             ( u2_col_out_165    ),
    .col_out_166             ( u2_col_out_166    ),
    .col_out_167             ( u2_col_out_167    ),
    .col_out_168             ( u2_col_out_168    ),
    .col_out_169             ( u2_col_out_169    ),
    .col_out_170             ( u2_col_out_170    ),
    .col_out_171             ( u2_col_out_171    ),
    .col_out_172             ( u2_col_out_172    ),
    .col_out_173             ( u2_col_out_173    ),
    .col_out_174             ( u2_col_out_174    ),
    .col_out_175             ( u2_col_out_175    ),
    .col_out_176             ( u2_col_out_176    ),
    .col_out_177             ( u2_col_out_177    ),
    .col_out_178             ( u2_col_out_178    ),
    .col_out_179             ( u2_col_out_179    ),
    .col_out_180             ( u2_col_out_180    ),
    .col_out_181             ( u2_col_out_181    ),
    .col_out_182             ( u2_col_out_182    ),
    .col_out_183             ( u2_col_out_183    ),
    .col_out_184             ( u2_col_out_184    ),
    .col_out_185             ( u2_col_out_185    ),
    .col_out_186             ( u2_col_out_186    ),
    .col_out_187             ( u2_col_out_187    ),
    .col_out_188             ( u2_col_out_188    ),
    .col_out_189             ( u2_col_out_189    ),
    .col_out_190             ( u2_col_out_190    ),
    .col_out_191             ( u2_col_out_191    ),
    .col_out_192             ( u2_col_out_192    ),
    .col_out_193             ( u2_col_out_193    ),
    .col_out_194             ( u2_col_out_194    ),
    .col_out_195             ( u2_col_out_195    ),
    .col_out_196             ( u2_col_out_196    ),
    .col_out_197             ( u2_col_out_197    ),
    .col_out_198             ( u2_col_out_198    ),
    .col_out_199             ( u2_col_out_199    ),
    .col_out_200             ( u2_col_out_200    ),
    .col_out_201             ( u2_col_out_201    ),
    .col_out_202             ( u2_col_out_202    ),
    .col_out_203             ( u2_col_out_203    ),
    .col_out_204             ( u2_col_out_204    ),
    .col_out_205             ( u2_col_out_205    ),
    .col_out_206             ( u2_col_out_206    ),
    .col_out_207             ( u2_col_out_207    ),
    .col_out_208             ( u2_col_out_208    ),
    .col_out_209             ( u2_col_out_209    ),
    .col_out_210             ( u2_col_out_210    ),
    .col_out_211             ( u2_col_out_211    ),
    .col_out_212             ( u2_col_out_212    ),
    .col_out_213             ( u2_col_out_213    ),
    .col_out_214             ( u2_col_out_214    ),
    .col_out_215             ( u2_col_out_215    ),
    .col_out_216             ( u2_col_out_216    ),
    .col_out_217             ( u2_col_out_217    ),
    .col_out_218             ( u2_col_out_218    ),
    .col_out_219             ( u2_col_out_219    ),
    .col_out_220             ( u2_col_out_220    ),
    .col_out_221             ( u2_col_out_221    ),
    .col_out_222             ( u2_col_out_222    ),
    .col_out_223             ( u2_col_out_223    ),
    .col_out_224             ( u2_col_out_224    ),
    .col_out_225             ( u2_col_out_225    ),
    .col_out_226             ( u2_col_out_226    ),
    .col_out_227             ( u2_col_out_227    ),
    .col_out_228             ( u2_col_out_228    ),
    .col_out_229             ( u2_col_out_229    ),
    .col_out_230             ( u2_col_out_230    ),
    .col_out_231             ( u2_col_out_231    ),
    .col_out_232             ( u2_col_out_232    ),
    .col_out_233             ( u2_col_out_233    ),
    .col_out_234             ( u2_col_out_234    ),
    .col_out_235             ( u2_col_out_235    ),
    .col_out_236             ( u2_col_out_236    ),
    .col_out_237             ( u2_col_out_237    ),
    .col_out_238             ( u2_col_out_238    ),
    .col_out_239             ( u2_col_out_239    ),
    .col_out_240             ( u2_col_out_240    ),
    .col_out_241             ( u2_col_out_241    ),
    .col_out_242             ( u2_col_out_242    ),
    .col_out_243             ( u2_col_out_243    ),
    .col_out_244             ( u2_col_out_244    ),
    .col_out_245             ( u2_col_out_245    ),
    .col_out_246             ( u2_col_out_246    ),
    .col_out_247             ( u2_col_out_247    ),
    .col_out_248             ( u2_col_out_248    ),
    .col_out_249             ( u2_col_out_249    ),
    .col_out_250             ( u2_col_out_250    ),
    .col_out_251             ( u2_col_out_251    ),
    .col_out_252             ( u2_col_out_252    ),
    .col_out_253             ( u2_col_out_253    ),
    .col_out_254             ( u2_col_out_254    ),
    .col_out_255             ( u2_col_out_255    ),
    .col_out_256             ( u2_col_out_256    ),
    .col_out_257             ( u2_col_out_257    ),
    .col_out_258             ( u2_col_out_258    ),
    .col_out_259             ( u2_col_out_259    ),
    .col_out_260             ( u2_col_out_260    ),
    .col_out_261             ( u2_col_out_261    ),
    .col_out_262             ( u2_col_out_262    ),
    .col_out_263             ( u2_col_out_263    ),
    .col_out_264             ( u2_col_out_264    ),
    .col_out_265             ( u2_col_out_265    ),
    .col_out_266             ( u2_col_out_266    ),
    .col_out_267             ( u2_col_out_267    ),
    .col_out_268             ( u2_col_out_268    ),
    .col_out_269             ( u2_col_out_269    ),
    .col_out_270             ( u2_col_out_270    ),
    .col_out_271             ( u2_col_out_271    ),
    .col_out_272             ( u2_col_out_272    ),
    .col_out_273             ( u2_col_out_273    ),
    .col_out_274             ( u2_col_out_274    ),
    .col_out_275             ( u2_col_out_275    ),
    .col_out_276             ( u2_col_out_276    ),
    .col_out_277             ( u2_col_out_277    ),
    .col_out_278             ( u2_col_out_278    ),
    .col_out_279             ( u2_col_out_279    ),
    .col_out_280             ( u2_col_out_280    ),
    .col_out_281             ( u2_col_out_281    ),
    .col_out_282             ( u2_col_out_282    ),
    .col_out_283             ( u2_col_out_283    ),
    .col_out_284             ( u2_col_out_284    ),
    .col_out_285             ( u2_col_out_285    ),
    .col_out_286             ( u2_col_out_286    ),
    .col_out_287             ( u2_col_out_287    ),
    .col_out_288             ( u2_col_out_288    ),
    .col_out_289             ( u2_col_out_289    ),
    .col_out_290             ( u2_col_out_290    ),
    .col_out_291             ( u2_col_out_291    ),
    .col_out_292             ( u2_col_out_292    ),
    .col_out_293             ( u2_col_out_293    ),
    .col_out_294             ( u2_col_out_294    ),
    .col_out_295             ( u2_col_out_295    ),
    .col_out_296             ( u2_col_out_296    ),
    .col_out_297             ( u2_col_out_297    ),
    .col_out_298             ( u2_col_out_298    ),
    .col_out_299             ( u2_col_out_299    ),
    .col_out_300             ( u2_col_out_300    ),
    .col_out_301             ( u2_col_out_301    ),
    .col_out_302             ( u2_col_out_302    ),
    .col_out_303             ( u2_col_out_303    ),
    .col_out_304             ( u2_col_out_304    ),
    .col_out_305             ( u2_col_out_305    ),
    .col_out_306             ( u2_col_out_306    ),
    .col_out_307             ( u2_col_out_307    ),
    .col_out_308             ( u2_col_out_308    ),
    .col_out_309             ( u2_col_out_309    ),
    .col_out_310             ( u2_col_out_310    ),
    .col_out_311             ( u2_col_out_311    ),
    .col_out_312             ( u2_col_out_312    ),
    .col_out_313             ( u2_col_out_313    ),
    .col_out_314             ( u2_col_out_314    ),
    .col_out_315             ( u2_col_out_315    ),
    .col_out_316             ( u2_col_out_316    ),
    .col_out_317             ( u2_col_out_317    ),
    .col_out_318             ( u2_col_out_318    ),
    .col_out_319             ( u2_col_out_319    ),
    .col_out_320             ( u2_col_out_320    ),
    .col_out_321             ( u2_col_out_321    ),
    .col_out_322             ( u2_col_out_322    ),
    .col_out_323             ( u2_col_out_323    ),
    .col_out_324             ( u2_col_out_324    ),
    .col_out_325             ( u2_col_out_325    ),
    .col_out_326             ( u2_col_out_326    ),
    .col_out_327             ( u2_col_out_327    ),
    .col_out_328             ( u2_col_out_328    ),
    .col_out_329             ( u2_col_out_329    ),
    .col_out_330             ( u2_col_out_330    ),
    .col_out_331             ( u2_col_out_331    ),
    .col_out_332             ( u2_col_out_332    ),
    .col_out_333             ( u2_col_out_333    ),
    .col_out_334             ( u2_col_out_334    ),
    .col_out_335             ( u2_col_out_335    ),
    .col_out_336             ( u2_col_out_336    ),
    .col_out_337             ( u2_col_out_337    ),
    .col_out_338             ( u2_col_out_338    ),
    .col_out_339             ( u2_col_out_339    ),
    .col_out_340             ( u2_col_out_340    ),
    .col_out_341             ( u2_col_out_341    ),
    .col_out_342             ( u2_col_out_342    ),
    .col_out_343             ( u2_col_out_343    ),
    .col_out_344             ( u2_col_out_344    ),
    .col_out_345             ( u2_col_out_345    ),
    .col_out_346             ( u2_col_out_346    ),
    .col_out_347             ( u2_col_out_347    ),
    .col_out_348             ( u2_col_out_348    ),
    .col_out_349             ( u2_col_out_349    ),
    .col_out_350             ( u2_col_out_350    ),
    .col_out_351             ( u2_col_out_351    ),
    .col_out_352             ( u2_col_out_352    ),
    .col_out_353             ( u2_col_out_353    ),
    .col_out_354             ( u2_col_out_354    ),
    .col_out_355             ( u2_col_out_355    ),
    .col_out_356             ( u2_col_out_356    ),
    .col_out_357             ( u2_col_out_357    ),
    .col_out_358             ( u2_col_out_358    ),
    .col_out_359             ( u2_col_out_359    ),
    .col_out_360             ( u2_col_out_360    ),
    .col_out_361             ( u2_col_out_361    ),
    .col_out_362             ( u2_col_out_362    ),
    .col_out_363             ( u2_col_out_363    ),
    .col_out_364             ( u2_col_out_364    ),
    .col_out_365             ( u2_col_out_365    ),
    .col_out_366             ( u2_col_out_366    ),
    .col_out_367             ( u2_col_out_367    ),
    .col_out_368             ( u2_col_out_368    ),
    .col_out_369             ( u2_col_out_369    ),
    .col_out_370             ( u2_col_out_370    ),
    .col_out_371             ( u2_col_out_371    ),
    .col_out_372             ( u2_col_out_372    ),
    .col_out_373             ( u2_col_out_373    ),
    .col_out_374             ( u2_col_out_374    ),
    .col_out_375             ( u2_col_out_375    ),
    .col_out_376             ( u2_col_out_376    ),
    .col_out_377             ( u2_col_out_377    ),
    .col_out_378             ( u2_col_out_378    ),
    .col_out_379             ( u2_col_out_379    ),
    .col_out_380             ( u2_col_out_380    ),
    .col_out_381             ( u2_col_out_381    ),
    .col_out_382             ( u2_col_out_382    ),
    .col_out_383             ( u2_col_out_383    ),
    .col_out_384             ( u2_col_out_384    ),
    .col_out_385             ( u2_col_out_385    ),
    .col_out_386             ( u2_col_out_386    ),
    .col_out_387             ( u2_col_out_387    ),
    .col_out_388             ( u2_col_out_388    ),
    .col_out_389             ( u2_col_out_389    ),
    .col_out_390             ( u2_col_out_390    ),
    .col_out_391             ( u2_col_out_391    ),
    .col_out_392             ( u2_col_out_392    ),
    .col_out_393             ( u2_col_out_393    ),
    .col_out_394             ( u2_col_out_394    ),
    .col_out_395             ( u2_col_out_395    ),
    .col_out_396             ( u2_col_out_396    ),
    .col_out_397             ( u2_col_out_397    ),
    .col_out_398             ( u2_col_out_398    ),
    .col_out_399             ( u2_col_out_399    ),
    .col_out_400             ( u2_col_out_400    ),
    .col_out_401             ( u2_col_out_401    ),
    .col_out_402             ( u2_col_out_402    ),
    .col_out_403             ( u2_col_out_403    ),
    .col_out_404             ( u2_col_out_404    ),
    .col_out_405             ( u2_col_out_405    ),
    .col_out_406             ( u2_col_out_406    ),
    .col_out_407             ( u2_col_out_407    ),
    .col_out_408             ( u2_col_out_408    ),
    .col_out_409             ( u2_col_out_409    ),
    .col_out_410             ( u2_col_out_410    ),
    .col_out_411             ( u2_col_out_411    ),
    .col_out_412             ( u2_col_out_412    ),
    .col_out_413             ( u2_col_out_413    ),
    .col_out_414             ( u2_col_out_414    ),
    .col_out_415             ( u2_col_out_415    ),
    .col_out_416             ( u2_col_out_416    ),
    .col_out_417             ( u2_col_out_417    ),
    .col_out_418             ( u2_col_out_418    ),
    .col_out_419             ( u2_col_out_419    ),
    .col_out_420             ( u2_col_out_420    ),
    .col_out_421             ( u2_col_out_421    ),
    .col_out_422             ( u2_col_out_422    ),
    .col_out_423             ( u2_col_out_423    ),
    .col_out_424             ( u2_col_out_424    ),
    .col_out_425             ( u2_col_out_425    ),
    .col_out_426             ( u2_col_out_426    ),
    .col_out_427             ( u2_col_out_427    ),
    .col_out_428             ( u2_col_out_428    ),
    .col_out_429             ( u2_col_out_429    ),
    .col_out_430             ( u2_col_out_430    ),
    .col_out_431             ( u2_col_out_431    ),
    .col_out_432             ( u2_col_out_432    ),
    .col_out_433             ( u2_col_out_433    ),
    .col_out_434             ( u2_col_out_434    ),
    .col_out_435             ( u2_col_out_435    ),
    .col_out_436             ( u2_col_out_436    ),
    .col_out_437             ( u2_col_out_437    ),
    .col_out_438             ( u2_col_out_438    ),
    .col_out_439             ( u2_col_out_439    ),
    .col_out_440             ( u2_col_out_440    ),
    .col_out_441             ( u2_col_out_441    ),
    .col_out_442             ( u2_col_out_442    ),
    .col_out_443             ( u2_col_out_443    ),
    .col_out_444             ( u2_col_out_444    ),
    .col_out_445             ( u2_col_out_445    ),
    .col_out_446             ( u2_col_out_446    ),
    .col_out_447             ( u2_col_out_447    ),
    .col_out_448             ( u2_col_out_448    ),
    .col_out_449             ( u2_col_out_449    ),
    .col_out_450             ( u2_col_out_450    ),
    .col_out_451             ( u2_col_out_451    ),
    .col_out_452             ( u2_col_out_452    ),
    .col_out_453             ( u2_col_out_453    ),
    .col_out_454             ( u2_col_out_454    ),
    .col_out_455             ( u2_col_out_455    ),
    .col_out_456             ( u2_col_out_456    ),
    .col_out_457             ( u2_col_out_457    ),
    .col_out_458             ( u2_col_out_458    ),
    .col_out_459             ( u2_col_out_459    ),
    .col_out_460             ( u2_col_out_460    ),
    .col_out_461             ( u2_col_out_461    ),
    .col_out_462             ( u2_col_out_462    ),
    .col_out_463             ( u2_col_out_463    ),
    .col_out_464             ( u2_col_out_464    ),
    .col_out_465             ( u2_col_out_465    ),
    .col_out_466             ( u2_col_out_466    ),
    .col_out_467             ( u2_col_out_467    ),
    .col_out_468             ( u2_col_out_468    ),
    .col_out_469             ( u2_col_out_469    ),
    .col_out_470             ( u2_col_out_470    ),
    .col_out_471             ( u2_col_out_471    ),
    .col_out_472             ( u2_col_out_472    ),
    .col_out_473             ( u2_col_out_473    ),
    .col_out_474             ( u2_col_out_474    ),
    .col_out_475             ( u2_col_out_475    ),
    .col_out_476             ( u2_col_out_476    ),
    .col_out_477             ( u2_col_out_477    ),
    .col_out_478             ( u2_col_out_478    ),
    .col_out_479             ( u2_col_out_479    ),
    .col_out_480             ( u2_col_out_480    ),
    .col_out_481             ( u2_col_out_481    ),
    .col_out_482             ( u2_col_out_482    ),
    .col_out_483             ( u2_col_out_483    ),
    .col_out_484             ( u2_col_out_484    ),
    .col_out_485             ( u2_col_out_485    ),
    .col_out_486             ( u2_col_out_486    ),
    .col_out_487             ( u2_col_out_487    ),
    .col_out_488             ( u2_col_out_488    ),
    .col_out_489             ( u2_col_out_489    ),
    .col_out_490             ( u2_col_out_490    ),
    .col_out_491             ( u2_col_out_491    ),
    .col_out_492             ( u2_col_out_492    ),
    .col_out_493             ( u2_col_out_493    ),
    .col_out_494             ( u2_col_out_494    ),
    .col_out_495             ( u2_col_out_495    ),
    .col_out_496             ( u2_col_out_496    ),
    .col_out_497             ( u2_col_out_497    ),
    .col_out_498             ( u2_col_out_498    ),
    .col_out_499             ( u2_col_out_499    ),
    .col_out_500             ( u2_col_out_500    ),
    .col_out_501             ( u2_col_out_501    ),
    .col_out_502             ( u2_col_out_502    ),
    .col_out_503             ( u2_col_out_503    ),
    .col_out_504             ( u2_col_out_504    ),
    .col_out_505             ( u2_col_out_505    ),
    .col_out_506             ( u2_col_out_506    ),
    .col_out_507             ( u2_col_out_507    ),
    .col_out_508             ( u2_col_out_508    ),
    .col_out_509             ( u2_col_out_509    ),
    .col_out_510             ( u2_col_out_510    ),
    .col_out_511             ( u2_col_out_511    ),
    .col_out_512             ( u2_col_out_512    ),
    .col_out_513             ( u2_col_out_513    ),
    .col_out_514             ( u2_col_out_514    ),
    .col_out_515             ( u2_col_out_515    ),
    .col_out_516             ( u2_col_out_516    ),
    .col_out_517             ( u2_col_out_517    ),
    .col_out_518             ( u2_col_out_518    ),
    .col_out_519             ( u2_col_out_519    ),
    .col_out_520             ( u2_col_out_520    ),
    .col_out_521             ( u2_col_out_521    ),
    .col_out_522             ( u2_col_out_522    ),
    .col_out_523             ( u2_col_out_523    ),
    .col_out_524             ( u2_col_out_524    ),
    .col_out_525             ( u2_col_out_525    ),
    .col_out_526             ( u2_col_out_526    ),
    .col_out_527             ( u2_col_out_527    ),
    .col_out_528             ( u2_col_out_528    ),
    .col_out_529             ( u2_col_out_529    ),
    .col_out_530             ( u2_col_out_530    ),
    .col_out_531             ( u2_col_out_531    ),
    .col_out_532             ( u2_col_out_532    ),
    .col_out_533             ( u2_col_out_533    ),
    .col_out_534             ( u2_col_out_534    ),
    .col_out_535             ( u2_col_out_535    ),
    .col_out_536             ( u2_col_out_536    ),
    .col_out_537             ( u2_col_out_537    ),
    .col_out_538             ( u2_col_out_538    ),
    .col_out_539             ( u2_col_out_539    ),
    .col_out_540             ( u2_col_out_540    ),
    .col_out_541             ( u2_col_out_541    ),
    .col_out_542             ( u2_col_out_542    ),
    .col_out_543             ( u2_col_out_543    ),
    .col_out_544             ( u2_col_out_544    ),
    .col_out_545             ( u2_col_out_545    ),
    .col_out_546             ( u2_col_out_546    ),
    .col_out_547             ( u2_col_out_547    ),
    .col_out_548             ( u2_col_out_548    ),
    .col_out_549             ( u2_col_out_549    ),
    .col_out_550             ( u2_col_out_550    ),
    .col_out_551             ( u2_col_out_551    ),
    .col_out_552             ( u2_col_out_552    ),
    .col_out_553             ( u2_col_out_553    ),
    .col_out_554             ( u2_col_out_554    ),
    .col_out_555             ( u2_col_out_555    ),
    .col_out_556             ( u2_col_out_556    ),
    .col_out_557             ( u2_col_out_557    ),
    .col_out_558             ( u2_col_out_558    ),
    .col_out_559             ( u2_col_out_559    ),
    .col_out_560             ( u2_col_out_560    ),
    .col_out_561             ( u2_col_out_561    ),
    .col_out_562             ( u2_col_out_562    ),
    .col_out_563             ( u2_col_out_563    ),
    .col_out_564             ( u2_col_out_564    ),
    .col_out_565             ( u2_col_out_565    ),
    .col_out_566             ( u2_col_out_566    ),
    .col_out_567             ( u2_col_out_567    ),
    .col_out_568             ( u2_col_out_568    ),
    .col_out_569             ( u2_col_out_569    ),
    .col_out_570             ( u2_col_out_570    ),
    .col_out_571             ( u2_col_out_571    ),
    .col_out_572             ( u2_col_out_572    ),
    .col_out_573             ( u2_col_out_573    ),
    .col_out_574             ( u2_col_out_574    ),
    .col_out_575             ( u2_col_out_575    ),
    .col_out_576             ( u2_col_out_576    ),
    .col_out_577             ( u2_col_out_577    ),
    .col_out_578             ( u2_col_out_578    ),
    .col_out_579             ( u2_col_out_579    ),
    .col_out_580             ( u2_col_out_580    ),
    .col_out_581             ( u2_col_out_581    ),
    .col_out_582             ( u2_col_out_582    ),
    .col_out_583             ( u2_col_out_583    ),
    .col_out_584             ( u2_col_out_584    ),
    .col_out_585             ( u2_col_out_585    ),
    .col_out_586             ( u2_col_out_586    ),
    .col_out_587             ( u2_col_out_587    ),
    .col_out_588             ( u2_col_out_588    ),
    .col_out_589             ( u2_col_out_589    ),
    .col_out_590             ( u2_col_out_590    ),
    .col_out_591             ( u2_col_out_591    ),
    .col_out_592             ( u2_col_out_592    ),
    .col_out_593             ( u2_col_out_593    ),
    .col_out_594             ( u2_col_out_594    ),
    .col_out_595             ( u2_col_out_595    ),
    .col_out_596             ( u2_col_out_596    ),
    .col_out_597             ( u2_col_out_597    ),
    .col_out_598             ( u2_col_out_598    ),
    .col_out_599             ( u2_col_out_599    ),
    .col_out_600             ( u2_col_out_600    ),
    .col_out_601             ( u2_col_out_601    ),
    .col_out_602             ( u2_col_out_602    ),
    .col_out_603             ( u2_col_out_603    ),
    .col_out_604             ( u2_col_out_604    ),
    .col_out_605             ( u2_col_out_605    ),
    .col_out_606             ( u2_col_out_606    ),
    .col_out_607             ( u2_col_out_607    ),
    .col_out_608             ( u2_col_out_608    ),
    .col_out_609             ( u2_col_out_609    ),
    .col_out_610             ( u2_col_out_610    ),
    .col_out_611             ( u2_col_out_611    ),
    .col_out_612             ( u2_col_out_612    ),
    .col_out_613             ( u2_col_out_613    ),
    .col_out_614             ( u2_col_out_614    ),
    .col_out_615             ( u2_col_out_615    ),
    .col_out_616             ( u2_col_out_616    ),
    .col_out_617             ( u2_col_out_617    ),
    .col_out_618             ( u2_col_out_618    ),
    .col_out_619             ( u2_col_out_619    ),
    .col_out_620             ( u2_col_out_620    ),
    .col_out_621             ( u2_col_out_621    ),
    .col_out_622             ( u2_col_out_622    ),
    .col_out_623             ( u2_col_out_623    ),
    .col_out_624             ( u2_col_out_624    ),
    .col_out_625             ( u2_col_out_625    ),
    .col_out_626             ( u2_col_out_626    ),
    .col_out_627             ( u2_col_out_627    ),
    .col_out_628             ( u2_col_out_628    ),
    .col_out_629             ( u2_col_out_629    ),
    .col_out_630             ( u2_col_out_630    ),
    .col_out_631             ( u2_col_out_631    ),
    .col_out_632             ( u2_col_out_632    ),
    .col_out_633             ( u2_col_out_633    ),
    .col_out_634             ( u2_col_out_634    ),
    .col_out_635             ( u2_col_out_635    ),
    .col_out_636             ( u2_col_out_636    ),
    .col_out_637             ( u2_col_out_637    ),
    .col_out_638             ( u2_col_out_638    ),
    .col_out_639             ( u2_col_out_639    ),
    .col_out_640             ( u2_col_out_640    ),
    .col_out_641             ( u2_col_out_641    ),
    .col_out_642             ( u2_col_out_642    ),
    .col_out_643             ( u2_col_out_643    ),
    .col_out_644             ( u2_col_out_644    ),
    .col_out_645             ( u2_col_out_645    ),
    .col_out_646             ( u2_col_out_646    ),
    .col_out_647             ( u2_col_out_647    ),
    .col_out_648             ( u2_col_out_648    ),
    .col_out_649             ( u2_col_out_649    ),
    .col_out_650             ( u2_col_out_650    ),
    .col_out_651             ( u2_col_out_651    ),
    .col_out_652             ( u2_col_out_652    ),
    .col_out_653             ( u2_col_out_653    ),
    .col_out_654             ( u2_col_out_654    ),
    .col_out_655             ( u2_col_out_655    ),
    .col_out_656             ( u2_col_out_656    ),
    .col_out_657             ( u2_col_out_657    ),
    .col_out_658             ( u2_col_out_658    ),
    .col_out_659             ( u2_col_out_659    ),
    .col_out_660             ( u2_col_out_660    ),
    .col_out_661             ( u2_col_out_661    ),
    .col_out_662             ( u2_col_out_662    ),
    .col_out_663             ( u2_col_out_663    ),
    .col_out_664             ( u2_col_out_664    ),
    .col_out_665             ( u2_col_out_665    ),
    .col_out_666             ( u2_col_out_666    ),
    .col_out_667             ( u2_col_out_667    ),
    .col_out_668             ( u2_col_out_668    ),
    .col_out_669             ( u2_col_out_669    ),
    .col_out_670             ( u2_col_out_670    ),
    .col_out_671             ( u2_col_out_671    ),
    .col_out_672             ( u2_col_out_672    ),
    .col_out_673             ( u2_col_out_673    ),
    .col_out_674             ( u2_col_out_674    ),
    .col_out_675             ( u2_col_out_675    ),
    .col_out_676             ( u2_col_out_676    ),
    .col_out_677             ( u2_col_out_677    ),
    .col_out_678             ( u2_col_out_678    ),
    .col_out_679             ( u2_col_out_679    ),
    .col_out_680             ( u2_col_out_680    ),
    .col_out_681             ( u2_col_out_681    ),
    .col_out_682             ( u2_col_out_682    ),
    .col_out_683             ( u2_col_out_683    ),
    .col_out_684             ( u2_col_out_684    ),
    .col_out_685             ( u2_col_out_685    ),
    .col_out_686             ( u2_col_out_686    ),
    .col_out_687             ( u2_col_out_687    ),
    .col_out_688             ( u2_col_out_688    ),
    .col_out_689             ( u2_col_out_689    ),
    .col_out_690             ( u2_col_out_690    ),
    .col_out_691             ( u2_col_out_691    ),
    .col_out_692             ( u2_col_out_692    ),
    .col_out_693             ( u2_col_out_693    ),
    .col_out_694             ( u2_col_out_694    ),
    .col_out_695             ( u2_col_out_695    ),
    .col_out_696             ( u2_col_out_696    ),
    .col_out_697             ( u2_col_out_697    ),
    .col_out_698             ( u2_col_out_698    ),
    .col_out_699             ( u2_col_out_699    ),
    .col_out_700             ( u2_col_out_700    ),
    .col_out_701             ( u2_col_out_701    ),
    .col_out_702             ( u2_col_out_702    ),
    .col_out_703             ( u2_col_out_703    ),
    .col_out_704             ( u2_col_out_704    ),
    .col_out_705             ( u2_col_out_705    ),
    .col_out_706             ( u2_col_out_706    ),
    .col_out_707             ( u2_col_out_707    ),
    .col_out_708             ( u2_col_out_708    ),
    .col_out_709             ( u2_col_out_709    ),
    .col_out_710             ( u2_col_out_710    ),
    .col_out_711             ( u2_col_out_711    ),
    .col_out_712             ( u2_col_out_712    ),
    .col_out_713             ( u2_col_out_713    ),
    .col_out_714             ( u2_col_out_714    ),
    .col_out_715             ( u2_col_out_715    ),
    .col_out_716             ( u2_col_out_716    ),
    .col_out_717             ( u2_col_out_717    ),
    .col_out_718             ( u2_col_out_718    ),
    .col_out_719             ( u2_col_out_719    ),
    .col_out_720             ( u2_col_out_720    ),
    .col_out_721             ( u2_col_out_721    ),
    .col_out_722             ( u2_col_out_722    ),
    .col_out_723             ( u2_col_out_723    ),
    .col_out_724             ( u2_col_out_724    ),
    .col_out_725             ( u2_col_out_725    ),
    .col_out_726             ( u2_col_out_726    ),
    .col_out_727             ( u2_col_out_727    ),
    .col_out_728             ( u2_col_out_728    ),
    .col_out_729             ( u2_col_out_729    ),
    .col_out_730             ( u2_col_out_730    ),
    .col_out_731             ( u2_col_out_731    ),
    .col_out_732             ( u2_col_out_732    ),
    .col_out_733             ( u2_col_out_733    ),
    .col_out_734             ( u2_col_out_734    ),
    .col_out_735             ( u2_col_out_735    ),
    .col_out_736             ( u2_col_out_736    ),
    .col_out_737             ( u2_col_out_737    ),
    .col_out_738             ( u2_col_out_738    ),
    .col_out_739             ( u2_col_out_739    ),
    .col_out_740             ( u2_col_out_740    ),
    .col_out_741             ( u2_col_out_741    ),
    .col_out_742             ( u2_col_out_742    ),
    .col_out_743             ( u2_col_out_743    ),
    .col_out_744             ( u2_col_out_744    ),
    .col_out_745             ( u2_col_out_745    ),
    .col_out_746             ( u2_col_out_746    ),
    .col_out_747             ( u2_col_out_747    ),
    .col_out_748             ( u2_col_out_748    ),
    .col_out_749             ( u2_col_out_749    ),
    .col_out_750             ( u2_col_out_750    ),
    .col_out_751             ( u2_col_out_751    ),
    .col_out_752             ( u2_col_out_752    ),
    .col_out_753             ( u2_col_out_753    ),
    .col_out_754             ( u2_col_out_754    ),
    .col_out_755             ( u2_col_out_755    ),
    .col_out_756             ( u2_col_out_756    ),
    .col_out_757             ( u2_col_out_757    ),
    .col_out_758             ( u2_col_out_758    ),
    .col_out_759             ( u2_col_out_759    ),
    .col_out_760             ( u2_col_out_760    ),
    .col_out_761             ( u2_col_out_761    ),
    .col_out_762             ( u2_col_out_762    ),
    .col_out_763             ( u2_col_out_763    ),
    .col_out_764             ( u2_col_out_764    ),
    .col_out_765             ( u2_col_out_765    ),
    .col_out_766             ( u2_col_out_766    ),
    .col_out_767             ( u2_col_out_767    ),
    .col_out_768             ( u2_col_out_768    ),
    .col_out_769             ( u2_col_out_769    ),
    .col_out_770             ( u2_col_out_770    ),
    .col_out_771             ( u2_col_out_771    ),
    .col_out_772             ( u2_col_out_772    ),
    .col_out_773             ( u2_col_out_773    ),
    .col_out_774             ( u2_col_out_774    ),
    .col_out_775             ( u2_col_out_775    ),
    .col_out_776             ( u2_col_out_776    ),
    .col_out_777             ( u2_col_out_777    ),
    .col_out_778             ( u2_col_out_778    ),
    .col_out_779             ( u2_col_out_779    ),
    .col_out_780             ( u2_col_out_780    ),
    .col_out_781             ( u2_col_out_781    ),
    .col_out_782             ( u2_col_out_782    ),
    .col_out_783             ( u2_col_out_783    ),
    .col_out_784             ( u2_col_out_784    ),
    .col_out_785             ( u2_col_out_785    ),
    .col_out_786             ( u2_col_out_786    ),
    .col_out_787             ( u2_col_out_787    ),
    .col_out_788             ( u2_col_out_788    ),
    .col_out_789             ( u2_col_out_789    ),
    .col_out_790             ( u2_col_out_790    ),
    .col_out_791             ( u2_col_out_791    ),
    .col_out_792             ( u2_col_out_792    ),
    .col_out_793             ( u2_col_out_793    ),
    .col_out_794             ( u2_col_out_794    ),
    .col_out_795             ( u2_col_out_795    ),
    .col_out_796             ( u2_col_out_796    ),
    .col_out_797             ( u2_col_out_797    ),
    .col_out_798             ( u2_col_out_798    ),
    .col_out_799             ( u2_col_out_799    ),
    .col_out_800             ( u2_col_out_800    ),
    .col_out_801             ( u2_col_out_801    ),
    .col_out_802             ( u2_col_out_802    ),
    .col_out_803             ( u2_col_out_803    ),
    .col_out_804             ( u2_col_out_804    ),
    .col_out_805             ( u2_col_out_805    ),
    .col_out_806             ( u2_col_out_806    ),
    .col_out_807             ( u2_col_out_807    ),
    .col_out_808             ( u2_col_out_808    ),
    .col_out_809             ( u2_col_out_809    ),
    .col_out_810             ( u2_col_out_810    ),
    .col_out_811             ( u2_col_out_811    ),
    .col_out_812             ( u2_col_out_812    ),
    .col_out_813             ( u2_col_out_813    ),
    .col_out_814             ( u2_col_out_814    ),
    .col_out_815             ( u2_col_out_815    ),
    .col_out_816             ( u2_col_out_816    ),
    .col_out_817             ( u2_col_out_817    ),
    .col_out_818             ( u2_col_out_818    ),
    .col_out_819             ( u2_col_out_819    ),
    .col_out_820             ( u2_col_out_820    ),
    .col_out_821             ( u2_col_out_821    ),
    .col_out_822             ( u2_col_out_822    ),
    .col_out_823             ( u2_col_out_823    ),
    .col_out_824             ( u2_col_out_824    ),
    .col_out_825             ( u2_col_out_825    ),
    .col_out_826             ( u2_col_out_826    ),
    .col_out_827             ( u2_col_out_827    ),
    .col_out_828             ( u2_col_out_828    ),
    .col_out_829             ( u2_col_out_829    ),
    .col_out_830             ( u2_col_out_830    ),
    .col_out_831             ( u2_col_out_831    ),
    .col_out_832             ( u2_col_out_832    ),
    .col_out_833             ( u2_col_out_833    ),
    .col_out_834             ( u2_col_out_834    ),
    .col_out_835             ( u2_col_out_835    ),
    .col_out_836             ( u2_col_out_836    ),
    .col_out_837             ( u2_col_out_837    ),
    .col_out_838             ( u2_col_out_838    ),
    .col_out_839             ( u2_col_out_839    ),
    .col_out_840             ( u2_col_out_840    ),
    .col_out_841             ( u2_col_out_841    ),
    .col_out_842             ( u2_col_out_842    ),
    .col_out_843             ( u2_col_out_843    ),
    .col_out_844             ( u2_col_out_844    ),
    .col_out_845             ( u2_col_out_845    ),
    .col_out_846             ( u2_col_out_846    ),
    .col_out_847             ( u2_col_out_847    ),
    .col_out_848             ( u2_col_out_848    ),
    .col_out_849             ( u2_col_out_849    ),
    .col_out_850             ( u2_col_out_850    ),
    .col_out_851             ( u2_col_out_851    ),
    .col_out_852             ( u2_col_out_852    ),
    .col_out_853             ( u2_col_out_853    ),
    .col_out_854             ( u2_col_out_854    ),
    .col_out_855             ( u2_col_out_855    ),
    .col_out_856             ( u2_col_out_856    ),
    .col_out_857             ( u2_col_out_857    ),
    .col_out_858             ( u2_col_out_858    ),
    .col_out_859             ( u2_col_out_859    ),
    .col_out_860             ( u2_col_out_860    ),
    .col_out_861             ( u2_col_out_861    ),
    .col_out_862             ( u2_col_out_862    ),
    .col_out_863             ( u2_col_out_863    ),
    .col_out_864             ( u2_col_out_864    ),
    .col_out_865             ( u2_col_out_865    ),
    .col_out_866             ( u2_col_out_866    ),
    .col_out_867             ( u2_col_out_867    ),
    .col_out_868             ( u2_col_out_868    ),
    .col_out_869             ( u2_col_out_869    ),
    .col_out_870             ( u2_col_out_870    ),
    .col_out_871             ( u2_col_out_871    ),
    .col_out_872             ( u2_col_out_872    ),
    .col_out_873             ( u2_col_out_873    ),
    .col_out_874             ( u2_col_out_874    ),
    .col_out_875             ( u2_col_out_875    ),
    .col_out_876             ( u2_col_out_876    ),
    .col_out_877             ( u2_col_out_877    ),
    .col_out_878             ( u2_col_out_878    ),
    .col_out_879             ( u2_col_out_879    ),
    .col_out_880             ( u2_col_out_880    ),
    .col_out_881             ( u2_col_out_881    ),
    .col_out_882             ( u2_col_out_882    ),
    .col_out_883             ( u2_col_out_883    ),
    .col_out_884             ( u2_col_out_884    ),
    .col_out_885             ( u2_col_out_885    ),
    .col_out_886             ( u2_col_out_886    ),
    .col_out_887             ( u2_col_out_887    ),
    .col_out_888             ( u2_col_out_888    ),
    .col_out_889             ( u2_col_out_889    ),
    .col_out_890             ( u2_col_out_890    ),
    .col_out_891             ( u2_col_out_891    ),
    .col_out_892             ( u2_col_out_892    ),
    .col_out_893             ( u2_col_out_893    ),
    .col_out_894             ( u2_col_out_894    ),
    .col_out_895             ( u2_col_out_895    ),
    .col_out_896             ( u2_col_out_896    ),
    .col_out_897             ( u2_col_out_897    ),
    .col_out_898             ( u2_col_out_898    ),
    .col_out_899             ( u2_col_out_899    ),
    .col_out_900             ( u2_col_out_900    ),
    .col_out_901             ( u2_col_out_901    ),
    .col_out_902             ( u2_col_out_902    ),
    .col_out_903             ( u2_col_out_903    ),
    .col_out_904             ( u2_col_out_904    ),
    .col_out_905             ( u2_col_out_905    ),
    .col_out_906             ( u2_col_out_906    ),
    .col_out_907             ( u2_col_out_907    ),
    .col_out_908             ( u2_col_out_908    ),
    .col_out_909             ( u2_col_out_909    ),
    .col_out_910             ( u2_col_out_910    ),
    .col_out_911             ( u2_col_out_911    ),
    .col_out_912             ( u2_col_out_912    ),
    .col_out_913             ( u2_col_out_913    ),
    .col_out_914             ( u2_col_out_914    ),
    .col_out_915             ( u2_col_out_915    ),
    .col_out_916             ( u2_col_out_916    ),
    .col_out_917             ( u2_col_out_917    ),
    .col_out_918             ( u2_col_out_918    ),
    .col_out_919             ( u2_col_out_919    ),
    .col_out_920             ( u2_col_out_920    ),
    .col_out_921             ( u2_col_out_921    ),
    .col_out_922             ( u2_col_out_922    ),
    .col_out_923             ( u2_col_out_923    ),
    .col_out_924             ( u2_col_out_924    ),
    .col_out_925             ( u2_col_out_925    ),
    .col_out_926             ( u2_col_out_926    ),
    .col_out_927             ( u2_col_out_927    ),
    .col_out_928             ( u2_col_out_928    ),
    .col_out_929             ( u2_col_out_929    ),
    .col_out_930             ( u2_col_out_930    ),
    .col_out_931             ( u2_col_out_931    ),
    .col_out_932             ( u2_col_out_932    ),
    .col_out_933             ( u2_col_out_933    ),
    .col_out_934             ( u2_col_out_934    ),
    .col_out_935             ( u2_col_out_935    ),
    .col_out_936             ( u2_col_out_936    ),
    .col_out_937             ( u2_col_out_937    ),
    .col_out_938             ( u2_col_out_938    ),
    .col_out_939             ( u2_col_out_939    ),
    .col_out_940             ( u2_col_out_940    ),
    .col_out_941             ( u2_col_out_941    ),
    .col_out_942             ( u2_col_out_942    ),
    .col_out_943             ( u2_col_out_943    ),
    .col_out_944             ( u2_col_out_944    ),
    .col_out_945             ( u2_col_out_945    ),
    .col_out_946             ( u2_col_out_946    ),
    .col_out_947             ( u2_col_out_947    ),
    .col_out_948             ( u2_col_out_948    ),
    .col_out_949             ( u2_col_out_949    ),
    .col_out_950             ( u2_col_out_950    ),
    .col_out_951             ( u2_col_out_951    ),
    .col_out_952             ( u2_col_out_952    ),
    .col_out_953             ( u2_col_out_953    ),
    .col_out_954             ( u2_col_out_954    ),
    .col_out_955             ( u2_col_out_955    ),
    .col_out_956             ( u2_col_out_956    ),
    .col_out_957             ( u2_col_out_957    ),
    .col_out_958             ( u2_col_out_958    ),
    .col_out_959             ( u2_col_out_959    ),
    .col_out_960             ( u2_col_out_960    ),
    .col_out_961             ( u2_col_out_961    ),
    .col_out_962             ( u2_col_out_962    ),
    .col_out_963             ( u2_col_out_963    ),
    .col_out_964             ( u2_col_out_964    ),
    .col_out_965             ( u2_col_out_965    ),
    .col_out_966             ( u2_col_out_966    ),
    .col_out_967             ( u2_col_out_967    ),
    .col_out_968             ( u2_col_out_968    ),
    .col_out_969             ( u2_col_out_969    ),
    .col_out_970             ( u2_col_out_970    ),
    .col_out_971             ( u2_col_out_971    ),
    .col_out_972             ( u2_col_out_972    ),
    .col_out_973             ( u2_col_out_973    ),
    .col_out_974             ( u2_col_out_974    ),
    .col_out_975             ( u2_col_out_975    ),
    .col_out_976             ( u2_col_out_976    ),
    .col_out_977             ( u2_col_out_977    ),
    .col_out_978             ( u2_col_out_978    ),
    .col_out_979             ( u2_col_out_979    ),
    .col_out_980             ( u2_col_out_980    ),
    .col_out_981             ( u2_col_out_981    ),
    .col_out_982             ( u2_col_out_982    ),
    .col_out_983             ( u2_col_out_983    ),
    .col_out_984             ( u2_col_out_984    ),
    .col_out_985             ( u2_col_out_985    ),
    .col_out_986             ( u2_col_out_986    ),
    .col_out_987             ( u2_col_out_987    ),
    .col_out_988             ( u2_col_out_988    ),
    .col_out_989             ( u2_col_out_989    ),
    .col_out_990             ( u2_col_out_990    ),
    .col_out_991             ( u2_col_out_991    ),
    .col_out_992             ( u2_col_out_992    ),
    .col_out_993             ( u2_col_out_993    ),
    .col_out_994             ( u2_col_out_994    ),
    .col_out_995             ( u2_col_out_995    ),
    .col_out_996             ( u2_col_out_996    ),
    .col_out_997             ( u2_col_out_997    ),
    .col_out_998             ( u2_col_out_998    ),
    .col_out_999             ( u2_col_out_999    ),
    .col_out_1000            ( u2_col_out_1000   ),
    .col_out_1001            ( u2_col_out_1001   ),
    .col_out_1002            ( u2_col_out_1002   ),
    .col_out_1003            ( u2_col_out_1003   ),
    .col_out_1004            ( u2_col_out_1004   ),
    .col_out_1005            ( u2_col_out_1005   ),
    .col_out_1006            ( u2_col_out_1006   ),
    .col_out_1007            ( u2_col_out_1007   ),
    .col_out_1008            ( u2_col_out_1008   ),
    .col_out_1009            ( u2_col_out_1009   ),
    .col_out_1010            ( u2_col_out_1010   ),
    .col_out_1011            ( u2_col_out_1011   ),
    .col_out_1012            ( u2_col_out_1012   ),
    .col_out_1013            ( u2_col_out_1013   ),
    .col_out_1014            ( u2_col_out_1014   ),
    .col_out_1015            ( u2_col_out_1015   ),
    .col_out_1016            ( u2_col_out_1016   ),
    .col_out_1017            ( u2_col_out_1017   ),
    .col_out_1018            ( u2_col_out_1018   ),
    .col_out_1019            ( u2_col_out_1019   ),
    .col_out_1020            ( u2_col_out_1020   ),
    .col_out_1021            ( u2_col_out_1021   ),
    .col_out_1022            ( u2_col_out_1022   ),
    .col_out_1023            ( u2_col_out_1023   ),
    .col_out_1024            ( u2_col_out_1024   ),
    .col_out_1025            ( u2_col_out_1025   ),
    .col_out_1026            ( u2_col_out_1026   ),
    .col_out_1027            ( u2_col_out_1027   ),
    .col_out_1028            ( u2_col_out_1028   ),
    .col_out_1029            ( u2_col_out_1029   ),
    .col_out_1030            ( u2_col_out_1030   ),
    .col_out_1031            ( u2_col_out_1031   ),
    .col_out_1032            ( u2_col_out_1032   ),
    .col_out_1033            ( u2_col_out_1033   )
);

































// compressor_array_6_4_1033 Outputs
wire  [3:0]  u3_col_out_0;
wire  [3:0]  u3_col_out_1;
wire  [3:0]  u3_col_out_2;
wire  [3:0]  u3_col_out_3;
wire  [3:0]  u3_col_out_4;
wire  [3:0]  u3_col_out_5;
wire  [3:0]  u3_col_out_6;
wire  [3:0]  u3_col_out_7;
wire  [3:0]  u3_col_out_8;
wire  [3:0]  u3_col_out_9;
wire  [3:0]  u3_col_out_10;
wire  [3:0]  u3_col_out_11;
wire  [3:0]  u3_col_out_12;
wire  [3:0]  u3_col_out_13;
wire  [3:0]  u3_col_out_14;
wire  [3:0]  u3_col_out_15;
wire  [3:0]  u3_col_out_16;
wire  [3:0]  u3_col_out_17;
wire  [3:0]  u3_col_out_18;
wire  [3:0]  u3_col_out_19;
wire  [3:0]  u3_col_out_20;
wire  [3:0]  u3_col_out_21;
wire  [3:0]  u3_col_out_22;
wire  [3:0]  u3_col_out_23;
wire  [3:0]  u3_col_out_24;
wire  [3:0]  u3_col_out_25;
wire  [3:0]  u3_col_out_26;
wire  [3:0]  u3_col_out_27;
wire  [3:0]  u3_col_out_28;
wire  [3:0]  u3_col_out_29;
wire  [3:0]  u3_col_out_30;
wire  [3:0]  u3_col_out_31;
wire  [3:0]  u3_col_out_32;
wire  [3:0]  u3_col_out_33;
wire  [3:0]  u3_col_out_34;
wire  [3:0]  u3_col_out_35;
wire  [3:0]  u3_col_out_36;
wire  [3:0]  u3_col_out_37;
wire  [3:0]  u3_col_out_38;
wire  [3:0]  u3_col_out_39;
wire  [3:0]  u3_col_out_40;
wire  [3:0]  u3_col_out_41;
wire  [3:0]  u3_col_out_42;
wire  [3:0]  u3_col_out_43;
wire  [3:0]  u3_col_out_44;
wire  [3:0]  u3_col_out_45;
wire  [3:0]  u3_col_out_46;
wire  [3:0]  u3_col_out_47;
wire  [3:0]  u3_col_out_48;
wire  [3:0]  u3_col_out_49;
wire  [3:0]  u3_col_out_50;
wire  [3:0]  u3_col_out_51;
wire  [3:0]  u3_col_out_52;
wire  [3:0]  u3_col_out_53;
wire  [3:0]  u3_col_out_54;
wire  [3:0]  u3_col_out_55;
wire  [3:0]  u3_col_out_56;
wire  [3:0]  u3_col_out_57;
wire  [3:0]  u3_col_out_58;
wire  [3:0]  u3_col_out_59;
wire  [3:0]  u3_col_out_60;
wire  [3:0]  u3_col_out_61;
wire  [3:0]  u3_col_out_62;
wire  [3:0]  u3_col_out_63;
wire  [3:0]  u3_col_out_64;
wire  [3:0]  u3_col_out_65;
wire  [3:0]  u3_col_out_66;
wire  [3:0]  u3_col_out_67;
wire  [3:0]  u3_col_out_68;
wire  [3:0]  u3_col_out_69;
wire  [3:0]  u3_col_out_70;
wire  [3:0]  u3_col_out_71;
wire  [3:0]  u3_col_out_72;
wire  [3:0]  u3_col_out_73;
wire  [3:0]  u3_col_out_74;
wire  [3:0]  u3_col_out_75;
wire  [3:0]  u3_col_out_76;
wire  [3:0]  u3_col_out_77;
wire  [3:0]  u3_col_out_78;
wire  [3:0]  u3_col_out_79;
wire  [3:0]  u3_col_out_80;
wire  [3:0]  u3_col_out_81;
wire  [3:0]  u3_col_out_82;
wire  [3:0]  u3_col_out_83;
wire  [3:0]  u3_col_out_84;
wire  [3:0]  u3_col_out_85;
wire  [3:0]  u3_col_out_86;
wire  [3:0]  u3_col_out_87;
wire  [3:0]  u3_col_out_88;
wire  [3:0]  u3_col_out_89;
wire  [3:0]  u3_col_out_90;
wire  [3:0]  u3_col_out_91;
wire  [3:0]  u3_col_out_92;
wire  [3:0]  u3_col_out_93;
wire  [3:0]  u3_col_out_94;
wire  [3:0]  u3_col_out_95;
wire  [3:0]  u3_col_out_96;
wire  [3:0]  u3_col_out_97;
wire  [3:0]  u3_col_out_98;
wire  [3:0]  u3_col_out_99;
wire  [3:0]  u3_col_out_100;
wire  [3:0]  u3_col_out_101;
wire  [3:0]  u3_col_out_102;
wire  [3:0]  u3_col_out_103;
wire  [3:0]  u3_col_out_104;
wire  [3:0]  u3_col_out_105;
wire  [3:0]  u3_col_out_106;
wire  [3:0]  u3_col_out_107;
wire  [3:0]  u3_col_out_108;
wire  [3:0]  u3_col_out_109;
wire  [3:0]  u3_col_out_110;
wire  [3:0]  u3_col_out_111;
wire  [3:0]  u3_col_out_112;
wire  [3:0]  u3_col_out_113;
wire  [3:0]  u3_col_out_114;
wire  [3:0]  u3_col_out_115;
wire  [3:0]  u3_col_out_116;
wire  [3:0]  u3_col_out_117;
wire  [3:0]  u3_col_out_118;
wire  [3:0]  u3_col_out_119;
wire  [3:0]  u3_col_out_120;
wire  [3:0]  u3_col_out_121;
wire  [3:0]  u3_col_out_122;
wire  [3:0]  u3_col_out_123;
wire  [3:0]  u3_col_out_124;
wire  [3:0]  u3_col_out_125;
wire  [3:0]  u3_col_out_126;
wire  [3:0]  u3_col_out_127;
wire  [3:0]  u3_col_out_128;
wire  [3:0]  u3_col_out_129;
wire  [3:0]  u3_col_out_130;
wire  [3:0]  u3_col_out_131;
wire  [3:0]  u3_col_out_132;
wire  [3:0]  u3_col_out_133;
wire  [3:0]  u3_col_out_134;
wire  [3:0]  u3_col_out_135;
wire  [3:0]  u3_col_out_136;
wire  [3:0]  u3_col_out_137;
wire  [3:0]  u3_col_out_138;
wire  [3:0]  u3_col_out_139;
wire  [3:0]  u3_col_out_140;
wire  [3:0]  u3_col_out_141;
wire  [3:0]  u3_col_out_142;
wire  [3:0]  u3_col_out_143;
wire  [3:0]  u3_col_out_144;
wire  [3:0]  u3_col_out_145;
wire  [3:0]  u3_col_out_146;
wire  [3:0]  u3_col_out_147;
wire  [3:0]  u3_col_out_148;
wire  [3:0]  u3_col_out_149;
wire  [3:0]  u3_col_out_150;
wire  [3:0]  u3_col_out_151;
wire  [3:0]  u3_col_out_152;
wire  [3:0]  u3_col_out_153;
wire  [3:0]  u3_col_out_154;
wire  [3:0]  u3_col_out_155;
wire  [3:0]  u3_col_out_156;
wire  [3:0]  u3_col_out_157;
wire  [3:0]  u3_col_out_158;
wire  [3:0]  u3_col_out_159;
wire  [3:0]  u3_col_out_160;
wire  [3:0]  u3_col_out_161;
wire  [3:0]  u3_col_out_162;
wire  [3:0]  u3_col_out_163;
wire  [3:0]  u3_col_out_164;
wire  [3:0]  u3_col_out_165;
wire  [3:0]  u3_col_out_166;
wire  [3:0]  u3_col_out_167;
wire  [3:0]  u3_col_out_168;
wire  [3:0]  u3_col_out_169;
wire  [3:0]  u3_col_out_170;
wire  [3:0]  u3_col_out_171;
wire  [3:0]  u3_col_out_172;
wire  [3:0]  u3_col_out_173;
wire  [3:0]  u3_col_out_174;
wire  [3:0]  u3_col_out_175;
wire  [3:0]  u3_col_out_176;
wire  [3:0]  u3_col_out_177;
wire  [3:0]  u3_col_out_178;
wire  [3:0]  u3_col_out_179;
wire  [3:0]  u3_col_out_180;
wire  [3:0]  u3_col_out_181;
wire  [3:0]  u3_col_out_182;
wire  [3:0]  u3_col_out_183;
wire  [3:0]  u3_col_out_184;
wire  [3:0]  u3_col_out_185;
wire  [3:0]  u3_col_out_186;
wire  [3:0]  u3_col_out_187;
wire  [3:0]  u3_col_out_188;
wire  [3:0]  u3_col_out_189;
wire  [3:0]  u3_col_out_190;
wire  [3:0]  u3_col_out_191;
wire  [3:0]  u3_col_out_192;
wire  [3:0]  u3_col_out_193;
wire  [3:0]  u3_col_out_194;
wire  [3:0]  u3_col_out_195;
wire  [3:0]  u3_col_out_196;
wire  [3:0]  u3_col_out_197;
wire  [3:0]  u3_col_out_198;
wire  [3:0]  u3_col_out_199;
wire  [3:0]  u3_col_out_200;
wire  [3:0]  u3_col_out_201;
wire  [3:0]  u3_col_out_202;
wire  [3:0]  u3_col_out_203;
wire  [3:0]  u3_col_out_204;
wire  [3:0]  u3_col_out_205;
wire  [3:0]  u3_col_out_206;
wire  [3:0]  u3_col_out_207;
wire  [3:0]  u3_col_out_208;
wire  [3:0]  u3_col_out_209;
wire  [3:0]  u3_col_out_210;
wire  [3:0]  u3_col_out_211;
wire  [3:0]  u3_col_out_212;
wire  [3:0]  u3_col_out_213;
wire  [3:0]  u3_col_out_214;
wire  [3:0]  u3_col_out_215;
wire  [3:0]  u3_col_out_216;
wire  [3:0]  u3_col_out_217;
wire  [3:0]  u3_col_out_218;
wire  [3:0]  u3_col_out_219;
wire  [3:0]  u3_col_out_220;
wire  [3:0]  u3_col_out_221;
wire  [3:0]  u3_col_out_222;
wire  [3:0]  u3_col_out_223;
wire  [3:0]  u3_col_out_224;
wire  [3:0]  u3_col_out_225;
wire  [3:0]  u3_col_out_226;
wire  [3:0]  u3_col_out_227;
wire  [3:0]  u3_col_out_228;
wire  [3:0]  u3_col_out_229;
wire  [3:0]  u3_col_out_230;
wire  [3:0]  u3_col_out_231;
wire  [3:0]  u3_col_out_232;
wire  [3:0]  u3_col_out_233;
wire  [3:0]  u3_col_out_234;
wire  [3:0]  u3_col_out_235;
wire  [3:0]  u3_col_out_236;
wire  [3:0]  u3_col_out_237;
wire  [3:0]  u3_col_out_238;
wire  [3:0]  u3_col_out_239;
wire  [3:0]  u3_col_out_240;
wire  [3:0]  u3_col_out_241;
wire  [3:0]  u3_col_out_242;
wire  [3:0]  u3_col_out_243;
wire  [3:0]  u3_col_out_244;
wire  [3:0]  u3_col_out_245;
wire  [3:0]  u3_col_out_246;
wire  [3:0]  u3_col_out_247;
wire  [3:0]  u3_col_out_248;
wire  [3:0]  u3_col_out_249;
wire  [3:0]  u3_col_out_250;
wire  [3:0]  u3_col_out_251;
wire  [3:0]  u3_col_out_252;
wire  [3:0]  u3_col_out_253;
wire  [3:0]  u3_col_out_254;
wire  [3:0]  u3_col_out_255;
wire  [3:0]  u3_col_out_256;
wire  [3:0]  u3_col_out_257;
wire  [3:0]  u3_col_out_258;
wire  [3:0]  u3_col_out_259;
wire  [3:0]  u3_col_out_260;
wire  [3:0]  u3_col_out_261;
wire  [3:0]  u3_col_out_262;
wire  [3:0]  u3_col_out_263;
wire  [3:0]  u3_col_out_264;
wire  [3:0]  u3_col_out_265;
wire  [3:0]  u3_col_out_266;
wire  [3:0]  u3_col_out_267;
wire  [3:0]  u3_col_out_268;
wire  [3:0]  u3_col_out_269;
wire  [3:0]  u3_col_out_270;
wire  [3:0]  u3_col_out_271;
wire  [3:0]  u3_col_out_272;
wire  [3:0]  u3_col_out_273;
wire  [3:0]  u3_col_out_274;
wire  [3:0]  u3_col_out_275;
wire  [3:0]  u3_col_out_276;
wire  [3:0]  u3_col_out_277;
wire  [3:0]  u3_col_out_278;
wire  [3:0]  u3_col_out_279;
wire  [3:0]  u3_col_out_280;
wire  [3:0]  u3_col_out_281;
wire  [3:0]  u3_col_out_282;
wire  [3:0]  u3_col_out_283;
wire  [3:0]  u3_col_out_284;
wire  [3:0]  u3_col_out_285;
wire  [3:0]  u3_col_out_286;
wire  [3:0]  u3_col_out_287;
wire  [3:0]  u3_col_out_288;
wire  [3:0]  u3_col_out_289;
wire  [3:0]  u3_col_out_290;
wire  [3:0]  u3_col_out_291;
wire  [3:0]  u3_col_out_292;
wire  [3:0]  u3_col_out_293;
wire  [3:0]  u3_col_out_294;
wire  [3:0]  u3_col_out_295;
wire  [3:0]  u3_col_out_296;
wire  [3:0]  u3_col_out_297;
wire  [3:0]  u3_col_out_298;
wire  [3:0]  u3_col_out_299;
wire  [3:0]  u3_col_out_300;
wire  [3:0]  u3_col_out_301;
wire  [3:0]  u3_col_out_302;
wire  [3:0]  u3_col_out_303;
wire  [3:0]  u3_col_out_304;
wire  [3:0]  u3_col_out_305;
wire  [3:0]  u3_col_out_306;
wire  [3:0]  u3_col_out_307;
wire  [3:0]  u3_col_out_308;
wire  [3:0]  u3_col_out_309;
wire  [3:0]  u3_col_out_310;
wire  [3:0]  u3_col_out_311;
wire  [3:0]  u3_col_out_312;
wire  [3:0]  u3_col_out_313;
wire  [3:0]  u3_col_out_314;
wire  [3:0]  u3_col_out_315;
wire  [3:0]  u3_col_out_316;
wire  [3:0]  u3_col_out_317;
wire  [3:0]  u3_col_out_318;
wire  [3:0]  u3_col_out_319;
wire  [3:0]  u3_col_out_320;
wire  [3:0]  u3_col_out_321;
wire  [3:0]  u3_col_out_322;
wire  [3:0]  u3_col_out_323;
wire  [3:0]  u3_col_out_324;
wire  [3:0]  u3_col_out_325;
wire  [3:0]  u3_col_out_326;
wire  [3:0]  u3_col_out_327;
wire  [3:0]  u3_col_out_328;
wire  [3:0]  u3_col_out_329;
wire  [3:0]  u3_col_out_330;
wire  [3:0]  u3_col_out_331;
wire  [3:0]  u3_col_out_332;
wire  [3:0]  u3_col_out_333;
wire  [3:0]  u3_col_out_334;
wire  [3:0]  u3_col_out_335;
wire  [3:0]  u3_col_out_336;
wire  [3:0]  u3_col_out_337;
wire  [3:0]  u3_col_out_338;
wire  [3:0]  u3_col_out_339;
wire  [3:0]  u3_col_out_340;
wire  [3:0]  u3_col_out_341;
wire  [3:0]  u3_col_out_342;
wire  [3:0]  u3_col_out_343;
wire  [3:0]  u3_col_out_344;
wire  [3:0]  u3_col_out_345;
wire  [3:0]  u3_col_out_346;
wire  [3:0]  u3_col_out_347;
wire  [3:0]  u3_col_out_348;
wire  [3:0]  u3_col_out_349;
wire  [3:0]  u3_col_out_350;
wire  [3:0]  u3_col_out_351;
wire  [3:0]  u3_col_out_352;
wire  [3:0]  u3_col_out_353;
wire  [3:0]  u3_col_out_354;
wire  [3:0]  u3_col_out_355;
wire  [3:0]  u3_col_out_356;
wire  [3:0]  u3_col_out_357;
wire  [3:0]  u3_col_out_358;
wire  [3:0]  u3_col_out_359;
wire  [3:0]  u3_col_out_360;
wire  [3:0]  u3_col_out_361;
wire  [3:0]  u3_col_out_362;
wire  [3:0]  u3_col_out_363;
wire  [3:0]  u3_col_out_364;
wire  [3:0]  u3_col_out_365;
wire  [3:0]  u3_col_out_366;
wire  [3:0]  u3_col_out_367;
wire  [3:0]  u3_col_out_368;
wire  [3:0]  u3_col_out_369;
wire  [3:0]  u3_col_out_370;
wire  [3:0]  u3_col_out_371;
wire  [3:0]  u3_col_out_372;
wire  [3:0]  u3_col_out_373;
wire  [3:0]  u3_col_out_374;
wire  [3:0]  u3_col_out_375;
wire  [3:0]  u3_col_out_376;
wire  [3:0]  u3_col_out_377;
wire  [3:0]  u3_col_out_378;
wire  [3:0]  u3_col_out_379;
wire  [3:0]  u3_col_out_380;
wire  [3:0]  u3_col_out_381;
wire  [3:0]  u3_col_out_382;
wire  [3:0]  u3_col_out_383;
wire  [3:0]  u3_col_out_384;
wire  [3:0]  u3_col_out_385;
wire  [3:0]  u3_col_out_386;
wire  [3:0]  u3_col_out_387;
wire  [3:0]  u3_col_out_388;
wire  [3:0]  u3_col_out_389;
wire  [3:0]  u3_col_out_390;
wire  [3:0]  u3_col_out_391;
wire  [3:0]  u3_col_out_392;
wire  [3:0]  u3_col_out_393;
wire  [3:0]  u3_col_out_394;
wire  [3:0]  u3_col_out_395;
wire  [3:0]  u3_col_out_396;
wire  [3:0]  u3_col_out_397;
wire  [3:0]  u3_col_out_398;
wire  [3:0]  u3_col_out_399;
wire  [3:0]  u3_col_out_400;
wire  [3:0]  u3_col_out_401;
wire  [3:0]  u3_col_out_402;
wire  [3:0]  u3_col_out_403;
wire  [3:0]  u3_col_out_404;
wire  [3:0]  u3_col_out_405;
wire  [3:0]  u3_col_out_406;
wire  [3:0]  u3_col_out_407;
wire  [3:0]  u3_col_out_408;
wire  [3:0]  u3_col_out_409;
wire  [3:0]  u3_col_out_410;
wire  [3:0]  u3_col_out_411;
wire  [3:0]  u3_col_out_412;
wire  [3:0]  u3_col_out_413;
wire  [3:0]  u3_col_out_414;
wire  [3:0]  u3_col_out_415;
wire  [3:0]  u3_col_out_416;
wire  [3:0]  u3_col_out_417;
wire  [3:0]  u3_col_out_418;
wire  [3:0]  u3_col_out_419;
wire  [3:0]  u3_col_out_420;
wire  [3:0]  u3_col_out_421;
wire  [3:0]  u3_col_out_422;
wire  [3:0]  u3_col_out_423;
wire  [3:0]  u3_col_out_424;
wire  [3:0]  u3_col_out_425;
wire  [3:0]  u3_col_out_426;
wire  [3:0]  u3_col_out_427;
wire  [3:0]  u3_col_out_428;
wire  [3:0]  u3_col_out_429;
wire  [3:0]  u3_col_out_430;
wire  [3:0]  u3_col_out_431;
wire  [3:0]  u3_col_out_432;
wire  [3:0]  u3_col_out_433;
wire  [3:0]  u3_col_out_434;
wire  [3:0]  u3_col_out_435;
wire  [3:0]  u3_col_out_436;
wire  [3:0]  u3_col_out_437;
wire  [3:0]  u3_col_out_438;
wire  [3:0]  u3_col_out_439;
wire  [3:0]  u3_col_out_440;
wire  [3:0]  u3_col_out_441;
wire  [3:0]  u3_col_out_442;
wire  [3:0]  u3_col_out_443;
wire  [3:0]  u3_col_out_444;
wire  [3:0]  u3_col_out_445;
wire  [3:0]  u3_col_out_446;
wire  [3:0]  u3_col_out_447;
wire  [3:0]  u3_col_out_448;
wire  [3:0]  u3_col_out_449;
wire  [3:0]  u3_col_out_450;
wire  [3:0]  u3_col_out_451;
wire  [3:0]  u3_col_out_452;
wire  [3:0]  u3_col_out_453;
wire  [3:0]  u3_col_out_454;
wire  [3:0]  u3_col_out_455;
wire  [3:0]  u3_col_out_456;
wire  [3:0]  u3_col_out_457;
wire  [3:0]  u3_col_out_458;
wire  [3:0]  u3_col_out_459;
wire  [3:0]  u3_col_out_460;
wire  [3:0]  u3_col_out_461;
wire  [3:0]  u3_col_out_462;
wire  [3:0]  u3_col_out_463;
wire  [3:0]  u3_col_out_464;
wire  [3:0]  u3_col_out_465;
wire  [3:0]  u3_col_out_466;
wire  [3:0]  u3_col_out_467;
wire  [3:0]  u3_col_out_468;
wire  [3:0]  u3_col_out_469;
wire  [3:0]  u3_col_out_470;
wire  [3:0]  u3_col_out_471;
wire  [3:0]  u3_col_out_472;
wire  [3:0]  u3_col_out_473;
wire  [3:0]  u3_col_out_474;
wire  [3:0]  u3_col_out_475;
wire  [3:0]  u3_col_out_476;
wire  [3:0]  u3_col_out_477;
wire  [3:0]  u3_col_out_478;
wire  [3:0]  u3_col_out_479;
wire  [3:0]  u3_col_out_480;
wire  [3:0]  u3_col_out_481;
wire  [3:0]  u3_col_out_482;
wire  [3:0]  u3_col_out_483;
wire  [3:0]  u3_col_out_484;
wire  [3:0]  u3_col_out_485;
wire  [3:0]  u3_col_out_486;
wire  [3:0]  u3_col_out_487;
wire  [3:0]  u3_col_out_488;
wire  [3:0]  u3_col_out_489;
wire  [3:0]  u3_col_out_490;
wire  [3:0]  u3_col_out_491;
wire  [3:0]  u3_col_out_492;
wire  [3:0]  u3_col_out_493;
wire  [3:0]  u3_col_out_494;
wire  [3:0]  u3_col_out_495;
wire  [3:0]  u3_col_out_496;
wire  [3:0]  u3_col_out_497;
wire  [3:0]  u3_col_out_498;
wire  [3:0]  u3_col_out_499;
wire  [3:0]  u3_col_out_500;
wire  [3:0]  u3_col_out_501;
wire  [3:0]  u3_col_out_502;
wire  [3:0]  u3_col_out_503;
wire  [3:0]  u3_col_out_504;
wire  [3:0]  u3_col_out_505;
wire  [3:0]  u3_col_out_506;
wire  [3:0]  u3_col_out_507;
wire  [3:0]  u3_col_out_508;
wire  [3:0]  u3_col_out_509;
wire  [3:0]  u3_col_out_510;
wire  [3:0]  u3_col_out_511;
wire  [3:0]  u3_col_out_512;
wire  [3:0]  u3_col_out_513;
wire  [3:0]  u3_col_out_514;
wire  [3:0]  u3_col_out_515;
wire  [3:0]  u3_col_out_516;
wire  [3:0]  u3_col_out_517;
wire  [3:0]  u3_col_out_518;
wire  [3:0]  u3_col_out_519;
wire  [3:0]  u3_col_out_520;
wire  [3:0]  u3_col_out_521;
wire  [3:0]  u3_col_out_522;
wire  [3:0]  u3_col_out_523;
wire  [3:0]  u3_col_out_524;
wire  [3:0]  u3_col_out_525;
wire  [3:0]  u3_col_out_526;
wire  [3:0]  u3_col_out_527;
wire  [3:0]  u3_col_out_528;
wire  [3:0]  u3_col_out_529;
wire  [3:0]  u3_col_out_530;
wire  [3:0]  u3_col_out_531;
wire  [3:0]  u3_col_out_532;
wire  [3:0]  u3_col_out_533;
wire  [3:0]  u3_col_out_534;
wire  [3:0]  u3_col_out_535;
wire  [3:0]  u3_col_out_536;
wire  [3:0]  u3_col_out_537;
wire  [3:0]  u3_col_out_538;
wire  [3:0]  u3_col_out_539;
wire  [3:0]  u3_col_out_540;
wire  [3:0]  u3_col_out_541;
wire  [3:0]  u3_col_out_542;
wire  [3:0]  u3_col_out_543;
wire  [3:0]  u3_col_out_544;
wire  [3:0]  u3_col_out_545;
wire  [3:0]  u3_col_out_546;
wire  [3:0]  u3_col_out_547;
wire  [3:0]  u3_col_out_548;
wire  [3:0]  u3_col_out_549;
wire  [3:0]  u3_col_out_550;
wire  [3:0]  u3_col_out_551;
wire  [3:0]  u3_col_out_552;
wire  [3:0]  u3_col_out_553;
wire  [3:0]  u3_col_out_554;
wire  [3:0]  u3_col_out_555;
wire  [3:0]  u3_col_out_556;
wire  [3:0]  u3_col_out_557;
wire  [3:0]  u3_col_out_558;
wire  [3:0]  u3_col_out_559;
wire  [3:0]  u3_col_out_560;
wire  [3:0]  u3_col_out_561;
wire  [3:0]  u3_col_out_562;
wire  [3:0]  u3_col_out_563;
wire  [3:0]  u3_col_out_564;
wire  [3:0]  u3_col_out_565;
wire  [3:0]  u3_col_out_566;
wire  [3:0]  u3_col_out_567;
wire  [3:0]  u3_col_out_568;
wire  [3:0]  u3_col_out_569;
wire  [3:0]  u3_col_out_570;
wire  [3:0]  u3_col_out_571;
wire  [3:0]  u3_col_out_572;
wire  [3:0]  u3_col_out_573;
wire  [3:0]  u3_col_out_574;
wire  [3:0]  u3_col_out_575;
wire  [3:0]  u3_col_out_576;
wire  [3:0]  u3_col_out_577;
wire  [3:0]  u3_col_out_578;
wire  [3:0]  u3_col_out_579;
wire  [3:0]  u3_col_out_580;
wire  [3:0]  u3_col_out_581;
wire  [3:0]  u3_col_out_582;
wire  [3:0]  u3_col_out_583;
wire  [3:0]  u3_col_out_584;
wire  [3:0]  u3_col_out_585;
wire  [3:0]  u3_col_out_586;
wire  [3:0]  u3_col_out_587;
wire  [3:0]  u3_col_out_588;
wire  [3:0]  u3_col_out_589;
wire  [3:0]  u3_col_out_590;
wire  [3:0]  u3_col_out_591;
wire  [3:0]  u3_col_out_592;
wire  [3:0]  u3_col_out_593;
wire  [3:0]  u3_col_out_594;
wire  [3:0]  u3_col_out_595;
wire  [3:0]  u3_col_out_596;
wire  [3:0]  u3_col_out_597;
wire  [3:0]  u3_col_out_598;
wire  [3:0]  u3_col_out_599;
wire  [3:0]  u3_col_out_600;
wire  [3:0]  u3_col_out_601;
wire  [3:0]  u3_col_out_602;
wire  [3:0]  u3_col_out_603;
wire  [3:0]  u3_col_out_604;
wire  [3:0]  u3_col_out_605;
wire  [3:0]  u3_col_out_606;
wire  [3:0]  u3_col_out_607;
wire  [3:0]  u3_col_out_608;
wire  [3:0]  u3_col_out_609;
wire  [3:0]  u3_col_out_610;
wire  [3:0]  u3_col_out_611;
wire  [3:0]  u3_col_out_612;
wire  [3:0]  u3_col_out_613;
wire  [3:0]  u3_col_out_614;
wire  [3:0]  u3_col_out_615;
wire  [3:0]  u3_col_out_616;
wire  [3:0]  u3_col_out_617;
wire  [3:0]  u3_col_out_618;
wire  [3:0]  u3_col_out_619;
wire  [3:0]  u3_col_out_620;
wire  [3:0]  u3_col_out_621;
wire  [3:0]  u3_col_out_622;
wire  [3:0]  u3_col_out_623;
wire  [3:0]  u3_col_out_624;
wire  [3:0]  u3_col_out_625;
wire  [3:0]  u3_col_out_626;
wire  [3:0]  u3_col_out_627;
wire  [3:0]  u3_col_out_628;
wire  [3:0]  u3_col_out_629;
wire  [3:0]  u3_col_out_630;
wire  [3:0]  u3_col_out_631;
wire  [3:0]  u3_col_out_632;
wire  [3:0]  u3_col_out_633;
wire  [3:0]  u3_col_out_634;
wire  [3:0]  u3_col_out_635;
wire  [3:0]  u3_col_out_636;
wire  [3:0]  u3_col_out_637;
wire  [3:0]  u3_col_out_638;
wire  [3:0]  u3_col_out_639;
wire  [3:0]  u3_col_out_640;
wire  [3:0]  u3_col_out_641;
wire  [3:0]  u3_col_out_642;
wire  [3:0]  u3_col_out_643;
wire  [3:0]  u3_col_out_644;
wire  [3:0]  u3_col_out_645;
wire  [3:0]  u3_col_out_646;
wire  [3:0]  u3_col_out_647;
wire  [3:0]  u3_col_out_648;
wire  [3:0]  u3_col_out_649;
wire  [3:0]  u3_col_out_650;
wire  [3:0]  u3_col_out_651;
wire  [3:0]  u3_col_out_652;
wire  [3:0]  u3_col_out_653;
wire  [3:0]  u3_col_out_654;
wire  [3:0]  u3_col_out_655;
wire  [3:0]  u3_col_out_656;
wire  [3:0]  u3_col_out_657;
wire  [3:0]  u3_col_out_658;
wire  [3:0]  u3_col_out_659;
wire  [3:0]  u3_col_out_660;
wire  [3:0]  u3_col_out_661;
wire  [3:0]  u3_col_out_662;
wire  [3:0]  u3_col_out_663;
wire  [3:0]  u3_col_out_664;
wire  [3:0]  u3_col_out_665;
wire  [3:0]  u3_col_out_666;
wire  [3:0]  u3_col_out_667;
wire  [3:0]  u3_col_out_668;
wire  [3:0]  u3_col_out_669;
wire  [3:0]  u3_col_out_670;
wire  [3:0]  u3_col_out_671;
wire  [3:0]  u3_col_out_672;
wire  [3:0]  u3_col_out_673;
wire  [3:0]  u3_col_out_674;
wire  [3:0]  u3_col_out_675;
wire  [3:0]  u3_col_out_676;
wire  [3:0]  u3_col_out_677;
wire  [3:0]  u3_col_out_678;
wire  [3:0]  u3_col_out_679;
wire  [3:0]  u3_col_out_680;
wire  [3:0]  u3_col_out_681;
wire  [3:0]  u3_col_out_682;
wire  [3:0]  u3_col_out_683;
wire  [3:0]  u3_col_out_684;
wire  [3:0]  u3_col_out_685;
wire  [3:0]  u3_col_out_686;
wire  [3:0]  u3_col_out_687;
wire  [3:0]  u3_col_out_688;
wire  [3:0]  u3_col_out_689;
wire  [3:0]  u3_col_out_690;
wire  [3:0]  u3_col_out_691;
wire  [3:0]  u3_col_out_692;
wire  [3:0]  u3_col_out_693;
wire  [3:0]  u3_col_out_694;
wire  [3:0]  u3_col_out_695;
wire  [3:0]  u3_col_out_696;
wire  [3:0]  u3_col_out_697;
wire  [3:0]  u3_col_out_698;
wire  [3:0]  u3_col_out_699;
wire  [3:0]  u3_col_out_700;
wire  [3:0]  u3_col_out_701;
wire  [3:0]  u3_col_out_702;
wire  [3:0]  u3_col_out_703;
wire  [3:0]  u3_col_out_704;
wire  [3:0]  u3_col_out_705;
wire  [3:0]  u3_col_out_706;
wire  [3:0]  u3_col_out_707;
wire  [3:0]  u3_col_out_708;
wire  [3:0]  u3_col_out_709;
wire  [3:0]  u3_col_out_710;
wire  [3:0]  u3_col_out_711;
wire  [3:0]  u3_col_out_712;
wire  [3:0]  u3_col_out_713;
wire  [3:0]  u3_col_out_714;
wire  [3:0]  u3_col_out_715;
wire  [3:0]  u3_col_out_716;
wire  [3:0]  u3_col_out_717;
wire  [3:0]  u3_col_out_718;
wire  [3:0]  u3_col_out_719;
wire  [3:0]  u3_col_out_720;
wire  [3:0]  u3_col_out_721;
wire  [3:0]  u3_col_out_722;
wire  [3:0]  u3_col_out_723;
wire  [3:0]  u3_col_out_724;
wire  [3:0]  u3_col_out_725;
wire  [3:0]  u3_col_out_726;
wire  [3:0]  u3_col_out_727;
wire  [3:0]  u3_col_out_728;
wire  [3:0]  u3_col_out_729;
wire  [3:0]  u3_col_out_730;
wire  [3:0]  u3_col_out_731;
wire  [3:0]  u3_col_out_732;
wire  [3:0]  u3_col_out_733;
wire  [3:0]  u3_col_out_734;
wire  [3:0]  u3_col_out_735;
wire  [3:0]  u3_col_out_736;
wire  [3:0]  u3_col_out_737;
wire  [3:0]  u3_col_out_738;
wire  [3:0]  u3_col_out_739;
wire  [3:0]  u3_col_out_740;
wire  [3:0]  u3_col_out_741;
wire  [3:0]  u3_col_out_742;
wire  [3:0]  u3_col_out_743;
wire  [3:0]  u3_col_out_744;
wire  [3:0]  u3_col_out_745;
wire  [3:0]  u3_col_out_746;
wire  [3:0]  u3_col_out_747;
wire  [3:0]  u3_col_out_748;
wire  [3:0]  u3_col_out_749;
wire  [3:0]  u3_col_out_750;
wire  [3:0]  u3_col_out_751;
wire  [3:0]  u3_col_out_752;
wire  [3:0]  u3_col_out_753;
wire  [3:0]  u3_col_out_754;
wire  [3:0]  u3_col_out_755;
wire  [3:0]  u3_col_out_756;
wire  [3:0]  u3_col_out_757;
wire  [3:0]  u3_col_out_758;
wire  [3:0]  u3_col_out_759;
wire  [3:0]  u3_col_out_760;
wire  [3:0]  u3_col_out_761;
wire  [3:0]  u3_col_out_762;
wire  [3:0]  u3_col_out_763;
wire  [3:0]  u3_col_out_764;
wire  [3:0]  u3_col_out_765;
wire  [3:0]  u3_col_out_766;
wire  [3:0]  u3_col_out_767;
wire  [3:0]  u3_col_out_768;
wire  [3:0]  u3_col_out_769;
wire  [3:0]  u3_col_out_770;
wire  [3:0]  u3_col_out_771;
wire  [3:0]  u3_col_out_772;
wire  [3:0]  u3_col_out_773;
wire  [3:0]  u3_col_out_774;
wire  [3:0]  u3_col_out_775;
wire  [3:0]  u3_col_out_776;
wire  [3:0]  u3_col_out_777;
wire  [3:0]  u3_col_out_778;
wire  [3:0]  u3_col_out_779;
wire  [3:0]  u3_col_out_780;
wire  [3:0]  u3_col_out_781;
wire  [3:0]  u3_col_out_782;
wire  [3:0]  u3_col_out_783;
wire  [3:0]  u3_col_out_784;
wire  [3:0]  u3_col_out_785;
wire  [3:0]  u3_col_out_786;
wire  [3:0]  u3_col_out_787;
wire  [3:0]  u3_col_out_788;
wire  [3:0]  u3_col_out_789;
wire  [3:0]  u3_col_out_790;
wire  [3:0]  u3_col_out_791;
wire  [3:0]  u3_col_out_792;
wire  [3:0]  u3_col_out_793;
wire  [3:0]  u3_col_out_794;
wire  [3:0]  u3_col_out_795;
wire  [3:0]  u3_col_out_796;
wire  [3:0]  u3_col_out_797;
wire  [3:0]  u3_col_out_798;
wire  [3:0]  u3_col_out_799;
wire  [3:0]  u3_col_out_800;
wire  [3:0]  u3_col_out_801;
wire  [3:0]  u3_col_out_802;
wire  [3:0]  u3_col_out_803;
wire  [3:0]  u3_col_out_804;
wire  [3:0]  u3_col_out_805;
wire  [3:0]  u3_col_out_806;
wire  [3:0]  u3_col_out_807;
wire  [3:0]  u3_col_out_808;
wire  [3:0]  u3_col_out_809;
wire  [3:0]  u3_col_out_810;
wire  [3:0]  u3_col_out_811;
wire  [3:0]  u3_col_out_812;
wire  [3:0]  u3_col_out_813;
wire  [3:0]  u3_col_out_814;
wire  [3:0]  u3_col_out_815;
wire  [3:0]  u3_col_out_816;
wire  [3:0]  u3_col_out_817;
wire  [3:0]  u3_col_out_818;
wire  [3:0]  u3_col_out_819;
wire  [3:0]  u3_col_out_820;
wire  [3:0]  u3_col_out_821;
wire  [3:0]  u3_col_out_822;
wire  [3:0]  u3_col_out_823;
wire  [3:0]  u3_col_out_824;
wire  [3:0]  u3_col_out_825;
wire  [3:0]  u3_col_out_826;
wire  [3:0]  u3_col_out_827;
wire  [3:0]  u3_col_out_828;
wire  [3:0]  u3_col_out_829;
wire  [3:0]  u3_col_out_830;
wire  [3:0]  u3_col_out_831;
wire  [3:0]  u3_col_out_832;
wire  [3:0]  u3_col_out_833;
wire  [3:0]  u3_col_out_834;
wire  [3:0]  u3_col_out_835;
wire  [3:0]  u3_col_out_836;
wire  [3:0]  u3_col_out_837;
wire  [3:0]  u3_col_out_838;
wire  [3:0]  u3_col_out_839;
wire  [3:0]  u3_col_out_840;
wire  [3:0]  u3_col_out_841;
wire  [3:0]  u3_col_out_842;
wire  [3:0]  u3_col_out_843;
wire  [3:0]  u3_col_out_844;
wire  [3:0]  u3_col_out_845;
wire  [3:0]  u3_col_out_846;
wire  [3:0]  u3_col_out_847;
wire  [3:0]  u3_col_out_848;
wire  [3:0]  u3_col_out_849;
wire  [3:0]  u3_col_out_850;
wire  [3:0]  u3_col_out_851;
wire  [3:0]  u3_col_out_852;
wire  [3:0]  u3_col_out_853;
wire  [3:0]  u3_col_out_854;
wire  [3:0]  u3_col_out_855;
wire  [3:0]  u3_col_out_856;
wire  [3:0]  u3_col_out_857;
wire  [3:0]  u3_col_out_858;
wire  [3:0]  u3_col_out_859;
wire  [3:0]  u3_col_out_860;
wire  [3:0]  u3_col_out_861;
wire  [3:0]  u3_col_out_862;
wire  [3:0]  u3_col_out_863;
wire  [3:0]  u3_col_out_864;
wire  [3:0]  u3_col_out_865;
wire  [3:0]  u3_col_out_866;
wire  [3:0]  u3_col_out_867;
wire  [3:0]  u3_col_out_868;
wire  [3:0]  u3_col_out_869;
wire  [3:0]  u3_col_out_870;
wire  [3:0]  u3_col_out_871;
wire  [3:0]  u3_col_out_872;
wire  [3:0]  u3_col_out_873;
wire  [3:0]  u3_col_out_874;
wire  [3:0]  u3_col_out_875;
wire  [3:0]  u3_col_out_876;
wire  [3:0]  u3_col_out_877;
wire  [3:0]  u3_col_out_878;
wire  [3:0]  u3_col_out_879;
wire  [3:0]  u3_col_out_880;
wire  [3:0]  u3_col_out_881;
wire  [3:0]  u3_col_out_882;
wire  [3:0]  u3_col_out_883;
wire  [3:0]  u3_col_out_884;
wire  [3:0]  u3_col_out_885;
wire  [3:0]  u3_col_out_886;
wire  [3:0]  u3_col_out_887;
wire  [3:0]  u3_col_out_888;
wire  [3:0]  u3_col_out_889;
wire  [3:0]  u3_col_out_890;
wire  [3:0]  u3_col_out_891;
wire  [3:0]  u3_col_out_892;
wire  [3:0]  u3_col_out_893;
wire  [3:0]  u3_col_out_894;
wire  [3:0]  u3_col_out_895;
wire  [3:0]  u3_col_out_896;
wire  [3:0]  u3_col_out_897;
wire  [3:0]  u3_col_out_898;
wire  [3:0]  u3_col_out_899;
wire  [3:0]  u3_col_out_900;
wire  [3:0]  u3_col_out_901;
wire  [3:0]  u3_col_out_902;
wire  [3:0]  u3_col_out_903;
wire  [3:0]  u3_col_out_904;
wire  [3:0]  u3_col_out_905;
wire  [3:0]  u3_col_out_906;
wire  [3:0]  u3_col_out_907;
wire  [3:0]  u3_col_out_908;
wire  [3:0]  u3_col_out_909;
wire  [3:0]  u3_col_out_910;
wire  [3:0]  u3_col_out_911;
wire  [3:0]  u3_col_out_912;
wire  [3:0]  u3_col_out_913;
wire  [3:0]  u3_col_out_914;
wire  [3:0]  u3_col_out_915;
wire  [3:0]  u3_col_out_916;
wire  [3:0]  u3_col_out_917;
wire  [3:0]  u3_col_out_918;
wire  [3:0]  u3_col_out_919;
wire  [3:0]  u3_col_out_920;
wire  [3:0]  u3_col_out_921;
wire  [3:0]  u3_col_out_922;
wire  [3:0]  u3_col_out_923;
wire  [3:0]  u3_col_out_924;
wire  [3:0]  u3_col_out_925;
wire  [3:0]  u3_col_out_926;
wire  [3:0]  u3_col_out_927;
wire  [3:0]  u3_col_out_928;
wire  [3:0]  u3_col_out_929;
wire  [3:0]  u3_col_out_930;
wire  [3:0]  u3_col_out_931;
wire  [3:0]  u3_col_out_932;
wire  [3:0]  u3_col_out_933;
wire  [3:0]  u3_col_out_934;
wire  [3:0]  u3_col_out_935;
wire  [3:0]  u3_col_out_936;
wire  [3:0]  u3_col_out_937;
wire  [3:0]  u3_col_out_938;
wire  [3:0]  u3_col_out_939;
wire  [3:0]  u3_col_out_940;
wire  [3:0]  u3_col_out_941;
wire  [3:0]  u3_col_out_942;
wire  [3:0]  u3_col_out_943;
wire  [3:0]  u3_col_out_944;
wire  [3:0]  u3_col_out_945;
wire  [3:0]  u3_col_out_946;
wire  [3:0]  u3_col_out_947;
wire  [3:0]  u3_col_out_948;
wire  [3:0]  u3_col_out_949;
wire  [3:0]  u3_col_out_950;
wire  [3:0]  u3_col_out_951;
wire  [3:0]  u3_col_out_952;
wire  [3:0]  u3_col_out_953;
wire  [3:0]  u3_col_out_954;
wire  [3:0]  u3_col_out_955;
wire  [3:0]  u3_col_out_956;
wire  [3:0]  u3_col_out_957;
wire  [3:0]  u3_col_out_958;
wire  [3:0]  u3_col_out_959;
wire  [3:0]  u3_col_out_960;
wire  [3:0]  u3_col_out_961;
wire  [3:0]  u3_col_out_962;
wire  [3:0]  u3_col_out_963;
wire  [3:0]  u3_col_out_964;
wire  [3:0]  u3_col_out_965;
wire  [3:0]  u3_col_out_966;
wire  [3:0]  u3_col_out_967;
wire  [3:0]  u3_col_out_968;
wire  [3:0]  u3_col_out_969;
wire  [3:0]  u3_col_out_970;
wire  [3:0]  u3_col_out_971;
wire  [3:0]  u3_col_out_972;
wire  [3:0]  u3_col_out_973;
wire  [3:0]  u3_col_out_974;
wire  [3:0]  u3_col_out_975;
wire  [3:0]  u3_col_out_976;
wire  [3:0]  u3_col_out_977;
wire  [3:0]  u3_col_out_978;
wire  [3:0]  u3_col_out_979;
wire  [3:0]  u3_col_out_980;
wire  [3:0]  u3_col_out_981;
wire  [3:0]  u3_col_out_982;
wire  [3:0]  u3_col_out_983;
wire  [3:0]  u3_col_out_984;
wire  [3:0]  u3_col_out_985;
wire  [3:0]  u3_col_out_986;
wire  [3:0]  u3_col_out_987;
wire  [3:0]  u3_col_out_988;
wire  [3:0]  u3_col_out_989;
wire  [3:0]  u3_col_out_990;
wire  [3:0]  u3_col_out_991;
wire  [3:0]  u3_col_out_992;
wire  [3:0]  u3_col_out_993;
wire  [3:0]  u3_col_out_994;
wire  [3:0]  u3_col_out_995;
wire  [3:0]  u3_col_out_996;
wire  [3:0]  u3_col_out_997;
wire  [3:0]  u3_col_out_998;
wire  [3:0]  u3_col_out_999;
wire  [3:0]  u3_col_out_1000;
wire  [3:0]  u3_col_out_1001;
wire  [3:0]  u3_col_out_1002;
wire  [3:0]  u3_col_out_1003;
wire  [3:0]  u3_col_out_1004;
wire  [3:0]  u3_col_out_1005;
wire  [3:0]  u3_col_out_1006;
wire  [3:0]  u3_col_out_1007;
wire  [3:0]  u3_col_out_1008;
wire  [3:0]  u3_col_out_1009;
wire  [3:0]  u3_col_out_1010;
wire  [3:0]  u3_col_out_1011;
wire  [3:0]  u3_col_out_1012;
wire  [3:0]  u3_col_out_1013;
wire  [3:0]  u3_col_out_1014;
wire  [3:0]  u3_col_out_1015;
wire  [3:0]  u3_col_out_1016;
wire  [3:0]  u3_col_out_1017;
wire  [3:0]  u3_col_out_1018;
wire  [3:0]  u3_col_out_1019;
wire  [3:0]  u3_col_out_1020;
wire  [3:0]  u3_col_out_1021;
wire  [3:0]  u3_col_out_1022;
wire  [3:0]  u3_col_out_1023;
wire  [3:0]  u3_col_out_1024;
wire  [3:0]  u3_col_out_1025;
wire  [3:0]  u3_col_out_1026;
wire  [3:0]  u3_col_out_1027;
wire  [3:0]  u3_col_out_1028;
wire  [3:0]  u3_col_out_1029;
wire  [3:0]  u3_col_out_1030;
wire  [3:0]  u3_col_out_1031;
wire  [3:0]  u3_col_out_1032;
wire  [3:0]  u3_col_out_1033;


compressor_array_6_4_1033  u3_compressor_array_6_4_1033 (
    .col_in_0                ( u2_col_out_0       ),
    .col_in_1                ( u2_col_out_1       ),
    .col_in_2                ( u2_col_out_2       ),
    .col_in_3                ( u2_col_out_3       ),
    .col_in_4                ( u2_col_out_4       ),
    .col_in_5                ( u2_col_out_5       ),
    .col_in_6                ( u2_col_out_6       ),
    .col_in_7                ( u2_col_out_7       ),
    .col_in_8                ( u2_col_out_8       ),
    .col_in_9                ( u2_col_out_9       ),
    .col_in_10               ( u2_col_out_10      ),
    .col_in_11               ( u2_col_out_11      ),
    .col_in_12               ( u2_col_out_12      ),
    .col_in_13               ( u2_col_out_13      ),
    .col_in_14               ( u2_col_out_14      ),
    .col_in_15               ( u2_col_out_15      ),
    .col_in_16               ( u2_col_out_16      ),
    .col_in_17               ( u2_col_out_17      ),
    .col_in_18               ( u2_col_out_18      ),
    .col_in_19               ( u2_col_out_19      ),
    .col_in_20               ( u2_col_out_20      ),
    .col_in_21               ( u2_col_out_21      ),
    .col_in_22               ( u2_col_out_22      ),
    .col_in_23               ( u2_col_out_23      ),
    .col_in_24               ( u2_col_out_24      ),
    .col_in_25               ( u2_col_out_25      ),
    .col_in_26               ( u2_col_out_26      ),
    .col_in_27               ( u2_col_out_27      ),
    .col_in_28               ( u2_col_out_28      ),
    .col_in_29               ( u2_col_out_29      ),
    .col_in_30               ( u2_col_out_30      ),
    .col_in_31               ( u2_col_out_31      ),
    .col_in_32               ( u2_col_out_32      ),
    .col_in_33               ( u2_col_out_33      ),
    .col_in_34               ( u2_col_out_34      ),
    .col_in_35               ( u2_col_out_35      ),
    .col_in_36               ( u2_col_out_36      ),
    .col_in_37               ( u2_col_out_37      ),
    .col_in_38               ( u2_col_out_38      ),
    .col_in_39               ( u2_col_out_39      ),
    .col_in_40               ( u2_col_out_40      ),
    .col_in_41               ( u2_col_out_41      ),
    .col_in_42               ( u2_col_out_42      ),
    .col_in_43               ( u2_col_out_43      ),
    .col_in_44               ( u2_col_out_44      ),
    .col_in_45               ( u2_col_out_45      ),
    .col_in_46               ( u2_col_out_46      ),
    .col_in_47               ( u2_col_out_47      ),
    .col_in_48               ( u2_col_out_48      ),
    .col_in_49               ( u2_col_out_49      ),
    .col_in_50               ( u2_col_out_50      ),
    .col_in_51               ( u2_col_out_51      ),
    .col_in_52               ( u2_col_out_52      ),
    .col_in_53               ( u2_col_out_53      ),
    .col_in_54               ( u2_col_out_54      ),
    .col_in_55               ( u2_col_out_55      ),
    .col_in_56               ( u2_col_out_56      ),
    .col_in_57               ( u2_col_out_57      ),
    .col_in_58               ( u2_col_out_58      ),
    .col_in_59               ( u2_col_out_59      ),
    .col_in_60               ( u2_col_out_60      ),
    .col_in_61               ( u2_col_out_61      ),
    .col_in_62               ( u2_col_out_62      ),
    .col_in_63               ( u2_col_out_63      ),
    .col_in_64               ( u2_col_out_64      ),
    .col_in_65               ( u2_col_out_65      ),
    .col_in_66               ( u2_col_out_66      ),
    .col_in_67               ( u2_col_out_67      ),
    .col_in_68               ( u2_col_out_68      ),
    .col_in_69               ( u2_col_out_69      ),
    .col_in_70               ( u2_col_out_70      ),
    .col_in_71               ( u2_col_out_71      ),
    .col_in_72               ( u2_col_out_72      ),
    .col_in_73               ( u2_col_out_73      ),
    .col_in_74               ( u2_col_out_74      ),
    .col_in_75               ( u2_col_out_75      ),
    .col_in_76               ( u2_col_out_76      ),
    .col_in_77               ( u2_col_out_77      ),
    .col_in_78               ( u2_col_out_78      ),
    .col_in_79               ( u2_col_out_79      ),
    .col_in_80               ( u2_col_out_80      ),
    .col_in_81               ( u2_col_out_81      ),
    .col_in_82               ( u2_col_out_82      ),
    .col_in_83               ( u2_col_out_83      ),
    .col_in_84               ( u2_col_out_84      ),
    .col_in_85               ( u2_col_out_85      ),
    .col_in_86               ( u2_col_out_86      ),
    .col_in_87               ( u2_col_out_87      ),
    .col_in_88               ( u2_col_out_88      ),
    .col_in_89               ( u2_col_out_89      ),
    .col_in_90               ( u2_col_out_90      ),
    .col_in_91               ( u2_col_out_91      ),
    .col_in_92               ( u2_col_out_92      ),
    .col_in_93               ( u2_col_out_93      ),
    .col_in_94               ( u2_col_out_94      ),
    .col_in_95               ( u2_col_out_95      ),
    .col_in_96               ( u2_col_out_96      ),
    .col_in_97               ( u2_col_out_97      ),
    .col_in_98               ( u2_col_out_98      ),
    .col_in_99               ( u2_col_out_99      ),
    .col_in_100              ( u2_col_out_100     ),
    .col_in_101              ( u2_col_out_101     ),
    .col_in_102              ( u2_col_out_102     ),
    .col_in_103              ( u2_col_out_103     ),
    .col_in_104              ( u2_col_out_104     ),
    .col_in_105              ( u2_col_out_105     ),
    .col_in_106              ( u2_col_out_106     ),
    .col_in_107              ( u2_col_out_107     ),
    .col_in_108              ( u2_col_out_108     ),
    .col_in_109              ( u2_col_out_109     ),
    .col_in_110              ( u2_col_out_110     ),
    .col_in_111              ( u2_col_out_111     ),
    .col_in_112              ( u2_col_out_112     ),
    .col_in_113              ( u2_col_out_113     ),
    .col_in_114              ( u2_col_out_114     ),
    .col_in_115              ( u2_col_out_115     ),
    .col_in_116              ( u2_col_out_116     ),
    .col_in_117              ( u2_col_out_117     ),
    .col_in_118              ( u2_col_out_118     ),
    .col_in_119              ( u2_col_out_119     ),
    .col_in_120              ( u2_col_out_120     ),
    .col_in_121              ( u2_col_out_121     ),
    .col_in_122              ( u2_col_out_122     ),
    .col_in_123              ( u2_col_out_123     ),
    .col_in_124              ( u2_col_out_124     ),
    .col_in_125              ( u2_col_out_125     ),
    .col_in_126              ( u2_col_out_126     ),
    .col_in_127              ( u2_col_out_127     ),
    .col_in_128              ( u2_col_out_128     ),
    .col_in_129              ( u2_col_out_129     ),
    .col_in_130              ( u2_col_out_130     ),
    .col_in_131              ( u2_col_out_131     ),
    .col_in_132              ( u2_col_out_132     ),
    .col_in_133              ( u2_col_out_133     ),
    .col_in_134              ( u2_col_out_134     ),
    .col_in_135              ( u2_col_out_135     ),
    .col_in_136              ( u2_col_out_136     ),
    .col_in_137              ( u2_col_out_137     ),
    .col_in_138              ( u2_col_out_138     ),
    .col_in_139              ( u2_col_out_139     ),
    .col_in_140              ( u2_col_out_140     ),
    .col_in_141              ( u2_col_out_141     ),
    .col_in_142              ( u2_col_out_142     ),
    .col_in_143              ( u2_col_out_143     ),
    .col_in_144              ( u2_col_out_144     ),
    .col_in_145              ( u2_col_out_145     ),
    .col_in_146              ( u2_col_out_146     ),
    .col_in_147              ( u2_col_out_147     ),
    .col_in_148              ( u2_col_out_148     ),
    .col_in_149              ( u2_col_out_149     ),
    .col_in_150              ( u2_col_out_150     ),
    .col_in_151              ( u2_col_out_151     ),
    .col_in_152              ( u2_col_out_152     ),
    .col_in_153              ( u2_col_out_153     ),
    .col_in_154              ( u2_col_out_154     ),
    .col_in_155              ( u2_col_out_155     ),
    .col_in_156              ( u2_col_out_156     ),
    .col_in_157              ( u2_col_out_157     ),
    .col_in_158              ( u2_col_out_158     ),
    .col_in_159              ( u2_col_out_159     ),
    .col_in_160              ( u2_col_out_160     ),
    .col_in_161              ( u2_col_out_161     ),
    .col_in_162              ( u2_col_out_162     ),
    .col_in_163              ( u2_col_out_163     ),
    .col_in_164              ( u2_col_out_164     ),
    .col_in_165              ( u2_col_out_165     ),
    .col_in_166              ( u2_col_out_166     ),
    .col_in_167              ( u2_col_out_167     ),
    .col_in_168              ( u2_col_out_168     ),
    .col_in_169              ( u2_col_out_169     ),
    .col_in_170              ( u2_col_out_170     ),
    .col_in_171              ( u2_col_out_171     ),
    .col_in_172              ( u2_col_out_172     ),
    .col_in_173              ( u2_col_out_173     ),
    .col_in_174              ( u2_col_out_174     ),
    .col_in_175              ( u2_col_out_175     ),
    .col_in_176              ( u2_col_out_176     ),
    .col_in_177              ( u2_col_out_177     ),
    .col_in_178              ( u2_col_out_178     ),
    .col_in_179              ( u2_col_out_179     ),
    .col_in_180              ( u2_col_out_180     ),
    .col_in_181              ( u2_col_out_181     ),
    .col_in_182              ( u2_col_out_182     ),
    .col_in_183              ( u2_col_out_183     ),
    .col_in_184              ( u2_col_out_184     ),
    .col_in_185              ( u2_col_out_185     ),
    .col_in_186              ( u2_col_out_186     ),
    .col_in_187              ( u2_col_out_187     ),
    .col_in_188              ( u2_col_out_188     ),
    .col_in_189              ( u2_col_out_189     ),
    .col_in_190              ( u2_col_out_190     ),
    .col_in_191              ( u2_col_out_191     ),
    .col_in_192              ( u2_col_out_192     ),
    .col_in_193              ( u2_col_out_193     ),
    .col_in_194              ( u2_col_out_194     ),
    .col_in_195              ( u2_col_out_195     ),
    .col_in_196              ( u2_col_out_196     ),
    .col_in_197              ( u2_col_out_197     ),
    .col_in_198              ( u2_col_out_198     ),
    .col_in_199              ( u2_col_out_199     ),
    .col_in_200              ( u2_col_out_200     ),
    .col_in_201              ( u2_col_out_201     ),
    .col_in_202              ( u2_col_out_202     ),
    .col_in_203              ( u2_col_out_203     ),
    .col_in_204              ( u2_col_out_204     ),
    .col_in_205              ( u2_col_out_205     ),
    .col_in_206              ( u2_col_out_206     ),
    .col_in_207              ( u2_col_out_207     ),
    .col_in_208              ( u2_col_out_208     ),
    .col_in_209              ( u2_col_out_209     ),
    .col_in_210              ( u2_col_out_210     ),
    .col_in_211              ( u2_col_out_211     ),
    .col_in_212              ( u2_col_out_212     ),
    .col_in_213              ( u2_col_out_213     ),
    .col_in_214              ( u2_col_out_214     ),
    .col_in_215              ( u2_col_out_215     ),
    .col_in_216              ( u2_col_out_216     ),
    .col_in_217              ( u2_col_out_217     ),
    .col_in_218              ( u2_col_out_218     ),
    .col_in_219              ( u2_col_out_219     ),
    .col_in_220              ( u2_col_out_220     ),
    .col_in_221              ( u2_col_out_221     ),
    .col_in_222              ( u2_col_out_222     ),
    .col_in_223              ( u2_col_out_223     ),
    .col_in_224              ( u2_col_out_224     ),
    .col_in_225              ( u2_col_out_225     ),
    .col_in_226              ( u2_col_out_226     ),
    .col_in_227              ( u2_col_out_227     ),
    .col_in_228              ( u2_col_out_228     ),
    .col_in_229              ( u2_col_out_229     ),
    .col_in_230              ( u2_col_out_230     ),
    .col_in_231              ( u2_col_out_231     ),
    .col_in_232              ( u2_col_out_232     ),
    .col_in_233              ( u2_col_out_233     ),
    .col_in_234              ( u2_col_out_234     ),
    .col_in_235              ( u2_col_out_235     ),
    .col_in_236              ( u2_col_out_236     ),
    .col_in_237              ( u2_col_out_237     ),
    .col_in_238              ( u2_col_out_238     ),
    .col_in_239              ( u2_col_out_239     ),
    .col_in_240              ( u2_col_out_240     ),
    .col_in_241              ( u2_col_out_241     ),
    .col_in_242              ( u2_col_out_242     ),
    .col_in_243              ( u2_col_out_243     ),
    .col_in_244              ( u2_col_out_244     ),
    .col_in_245              ( u2_col_out_245     ),
    .col_in_246              ( u2_col_out_246     ),
    .col_in_247              ( u2_col_out_247     ),
    .col_in_248              ( u2_col_out_248     ),
    .col_in_249              ( u2_col_out_249     ),
    .col_in_250              ( u2_col_out_250     ),
    .col_in_251              ( u2_col_out_251     ),
    .col_in_252              ( u2_col_out_252     ),
    .col_in_253              ( u2_col_out_253     ),
    .col_in_254              ( u2_col_out_254     ),
    .col_in_255              ( u2_col_out_255     ),
    .col_in_256              ( u2_col_out_256     ),
    .col_in_257              ( u2_col_out_257     ),
    .col_in_258              ( u2_col_out_258     ),
    .col_in_259              ( u2_col_out_259     ),
    .col_in_260              ( u2_col_out_260     ),
    .col_in_261              ( u2_col_out_261     ),
    .col_in_262              ( u2_col_out_262     ),
    .col_in_263              ( u2_col_out_263     ),
    .col_in_264              ( u2_col_out_264     ),
    .col_in_265              ( u2_col_out_265     ),
    .col_in_266              ( u2_col_out_266     ),
    .col_in_267              ( u2_col_out_267     ),
    .col_in_268              ( u2_col_out_268     ),
    .col_in_269              ( u2_col_out_269     ),
    .col_in_270              ( u2_col_out_270     ),
    .col_in_271              ( u2_col_out_271     ),
    .col_in_272              ( u2_col_out_272     ),
    .col_in_273              ( u2_col_out_273     ),
    .col_in_274              ( u2_col_out_274     ),
    .col_in_275              ( u2_col_out_275     ),
    .col_in_276              ( u2_col_out_276     ),
    .col_in_277              ( u2_col_out_277     ),
    .col_in_278              ( u2_col_out_278     ),
    .col_in_279              ( u2_col_out_279     ),
    .col_in_280              ( u2_col_out_280     ),
    .col_in_281              ( u2_col_out_281     ),
    .col_in_282              ( u2_col_out_282     ),
    .col_in_283              ( u2_col_out_283     ),
    .col_in_284              ( u2_col_out_284     ),
    .col_in_285              ( u2_col_out_285     ),
    .col_in_286              ( u2_col_out_286     ),
    .col_in_287              ( u2_col_out_287     ),
    .col_in_288              ( u2_col_out_288     ),
    .col_in_289              ( u2_col_out_289     ),
    .col_in_290              ( u2_col_out_290     ),
    .col_in_291              ( u2_col_out_291     ),
    .col_in_292              ( u2_col_out_292     ),
    .col_in_293              ( u2_col_out_293     ),
    .col_in_294              ( u2_col_out_294     ),
    .col_in_295              ( u2_col_out_295     ),
    .col_in_296              ( u2_col_out_296     ),
    .col_in_297              ( u2_col_out_297     ),
    .col_in_298              ( u2_col_out_298     ),
    .col_in_299              ( u2_col_out_299     ),
    .col_in_300              ( u2_col_out_300     ),
    .col_in_301              ( u2_col_out_301     ),
    .col_in_302              ( u2_col_out_302     ),
    .col_in_303              ( u2_col_out_303     ),
    .col_in_304              ( u2_col_out_304     ),
    .col_in_305              ( u2_col_out_305     ),
    .col_in_306              ( u2_col_out_306     ),
    .col_in_307              ( u2_col_out_307     ),
    .col_in_308              ( u2_col_out_308     ),
    .col_in_309              ( u2_col_out_309     ),
    .col_in_310              ( u2_col_out_310     ),
    .col_in_311              ( u2_col_out_311     ),
    .col_in_312              ( u2_col_out_312     ),
    .col_in_313              ( u2_col_out_313     ),
    .col_in_314              ( u2_col_out_314     ),
    .col_in_315              ( u2_col_out_315     ),
    .col_in_316              ( u2_col_out_316     ),
    .col_in_317              ( u2_col_out_317     ),
    .col_in_318              ( u2_col_out_318     ),
    .col_in_319              ( u2_col_out_319     ),
    .col_in_320              ( u2_col_out_320     ),
    .col_in_321              ( u2_col_out_321     ),
    .col_in_322              ( u2_col_out_322     ),
    .col_in_323              ( u2_col_out_323     ),
    .col_in_324              ( u2_col_out_324     ),
    .col_in_325              ( u2_col_out_325     ),
    .col_in_326              ( u2_col_out_326     ),
    .col_in_327              ( u2_col_out_327     ),
    .col_in_328              ( u2_col_out_328     ),
    .col_in_329              ( u2_col_out_329     ),
    .col_in_330              ( u2_col_out_330     ),
    .col_in_331              ( u2_col_out_331     ),
    .col_in_332              ( u2_col_out_332     ),
    .col_in_333              ( u2_col_out_333     ),
    .col_in_334              ( u2_col_out_334     ),
    .col_in_335              ( u2_col_out_335     ),
    .col_in_336              ( u2_col_out_336     ),
    .col_in_337              ( u2_col_out_337     ),
    .col_in_338              ( u2_col_out_338     ),
    .col_in_339              ( u2_col_out_339     ),
    .col_in_340              ( u2_col_out_340     ),
    .col_in_341              ( u2_col_out_341     ),
    .col_in_342              ( u2_col_out_342     ),
    .col_in_343              ( u2_col_out_343     ),
    .col_in_344              ( u2_col_out_344     ),
    .col_in_345              ( u2_col_out_345     ),
    .col_in_346              ( u2_col_out_346     ),
    .col_in_347              ( u2_col_out_347     ),
    .col_in_348              ( u2_col_out_348     ),
    .col_in_349              ( u2_col_out_349     ),
    .col_in_350              ( u2_col_out_350     ),
    .col_in_351              ( u2_col_out_351     ),
    .col_in_352              ( u2_col_out_352     ),
    .col_in_353              ( u2_col_out_353     ),
    .col_in_354              ( u2_col_out_354     ),
    .col_in_355              ( u2_col_out_355     ),
    .col_in_356              ( u2_col_out_356     ),
    .col_in_357              ( u2_col_out_357     ),
    .col_in_358              ( u2_col_out_358     ),
    .col_in_359              ( u2_col_out_359     ),
    .col_in_360              ( u2_col_out_360     ),
    .col_in_361              ( u2_col_out_361     ),
    .col_in_362              ( u2_col_out_362     ),
    .col_in_363              ( u2_col_out_363     ),
    .col_in_364              ( u2_col_out_364     ),
    .col_in_365              ( u2_col_out_365     ),
    .col_in_366              ( u2_col_out_366     ),
    .col_in_367              ( u2_col_out_367     ),
    .col_in_368              ( u2_col_out_368     ),
    .col_in_369              ( u2_col_out_369     ),
    .col_in_370              ( u2_col_out_370     ),
    .col_in_371              ( u2_col_out_371     ),
    .col_in_372              ( u2_col_out_372     ),
    .col_in_373              ( u2_col_out_373     ),
    .col_in_374              ( u2_col_out_374     ),
    .col_in_375              ( u2_col_out_375     ),
    .col_in_376              ( u2_col_out_376     ),
    .col_in_377              ( u2_col_out_377     ),
    .col_in_378              ( u2_col_out_378     ),
    .col_in_379              ( u2_col_out_379     ),
    .col_in_380              ( u2_col_out_380     ),
    .col_in_381              ( u2_col_out_381     ),
    .col_in_382              ( u2_col_out_382     ),
    .col_in_383              ( u2_col_out_383     ),
    .col_in_384              ( u2_col_out_384     ),
    .col_in_385              ( u2_col_out_385     ),
    .col_in_386              ( u2_col_out_386     ),
    .col_in_387              ( u2_col_out_387     ),
    .col_in_388              ( u2_col_out_388     ),
    .col_in_389              ( u2_col_out_389     ),
    .col_in_390              ( u2_col_out_390     ),
    .col_in_391              ( u2_col_out_391     ),
    .col_in_392              ( u2_col_out_392     ),
    .col_in_393              ( u2_col_out_393     ),
    .col_in_394              ( u2_col_out_394     ),
    .col_in_395              ( u2_col_out_395     ),
    .col_in_396              ( u2_col_out_396     ),
    .col_in_397              ( u2_col_out_397     ),
    .col_in_398              ( u2_col_out_398     ),
    .col_in_399              ( u2_col_out_399     ),
    .col_in_400              ( u2_col_out_400     ),
    .col_in_401              ( u2_col_out_401     ),
    .col_in_402              ( u2_col_out_402     ),
    .col_in_403              ( u2_col_out_403     ),
    .col_in_404              ( u2_col_out_404     ),
    .col_in_405              ( u2_col_out_405     ),
    .col_in_406              ( u2_col_out_406     ),
    .col_in_407              ( u2_col_out_407     ),
    .col_in_408              ( u2_col_out_408     ),
    .col_in_409              ( u2_col_out_409     ),
    .col_in_410              ( u2_col_out_410     ),
    .col_in_411              ( u2_col_out_411     ),
    .col_in_412              ( u2_col_out_412     ),
    .col_in_413              ( u2_col_out_413     ),
    .col_in_414              ( u2_col_out_414     ),
    .col_in_415              ( u2_col_out_415     ),
    .col_in_416              ( u2_col_out_416     ),
    .col_in_417              ( u2_col_out_417     ),
    .col_in_418              ( u2_col_out_418     ),
    .col_in_419              ( u2_col_out_419     ),
    .col_in_420              ( u2_col_out_420     ),
    .col_in_421              ( u2_col_out_421     ),
    .col_in_422              ( u2_col_out_422     ),
    .col_in_423              ( u2_col_out_423     ),
    .col_in_424              ( u2_col_out_424     ),
    .col_in_425              ( u2_col_out_425     ),
    .col_in_426              ( u2_col_out_426     ),
    .col_in_427              ( u2_col_out_427     ),
    .col_in_428              ( u2_col_out_428     ),
    .col_in_429              ( u2_col_out_429     ),
    .col_in_430              ( u2_col_out_430     ),
    .col_in_431              ( u2_col_out_431     ),
    .col_in_432              ( u2_col_out_432     ),
    .col_in_433              ( u2_col_out_433     ),
    .col_in_434              ( u2_col_out_434     ),
    .col_in_435              ( u2_col_out_435     ),
    .col_in_436              ( u2_col_out_436     ),
    .col_in_437              ( u2_col_out_437     ),
    .col_in_438              ( u2_col_out_438     ),
    .col_in_439              ( u2_col_out_439     ),
    .col_in_440              ( u2_col_out_440     ),
    .col_in_441              ( u2_col_out_441     ),
    .col_in_442              ( u2_col_out_442     ),
    .col_in_443              ( u2_col_out_443     ),
    .col_in_444              ( u2_col_out_444     ),
    .col_in_445              ( u2_col_out_445     ),
    .col_in_446              ( u2_col_out_446     ),
    .col_in_447              ( u2_col_out_447     ),
    .col_in_448              ( u2_col_out_448     ),
    .col_in_449              ( u2_col_out_449     ),
    .col_in_450              ( u2_col_out_450     ),
    .col_in_451              ( u2_col_out_451     ),
    .col_in_452              ( u2_col_out_452     ),
    .col_in_453              ( u2_col_out_453     ),
    .col_in_454              ( u2_col_out_454     ),
    .col_in_455              ( u2_col_out_455     ),
    .col_in_456              ( u2_col_out_456     ),
    .col_in_457              ( u2_col_out_457     ),
    .col_in_458              ( u2_col_out_458     ),
    .col_in_459              ( u2_col_out_459     ),
    .col_in_460              ( u2_col_out_460     ),
    .col_in_461              ( u2_col_out_461     ),
    .col_in_462              ( u2_col_out_462     ),
    .col_in_463              ( u2_col_out_463     ),
    .col_in_464              ( u2_col_out_464     ),
    .col_in_465              ( u2_col_out_465     ),
    .col_in_466              ( u2_col_out_466     ),
    .col_in_467              ( u2_col_out_467     ),
    .col_in_468              ( u2_col_out_468     ),
    .col_in_469              ( u2_col_out_469     ),
    .col_in_470              ( u2_col_out_470     ),
    .col_in_471              ( u2_col_out_471     ),
    .col_in_472              ( u2_col_out_472     ),
    .col_in_473              ( u2_col_out_473     ),
    .col_in_474              ( u2_col_out_474     ),
    .col_in_475              ( u2_col_out_475     ),
    .col_in_476              ( u2_col_out_476     ),
    .col_in_477              ( u2_col_out_477     ),
    .col_in_478              ( u2_col_out_478     ),
    .col_in_479              ( u2_col_out_479     ),
    .col_in_480              ( u2_col_out_480     ),
    .col_in_481              ( u2_col_out_481     ),
    .col_in_482              ( u2_col_out_482     ),
    .col_in_483              ( u2_col_out_483     ),
    .col_in_484              ( u2_col_out_484     ),
    .col_in_485              ( u2_col_out_485     ),
    .col_in_486              ( u2_col_out_486     ),
    .col_in_487              ( u2_col_out_487     ),
    .col_in_488              ( u2_col_out_488     ),
    .col_in_489              ( u2_col_out_489     ),
    .col_in_490              ( u2_col_out_490     ),
    .col_in_491              ( u2_col_out_491     ),
    .col_in_492              ( u2_col_out_492     ),
    .col_in_493              ( u2_col_out_493     ),
    .col_in_494              ( u2_col_out_494     ),
    .col_in_495              ( u2_col_out_495     ),
    .col_in_496              ( u2_col_out_496     ),
    .col_in_497              ( u2_col_out_497     ),
    .col_in_498              ( u2_col_out_498     ),
    .col_in_499              ( u2_col_out_499     ),
    .col_in_500              ( u2_col_out_500     ),
    .col_in_501              ( u2_col_out_501     ),
    .col_in_502              ( u2_col_out_502     ),
    .col_in_503              ( u2_col_out_503     ),
    .col_in_504              ( u2_col_out_504     ),
    .col_in_505              ( u2_col_out_505     ),
    .col_in_506              ( u2_col_out_506     ),
    .col_in_507              ( u2_col_out_507     ),
    .col_in_508              ( u2_col_out_508     ),
    .col_in_509              ( u2_col_out_509     ),
    .col_in_510              ( u2_col_out_510     ),
    .col_in_511              ( u2_col_out_511     ),
    .col_in_512              ( u2_col_out_512     ),
    .col_in_513              ( u2_col_out_513     ),
    .col_in_514              ( u2_col_out_514     ),
    .col_in_515              ( u2_col_out_515     ),
    .col_in_516              ( u2_col_out_516     ),
    .col_in_517              ( u2_col_out_517     ),
    .col_in_518              ( u2_col_out_518     ),
    .col_in_519              ( u2_col_out_519     ),
    .col_in_520              ( u2_col_out_520     ),
    .col_in_521              ( u2_col_out_521     ),
    .col_in_522              ( u2_col_out_522     ),
    .col_in_523              ( u2_col_out_523     ),
    .col_in_524              ( u2_col_out_524     ),
    .col_in_525              ( u2_col_out_525     ),
    .col_in_526              ( u2_col_out_526     ),
    .col_in_527              ( u2_col_out_527     ),
    .col_in_528              ( u2_col_out_528     ),
    .col_in_529              ( u2_col_out_529     ),
    .col_in_530              ( u2_col_out_530     ),
    .col_in_531              ( u2_col_out_531     ),
    .col_in_532              ( u2_col_out_532     ),
    .col_in_533              ( u2_col_out_533     ),
    .col_in_534              ( u2_col_out_534     ),
    .col_in_535              ( u2_col_out_535     ),
    .col_in_536              ( u2_col_out_536     ),
    .col_in_537              ( u2_col_out_537     ),
    .col_in_538              ( u2_col_out_538     ),
    .col_in_539              ( u2_col_out_539     ),
    .col_in_540              ( u2_col_out_540     ),
    .col_in_541              ( u2_col_out_541     ),
    .col_in_542              ( u2_col_out_542     ),
    .col_in_543              ( u2_col_out_543     ),
    .col_in_544              ( u2_col_out_544     ),
    .col_in_545              ( u2_col_out_545     ),
    .col_in_546              ( u2_col_out_546     ),
    .col_in_547              ( u2_col_out_547     ),
    .col_in_548              ( u2_col_out_548     ),
    .col_in_549              ( u2_col_out_549     ),
    .col_in_550              ( u2_col_out_550     ),
    .col_in_551              ( u2_col_out_551     ),
    .col_in_552              ( u2_col_out_552     ),
    .col_in_553              ( u2_col_out_553     ),
    .col_in_554              ( u2_col_out_554     ),
    .col_in_555              ( u2_col_out_555     ),
    .col_in_556              ( u2_col_out_556     ),
    .col_in_557              ( u2_col_out_557     ),
    .col_in_558              ( u2_col_out_558     ),
    .col_in_559              ( u2_col_out_559     ),
    .col_in_560              ( u2_col_out_560     ),
    .col_in_561              ( u2_col_out_561     ),
    .col_in_562              ( u2_col_out_562     ),
    .col_in_563              ( u2_col_out_563     ),
    .col_in_564              ( u2_col_out_564     ),
    .col_in_565              ( u2_col_out_565     ),
    .col_in_566              ( u2_col_out_566     ),
    .col_in_567              ( u2_col_out_567     ),
    .col_in_568              ( u2_col_out_568     ),
    .col_in_569              ( u2_col_out_569     ),
    .col_in_570              ( u2_col_out_570     ),
    .col_in_571              ( u2_col_out_571     ),
    .col_in_572              ( u2_col_out_572     ),
    .col_in_573              ( u2_col_out_573     ),
    .col_in_574              ( u2_col_out_574     ),
    .col_in_575              ( u2_col_out_575     ),
    .col_in_576              ( u2_col_out_576     ),
    .col_in_577              ( u2_col_out_577     ),
    .col_in_578              ( u2_col_out_578     ),
    .col_in_579              ( u2_col_out_579     ),
    .col_in_580              ( u2_col_out_580     ),
    .col_in_581              ( u2_col_out_581     ),
    .col_in_582              ( u2_col_out_582     ),
    .col_in_583              ( u2_col_out_583     ),
    .col_in_584              ( u2_col_out_584     ),
    .col_in_585              ( u2_col_out_585     ),
    .col_in_586              ( u2_col_out_586     ),
    .col_in_587              ( u2_col_out_587     ),
    .col_in_588              ( u2_col_out_588     ),
    .col_in_589              ( u2_col_out_589     ),
    .col_in_590              ( u2_col_out_590     ),
    .col_in_591              ( u2_col_out_591     ),
    .col_in_592              ( u2_col_out_592     ),
    .col_in_593              ( u2_col_out_593     ),
    .col_in_594              ( u2_col_out_594     ),
    .col_in_595              ( u2_col_out_595     ),
    .col_in_596              ( u2_col_out_596     ),
    .col_in_597              ( u2_col_out_597     ),
    .col_in_598              ( u2_col_out_598     ),
    .col_in_599              ( u2_col_out_599     ),
    .col_in_600              ( u2_col_out_600     ),
    .col_in_601              ( u2_col_out_601     ),
    .col_in_602              ( u2_col_out_602     ),
    .col_in_603              ( u2_col_out_603     ),
    .col_in_604              ( u2_col_out_604     ),
    .col_in_605              ( u2_col_out_605     ),
    .col_in_606              ( u2_col_out_606     ),
    .col_in_607              ( u2_col_out_607     ),
    .col_in_608              ( u2_col_out_608     ),
    .col_in_609              ( u2_col_out_609     ),
    .col_in_610              ( u2_col_out_610     ),
    .col_in_611              ( u2_col_out_611     ),
    .col_in_612              ( u2_col_out_612     ),
    .col_in_613              ( u2_col_out_613     ),
    .col_in_614              ( u2_col_out_614     ),
    .col_in_615              ( u2_col_out_615     ),
    .col_in_616              ( u2_col_out_616     ),
    .col_in_617              ( u2_col_out_617     ),
    .col_in_618              ( u2_col_out_618     ),
    .col_in_619              ( u2_col_out_619     ),
    .col_in_620              ( u2_col_out_620     ),
    .col_in_621              ( u2_col_out_621     ),
    .col_in_622              ( u2_col_out_622     ),
    .col_in_623              ( u2_col_out_623     ),
    .col_in_624              ( u2_col_out_624     ),
    .col_in_625              ( u2_col_out_625     ),
    .col_in_626              ( u2_col_out_626     ),
    .col_in_627              ( u2_col_out_627     ),
    .col_in_628              ( u2_col_out_628     ),
    .col_in_629              ( u2_col_out_629     ),
    .col_in_630              ( u2_col_out_630     ),
    .col_in_631              ( u2_col_out_631     ),
    .col_in_632              ( u2_col_out_632     ),
    .col_in_633              ( u2_col_out_633     ),
    .col_in_634              ( u2_col_out_634     ),
    .col_in_635              ( u2_col_out_635     ),
    .col_in_636              ( u2_col_out_636     ),
    .col_in_637              ( u2_col_out_637     ),
    .col_in_638              ( u2_col_out_638     ),
    .col_in_639              ( u2_col_out_639     ),
    .col_in_640              ( u2_col_out_640     ),
    .col_in_641              ( u2_col_out_641     ),
    .col_in_642              ( u2_col_out_642     ),
    .col_in_643              ( u2_col_out_643     ),
    .col_in_644              ( u2_col_out_644     ),
    .col_in_645              ( u2_col_out_645     ),
    .col_in_646              ( u2_col_out_646     ),
    .col_in_647              ( u2_col_out_647     ),
    .col_in_648              ( u2_col_out_648     ),
    .col_in_649              ( u2_col_out_649     ),
    .col_in_650              ( u2_col_out_650     ),
    .col_in_651              ( u2_col_out_651     ),
    .col_in_652              ( u2_col_out_652     ),
    .col_in_653              ( u2_col_out_653     ),
    .col_in_654              ( u2_col_out_654     ),
    .col_in_655              ( u2_col_out_655     ),
    .col_in_656              ( u2_col_out_656     ),
    .col_in_657              ( u2_col_out_657     ),
    .col_in_658              ( u2_col_out_658     ),
    .col_in_659              ( u2_col_out_659     ),
    .col_in_660              ( u2_col_out_660     ),
    .col_in_661              ( u2_col_out_661     ),
    .col_in_662              ( u2_col_out_662     ),
    .col_in_663              ( u2_col_out_663     ),
    .col_in_664              ( u2_col_out_664     ),
    .col_in_665              ( u2_col_out_665     ),
    .col_in_666              ( u2_col_out_666     ),
    .col_in_667              ( u2_col_out_667     ),
    .col_in_668              ( u2_col_out_668     ),
    .col_in_669              ( u2_col_out_669     ),
    .col_in_670              ( u2_col_out_670     ),
    .col_in_671              ( u2_col_out_671     ),
    .col_in_672              ( u2_col_out_672     ),
    .col_in_673              ( u2_col_out_673     ),
    .col_in_674              ( u2_col_out_674     ),
    .col_in_675              ( u2_col_out_675     ),
    .col_in_676              ( u2_col_out_676     ),
    .col_in_677              ( u2_col_out_677     ),
    .col_in_678              ( u2_col_out_678     ),
    .col_in_679              ( u2_col_out_679     ),
    .col_in_680              ( u2_col_out_680     ),
    .col_in_681              ( u2_col_out_681     ),
    .col_in_682              ( u2_col_out_682     ),
    .col_in_683              ( u2_col_out_683     ),
    .col_in_684              ( u2_col_out_684     ),
    .col_in_685              ( u2_col_out_685     ),
    .col_in_686              ( u2_col_out_686     ),
    .col_in_687              ( u2_col_out_687     ),
    .col_in_688              ( u2_col_out_688     ),
    .col_in_689              ( u2_col_out_689     ),
    .col_in_690              ( u2_col_out_690     ),
    .col_in_691              ( u2_col_out_691     ),
    .col_in_692              ( u2_col_out_692     ),
    .col_in_693              ( u2_col_out_693     ),
    .col_in_694              ( u2_col_out_694     ),
    .col_in_695              ( u2_col_out_695     ),
    .col_in_696              ( u2_col_out_696     ),
    .col_in_697              ( u2_col_out_697     ),
    .col_in_698              ( u2_col_out_698     ),
    .col_in_699              ( u2_col_out_699     ),
    .col_in_700              ( u2_col_out_700     ),
    .col_in_701              ( u2_col_out_701     ),
    .col_in_702              ( u2_col_out_702     ),
    .col_in_703              ( u2_col_out_703     ),
    .col_in_704              ( u2_col_out_704     ),
    .col_in_705              ( u2_col_out_705     ),
    .col_in_706              ( u2_col_out_706     ),
    .col_in_707              ( u2_col_out_707     ),
    .col_in_708              ( u2_col_out_708     ),
    .col_in_709              ( u2_col_out_709     ),
    .col_in_710              ( u2_col_out_710     ),
    .col_in_711              ( u2_col_out_711     ),
    .col_in_712              ( u2_col_out_712     ),
    .col_in_713              ( u2_col_out_713     ),
    .col_in_714              ( u2_col_out_714     ),
    .col_in_715              ( u2_col_out_715     ),
    .col_in_716              ( u2_col_out_716     ),
    .col_in_717              ( u2_col_out_717     ),
    .col_in_718              ( u2_col_out_718     ),
    .col_in_719              ( u2_col_out_719     ),
    .col_in_720              ( u2_col_out_720     ),
    .col_in_721              ( u2_col_out_721     ),
    .col_in_722              ( u2_col_out_722     ),
    .col_in_723              ( u2_col_out_723     ),
    .col_in_724              ( u2_col_out_724     ),
    .col_in_725              ( u2_col_out_725     ),
    .col_in_726              ( u2_col_out_726     ),
    .col_in_727              ( u2_col_out_727     ),
    .col_in_728              ( u2_col_out_728     ),
    .col_in_729              ( u2_col_out_729     ),
    .col_in_730              ( u2_col_out_730     ),
    .col_in_731              ( u2_col_out_731     ),
    .col_in_732              ( u2_col_out_732     ),
    .col_in_733              ( u2_col_out_733     ),
    .col_in_734              ( u2_col_out_734     ),
    .col_in_735              ( u2_col_out_735     ),
    .col_in_736              ( u2_col_out_736     ),
    .col_in_737              ( u2_col_out_737     ),
    .col_in_738              ( u2_col_out_738     ),
    .col_in_739              ( u2_col_out_739     ),
    .col_in_740              ( u2_col_out_740     ),
    .col_in_741              ( u2_col_out_741     ),
    .col_in_742              ( u2_col_out_742     ),
    .col_in_743              ( u2_col_out_743     ),
    .col_in_744              ( u2_col_out_744     ),
    .col_in_745              ( u2_col_out_745     ),
    .col_in_746              ( u2_col_out_746     ),
    .col_in_747              ( u2_col_out_747     ),
    .col_in_748              ( u2_col_out_748     ),
    .col_in_749              ( u2_col_out_749     ),
    .col_in_750              ( u2_col_out_750     ),
    .col_in_751              ( u2_col_out_751     ),
    .col_in_752              ( u2_col_out_752     ),
    .col_in_753              ( u2_col_out_753     ),
    .col_in_754              ( u2_col_out_754     ),
    .col_in_755              ( u2_col_out_755     ),
    .col_in_756              ( u2_col_out_756     ),
    .col_in_757              ( u2_col_out_757     ),
    .col_in_758              ( u2_col_out_758     ),
    .col_in_759              ( u2_col_out_759     ),
    .col_in_760              ( u2_col_out_760     ),
    .col_in_761              ( u2_col_out_761     ),
    .col_in_762              ( u2_col_out_762     ),
    .col_in_763              ( u2_col_out_763     ),
    .col_in_764              ( u2_col_out_764     ),
    .col_in_765              ( u2_col_out_765     ),
    .col_in_766              ( u2_col_out_766     ),
    .col_in_767              ( u2_col_out_767     ),
    .col_in_768              ( u2_col_out_768     ),
    .col_in_769              ( u2_col_out_769     ),
    .col_in_770              ( u2_col_out_770     ),
    .col_in_771              ( u2_col_out_771     ),
    .col_in_772              ( u2_col_out_772     ),
    .col_in_773              ( u2_col_out_773     ),
    .col_in_774              ( u2_col_out_774     ),
    .col_in_775              ( u2_col_out_775     ),
    .col_in_776              ( u2_col_out_776     ),
    .col_in_777              ( u2_col_out_777     ),
    .col_in_778              ( u2_col_out_778     ),
    .col_in_779              ( u2_col_out_779     ),
    .col_in_780              ( u2_col_out_780     ),
    .col_in_781              ( u2_col_out_781     ),
    .col_in_782              ( u2_col_out_782     ),
    .col_in_783              ( u2_col_out_783     ),
    .col_in_784              ( u2_col_out_784     ),
    .col_in_785              ( u2_col_out_785     ),
    .col_in_786              ( u2_col_out_786     ),
    .col_in_787              ( u2_col_out_787     ),
    .col_in_788              ( u2_col_out_788     ),
    .col_in_789              ( u2_col_out_789     ),
    .col_in_790              ( u2_col_out_790     ),
    .col_in_791              ( u2_col_out_791     ),
    .col_in_792              ( u2_col_out_792     ),
    .col_in_793              ( u2_col_out_793     ),
    .col_in_794              ( u2_col_out_794     ),
    .col_in_795              ( u2_col_out_795     ),
    .col_in_796              ( u2_col_out_796     ),
    .col_in_797              ( u2_col_out_797     ),
    .col_in_798              ( u2_col_out_798     ),
    .col_in_799              ( u2_col_out_799     ),
    .col_in_800              ( u2_col_out_800     ),
    .col_in_801              ( u2_col_out_801     ),
    .col_in_802              ( u2_col_out_802     ),
    .col_in_803              ( u2_col_out_803     ),
    .col_in_804              ( u2_col_out_804     ),
    .col_in_805              ( u2_col_out_805     ),
    .col_in_806              ( u2_col_out_806     ),
    .col_in_807              ( u2_col_out_807     ),
    .col_in_808              ( u2_col_out_808     ),
    .col_in_809              ( u2_col_out_809     ),
    .col_in_810              ( u2_col_out_810     ),
    .col_in_811              ( u2_col_out_811     ),
    .col_in_812              ( u2_col_out_812     ),
    .col_in_813              ( u2_col_out_813     ),
    .col_in_814              ( u2_col_out_814     ),
    .col_in_815              ( u2_col_out_815     ),
    .col_in_816              ( u2_col_out_816     ),
    .col_in_817              ( u2_col_out_817     ),
    .col_in_818              ( u2_col_out_818     ),
    .col_in_819              ( u2_col_out_819     ),
    .col_in_820              ( u2_col_out_820     ),
    .col_in_821              ( u2_col_out_821     ),
    .col_in_822              ( u2_col_out_822     ),
    .col_in_823              ( u2_col_out_823     ),
    .col_in_824              ( u2_col_out_824     ),
    .col_in_825              ( u2_col_out_825     ),
    .col_in_826              ( u2_col_out_826     ),
    .col_in_827              ( u2_col_out_827     ),
    .col_in_828              ( u2_col_out_828     ),
    .col_in_829              ( u2_col_out_829     ),
    .col_in_830              ( u2_col_out_830     ),
    .col_in_831              ( u2_col_out_831     ),
    .col_in_832              ( u2_col_out_832     ),
    .col_in_833              ( u2_col_out_833     ),
    .col_in_834              ( u2_col_out_834     ),
    .col_in_835              ( u2_col_out_835     ),
    .col_in_836              ( u2_col_out_836     ),
    .col_in_837              ( u2_col_out_837     ),
    .col_in_838              ( u2_col_out_838     ),
    .col_in_839              ( u2_col_out_839     ),
    .col_in_840              ( u2_col_out_840     ),
    .col_in_841              ( u2_col_out_841     ),
    .col_in_842              ( u2_col_out_842     ),
    .col_in_843              ( u2_col_out_843     ),
    .col_in_844              ( u2_col_out_844     ),
    .col_in_845              ( u2_col_out_845     ),
    .col_in_846              ( u2_col_out_846     ),
    .col_in_847              ( u2_col_out_847     ),
    .col_in_848              ( u2_col_out_848     ),
    .col_in_849              ( u2_col_out_849     ),
    .col_in_850              ( u2_col_out_850     ),
    .col_in_851              ( u2_col_out_851     ),
    .col_in_852              ( u2_col_out_852     ),
    .col_in_853              ( u2_col_out_853     ),
    .col_in_854              ( u2_col_out_854     ),
    .col_in_855              ( u2_col_out_855     ),
    .col_in_856              ( u2_col_out_856     ),
    .col_in_857              ( u2_col_out_857     ),
    .col_in_858              ( u2_col_out_858     ),
    .col_in_859              ( u2_col_out_859     ),
    .col_in_860              ( u2_col_out_860     ),
    .col_in_861              ( u2_col_out_861     ),
    .col_in_862              ( u2_col_out_862     ),
    .col_in_863              ( u2_col_out_863     ),
    .col_in_864              ( u2_col_out_864     ),
    .col_in_865              ( u2_col_out_865     ),
    .col_in_866              ( u2_col_out_866     ),
    .col_in_867              ( u2_col_out_867     ),
    .col_in_868              ( u2_col_out_868     ),
    .col_in_869              ( u2_col_out_869     ),
    .col_in_870              ( u2_col_out_870     ),
    .col_in_871              ( u2_col_out_871     ),
    .col_in_872              ( u2_col_out_872     ),
    .col_in_873              ( u2_col_out_873     ),
    .col_in_874              ( u2_col_out_874     ),
    .col_in_875              ( u2_col_out_875     ),
    .col_in_876              ( u2_col_out_876     ),
    .col_in_877              ( u2_col_out_877     ),
    .col_in_878              ( u2_col_out_878     ),
    .col_in_879              ( u2_col_out_879     ),
    .col_in_880              ( u2_col_out_880     ),
    .col_in_881              ( u2_col_out_881     ),
    .col_in_882              ( u2_col_out_882     ),
    .col_in_883              ( u2_col_out_883     ),
    .col_in_884              ( u2_col_out_884     ),
    .col_in_885              ( u2_col_out_885     ),
    .col_in_886              ( u2_col_out_886     ),
    .col_in_887              ( u2_col_out_887     ),
    .col_in_888              ( u2_col_out_888     ),
    .col_in_889              ( u2_col_out_889     ),
    .col_in_890              ( u2_col_out_890     ),
    .col_in_891              ( u2_col_out_891     ),
    .col_in_892              ( u2_col_out_892     ),
    .col_in_893              ( u2_col_out_893     ),
    .col_in_894              ( u2_col_out_894     ),
    .col_in_895              ( u2_col_out_895     ),
    .col_in_896              ( u2_col_out_896     ),
    .col_in_897              ( u2_col_out_897     ),
    .col_in_898              ( u2_col_out_898     ),
    .col_in_899              ( u2_col_out_899     ),
    .col_in_900              ( u2_col_out_900     ),
    .col_in_901              ( u2_col_out_901     ),
    .col_in_902              ( u2_col_out_902     ),
    .col_in_903              ( u2_col_out_903     ),
    .col_in_904              ( u2_col_out_904     ),
    .col_in_905              ( u2_col_out_905     ),
    .col_in_906              ( u2_col_out_906     ),
    .col_in_907              ( u2_col_out_907     ),
    .col_in_908              ( u2_col_out_908     ),
    .col_in_909              ( u2_col_out_909     ),
    .col_in_910              ( u2_col_out_910     ),
    .col_in_911              ( u2_col_out_911     ),
    .col_in_912              ( u2_col_out_912     ),
    .col_in_913              ( u2_col_out_913     ),
    .col_in_914              ( u2_col_out_914     ),
    .col_in_915              ( u2_col_out_915     ),
    .col_in_916              ( u2_col_out_916     ),
    .col_in_917              ( u2_col_out_917     ),
    .col_in_918              ( u2_col_out_918     ),
    .col_in_919              ( u2_col_out_919     ),
    .col_in_920              ( u2_col_out_920     ),
    .col_in_921              ( u2_col_out_921     ),
    .col_in_922              ( u2_col_out_922     ),
    .col_in_923              ( u2_col_out_923     ),
    .col_in_924              ( u2_col_out_924     ),
    .col_in_925              ( u2_col_out_925     ),
    .col_in_926              ( u2_col_out_926     ),
    .col_in_927              ( u2_col_out_927     ),
    .col_in_928              ( u2_col_out_928     ),
    .col_in_929              ( u2_col_out_929     ),
    .col_in_930              ( u2_col_out_930     ),
    .col_in_931              ( u2_col_out_931     ),
    .col_in_932              ( u2_col_out_932     ),
    .col_in_933              ( u2_col_out_933     ),
    .col_in_934              ( u2_col_out_934     ),
    .col_in_935              ( u2_col_out_935     ),
    .col_in_936              ( u2_col_out_936     ),
    .col_in_937              ( u2_col_out_937     ),
    .col_in_938              ( u2_col_out_938     ),
    .col_in_939              ( u2_col_out_939     ),
    .col_in_940              ( u2_col_out_940     ),
    .col_in_941              ( u2_col_out_941     ),
    .col_in_942              ( u2_col_out_942     ),
    .col_in_943              ( u2_col_out_943     ),
    .col_in_944              ( u2_col_out_944     ),
    .col_in_945              ( u2_col_out_945     ),
    .col_in_946              ( u2_col_out_946     ),
    .col_in_947              ( u2_col_out_947     ),
    .col_in_948              ( u2_col_out_948     ),
    .col_in_949              ( u2_col_out_949     ),
    .col_in_950              ( u2_col_out_950     ),
    .col_in_951              ( u2_col_out_951     ),
    .col_in_952              ( u2_col_out_952     ),
    .col_in_953              ( u2_col_out_953     ),
    .col_in_954              ( u2_col_out_954     ),
    .col_in_955              ( u2_col_out_955     ),
    .col_in_956              ( u2_col_out_956     ),
    .col_in_957              ( u2_col_out_957     ),
    .col_in_958              ( u2_col_out_958     ),
    .col_in_959              ( u2_col_out_959     ),
    .col_in_960              ( u2_col_out_960     ),
    .col_in_961              ( u2_col_out_961     ),
    .col_in_962              ( u2_col_out_962     ),
    .col_in_963              ( u2_col_out_963     ),
    .col_in_964              ( u2_col_out_964     ),
    .col_in_965              ( u2_col_out_965     ),
    .col_in_966              ( u2_col_out_966     ),
    .col_in_967              ( u2_col_out_967     ),
    .col_in_968              ( u2_col_out_968     ),
    .col_in_969              ( u2_col_out_969     ),
    .col_in_970              ( u2_col_out_970     ),
    .col_in_971              ( u2_col_out_971     ),
    .col_in_972              ( u2_col_out_972     ),
    .col_in_973              ( u2_col_out_973     ),
    .col_in_974              ( u2_col_out_974     ),
    .col_in_975              ( u2_col_out_975     ),
    .col_in_976              ( u2_col_out_976     ),
    .col_in_977              ( u2_col_out_977     ),
    .col_in_978              ( u2_col_out_978     ),
    .col_in_979              ( u2_col_out_979     ),
    .col_in_980              ( u2_col_out_980     ),
    .col_in_981              ( u2_col_out_981     ),
    .col_in_982              ( u2_col_out_982     ),
    .col_in_983              ( u2_col_out_983     ),
    .col_in_984              ( u2_col_out_984     ),
    .col_in_985              ( u2_col_out_985     ),
    .col_in_986              ( u2_col_out_986     ),
    .col_in_987              ( u2_col_out_987     ),
    .col_in_988              ( u2_col_out_988     ),
    .col_in_989              ( u2_col_out_989     ),
    .col_in_990              ( u2_col_out_990     ),
    .col_in_991              ( u2_col_out_991     ),
    .col_in_992              ( u2_col_out_992     ),
    .col_in_993              ( u2_col_out_993     ),
    .col_in_994              ( u2_col_out_994     ),
    .col_in_995              ( u2_col_out_995     ),
    .col_in_996              ( u2_col_out_996     ),
    .col_in_997              ( u2_col_out_997     ),
    .col_in_998              ( u2_col_out_998     ),
    .col_in_999              ( u2_col_out_999     ),
    .col_in_1000             ( u2_col_out_1000    ),
    .col_in_1001             ( u2_col_out_1001    ),
    .col_in_1002             ( u2_col_out_1002    ),
    .col_in_1003             ( u2_col_out_1003    ),
    .col_in_1004             ( u2_col_out_1004    ),
    .col_in_1005             ( u2_col_out_1005    ),
    .col_in_1006             ( u2_col_out_1006    ),
    .col_in_1007             ( u2_col_out_1007    ),
    .col_in_1008             ( u2_col_out_1008    ),
    .col_in_1009             ( u2_col_out_1009    ),
    .col_in_1010             ( u2_col_out_1010    ),
    .col_in_1011             ( u2_col_out_1011    ),
    .col_in_1012             ( u2_col_out_1012    ),
    .col_in_1013             ( u2_col_out_1013    ),
    .col_in_1014             ( u2_col_out_1014    ),
    .col_in_1015             ( u2_col_out_1015    ),
    .col_in_1016             ( u2_col_out_1016    ),
    .col_in_1017             ( u2_col_out_1017    ),
    .col_in_1018             ( u2_col_out_1018    ),
    .col_in_1019             ( u2_col_out_1019    ),
    .col_in_1020             ( u2_col_out_1020    ),
    .col_in_1021             ( u2_col_out_1021    ),
    .col_in_1022             ( u2_col_out_1022    ),
    .col_in_1023             ( u2_col_out_1023    ),
    .col_in_1024             ( u2_col_out_1024    ),
    .col_in_1025             ( u2_col_out_1025    ),
    .col_in_1026             ( u2_col_out_1026    ),
    .col_in_1027             ( u2_col_out_1027    ),
    .col_in_1028             ( u2_col_out_1028    ),
    .col_in_1029             ( u2_col_out_1029    ),
    .col_in_1030             ( u2_col_out_1030    ),
    .col_in_1031             ( u2_col_out_1031    ),
    .col_in_1032             ( u2_col_out_1032    ),


    .col_out_0               ( u3_col_out_0      ),
    .col_out_1               ( u3_col_out_1      ),
    .col_out_2               ( u3_col_out_2      ),
    .col_out_3               ( u3_col_out_3      ),
    .col_out_4               ( u3_col_out_4      ),
    .col_out_5               ( u3_col_out_5      ),
    .col_out_6               ( u3_col_out_6      ),
    .col_out_7               ( u3_col_out_7      ),
    .col_out_8               ( u3_col_out_8      ),
    .col_out_9               ( u3_col_out_9      ),
    .col_out_10              ( u3_col_out_10     ),
    .col_out_11              ( u3_col_out_11     ),
    .col_out_12              ( u3_col_out_12     ),
    .col_out_13              ( u3_col_out_13     ),
    .col_out_14              ( u3_col_out_14     ),
    .col_out_15              ( u3_col_out_15     ),
    .col_out_16              ( u3_col_out_16     ),
    .col_out_17              ( u3_col_out_17     ),
    .col_out_18              ( u3_col_out_18     ),
    .col_out_19              ( u3_col_out_19     ),
    .col_out_20              ( u3_col_out_20     ),
    .col_out_21              ( u3_col_out_21     ),
    .col_out_22              ( u3_col_out_22     ),
    .col_out_23              ( u3_col_out_23     ),
    .col_out_24              ( u3_col_out_24     ),
    .col_out_25              ( u3_col_out_25     ),
    .col_out_26              ( u3_col_out_26     ),
    .col_out_27              ( u3_col_out_27     ),
    .col_out_28              ( u3_col_out_28     ),
    .col_out_29              ( u3_col_out_29     ),
    .col_out_30              ( u3_col_out_30     ),
    .col_out_31              ( u3_col_out_31     ),
    .col_out_32              ( u3_col_out_32     ),
    .col_out_33              ( u3_col_out_33     ),
    .col_out_34              ( u3_col_out_34     ),
    .col_out_35              ( u3_col_out_35     ),
    .col_out_36              ( u3_col_out_36     ),
    .col_out_37              ( u3_col_out_37     ),
    .col_out_38              ( u3_col_out_38     ),
    .col_out_39              ( u3_col_out_39     ),
    .col_out_40              ( u3_col_out_40     ),
    .col_out_41              ( u3_col_out_41     ),
    .col_out_42              ( u3_col_out_42     ),
    .col_out_43              ( u3_col_out_43     ),
    .col_out_44              ( u3_col_out_44     ),
    .col_out_45              ( u3_col_out_45     ),
    .col_out_46              ( u3_col_out_46     ),
    .col_out_47              ( u3_col_out_47     ),
    .col_out_48              ( u3_col_out_48     ),
    .col_out_49              ( u3_col_out_49     ),
    .col_out_50              ( u3_col_out_50     ),
    .col_out_51              ( u3_col_out_51     ),
    .col_out_52              ( u3_col_out_52     ),
    .col_out_53              ( u3_col_out_53     ),
    .col_out_54              ( u3_col_out_54     ),
    .col_out_55              ( u3_col_out_55     ),
    .col_out_56              ( u3_col_out_56     ),
    .col_out_57              ( u3_col_out_57     ),
    .col_out_58              ( u3_col_out_58     ),
    .col_out_59              ( u3_col_out_59     ),
    .col_out_60              ( u3_col_out_60     ),
    .col_out_61              ( u3_col_out_61     ),
    .col_out_62              ( u3_col_out_62     ),
    .col_out_63              ( u3_col_out_63     ),
    .col_out_64              ( u3_col_out_64     ),
    .col_out_65              ( u3_col_out_65     ),
    .col_out_66              ( u3_col_out_66     ),
    .col_out_67              ( u3_col_out_67     ),
    .col_out_68              ( u3_col_out_68     ),
    .col_out_69              ( u3_col_out_69     ),
    .col_out_70              ( u3_col_out_70     ),
    .col_out_71              ( u3_col_out_71     ),
    .col_out_72              ( u3_col_out_72     ),
    .col_out_73              ( u3_col_out_73     ),
    .col_out_74              ( u3_col_out_74     ),
    .col_out_75              ( u3_col_out_75     ),
    .col_out_76              ( u3_col_out_76     ),
    .col_out_77              ( u3_col_out_77     ),
    .col_out_78              ( u3_col_out_78     ),
    .col_out_79              ( u3_col_out_79     ),
    .col_out_80              ( u3_col_out_80     ),
    .col_out_81              ( u3_col_out_81     ),
    .col_out_82              ( u3_col_out_82     ),
    .col_out_83              ( u3_col_out_83     ),
    .col_out_84              ( u3_col_out_84     ),
    .col_out_85              ( u3_col_out_85     ),
    .col_out_86              ( u3_col_out_86     ),
    .col_out_87              ( u3_col_out_87     ),
    .col_out_88              ( u3_col_out_88     ),
    .col_out_89              ( u3_col_out_89     ),
    .col_out_90              ( u3_col_out_90     ),
    .col_out_91              ( u3_col_out_91     ),
    .col_out_92              ( u3_col_out_92     ),
    .col_out_93              ( u3_col_out_93     ),
    .col_out_94              ( u3_col_out_94     ),
    .col_out_95              ( u3_col_out_95     ),
    .col_out_96              ( u3_col_out_96     ),
    .col_out_97              ( u3_col_out_97     ),
    .col_out_98              ( u3_col_out_98     ),
    .col_out_99              ( u3_col_out_99     ),
    .col_out_100             ( u3_col_out_100    ),
    .col_out_101             ( u3_col_out_101    ),
    .col_out_102             ( u3_col_out_102    ),
    .col_out_103             ( u3_col_out_103    ),
    .col_out_104             ( u3_col_out_104    ),
    .col_out_105             ( u3_col_out_105    ),
    .col_out_106             ( u3_col_out_106    ),
    .col_out_107             ( u3_col_out_107    ),
    .col_out_108             ( u3_col_out_108    ),
    .col_out_109             ( u3_col_out_109    ),
    .col_out_110             ( u3_col_out_110    ),
    .col_out_111             ( u3_col_out_111    ),
    .col_out_112             ( u3_col_out_112    ),
    .col_out_113             ( u3_col_out_113    ),
    .col_out_114             ( u3_col_out_114    ),
    .col_out_115             ( u3_col_out_115    ),
    .col_out_116             ( u3_col_out_116    ),
    .col_out_117             ( u3_col_out_117    ),
    .col_out_118             ( u3_col_out_118    ),
    .col_out_119             ( u3_col_out_119    ),
    .col_out_120             ( u3_col_out_120    ),
    .col_out_121             ( u3_col_out_121    ),
    .col_out_122             ( u3_col_out_122    ),
    .col_out_123             ( u3_col_out_123    ),
    .col_out_124             ( u3_col_out_124    ),
    .col_out_125             ( u3_col_out_125    ),
    .col_out_126             ( u3_col_out_126    ),
    .col_out_127             ( u3_col_out_127    ),
    .col_out_128             ( u3_col_out_128    ),
    .col_out_129             ( u3_col_out_129    ),
    .col_out_130             ( u3_col_out_130    ),
    .col_out_131             ( u3_col_out_131    ),
    .col_out_132             ( u3_col_out_132    ),
    .col_out_133             ( u3_col_out_133    ),
    .col_out_134             ( u3_col_out_134    ),
    .col_out_135             ( u3_col_out_135    ),
    .col_out_136             ( u3_col_out_136    ),
    .col_out_137             ( u3_col_out_137    ),
    .col_out_138             ( u3_col_out_138    ),
    .col_out_139             ( u3_col_out_139    ),
    .col_out_140             ( u3_col_out_140    ),
    .col_out_141             ( u3_col_out_141    ),
    .col_out_142             ( u3_col_out_142    ),
    .col_out_143             ( u3_col_out_143    ),
    .col_out_144             ( u3_col_out_144    ),
    .col_out_145             ( u3_col_out_145    ),
    .col_out_146             ( u3_col_out_146    ),
    .col_out_147             ( u3_col_out_147    ),
    .col_out_148             ( u3_col_out_148    ),
    .col_out_149             ( u3_col_out_149    ),
    .col_out_150             ( u3_col_out_150    ),
    .col_out_151             ( u3_col_out_151    ),
    .col_out_152             ( u3_col_out_152    ),
    .col_out_153             ( u3_col_out_153    ),
    .col_out_154             ( u3_col_out_154    ),
    .col_out_155             ( u3_col_out_155    ),
    .col_out_156             ( u3_col_out_156    ),
    .col_out_157             ( u3_col_out_157    ),
    .col_out_158             ( u3_col_out_158    ),
    .col_out_159             ( u3_col_out_159    ),
    .col_out_160             ( u3_col_out_160    ),
    .col_out_161             ( u3_col_out_161    ),
    .col_out_162             ( u3_col_out_162    ),
    .col_out_163             ( u3_col_out_163    ),
    .col_out_164             ( u3_col_out_164    ),
    .col_out_165             ( u3_col_out_165    ),
    .col_out_166             ( u3_col_out_166    ),
    .col_out_167             ( u3_col_out_167    ),
    .col_out_168             ( u3_col_out_168    ),
    .col_out_169             ( u3_col_out_169    ),
    .col_out_170             ( u3_col_out_170    ),
    .col_out_171             ( u3_col_out_171    ),
    .col_out_172             ( u3_col_out_172    ),
    .col_out_173             ( u3_col_out_173    ),
    .col_out_174             ( u3_col_out_174    ),
    .col_out_175             ( u3_col_out_175    ),
    .col_out_176             ( u3_col_out_176    ),
    .col_out_177             ( u3_col_out_177    ),
    .col_out_178             ( u3_col_out_178    ),
    .col_out_179             ( u3_col_out_179    ),
    .col_out_180             ( u3_col_out_180    ),
    .col_out_181             ( u3_col_out_181    ),
    .col_out_182             ( u3_col_out_182    ),
    .col_out_183             ( u3_col_out_183    ),
    .col_out_184             ( u3_col_out_184    ),
    .col_out_185             ( u3_col_out_185    ),
    .col_out_186             ( u3_col_out_186    ),
    .col_out_187             ( u3_col_out_187    ),
    .col_out_188             ( u3_col_out_188    ),
    .col_out_189             ( u3_col_out_189    ),
    .col_out_190             ( u3_col_out_190    ),
    .col_out_191             ( u3_col_out_191    ),
    .col_out_192             ( u3_col_out_192    ),
    .col_out_193             ( u3_col_out_193    ),
    .col_out_194             ( u3_col_out_194    ),
    .col_out_195             ( u3_col_out_195    ),
    .col_out_196             ( u3_col_out_196    ),
    .col_out_197             ( u3_col_out_197    ),
    .col_out_198             ( u3_col_out_198    ),
    .col_out_199             ( u3_col_out_199    ),
    .col_out_200             ( u3_col_out_200    ),
    .col_out_201             ( u3_col_out_201    ),
    .col_out_202             ( u3_col_out_202    ),
    .col_out_203             ( u3_col_out_203    ),
    .col_out_204             ( u3_col_out_204    ),
    .col_out_205             ( u3_col_out_205    ),
    .col_out_206             ( u3_col_out_206    ),
    .col_out_207             ( u3_col_out_207    ),
    .col_out_208             ( u3_col_out_208    ),
    .col_out_209             ( u3_col_out_209    ),
    .col_out_210             ( u3_col_out_210    ),
    .col_out_211             ( u3_col_out_211    ),
    .col_out_212             ( u3_col_out_212    ),
    .col_out_213             ( u3_col_out_213    ),
    .col_out_214             ( u3_col_out_214    ),
    .col_out_215             ( u3_col_out_215    ),
    .col_out_216             ( u3_col_out_216    ),
    .col_out_217             ( u3_col_out_217    ),
    .col_out_218             ( u3_col_out_218    ),
    .col_out_219             ( u3_col_out_219    ),
    .col_out_220             ( u3_col_out_220    ),
    .col_out_221             ( u3_col_out_221    ),
    .col_out_222             ( u3_col_out_222    ),
    .col_out_223             ( u3_col_out_223    ),
    .col_out_224             ( u3_col_out_224    ),
    .col_out_225             ( u3_col_out_225    ),
    .col_out_226             ( u3_col_out_226    ),
    .col_out_227             ( u3_col_out_227    ),
    .col_out_228             ( u3_col_out_228    ),
    .col_out_229             ( u3_col_out_229    ),
    .col_out_230             ( u3_col_out_230    ),
    .col_out_231             ( u3_col_out_231    ),
    .col_out_232             ( u3_col_out_232    ),
    .col_out_233             ( u3_col_out_233    ),
    .col_out_234             ( u3_col_out_234    ),
    .col_out_235             ( u3_col_out_235    ),
    .col_out_236             ( u3_col_out_236    ),
    .col_out_237             ( u3_col_out_237    ),
    .col_out_238             ( u3_col_out_238    ),
    .col_out_239             ( u3_col_out_239    ),
    .col_out_240             ( u3_col_out_240    ),
    .col_out_241             ( u3_col_out_241    ),
    .col_out_242             ( u3_col_out_242    ),
    .col_out_243             ( u3_col_out_243    ),
    .col_out_244             ( u3_col_out_244    ),
    .col_out_245             ( u3_col_out_245    ),
    .col_out_246             ( u3_col_out_246    ),
    .col_out_247             ( u3_col_out_247    ),
    .col_out_248             ( u3_col_out_248    ),
    .col_out_249             ( u3_col_out_249    ),
    .col_out_250             ( u3_col_out_250    ),
    .col_out_251             ( u3_col_out_251    ),
    .col_out_252             ( u3_col_out_252    ),
    .col_out_253             ( u3_col_out_253    ),
    .col_out_254             ( u3_col_out_254    ),
    .col_out_255             ( u3_col_out_255    ),
    .col_out_256             ( u3_col_out_256    ),
    .col_out_257             ( u3_col_out_257    ),
    .col_out_258             ( u3_col_out_258    ),
    .col_out_259             ( u3_col_out_259    ),
    .col_out_260             ( u3_col_out_260    ),
    .col_out_261             ( u3_col_out_261    ),
    .col_out_262             ( u3_col_out_262    ),
    .col_out_263             ( u3_col_out_263    ),
    .col_out_264             ( u3_col_out_264    ),
    .col_out_265             ( u3_col_out_265    ),
    .col_out_266             ( u3_col_out_266    ),
    .col_out_267             ( u3_col_out_267    ),
    .col_out_268             ( u3_col_out_268    ),
    .col_out_269             ( u3_col_out_269    ),
    .col_out_270             ( u3_col_out_270    ),
    .col_out_271             ( u3_col_out_271    ),
    .col_out_272             ( u3_col_out_272    ),
    .col_out_273             ( u3_col_out_273    ),
    .col_out_274             ( u3_col_out_274    ),
    .col_out_275             ( u3_col_out_275    ),
    .col_out_276             ( u3_col_out_276    ),
    .col_out_277             ( u3_col_out_277    ),
    .col_out_278             ( u3_col_out_278    ),
    .col_out_279             ( u3_col_out_279    ),
    .col_out_280             ( u3_col_out_280    ),
    .col_out_281             ( u3_col_out_281    ),
    .col_out_282             ( u3_col_out_282    ),
    .col_out_283             ( u3_col_out_283    ),
    .col_out_284             ( u3_col_out_284    ),
    .col_out_285             ( u3_col_out_285    ),
    .col_out_286             ( u3_col_out_286    ),
    .col_out_287             ( u3_col_out_287    ),
    .col_out_288             ( u3_col_out_288    ),
    .col_out_289             ( u3_col_out_289    ),
    .col_out_290             ( u3_col_out_290    ),
    .col_out_291             ( u3_col_out_291    ),
    .col_out_292             ( u3_col_out_292    ),
    .col_out_293             ( u3_col_out_293    ),
    .col_out_294             ( u3_col_out_294    ),
    .col_out_295             ( u3_col_out_295    ),
    .col_out_296             ( u3_col_out_296    ),
    .col_out_297             ( u3_col_out_297    ),
    .col_out_298             ( u3_col_out_298    ),
    .col_out_299             ( u3_col_out_299    ),
    .col_out_300             ( u3_col_out_300    ),
    .col_out_301             ( u3_col_out_301    ),
    .col_out_302             ( u3_col_out_302    ),
    .col_out_303             ( u3_col_out_303    ),
    .col_out_304             ( u3_col_out_304    ),
    .col_out_305             ( u3_col_out_305    ),
    .col_out_306             ( u3_col_out_306    ),
    .col_out_307             ( u3_col_out_307    ),
    .col_out_308             ( u3_col_out_308    ),
    .col_out_309             ( u3_col_out_309    ),
    .col_out_310             ( u3_col_out_310    ),
    .col_out_311             ( u3_col_out_311    ),
    .col_out_312             ( u3_col_out_312    ),
    .col_out_313             ( u3_col_out_313    ),
    .col_out_314             ( u3_col_out_314    ),
    .col_out_315             ( u3_col_out_315    ),
    .col_out_316             ( u3_col_out_316    ),
    .col_out_317             ( u3_col_out_317    ),
    .col_out_318             ( u3_col_out_318    ),
    .col_out_319             ( u3_col_out_319    ),
    .col_out_320             ( u3_col_out_320    ),
    .col_out_321             ( u3_col_out_321    ),
    .col_out_322             ( u3_col_out_322    ),
    .col_out_323             ( u3_col_out_323    ),
    .col_out_324             ( u3_col_out_324    ),
    .col_out_325             ( u3_col_out_325    ),
    .col_out_326             ( u3_col_out_326    ),
    .col_out_327             ( u3_col_out_327    ),
    .col_out_328             ( u3_col_out_328    ),
    .col_out_329             ( u3_col_out_329    ),
    .col_out_330             ( u3_col_out_330    ),
    .col_out_331             ( u3_col_out_331    ),
    .col_out_332             ( u3_col_out_332    ),
    .col_out_333             ( u3_col_out_333    ),
    .col_out_334             ( u3_col_out_334    ),
    .col_out_335             ( u3_col_out_335    ),
    .col_out_336             ( u3_col_out_336    ),
    .col_out_337             ( u3_col_out_337    ),
    .col_out_338             ( u3_col_out_338    ),
    .col_out_339             ( u3_col_out_339    ),
    .col_out_340             ( u3_col_out_340    ),
    .col_out_341             ( u3_col_out_341    ),
    .col_out_342             ( u3_col_out_342    ),
    .col_out_343             ( u3_col_out_343    ),
    .col_out_344             ( u3_col_out_344    ),
    .col_out_345             ( u3_col_out_345    ),
    .col_out_346             ( u3_col_out_346    ),
    .col_out_347             ( u3_col_out_347    ),
    .col_out_348             ( u3_col_out_348    ),
    .col_out_349             ( u3_col_out_349    ),
    .col_out_350             ( u3_col_out_350    ),
    .col_out_351             ( u3_col_out_351    ),
    .col_out_352             ( u3_col_out_352    ),
    .col_out_353             ( u3_col_out_353    ),
    .col_out_354             ( u3_col_out_354    ),
    .col_out_355             ( u3_col_out_355    ),
    .col_out_356             ( u3_col_out_356    ),
    .col_out_357             ( u3_col_out_357    ),
    .col_out_358             ( u3_col_out_358    ),
    .col_out_359             ( u3_col_out_359    ),
    .col_out_360             ( u3_col_out_360    ),
    .col_out_361             ( u3_col_out_361    ),
    .col_out_362             ( u3_col_out_362    ),
    .col_out_363             ( u3_col_out_363    ),
    .col_out_364             ( u3_col_out_364    ),
    .col_out_365             ( u3_col_out_365    ),
    .col_out_366             ( u3_col_out_366    ),
    .col_out_367             ( u3_col_out_367    ),
    .col_out_368             ( u3_col_out_368    ),
    .col_out_369             ( u3_col_out_369    ),
    .col_out_370             ( u3_col_out_370    ),
    .col_out_371             ( u3_col_out_371    ),
    .col_out_372             ( u3_col_out_372    ),
    .col_out_373             ( u3_col_out_373    ),
    .col_out_374             ( u3_col_out_374    ),
    .col_out_375             ( u3_col_out_375    ),
    .col_out_376             ( u3_col_out_376    ),
    .col_out_377             ( u3_col_out_377    ),
    .col_out_378             ( u3_col_out_378    ),
    .col_out_379             ( u3_col_out_379    ),
    .col_out_380             ( u3_col_out_380    ),
    .col_out_381             ( u3_col_out_381    ),
    .col_out_382             ( u3_col_out_382    ),
    .col_out_383             ( u3_col_out_383    ),
    .col_out_384             ( u3_col_out_384    ),
    .col_out_385             ( u3_col_out_385    ),
    .col_out_386             ( u3_col_out_386    ),
    .col_out_387             ( u3_col_out_387    ),
    .col_out_388             ( u3_col_out_388    ),
    .col_out_389             ( u3_col_out_389    ),
    .col_out_390             ( u3_col_out_390    ),
    .col_out_391             ( u3_col_out_391    ),
    .col_out_392             ( u3_col_out_392    ),
    .col_out_393             ( u3_col_out_393    ),
    .col_out_394             ( u3_col_out_394    ),
    .col_out_395             ( u3_col_out_395    ),
    .col_out_396             ( u3_col_out_396    ),
    .col_out_397             ( u3_col_out_397    ),
    .col_out_398             ( u3_col_out_398    ),
    .col_out_399             ( u3_col_out_399    ),
    .col_out_400             ( u3_col_out_400    ),
    .col_out_401             ( u3_col_out_401    ),
    .col_out_402             ( u3_col_out_402    ),
    .col_out_403             ( u3_col_out_403    ),
    .col_out_404             ( u3_col_out_404    ),
    .col_out_405             ( u3_col_out_405    ),
    .col_out_406             ( u3_col_out_406    ),
    .col_out_407             ( u3_col_out_407    ),
    .col_out_408             ( u3_col_out_408    ),
    .col_out_409             ( u3_col_out_409    ),
    .col_out_410             ( u3_col_out_410    ),
    .col_out_411             ( u3_col_out_411    ),
    .col_out_412             ( u3_col_out_412    ),
    .col_out_413             ( u3_col_out_413    ),
    .col_out_414             ( u3_col_out_414    ),
    .col_out_415             ( u3_col_out_415    ),
    .col_out_416             ( u3_col_out_416    ),
    .col_out_417             ( u3_col_out_417    ),
    .col_out_418             ( u3_col_out_418    ),
    .col_out_419             ( u3_col_out_419    ),
    .col_out_420             ( u3_col_out_420    ),
    .col_out_421             ( u3_col_out_421    ),
    .col_out_422             ( u3_col_out_422    ),
    .col_out_423             ( u3_col_out_423    ),
    .col_out_424             ( u3_col_out_424    ),
    .col_out_425             ( u3_col_out_425    ),
    .col_out_426             ( u3_col_out_426    ),
    .col_out_427             ( u3_col_out_427    ),
    .col_out_428             ( u3_col_out_428    ),
    .col_out_429             ( u3_col_out_429    ),
    .col_out_430             ( u3_col_out_430    ),
    .col_out_431             ( u3_col_out_431    ),
    .col_out_432             ( u3_col_out_432    ),
    .col_out_433             ( u3_col_out_433    ),
    .col_out_434             ( u3_col_out_434    ),
    .col_out_435             ( u3_col_out_435    ),
    .col_out_436             ( u3_col_out_436    ),
    .col_out_437             ( u3_col_out_437    ),
    .col_out_438             ( u3_col_out_438    ),
    .col_out_439             ( u3_col_out_439    ),
    .col_out_440             ( u3_col_out_440    ),
    .col_out_441             ( u3_col_out_441    ),
    .col_out_442             ( u3_col_out_442    ),
    .col_out_443             ( u3_col_out_443    ),
    .col_out_444             ( u3_col_out_444    ),
    .col_out_445             ( u3_col_out_445    ),
    .col_out_446             ( u3_col_out_446    ),
    .col_out_447             ( u3_col_out_447    ),
    .col_out_448             ( u3_col_out_448    ),
    .col_out_449             ( u3_col_out_449    ),
    .col_out_450             ( u3_col_out_450    ),
    .col_out_451             ( u3_col_out_451    ),
    .col_out_452             ( u3_col_out_452    ),
    .col_out_453             ( u3_col_out_453    ),
    .col_out_454             ( u3_col_out_454    ),
    .col_out_455             ( u3_col_out_455    ),
    .col_out_456             ( u3_col_out_456    ),
    .col_out_457             ( u3_col_out_457    ),
    .col_out_458             ( u3_col_out_458    ),
    .col_out_459             ( u3_col_out_459    ),
    .col_out_460             ( u3_col_out_460    ),
    .col_out_461             ( u3_col_out_461    ),
    .col_out_462             ( u3_col_out_462    ),
    .col_out_463             ( u3_col_out_463    ),
    .col_out_464             ( u3_col_out_464    ),
    .col_out_465             ( u3_col_out_465    ),
    .col_out_466             ( u3_col_out_466    ),
    .col_out_467             ( u3_col_out_467    ),
    .col_out_468             ( u3_col_out_468    ),
    .col_out_469             ( u3_col_out_469    ),
    .col_out_470             ( u3_col_out_470    ),
    .col_out_471             ( u3_col_out_471    ),
    .col_out_472             ( u3_col_out_472    ),
    .col_out_473             ( u3_col_out_473    ),
    .col_out_474             ( u3_col_out_474    ),
    .col_out_475             ( u3_col_out_475    ),
    .col_out_476             ( u3_col_out_476    ),
    .col_out_477             ( u3_col_out_477    ),
    .col_out_478             ( u3_col_out_478    ),
    .col_out_479             ( u3_col_out_479    ),
    .col_out_480             ( u3_col_out_480    ),
    .col_out_481             ( u3_col_out_481    ),
    .col_out_482             ( u3_col_out_482    ),
    .col_out_483             ( u3_col_out_483    ),
    .col_out_484             ( u3_col_out_484    ),
    .col_out_485             ( u3_col_out_485    ),
    .col_out_486             ( u3_col_out_486    ),
    .col_out_487             ( u3_col_out_487    ),
    .col_out_488             ( u3_col_out_488    ),
    .col_out_489             ( u3_col_out_489    ),
    .col_out_490             ( u3_col_out_490    ),
    .col_out_491             ( u3_col_out_491    ),
    .col_out_492             ( u3_col_out_492    ),
    .col_out_493             ( u3_col_out_493    ),
    .col_out_494             ( u3_col_out_494    ),
    .col_out_495             ( u3_col_out_495    ),
    .col_out_496             ( u3_col_out_496    ),
    .col_out_497             ( u3_col_out_497    ),
    .col_out_498             ( u3_col_out_498    ),
    .col_out_499             ( u3_col_out_499    ),
    .col_out_500             ( u3_col_out_500    ),
    .col_out_501             ( u3_col_out_501    ),
    .col_out_502             ( u3_col_out_502    ),
    .col_out_503             ( u3_col_out_503    ),
    .col_out_504             ( u3_col_out_504    ),
    .col_out_505             ( u3_col_out_505    ),
    .col_out_506             ( u3_col_out_506    ),
    .col_out_507             ( u3_col_out_507    ),
    .col_out_508             ( u3_col_out_508    ),
    .col_out_509             ( u3_col_out_509    ),
    .col_out_510             ( u3_col_out_510    ),
    .col_out_511             ( u3_col_out_511    ),
    .col_out_512             ( u3_col_out_512    ),
    .col_out_513             ( u3_col_out_513    ),
    .col_out_514             ( u3_col_out_514    ),
    .col_out_515             ( u3_col_out_515    ),
    .col_out_516             ( u3_col_out_516    ),
    .col_out_517             ( u3_col_out_517    ),
    .col_out_518             ( u3_col_out_518    ),
    .col_out_519             ( u3_col_out_519    ),
    .col_out_520             ( u3_col_out_520    ),
    .col_out_521             ( u3_col_out_521    ),
    .col_out_522             ( u3_col_out_522    ),
    .col_out_523             ( u3_col_out_523    ),
    .col_out_524             ( u3_col_out_524    ),
    .col_out_525             ( u3_col_out_525    ),
    .col_out_526             ( u3_col_out_526    ),
    .col_out_527             ( u3_col_out_527    ),
    .col_out_528             ( u3_col_out_528    ),
    .col_out_529             ( u3_col_out_529    ),
    .col_out_530             ( u3_col_out_530    ),
    .col_out_531             ( u3_col_out_531    ),
    .col_out_532             ( u3_col_out_532    ),
    .col_out_533             ( u3_col_out_533    ),
    .col_out_534             ( u3_col_out_534    ),
    .col_out_535             ( u3_col_out_535    ),
    .col_out_536             ( u3_col_out_536    ),
    .col_out_537             ( u3_col_out_537    ),
    .col_out_538             ( u3_col_out_538    ),
    .col_out_539             ( u3_col_out_539    ),
    .col_out_540             ( u3_col_out_540    ),
    .col_out_541             ( u3_col_out_541    ),
    .col_out_542             ( u3_col_out_542    ),
    .col_out_543             ( u3_col_out_543    ),
    .col_out_544             ( u3_col_out_544    ),
    .col_out_545             ( u3_col_out_545    ),
    .col_out_546             ( u3_col_out_546    ),
    .col_out_547             ( u3_col_out_547    ),
    .col_out_548             ( u3_col_out_548    ),
    .col_out_549             ( u3_col_out_549    ),
    .col_out_550             ( u3_col_out_550    ),
    .col_out_551             ( u3_col_out_551    ),
    .col_out_552             ( u3_col_out_552    ),
    .col_out_553             ( u3_col_out_553    ),
    .col_out_554             ( u3_col_out_554    ),
    .col_out_555             ( u3_col_out_555    ),
    .col_out_556             ( u3_col_out_556    ),
    .col_out_557             ( u3_col_out_557    ),
    .col_out_558             ( u3_col_out_558    ),
    .col_out_559             ( u3_col_out_559    ),
    .col_out_560             ( u3_col_out_560    ),
    .col_out_561             ( u3_col_out_561    ),
    .col_out_562             ( u3_col_out_562    ),
    .col_out_563             ( u3_col_out_563    ),
    .col_out_564             ( u3_col_out_564    ),
    .col_out_565             ( u3_col_out_565    ),
    .col_out_566             ( u3_col_out_566    ),
    .col_out_567             ( u3_col_out_567    ),
    .col_out_568             ( u3_col_out_568    ),
    .col_out_569             ( u3_col_out_569    ),
    .col_out_570             ( u3_col_out_570    ),
    .col_out_571             ( u3_col_out_571    ),
    .col_out_572             ( u3_col_out_572    ),
    .col_out_573             ( u3_col_out_573    ),
    .col_out_574             ( u3_col_out_574    ),
    .col_out_575             ( u3_col_out_575    ),
    .col_out_576             ( u3_col_out_576    ),
    .col_out_577             ( u3_col_out_577    ),
    .col_out_578             ( u3_col_out_578    ),
    .col_out_579             ( u3_col_out_579    ),
    .col_out_580             ( u3_col_out_580    ),
    .col_out_581             ( u3_col_out_581    ),
    .col_out_582             ( u3_col_out_582    ),
    .col_out_583             ( u3_col_out_583    ),
    .col_out_584             ( u3_col_out_584    ),
    .col_out_585             ( u3_col_out_585    ),
    .col_out_586             ( u3_col_out_586    ),
    .col_out_587             ( u3_col_out_587    ),
    .col_out_588             ( u3_col_out_588    ),
    .col_out_589             ( u3_col_out_589    ),
    .col_out_590             ( u3_col_out_590    ),
    .col_out_591             ( u3_col_out_591    ),
    .col_out_592             ( u3_col_out_592    ),
    .col_out_593             ( u3_col_out_593    ),
    .col_out_594             ( u3_col_out_594    ),
    .col_out_595             ( u3_col_out_595    ),
    .col_out_596             ( u3_col_out_596    ),
    .col_out_597             ( u3_col_out_597    ),
    .col_out_598             ( u3_col_out_598    ),
    .col_out_599             ( u3_col_out_599    ),
    .col_out_600             ( u3_col_out_600    ),
    .col_out_601             ( u3_col_out_601    ),
    .col_out_602             ( u3_col_out_602    ),
    .col_out_603             ( u3_col_out_603    ),
    .col_out_604             ( u3_col_out_604    ),
    .col_out_605             ( u3_col_out_605    ),
    .col_out_606             ( u3_col_out_606    ),
    .col_out_607             ( u3_col_out_607    ),
    .col_out_608             ( u3_col_out_608    ),
    .col_out_609             ( u3_col_out_609    ),
    .col_out_610             ( u3_col_out_610    ),
    .col_out_611             ( u3_col_out_611    ),
    .col_out_612             ( u3_col_out_612    ),
    .col_out_613             ( u3_col_out_613    ),
    .col_out_614             ( u3_col_out_614    ),
    .col_out_615             ( u3_col_out_615    ),
    .col_out_616             ( u3_col_out_616    ),
    .col_out_617             ( u3_col_out_617    ),
    .col_out_618             ( u3_col_out_618    ),
    .col_out_619             ( u3_col_out_619    ),
    .col_out_620             ( u3_col_out_620    ),
    .col_out_621             ( u3_col_out_621    ),
    .col_out_622             ( u3_col_out_622    ),
    .col_out_623             ( u3_col_out_623    ),
    .col_out_624             ( u3_col_out_624    ),
    .col_out_625             ( u3_col_out_625    ),
    .col_out_626             ( u3_col_out_626    ),
    .col_out_627             ( u3_col_out_627    ),
    .col_out_628             ( u3_col_out_628    ),
    .col_out_629             ( u3_col_out_629    ),
    .col_out_630             ( u3_col_out_630    ),
    .col_out_631             ( u3_col_out_631    ),
    .col_out_632             ( u3_col_out_632    ),
    .col_out_633             ( u3_col_out_633    ),
    .col_out_634             ( u3_col_out_634    ),
    .col_out_635             ( u3_col_out_635    ),
    .col_out_636             ( u3_col_out_636    ),
    .col_out_637             ( u3_col_out_637    ),
    .col_out_638             ( u3_col_out_638    ),
    .col_out_639             ( u3_col_out_639    ),
    .col_out_640             ( u3_col_out_640    ),
    .col_out_641             ( u3_col_out_641    ),
    .col_out_642             ( u3_col_out_642    ),
    .col_out_643             ( u3_col_out_643    ),
    .col_out_644             ( u3_col_out_644    ),
    .col_out_645             ( u3_col_out_645    ),
    .col_out_646             ( u3_col_out_646    ),
    .col_out_647             ( u3_col_out_647    ),
    .col_out_648             ( u3_col_out_648    ),
    .col_out_649             ( u3_col_out_649    ),
    .col_out_650             ( u3_col_out_650    ),
    .col_out_651             ( u3_col_out_651    ),
    .col_out_652             ( u3_col_out_652    ),
    .col_out_653             ( u3_col_out_653    ),
    .col_out_654             ( u3_col_out_654    ),
    .col_out_655             ( u3_col_out_655    ),
    .col_out_656             ( u3_col_out_656    ),
    .col_out_657             ( u3_col_out_657    ),
    .col_out_658             ( u3_col_out_658    ),
    .col_out_659             ( u3_col_out_659    ),
    .col_out_660             ( u3_col_out_660    ),
    .col_out_661             ( u3_col_out_661    ),
    .col_out_662             ( u3_col_out_662    ),
    .col_out_663             ( u3_col_out_663    ),
    .col_out_664             ( u3_col_out_664    ),
    .col_out_665             ( u3_col_out_665    ),
    .col_out_666             ( u3_col_out_666    ),
    .col_out_667             ( u3_col_out_667    ),
    .col_out_668             ( u3_col_out_668    ),
    .col_out_669             ( u3_col_out_669    ),
    .col_out_670             ( u3_col_out_670    ),
    .col_out_671             ( u3_col_out_671    ),
    .col_out_672             ( u3_col_out_672    ),
    .col_out_673             ( u3_col_out_673    ),
    .col_out_674             ( u3_col_out_674    ),
    .col_out_675             ( u3_col_out_675    ),
    .col_out_676             ( u3_col_out_676    ),
    .col_out_677             ( u3_col_out_677    ),
    .col_out_678             ( u3_col_out_678    ),
    .col_out_679             ( u3_col_out_679    ),
    .col_out_680             ( u3_col_out_680    ),
    .col_out_681             ( u3_col_out_681    ),
    .col_out_682             ( u3_col_out_682    ),
    .col_out_683             ( u3_col_out_683    ),
    .col_out_684             ( u3_col_out_684    ),
    .col_out_685             ( u3_col_out_685    ),
    .col_out_686             ( u3_col_out_686    ),
    .col_out_687             ( u3_col_out_687    ),
    .col_out_688             ( u3_col_out_688    ),
    .col_out_689             ( u3_col_out_689    ),
    .col_out_690             ( u3_col_out_690    ),
    .col_out_691             ( u3_col_out_691    ),
    .col_out_692             ( u3_col_out_692    ),
    .col_out_693             ( u3_col_out_693    ),
    .col_out_694             ( u3_col_out_694    ),
    .col_out_695             ( u3_col_out_695    ),
    .col_out_696             ( u3_col_out_696    ),
    .col_out_697             ( u3_col_out_697    ),
    .col_out_698             ( u3_col_out_698    ),
    .col_out_699             ( u3_col_out_699    ),
    .col_out_700             ( u3_col_out_700    ),
    .col_out_701             ( u3_col_out_701    ),
    .col_out_702             ( u3_col_out_702    ),
    .col_out_703             ( u3_col_out_703    ),
    .col_out_704             ( u3_col_out_704    ),
    .col_out_705             ( u3_col_out_705    ),
    .col_out_706             ( u3_col_out_706    ),
    .col_out_707             ( u3_col_out_707    ),
    .col_out_708             ( u3_col_out_708    ),
    .col_out_709             ( u3_col_out_709    ),
    .col_out_710             ( u3_col_out_710    ),
    .col_out_711             ( u3_col_out_711    ),
    .col_out_712             ( u3_col_out_712    ),
    .col_out_713             ( u3_col_out_713    ),
    .col_out_714             ( u3_col_out_714    ),
    .col_out_715             ( u3_col_out_715    ),
    .col_out_716             ( u3_col_out_716    ),
    .col_out_717             ( u3_col_out_717    ),
    .col_out_718             ( u3_col_out_718    ),
    .col_out_719             ( u3_col_out_719    ),
    .col_out_720             ( u3_col_out_720    ),
    .col_out_721             ( u3_col_out_721    ),
    .col_out_722             ( u3_col_out_722    ),
    .col_out_723             ( u3_col_out_723    ),
    .col_out_724             ( u3_col_out_724    ),
    .col_out_725             ( u3_col_out_725    ),
    .col_out_726             ( u3_col_out_726    ),
    .col_out_727             ( u3_col_out_727    ),
    .col_out_728             ( u3_col_out_728    ),
    .col_out_729             ( u3_col_out_729    ),
    .col_out_730             ( u3_col_out_730    ),
    .col_out_731             ( u3_col_out_731    ),
    .col_out_732             ( u3_col_out_732    ),
    .col_out_733             ( u3_col_out_733    ),
    .col_out_734             ( u3_col_out_734    ),
    .col_out_735             ( u3_col_out_735    ),
    .col_out_736             ( u3_col_out_736    ),
    .col_out_737             ( u3_col_out_737    ),
    .col_out_738             ( u3_col_out_738    ),
    .col_out_739             ( u3_col_out_739    ),
    .col_out_740             ( u3_col_out_740    ),
    .col_out_741             ( u3_col_out_741    ),
    .col_out_742             ( u3_col_out_742    ),
    .col_out_743             ( u3_col_out_743    ),
    .col_out_744             ( u3_col_out_744    ),
    .col_out_745             ( u3_col_out_745    ),
    .col_out_746             ( u3_col_out_746    ),
    .col_out_747             ( u3_col_out_747    ),
    .col_out_748             ( u3_col_out_748    ),
    .col_out_749             ( u3_col_out_749    ),
    .col_out_750             ( u3_col_out_750    ),
    .col_out_751             ( u3_col_out_751    ),
    .col_out_752             ( u3_col_out_752    ),
    .col_out_753             ( u3_col_out_753    ),
    .col_out_754             ( u3_col_out_754    ),
    .col_out_755             ( u3_col_out_755    ),
    .col_out_756             ( u3_col_out_756    ),
    .col_out_757             ( u3_col_out_757    ),
    .col_out_758             ( u3_col_out_758    ),
    .col_out_759             ( u3_col_out_759    ),
    .col_out_760             ( u3_col_out_760    ),
    .col_out_761             ( u3_col_out_761    ),
    .col_out_762             ( u3_col_out_762    ),
    .col_out_763             ( u3_col_out_763    ),
    .col_out_764             ( u3_col_out_764    ),
    .col_out_765             ( u3_col_out_765    ),
    .col_out_766             ( u3_col_out_766    ),
    .col_out_767             ( u3_col_out_767    ),
    .col_out_768             ( u3_col_out_768    ),
    .col_out_769             ( u3_col_out_769    ),
    .col_out_770             ( u3_col_out_770    ),
    .col_out_771             ( u3_col_out_771    ),
    .col_out_772             ( u3_col_out_772    ),
    .col_out_773             ( u3_col_out_773    ),
    .col_out_774             ( u3_col_out_774    ),
    .col_out_775             ( u3_col_out_775    ),
    .col_out_776             ( u3_col_out_776    ),
    .col_out_777             ( u3_col_out_777    ),
    .col_out_778             ( u3_col_out_778    ),
    .col_out_779             ( u3_col_out_779    ),
    .col_out_780             ( u3_col_out_780    ),
    .col_out_781             ( u3_col_out_781    ),
    .col_out_782             ( u3_col_out_782    ),
    .col_out_783             ( u3_col_out_783    ),
    .col_out_784             ( u3_col_out_784    ),
    .col_out_785             ( u3_col_out_785    ),
    .col_out_786             ( u3_col_out_786    ),
    .col_out_787             ( u3_col_out_787    ),
    .col_out_788             ( u3_col_out_788    ),
    .col_out_789             ( u3_col_out_789    ),
    .col_out_790             ( u3_col_out_790    ),
    .col_out_791             ( u3_col_out_791    ),
    .col_out_792             ( u3_col_out_792    ),
    .col_out_793             ( u3_col_out_793    ),
    .col_out_794             ( u3_col_out_794    ),
    .col_out_795             ( u3_col_out_795    ),
    .col_out_796             ( u3_col_out_796    ),
    .col_out_797             ( u3_col_out_797    ),
    .col_out_798             ( u3_col_out_798    ),
    .col_out_799             ( u3_col_out_799    ),
    .col_out_800             ( u3_col_out_800    ),
    .col_out_801             ( u3_col_out_801    ),
    .col_out_802             ( u3_col_out_802    ),
    .col_out_803             ( u3_col_out_803    ),
    .col_out_804             ( u3_col_out_804    ),
    .col_out_805             ( u3_col_out_805    ),
    .col_out_806             ( u3_col_out_806    ),
    .col_out_807             ( u3_col_out_807    ),
    .col_out_808             ( u3_col_out_808    ),
    .col_out_809             ( u3_col_out_809    ),
    .col_out_810             ( u3_col_out_810    ),
    .col_out_811             ( u3_col_out_811    ),
    .col_out_812             ( u3_col_out_812    ),
    .col_out_813             ( u3_col_out_813    ),
    .col_out_814             ( u3_col_out_814    ),
    .col_out_815             ( u3_col_out_815    ),
    .col_out_816             ( u3_col_out_816    ),
    .col_out_817             ( u3_col_out_817    ),
    .col_out_818             ( u3_col_out_818    ),
    .col_out_819             ( u3_col_out_819    ),
    .col_out_820             ( u3_col_out_820    ),
    .col_out_821             ( u3_col_out_821    ),
    .col_out_822             ( u3_col_out_822    ),
    .col_out_823             ( u3_col_out_823    ),
    .col_out_824             ( u3_col_out_824    ),
    .col_out_825             ( u3_col_out_825    ),
    .col_out_826             ( u3_col_out_826    ),
    .col_out_827             ( u3_col_out_827    ),
    .col_out_828             ( u3_col_out_828    ),
    .col_out_829             ( u3_col_out_829    ),
    .col_out_830             ( u3_col_out_830    ),
    .col_out_831             ( u3_col_out_831    ),
    .col_out_832             ( u3_col_out_832    ),
    .col_out_833             ( u3_col_out_833    ),
    .col_out_834             ( u3_col_out_834    ),
    .col_out_835             ( u3_col_out_835    ),
    .col_out_836             ( u3_col_out_836    ),
    .col_out_837             ( u3_col_out_837    ),
    .col_out_838             ( u3_col_out_838    ),
    .col_out_839             ( u3_col_out_839    ),
    .col_out_840             ( u3_col_out_840    ),
    .col_out_841             ( u3_col_out_841    ),
    .col_out_842             ( u3_col_out_842    ),
    .col_out_843             ( u3_col_out_843    ),
    .col_out_844             ( u3_col_out_844    ),
    .col_out_845             ( u3_col_out_845    ),
    .col_out_846             ( u3_col_out_846    ),
    .col_out_847             ( u3_col_out_847    ),
    .col_out_848             ( u3_col_out_848    ),
    .col_out_849             ( u3_col_out_849    ),
    .col_out_850             ( u3_col_out_850    ),
    .col_out_851             ( u3_col_out_851    ),
    .col_out_852             ( u3_col_out_852    ),
    .col_out_853             ( u3_col_out_853    ),
    .col_out_854             ( u3_col_out_854    ),
    .col_out_855             ( u3_col_out_855    ),
    .col_out_856             ( u3_col_out_856    ),
    .col_out_857             ( u3_col_out_857    ),
    .col_out_858             ( u3_col_out_858    ),
    .col_out_859             ( u3_col_out_859    ),
    .col_out_860             ( u3_col_out_860    ),
    .col_out_861             ( u3_col_out_861    ),
    .col_out_862             ( u3_col_out_862    ),
    .col_out_863             ( u3_col_out_863    ),
    .col_out_864             ( u3_col_out_864    ),
    .col_out_865             ( u3_col_out_865    ),
    .col_out_866             ( u3_col_out_866    ),
    .col_out_867             ( u3_col_out_867    ),
    .col_out_868             ( u3_col_out_868    ),
    .col_out_869             ( u3_col_out_869    ),
    .col_out_870             ( u3_col_out_870    ),
    .col_out_871             ( u3_col_out_871    ),
    .col_out_872             ( u3_col_out_872    ),
    .col_out_873             ( u3_col_out_873    ),
    .col_out_874             ( u3_col_out_874    ),
    .col_out_875             ( u3_col_out_875    ),
    .col_out_876             ( u3_col_out_876    ),
    .col_out_877             ( u3_col_out_877    ),
    .col_out_878             ( u3_col_out_878    ),
    .col_out_879             ( u3_col_out_879    ),
    .col_out_880             ( u3_col_out_880    ),
    .col_out_881             ( u3_col_out_881    ),
    .col_out_882             ( u3_col_out_882    ),
    .col_out_883             ( u3_col_out_883    ),
    .col_out_884             ( u3_col_out_884    ),
    .col_out_885             ( u3_col_out_885    ),
    .col_out_886             ( u3_col_out_886    ),
    .col_out_887             ( u3_col_out_887    ),
    .col_out_888             ( u3_col_out_888    ),
    .col_out_889             ( u3_col_out_889    ),
    .col_out_890             ( u3_col_out_890    ),
    .col_out_891             ( u3_col_out_891    ),
    .col_out_892             ( u3_col_out_892    ),
    .col_out_893             ( u3_col_out_893    ),
    .col_out_894             ( u3_col_out_894    ),
    .col_out_895             ( u3_col_out_895    ),
    .col_out_896             ( u3_col_out_896    ),
    .col_out_897             ( u3_col_out_897    ),
    .col_out_898             ( u3_col_out_898    ),
    .col_out_899             ( u3_col_out_899    ),
    .col_out_900             ( u3_col_out_900    ),
    .col_out_901             ( u3_col_out_901    ),
    .col_out_902             ( u3_col_out_902    ),
    .col_out_903             ( u3_col_out_903    ),
    .col_out_904             ( u3_col_out_904    ),
    .col_out_905             ( u3_col_out_905    ),
    .col_out_906             ( u3_col_out_906    ),
    .col_out_907             ( u3_col_out_907    ),
    .col_out_908             ( u3_col_out_908    ),
    .col_out_909             ( u3_col_out_909    ),
    .col_out_910             ( u3_col_out_910    ),
    .col_out_911             ( u3_col_out_911    ),
    .col_out_912             ( u3_col_out_912    ),
    .col_out_913             ( u3_col_out_913    ),
    .col_out_914             ( u3_col_out_914    ),
    .col_out_915             ( u3_col_out_915    ),
    .col_out_916             ( u3_col_out_916    ),
    .col_out_917             ( u3_col_out_917    ),
    .col_out_918             ( u3_col_out_918    ),
    .col_out_919             ( u3_col_out_919    ),
    .col_out_920             ( u3_col_out_920    ),
    .col_out_921             ( u3_col_out_921    ),
    .col_out_922             ( u3_col_out_922    ),
    .col_out_923             ( u3_col_out_923    ),
    .col_out_924             ( u3_col_out_924    ),
    .col_out_925             ( u3_col_out_925    ),
    .col_out_926             ( u3_col_out_926    ),
    .col_out_927             ( u3_col_out_927    ),
    .col_out_928             ( u3_col_out_928    ),
    .col_out_929             ( u3_col_out_929    ),
    .col_out_930             ( u3_col_out_930    ),
    .col_out_931             ( u3_col_out_931    ),
    .col_out_932             ( u3_col_out_932    ),
    .col_out_933             ( u3_col_out_933    ),
    .col_out_934             ( u3_col_out_934    ),
    .col_out_935             ( u3_col_out_935    ),
    .col_out_936             ( u3_col_out_936    ),
    .col_out_937             ( u3_col_out_937    ),
    .col_out_938             ( u3_col_out_938    ),
    .col_out_939             ( u3_col_out_939    ),
    .col_out_940             ( u3_col_out_940    ),
    .col_out_941             ( u3_col_out_941    ),
    .col_out_942             ( u3_col_out_942    ),
    .col_out_943             ( u3_col_out_943    ),
    .col_out_944             ( u3_col_out_944    ),
    .col_out_945             ( u3_col_out_945    ),
    .col_out_946             ( u3_col_out_946    ),
    .col_out_947             ( u3_col_out_947    ),
    .col_out_948             ( u3_col_out_948    ),
    .col_out_949             ( u3_col_out_949    ),
    .col_out_950             ( u3_col_out_950    ),
    .col_out_951             ( u3_col_out_951    ),
    .col_out_952             ( u3_col_out_952    ),
    .col_out_953             ( u3_col_out_953    ),
    .col_out_954             ( u3_col_out_954    ),
    .col_out_955             ( u3_col_out_955    ),
    .col_out_956             ( u3_col_out_956    ),
    .col_out_957             ( u3_col_out_957    ),
    .col_out_958             ( u3_col_out_958    ),
    .col_out_959             ( u3_col_out_959    ),
    .col_out_960             ( u3_col_out_960    ),
    .col_out_961             ( u3_col_out_961    ),
    .col_out_962             ( u3_col_out_962    ),
    .col_out_963             ( u3_col_out_963    ),
    .col_out_964             ( u3_col_out_964    ),
    .col_out_965             ( u3_col_out_965    ),
    .col_out_966             ( u3_col_out_966    ),
    .col_out_967             ( u3_col_out_967    ),
    .col_out_968             ( u3_col_out_968    ),
    .col_out_969             ( u3_col_out_969    ),
    .col_out_970             ( u3_col_out_970    ),
    .col_out_971             ( u3_col_out_971    ),
    .col_out_972             ( u3_col_out_972    ),
    .col_out_973             ( u3_col_out_973    ),
    .col_out_974             ( u3_col_out_974    ),
    .col_out_975             ( u3_col_out_975    ),
    .col_out_976             ( u3_col_out_976    ),
    .col_out_977             ( u3_col_out_977    ),
    .col_out_978             ( u3_col_out_978    ),
    .col_out_979             ( u3_col_out_979    ),
    .col_out_980             ( u3_col_out_980    ),
    .col_out_981             ( u3_col_out_981    ),
    .col_out_982             ( u3_col_out_982    ),
    .col_out_983             ( u3_col_out_983    ),
    .col_out_984             ( u3_col_out_984    ),
    .col_out_985             ( u3_col_out_985    ),
    .col_out_986             ( u3_col_out_986    ),
    .col_out_987             ( u3_col_out_987    ),
    .col_out_988             ( u3_col_out_988    ),
    .col_out_989             ( u3_col_out_989    ),
    .col_out_990             ( u3_col_out_990    ),
    .col_out_991             ( u3_col_out_991    ),
    .col_out_992             ( u3_col_out_992    ),
    .col_out_993             ( u3_col_out_993    ),
    .col_out_994             ( u3_col_out_994    ),
    .col_out_995             ( u3_col_out_995    ),
    .col_out_996             ( u3_col_out_996    ),
    .col_out_997             ( u3_col_out_997    ),
    .col_out_998             ( u3_col_out_998    ),
    .col_out_999             ( u3_col_out_999    ),
    .col_out_1000            ( u3_col_out_1000   ),
    .col_out_1001            ( u3_col_out_1001   ),
    .col_out_1002            ( u3_col_out_1002   ),
    .col_out_1003            ( u3_col_out_1003   ),
    .col_out_1004            ( u3_col_out_1004   ),
    .col_out_1005            ( u3_col_out_1005   ),
    .col_out_1006            ( u3_col_out_1006   ),
    .col_out_1007            ( u3_col_out_1007   ),
    .col_out_1008            ( u3_col_out_1008   ),
    .col_out_1009            ( u3_col_out_1009   ),
    .col_out_1010            ( u3_col_out_1010   ),
    .col_out_1011            ( u3_col_out_1011   ),
    .col_out_1012            ( u3_col_out_1012   ),
    .col_out_1013            ( u3_col_out_1013   ),
    .col_out_1014            ( u3_col_out_1014   ),
    .col_out_1015            ( u3_col_out_1015   ),
    .col_out_1016            ( u3_col_out_1016   ),
    .col_out_1017            ( u3_col_out_1017   ),
    .col_out_1018            ( u3_col_out_1018   ),
    .col_out_1019            ( u3_col_out_1019   ),
    .col_out_1020            ( u3_col_out_1020   ),
    .col_out_1021            ( u3_col_out_1021   ),
    .col_out_1022            ( u3_col_out_1022   ),
    .col_out_1023            ( u3_col_out_1023   ),
    .col_out_1024            ( u3_col_out_1024   ),
    .col_out_1025            ( u3_col_out_1025   ),
    .col_out_1026            ( u3_col_out_1026   ),
    .col_out_1027            ( u3_col_out_1027   ),
    .col_out_1028            ( u3_col_out_1028   ),
    .col_out_1029            ( u3_col_out_1029   ),
    .col_out_1030            ( u3_col_out_1030   ),
    .col_out_1031            ( u3_col_out_1031   ),
    .col_out_1032            ( u3_col_out_1032   ),
    .col_out_1033            ( u3_col_out_1033   )
);





















// compressor_array_4_3_1033 Outputs
wire  [2:0]  u4_col_out_0;
wire  [2:0]  u4_col_out_1;
wire  [2:0]  u4_col_out_2;
wire  [2:0]  u4_col_out_3;
wire  [2:0]  u4_col_out_4;
wire  [2:0]  u4_col_out_5;
wire  [2:0]  u4_col_out_6;
wire  [2:0]  u4_col_out_7;
wire  [2:0]  u4_col_out_8;
wire  [2:0]  u4_col_out_9;
wire  [2:0]  u4_col_out_10;
wire  [2:0]  u4_col_out_11;
wire  [2:0]  u4_col_out_12;
wire  [2:0]  u4_col_out_13;
wire  [2:0]  u4_col_out_14;
wire  [2:0]  u4_col_out_15;
wire  [2:0]  u4_col_out_16;
wire  [2:0]  u4_col_out_17;
wire  [2:0]  u4_col_out_18;
wire  [2:0]  u4_col_out_19;
wire  [2:0]  u4_col_out_20;
wire  [2:0]  u4_col_out_21;
wire  [2:0]  u4_col_out_22;
wire  [2:0]  u4_col_out_23;
wire  [2:0]  u4_col_out_24;
wire  [2:0]  u4_col_out_25;
wire  [2:0]  u4_col_out_26;
wire  [2:0]  u4_col_out_27;
wire  [2:0]  u4_col_out_28;
wire  [2:0]  u4_col_out_29;
wire  [2:0]  u4_col_out_30;
wire  [2:0]  u4_col_out_31;
wire  [2:0]  u4_col_out_32;
wire  [2:0]  u4_col_out_33;
wire  [2:0]  u4_col_out_34;
wire  [2:0]  u4_col_out_35;
wire  [2:0]  u4_col_out_36;
wire  [2:0]  u4_col_out_37;
wire  [2:0]  u4_col_out_38;
wire  [2:0]  u4_col_out_39;
wire  [2:0]  u4_col_out_40;
wire  [2:0]  u4_col_out_41;
wire  [2:0]  u4_col_out_42;
wire  [2:0]  u4_col_out_43;
wire  [2:0]  u4_col_out_44;
wire  [2:0]  u4_col_out_45;
wire  [2:0]  u4_col_out_46;
wire  [2:0]  u4_col_out_47;
wire  [2:0]  u4_col_out_48;
wire  [2:0]  u4_col_out_49;
wire  [2:0]  u4_col_out_50;
wire  [2:0]  u4_col_out_51;
wire  [2:0]  u4_col_out_52;
wire  [2:0]  u4_col_out_53;
wire  [2:0]  u4_col_out_54;
wire  [2:0]  u4_col_out_55;
wire  [2:0]  u4_col_out_56;
wire  [2:0]  u4_col_out_57;
wire  [2:0]  u4_col_out_58;
wire  [2:0]  u4_col_out_59;
wire  [2:0]  u4_col_out_60;
wire  [2:0]  u4_col_out_61;
wire  [2:0]  u4_col_out_62;
wire  [2:0]  u4_col_out_63;
wire  [2:0]  u4_col_out_64;
wire  [2:0]  u4_col_out_65;
wire  [2:0]  u4_col_out_66;
wire  [2:0]  u4_col_out_67;
wire  [2:0]  u4_col_out_68;
wire  [2:0]  u4_col_out_69;
wire  [2:0]  u4_col_out_70;
wire  [2:0]  u4_col_out_71;
wire  [2:0]  u4_col_out_72;
wire  [2:0]  u4_col_out_73;
wire  [2:0]  u4_col_out_74;
wire  [2:0]  u4_col_out_75;
wire  [2:0]  u4_col_out_76;
wire  [2:0]  u4_col_out_77;
wire  [2:0]  u4_col_out_78;
wire  [2:0]  u4_col_out_79;
wire  [2:0]  u4_col_out_80;
wire  [2:0]  u4_col_out_81;
wire  [2:0]  u4_col_out_82;
wire  [2:0]  u4_col_out_83;
wire  [2:0]  u4_col_out_84;
wire  [2:0]  u4_col_out_85;
wire  [2:0]  u4_col_out_86;
wire  [2:0]  u4_col_out_87;
wire  [2:0]  u4_col_out_88;
wire  [2:0]  u4_col_out_89;
wire  [2:0]  u4_col_out_90;
wire  [2:0]  u4_col_out_91;
wire  [2:0]  u4_col_out_92;
wire  [2:0]  u4_col_out_93;
wire  [2:0]  u4_col_out_94;
wire  [2:0]  u4_col_out_95;
wire  [2:0]  u4_col_out_96;
wire  [2:0]  u4_col_out_97;
wire  [2:0]  u4_col_out_98;
wire  [2:0]  u4_col_out_99;
wire  [2:0]  u4_col_out_100;
wire  [2:0]  u4_col_out_101;
wire  [2:0]  u4_col_out_102;
wire  [2:0]  u4_col_out_103;
wire  [2:0]  u4_col_out_104;
wire  [2:0]  u4_col_out_105;
wire  [2:0]  u4_col_out_106;
wire  [2:0]  u4_col_out_107;
wire  [2:0]  u4_col_out_108;
wire  [2:0]  u4_col_out_109;
wire  [2:0]  u4_col_out_110;
wire  [2:0]  u4_col_out_111;
wire  [2:0]  u4_col_out_112;
wire  [2:0]  u4_col_out_113;
wire  [2:0]  u4_col_out_114;
wire  [2:0]  u4_col_out_115;
wire  [2:0]  u4_col_out_116;
wire  [2:0]  u4_col_out_117;
wire  [2:0]  u4_col_out_118;
wire  [2:0]  u4_col_out_119;
wire  [2:0]  u4_col_out_120;
wire  [2:0]  u4_col_out_121;
wire  [2:0]  u4_col_out_122;
wire  [2:0]  u4_col_out_123;
wire  [2:0]  u4_col_out_124;
wire  [2:0]  u4_col_out_125;
wire  [2:0]  u4_col_out_126;
wire  [2:0]  u4_col_out_127;
wire  [2:0]  u4_col_out_128;
wire  [2:0]  u4_col_out_129;
wire  [2:0]  u4_col_out_130;
wire  [2:0]  u4_col_out_131;
wire  [2:0]  u4_col_out_132;
wire  [2:0]  u4_col_out_133;
wire  [2:0]  u4_col_out_134;
wire  [2:0]  u4_col_out_135;
wire  [2:0]  u4_col_out_136;
wire  [2:0]  u4_col_out_137;
wire  [2:0]  u4_col_out_138;
wire  [2:0]  u4_col_out_139;
wire  [2:0]  u4_col_out_140;
wire  [2:0]  u4_col_out_141;
wire  [2:0]  u4_col_out_142;
wire  [2:0]  u4_col_out_143;
wire  [2:0]  u4_col_out_144;
wire  [2:0]  u4_col_out_145;
wire  [2:0]  u4_col_out_146;
wire  [2:0]  u4_col_out_147;
wire  [2:0]  u4_col_out_148;
wire  [2:0]  u4_col_out_149;
wire  [2:0]  u4_col_out_150;
wire  [2:0]  u4_col_out_151;
wire  [2:0]  u4_col_out_152;
wire  [2:0]  u4_col_out_153;
wire  [2:0]  u4_col_out_154;
wire  [2:0]  u4_col_out_155;
wire  [2:0]  u4_col_out_156;
wire  [2:0]  u4_col_out_157;
wire  [2:0]  u4_col_out_158;
wire  [2:0]  u4_col_out_159;
wire  [2:0]  u4_col_out_160;
wire  [2:0]  u4_col_out_161;
wire  [2:0]  u4_col_out_162;
wire  [2:0]  u4_col_out_163;
wire  [2:0]  u4_col_out_164;
wire  [2:0]  u4_col_out_165;
wire  [2:0]  u4_col_out_166;
wire  [2:0]  u4_col_out_167;
wire  [2:0]  u4_col_out_168;
wire  [2:0]  u4_col_out_169;
wire  [2:0]  u4_col_out_170;
wire  [2:0]  u4_col_out_171;
wire  [2:0]  u4_col_out_172;
wire  [2:0]  u4_col_out_173;
wire  [2:0]  u4_col_out_174;
wire  [2:0]  u4_col_out_175;
wire  [2:0]  u4_col_out_176;
wire  [2:0]  u4_col_out_177;
wire  [2:0]  u4_col_out_178;
wire  [2:0]  u4_col_out_179;
wire  [2:0]  u4_col_out_180;
wire  [2:0]  u4_col_out_181;
wire  [2:0]  u4_col_out_182;
wire  [2:0]  u4_col_out_183;
wire  [2:0]  u4_col_out_184;
wire  [2:0]  u4_col_out_185;
wire  [2:0]  u4_col_out_186;
wire  [2:0]  u4_col_out_187;
wire  [2:0]  u4_col_out_188;
wire  [2:0]  u4_col_out_189;
wire  [2:0]  u4_col_out_190;
wire  [2:0]  u4_col_out_191;
wire  [2:0]  u4_col_out_192;
wire  [2:0]  u4_col_out_193;
wire  [2:0]  u4_col_out_194;
wire  [2:0]  u4_col_out_195;
wire  [2:0]  u4_col_out_196;
wire  [2:0]  u4_col_out_197;
wire  [2:0]  u4_col_out_198;
wire  [2:0]  u4_col_out_199;
wire  [2:0]  u4_col_out_200;
wire  [2:0]  u4_col_out_201;
wire  [2:0]  u4_col_out_202;
wire  [2:0]  u4_col_out_203;
wire  [2:0]  u4_col_out_204;
wire  [2:0]  u4_col_out_205;
wire  [2:0]  u4_col_out_206;
wire  [2:0]  u4_col_out_207;
wire  [2:0]  u4_col_out_208;
wire  [2:0]  u4_col_out_209;
wire  [2:0]  u4_col_out_210;
wire  [2:0]  u4_col_out_211;
wire  [2:0]  u4_col_out_212;
wire  [2:0]  u4_col_out_213;
wire  [2:0]  u4_col_out_214;
wire  [2:0]  u4_col_out_215;
wire  [2:0]  u4_col_out_216;
wire  [2:0]  u4_col_out_217;
wire  [2:0]  u4_col_out_218;
wire  [2:0]  u4_col_out_219;
wire  [2:0]  u4_col_out_220;
wire  [2:0]  u4_col_out_221;
wire  [2:0]  u4_col_out_222;
wire  [2:0]  u4_col_out_223;
wire  [2:0]  u4_col_out_224;
wire  [2:0]  u4_col_out_225;
wire  [2:0]  u4_col_out_226;
wire  [2:0]  u4_col_out_227;
wire  [2:0]  u4_col_out_228;
wire  [2:0]  u4_col_out_229;
wire  [2:0]  u4_col_out_230;
wire  [2:0]  u4_col_out_231;
wire  [2:0]  u4_col_out_232;
wire  [2:0]  u4_col_out_233;
wire  [2:0]  u4_col_out_234;
wire  [2:0]  u4_col_out_235;
wire  [2:0]  u4_col_out_236;
wire  [2:0]  u4_col_out_237;
wire  [2:0]  u4_col_out_238;
wire  [2:0]  u4_col_out_239;
wire  [2:0]  u4_col_out_240;
wire  [2:0]  u4_col_out_241;
wire  [2:0]  u4_col_out_242;
wire  [2:0]  u4_col_out_243;
wire  [2:0]  u4_col_out_244;
wire  [2:0]  u4_col_out_245;
wire  [2:0]  u4_col_out_246;
wire  [2:0]  u4_col_out_247;
wire  [2:0]  u4_col_out_248;
wire  [2:0]  u4_col_out_249;
wire  [2:0]  u4_col_out_250;
wire  [2:0]  u4_col_out_251;
wire  [2:0]  u4_col_out_252;
wire  [2:0]  u4_col_out_253;
wire  [2:0]  u4_col_out_254;
wire  [2:0]  u4_col_out_255;
wire  [2:0]  u4_col_out_256;
wire  [2:0]  u4_col_out_257;
wire  [2:0]  u4_col_out_258;
wire  [2:0]  u4_col_out_259;
wire  [2:0]  u4_col_out_260;
wire  [2:0]  u4_col_out_261;
wire  [2:0]  u4_col_out_262;
wire  [2:0]  u4_col_out_263;
wire  [2:0]  u4_col_out_264;
wire  [2:0]  u4_col_out_265;
wire  [2:0]  u4_col_out_266;
wire  [2:0]  u4_col_out_267;
wire  [2:0]  u4_col_out_268;
wire  [2:0]  u4_col_out_269;
wire  [2:0]  u4_col_out_270;
wire  [2:0]  u4_col_out_271;
wire  [2:0]  u4_col_out_272;
wire  [2:0]  u4_col_out_273;
wire  [2:0]  u4_col_out_274;
wire  [2:0]  u4_col_out_275;
wire  [2:0]  u4_col_out_276;
wire  [2:0]  u4_col_out_277;
wire  [2:0]  u4_col_out_278;
wire  [2:0]  u4_col_out_279;
wire  [2:0]  u4_col_out_280;
wire  [2:0]  u4_col_out_281;
wire  [2:0]  u4_col_out_282;
wire  [2:0]  u4_col_out_283;
wire  [2:0]  u4_col_out_284;
wire  [2:0]  u4_col_out_285;
wire  [2:0]  u4_col_out_286;
wire  [2:0]  u4_col_out_287;
wire  [2:0]  u4_col_out_288;
wire  [2:0]  u4_col_out_289;
wire  [2:0]  u4_col_out_290;
wire  [2:0]  u4_col_out_291;
wire  [2:0]  u4_col_out_292;
wire  [2:0]  u4_col_out_293;
wire  [2:0]  u4_col_out_294;
wire  [2:0]  u4_col_out_295;
wire  [2:0]  u4_col_out_296;
wire  [2:0]  u4_col_out_297;
wire  [2:0]  u4_col_out_298;
wire  [2:0]  u4_col_out_299;
wire  [2:0]  u4_col_out_300;
wire  [2:0]  u4_col_out_301;
wire  [2:0]  u4_col_out_302;
wire  [2:0]  u4_col_out_303;
wire  [2:0]  u4_col_out_304;
wire  [2:0]  u4_col_out_305;
wire  [2:0]  u4_col_out_306;
wire  [2:0]  u4_col_out_307;
wire  [2:0]  u4_col_out_308;
wire  [2:0]  u4_col_out_309;
wire  [2:0]  u4_col_out_310;
wire  [2:0]  u4_col_out_311;
wire  [2:0]  u4_col_out_312;
wire  [2:0]  u4_col_out_313;
wire  [2:0]  u4_col_out_314;
wire  [2:0]  u4_col_out_315;
wire  [2:0]  u4_col_out_316;
wire  [2:0]  u4_col_out_317;
wire  [2:0]  u4_col_out_318;
wire  [2:0]  u4_col_out_319;
wire  [2:0]  u4_col_out_320;
wire  [2:0]  u4_col_out_321;
wire  [2:0]  u4_col_out_322;
wire  [2:0]  u4_col_out_323;
wire  [2:0]  u4_col_out_324;
wire  [2:0]  u4_col_out_325;
wire  [2:0]  u4_col_out_326;
wire  [2:0]  u4_col_out_327;
wire  [2:0]  u4_col_out_328;
wire  [2:0]  u4_col_out_329;
wire  [2:0]  u4_col_out_330;
wire  [2:0]  u4_col_out_331;
wire  [2:0]  u4_col_out_332;
wire  [2:0]  u4_col_out_333;
wire  [2:0]  u4_col_out_334;
wire  [2:0]  u4_col_out_335;
wire  [2:0]  u4_col_out_336;
wire  [2:0]  u4_col_out_337;
wire  [2:0]  u4_col_out_338;
wire  [2:0]  u4_col_out_339;
wire  [2:0]  u4_col_out_340;
wire  [2:0]  u4_col_out_341;
wire  [2:0]  u4_col_out_342;
wire  [2:0]  u4_col_out_343;
wire  [2:0]  u4_col_out_344;
wire  [2:0]  u4_col_out_345;
wire  [2:0]  u4_col_out_346;
wire  [2:0]  u4_col_out_347;
wire  [2:0]  u4_col_out_348;
wire  [2:0]  u4_col_out_349;
wire  [2:0]  u4_col_out_350;
wire  [2:0]  u4_col_out_351;
wire  [2:0]  u4_col_out_352;
wire  [2:0]  u4_col_out_353;
wire  [2:0]  u4_col_out_354;
wire  [2:0]  u4_col_out_355;
wire  [2:0]  u4_col_out_356;
wire  [2:0]  u4_col_out_357;
wire  [2:0]  u4_col_out_358;
wire  [2:0]  u4_col_out_359;
wire  [2:0]  u4_col_out_360;
wire  [2:0]  u4_col_out_361;
wire  [2:0]  u4_col_out_362;
wire  [2:0]  u4_col_out_363;
wire  [2:0]  u4_col_out_364;
wire  [2:0]  u4_col_out_365;
wire  [2:0]  u4_col_out_366;
wire  [2:0]  u4_col_out_367;
wire  [2:0]  u4_col_out_368;
wire  [2:0]  u4_col_out_369;
wire  [2:0]  u4_col_out_370;
wire  [2:0]  u4_col_out_371;
wire  [2:0]  u4_col_out_372;
wire  [2:0]  u4_col_out_373;
wire  [2:0]  u4_col_out_374;
wire  [2:0]  u4_col_out_375;
wire  [2:0]  u4_col_out_376;
wire  [2:0]  u4_col_out_377;
wire  [2:0]  u4_col_out_378;
wire  [2:0]  u4_col_out_379;
wire  [2:0]  u4_col_out_380;
wire  [2:0]  u4_col_out_381;
wire  [2:0]  u4_col_out_382;
wire  [2:0]  u4_col_out_383;
wire  [2:0]  u4_col_out_384;
wire  [2:0]  u4_col_out_385;
wire  [2:0]  u4_col_out_386;
wire  [2:0]  u4_col_out_387;
wire  [2:0]  u4_col_out_388;
wire  [2:0]  u4_col_out_389;
wire  [2:0]  u4_col_out_390;
wire  [2:0]  u4_col_out_391;
wire  [2:0]  u4_col_out_392;
wire  [2:0]  u4_col_out_393;
wire  [2:0]  u4_col_out_394;
wire  [2:0]  u4_col_out_395;
wire  [2:0]  u4_col_out_396;
wire  [2:0]  u4_col_out_397;
wire  [2:0]  u4_col_out_398;
wire  [2:0]  u4_col_out_399;
wire  [2:0]  u4_col_out_400;
wire  [2:0]  u4_col_out_401;
wire  [2:0]  u4_col_out_402;
wire  [2:0]  u4_col_out_403;
wire  [2:0]  u4_col_out_404;
wire  [2:0]  u4_col_out_405;
wire  [2:0]  u4_col_out_406;
wire  [2:0]  u4_col_out_407;
wire  [2:0]  u4_col_out_408;
wire  [2:0]  u4_col_out_409;
wire  [2:0]  u4_col_out_410;
wire  [2:0]  u4_col_out_411;
wire  [2:0]  u4_col_out_412;
wire  [2:0]  u4_col_out_413;
wire  [2:0]  u4_col_out_414;
wire  [2:0]  u4_col_out_415;
wire  [2:0]  u4_col_out_416;
wire  [2:0]  u4_col_out_417;
wire  [2:0]  u4_col_out_418;
wire  [2:0]  u4_col_out_419;
wire  [2:0]  u4_col_out_420;
wire  [2:0]  u4_col_out_421;
wire  [2:0]  u4_col_out_422;
wire  [2:0]  u4_col_out_423;
wire  [2:0]  u4_col_out_424;
wire  [2:0]  u4_col_out_425;
wire  [2:0]  u4_col_out_426;
wire  [2:0]  u4_col_out_427;
wire  [2:0]  u4_col_out_428;
wire  [2:0]  u4_col_out_429;
wire  [2:0]  u4_col_out_430;
wire  [2:0]  u4_col_out_431;
wire  [2:0]  u4_col_out_432;
wire  [2:0]  u4_col_out_433;
wire  [2:0]  u4_col_out_434;
wire  [2:0]  u4_col_out_435;
wire  [2:0]  u4_col_out_436;
wire  [2:0]  u4_col_out_437;
wire  [2:0]  u4_col_out_438;
wire  [2:0]  u4_col_out_439;
wire  [2:0]  u4_col_out_440;
wire  [2:0]  u4_col_out_441;
wire  [2:0]  u4_col_out_442;
wire  [2:0]  u4_col_out_443;
wire  [2:0]  u4_col_out_444;
wire  [2:0]  u4_col_out_445;
wire  [2:0]  u4_col_out_446;
wire  [2:0]  u4_col_out_447;
wire  [2:0]  u4_col_out_448;
wire  [2:0]  u4_col_out_449;
wire  [2:0]  u4_col_out_450;
wire  [2:0]  u4_col_out_451;
wire  [2:0]  u4_col_out_452;
wire  [2:0]  u4_col_out_453;
wire  [2:0]  u4_col_out_454;
wire  [2:0]  u4_col_out_455;
wire  [2:0]  u4_col_out_456;
wire  [2:0]  u4_col_out_457;
wire  [2:0]  u4_col_out_458;
wire  [2:0]  u4_col_out_459;
wire  [2:0]  u4_col_out_460;
wire  [2:0]  u4_col_out_461;
wire  [2:0]  u4_col_out_462;
wire  [2:0]  u4_col_out_463;
wire  [2:0]  u4_col_out_464;
wire  [2:0]  u4_col_out_465;
wire  [2:0]  u4_col_out_466;
wire  [2:0]  u4_col_out_467;
wire  [2:0]  u4_col_out_468;
wire  [2:0]  u4_col_out_469;
wire  [2:0]  u4_col_out_470;
wire  [2:0]  u4_col_out_471;
wire  [2:0]  u4_col_out_472;
wire  [2:0]  u4_col_out_473;
wire  [2:0]  u4_col_out_474;
wire  [2:0]  u4_col_out_475;
wire  [2:0]  u4_col_out_476;
wire  [2:0]  u4_col_out_477;
wire  [2:0]  u4_col_out_478;
wire  [2:0]  u4_col_out_479;
wire  [2:0]  u4_col_out_480;
wire  [2:0]  u4_col_out_481;
wire  [2:0]  u4_col_out_482;
wire  [2:0]  u4_col_out_483;
wire  [2:0]  u4_col_out_484;
wire  [2:0]  u4_col_out_485;
wire  [2:0]  u4_col_out_486;
wire  [2:0]  u4_col_out_487;
wire  [2:0]  u4_col_out_488;
wire  [2:0]  u4_col_out_489;
wire  [2:0]  u4_col_out_490;
wire  [2:0]  u4_col_out_491;
wire  [2:0]  u4_col_out_492;
wire  [2:0]  u4_col_out_493;
wire  [2:0]  u4_col_out_494;
wire  [2:0]  u4_col_out_495;
wire  [2:0]  u4_col_out_496;
wire  [2:0]  u4_col_out_497;
wire  [2:0]  u4_col_out_498;
wire  [2:0]  u4_col_out_499;
wire  [2:0]  u4_col_out_500;
wire  [2:0]  u4_col_out_501;
wire  [2:0]  u4_col_out_502;
wire  [2:0]  u4_col_out_503;
wire  [2:0]  u4_col_out_504;
wire  [2:0]  u4_col_out_505;
wire  [2:0]  u4_col_out_506;
wire  [2:0]  u4_col_out_507;
wire  [2:0]  u4_col_out_508;
wire  [2:0]  u4_col_out_509;
wire  [2:0]  u4_col_out_510;
wire  [2:0]  u4_col_out_511;
wire  [2:0]  u4_col_out_512;
wire  [2:0]  u4_col_out_513;
wire  [2:0]  u4_col_out_514;
wire  [2:0]  u4_col_out_515;
wire  [2:0]  u4_col_out_516;
wire  [2:0]  u4_col_out_517;
wire  [2:0]  u4_col_out_518;
wire  [2:0]  u4_col_out_519;
wire  [2:0]  u4_col_out_520;
wire  [2:0]  u4_col_out_521;
wire  [2:0]  u4_col_out_522;
wire  [2:0]  u4_col_out_523;
wire  [2:0]  u4_col_out_524;
wire  [2:0]  u4_col_out_525;
wire  [2:0]  u4_col_out_526;
wire  [2:0]  u4_col_out_527;
wire  [2:0]  u4_col_out_528;
wire  [2:0]  u4_col_out_529;
wire  [2:0]  u4_col_out_530;
wire  [2:0]  u4_col_out_531;
wire  [2:0]  u4_col_out_532;
wire  [2:0]  u4_col_out_533;
wire  [2:0]  u4_col_out_534;
wire  [2:0]  u4_col_out_535;
wire  [2:0]  u4_col_out_536;
wire  [2:0]  u4_col_out_537;
wire  [2:0]  u4_col_out_538;
wire  [2:0]  u4_col_out_539;
wire  [2:0]  u4_col_out_540;
wire  [2:0]  u4_col_out_541;
wire  [2:0]  u4_col_out_542;
wire  [2:0]  u4_col_out_543;
wire  [2:0]  u4_col_out_544;
wire  [2:0]  u4_col_out_545;
wire  [2:0]  u4_col_out_546;
wire  [2:0]  u4_col_out_547;
wire  [2:0]  u4_col_out_548;
wire  [2:0]  u4_col_out_549;
wire  [2:0]  u4_col_out_550;
wire  [2:0]  u4_col_out_551;
wire  [2:0]  u4_col_out_552;
wire  [2:0]  u4_col_out_553;
wire  [2:0]  u4_col_out_554;
wire  [2:0]  u4_col_out_555;
wire  [2:0]  u4_col_out_556;
wire  [2:0]  u4_col_out_557;
wire  [2:0]  u4_col_out_558;
wire  [2:0]  u4_col_out_559;
wire  [2:0]  u4_col_out_560;
wire  [2:0]  u4_col_out_561;
wire  [2:0]  u4_col_out_562;
wire  [2:0]  u4_col_out_563;
wire  [2:0]  u4_col_out_564;
wire  [2:0]  u4_col_out_565;
wire  [2:0]  u4_col_out_566;
wire  [2:0]  u4_col_out_567;
wire  [2:0]  u4_col_out_568;
wire  [2:0]  u4_col_out_569;
wire  [2:0]  u4_col_out_570;
wire  [2:0]  u4_col_out_571;
wire  [2:0]  u4_col_out_572;
wire  [2:0]  u4_col_out_573;
wire  [2:0]  u4_col_out_574;
wire  [2:0]  u4_col_out_575;
wire  [2:0]  u4_col_out_576;
wire  [2:0]  u4_col_out_577;
wire  [2:0]  u4_col_out_578;
wire  [2:0]  u4_col_out_579;
wire  [2:0]  u4_col_out_580;
wire  [2:0]  u4_col_out_581;
wire  [2:0]  u4_col_out_582;
wire  [2:0]  u4_col_out_583;
wire  [2:0]  u4_col_out_584;
wire  [2:0]  u4_col_out_585;
wire  [2:0]  u4_col_out_586;
wire  [2:0]  u4_col_out_587;
wire  [2:0]  u4_col_out_588;
wire  [2:0]  u4_col_out_589;
wire  [2:0]  u4_col_out_590;
wire  [2:0]  u4_col_out_591;
wire  [2:0]  u4_col_out_592;
wire  [2:0]  u4_col_out_593;
wire  [2:0]  u4_col_out_594;
wire  [2:0]  u4_col_out_595;
wire  [2:0]  u4_col_out_596;
wire  [2:0]  u4_col_out_597;
wire  [2:0]  u4_col_out_598;
wire  [2:0]  u4_col_out_599;
wire  [2:0]  u4_col_out_600;
wire  [2:0]  u4_col_out_601;
wire  [2:0]  u4_col_out_602;
wire  [2:0]  u4_col_out_603;
wire  [2:0]  u4_col_out_604;
wire  [2:0]  u4_col_out_605;
wire  [2:0]  u4_col_out_606;
wire  [2:0]  u4_col_out_607;
wire  [2:0]  u4_col_out_608;
wire  [2:0]  u4_col_out_609;
wire  [2:0]  u4_col_out_610;
wire  [2:0]  u4_col_out_611;
wire  [2:0]  u4_col_out_612;
wire  [2:0]  u4_col_out_613;
wire  [2:0]  u4_col_out_614;
wire  [2:0]  u4_col_out_615;
wire  [2:0]  u4_col_out_616;
wire  [2:0]  u4_col_out_617;
wire  [2:0]  u4_col_out_618;
wire  [2:0]  u4_col_out_619;
wire  [2:0]  u4_col_out_620;
wire  [2:0]  u4_col_out_621;
wire  [2:0]  u4_col_out_622;
wire  [2:0]  u4_col_out_623;
wire  [2:0]  u4_col_out_624;
wire  [2:0]  u4_col_out_625;
wire  [2:0]  u4_col_out_626;
wire  [2:0]  u4_col_out_627;
wire  [2:0]  u4_col_out_628;
wire  [2:0]  u4_col_out_629;
wire  [2:0]  u4_col_out_630;
wire  [2:0]  u4_col_out_631;
wire  [2:0]  u4_col_out_632;
wire  [2:0]  u4_col_out_633;
wire  [2:0]  u4_col_out_634;
wire  [2:0]  u4_col_out_635;
wire  [2:0]  u4_col_out_636;
wire  [2:0]  u4_col_out_637;
wire  [2:0]  u4_col_out_638;
wire  [2:0]  u4_col_out_639;
wire  [2:0]  u4_col_out_640;
wire  [2:0]  u4_col_out_641;
wire  [2:0]  u4_col_out_642;
wire  [2:0]  u4_col_out_643;
wire  [2:0]  u4_col_out_644;
wire  [2:0]  u4_col_out_645;
wire  [2:0]  u4_col_out_646;
wire  [2:0]  u4_col_out_647;
wire  [2:0]  u4_col_out_648;
wire  [2:0]  u4_col_out_649;
wire  [2:0]  u4_col_out_650;
wire  [2:0]  u4_col_out_651;
wire  [2:0]  u4_col_out_652;
wire  [2:0]  u4_col_out_653;
wire  [2:0]  u4_col_out_654;
wire  [2:0]  u4_col_out_655;
wire  [2:0]  u4_col_out_656;
wire  [2:0]  u4_col_out_657;
wire  [2:0]  u4_col_out_658;
wire  [2:0]  u4_col_out_659;
wire  [2:0]  u4_col_out_660;
wire  [2:0]  u4_col_out_661;
wire  [2:0]  u4_col_out_662;
wire  [2:0]  u4_col_out_663;
wire  [2:0]  u4_col_out_664;
wire  [2:0]  u4_col_out_665;
wire  [2:0]  u4_col_out_666;
wire  [2:0]  u4_col_out_667;
wire  [2:0]  u4_col_out_668;
wire  [2:0]  u4_col_out_669;
wire  [2:0]  u4_col_out_670;
wire  [2:0]  u4_col_out_671;
wire  [2:0]  u4_col_out_672;
wire  [2:0]  u4_col_out_673;
wire  [2:0]  u4_col_out_674;
wire  [2:0]  u4_col_out_675;
wire  [2:0]  u4_col_out_676;
wire  [2:0]  u4_col_out_677;
wire  [2:0]  u4_col_out_678;
wire  [2:0]  u4_col_out_679;
wire  [2:0]  u4_col_out_680;
wire  [2:0]  u4_col_out_681;
wire  [2:0]  u4_col_out_682;
wire  [2:0]  u4_col_out_683;
wire  [2:0]  u4_col_out_684;
wire  [2:0]  u4_col_out_685;
wire  [2:0]  u4_col_out_686;
wire  [2:0]  u4_col_out_687;
wire  [2:0]  u4_col_out_688;
wire  [2:0]  u4_col_out_689;
wire  [2:0]  u4_col_out_690;
wire  [2:0]  u4_col_out_691;
wire  [2:0]  u4_col_out_692;
wire  [2:0]  u4_col_out_693;
wire  [2:0]  u4_col_out_694;
wire  [2:0]  u4_col_out_695;
wire  [2:0]  u4_col_out_696;
wire  [2:0]  u4_col_out_697;
wire  [2:0]  u4_col_out_698;
wire  [2:0]  u4_col_out_699;
wire  [2:0]  u4_col_out_700;
wire  [2:0]  u4_col_out_701;
wire  [2:0]  u4_col_out_702;
wire  [2:0]  u4_col_out_703;
wire  [2:0]  u4_col_out_704;
wire  [2:0]  u4_col_out_705;
wire  [2:0]  u4_col_out_706;
wire  [2:0]  u4_col_out_707;
wire  [2:0]  u4_col_out_708;
wire  [2:0]  u4_col_out_709;
wire  [2:0]  u4_col_out_710;
wire  [2:0]  u4_col_out_711;
wire  [2:0]  u4_col_out_712;
wire  [2:0]  u4_col_out_713;
wire  [2:0]  u4_col_out_714;
wire  [2:0]  u4_col_out_715;
wire  [2:0]  u4_col_out_716;
wire  [2:0]  u4_col_out_717;
wire  [2:0]  u4_col_out_718;
wire  [2:0]  u4_col_out_719;
wire  [2:0]  u4_col_out_720;
wire  [2:0]  u4_col_out_721;
wire  [2:0]  u4_col_out_722;
wire  [2:0]  u4_col_out_723;
wire  [2:0]  u4_col_out_724;
wire  [2:0]  u4_col_out_725;
wire  [2:0]  u4_col_out_726;
wire  [2:0]  u4_col_out_727;
wire  [2:0]  u4_col_out_728;
wire  [2:0]  u4_col_out_729;
wire  [2:0]  u4_col_out_730;
wire  [2:0]  u4_col_out_731;
wire  [2:0]  u4_col_out_732;
wire  [2:0]  u4_col_out_733;
wire  [2:0]  u4_col_out_734;
wire  [2:0]  u4_col_out_735;
wire  [2:0]  u4_col_out_736;
wire  [2:0]  u4_col_out_737;
wire  [2:0]  u4_col_out_738;
wire  [2:0]  u4_col_out_739;
wire  [2:0]  u4_col_out_740;
wire  [2:0]  u4_col_out_741;
wire  [2:0]  u4_col_out_742;
wire  [2:0]  u4_col_out_743;
wire  [2:0]  u4_col_out_744;
wire  [2:0]  u4_col_out_745;
wire  [2:0]  u4_col_out_746;
wire  [2:0]  u4_col_out_747;
wire  [2:0]  u4_col_out_748;
wire  [2:0]  u4_col_out_749;
wire  [2:0]  u4_col_out_750;
wire  [2:0]  u4_col_out_751;
wire  [2:0]  u4_col_out_752;
wire  [2:0]  u4_col_out_753;
wire  [2:0]  u4_col_out_754;
wire  [2:0]  u4_col_out_755;
wire  [2:0]  u4_col_out_756;
wire  [2:0]  u4_col_out_757;
wire  [2:0]  u4_col_out_758;
wire  [2:0]  u4_col_out_759;
wire  [2:0]  u4_col_out_760;
wire  [2:0]  u4_col_out_761;
wire  [2:0]  u4_col_out_762;
wire  [2:0]  u4_col_out_763;
wire  [2:0]  u4_col_out_764;
wire  [2:0]  u4_col_out_765;
wire  [2:0]  u4_col_out_766;
wire  [2:0]  u4_col_out_767;
wire  [2:0]  u4_col_out_768;
wire  [2:0]  u4_col_out_769;
wire  [2:0]  u4_col_out_770;
wire  [2:0]  u4_col_out_771;
wire  [2:0]  u4_col_out_772;
wire  [2:0]  u4_col_out_773;
wire  [2:0]  u4_col_out_774;
wire  [2:0]  u4_col_out_775;
wire  [2:0]  u4_col_out_776;
wire  [2:0]  u4_col_out_777;
wire  [2:0]  u4_col_out_778;
wire  [2:0]  u4_col_out_779;
wire  [2:0]  u4_col_out_780;
wire  [2:0]  u4_col_out_781;
wire  [2:0]  u4_col_out_782;
wire  [2:0]  u4_col_out_783;
wire  [2:0]  u4_col_out_784;
wire  [2:0]  u4_col_out_785;
wire  [2:0]  u4_col_out_786;
wire  [2:0]  u4_col_out_787;
wire  [2:0]  u4_col_out_788;
wire  [2:0]  u4_col_out_789;
wire  [2:0]  u4_col_out_790;
wire  [2:0]  u4_col_out_791;
wire  [2:0]  u4_col_out_792;
wire  [2:0]  u4_col_out_793;
wire  [2:0]  u4_col_out_794;
wire  [2:0]  u4_col_out_795;
wire  [2:0]  u4_col_out_796;
wire  [2:0]  u4_col_out_797;
wire  [2:0]  u4_col_out_798;
wire  [2:0]  u4_col_out_799;
wire  [2:0]  u4_col_out_800;
wire  [2:0]  u4_col_out_801;
wire  [2:0]  u4_col_out_802;
wire  [2:0]  u4_col_out_803;
wire  [2:0]  u4_col_out_804;
wire  [2:0]  u4_col_out_805;
wire  [2:0]  u4_col_out_806;
wire  [2:0]  u4_col_out_807;
wire  [2:0]  u4_col_out_808;
wire  [2:0]  u4_col_out_809;
wire  [2:0]  u4_col_out_810;
wire  [2:0]  u4_col_out_811;
wire  [2:0]  u4_col_out_812;
wire  [2:0]  u4_col_out_813;
wire  [2:0]  u4_col_out_814;
wire  [2:0]  u4_col_out_815;
wire  [2:0]  u4_col_out_816;
wire  [2:0]  u4_col_out_817;
wire  [2:0]  u4_col_out_818;
wire  [2:0]  u4_col_out_819;
wire  [2:0]  u4_col_out_820;
wire  [2:0]  u4_col_out_821;
wire  [2:0]  u4_col_out_822;
wire  [2:0]  u4_col_out_823;
wire  [2:0]  u4_col_out_824;
wire  [2:0]  u4_col_out_825;
wire  [2:0]  u4_col_out_826;
wire  [2:0]  u4_col_out_827;
wire  [2:0]  u4_col_out_828;
wire  [2:0]  u4_col_out_829;
wire  [2:0]  u4_col_out_830;
wire  [2:0]  u4_col_out_831;
wire  [2:0]  u4_col_out_832;
wire  [2:0]  u4_col_out_833;
wire  [2:0]  u4_col_out_834;
wire  [2:0]  u4_col_out_835;
wire  [2:0]  u4_col_out_836;
wire  [2:0]  u4_col_out_837;
wire  [2:0]  u4_col_out_838;
wire  [2:0]  u4_col_out_839;
wire  [2:0]  u4_col_out_840;
wire  [2:0]  u4_col_out_841;
wire  [2:0]  u4_col_out_842;
wire  [2:0]  u4_col_out_843;
wire  [2:0]  u4_col_out_844;
wire  [2:0]  u4_col_out_845;
wire  [2:0]  u4_col_out_846;
wire  [2:0]  u4_col_out_847;
wire  [2:0]  u4_col_out_848;
wire  [2:0]  u4_col_out_849;
wire  [2:0]  u4_col_out_850;
wire  [2:0]  u4_col_out_851;
wire  [2:0]  u4_col_out_852;
wire  [2:0]  u4_col_out_853;
wire  [2:0]  u4_col_out_854;
wire  [2:0]  u4_col_out_855;
wire  [2:0]  u4_col_out_856;
wire  [2:0]  u4_col_out_857;
wire  [2:0]  u4_col_out_858;
wire  [2:0]  u4_col_out_859;
wire  [2:0]  u4_col_out_860;
wire  [2:0]  u4_col_out_861;
wire  [2:0]  u4_col_out_862;
wire  [2:0]  u4_col_out_863;
wire  [2:0]  u4_col_out_864;
wire  [2:0]  u4_col_out_865;
wire  [2:0]  u4_col_out_866;
wire  [2:0]  u4_col_out_867;
wire  [2:0]  u4_col_out_868;
wire  [2:0]  u4_col_out_869;
wire  [2:0]  u4_col_out_870;
wire  [2:0]  u4_col_out_871;
wire  [2:0]  u4_col_out_872;
wire  [2:0]  u4_col_out_873;
wire  [2:0]  u4_col_out_874;
wire  [2:0]  u4_col_out_875;
wire  [2:0]  u4_col_out_876;
wire  [2:0]  u4_col_out_877;
wire  [2:0]  u4_col_out_878;
wire  [2:0]  u4_col_out_879;
wire  [2:0]  u4_col_out_880;
wire  [2:0]  u4_col_out_881;
wire  [2:0]  u4_col_out_882;
wire  [2:0]  u4_col_out_883;
wire  [2:0]  u4_col_out_884;
wire  [2:0]  u4_col_out_885;
wire  [2:0]  u4_col_out_886;
wire  [2:0]  u4_col_out_887;
wire  [2:0]  u4_col_out_888;
wire  [2:0]  u4_col_out_889;
wire  [2:0]  u4_col_out_890;
wire  [2:0]  u4_col_out_891;
wire  [2:0]  u4_col_out_892;
wire  [2:0]  u4_col_out_893;
wire  [2:0]  u4_col_out_894;
wire  [2:0]  u4_col_out_895;
wire  [2:0]  u4_col_out_896;
wire  [2:0]  u4_col_out_897;
wire  [2:0]  u4_col_out_898;
wire  [2:0]  u4_col_out_899;
wire  [2:0]  u4_col_out_900;
wire  [2:0]  u4_col_out_901;
wire  [2:0]  u4_col_out_902;
wire  [2:0]  u4_col_out_903;
wire  [2:0]  u4_col_out_904;
wire  [2:0]  u4_col_out_905;
wire  [2:0]  u4_col_out_906;
wire  [2:0]  u4_col_out_907;
wire  [2:0]  u4_col_out_908;
wire  [2:0]  u4_col_out_909;
wire  [2:0]  u4_col_out_910;
wire  [2:0]  u4_col_out_911;
wire  [2:0]  u4_col_out_912;
wire  [2:0]  u4_col_out_913;
wire  [2:0]  u4_col_out_914;
wire  [2:0]  u4_col_out_915;
wire  [2:0]  u4_col_out_916;
wire  [2:0]  u4_col_out_917;
wire  [2:0]  u4_col_out_918;
wire  [2:0]  u4_col_out_919;
wire  [2:0]  u4_col_out_920;
wire  [2:0]  u4_col_out_921;
wire  [2:0]  u4_col_out_922;
wire  [2:0]  u4_col_out_923;
wire  [2:0]  u4_col_out_924;
wire  [2:0]  u4_col_out_925;
wire  [2:0]  u4_col_out_926;
wire  [2:0]  u4_col_out_927;
wire  [2:0]  u4_col_out_928;
wire  [2:0]  u4_col_out_929;
wire  [2:0]  u4_col_out_930;
wire  [2:0]  u4_col_out_931;
wire  [2:0]  u4_col_out_932;
wire  [2:0]  u4_col_out_933;
wire  [2:0]  u4_col_out_934;
wire  [2:0]  u4_col_out_935;
wire  [2:0]  u4_col_out_936;
wire  [2:0]  u4_col_out_937;
wire  [2:0]  u4_col_out_938;
wire  [2:0]  u4_col_out_939;
wire  [2:0]  u4_col_out_940;
wire  [2:0]  u4_col_out_941;
wire  [2:0]  u4_col_out_942;
wire  [2:0]  u4_col_out_943;
wire  [2:0]  u4_col_out_944;
wire  [2:0]  u4_col_out_945;
wire  [2:0]  u4_col_out_946;
wire  [2:0]  u4_col_out_947;
wire  [2:0]  u4_col_out_948;
wire  [2:0]  u4_col_out_949;
wire  [2:0]  u4_col_out_950;
wire  [2:0]  u4_col_out_951;
wire  [2:0]  u4_col_out_952;
wire  [2:0]  u4_col_out_953;
wire  [2:0]  u4_col_out_954;
wire  [2:0]  u4_col_out_955;
wire  [2:0]  u4_col_out_956;
wire  [2:0]  u4_col_out_957;
wire  [2:0]  u4_col_out_958;
wire  [2:0]  u4_col_out_959;
wire  [2:0]  u4_col_out_960;
wire  [2:0]  u4_col_out_961;
wire  [2:0]  u4_col_out_962;
wire  [2:0]  u4_col_out_963;
wire  [2:0]  u4_col_out_964;
wire  [2:0]  u4_col_out_965;
wire  [2:0]  u4_col_out_966;
wire  [2:0]  u4_col_out_967;
wire  [2:0]  u4_col_out_968;
wire  [2:0]  u4_col_out_969;
wire  [2:0]  u4_col_out_970;
wire  [2:0]  u4_col_out_971;
wire  [2:0]  u4_col_out_972;
wire  [2:0]  u4_col_out_973;
wire  [2:0]  u4_col_out_974;
wire  [2:0]  u4_col_out_975;
wire  [2:0]  u4_col_out_976;
wire  [2:0]  u4_col_out_977;
wire  [2:0]  u4_col_out_978;
wire  [2:0]  u4_col_out_979;
wire  [2:0]  u4_col_out_980;
wire  [2:0]  u4_col_out_981;
wire  [2:0]  u4_col_out_982;
wire  [2:0]  u4_col_out_983;
wire  [2:0]  u4_col_out_984;
wire  [2:0]  u4_col_out_985;
wire  [2:0]  u4_col_out_986;
wire  [2:0]  u4_col_out_987;
wire  [2:0]  u4_col_out_988;
wire  [2:0]  u4_col_out_989;
wire  [2:0]  u4_col_out_990;
wire  [2:0]  u4_col_out_991;
wire  [2:0]  u4_col_out_992;
wire  [2:0]  u4_col_out_993;
wire  [2:0]  u4_col_out_994;
wire  [2:0]  u4_col_out_995;
wire  [2:0]  u4_col_out_996;
wire  [2:0]  u4_col_out_997;
wire  [2:0]  u4_col_out_998;
wire  [2:0]  u4_col_out_999;
wire  [2:0]  u4_col_out_1000;
wire  [2:0]  u4_col_out_1001;
wire  [2:0]  u4_col_out_1002;
wire  [2:0]  u4_col_out_1003;
wire  [2:0]  u4_col_out_1004;
wire  [2:0]  u4_col_out_1005;
wire  [2:0]  u4_col_out_1006;
wire  [2:0]  u4_col_out_1007;
wire  [2:0]  u4_col_out_1008;
wire  [2:0]  u4_col_out_1009;
wire  [2:0]  u4_col_out_1010;
wire  [2:0]  u4_col_out_1011;
wire  [2:0]  u4_col_out_1012;
wire  [2:0]  u4_col_out_1013;
wire  [2:0]  u4_col_out_1014;
wire  [2:0]  u4_col_out_1015;
wire  [2:0]  u4_col_out_1016;
wire  [2:0]  u4_col_out_1017;
wire  [2:0]  u4_col_out_1018;
wire  [2:0]  u4_col_out_1019;
wire  [2:0]  u4_col_out_1020;
wire  [2:0]  u4_col_out_1021;
wire  [2:0]  u4_col_out_1022;
wire  [2:0]  u4_col_out_1023;
wire  [2:0]  u4_col_out_1024;
wire  [2:0]  u4_col_out_1025;
wire  [2:0]  u4_col_out_1026;
wire  [2:0]  u4_col_out_1027;
wire  [2:0]  u4_col_out_1028;
wire  [2:0]  u4_col_out_1029;
wire  [2:0]  u4_col_out_1030;
wire  [2:0]  u4_col_out_1031;
wire  [2:0]  u4_col_out_1032;
wire  [2:0]  u4_col_out_1033;

compressor_array_4_3_1033  u4_compressor_array_4_3_1033 (
    .col_in_0                ( u3_col_out_0       ),
    .col_in_1                ( u3_col_out_1       ),
    .col_in_2                ( u3_col_out_2       ),
    .col_in_3                ( u3_col_out_3       ),
    .col_in_4                ( u3_col_out_4       ),
    .col_in_5                ( u3_col_out_5       ),
    .col_in_6                ( u3_col_out_6       ),
    .col_in_7                ( u3_col_out_7       ),
    .col_in_8                ( u3_col_out_8       ),
    .col_in_9                ( u3_col_out_9       ),
    .col_in_10               ( u3_col_out_10      ),
    .col_in_11               ( u3_col_out_11      ),
    .col_in_12               ( u3_col_out_12      ),
    .col_in_13               ( u3_col_out_13      ),
    .col_in_14               ( u3_col_out_14      ),
    .col_in_15               ( u3_col_out_15      ),
    .col_in_16               ( u3_col_out_16      ),
    .col_in_17               ( u3_col_out_17      ),
    .col_in_18               ( u3_col_out_18      ),
    .col_in_19               ( u3_col_out_19      ),
    .col_in_20               ( u3_col_out_20      ),
    .col_in_21               ( u3_col_out_21      ),
    .col_in_22               ( u3_col_out_22      ),
    .col_in_23               ( u3_col_out_23      ),
    .col_in_24               ( u3_col_out_24      ),
    .col_in_25               ( u3_col_out_25      ),
    .col_in_26               ( u3_col_out_26      ),
    .col_in_27               ( u3_col_out_27      ),
    .col_in_28               ( u3_col_out_28      ),
    .col_in_29               ( u3_col_out_29      ),
    .col_in_30               ( u3_col_out_30      ),
    .col_in_31               ( u3_col_out_31      ),
    .col_in_32               ( u3_col_out_32      ),
    .col_in_33               ( u3_col_out_33      ),
    .col_in_34               ( u3_col_out_34      ),
    .col_in_35               ( u3_col_out_35      ),
    .col_in_36               ( u3_col_out_36      ),
    .col_in_37               ( u3_col_out_37      ),
    .col_in_38               ( u3_col_out_38      ),
    .col_in_39               ( u3_col_out_39      ),
    .col_in_40               ( u3_col_out_40      ),
    .col_in_41               ( u3_col_out_41      ),
    .col_in_42               ( u3_col_out_42      ),
    .col_in_43               ( u3_col_out_43      ),
    .col_in_44               ( u3_col_out_44      ),
    .col_in_45               ( u3_col_out_45      ),
    .col_in_46               ( u3_col_out_46      ),
    .col_in_47               ( u3_col_out_47      ),
    .col_in_48               ( u3_col_out_48      ),
    .col_in_49               ( u3_col_out_49      ),
    .col_in_50               ( u3_col_out_50      ),
    .col_in_51               ( u3_col_out_51      ),
    .col_in_52               ( u3_col_out_52      ),
    .col_in_53               ( u3_col_out_53      ),
    .col_in_54               ( u3_col_out_54      ),
    .col_in_55               ( u3_col_out_55      ),
    .col_in_56               ( u3_col_out_56      ),
    .col_in_57               ( u3_col_out_57      ),
    .col_in_58               ( u3_col_out_58      ),
    .col_in_59               ( u3_col_out_59      ),
    .col_in_60               ( u3_col_out_60      ),
    .col_in_61               ( u3_col_out_61      ),
    .col_in_62               ( u3_col_out_62      ),
    .col_in_63               ( u3_col_out_63      ),
    .col_in_64               ( u3_col_out_64      ),
    .col_in_65               ( u3_col_out_65      ),
    .col_in_66               ( u3_col_out_66      ),
    .col_in_67               ( u3_col_out_67      ),
    .col_in_68               ( u3_col_out_68      ),
    .col_in_69               ( u3_col_out_69      ),
    .col_in_70               ( u3_col_out_70      ),
    .col_in_71               ( u3_col_out_71      ),
    .col_in_72               ( u3_col_out_72      ),
    .col_in_73               ( u3_col_out_73      ),
    .col_in_74               ( u3_col_out_74      ),
    .col_in_75               ( u3_col_out_75      ),
    .col_in_76               ( u3_col_out_76      ),
    .col_in_77               ( u3_col_out_77      ),
    .col_in_78               ( u3_col_out_78      ),
    .col_in_79               ( u3_col_out_79      ),
    .col_in_80               ( u3_col_out_80      ),
    .col_in_81               ( u3_col_out_81      ),
    .col_in_82               ( u3_col_out_82      ),
    .col_in_83               ( u3_col_out_83      ),
    .col_in_84               ( u3_col_out_84      ),
    .col_in_85               ( u3_col_out_85      ),
    .col_in_86               ( u3_col_out_86      ),
    .col_in_87               ( u3_col_out_87      ),
    .col_in_88               ( u3_col_out_88      ),
    .col_in_89               ( u3_col_out_89      ),
    .col_in_90               ( u3_col_out_90      ),
    .col_in_91               ( u3_col_out_91      ),
    .col_in_92               ( u3_col_out_92      ),
    .col_in_93               ( u3_col_out_93      ),
    .col_in_94               ( u3_col_out_94      ),
    .col_in_95               ( u3_col_out_95      ),
    .col_in_96               ( u3_col_out_96      ),
    .col_in_97               ( u3_col_out_97      ),
    .col_in_98               ( u3_col_out_98      ),
    .col_in_99               ( u3_col_out_99      ),
    .col_in_100              ( u3_col_out_100     ),
    .col_in_101              ( u3_col_out_101     ),
    .col_in_102              ( u3_col_out_102     ),
    .col_in_103              ( u3_col_out_103     ),
    .col_in_104              ( u3_col_out_104     ),
    .col_in_105              ( u3_col_out_105     ),
    .col_in_106              ( u3_col_out_106     ),
    .col_in_107              ( u3_col_out_107     ),
    .col_in_108              ( u3_col_out_108     ),
    .col_in_109              ( u3_col_out_109     ),
    .col_in_110              ( u3_col_out_110     ),
    .col_in_111              ( u3_col_out_111     ),
    .col_in_112              ( u3_col_out_112     ),
    .col_in_113              ( u3_col_out_113     ),
    .col_in_114              ( u3_col_out_114     ),
    .col_in_115              ( u3_col_out_115     ),
    .col_in_116              ( u3_col_out_116     ),
    .col_in_117              ( u3_col_out_117     ),
    .col_in_118              ( u3_col_out_118     ),
    .col_in_119              ( u3_col_out_119     ),
    .col_in_120              ( u3_col_out_120     ),
    .col_in_121              ( u3_col_out_121     ),
    .col_in_122              ( u3_col_out_122     ),
    .col_in_123              ( u3_col_out_123     ),
    .col_in_124              ( u3_col_out_124     ),
    .col_in_125              ( u3_col_out_125     ),
    .col_in_126              ( u3_col_out_126     ),
    .col_in_127              ( u3_col_out_127     ),
    .col_in_128              ( u3_col_out_128     ),
    .col_in_129              ( u3_col_out_129     ),
    .col_in_130              ( u3_col_out_130     ),
    .col_in_131              ( u3_col_out_131     ),
    .col_in_132              ( u3_col_out_132     ),
    .col_in_133              ( u3_col_out_133     ),
    .col_in_134              ( u3_col_out_134     ),
    .col_in_135              ( u3_col_out_135     ),
    .col_in_136              ( u3_col_out_136     ),
    .col_in_137              ( u3_col_out_137     ),
    .col_in_138              ( u3_col_out_138     ),
    .col_in_139              ( u3_col_out_139     ),
    .col_in_140              ( u3_col_out_140     ),
    .col_in_141              ( u3_col_out_141     ),
    .col_in_142              ( u3_col_out_142     ),
    .col_in_143              ( u3_col_out_143     ),
    .col_in_144              ( u3_col_out_144     ),
    .col_in_145              ( u3_col_out_145     ),
    .col_in_146              ( u3_col_out_146     ),
    .col_in_147              ( u3_col_out_147     ),
    .col_in_148              ( u3_col_out_148     ),
    .col_in_149              ( u3_col_out_149     ),
    .col_in_150              ( u3_col_out_150     ),
    .col_in_151              ( u3_col_out_151     ),
    .col_in_152              ( u3_col_out_152     ),
    .col_in_153              ( u3_col_out_153     ),
    .col_in_154              ( u3_col_out_154     ),
    .col_in_155              ( u3_col_out_155     ),
    .col_in_156              ( u3_col_out_156     ),
    .col_in_157              ( u3_col_out_157     ),
    .col_in_158              ( u3_col_out_158     ),
    .col_in_159              ( u3_col_out_159     ),
    .col_in_160              ( u3_col_out_160     ),
    .col_in_161              ( u3_col_out_161     ),
    .col_in_162              ( u3_col_out_162     ),
    .col_in_163              ( u3_col_out_163     ),
    .col_in_164              ( u3_col_out_164     ),
    .col_in_165              ( u3_col_out_165     ),
    .col_in_166              ( u3_col_out_166     ),
    .col_in_167              ( u3_col_out_167     ),
    .col_in_168              ( u3_col_out_168     ),
    .col_in_169              ( u3_col_out_169     ),
    .col_in_170              ( u3_col_out_170     ),
    .col_in_171              ( u3_col_out_171     ),
    .col_in_172              ( u3_col_out_172     ),
    .col_in_173              ( u3_col_out_173     ),
    .col_in_174              ( u3_col_out_174     ),
    .col_in_175              ( u3_col_out_175     ),
    .col_in_176              ( u3_col_out_176     ),
    .col_in_177              ( u3_col_out_177     ),
    .col_in_178              ( u3_col_out_178     ),
    .col_in_179              ( u3_col_out_179     ),
    .col_in_180              ( u3_col_out_180     ),
    .col_in_181              ( u3_col_out_181     ),
    .col_in_182              ( u3_col_out_182     ),
    .col_in_183              ( u3_col_out_183     ),
    .col_in_184              ( u3_col_out_184     ),
    .col_in_185              ( u3_col_out_185     ),
    .col_in_186              ( u3_col_out_186     ),
    .col_in_187              ( u3_col_out_187     ),
    .col_in_188              ( u3_col_out_188     ),
    .col_in_189              ( u3_col_out_189     ),
    .col_in_190              ( u3_col_out_190     ),
    .col_in_191              ( u3_col_out_191     ),
    .col_in_192              ( u3_col_out_192     ),
    .col_in_193              ( u3_col_out_193     ),
    .col_in_194              ( u3_col_out_194     ),
    .col_in_195              ( u3_col_out_195     ),
    .col_in_196              ( u3_col_out_196     ),
    .col_in_197              ( u3_col_out_197     ),
    .col_in_198              ( u3_col_out_198     ),
    .col_in_199              ( u3_col_out_199     ),
    .col_in_200              ( u3_col_out_200     ),
    .col_in_201              ( u3_col_out_201     ),
    .col_in_202              ( u3_col_out_202     ),
    .col_in_203              ( u3_col_out_203     ),
    .col_in_204              ( u3_col_out_204     ),
    .col_in_205              ( u3_col_out_205     ),
    .col_in_206              ( u3_col_out_206     ),
    .col_in_207              ( u3_col_out_207     ),
    .col_in_208              ( u3_col_out_208     ),
    .col_in_209              ( u3_col_out_209     ),
    .col_in_210              ( u3_col_out_210     ),
    .col_in_211              ( u3_col_out_211     ),
    .col_in_212              ( u3_col_out_212     ),
    .col_in_213              ( u3_col_out_213     ),
    .col_in_214              ( u3_col_out_214     ),
    .col_in_215              ( u3_col_out_215     ),
    .col_in_216              ( u3_col_out_216     ),
    .col_in_217              ( u3_col_out_217     ),
    .col_in_218              ( u3_col_out_218     ),
    .col_in_219              ( u3_col_out_219     ),
    .col_in_220              ( u3_col_out_220     ),
    .col_in_221              ( u3_col_out_221     ),
    .col_in_222              ( u3_col_out_222     ),
    .col_in_223              ( u3_col_out_223     ),
    .col_in_224              ( u3_col_out_224     ),
    .col_in_225              ( u3_col_out_225     ),
    .col_in_226              ( u3_col_out_226     ),
    .col_in_227              ( u3_col_out_227     ),
    .col_in_228              ( u3_col_out_228     ),
    .col_in_229              ( u3_col_out_229     ),
    .col_in_230              ( u3_col_out_230     ),
    .col_in_231              ( u3_col_out_231     ),
    .col_in_232              ( u3_col_out_232     ),
    .col_in_233              ( u3_col_out_233     ),
    .col_in_234              ( u3_col_out_234     ),
    .col_in_235              ( u3_col_out_235     ),
    .col_in_236              ( u3_col_out_236     ),
    .col_in_237              ( u3_col_out_237     ),
    .col_in_238              ( u3_col_out_238     ),
    .col_in_239              ( u3_col_out_239     ),
    .col_in_240              ( u3_col_out_240     ),
    .col_in_241              ( u3_col_out_241     ),
    .col_in_242              ( u3_col_out_242     ),
    .col_in_243              ( u3_col_out_243     ),
    .col_in_244              ( u3_col_out_244     ),
    .col_in_245              ( u3_col_out_245     ),
    .col_in_246              ( u3_col_out_246     ),
    .col_in_247              ( u3_col_out_247     ),
    .col_in_248              ( u3_col_out_248     ),
    .col_in_249              ( u3_col_out_249     ),
    .col_in_250              ( u3_col_out_250     ),
    .col_in_251              ( u3_col_out_251     ),
    .col_in_252              ( u3_col_out_252     ),
    .col_in_253              ( u3_col_out_253     ),
    .col_in_254              ( u3_col_out_254     ),
    .col_in_255              ( u3_col_out_255     ),
    .col_in_256              ( u3_col_out_256     ),
    .col_in_257              ( u3_col_out_257     ),
    .col_in_258              ( u3_col_out_258     ),
    .col_in_259              ( u3_col_out_259     ),
    .col_in_260              ( u3_col_out_260     ),
    .col_in_261              ( u3_col_out_261     ),
    .col_in_262              ( u3_col_out_262     ),
    .col_in_263              ( u3_col_out_263     ),
    .col_in_264              ( u3_col_out_264     ),
    .col_in_265              ( u3_col_out_265     ),
    .col_in_266              ( u3_col_out_266     ),
    .col_in_267              ( u3_col_out_267     ),
    .col_in_268              ( u3_col_out_268     ),
    .col_in_269              ( u3_col_out_269     ),
    .col_in_270              ( u3_col_out_270     ),
    .col_in_271              ( u3_col_out_271     ),
    .col_in_272              ( u3_col_out_272     ),
    .col_in_273              ( u3_col_out_273     ),
    .col_in_274              ( u3_col_out_274     ),
    .col_in_275              ( u3_col_out_275     ),
    .col_in_276              ( u3_col_out_276     ),
    .col_in_277              ( u3_col_out_277     ),
    .col_in_278              ( u3_col_out_278     ),
    .col_in_279              ( u3_col_out_279     ),
    .col_in_280              ( u3_col_out_280     ),
    .col_in_281              ( u3_col_out_281     ),
    .col_in_282              ( u3_col_out_282     ),
    .col_in_283              ( u3_col_out_283     ),
    .col_in_284              ( u3_col_out_284     ),
    .col_in_285              ( u3_col_out_285     ),
    .col_in_286              ( u3_col_out_286     ),
    .col_in_287              ( u3_col_out_287     ),
    .col_in_288              ( u3_col_out_288     ),
    .col_in_289              ( u3_col_out_289     ),
    .col_in_290              ( u3_col_out_290     ),
    .col_in_291              ( u3_col_out_291     ),
    .col_in_292              ( u3_col_out_292     ),
    .col_in_293              ( u3_col_out_293     ),
    .col_in_294              ( u3_col_out_294     ),
    .col_in_295              ( u3_col_out_295     ),
    .col_in_296              ( u3_col_out_296     ),
    .col_in_297              ( u3_col_out_297     ),
    .col_in_298              ( u3_col_out_298     ),
    .col_in_299              ( u3_col_out_299     ),
    .col_in_300              ( u3_col_out_300     ),
    .col_in_301              ( u3_col_out_301     ),
    .col_in_302              ( u3_col_out_302     ),
    .col_in_303              ( u3_col_out_303     ),
    .col_in_304              ( u3_col_out_304     ),
    .col_in_305              ( u3_col_out_305     ),
    .col_in_306              ( u3_col_out_306     ),
    .col_in_307              ( u3_col_out_307     ),
    .col_in_308              ( u3_col_out_308     ),
    .col_in_309              ( u3_col_out_309     ),
    .col_in_310              ( u3_col_out_310     ),
    .col_in_311              ( u3_col_out_311     ),
    .col_in_312              ( u3_col_out_312     ),
    .col_in_313              ( u3_col_out_313     ),
    .col_in_314              ( u3_col_out_314     ),
    .col_in_315              ( u3_col_out_315     ),
    .col_in_316              ( u3_col_out_316     ),
    .col_in_317              ( u3_col_out_317     ),
    .col_in_318              ( u3_col_out_318     ),
    .col_in_319              ( u3_col_out_319     ),
    .col_in_320              ( u3_col_out_320     ),
    .col_in_321              ( u3_col_out_321     ),
    .col_in_322              ( u3_col_out_322     ),
    .col_in_323              ( u3_col_out_323     ),
    .col_in_324              ( u3_col_out_324     ),
    .col_in_325              ( u3_col_out_325     ),
    .col_in_326              ( u3_col_out_326     ),
    .col_in_327              ( u3_col_out_327     ),
    .col_in_328              ( u3_col_out_328     ),
    .col_in_329              ( u3_col_out_329     ),
    .col_in_330              ( u3_col_out_330     ),
    .col_in_331              ( u3_col_out_331     ),
    .col_in_332              ( u3_col_out_332     ),
    .col_in_333              ( u3_col_out_333     ),
    .col_in_334              ( u3_col_out_334     ),
    .col_in_335              ( u3_col_out_335     ),
    .col_in_336              ( u3_col_out_336     ),
    .col_in_337              ( u3_col_out_337     ),
    .col_in_338              ( u3_col_out_338     ),
    .col_in_339              ( u3_col_out_339     ),
    .col_in_340              ( u3_col_out_340     ),
    .col_in_341              ( u3_col_out_341     ),
    .col_in_342              ( u3_col_out_342     ),
    .col_in_343              ( u3_col_out_343     ),
    .col_in_344              ( u3_col_out_344     ),
    .col_in_345              ( u3_col_out_345     ),
    .col_in_346              ( u3_col_out_346     ),
    .col_in_347              ( u3_col_out_347     ),
    .col_in_348              ( u3_col_out_348     ),
    .col_in_349              ( u3_col_out_349     ),
    .col_in_350              ( u3_col_out_350     ),
    .col_in_351              ( u3_col_out_351     ),
    .col_in_352              ( u3_col_out_352     ),
    .col_in_353              ( u3_col_out_353     ),
    .col_in_354              ( u3_col_out_354     ),
    .col_in_355              ( u3_col_out_355     ),
    .col_in_356              ( u3_col_out_356     ),
    .col_in_357              ( u3_col_out_357     ),
    .col_in_358              ( u3_col_out_358     ),
    .col_in_359              ( u3_col_out_359     ),
    .col_in_360              ( u3_col_out_360     ),
    .col_in_361              ( u3_col_out_361     ),
    .col_in_362              ( u3_col_out_362     ),
    .col_in_363              ( u3_col_out_363     ),
    .col_in_364              ( u3_col_out_364     ),
    .col_in_365              ( u3_col_out_365     ),
    .col_in_366              ( u3_col_out_366     ),
    .col_in_367              ( u3_col_out_367     ),
    .col_in_368              ( u3_col_out_368     ),
    .col_in_369              ( u3_col_out_369     ),
    .col_in_370              ( u3_col_out_370     ),
    .col_in_371              ( u3_col_out_371     ),
    .col_in_372              ( u3_col_out_372     ),
    .col_in_373              ( u3_col_out_373     ),
    .col_in_374              ( u3_col_out_374     ),
    .col_in_375              ( u3_col_out_375     ),
    .col_in_376              ( u3_col_out_376     ),
    .col_in_377              ( u3_col_out_377     ),
    .col_in_378              ( u3_col_out_378     ),
    .col_in_379              ( u3_col_out_379     ),
    .col_in_380              ( u3_col_out_380     ),
    .col_in_381              ( u3_col_out_381     ),
    .col_in_382              ( u3_col_out_382     ),
    .col_in_383              ( u3_col_out_383     ),
    .col_in_384              ( u3_col_out_384     ),
    .col_in_385              ( u3_col_out_385     ),
    .col_in_386              ( u3_col_out_386     ),
    .col_in_387              ( u3_col_out_387     ),
    .col_in_388              ( u3_col_out_388     ),
    .col_in_389              ( u3_col_out_389     ),
    .col_in_390              ( u3_col_out_390     ),
    .col_in_391              ( u3_col_out_391     ),
    .col_in_392              ( u3_col_out_392     ),
    .col_in_393              ( u3_col_out_393     ),
    .col_in_394              ( u3_col_out_394     ),
    .col_in_395              ( u3_col_out_395     ),
    .col_in_396              ( u3_col_out_396     ),
    .col_in_397              ( u3_col_out_397     ),
    .col_in_398              ( u3_col_out_398     ),
    .col_in_399              ( u3_col_out_399     ),
    .col_in_400              ( u3_col_out_400     ),
    .col_in_401              ( u3_col_out_401     ),
    .col_in_402              ( u3_col_out_402     ),
    .col_in_403              ( u3_col_out_403     ),
    .col_in_404              ( u3_col_out_404     ),
    .col_in_405              ( u3_col_out_405     ),
    .col_in_406              ( u3_col_out_406     ),
    .col_in_407              ( u3_col_out_407     ),
    .col_in_408              ( u3_col_out_408     ),
    .col_in_409              ( u3_col_out_409     ),
    .col_in_410              ( u3_col_out_410     ),
    .col_in_411              ( u3_col_out_411     ),
    .col_in_412              ( u3_col_out_412     ),
    .col_in_413              ( u3_col_out_413     ),
    .col_in_414              ( u3_col_out_414     ),
    .col_in_415              ( u3_col_out_415     ),
    .col_in_416              ( u3_col_out_416     ),
    .col_in_417              ( u3_col_out_417     ),
    .col_in_418              ( u3_col_out_418     ),
    .col_in_419              ( u3_col_out_419     ),
    .col_in_420              ( u3_col_out_420     ),
    .col_in_421              ( u3_col_out_421     ),
    .col_in_422              ( u3_col_out_422     ),
    .col_in_423              ( u3_col_out_423     ),
    .col_in_424              ( u3_col_out_424     ),
    .col_in_425              ( u3_col_out_425     ),
    .col_in_426              ( u3_col_out_426     ),
    .col_in_427              ( u3_col_out_427     ),
    .col_in_428              ( u3_col_out_428     ),
    .col_in_429              ( u3_col_out_429     ),
    .col_in_430              ( u3_col_out_430     ),
    .col_in_431              ( u3_col_out_431     ),
    .col_in_432              ( u3_col_out_432     ),
    .col_in_433              ( u3_col_out_433     ),
    .col_in_434              ( u3_col_out_434     ),
    .col_in_435              ( u3_col_out_435     ),
    .col_in_436              ( u3_col_out_436     ),
    .col_in_437              ( u3_col_out_437     ),
    .col_in_438              ( u3_col_out_438     ),
    .col_in_439              ( u3_col_out_439     ),
    .col_in_440              ( u3_col_out_440     ),
    .col_in_441              ( u3_col_out_441     ),
    .col_in_442              ( u3_col_out_442     ),
    .col_in_443              ( u3_col_out_443     ),
    .col_in_444              ( u3_col_out_444     ),
    .col_in_445              ( u3_col_out_445     ),
    .col_in_446              ( u3_col_out_446     ),
    .col_in_447              ( u3_col_out_447     ),
    .col_in_448              ( u3_col_out_448     ),
    .col_in_449              ( u3_col_out_449     ),
    .col_in_450              ( u3_col_out_450     ),
    .col_in_451              ( u3_col_out_451     ),
    .col_in_452              ( u3_col_out_452     ),
    .col_in_453              ( u3_col_out_453     ),
    .col_in_454              ( u3_col_out_454     ),
    .col_in_455              ( u3_col_out_455     ),
    .col_in_456              ( u3_col_out_456     ),
    .col_in_457              ( u3_col_out_457     ),
    .col_in_458              ( u3_col_out_458     ),
    .col_in_459              ( u3_col_out_459     ),
    .col_in_460              ( u3_col_out_460     ),
    .col_in_461              ( u3_col_out_461     ),
    .col_in_462              ( u3_col_out_462     ),
    .col_in_463              ( u3_col_out_463     ),
    .col_in_464              ( u3_col_out_464     ),
    .col_in_465              ( u3_col_out_465     ),
    .col_in_466              ( u3_col_out_466     ),
    .col_in_467              ( u3_col_out_467     ),
    .col_in_468              ( u3_col_out_468     ),
    .col_in_469              ( u3_col_out_469     ),
    .col_in_470              ( u3_col_out_470     ),
    .col_in_471              ( u3_col_out_471     ),
    .col_in_472              ( u3_col_out_472     ),
    .col_in_473              ( u3_col_out_473     ),
    .col_in_474              ( u3_col_out_474     ),
    .col_in_475              ( u3_col_out_475     ),
    .col_in_476              ( u3_col_out_476     ),
    .col_in_477              ( u3_col_out_477     ),
    .col_in_478              ( u3_col_out_478     ),
    .col_in_479              ( u3_col_out_479     ),
    .col_in_480              ( u3_col_out_480     ),
    .col_in_481              ( u3_col_out_481     ),
    .col_in_482              ( u3_col_out_482     ),
    .col_in_483              ( u3_col_out_483     ),
    .col_in_484              ( u3_col_out_484     ),
    .col_in_485              ( u3_col_out_485     ),
    .col_in_486              ( u3_col_out_486     ),
    .col_in_487              ( u3_col_out_487     ),
    .col_in_488              ( u3_col_out_488     ),
    .col_in_489              ( u3_col_out_489     ),
    .col_in_490              ( u3_col_out_490     ),
    .col_in_491              ( u3_col_out_491     ),
    .col_in_492              ( u3_col_out_492     ),
    .col_in_493              ( u3_col_out_493     ),
    .col_in_494              ( u3_col_out_494     ),
    .col_in_495              ( u3_col_out_495     ),
    .col_in_496              ( u3_col_out_496     ),
    .col_in_497              ( u3_col_out_497     ),
    .col_in_498              ( u3_col_out_498     ),
    .col_in_499              ( u3_col_out_499     ),
    .col_in_500              ( u3_col_out_500     ),
    .col_in_501              ( u3_col_out_501     ),
    .col_in_502              ( u3_col_out_502     ),
    .col_in_503              ( u3_col_out_503     ),
    .col_in_504              ( u3_col_out_504     ),
    .col_in_505              ( u3_col_out_505     ),
    .col_in_506              ( u3_col_out_506     ),
    .col_in_507              ( u3_col_out_507     ),
    .col_in_508              ( u3_col_out_508     ),
    .col_in_509              ( u3_col_out_509     ),
    .col_in_510              ( u3_col_out_510     ),
    .col_in_511              ( u3_col_out_511     ),
    .col_in_512              ( u3_col_out_512     ),
    .col_in_513              ( u3_col_out_513     ),
    .col_in_514              ( u3_col_out_514     ),
    .col_in_515              ( u3_col_out_515     ),
    .col_in_516              ( u3_col_out_516     ),
    .col_in_517              ( u3_col_out_517     ),
    .col_in_518              ( u3_col_out_518     ),
    .col_in_519              ( u3_col_out_519     ),
    .col_in_520              ( u3_col_out_520     ),
    .col_in_521              ( u3_col_out_521     ),
    .col_in_522              ( u3_col_out_522     ),
    .col_in_523              ( u3_col_out_523     ),
    .col_in_524              ( u3_col_out_524     ),
    .col_in_525              ( u3_col_out_525     ),
    .col_in_526              ( u3_col_out_526     ),
    .col_in_527              ( u3_col_out_527     ),
    .col_in_528              ( u3_col_out_528     ),
    .col_in_529              ( u3_col_out_529     ),
    .col_in_530              ( u3_col_out_530     ),
    .col_in_531              ( u3_col_out_531     ),
    .col_in_532              ( u3_col_out_532     ),
    .col_in_533              ( u3_col_out_533     ),
    .col_in_534              ( u3_col_out_534     ),
    .col_in_535              ( u3_col_out_535     ),
    .col_in_536              ( u3_col_out_536     ),
    .col_in_537              ( u3_col_out_537     ),
    .col_in_538              ( u3_col_out_538     ),
    .col_in_539              ( u3_col_out_539     ),
    .col_in_540              ( u3_col_out_540     ),
    .col_in_541              ( u3_col_out_541     ),
    .col_in_542              ( u3_col_out_542     ),
    .col_in_543              ( u3_col_out_543     ),
    .col_in_544              ( u3_col_out_544     ),
    .col_in_545              ( u3_col_out_545     ),
    .col_in_546              ( u3_col_out_546     ),
    .col_in_547              ( u3_col_out_547     ),
    .col_in_548              ( u3_col_out_548     ),
    .col_in_549              ( u3_col_out_549     ),
    .col_in_550              ( u3_col_out_550     ),
    .col_in_551              ( u3_col_out_551     ),
    .col_in_552              ( u3_col_out_552     ),
    .col_in_553              ( u3_col_out_553     ),
    .col_in_554              ( u3_col_out_554     ),
    .col_in_555              ( u3_col_out_555     ),
    .col_in_556              ( u3_col_out_556     ),
    .col_in_557              ( u3_col_out_557     ),
    .col_in_558              ( u3_col_out_558     ),
    .col_in_559              ( u3_col_out_559     ),
    .col_in_560              ( u3_col_out_560     ),
    .col_in_561              ( u3_col_out_561     ),
    .col_in_562              ( u3_col_out_562     ),
    .col_in_563              ( u3_col_out_563     ),
    .col_in_564              ( u3_col_out_564     ),
    .col_in_565              ( u3_col_out_565     ),
    .col_in_566              ( u3_col_out_566     ),
    .col_in_567              ( u3_col_out_567     ),
    .col_in_568              ( u3_col_out_568     ),
    .col_in_569              ( u3_col_out_569     ),
    .col_in_570              ( u3_col_out_570     ),
    .col_in_571              ( u3_col_out_571     ),
    .col_in_572              ( u3_col_out_572     ),
    .col_in_573              ( u3_col_out_573     ),
    .col_in_574              ( u3_col_out_574     ),
    .col_in_575              ( u3_col_out_575     ),
    .col_in_576              ( u3_col_out_576     ),
    .col_in_577              ( u3_col_out_577     ),
    .col_in_578              ( u3_col_out_578     ),
    .col_in_579              ( u3_col_out_579     ),
    .col_in_580              ( u3_col_out_580     ),
    .col_in_581              ( u3_col_out_581     ),
    .col_in_582              ( u3_col_out_582     ),
    .col_in_583              ( u3_col_out_583     ),
    .col_in_584              ( u3_col_out_584     ),
    .col_in_585              ( u3_col_out_585     ),
    .col_in_586              ( u3_col_out_586     ),
    .col_in_587              ( u3_col_out_587     ),
    .col_in_588              ( u3_col_out_588     ),
    .col_in_589              ( u3_col_out_589     ),
    .col_in_590              ( u3_col_out_590     ),
    .col_in_591              ( u3_col_out_591     ),
    .col_in_592              ( u3_col_out_592     ),
    .col_in_593              ( u3_col_out_593     ),
    .col_in_594              ( u3_col_out_594     ),
    .col_in_595              ( u3_col_out_595     ),
    .col_in_596              ( u3_col_out_596     ),
    .col_in_597              ( u3_col_out_597     ),
    .col_in_598              ( u3_col_out_598     ),
    .col_in_599              ( u3_col_out_599     ),
    .col_in_600              ( u3_col_out_600     ),
    .col_in_601              ( u3_col_out_601     ),
    .col_in_602              ( u3_col_out_602     ),
    .col_in_603              ( u3_col_out_603     ),
    .col_in_604              ( u3_col_out_604     ),
    .col_in_605              ( u3_col_out_605     ),
    .col_in_606              ( u3_col_out_606     ),
    .col_in_607              ( u3_col_out_607     ),
    .col_in_608              ( u3_col_out_608     ),
    .col_in_609              ( u3_col_out_609     ),
    .col_in_610              ( u3_col_out_610     ),
    .col_in_611              ( u3_col_out_611     ),
    .col_in_612              ( u3_col_out_612     ),
    .col_in_613              ( u3_col_out_613     ),
    .col_in_614              ( u3_col_out_614     ),
    .col_in_615              ( u3_col_out_615     ),
    .col_in_616              ( u3_col_out_616     ),
    .col_in_617              ( u3_col_out_617     ),
    .col_in_618              ( u3_col_out_618     ),
    .col_in_619              ( u3_col_out_619     ),
    .col_in_620              ( u3_col_out_620     ),
    .col_in_621              ( u3_col_out_621     ),
    .col_in_622              ( u3_col_out_622     ),
    .col_in_623              ( u3_col_out_623     ),
    .col_in_624              ( u3_col_out_624     ),
    .col_in_625              ( u3_col_out_625     ),
    .col_in_626              ( u3_col_out_626     ),
    .col_in_627              ( u3_col_out_627     ),
    .col_in_628              ( u3_col_out_628     ),
    .col_in_629              ( u3_col_out_629     ),
    .col_in_630              ( u3_col_out_630     ),
    .col_in_631              ( u3_col_out_631     ),
    .col_in_632              ( u3_col_out_632     ),
    .col_in_633              ( u3_col_out_633     ),
    .col_in_634              ( u3_col_out_634     ),
    .col_in_635              ( u3_col_out_635     ),
    .col_in_636              ( u3_col_out_636     ),
    .col_in_637              ( u3_col_out_637     ),
    .col_in_638              ( u3_col_out_638     ),
    .col_in_639              ( u3_col_out_639     ),
    .col_in_640              ( u3_col_out_640     ),
    .col_in_641              ( u3_col_out_641     ),
    .col_in_642              ( u3_col_out_642     ),
    .col_in_643              ( u3_col_out_643     ),
    .col_in_644              ( u3_col_out_644     ),
    .col_in_645              ( u3_col_out_645     ),
    .col_in_646              ( u3_col_out_646     ),
    .col_in_647              ( u3_col_out_647     ),
    .col_in_648              ( u3_col_out_648     ),
    .col_in_649              ( u3_col_out_649     ),
    .col_in_650              ( u3_col_out_650     ),
    .col_in_651              ( u3_col_out_651     ),
    .col_in_652              ( u3_col_out_652     ),
    .col_in_653              ( u3_col_out_653     ),
    .col_in_654              ( u3_col_out_654     ),
    .col_in_655              ( u3_col_out_655     ),
    .col_in_656              ( u3_col_out_656     ),
    .col_in_657              ( u3_col_out_657     ),
    .col_in_658              ( u3_col_out_658     ),
    .col_in_659              ( u3_col_out_659     ),
    .col_in_660              ( u3_col_out_660     ),
    .col_in_661              ( u3_col_out_661     ),
    .col_in_662              ( u3_col_out_662     ),
    .col_in_663              ( u3_col_out_663     ),
    .col_in_664              ( u3_col_out_664     ),
    .col_in_665              ( u3_col_out_665     ),
    .col_in_666              ( u3_col_out_666     ),
    .col_in_667              ( u3_col_out_667     ),
    .col_in_668              ( u3_col_out_668     ),
    .col_in_669              ( u3_col_out_669     ),
    .col_in_670              ( u3_col_out_670     ),
    .col_in_671              ( u3_col_out_671     ),
    .col_in_672              ( u3_col_out_672     ),
    .col_in_673              ( u3_col_out_673     ),
    .col_in_674              ( u3_col_out_674     ),
    .col_in_675              ( u3_col_out_675     ),
    .col_in_676              ( u3_col_out_676     ),
    .col_in_677              ( u3_col_out_677     ),
    .col_in_678              ( u3_col_out_678     ),
    .col_in_679              ( u3_col_out_679     ),
    .col_in_680              ( u3_col_out_680     ),
    .col_in_681              ( u3_col_out_681     ),
    .col_in_682              ( u3_col_out_682     ),
    .col_in_683              ( u3_col_out_683     ),
    .col_in_684              ( u3_col_out_684     ),
    .col_in_685              ( u3_col_out_685     ),
    .col_in_686              ( u3_col_out_686     ),
    .col_in_687              ( u3_col_out_687     ),
    .col_in_688              ( u3_col_out_688     ),
    .col_in_689              ( u3_col_out_689     ),
    .col_in_690              ( u3_col_out_690     ),
    .col_in_691              ( u3_col_out_691     ),
    .col_in_692              ( u3_col_out_692     ),
    .col_in_693              ( u3_col_out_693     ),
    .col_in_694              ( u3_col_out_694     ),
    .col_in_695              ( u3_col_out_695     ),
    .col_in_696              ( u3_col_out_696     ),
    .col_in_697              ( u3_col_out_697     ),
    .col_in_698              ( u3_col_out_698     ),
    .col_in_699              ( u3_col_out_699     ),
    .col_in_700              ( u3_col_out_700     ),
    .col_in_701              ( u3_col_out_701     ),
    .col_in_702              ( u3_col_out_702     ),
    .col_in_703              ( u3_col_out_703     ),
    .col_in_704              ( u3_col_out_704     ),
    .col_in_705              ( u3_col_out_705     ),
    .col_in_706              ( u3_col_out_706     ),
    .col_in_707              ( u3_col_out_707     ),
    .col_in_708              ( u3_col_out_708     ),
    .col_in_709              ( u3_col_out_709     ),
    .col_in_710              ( u3_col_out_710     ),
    .col_in_711              ( u3_col_out_711     ),
    .col_in_712              ( u3_col_out_712     ),
    .col_in_713              ( u3_col_out_713     ),
    .col_in_714              ( u3_col_out_714     ),
    .col_in_715              ( u3_col_out_715     ),
    .col_in_716              ( u3_col_out_716     ),
    .col_in_717              ( u3_col_out_717     ),
    .col_in_718              ( u3_col_out_718     ),
    .col_in_719              ( u3_col_out_719     ),
    .col_in_720              ( u3_col_out_720     ),
    .col_in_721              ( u3_col_out_721     ),
    .col_in_722              ( u3_col_out_722     ),
    .col_in_723              ( u3_col_out_723     ),
    .col_in_724              ( u3_col_out_724     ),
    .col_in_725              ( u3_col_out_725     ),
    .col_in_726              ( u3_col_out_726     ),
    .col_in_727              ( u3_col_out_727     ),
    .col_in_728              ( u3_col_out_728     ),
    .col_in_729              ( u3_col_out_729     ),
    .col_in_730              ( u3_col_out_730     ),
    .col_in_731              ( u3_col_out_731     ),
    .col_in_732              ( u3_col_out_732     ),
    .col_in_733              ( u3_col_out_733     ),
    .col_in_734              ( u3_col_out_734     ),
    .col_in_735              ( u3_col_out_735     ),
    .col_in_736              ( u3_col_out_736     ),
    .col_in_737              ( u3_col_out_737     ),
    .col_in_738              ( u3_col_out_738     ),
    .col_in_739              ( u3_col_out_739     ),
    .col_in_740              ( u3_col_out_740     ),
    .col_in_741              ( u3_col_out_741     ),
    .col_in_742              ( u3_col_out_742     ),
    .col_in_743              ( u3_col_out_743     ),
    .col_in_744              ( u3_col_out_744     ),
    .col_in_745              ( u3_col_out_745     ),
    .col_in_746              ( u3_col_out_746     ),
    .col_in_747              ( u3_col_out_747     ),
    .col_in_748              ( u3_col_out_748     ),
    .col_in_749              ( u3_col_out_749     ),
    .col_in_750              ( u3_col_out_750     ),
    .col_in_751              ( u3_col_out_751     ),
    .col_in_752              ( u3_col_out_752     ),
    .col_in_753              ( u3_col_out_753     ),
    .col_in_754              ( u3_col_out_754     ),
    .col_in_755              ( u3_col_out_755     ),
    .col_in_756              ( u3_col_out_756     ),
    .col_in_757              ( u3_col_out_757     ),
    .col_in_758              ( u3_col_out_758     ),
    .col_in_759              ( u3_col_out_759     ),
    .col_in_760              ( u3_col_out_760     ),
    .col_in_761              ( u3_col_out_761     ),
    .col_in_762              ( u3_col_out_762     ),
    .col_in_763              ( u3_col_out_763     ),
    .col_in_764              ( u3_col_out_764     ),
    .col_in_765              ( u3_col_out_765     ),
    .col_in_766              ( u3_col_out_766     ),
    .col_in_767              ( u3_col_out_767     ),
    .col_in_768              ( u3_col_out_768     ),
    .col_in_769              ( u3_col_out_769     ),
    .col_in_770              ( u3_col_out_770     ),
    .col_in_771              ( u3_col_out_771     ),
    .col_in_772              ( u3_col_out_772     ),
    .col_in_773              ( u3_col_out_773     ),
    .col_in_774              ( u3_col_out_774     ),
    .col_in_775              ( u3_col_out_775     ),
    .col_in_776              ( u3_col_out_776     ),
    .col_in_777              ( u3_col_out_777     ),
    .col_in_778              ( u3_col_out_778     ),
    .col_in_779              ( u3_col_out_779     ),
    .col_in_780              ( u3_col_out_780     ),
    .col_in_781              ( u3_col_out_781     ),
    .col_in_782              ( u3_col_out_782     ),
    .col_in_783              ( u3_col_out_783     ),
    .col_in_784              ( u3_col_out_784     ),
    .col_in_785              ( u3_col_out_785     ),
    .col_in_786              ( u3_col_out_786     ),
    .col_in_787              ( u3_col_out_787     ),
    .col_in_788              ( u3_col_out_788     ),
    .col_in_789              ( u3_col_out_789     ),
    .col_in_790              ( u3_col_out_790     ),
    .col_in_791              ( u3_col_out_791     ),
    .col_in_792              ( u3_col_out_792     ),
    .col_in_793              ( u3_col_out_793     ),
    .col_in_794              ( u3_col_out_794     ),
    .col_in_795              ( u3_col_out_795     ),
    .col_in_796              ( u3_col_out_796     ),
    .col_in_797              ( u3_col_out_797     ),
    .col_in_798              ( u3_col_out_798     ),
    .col_in_799              ( u3_col_out_799     ),
    .col_in_800              ( u3_col_out_800     ),
    .col_in_801              ( u3_col_out_801     ),
    .col_in_802              ( u3_col_out_802     ),
    .col_in_803              ( u3_col_out_803     ),
    .col_in_804              ( u3_col_out_804     ),
    .col_in_805              ( u3_col_out_805     ),
    .col_in_806              ( u3_col_out_806     ),
    .col_in_807              ( u3_col_out_807     ),
    .col_in_808              ( u3_col_out_808     ),
    .col_in_809              ( u3_col_out_809     ),
    .col_in_810              ( u3_col_out_810     ),
    .col_in_811              ( u3_col_out_811     ),
    .col_in_812              ( u3_col_out_812     ),
    .col_in_813              ( u3_col_out_813     ),
    .col_in_814              ( u3_col_out_814     ),
    .col_in_815              ( u3_col_out_815     ),
    .col_in_816              ( u3_col_out_816     ),
    .col_in_817              ( u3_col_out_817     ),
    .col_in_818              ( u3_col_out_818     ),
    .col_in_819              ( u3_col_out_819     ),
    .col_in_820              ( u3_col_out_820     ),
    .col_in_821              ( u3_col_out_821     ),
    .col_in_822              ( u3_col_out_822     ),
    .col_in_823              ( u3_col_out_823     ),
    .col_in_824              ( u3_col_out_824     ),
    .col_in_825              ( u3_col_out_825     ),
    .col_in_826              ( u3_col_out_826     ),
    .col_in_827              ( u3_col_out_827     ),
    .col_in_828              ( u3_col_out_828     ),
    .col_in_829              ( u3_col_out_829     ),
    .col_in_830              ( u3_col_out_830     ),
    .col_in_831              ( u3_col_out_831     ),
    .col_in_832              ( u3_col_out_832     ),
    .col_in_833              ( u3_col_out_833     ),
    .col_in_834              ( u3_col_out_834     ),
    .col_in_835              ( u3_col_out_835     ),
    .col_in_836              ( u3_col_out_836     ),
    .col_in_837              ( u3_col_out_837     ),
    .col_in_838              ( u3_col_out_838     ),
    .col_in_839              ( u3_col_out_839     ),
    .col_in_840              ( u3_col_out_840     ),
    .col_in_841              ( u3_col_out_841     ),
    .col_in_842              ( u3_col_out_842     ),
    .col_in_843              ( u3_col_out_843     ),
    .col_in_844              ( u3_col_out_844     ),
    .col_in_845              ( u3_col_out_845     ),
    .col_in_846              ( u3_col_out_846     ),
    .col_in_847              ( u3_col_out_847     ),
    .col_in_848              ( u3_col_out_848     ),
    .col_in_849              ( u3_col_out_849     ),
    .col_in_850              ( u3_col_out_850     ),
    .col_in_851              ( u3_col_out_851     ),
    .col_in_852              ( u3_col_out_852     ),
    .col_in_853              ( u3_col_out_853     ),
    .col_in_854              ( u3_col_out_854     ),
    .col_in_855              ( u3_col_out_855     ),
    .col_in_856              ( u3_col_out_856     ),
    .col_in_857              ( u3_col_out_857     ),
    .col_in_858              ( u3_col_out_858     ),
    .col_in_859              ( u3_col_out_859     ),
    .col_in_860              ( u3_col_out_860     ),
    .col_in_861              ( u3_col_out_861     ),
    .col_in_862              ( u3_col_out_862     ),
    .col_in_863              ( u3_col_out_863     ),
    .col_in_864              ( u3_col_out_864     ),
    .col_in_865              ( u3_col_out_865     ),
    .col_in_866              ( u3_col_out_866     ),
    .col_in_867              ( u3_col_out_867     ),
    .col_in_868              ( u3_col_out_868     ),
    .col_in_869              ( u3_col_out_869     ),
    .col_in_870              ( u3_col_out_870     ),
    .col_in_871              ( u3_col_out_871     ),
    .col_in_872              ( u3_col_out_872     ),
    .col_in_873              ( u3_col_out_873     ),
    .col_in_874              ( u3_col_out_874     ),
    .col_in_875              ( u3_col_out_875     ),
    .col_in_876              ( u3_col_out_876     ),
    .col_in_877              ( u3_col_out_877     ),
    .col_in_878              ( u3_col_out_878     ),
    .col_in_879              ( u3_col_out_879     ),
    .col_in_880              ( u3_col_out_880     ),
    .col_in_881              ( u3_col_out_881     ),
    .col_in_882              ( u3_col_out_882     ),
    .col_in_883              ( u3_col_out_883     ),
    .col_in_884              ( u3_col_out_884     ),
    .col_in_885              ( u3_col_out_885     ),
    .col_in_886              ( u3_col_out_886     ),
    .col_in_887              ( u3_col_out_887     ),
    .col_in_888              ( u3_col_out_888     ),
    .col_in_889              ( u3_col_out_889     ),
    .col_in_890              ( u3_col_out_890     ),
    .col_in_891              ( u3_col_out_891     ),
    .col_in_892              ( u3_col_out_892     ),
    .col_in_893              ( u3_col_out_893     ),
    .col_in_894              ( u3_col_out_894     ),
    .col_in_895              ( u3_col_out_895     ),
    .col_in_896              ( u3_col_out_896     ),
    .col_in_897              ( u3_col_out_897     ),
    .col_in_898              ( u3_col_out_898     ),
    .col_in_899              ( u3_col_out_899     ),
    .col_in_900              ( u3_col_out_900     ),
    .col_in_901              ( u3_col_out_901     ),
    .col_in_902              ( u3_col_out_902     ),
    .col_in_903              ( u3_col_out_903     ),
    .col_in_904              ( u3_col_out_904     ),
    .col_in_905              ( u3_col_out_905     ),
    .col_in_906              ( u3_col_out_906     ),
    .col_in_907              ( u3_col_out_907     ),
    .col_in_908              ( u3_col_out_908     ),
    .col_in_909              ( u3_col_out_909     ),
    .col_in_910              ( u3_col_out_910     ),
    .col_in_911              ( u3_col_out_911     ),
    .col_in_912              ( u3_col_out_912     ),
    .col_in_913              ( u3_col_out_913     ),
    .col_in_914              ( u3_col_out_914     ),
    .col_in_915              ( u3_col_out_915     ),
    .col_in_916              ( u3_col_out_916     ),
    .col_in_917              ( u3_col_out_917     ),
    .col_in_918              ( u3_col_out_918     ),
    .col_in_919              ( u3_col_out_919     ),
    .col_in_920              ( u3_col_out_920     ),
    .col_in_921              ( u3_col_out_921     ),
    .col_in_922              ( u3_col_out_922     ),
    .col_in_923              ( u3_col_out_923     ),
    .col_in_924              ( u3_col_out_924     ),
    .col_in_925              ( u3_col_out_925     ),
    .col_in_926              ( u3_col_out_926     ),
    .col_in_927              ( u3_col_out_927     ),
    .col_in_928              ( u3_col_out_928     ),
    .col_in_929              ( u3_col_out_929     ),
    .col_in_930              ( u3_col_out_930     ),
    .col_in_931              ( u3_col_out_931     ),
    .col_in_932              ( u3_col_out_932     ),
    .col_in_933              ( u3_col_out_933     ),
    .col_in_934              ( u3_col_out_934     ),
    .col_in_935              ( u3_col_out_935     ),
    .col_in_936              ( u3_col_out_936     ),
    .col_in_937              ( u3_col_out_937     ),
    .col_in_938              ( u3_col_out_938     ),
    .col_in_939              ( u3_col_out_939     ),
    .col_in_940              ( u3_col_out_940     ),
    .col_in_941              ( u3_col_out_941     ),
    .col_in_942              ( u3_col_out_942     ),
    .col_in_943              ( u3_col_out_943     ),
    .col_in_944              ( u3_col_out_944     ),
    .col_in_945              ( u3_col_out_945     ),
    .col_in_946              ( u3_col_out_946     ),
    .col_in_947              ( u3_col_out_947     ),
    .col_in_948              ( u3_col_out_948     ),
    .col_in_949              ( u3_col_out_949     ),
    .col_in_950              ( u3_col_out_950     ),
    .col_in_951              ( u3_col_out_951     ),
    .col_in_952              ( u3_col_out_952     ),
    .col_in_953              ( u3_col_out_953     ),
    .col_in_954              ( u3_col_out_954     ),
    .col_in_955              ( u3_col_out_955     ),
    .col_in_956              ( u3_col_out_956     ),
    .col_in_957              ( u3_col_out_957     ),
    .col_in_958              ( u3_col_out_958     ),
    .col_in_959              ( u3_col_out_959     ),
    .col_in_960              ( u3_col_out_960     ),
    .col_in_961              ( u3_col_out_961     ),
    .col_in_962              ( u3_col_out_962     ),
    .col_in_963              ( u3_col_out_963     ),
    .col_in_964              ( u3_col_out_964     ),
    .col_in_965              ( u3_col_out_965     ),
    .col_in_966              ( u3_col_out_966     ),
    .col_in_967              ( u3_col_out_967     ),
    .col_in_968              ( u3_col_out_968     ),
    .col_in_969              ( u3_col_out_969     ),
    .col_in_970              ( u3_col_out_970     ),
    .col_in_971              ( u3_col_out_971     ),
    .col_in_972              ( u3_col_out_972     ),
    .col_in_973              ( u3_col_out_973     ),
    .col_in_974              ( u3_col_out_974     ),
    .col_in_975              ( u3_col_out_975     ),
    .col_in_976              ( u3_col_out_976     ),
    .col_in_977              ( u3_col_out_977     ),
    .col_in_978              ( u3_col_out_978     ),
    .col_in_979              ( u3_col_out_979     ),
    .col_in_980              ( u3_col_out_980     ),
    .col_in_981              ( u3_col_out_981     ),
    .col_in_982              ( u3_col_out_982     ),
    .col_in_983              ( u3_col_out_983     ),
    .col_in_984              ( u3_col_out_984     ),
    .col_in_985              ( u3_col_out_985     ),
    .col_in_986              ( u3_col_out_986     ),
    .col_in_987              ( u3_col_out_987     ),
    .col_in_988              ( u3_col_out_988     ),
    .col_in_989              ( u3_col_out_989     ),
    .col_in_990              ( u3_col_out_990     ),
    .col_in_991              ( u3_col_out_991     ),
    .col_in_992              ( u3_col_out_992     ),
    .col_in_993              ( u3_col_out_993     ),
    .col_in_994              ( u3_col_out_994     ),
    .col_in_995              ( u3_col_out_995     ),
    .col_in_996              ( u3_col_out_996     ),
    .col_in_997              ( u3_col_out_997     ),
    .col_in_998              ( u3_col_out_998     ),
    .col_in_999              ( u3_col_out_999     ),
    .col_in_1000             ( u3_col_out_1000    ),
    .col_in_1001             ( u3_col_out_1001    ),
    .col_in_1002             ( u3_col_out_1002    ),
    .col_in_1003             ( u3_col_out_1003    ),
    .col_in_1004             ( u3_col_out_1004    ),
    .col_in_1005             ( u3_col_out_1005    ),
    .col_in_1006             ( u3_col_out_1006    ),
    .col_in_1007             ( u3_col_out_1007    ),
    .col_in_1008             ( u3_col_out_1008    ),
    .col_in_1009             ( u3_col_out_1009    ),
    .col_in_1010             ( u3_col_out_1010    ),
    .col_in_1011             ( u3_col_out_1011    ),
    .col_in_1012             ( u3_col_out_1012    ),
    .col_in_1013             ( u3_col_out_1013    ),
    .col_in_1014             ( u3_col_out_1014    ),
    .col_in_1015             ( u3_col_out_1015    ),
    .col_in_1016             ( u3_col_out_1016    ),
    .col_in_1017             ( u3_col_out_1017    ),
    .col_in_1018             ( u3_col_out_1018    ),
    .col_in_1019             ( u3_col_out_1019    ),
    .col_in_1020             ( u3_col_out_1020    ),
    .col_in_1021             ( u3_col_out_1021    ),
    .col_in_1022             ( u3_col_out_1022    ),
    .col_in_1023             ( u3_col_out_1023    ),
    .col_in_1024             ( u3_col_out_1024    ),
    .col_in_1025             ( u3_col_out_1025    ),
    .col_in_1026             ( u3_col_out_1026    ),
    .col_in_1027             ( u3_col_out_1027    ),
    .col_in_1028             ( u3_col_out_1028    ),
    .col_in_1029             ( u3_col_out_1029    ),
    .col_in_1030             ( u3_col_out_1030    ),
    .col_in_1031             ( u3_col_out_1031    ),
    .col_in_1032             ( u3_col_out_1032    ),


    .col_out_0               ( u4_col_out_0      ),
    .col_out_1               ( u4_col_out_1      ),
    .col_out_2               ( u4_col_out_2      ),
    .col_out_3               ( u4_col_out_3      ),
    .col_out_4               ( u4_col_out_4      ),
    .col_out_5               ( u4_col_out_5      ),
    .col_out_6               ( u4_col_out_6      ),
    .col_out_7               ( u4_col_out_7      ),
    .col_out_8               ( u4_col_out_8      ),
    .col_out_9               ( u4_col_out_9      ),
    .col_out_10              ( u4_col_out_10     ),
    .col_out_11              ( u4_col_out_11     ),
    .col_out_12              ( u4_col_out_12     ),
    .col_out_13              ( u4_col_out_13     ),
    .col_out_14              ( u4_col_out_14     ),
    .col_out_15              ( u4_col_out_15     ),
    .col_out_16              ( u4_col_out_16     ),
    .col_out_17              ( u4_col_out_17     ),
    .col_out_18              ( u4_col_out_18     ),
    .col_out_19              ( u4_col_out_19     ),
    .col_out_20              ( u4_col_out_20     ),
    .col_out_21              ( u4_col_out_21     ),
    .col_out_22              ( u4_col_out_22     ),
    .col_out_23              ( u4_col_out_23     ),
    .col_out_24              ( u4_col_out_24     ),
    .col_out_25              ( u4_col_out_25     ),
    .col_out_26              ( u4_col_out_26     ),
    .col_out_27              ( u4_col_out_27     ),
    .col_out_28              ( u4_col_out_28     ),
    .col_out_29              ( u4_col_out_29     ),
    .col_out_30              ( u4_col_out_30     ),
    .col_out_31              ( u4_col_out_31     ),
    .col_out_32              ( u4_col_out_32     ),
    .col_out_33              ( u4_col_out_33     ),
    .col_out_34              ( u4_col_out_34     ),
    .col_out_35              ( u4_col_out_35     ),
    .col_out_36              ( u4_col_out_36     ),
    .col_out_37              ( u4_col_out_37     ),
    .col_out_38              ( u4_col_out_38     ),
    .col_out_39              ( u4_col_out_39     ),
    .col_out_40              ( u4_col_out_40     ),
    .col_out_41              ( u4_col_out_41     ),
    .col_out_42              ( u4_col_out_42     ),
    .col_out_43              ( u4_col_out_43     ),
    .col_out_44              ( u4_col_out_44     ),
    .col_out_45              ( u4_col_out_45     ),
    .col_out_46              ( u4_col_out_46     ),
    .col_out_47              ( u4_col_out_47     ),
    .col_out_48              ( u4_col_out_48     ),
    .col_out_49              ( u4_col_out_49     ),
    .col_out_50              ( u4_col_out_50     ),
    .col_out_51              ( u4_col_out_51     ),
    .col_out_52              ( u4_col_out_52     ),
    .col_out_53              ( u4_col_out_53     ),
    .col_out_54              ( u4_col_out_54     ),
    .col_out_55              ( u4_col_out_55     ),
    .col_out_56              ( u4_col_out_56     ),
    .col_out_57              ( u4_col_out_57     ),
    .col_out_58              ( u4_col_out_58     ),
    .col_out_59              ( u4_col_out_59     ),
    .col_out_60              ( u4_col_out_60     ),
    .col_out_61              ( u4_col_out_61     ),
    .col_out_62              ( u4_col_out_62     ),
    .col_out_63              ( u4_col_out_63     ),
    .col_out_64              ( u4_col_out_64     ),
    .col_out_65              ( u4_col_out_65     ),
    .col_out_66              ( u4_col_out_66     ),
    .col_out_67              ( u4_col_out_67     ),
    .col_out_68              ( u4_col_out_68     ),
    .col_out_69              ( u4_col_out_69     ),
    .col_out_70              ( u4_col_out_70     ),
    .col_out_71              ( u4_col_out_71     ),
    .col_out_72              ( u4_col_out_72     ),
    .col_out_73              ( u4_col_out_73     ),
    .col_out_74              ( u4_col_out_74     ),
    .col_out_75              ( u4_col_out_75     ),
    .col_out_76              ( u4_col_out_76     ),
    .col_out_77              ( u4_col_out_77     ),
    .col_out_78              ( u4_col_out_78     ),
    .col_out_79              ( u4_col_out_79     ),
    .col_out_80              ( u4_col_out_80     ),
    .col_out_81              ( u4_col_out_81     ),
    .col_out_82              ( u4_col_out_82     ),
    .col_out_83              ( u4_col_out_83     ),
    .col_out_84              ( u4_col_out_84     ),
    .col_out_85              ( u4_col_out_85     ),
    .col_out_86              ( u4_col_out_86     ),
    .col_out_87              ( u4_col_out_87     ),
    .col_out_88              ( u4_col_out_88     ),
    .col_out_89              ( u4_col_out_89     ),
    .col_out_90              ( u4_col_out_90     ),
    .col_out_91              ( u4_col_out_91     ),
    .col_out_92              ( u4_col_out_92     ),
    .col_out_93              ( u4_col_out_93     ),
    .col_out_94              ( u4_col_out_94     ),
    .col_out_95              ( u4_col_out_95     ),
    .col_out_96              ( u4_col_out_96     ),
    .col_out_97              ( u4_col_out_97     ),
    .col_out_98              ( u4_col_out_98     ),
    .col_out_99              ( u4_col_out_99     ),
    .col_out_100             ( u4_col_out_100    ),
    .col_out_101             ( u4_col_out_101    ),
    .col_out_102             ( u4_col_out_102    ),
    .col_out_103             ( u4_col_out_103    ),
    .col_out_104             ( u4_col_out_104    ),
    .col_out_105             ( u4_col_out_105    ),
    .col_out_106             ( u4_col_out_106    ),
    .col_out_107             ( u4_col_out_107    ),
    .col_out_108             ( u4_col_out_108    ),
    .col_out_109             ( u4_col_out_109    ),
    .col_out_110             ( u4_col_out_110    ),
    .col_out_111             ( u4_col_out_111    ),
    .col_out_112             ( u4_col_out_112    ),
    .col_out_113             ( u4_col_out_113    ),
    .col_out_114             ( u4_col_out_114    ),
    .col_out_115             ( u4_col_out_115    ),
    .col_out_116             ( u4_col_out_116    ),
    .col_out_117             ( u4_col_out_117    ),
    .col_out_118             ( u4_col_out_118    ),
    .col_out_119             ( u4_col_out_119    ),
    .col_out_120             ( u4_col_out_120    ),
    .col_out_121             ( u4_col_out_121    ),
    .col_out_122             ( u4_col_out_122    ),
    .col_out_123             ( u4_col_out_123    ),
    .col_out_124             ( u4_col_out_124    ),
    .col_out_125             ( u4_col_out_125    ),
    .col_out_126             ( u4_col_out_126    ),
    .col_out_127             ( u4_col_out_127    ),
    .col_out_128             ( u4_col_out_128    ),
    .col_out_129             ( u4_col_out_129    ),
    .col_out_130             ( u4_col_out_130    ),
    .col_out_131             ( u4_col_out_131    ),
    .col_out_132             ( u4_col_out_132    ),
    .col_out_133             ( u4_col_out_133    ),
    .col_out_134             ( u4_col_out_134    ),
    .col_out_135             ( u4_col_out_135    ),
    .col_out_136             ( u4_col_out_136    ),
    .col_out_137             ( u4_col_out_137    ),
    .col_out_138             ( u4_col_out_138    ),
    .col_out_139             ( u4_col_out_139    ),
    .col_out_140             ( u4_col_out_140    ),
    .col_out_141             ( u4_col_out_141    ),
    .col_out_142             ( u4_col_out_142    ),
    .col_out_143             ( u4_col_out_143    ),
    .col_out_144             ( u4_col_out_144    ),
    .col_out_145             ( u4_col_out_145    ),
    .col_out_146             ( u4_col_out_146    ),
    .col_out_147             ( u4_col_out_147    ),
    .col_out_148             ( u4_col_out_148    ),
    .col_out_149             ( u4_col_out_149    ),
    .col_out_150             ( u4_col_out_150    ),
    .col_out_151             ( u4_col_out_151    ),
    .col_out_152             ( u4_col_out_152    ),
    .col_out_153             ( u4_col_out_153    ),
    .col_out_154             ( u4_col_out_154    ),
    .col_out_155             ( u4_col_out_155    ),
    .col_out_156             ( u4_col_out_156    ),
    .col_out_157             ( u4_col_out_157    ),
    .col_out_158             ( u4_col_out_158    ),
    .col_out_159             ( u4_col_out_159    ),
    .col_out_160             ( u4_col_out_160    ),
    .col_out_161             ( u4_col_out_161    ),
    .col_out_162             ( u4_col_out_162    ),
    .col_out_163             ( u4_col_out_163    ),
    .col_out_164             ( u4_col_out_164    ),
    .col_out_165             ( u4_col_out_165    ),
    .col_out_166             ( u4_col_out_166    ),
    .col_out_167             ( u4_col_out_167    ),
    .col_out_168             ( u4_col_out_168    ),
    .col_out_169             ( u4_col_out_169    ),
    .col_out_170             ( u4_col_out_170    ),
    .col_out_171             ( u4_col_out_171    ),
    .col_out_172             ( u4_col_out_172    ),
    .col_out_173             ( u4_col_out_173    ),
    .col_out_174             ( u4_col_out_174    ),
    .col_out_175             ( u4_col_out_175    ),
    .col_out_176             ( u4_col_out_176    ),
    .col_out_177             ( u4_col_out_177    ),
    .col_out_178             ( u4_col_out_178    ),
    .col_out_179             ( u4_col_out_179    ),
    .col_out_180             ( u4_col_out_180    ),
    .col_out_181             ( u4_col_out_181    ),
    .col_out_182             ( u4_col_out_182    ),
    .col_out_183             ( u4_col_out_183    ),
    .col_out_184             ( u4_col_out_184    ),
    .col_out_185             ( u4_col_out_185    ),
    .col_out_186             ( u4_col_out_186    ),
    .col_out_187             ( u4_col_out_187    ),
    .col_out_188             ( u4_col_out_188    ),
    .col_out_189             ( u4_col_out_189    ),
    .col_out_190             ( u4_col_out_190    ),
    .col_out_191             ( u4_col_out_191    ),
    .col_out_192             ( u4_col_out_192    ),
    .col_out_193             ( u4_col_out_193    ),
    .col_out_194             ( u4_col_out_194    ),
    .col_out_195             ( u4_col_out_195    ),
    .col_out_196             ( u4_col_out_196    ),
    .col_out_197             ( u4_col_out_197    ),
    .col_out_198             ( u4_col_out_198    ),
    .col_out_199             ( u4_col_out_199    ),
    .col_out_200             ( u4_col_out_200    ),
    .col_out_201             ( u4_col_out_201    ),
    .col_out_202             ( u4_col_out_202    ),
    .col_out_203             ( u4_col_out_203    ),
    .col_out_204             ( u4_col_out_204    ),
    .col_out_205             ( u4_col_out_205    ),
    .col_out_206             ( u4_col_out_206    ),
    .col_out_207             ( u4_col_out_207    ),
    .col_out_208             ( u4_col_out_208    ),
    .col_out_209             ( u4_col_out_209    ),
    .col_out_210             ( u4_col_out_210    ),
    .col_out_211             ( u4_col_out_211    ),
    .col_out_212             ( u4_col_out_212    ),
    .col_out_213             ( u4_col_out_213    ),
    .col_out_214             ( u4_col_out_214    ),
    .col_out_215             ( u4_col_out_215    ),
    .col_out_216             ( u4_col_out_216    ),
    .col_out_217             ( u4_col_out_217    ),
    .col_out_218             ( u4_col_out_218    ),
    .col_out_219             ( u4_col_out_219    ),
    .col_out_220             ( u4_col_out_220    ),
    .col_out_221             ( u4_col_out_221    ),
    .col_out_222             ( u4_col_out_222    ),
    .col_out_223             ( u4_col_out_223    ),
    .col_out_224             ( u4_col_out_224    ),
    .col_out_225             ( u4_col_out_225    ),
    .col_out_226             ( u4_col_out_226    ),
    .col_out_227             ( u4_col_out_227    ),
    .col_out_228             ( u4_col_out_228    ),
    .col_out_229             ( u4_col_out_229    ),
    .col_out_230             ( u4_col_out_230    ),
    .col_out_231             ( u4_col_out_231    ),
    .col_out_232             ( u4_col_out_232    ),
    .col_out_233             ( u4_col_out_233    ),
    .col_out_234             ( u4_col_out_234    ),
    .col_out_235             ( u4_col_out_235    ),
    .col_out_236             ( u4_col_out_236    ),
    .col_out_237             ( u4_col_out_237    ),
    .col_out_238             ( u4_col_out_238    ),
    .col_out_239             ( u4_col_out_239    ),
    .col_out_240             ( u4_col_out_240    ),
    .col_out_241             ( u4_col_out_241    ),
    .col_out_242             ( u4_col_out_242    ),
    .col_out_243             ( u4_col_out_243    ),
    .col_out_244             ( u4_col_out_244    ),
    .col_out_245             ( u4_col_out_245    ),
    .col_out_246             ( u4_col_out_246    ),
    .col_out_247             ( u4_col_out_247    ),
    .col_out_248             ( u4_col_out_248    ),
    .col_out_249             ( u4_col_out_249    ),
    .col_out_250             ( u4_col_out_250    ),
    .col_out_251             ( u4_col_out_251    ),
    .col_out_252             ( u4_col_out_252    ),
    .col_out_253             ( u4_col_out_253    ),
    .col_out_254             ( u4_col_out_254    ),
    .col_out_255             ( u4_col_out_255    ),
    .col_out_256             ( u4_col_out_256    ),
    .col_out_257             ( u4_col_out_257    ),
    .col_out_258             ( u4_col_out_258    ),
    .col_out_259             ( u4_col_out_259    ),
    .col_out_260             ( u4_col_out_260    ),
    .col_out_261             ( u4_col_out_261    ),
    .col_out_262             ( u4_col_out_262    ),
    .col_out_263             ( u4_col_out_263    ),
    .col_out_264             ( u4_col_out_264    ),
    .col_out_265             ( u4_col_out_265    ),
    .col_out_266             ( u4_col_out_266    ),
    .col_out_267             ( u4_col_out_267    ),
    .col_out_268             ( u4_col_out_268    ),
    .col_out_269             ( u4_col_out_269    ),
    .col_out_270             ( u4_col_out_270    ),
    .col_out_271             ( u4_col_out_271    ),
    .col_out_272             ( u4_col_out_272    ),
    .col_out_273             ( u4_col_out_273    ),
    .col_out_274             ( u4_col_out_274    ),
    .col_out_275             ( u4_col_out_275    ),
    .col_out_276             ( u4_col_out_276    ),
    .col_out_277             ( u4_col_out_277    ),
    .col_out_278             ( u4_col_out_278    ),
    .col_out_279             ( u4_col_out_279    ),
    .col_out_280             ( u4_col_out_280    ),
    .col_out_281             ( u4_col_out_281    ),
    .col_out_282             ( u4_col_out_282    ),
    .col_out_283             ( u4_col_out_283    ),
    .col_out_284             ( u4_col_out_284    ),
    .col_out_285             ( u4_col_out_285    ),
    .col_out_286             ( u4_col_out_286    ),
    .col_out_287             ( u4_col_out_287    ),
    .col_out_288             ( u4_col_out_288    ),
    .col_out_289             ( u4_col_out_289    ),
    .col_out_290             ( u4_col_out_290    ),
    .col_out_291             ( u4_col_out_291    ),
    .col_out_292             ( u4_col_out_292    ),
    .col_out_293             ( u4_col_out_293    ),
    .col_out_294             ( u4_col_out_294    ),
    .col_out_295             ( u4_col_out_295    ),
    .col_out_296             ( u4_col_out_296    ),
    .col_out_297             ( u4_col_out_297    ),
    .col_out_298             ( u4_col_out_298    ),
    .col_out_299             ( u4_col_out_299    ),
    .col_out_300             ( u4_col_out_300    ),
    .col_out_301             ( u4_col_out_301    ),
    .col_out_302             ( u4_col_out_302    ),
    .col_out_303             ( u4_col_out_303    ),
    .col_out_304             ( u4_col_out_304    ),
    .col_out_305             ( u4_col_out_305    ),
    .col_out_306             ( u4_col_out_306    ),
    .col_out_307             ( u4_col_out_307    ),
    .col_out_308             ( u4_col_out_308    ),
    .col_out_309             ( u4_col_out_309    ),
    .col_out_310             ( u4_col_out_310    ),
    .col_out_311             ( u4_col_out_311    ),
    .col_out_312             ( u4_col_out_312    ),
    .col_out_313             ( u4_col_out_313    ),
    .col_out_314             ( u4_col_out_314    ),
    .col_out_315             ( u4_col_out_315    ),
    .col_out_316             ( u4_col_out_316    ),
    .col_out_317             ( u4_col_out_317    ),
    .col_out_318             ( u4_col_out_318    ),
    .col_out_319             ( u4_col_out_319    ),
    .col_out_320             ( u4_col_out_320    ),
    .col_out_321             ( u4_col_out_321    ),
    .col_out_322             ( u4_col_out_322    ),
    .col_out_323             ( u4_col_out_323    ),
    .col_out_324             ( u4_col_out_324    ),
    .col_out_325             ( u4_col_out_325    ),
    .col_out_326             ( u4_col_out_326    ),
    .col_out_327             ( u4_col_out_327    ),
    .col_out_328             ( u4_col_out_328    ),
    .col_out_329             ( u4_col_out_329    ),
    .col_out_330             ( u4_col_out_330    ),
    .col_out_331             ( u4_col_out_331    ),
    .col_out_332             ( u4_col_out_332    ),
    .col_out_333             ( u4_col_out_333    ),
    .col_out_334             ( u4_col_out_334    ),
    .col_out_335             ( u4_col_out_335    ),
    .col_out_336             ( u4_col_out_336    ),
    .col_out_337             ( u4_col_out_337    ),
    .col_out_338             ( u4_col_out_338    ),
    .col_out_339             ( u4_col_out_339    ),
    .col_out_340             ( u4_col_out_340    ),
    .col_out_341             ( u4_col_out_341    ),
    .col_out_342             ( u4_col_out_342    ),
    .col_out_343             ( u4_col_out_343    ),
    .col_out_344             ( u4_col_out_344    ),
    .col_out_345             ( u4_col_out_345    ),
    .col_out_346             ( u4_col_out_346    ),
    .col_out_347             ( u4_col_out_347    ),
    .col_out_348             ( u4_col_out_348    ),
    .col_out_349             ( u4_col_out_349    ),
    .col_out_350             ( u4_col_out_350    ),
    .col_out_351             ( u4_col_out_351    ),
    .col_out_352             ( u4_col_out_352    ),
    .col_out_353             ( u4_col_out_353    ),
    .col_out_354             ( u4_col_out_354    ),
    .col_out_355             ( u4_col_out_355    ),
    .col_out_356             ( u4_col_out_356    ),
    .col_out_357             ( u4_col_out_357    ),
    .col_out_358             ( u4_col_out_358    ),
    .col_out_359             ( u4_col_out_359    ),
    .col_out_360             ( u4_col_out_360    ),
    .col_out_361             ( u4_col_out_361    ),
    .col_out_362             ( u4_col_out_362    ),
    .col_out_363             ( u4_col_out_363    ),
    .col_out_364             ( u4_col_out_364    ),
    .col_out_365             ( u4_col_out_365    ),
    .col_out_366             ( u4_col_out_366    ),
    .col_out_367             ( u4_col_out_367    ),
    .col_out_368             ( u4_col_out_368    ),
    .col_out_369             ( u4_col_out_369    ),
    .col_out_370             ( u4_col_out_370    ),
    .col_out_371             ( u4_col_out_371    ),
    .col_out_372             ( u4_col_out_372    ),
    .col_out_373             ( u4_col_out_373    ),
    .col_out_374             ( u4_col_out_374    ),
    .col_out_375             ( u4_col_out_375    ),
    .col_out_376             ( u4_col_out_376    ),
    .col_out_377             ( u4_col_out_377    ),
    .col_out_378             ( u4_col_out_378    ),
    .col_out_379             ( u4_col_out_379    ),
    .col_out_380             ( u4_col_out_380    ),
    .col_out_381             ( u4_col_out_381    ),
    .col_out_382             ( u4_col_out_382    ),
    .col_out_383             ( u4_col_out_383    ),
    .col_out_384             ( u4_col_out_384    ),
    .col_out_385             ( u4_col_out_385    ),
    .col_out_386             ( u4_col_out_386    ),
    .col_out_387             ( u4_col_out_387    ),
    .col_out_388             ( u4_col_out_388    ),
    .col_out_389             ( u4_col_out_389    ),
    .col_out_390             ( u4_col_out_390    ),
    .col_out_391             ( u4_col_out_391    ),
    .col_out_392             ( u4_col_out_392    ),
    .col_out_393             ( u4_col_out_393    ),
    .col_out_394             ( u4_col_out_394    ),
    .col_out_395             ( u4_col_out_395    ),
    .col_out_396             ( u4_col_out_396    ),
    .col_out_397             ( u4_col_out_397    ),
    .col_out_398             ( u4_col_out_398    ),
    .col_out_399             ( u4_col_out_399    ),
    .col_out_400             ( u4_col_out_400    ),
    .col_out_401             ( u4_col_out_401    ),
    .col_out_402             ( u4_col_out_402    ),
    .col_out_403             ( u4_col_out_403    ),
    .col_out_404             ( u4_col_out_404    ),
    .col_out_405             ( u4_col_out_405    ),
    .col_out_406             ( u4_col_out_406    ),
    .col_out_407             ( u4_col_out_407    ),
    .col_out_408             ( u4_col_out_408    ),
    .col_out_409             ( u4_col_out_409    ),
    .col_out_410             ( u4_col_out_410    ),
    .col_out_411             ( u4_col_out_411    ),
    .col_out_412             ( u4_col_out_412    ),
    .col_out_413             ( u4_col_out_413    ),
    .col_out_414             ( u4_col_out_414    ),
    .col_out_415             ( u4_col_out_415    ),
    .col_out_416             ( u4_col_out_416    ),
    .col_out_417             ( u4_col_out_417    ),
    .col_out_418             ( u4_col_out_418    ),
    .col_out_419             ( u4_col_out_419    ),
    .col_out_420             ( u4_col_out_420    ),
    .col_out_421             ( u4_col_out_421    ),
    .col_out_422             ( u4_col_out_422    ),
    .col_out_423             ( u4_col_out_423    ),
    .col_out_424             ( u4_col_out_424    ),
    .col_out_425             ( u4_col_out_425    ),
    .col_out_426             ( u4_col_out_426    ),
    .col_out_427             ( u4_col_out_427    ),
    .col_out_428             ( u4_col_out_428    ),
    .col_out_429             ( u4_col_out_429    ),
    .col_out_430             ( u4_col_out_430    ),
    .col_out_431             ( u4_col_out_431    ),
    .col_out_432             ( u4_col_out_432    ),
    .col_out_433             ( u4_col_out_433    ),
    .col_out_434             ( u4_col_out_434    ),
    .col_out_435             ( u4_col_out_435    ),
    .col_out_436             ( u4_col_out_436    ),
    .col_out_437             ( u4_col_out_437    ),
    .col_out_438             ( u4_col_out_438    ),
    .col_out_439             ( u4_col_out_439    ),
    .col_out_440             ( u4_col_out_440    ),
    .col_out_441             ( u4_col_out_441    ),
    .col_out_442             ( u4_col_out_442    ),
    .col_out_443             ( u4_col_out_443    ),
    .col_out_444             ( u4_col_out_444    ),
    .col_out_445             ( u4_col_out_445    ),
    .col_out_446             ( u4_col_out_446    ),
    .col_out_447             ( u4_col_out_447    ),
    .col_out_448             ( u4_col_out_448    ),
    .col_out_449             ( u4_col_out_449    ),
    .col_out_450             ( u4_col_out_450    ),
    .col_out_451             ( u4_col_out_451    ),
    .col_out_452             ( u4_col_out_452    ),
    .col_out_453             ( u4_col_out_453    ),
    .col_out_454             ( u4_col_out_454    ),
    .col_out_455             ( u4_col_out_455    ),
    .col_out_456             ( u4_col_out_456    ),
    .col_out_457             ( u4_col_out_457    ),
    .col_out_458             ( u4_col_out_458    ),
    .col_out_459             ( u4_col_out_459    ),
    .col_out_460             ( u4_col_out_460    ),
    .col_out_461             ( u4_col_out_461    ),
    .col_out_462             ( u4_col_out_462    ),
    .col_out_463             ( u4_col_out_463    ),
    .col_out_464             ( u4_col_out_464    ),
    .col_out_465             ( u4_col_out_465    ),
    .col_out_466             ( u4_col_out_466    ),
    .col_out_467             ( u4_col_out_467    ),
    .col_out_468             ( u4_col_out_468    ),
    .col_out_469             ( u4_col_out_469    ),
    .col_out_470             ( u4_col_out_470    ),
    .col_out_471             ( u4_col_out_471    ),
    .col_out_472             ( u4_col_out_472    ),
    .col_out_473             ( u4_col_out_473    ),
    .col_out_474             ( u4_col_out_474    ),
    .col_out_475             ( u4_col_out_475    ),
    .col_out_476             ( u4_col_out_476    ),
    .col_out_477             ( u4_col_out_477    ),
    .col_out_478             ( u4_col_out_478    ),
    .col_out_479             ( u4_col_out_479    ),
    .col_out_480             ( u4_col_out_480    ),
    .col_out_481             ( u4_col_out_481    ),
    .col_out_482             ( u4_col_out_482    ),
    .col_out_483             ( u4_col_out_483    ),
    .col_out_484             ( u4_col_out_484    ),
    .col_out_485             ( u4_col_out_485    ),
    .col_out_486             ( u4_col_out_486    ),
    .col_out_487             ( u4_col_out_487    ),
    .col_out_488             ( u4_col_out_488    ),
    .col_out_489             ( u4_col_out_489    ),
    .col_out_490             ( u4_col_out_490    ),
    .col_out_491             ( u4_col_out_491    ),
    .col_out_492             ( u4_col_out_492    ),
    .col_out_493             ( u4_col_out_493    ),
    .col_out_494             ( u4_col_out_494    ),
    .col_out_495             ( u4_col_out_495    ),
    .col_out_496             ( u4_col_out_496    ),
    .col_out_497             ( u4_col_out_497    ),
    .col_out_498             ( u4_col_out_498    ),
    .col_out_499             ( u4_col_out_499    ),
    .col_out_500             ( u4_col_out_500    ),
    .col_out_501             ( u4_col_out_501    ),
    .col_out_502             ( u4_col_out_502    ),
    .col_out_503             ( u4_col_out_503    ),
    .col_out_504             ( u4_col_out_504    ),
    .col_out_505             ( u4_col_out_505    ),
    .col_out_506             ( u4_col_out_506    ),
    .col_out_507             ( u4_col_out_507    ),
    .col_out_508             ( u4_col_out_508    ),
    .col_out_509             ( u4_col_out_509    ),
    .col_out_510             ( u4_col_out_510    ),
    .col_out_511             ( u4_col_out_511    ),
    .col_out_512             ( u4_col_out_512    ),
    .col_out_513             ( u4_col_out_513    ),
    .col_out_514             ( u4_col_out_514    ),
    .col_out_515             ( u4_col_out_515    ),
    .col_out_516             ( u4_col_out_516    ),
    .col_out_517             ( u4_col_out_517    ),
    .col_out_518             ( u4_col_out_518    ),
    .col_out_519             ( u4_col_out_519    ),
    .col_out_520             ( u4_col_out_520    ),
    .col_out_521             ( u4_col_out_521    ),
    .col_out_522             ( u4_col_out_522    ),
    .col_out_523             ( u4_col_out_523    ),
    .col_out_524             ( u4_col_out_524    ),
    .col_out_525             ( u4_col_out_525    ),
    .col_out_526             ( u4_col_out_526    ),
    .col_out_527             ( u4_col_out_527    ),
    .col_out_528             ( u4_col_out_528    ),
    .col_out_529             ( u4_col_out_529    ),
    .col_out_530             ( u4_col_out_530    ),
    .col_out_531             ( u4_col_out_531    ),
    .col_out_532             ( u4_col_out_532    ),
    .col_out_533             ( u4_col_out_533    ),
    .col_out_534             ( u4_col_out_534    ),
    .col_out_535             ( u4_col_out_535    ),
    .col_out_536             ( u4_col_out_536    ),
    .col_out_537             ( u4_col_out_537    ),
    .col_out_538             ( u4_col_out_538    ),
    .col_out_539             ( u4_col_out_539    ),
    .col_out_540             ( u4_col_out_540    ),
    .col_out_541             ( u4_col_out_541    ),
    .col_out_542             ( u4_col_out_542    ),
    .col_out_543             ( u4_col_out_543    ),
    .col_out_544             ( u4_col_out_544    ),
    .col_out_545             ( u4_col_out_545    ),
    .col_out_546             ( u4_col_out_546    ),
    .col_out_547             ( u4_col_out_547    ),
    .col_out_548             ( u4_col_out_548    ),
    .col_out_549             ( u4_col_out_549    ),
    .col_out_550             ( u4_col_out_550    ),
    .col_out_551             ( u4_col_out_551    ),
    .col_out_552             ( u4_col_out_552    ),
    .col_out_553             ( u4_col_out_553    ),
    .col_out_554             ( u4_col_out_554    ),
    .col_out_555             ( u4_col_out_555    ),
    .col_out_556             ( u4_col_out_556    ),
    .col_out_557             ( u4_col_out_557    ),
    .col_out_558             ( u4_col_out_558    ),
    .col_out_559             ( u4_col_out_559    ),
    .col_out_560             ( u4_col_out_560    ),
    .col_out_561             ( u4_col_out_561    ),
    .col_out_562             ( u4_col_out_562    ),
    .col_out_563             ( u4_col_out_563    ),
    .col_out_564             ( u4_col_out_564    ),
    .col_out_565             ( u4_col_out_565    ),
    .col_out_566             ( u4_col_out_566    ),
    .col_out_567             ( u4_col_out_567    ),
    .col_out_568             ( u4_col_out_568    ),
    .col_out_569             ( u4_col_out_569    ),
    .col_out_570             ( u4_col_out_570    ),
    .col_out_571             ( u4_col_out_571    ),
    .col_out_572             ( u4_col_out_572    ),
    .col_out_573             ( u4_col_out_573    ),
    .col_out_574             ( u4_col_out_574    ),
    .col_out_575             ( u4_col_out_575    ),
    .col_out_576             ( u4_col_out_576    ),
    .col_out_577             ( u4_col_out_577    ),
    .col_out_578             ( u4_col_out_578    ),
    .col_out_579             ( u4_col_out_579    ),
    .col_out_580             ( u4_col_out_580    ),
    .col_out_581             ( u4_col_out_581    ),
    .col_out_582             ( u4_col_out_582    ),
    .col_out_583             ( u4_col_out_583    ),
    .col_out_584             ( u4_col_out_584    ),
    .col_out_585             ( u4_col_out_585    ),
    .col_out_586             ( u4_col_out_586    ),
    .col_out_587             ( u4_col_out_587    ),
    .col_out_588             ( u4_col_out_588    ),
    .col_out_589             ( u4_col_out_589    ),
    .col_out_590             ( u4_col_out_590    ),
    .col_out_591             ( u4_col_out_591    ),
    .col_out_592             ( u4_col_out_592    ),
    .col_out_593             ( u4_col_out_593    ),
    .col_out_594             ( u4_col_out_594    ),
    .col_out_595             ( u4_col_out_595    ),
    .col_out_596             ( u4_col_out_596    ),
    .col_out_597             ( u4_col_out_597    ),
    .col_out_598             ( u4_col_out_598    ),
    .col_out_599             ( u4_col_out_599    ),
    .col_out_600             ( u4_col_out_600    ),
    .col_out_601             ( u4_col_out_601    ),
    .col_out_602             ( u4_col_out_602    ),
    .col_out_603             ( u4_col_out_603    ),
    .col_out_604             ( u4_col_out_604    ),
    .col_out_605             ( u4_col_out_605    ),
    .col_out_606             ( u4_col_out_606    ),
    .col_out_607             ( u4_col_out_607    ),
    .col_out_608             ( u4_col_out_608    ),
    .col_out_609             ( u4_col_out_609    ),
    .col_out_610             ( u4_col_out_610    ),
    .col_out_611             ( u4_col_out_611    ),
    .col_out_612             ( u4_col_out_612    ),
    .col_out_613             ( u4_col_out_613    ),
    .col_out_614             ( u4_col_out_614    ),
    .col_out_615             ( u4_col_out_615    ),
    .col_out_616             ( u4_col_out_616    ),
    .col_out_617             ( u4_col_out_617    ),
    .col_out_618             ( u4_col_out_618    ),
    .col_out_619             ( u4_col_out_619    ),
    .col_out_620             ( u4_col_out_620    ),
    .col_out_621             ( u4_col_out_621    ),
    .col_out_622             ( u4_col_out_622    ),
    .col_out_623             ( u4_col_out_623    ),
    .col_out_624             ( u4_col_out_624    ),
    .col_out_625             ( u4_col_out_625    ),
    .col_out_626             ( u4_col_out_626    ),
    .col_out_627             ( u4_col_out_627    ),
    .col_out_628             ( u4_col_out_628    ),
    .col_out_629             ( u4_col_out_629    ),
    .col_out_630             ( u4_col_out_630    ),
    .col_out_631             ( u4_col_out_631    ),
    .col_out_632             ( u4_col_out_632    ),
    .col_out_633             ( u4_col_out_633    ),
    .col_out_634             ( u4_col_out_634    ),
    .col_out_635             ( u4_col_out_635    ),
    .col_out_636             ( u4_col_out_636    ),
    .col_out_637             ( u4_col_out_637    ),
    .col_out_638             ( u4_col_out_638    ),
    .col_out_639             ( u4_col_out_639    ),
    .col_out_640             ( u4_col_out_640    ),
    .col_out_641             ( u4_col_out_641    ),
    .col_out_642             ( u4_col_out_642    ),
    .col_out_643             ( u4_col_out_643    ),
    .col_out_644             ( u4_col_out_644    ),
    .col_out_645             ( u4_col_out_645    ),
    .col_out_646             ( u4_col_out_646    ),
    .col_out_647             ( u4_col_out_647    ),
    .col_out_648             ( u4_col_out_648    ),
    .col_out_649             ( u4_col_out_649    ),
    .col_out_650             ( u4_col_out_650    ),
    .col_out_651             ( u4_col_out_651    ),
    .col_out_652             ( u4_col_out_652    ),
    .col_out_653             ( u4_col_out_653    ),
    .col_out_654             ( u4_col_out_654    ),
    .col_out_655             ( u4_col_out_655    ),
    .col_out_656             ( u4_col_out_656    ),
    .col_out_657             ( u4_col_out_657    ),
    .col_out_658             ( u4_col_out_658    ),
    .col_out_659             ( u4_col_out_659    ),
    .col_out_660             ( u4_col_out_660    ),
    .col_out_661             ( u4_col_out_661    ),
    .col_out_662             ( u4_col_out_662    ),
    .col_out_663             ( u4_col_out_663    ),
    .col_out_664             ( u4_col_out_664    ),
    .col_out_665             ( u4_col_out_665    ),
    .col_out_666             ( u4_col_out_666    ),
    .col_out_667             ( u4_col_out_667    ),
    .col_out_668             ( u4_col_out_668    ),
    .col_out_669             ( u4_col_out_669    ),
    .col_out_670             ( u4_col_out_670    ),
    .col_out_671             ( u4_col_out_671    ),
    .col_out_672             ( u4_col_out_672    ),
    .col_out_673             ( u4_col_out_673    ),
    .col_out_674             ( u4_col_out_674    ),
    .col_out_675             ( u4_col_out_675    ),
    .col_out_676             ( u4_col_out_676    ),
    .col_out_677             ( u4_col_out_677    ),
    .col_out_678             ( u4_col_out_678    ),
    .col_out_679             ( u4_col_out_679    ),
    .col_out_680             ( u4_col_out_680    ),
    .col_out_681             ( u4_col_out_681    ),
    .col_out_682             ( u4_col_out_682    ),
    .col_out_683             ( u4_col_out_683    ),
    .col_out_684             ( u4_col_out_684    ),
    .col_out_685             ( u4_col_out_685    ),
    .col_out_686             ( u4_col_out_686    ),
    .col_out_687             ( u4_col_out_687    ),
    .col_out_688             ( u4_col_out_688    ),
    .col_out_689             ( u4_col_out_689    ),
    .col_out_690             ( u4_col_out_690    ),
    .col_out_691             ( u4_col_out_691    ),
    .col_out_692             ( u4_col_out_692    ),
    .col_out_693             ( u4_col_out_693    ),
    .col_out_694             ( u4_col_out_694    ),
    .col_out_695             ( u4_col_out_695    ),
    .col_out_696             ( u4_col_out_696    ),
    .col_out_697             ( u4_col_out_697    ),
    .col_out_698             ( u4_col_out_698    ),
    .col_out_699             ( u4_col_out_699    ),
    .col_out_700             ( u4_col_out_700    ),
    .col_out_701             ( u4_col_out_701    ),
    .col_out_702             ( u4_col_out_702    ),
    .col_out_703             ( u4_col_out_703    ),
    .col_out_704             ( u4_col_out_704    ),
    .col_out_705             ( u4_col_out_705    ),
    .col_out_706             ( u4_col_out_706    ),
    .col_out_707             ( u4_col_out_707    ),
    .col_out_708             ( u4_col_out_708    ),
    .col_out_709             ( u4_col_out_709    ),
    .col_out_710             ( u4_col_out_710    ),
    .col_out_711             ( u4_col_out_711    ),
    .col_out_712             ( u4_col_out_712    ),
    .col_out_713             ( u4_col_out_713    ),
    .col_out_714             ( u4_col_out_714    ),
    .col_out_715             ( u4_col_out_715    ),
    .col_out_716             ( u4_col_out_716    ),
    .col_out_717             ( u4_col_out_717    ),
    .col_out_718             ( u4_col_out_718    ),
    .col_out_719             ( u4_col_out_719    ),
    .col_out_720             ( u4_col_out_720    ),
    .col_out_721             ( u4_col_out_721    ),
    .col_out_722             ( u4_col_out_722    ),
    .col_out_723             ( u4_col_out_723    ),
    .col_out_724             ( u4_col_out_724    ),
    .col_out_725             ( u4_col_out_725    ),
    .col_out_726             ( u4_col_out_726    ),
    .col_out_727             ( u4_col_out_727    ),
    .col_out_728             ( u4_col_out_728    ),
    .col_out_729             ( u4_col_out_729    ),
    .col_out_730             ( u4_col_out_730    ),
    .col_out_731             ( u4_col_out_731    ),
    .col_out_732             ( u4_col_out_732    ),
    .col_out_733             ( u4_col_out_733    ),
    .col_out_734             ( u4_col_out_734    ),
    .col_out_735             ( u4_col_out_735    ),
    .col_out_736             ( u4_col_out_736    ),
    .col_out_737             ( u4_col_out_737    ),
    .col_out_738             ( u4_col_out_738    ),
    .col_out_739             ( u4_col_out_739    ),
    .col_out_740             ( u4_col_out_740    ),
    .col_out_741             ( u4_col_out_741    ),
    .col_out_742             ( u4_col_out_742    ),
    .col_out_743             ( u4_col_out_743    ),
    .col_out_744             ( u4_col_out_744    ),
    .col_out_745             ( u4_col_out_745    ),
    .col_out_746             ( u4_col_out_746    ),
    .col_out_747             ( u4_col_out_747    ),
    .col_out_748             ( u4_col_out_748    ),
    .col_out_749             ( u4_col_out_749    ),
    .col_out_750             ( u4_col_out_750    ),
    .col_out_751             ( u4_col_out_751    ),
    .col_out_752             ( u4_col_out_752    ),
    .col_out_753             ( u4_col_out_753    ),
    .col_out_754             ( u4_col_out_754    ),
    .col_out_755             ( u4_col_out_755    ),
    .col_out_756             ( u4_col_out_756    ),
    .col_out_757             ( u4_col_out_757    ),
    .col_out_758             ( u4_col_out_758    ),
    .col_out_759             ( u4_col_out_759    ),
    .col_out_760             ( u4_col_out_760    ),
    .col_out_761             ( u4_col_out_761    ),
    .col_out_762             ( u4_col_out_762    ),
    .col_out_763             ( u4_col_out_763    ),
    .col_out_764             ( u4_col_out_764    ),
    .col_out_765             ( u4_col_out_765    ),
    .col_out_766             ( u4_col_out_766    ),
    .col_out_767             ( u4_col_out_767    ),
    .col_out_768             ( u4_col_out_768    ),
    .col_out_769             ( u4_col_out_769    ),
    .col_out_770             ( u4_col_out_770    ),
    .col_out_771             ( u4_col_out_771    ),
    .col_out_772             ( u4_col_out_772    ),
    .col_out_773             ( u4_col_out_773    ),
    .col_out_774             ( u4_col_out_774    ),
    .col_out_775             ( u4_col_out_775    ),
    .col_out_776             ( u4_col_out_776    ),
    .col_out_777             ( u4_col_out_777    ),
    .col_out_778             ( u4_col_out_778    ),
    .col_out_779             ( u4_col_out_779    ),
    .col_out_780             ( u4_col_out_780    ),
    .col_out_781             ( u4_col_out_781    ),
    .col_out_782             ( u4_col_out_782    ),
    .col_out_783             ( u4_col_out_783    ),
    .col_out_784             ( u4_col_out_784    ),
    .col_out_785             ( u4_col_out_785    ),
    .col_out_786             ( u4_col_out_786    ),
    .col_out_787             ( u4_col_out_787    ),
    .col_out_788             ( u4_col_out_788    ),
    .col_out_789             ( u4_col_out_789    ),
    .col_out_790             ( u4_col_out_790    ),
    .col_out_791             ( u4_col_out_791    ),
    .col_out_792             ( u4_col_out_792    ),
    .col_out_793             ( u4_col_out_793    ),
    .col_out_794             ( u4_col_out_794    ),
    .col_out_795             ( u4_col_out_795    ),
    .col_out_796             ( u4_col_out_796    ),
    .col_out_797             ( u4_col_out_797    ),
    .col_out_798             ( u4_col_out_798    ),
    .col_out_799             ( u4_col_out_799    ),
    .col_out_800             ( u4_col_out_800    ),
    .col_out_801             ( u4_col_out_801    ),
    .col_out_802             ( u4_col_out_802    ),
    .col_out_803             ( u4_col_out_803    ),
    .col_out_804             ( u4_col_out_804    ),
    .col_out_805             ( u4_col_out_805    ),
    .col_out_806             ( u4_col_out_806    ),
    .col_out_807             ( u4_col_out_807    ),
    .col_out_808             ( u4_col_out_808    ),
    .col_out_809             ( u4_col_out_809    ),
    .col_out_810             ( u4_col_out_810    ),
    .col_out_811             ( u4_col_out_811    ),
    .col_out_812             ( u4_col_out_812    ),
    .col_out_813             ( u4_col_out_813    ),
    .col_out_814             ( u4_col_out_814    ),
    .col_out_815             ( u4_col_out_815    ),
    .col_out_816             ( u4_col_out_816    ),
    .col_out_817             ( u4_col_out_817    ),
    .col_out_818             ( u4_col_out_818    ),
    .col_out_819             ( u4_col_out_819    ),
    .col_out_820             ( u4_col_out_820    ),
    .col_out_821             ( u4_col_out_821    ),
    .col_out_822             ( u4_col_out_822    ),
    .col_out_823             ( u4_col_out_823    ),
    .col_out_824             ( u4_col_out_824    ),
    .col_out_825             ( u4_col_out_825    ),
    .col_out_826             ( u4_col_out_826    ),
    .col_out_827             ( u4_col_out_827    ),
    .col_out_828             ( u4_col_out_828    ),
    .col_out_829             ( u4_col_out_829    ),
    .col_out_830             ( u4_col_out_830    ),
    .col_out_831             ( u4_col_out_831    ),
    .col_out_832             ( u4_col_out_832    ),
    .col_out_833             ( u4_col_out_833    ),
    .col_out_834             ( u4_col_out_834    ),
    .col_out_835             ( u4_col_out_835    ),
    .col_out_836             ( u4_col_out_836    ),
    .col_out_837             ( u4_col_out_837    ),
    .col_out_838             ( u4_col_out_838    ),
    .col_out_839             ( u4_col_out_839    ),
    .col_out_840             ( u4_col_out_840    ),
    .col_out_841             ( u4_col_out_841    ),
    .col_out_842             ( u4_col_out_842    ),
    .col_out_843             ( u4_col_out_843    ),
    .col_out_844             ( u4_col_out_844    ),
    .col_out_845             ( u4_col_out_845    ),
    .col_out_846             ( u4_col_out_846    ),
    .col_out_847             ( u4_col_out_847    ),
    .col_out_848             ( u4_col_out_848    ),
    .col_out_849             ( u4_col_out_849    ),
    .col_out_850             ( u4_col_out_850    ),
    .col_out_851             ( u4_col_out_851    ),
    .col_out_852             ( u4_col_out_852    ),
    .col_out_853             ( u4_col_out_853    ),
    .col_out_854             ( u4_col_out_854    ),
    .col_out_855             ( u4_col_out_855    ),
    .col_out_856             ( u4_col_out_856    ),
    .col_out_857             ( u4_col_out_857    ),
    .col_out_858             ( u4_col_out_858    ),
    .col_out_859             ( u4_col_out_859    ),
    .col_out_860             ( u4_col_out_860    ),
    .col_out_861             ( u4_col_out_861    ),
    .col_out_862             ( u4_col_out_862    ),
    .col_out_863             ( u4_col_out_863    ),
    .col_out_864             ( u4_col_out_864    ),
    .col_out_865             ( u4_col_out_865    ),
    .col_out_866             ( u4_col_out_866    ),
    .col_out_867             ( u4_col_out_867    ),
    .col_out_868             ( u4_col_out_868    ),
    .col_out_869             ( u4_col_out_869    ),
    .col_out_870             ( u4_col_out_870    ),
    .col_out_871             ( u4_col_out_871    ),
    .col_out_872             ( u4_col_out_872    ),
    .col_out_873             ( u4_col_out_873    ),
    .col_out_874             ( u4_col_out_874    ),
    .col_out_875             ( u4_col_out_875    ),
    .col_out_876             ( u4_col_out_876    ),
    .col_out_877             ( u4_col_out_877    ),
    .col_out_878             ( u4_col_out_878    ),
    .col_out_879             ( u4_col_out_879    ),
    .col_out_880             ( u4_col_out_880    ),
    .col_out_881             ( u4_col_out_881    ),
    .col_out_882             ( u4_col_out_882    ),
    .col_out_883             ( u4_col_out_883    ),
    .col_out_884             ( u4_col_out_884    ),
    .col_out_885             ( u4_col_out_885    ),
    .col_out_886             ( u4_col_out_886    ),
    .col_out_887             ( u4_col_out_887    ),
    .col_out_888             ( u4_col_out_888    ),
    .col_out_889             ( u4_col_out_889    ),
    .col_out_890             ( u4_col_out_890    ),
    .col_out_891             ( u4_col_out_891    ),
    .col_out_892             ( u4_col_out_892    ),
    .col_out_893             ( u4_col_out_893    ),
    .col_out_894             ( u4_col_out_894    ),
    .col_out_895             ( u4_col_out_895    ),
    .col_out_896             ( u4_col_out_896    ),
    .col_out_897             ( u4_col_out_897    ),
    .col_out_898             ( u4_col_out_898    ),
    .col_out_899             ( u4_col_out_899    ),
    .col_out_900             ( u4_col_out_900    ),
    .col_out_901             ( u4_col_out_901    ),
    .col_out_902             ( u4_col_out_902    ),
    .col_out_903             ( u4_col_out_903    ),
    .col_out_904             ( u4_col_out_904    ),
    .col_out_905             ( u4_col_out_905    ),
    .col_out_906             ( u4_col_out_906    ),
    .col_out_907             ( u4_col_out_907    ),
    .col_out_908             ( u4_col_out_908    ),
    .col_out_909             ( u4_col_out_909    ),
    .col_out_910             ( u4_col_out_910    ),
    .col_out_911             ( u4_col_out_911    ),
    .col_out_912             ( u4_col_out_912    ),
    .col_out_913             ( u4_col_out_913    ),
    .col_out_914             ( u4_col_out_914    ),
    .col_out_915             ( u4_col_out_915    ),
    .col_out_916             ( u4_col_out_916    ),
    .col_out_917             ( u4_col_out_917    ),
    .col_out_918             ( u4_col_out_918    ),
    .col_out_919             ( u4_col_out_919    ),
    .col_out_920             ( u4_col_out_920    ),
    .col_out_921             ( u4_col_out_921    ),
    .col_out_922             ( u4_col_out_922    ),
    .col_out_923             ( u4_col_out_923    ),
    .col_out_924             ( u4_col_out_924    ),
    .col_out_925             ( u4_col_out_925    ),
    .col_out_926             ( u4_col_out_926    ),
    .col_out_927             ( u4_col_out_927    ),
    .col_out_928             ( u4_col_out_928    ),
    .col_out_929             ( u4_col_out_929    ),
    .col_out_930             ( u4_col_out_930    ),
    .col_out_931             ( u4_col_out_931    ),
    .col_out_932             ( u4_col_out_932    ),
    .col_out_933             ( u4_col_out_933    ),
    .col_out_934             ( u4_col_out_934    ),
    .col_out_935             ( u4_col_out_935    ),
    .col_out_936             ( u4_col_out_936    ),
    .col_out_937             ( u4_col_out_937    ),
    .col_out_938             ( u4_col_out_938    ),
    .col_out_939             ( u4_col_out_939    ),
    .col_out_940             ( u4_col_out_940    ),
    .col_out_941             ( u4_col_out_941    ),
    .col_out_942             ( u4_col_out_942    ),
    .col_out_943             ( u4_col_out_943    ),
    .col_out_944             ( u4_col_out_944    ),
    .col_out_945             ( u4_col_out_945    ),
    .col_out_946             ( u4_col_out_946    ),
    .col_out_947             ( u4_col_out_947    ),
    .col_out_948             ( u4_col_out_948    ),
    .col_out_949             ( u4_col_out_949    ),
    .col_out_950             ( u4_col_out_950    ),
    .col_out_951             ( u4_col_out_951    ),
    .col_out_952             ( u4_col_out_952    ),
    .col_out_953             ( u4_col_out_953    ),
    .col_out_954             ( u4_col_out_954    ),
    .col_out_955             ( u4_col_out_955    ),
    .col_out_956             ( u4_col_out_956    ),
    .col_out_957             ( u4_col_out_957    ),
    .col_out_958             ( u4_col_out_958    ),
    .col_out_959             ( u4_col_out_959    ),
    .col_out_960             ( u4_col_out_960    ),
    .col_out_961             ( u4_col_out_961    ),
    .col_out_962             ( u4_col_out_962    ),
    .col_out_963             ( u4_col_out_963    ),
    .col_out_964             ( u4_col_out_964    ),
    .col_out_965             ( u4_col_out_965    ),
    .col_out_966             ( u4_col_out_966    ),
    .col_out_967             ( u4_col_out_967    ),
    .col_out_968             ( u4_col_out_968    ),
    .col_out_969             ( u4_col_out_969    ),
    .col_out_970             ( u4_col_out_970    ),
    .col_out_971             ( u4_col_out_971    ),
    .col_out_972             ( u4_col_out_972    ),
    .col_out_973             ( u4_col_out_973    ),
    .col_out_974             ( u4_col_out_974    ),
    .col_out_975             ( u4_col_out_975    ),
    .col_out_976             ( u4_col_out_976    ),
    .col_out_977             ( u4_col_out_977    ),
    .col_out_978             ( u4_col_out_978    ),
    .col_out_979             ( u4_col_out_979    ),
    .col_out_980             ( u4_col_out_980    ),
    .col_out_981             ( u4_col_out_981    ),
    .col_out_982             ( u4_col_out_982    ),
    .col_out_983             ( u4_col_out_983    ),
    .col_out_984             ( u4_col_out_984    ),
    .col_out_985             ( u4_col_out_985    ),
    .col_out_986             ( u4_col_out_986    ),
    .col_out_987             ( u4_col_out_987    ),
    .col_out_988             ( u4_col_out_988    ),
    .col_out_989             ( u4_col_out_989    ),
    .col_out_990             ( u4_col_out_990    ),
    .col_out_991             ( u4_col_out_991    ),
    .col_out_992             ( u4_col_out_992    ),
    .col_out_993             ( u4_col_out_993    ),
    .col_out_994             ( u4_col_out_994    ),
    .col_out_995             ( u4_col_out_995    ),
    .col_out_996             ( u4_col_out_996    ),
    .col_out_997             ( u4_col_out_997    ),
    .col_out_998             ( u4_col_out_998    ),
    .col_out_999             ( u4_col_out_999    ),
    .col_out_1000            ( u4_col_out_1000   ),
    .col_out_1001            ( u4_col_out_1001   ),
    .col_out_1002            ( u4_col_out_1002   ),
    .col_out_1003            ( u4_col_out_1003   ),
    .col_out_1004            ( u4_col_out_1004   ),
    .col_out_1005            ( u4_col_out_1005   ),
    .col_out_1006            ( u4_col_out_1006   ),
    .col_out_1007            ( u4_col_out_1007   ),
    .col_out_1008            ( u4_col_out_1008   ),
    .col_out_1009            ( u4_col_out_1009   ),
    .col_out_1010            ( u4_col_out_1010   ),
    .col_out_1011            ( u4_col_out_1011   ),
    .col_out_1012            ( u4_col_out_1012   ),
    .col_out_1013            ( u4_col_out_1013   ),
    .col_out_1014            ( u4_col_out_1014   ),
    .col_out_1015            ( u4_col_out_1015   ),
    .col_out_1016            ( u4_col_out_1016   ),
    .col_out_1017            ( u4_col_out_1017   ),
    .col_out_1018            ( u4_col_out_1018   ),
    .col_out_1019            ( u4_col_out_1019   ),
    .col_out_1020            ( u4_col_out_1020   ),
    .col_out_1021            ( u4_col_out_1021   ),
    .col_out_1022            ( u4_col_out_1022   ),
    .col_out_1023            ( u4_col_out_1023   ),
    .col_out_1024            ( u4_col_out_1024   ),
    .col_out_1025            ( u4_col_out_1025   ),
    .col_out_1026            ( u4_col_out_1026   ),
    .col_out_1027            ( u4_col_out_1027   ),
    .col_out_1028            ( u4_col_out_1028   ),
    .col_out_1029            ( u4_col_out_1029   ),
    .col_out_1030            ( u4_col_out_1030   ),
    .col_out_1031            ( u4_col_out_1031   ),
    .col_out_1032            ( u4_col_out_1032   ),
    .col_out_1033            ( u4_col_out_1033   )
);




// compressor_array_3_2_1033 Outputs
wire  [1:0]  u5_col_out_0;
wire  [1:0]  u5_col_out_1;
wire  [1:0]  u5_col_out_2;
wire  [1:0]  u5_col_out_3;
wire  [1:0]  u5_col_out_4;
wire  [1:0]  u5_col_out_5;
wire  [1:0]  u5_col_out_6;
wire  [1:0]  u5_col_out_7;
wire  [1:0]  u5_col_out_8;
wire  [1:0]  u5_col_out_9;
wire  [1:0]  u5_col_out_10;
wire  [1:0]  u5_col_out_11;
wire  [1:0]  u5_col_out_12;
wire  [1:0]  u5_col_out_13;
wire  [1:0]  u5_col_out_14;
wire  [1:0]  u5_col_out_15;
wire  [1:0]  u5_col_out_16;
wire  [1:0]  u5_col_out_17;
wire  [1:0]  u5_col_out_18;
wire  [1:0]  u5_col_out_19;
wire  [1:0]  u5_col_out_20;
wire  [1:0]  u5_col_out_21;
wire  [1:0]  u5_col_out_22;
wire  [1:0]  u5_col_out_23;
wire  [1:0]  u5_col_out_24;
wire  [1:0]  u5_col_out_25;
wire  [1:0]  u5_col_out_26;
wire  [1:0]  u5_col_out_27;
wire  [1:0]  u5_col_out_28;
wire  [1:0]  u5_col_out_29;
wire  [1:0]  u5_col_out_30;
wire  [1:0]  u5_col_out_31;
wire  [1:0]  u5_col_out_32;
wire  [1:0]  u5_col_out_33;
wire  [1:0]  u5_col_out_34;
wire  [1:0]  u5_col_out_35;
wire  [1:0]  u5_col_out_36;
wire  [1:0]  u5_col_out_37;
wire  [1:0]  u5_col_out_38;
wire  [1:0]  u5_col_out_39;
wire  [1:0]  u5_col_out_40;
wire  [1:0]  u5_col_out_41;
wire  [1:0]  u5_col_out_42;
wire  [1:0]  u5_col_out_43;
wire  [1:0]  u5_col_out_44;
wire  [1:0]  u5_col_out_45;
wire  [1:0]  u5_col_out_46;
wire  [1:0]  u5_col_out_47;
wire  [1:0]  u5_col_out_48;
wire  [1:0]  u5_col_out_49;
wire  [1:0]  u5_col_out_50;
wire  [1:0]  u5_col_out_51;
wire  [1:0]  u5_col_out_52;
wire  [1:0]  u5_col_out_53;
wire  [1:0]  u5_col_out_54;
wire  [1:0]  u5_col_out_55;
wire  [1:0]  u5_col_out_56;
wire  [1:0]  u5_col_out_57;
wire  [1:0]  u5_col_out_58;
wire  [1:0]  u5_col_out_59;
wire  [1:0]  u5_col_out_60;
wire  [1:0]  u5_col_out_61;
wire  [1:0]  u5_col_out_62;
wire  [1:0]  u5_col_out_63;
wire  [1:0]  u5_col_out_64;
wire  [1:0]  u5_col_out_65;
wire  [1:0]  u5_col_out_66;
wire  [1:0]  u5_col_out_67;
wire  [1:0]  u5_col_out_68;
wire  [1:0]  u5_col_out_69;
wire  [1:0]  u5_col_out_70;
wire  [1:0]  u5_col_out_71;
wire  [1:0]  u5_col_out_72;
wire  [1:0]  u5_col_out_73;
wire  [1:0]  u5_col_out_74;
wire  [1:0]  u5_col_out_75;
wire  [1:0]  u5_col_out_76;
wire  [1:0]  u5_col_out_77;
wire  [1:0]  u5_col_out_78;
wire  [1:0]  u5_col_out_79;
wire  [1:0]  u5_col_out_80;
wire  [1:0]  u5_col_out_81;
wire  [1:0]  u5_col_out_82;
wire  [1:0]  u5_col_out_83;
wire  [1:0]  u5_col_out_84;
wire  [1:0]  u5_col_out_85;
wire  [1:0]  u5_col_out_86;
wire  [1:0]  u5_col_out_87;
wire  [1:0]  u5_col_out_88;
wire  [1:0]  u5_col_out_89;
wire  [1:0]  u5_col_out_90;
wire  [1:0]  u5_col_out_91;
wire  [1:0]  u5_col_out_92;
wire  [1:0]  u5_col_out_93;
wire  [1:0]  u5_col_out_94;
wire  [1:0]  u5_col_out_95;
wire  [1:0]  u5_col_out_96;
wire  [1:0]  u5_col_out_97;
wire  [1:0]  u5_col_out_98;
wire  [1:0]  u5_col_out_99;
wire  [1:0]  u5_col_out_100;
wire  [1:0]  u5_col_out_101;
wire  [1:0]  u5_col_out_102;
wire  [1:0]  u5_col_out_103;
wire  [1:0]  u5_col_out_104;
wire  [1:0]  u5_col_out_105;
wire  [1:0]  u5_col_out_106;
wire  [1:0]  u5_col_out_107;
wire  [1:0]  u5_col_out_108;
wire  [1:0]  u5_col_out_109;
wire  [1:0]  u5_col_out_110;
wire  [1:0]  u5_col_out_111;
wire  [1:0]  u5_col_out_112;
wire  [1:0]  u5_col_out_113;
wire  [1:0]  u5_col_out_114;
wire  [1:0]  u5_col_out_115;
wire  [1:0]  u5_col_out_116;
wire  [1:0]  u5_col_out_117;
wire  [1:0]  u5_col_out_118;
wire  [1:0]  u5_col_out_119;
wire  [1:0]  u5_col_out_120;
wire  [1:0]  u5_col_out_121;
wire  [1:0]  u5_col_out_122;
wire  [1:0]  u5_col_out_123;
wire  [1:0]  u5_col_out_124;
wire  [1:0]  u5_col_out_125;
wire  [1:0]  u5_col_out_126;
wire  [1:0]  u5_col_out_127;
wire  [1:0]  u5_col_out_128;
wire  [1:0]  u5_col_out_129;
wire  [1:0]  u5_col_out_130;
wire  [1:0]  u5_col_out_131;
wire  [1:0]  u5_col_out_132;
wire  [1:0]  u5_col_out_133;
wire  [1:0]  u5_col_out_134;
wire  [1:0]  u5_col_out_135;
wire  [1:0]  u5_col_out_136;
wire  [1:0]  u5_col_out_137;
wire  [1:0]  u5_col_out_138;
wire  [1:0]  u5_col_out_139;
wire  [1:0]  u5_col_out_140;
wire  [1:0]  u5_col_out_141;
wire  [1:0]  u5_col_out_142;
wire  [1:0]  u5_col_out_143;
wire  [1:0]  u5_col_out_144;
wire  [1:0]  u5_col_out_145;
wire  [1:0]  u5_col_out_146;
wire  [1:0]  u5_col_out_147;
wire  [1:0]  u5_col_out_148;
wire  [1:0]  u5_col_out_149;
wire  [1:0]  u5_col_out_150;
wire  [1:0]  u5_col_out_151;
wire  [1:0]  u5_col_out_152;
wire  [1:0]  u5_col_out_153;
wire  [1:0]  u5_col_out_154;
wire  [1:0]  u5_col_out_155;
wire  [1:0]  u5_col_out_156;
wire  [1:0]  u5_col_out_157;
wire  [1:0]  u5_col_out_158;
wire  [1:0]  u5_col_out_159;
wire  [1:0]  u5_col_out_160;
wire  [1:0]  u5_col_out_161;
wire  [1:0]  u5_col_out_162;
wire  [1:0]  u5_col_out_163;
wire  [1:0]  u5_col_out_164;
wire  [1:0]  u5_col_out_165;
wire  [1:0]  u5_col_out_166;
wire  [1:0]  u5_col_out_167;
wire  [1:0]  u5_col_out_168;
wire  [1:0]  u5_col_out_169;
wire  [1:0]  u5_col_out_170;
wire  [1:0]  u5_col_out_171;
wire  [1:0]  u5_col_out_172;
wire  [1:0]  u5_col_out_173;
wire  [1:0]  u5_col_out_174;
wire  [1:0]  u5_col_out_175;
wire  [1:0]  u5_col_out_176;
wire  [1:0]  u5_col_out_177;
wire  [1:0]  u5_col_out_178;
wire  [1:0]  u5_col_out_179;
wire  [1:0]  u5_col_out_180;
wire  [1:0]  u5_col_out_181;
wire  [1:0]  u5_col_out_182;
wire  [1:0]  u5_col_out_183;
wire  [1:0]  u5_col_out_184;
wire  [1:0]  u5_col_out_185;
wire  [1:0]  u5_col_out_186;
wire  [1:0]  u5_col_out_187;
wire  [1:0]  u5_col_out_188;
wire  [1:0]  u5_col_out_189;
wire  [1:0]  u5_col_out_190;
wire  [1:0]  u5_col_out_191;
wire  [1:0]  u5_col_out_192;
wire  [1:0]  u5_col_out_193;
wire  [1:0]  u5_col_out_194;
wire  [1:0]  u5_col_out_195;
wire  [1:0]  u5_col_out_196;
wire  [1:0]  u5_col_out_197;
wire  [1:0]  u5_col_out_198;
wire  [1:0]  u5_col_out_199;
wire  [1:0]  u5_col_out_200;
wire  [1:0]  u5_col_out_201;
wire  [1:0]  u5_col_out_202;
wire  [1:0]  u5_col_out_203;
wire  [1:0]  u5_col_out_204;
wire  [1:0]  u5_col_out_205;
wire  [1:0]  u5_col_out_206;
wire  [1:0]  u5_col_out_207;
wire  [1:0]  u5_col_out_208;
wire  [1:0]  u5_col_out_209;
wire  [1:0]  u5_col_out_210;
wire  [1:0]  u5_col_out_211;
wire  [1:0]  u5_col_out_212;
wire  [1:0]  u5_col_out_213;
wire  [1:0]  u5_col_out_214;
wire  [1:0]  u5_col_out_215;
wire  [1:0]  u5_col_out_216;
wire  [1:0]  u5_col_out_217;
wire  [1:0]  u5_col_out_218;
wire  [1:0]  u5_col_out_219;
wire  [1:0]  u5_col_out_220;
wire  [1:0]  u5_col_out_221;
wire  [1:0]  u5_col_out_222;
wire  [1:0]  u5_col_out_223;
wire  [1:0]  u5_col_out_224;
wire  [1:0]  u5_col_out_225;
wire  [1:0]  u5_col_out_226;
wire  [1:0]  u5_col_out_227;
wire  [1:0]  u5_col_out_228;
wire  [1:0]  u5_col_out_229;
wire  [1:0]  u5_col_out_230;
wire  [1:0]  u5_col_out_231;
wire  [1:0]  u5_col_out_232;
wire  [1:0]  u5_col_out_233;
wire  [1:0]  u5_col_out_234;
wire  [1:0]  u5_col_out_235;
wire  [1:0]  u5_col_out_236;
wire  [1:0]  u5_col_out_237;
wire  [1:0]  u5_col_out_238;
wire  [1:0]  u5_col_out_239;
wire  [1:0]  u5_col_out_240;
wire  [1:0]  u5_col_out_241;
wire  [1:0]  u5_col_out_242;
wire  [1:0]  u5_col_out_243;
wire  [1:0]  u5_col_out_244;
wire  [1:0]  u5_col_out_245;
wire  [1:0]  u5_col_out_246;
wire  [1:0]  u5_col_out_247;
wire  [1:0]  u5_col_out_248;
wire  [1:0]  u5_col_out_249;
wire  [1:0]  u5_col_out_250;
wire  [1:0]  u5_col_out_251;
wire  [1:0]  u5_col_out_252;
wire  [1:0]  u5_col_out_253;
wire  [1:0]  u5_col_out_254;
wire  [1:0]  u5_col_out_255;
wire  [1:0]  u5_col_out_256;
wire  [1:0]  u5_col_out_257;
wire  [1:0]  u5_col_out_258;
wire  [1:0]  u5_col_out_259;
wire  [1:0]  u5_col_out_260;
wire  [1:0]  u5_col_out_261;
wire  [1:0]  u5_col_out_262;
wire  [1:0]  u5_col_out_263;
wire  [1:0]  u5_col_out_264;
wire  [1:0]  u5_col_out_265;
wire  [1:0]  u5_col_out_266;
wire  [1:0]  u5_col_out_267;
wire  [1:0]  u5_col_out_268;
wire  [1:0]  u5_col_out_269;
wire  [1:0]  u5_col_out_270;
wire  [1:0]  u5_col_out_271;
wire  [1:0]  u5_col_out_272;
wire  [1:0]  u5_col_out_273;
wire  [1:0]  u5_col_out_274;
wire  [1:0]  u5_col_out_275;
wire  [1:0]  u5_col_out_276;
wire  [1:0]  u5_col_out_277;
wire  [1:0]  u5_col_out_278;
wire  [1:0]  u5_col_out_279;
wire  [1:0]  u5_col_out_280;
wire  [1:0]  u5_col_out_281;
wire  [1:0]  u5_col_out_282;
wire  [1:0]  u5_col_out_283;
wire  [1:0]  u5_col_out_284;
wire  [1:0]  u5_col_out_285;
wire  [1:0]  u5_col_out_286;
wire  [1:0]  u5_col_out_287;
wire  [1:0]  u5_col_out_288;
wire  [1:0]  u5_col_out_289;
wire  [1:0]  u5_col_out_290;
wire  [1:0]  u5_col_out_291;
wire  [1:0]  u5_col_out_292;
wire  [1:0]  u5_col_out_293;
wire  [1:0]  u5_col_out_294;
wire  [1:0]  u5_col_out_295;
wire  [1:0]  u5_col_out_296;
wire  [1:0]  u5_col_out_297;
wire  [1:0]  u5_col_out_298;
wire  [1:0]  u5_col_out_299;
wire  [1:0]  u5_col_out_300;
wire  [1:0]  u5_col_out_301;
wire  [1:0]  u5_col_out_302;
wire  [1:0]  u5_col_out_303;
wire  [1:0]  u5_col_out_304;
wire  [1:0]  u5_col_out_305;
wire  [1:0]  u5_col_out_306;
wire  [1:0]  u5_col_out_307;
wire  [1:0]  u5_col_out_308;
wire  [1:0]  u5_col_out_309;
wire  [1:0]  u5_col_out_310;
wire  [1:0]  u5_col_out_311;
wire  [1:0]  u5_col_out_312;
wire  [1:0]  u5_col_out_313;
wire  [1:0]  u5_col_out_314;
wire  [1:0]  u5_col_out_315;
wire  [1:0]  u5_col_out_316;
wire  [1:0]  u5_col_out_317;
wire  [1:0]  u5_col_out_318;
wire  [1:0]  u5_col_out_319;
wire  [1:0]  u5_col_out_320;
wire  [1:0]  u5_col_out_321;
wire  [1:0]  u5_col_out_322;
wire  [1:0]  u5_col_out_323;
wire  [1:0]  u5_col_out_324;
wire  [1:0]  u5_col_out_325;
wire  [1:0]  u5_col_out_326;
wire  [1:0]  u5_col_out_327;
wire  [1:0]  u5_col_out_328;
wire  [1:0]  u5_col_out_329;
wire  [1:0]  u5_col_out_330;
wire  [1:0]  u5_col_out_331;
wire  [1:0]  u5_col_out_332;
wire  [1:0]  u5_col_out_333;
wire  [1:0]  u5_col_out_334;
wire  [1:0]  u5_col_out_335;
wire  [1:0]  u5_col_out_336;
wire  [1:0]  u5_col_out_337;
wire  [1:0]  u5_col_out_338;
wire  [1:0]  u5_col_out_339;
wire  [1:0]  u5_col_out_340;
wire  [1:0]  u5_col_out_341;
wire  [1:0]  u5_col_out_342;
wire  [1:0]  u5_col_out_343;
wire  [1:0]  u5_col_out_344;
wire  [1:0]  u5_col_out_345;
wire  [1:0]  u5_col_out_346;
wire  [1:0]  u5_col_out_347;
wire  [1:0]  u5_col_out_348;
wire  [1:0]  u5_col_out_349;
wire  [1:0]  u5_col_out_350;
wire  [1:0]  u5_col_out_351;
wire  [1:0]  u5_col_out_352;
wire  [1:0]  u5_col_out_353;
wire  [1:0]  u5_col_out_354;
wire  [1:0]  u5_col_out_355;
wire  [1:0]  u5_col_out_356;
wire  [1:0]  u5_col_out_357;
wire  [1:0]  u5_col_out_358;
wire  [1:0]  u5_col_out_359;
wire  [1:0]  u5_col_out_360;
wire  [1:0]  u5_col_out_361;
wire  [1:0]  u5_col_out_362;
wire  [1:0]  u5_col_out_363;
wire  [1:0]  u5_col_out_364;
wire  [1:0]  u5_col_out_365;
wire  [1:0]  u5_col_out_366;
wire  [1:0]  u5_col_out_367;
wire  [1:0]  u5_col_out_368;
wire  [1:0]  u5_col_out_369;
wire  [1:0]  u5_col_out_370;
wire  [1:0]  u5_col_out_371;
wire  [1:0]  u5_col_out_372;
wire  [1:0]  u5_col_out_373;
wire  [1:0]  u5_col_out_374;
wire  [1:0]  u5_col_out_375;
wire  [1:0]  u5_col_out_376;
wire  [1:0]  u5_col_out_377;
wire  [1:0]  u5_col_out_378;
wire  [1:0]  u5_col_out_379;
wire  [1:0]  u5_col_out_380;
wire  [1:0]  u5_col_out_381;
wire  [1:0]  u5_col_out_382;
wire  [1:0]  u5_col_out_383;
wire  [1:0]  u5_col_out_384;
wire  [1:0]  u5_col_out_385;
wire  [1:0]  u5_col_out_386;
wire  [1:0]  u5_col_out_387;
wire  [1:0]  u5_col_out_388;
wire  [1:0]  u5_col_out_389;
wire  [1:0]  u5_col_out_390;
wire  [1:0]  u5_col_out_391;
wire  [1:0]  u5_col_out_392;
wire  [1:0]  u5_col_out_393;
wire  [1:0]  u5_col_out_394;
wire  [1:0]  u5_col_out_395;
wire  [1:0]  u5_col_out_396;
wire  [1:0]  u5_col_out_397;
wire  [1:0]  u5_col_out_398;
wire  [1:0]  u5_col_out_399;
wire  [1:0]  u5_col_out_400;
wire  [1:0]  u5_col_out_401;
wire  [1:0]  u5_col_out_402;
wire  [1:0]  u5_col_out_403;
wire  [1:0]  u5_col_out_404;
wire  [1:0]  u5_col_out_405;
wire  [1:0]  u5_col_out_406;
wire  [1:0]  u5_col_out_407;
wire  [1:0]  u5_col_out_408;
wire  [1:0]  u5_col_out_409;
wire  [1:0]  u5_col_out_410;
wire  [1:0]  u5_col_out_411;
wire  [1:0]  u5_col_out_412;
wire  [1:0]  u5_col_out_413;
wire  [1:0]  u5_col_out_414;
wire  [1:0]  u5_col_out_415;
wire  [1:0]  u5_col_out_416;
wire  [1:0]  u5_col_out_417;
wire  [1:0]  u5_col_out_418;
wire  [1:0]  u5_col_out_419;
wire  [1:0]  u5_col_out_420;
wire  [1:0]  u5_col_out_421;
wire  [1:0]  u5_col_out_422;
wire  [1:0]  u5_col_out_423;
wire  [1:0]  u5_col_out_424;
wire  [1:0]  u5_col_out_425;
wire  [1:0]  u5_col_out_426;
wire  [1:0]  u5_col_out_427;
wire  [1:0]  u5_col_out_428;
wire  [1:0]  u5_col_out_429;
wire  [1:0]  u5_col_out_430;
wire  [1:0]  u5_col_out_431;
wire  [1:0]  u5_col_out_432;
wire  [1:0]  u5_col_out_433;
wire  [1:0]  u5_col_out_434;
wire  [1:0]  u5_col_out_435;
wire  [1:0]  u5_col_out_436;
wire  [1:0]  u5_col_out_437;
wire  [1:0]  u5_col_out_438;
wire  [1:0]  u5_col_out_439;
wire  [1:0]  u5_col_out_440;
wire  [1:0]  u5_col_out_441;
wire  [1:0]  u5_col_out_442;
wire  [1:0]  u5_col_out_443;
wire  [1:0]  u5_col_out_444;
wire  [1:0]  u5_col_out_445;
wire  [1:0]  u5_col_out_446;
wire  [1:0]  u5_col_out_447;
wire  [1:0]  u5_col_out_448;
wire  [1:0]  u5_col_out_449;
wire  [1:0]  u5_col_out_450;
wire  [1:0]  u5_col_out_451;
wire  [1:0]  u5_col_out_452;
wire  [1:0]  u5_col_out_453;
wire  [1:0]  u5_col_out_454;
wire  [1:0]  u5_col_out_455;
wire  [1:0]  u5_col_out_456;
wire  [1:0]  u5_col_out_457;
wire  [1:0]  u5_col_out_458;
wire  [1:0]  u5_col_out_459;
wire  [1:0]  u5_col_out_460;
wire  [1:0]  u5_col_out_461;
wire  [1:0]  u5_col_out_462;
wire  [1:0]  u5_col_out_463;
wire  [1:0]  u5_col_out_464;
wire  [1:0]  u5_col_out_465;
wire  [1:0]  u5_col_out_466;
wire  [1:0]  u5_col_out_467;
wire  [1:0]  u5_col_out_468;
wire  [1:0]  u5_col_out_469;
wire  [1:0]  u5_col_out_470;
wire  [1:0]  u5_col_out_471;
wire  [1:0]  u5_col_out_472;
wire  [1:0]  u5_col_out_473;
wire  [1:0]  u5_col_out_474;
wire  [1:0]  u5_col_out_475;
wire  [1:0]  u5_col_out_476;
wire  [1:0]  u5_col_out_477;
wire  [1:0]  u5_col_out_478;
wire  [1:0]  u5_col_out_479;
wire  [1:0]  u5_col_out_480;
wire  [1:0]  u5_col_out_481;
wire  [1:0]  u5_col_out_482;
wire  [1:0]  u5_col_out_483;
wire  [1:0]  u5_col_out_484;
wire  [1:0]  u5_col_out_485;
wire  [1:0]  u5_col_out_486;
wire  [1:0]  u5_col_out_487;
wire  [1:0]  u5_col_out_488;
wire  [1:0]  u5_col_out_489;
wire  [1:0]  u5_col_out_490;
wire  [1:0]  u5_col_out_491;
wire  [1:0]  u5_col_out_492;
wire  [1:0]  u5_col_out_493;
wire  [1:0]  u5_col_out_494;
wire  [1:0]  u5_col_out_495;
wire  [1:0]  u5_col_out_496;
wire  [1:0]  u5_col_out_497;
wire  [1:0]  u5_col_out_498;
wire  [1:0]  u5_col_out_499;
wire  [1:0]  u5_col_out_500;
wire  [1:0]  u5_col_out_501;
wire  [1:0]  u5_col_out_502;
wire  [1:0]  u5_col_out_503;
wire  [1:0]  u5_col_out_504;
wire  [1:0]  u5_col_out_505;
wire  [1:0]  u5_col_out_506;
wire  [1:0]  u5_col_out_507;
wire  [1:0]  u5_col_out_508;
wire  [1:0]  u5_col_out_509;
wire  [1:0]  u5_col_out_510;
wire  [1:0]  u5_col_out_511;
wire  [1:0]  u5_col_out_512;
wire  [1:0]  u5_col_out_513;
wire  [1:0]  u5_col_out_514;
wire  [1:0]  u5_col_out_515;
wire  [1:0]  u5_col_out_516;
wire  [1:0]  u5_col_out_517;
wire  [1:0]  u5_col_out_518;
wire  [1:0]  u5_col_out_519;
wire  [1:0]  u5_col_out_520;
wire  [1:0]  u5_col_out_521;
wire  [1:0]  u5_col_out_522;
wire  [1:0]  u5_col_out_523;
wire  [1:0]  u5_col_out_524;
wire  [1:0]  u5_col_out_525;
wire  [1:0]  u5_col_out_526;
wire  [1:0]  u5_col_out_527;
wire  [1:0]  u5_col_out_528;
wire  [1:0]  u5_col_out_529;
wire  [1:0]  u5_col_out_530;
wire  [1:0]  u5_col_out_531;
wire  [1:0]  u5_col_out_532;
wire  [1:0]  u5_col_out_533;
wire  [1:0]  u5_col_out_534;
wire  [1:0]  u5_col_out_535;
wire  [1:0]  u5_col_out_536;
wire  [1:0]  u5_col_out_537;
wire  [1:0]  u5_col_out_538;
wire  [1:0]  u5_col_out_539;
wire  [1:0]  u5_col_out_540;
wire  [1:0]  u5_col_out_541;
wire  [1:0]  u5_col_out_542;
wire  [1:0]  u5_col_out_543;
wire  [1:0]  u5_col_out_544;
wire  [1:0]  u5_col_out_545;
wire  [1:0]  u5_col_out_546;
wire  [1:0]  u5_col_out_547;
wire  [1:0]  u5_col_out_548;
wire  [1:0]  u5_col_out_549;
wire  [1:0]  u5_col_out_550;
wire  [1:0]  u5_col_out_551;
wire  [1:0]  u5_col_out_552;
wire  [1:0]  u5_col_out_553;
wire  [1:0]  u5_col_out_554;
wire  [1:0]  u5_col_out_555;
wire  [1:0]  u5_col_out_556;
wire  [1:0]  u5_col_out_557;
wire  [1:0]  u5_col_out_558;
wire  [1:0]  u5_col_out_559;
wire  [1:0]  u5_col_out_560;
wire  [1:0]  u5_col_out_561;
wire  [1:0]  u5_col_out_562;
wire  [1:0]  u5_col_out_563;
wire  [1:0]  u5_col_out_564;
wire  [1:0]  u5_col_out_565;
wire  [1:0]  u5_col_out_566;
wire  [1:0]  u5_col_out_567;
wire  [1:0]  u5_col_out_568;
wire  [1:0]  u5_col_out_569;
wire  [1:0]  u5_col_out_570;
wire  [1:0]  u5_col_out_571;
wire  [1:0]  u5_col_out_572;
wire  [1:0]  u5_col_out_573;
wire  [1:0]  u5_col_out_574;
wire  [1:0]  u5_col_out_575;
wire  [1:0]  u5_col_out_576;
wire  [1:0]  u5_col_out_577;
wire  [1:0]  u5_col_out_578;
wire  [1:0]  u5_col_out_579;
wire  [1:0]  u5_col_out_580;
wire  [1:0]  u5_col_out_581;
wire  [1:0]  u5_col_out_582;
wire  [1:0]  u5_col_out_583;
wire  [1:0]  u5_col_out_584;
wire  [1:0]  u5_col_out_585;
wire  [1:0]  u5_col_out_586;
wire  [1:0]  u5_col_out_587;
wire  [1:0]  u5_col_out_588;
wire  [1:0]  u5_col_out_589;
wire  [1:0]  u5_col_out_590;
wire  [1:0]  u5_col_out_591;
wire  [1:0]  u5_col_out_592;
wire  [1:0]  u5_col_out_593;
wire  [1:0]  u5_col_out_594;
wire  [1:0]  u5_col_out_595;
wire  [1:0]  u5_col_out_596;
wire  [1:0]  u5_col_out_597;
wire  [1:0]  u5_col_out_598;
wire  [1:0]  u5_col_out_599;
wire  [1:0]  u5_col_out_600;
wire  [1:0]  u5_col_out_601;
wire  [1:0]  u5_col_out_602;
wire  [1:0]  u5_col_out_603;
wire  [1:0]  u5_col_out_604;
wire  [1:0]  u5_col_out_605;
wire  [1:0]  u5_col_out_606;
wire  [1:0]  u5_col_out_607;
wire  [1:0]  u5_col_out_608;
wire  [1:0]  u5_col_out_609;
wire  [1:0]  u5_col_out_610;
wire  [1:0]  u5_col_out_611;
wire  [1:0]  u5_col_out_612;
wire  [1:0]  u5_col_out_613;
wire  [1:0]  u5_col_out_614;
wire  [1:0]  u5_col_out_615;
wire  [1:0]  u5_col_out_616;
wire  [1:0]  u5_col_out_617;
wire  [1:0]  u5_col_out_618;
wire  [1:0]  u5_col_out_619;
wire  [1:0]  u5_col_out_620;
wire  [1:0]  u5_col_out_621;
wire  [1:0]  u5_col_out_622;
wire  [1:0]  u5_col_out_623;
wire  [1:0]  u5_col_out_624;
wire  [1:0]  u5_col_out_625;
wire  [1:0]  u5_col_out_626;
wire  [1:0]  u5_col_out_627;
wire  [1:0]  u5_col_out_628;
wire  [1:0]  u5_col_out_629;
wire  [1:0]  u5_col_out_630;
wire  [1:0]  u5_col_out_631;
wire  [1:0]  u5_col_out_632;
wire  [1:0]  u5_col_out_633;
wire  [1:0]  u5_col_out_634;
wire  [1:0]  u5_col_out_635;
wire  [1:0]  u5_col_out_636;
wire  [1:0]  u5_col_out_637;
wire  [1:0]  u5_col_out_638;
wire  [1:0]  u5_col_out_639;
wire  [1:0]  u5_col_out_640;
wire  [1:0]  u5_col_out_641;
wire  [1:0]  u5_col_out_642;
wire  [1:0]  u5_col_out_643;
wire  [1:0]  u5_col_out_644;
wire  [1:0]  u5_col_out_645;
wire  [1:0]  u5_col_out_646;
wire  [1:0]  u5_col_out_647;
wire  [1:0]  u5_col_out_648;
wire  [1:0]  u5_col_out_649;
wire  [1:0]  u5_col_out_650;
wire  [1:0]  u5_col_out_651;
wire  [1:0]  u5_col_out_652;
wire  [1:0]  u5_col_out_653;
wire  [1:0]  u5_col_out_654;
wire  [1:0]  u5_col_out_655;
wire  [1:0]  u5_col_out_656;
wire  [1:0]  u5_col_out_657;
wire  [1:0]  u5_col_out_658;
wire  [1:0]  u5_col_out_659;
wire  [1:0]  u5_col_out_660;
wire  [1:0]  u5_col_out_661;
wire  [1:0]  u5_col_out_662;
wire  [1:0]  u5_col_out_663;
wire  [1:0]  u5_col_out_664;
wire  [1:0]  u5_col_out_665;
wire  [1:0]  u5_col_out_666;
wire  [1:0]  u5_col_out_667;
wire  [1:0]  u5_col_out_668;
wire  [1:0]  u5_col_out_669;
wire  [1:0]  u5_col_out_670;
wire  [1:0]  u5_col_out_671;
wire  [1:0]  u5_col_out_672;
wire  [1:0]  u5_col_out_673;
wire  [1:0]  u5_col_out_674;
wire  [1:0]  u5_col_out_675;
wire  [1:0]  u5_col_out_676;
wire  [1:0]  u5_col_out_677;
wire  [1:0]  u5_col_out_678;
wire  [1:0]  u5_col_out_679;
wire  [1:0]  u5_col_out_680;
wire  [1:0]  u5_col_out_681;
wire  [1:0]  u5_col_out_682;
wire  [1:0]  u5_col_out_683;
wire  [1:0]  u5_col_out_684;
wire  [1:0]  u5_col_out_685;
wire  [1:0]  u5_col_out_686;
wire  [1:0]  u5_col_out_687;
wire  [1:0]  u5_col_out_688;
wire  [1:0]  u5_col_out_689;
wire  [1:0]  u5_col_out_690;
wire  [1:0]  u5_col_out_691;
wire  [1:0]  u5_col_out_692;
wire  [1:0]  u5_col_out_693;
wire  [1:0]  u5_col_out_694;
wire  [1:0]  u5_col_out_695;
wire  [1:0]  u5_col_out_696;
wire  [1:0]  u5_col_out_697;
wire  [1:0]  u5_col_out_698;
wire  [1:0]  u5_col_out_699;
wire  [1:0]  u5_col_out_700;
wire  [1:0]  u5_col_out_701;
wire  [1:0]  u5_col_out_702;
wire  [1:0]  u5_col_out_703;
wire  [1:0]  u5_col_out_704;
wire  [1:0]  u5_col_out_705;
wire  [1:0]  u5_col_out_706;
wire  [1:0]  u5_col_out_707;
wire  [1:0]  u5_col_out_708;
wire  [1:0]  u5_col_out_709;
wire  [1:0]  u5_col_out_710;
wire  [1:0]  u5_col_out_711;
wire  [1:0]  u5_col_out_712;
wire  [1:0]  u5_col_out_713;
wire  [1:0]  u5_col_out_714;
wire  [1:0]  u5_col_out_715;
wire  [1:0]  u5_col_out_716;
wire  [1:0]  u5_col_out_717;
wire  [1:0]  u5_col_out_718;
wire  [1:0]  u5_col_out_719;
wire  [1:0]  u5_col_out_720;
wire  [1:0]  u5_col_out_721;
wire  [1:0]  u5_col_out_722;
wire  [1:0]  u5_col_out_723;
wire  [1:0]  u5_col_out_724;
wire  [1:0]  u5_col_out_725;
wire  [1:0]  u5_col_out_726;
wire  [1:0]  u5_col_out_727;
wire  [1:0]  u5_col_out_728;
wire  [1:0]  u5_col_out_729;
wire  [1:0]  u5_col_out_730;
wire  [1:0]  u5_col_out_731;
wire  [1:0]  u5_col_out_732;
wire  [1:0]  u5_col_out_733;
wire  [1:0]  u5_col_out_734;
wire  [1:0]  u5_col_out_735;
wire  [1:0]  u5_col_out_736;
wire  [1:0]  u5_col_out_737;
wire  [1:0]  u5_col_out_738;
wire  [1:0]  u5_col_out_739;
wire  [1:0]  u5_col_out_740;
wire  [1:0]  u5_col_out_741;
wire  [1:0]  u5_col_out_742;
wire  [1:0]  u5_col_out_743;
wire  [1:0]  u5_col_out_744;
wire  [1:0]  u5_col_out_745;
wire  [1:0]  u5_col_out_746;
wire  [1:0]  u5_col_out_747;
wire  [1:0]  u5_col_out_748;
wire  [1:0]  u5_col_out_749;
wire  [1:0]  u5_col_out_750;
wire  [1:0]  u5_col_out_751;
wire  [1:0]  u5_col_out_752;
wire  [1:0]  u5_col_out_753;
wire  [1:0]  u5_col_out_754;
wire  [1:0]  u5_col_out_755;
wire  [1:0]  u5_col_out_756;
wire  [1:0]  u5_col_out_757;
wire  [1:0]  u5_col_out_758;
wire  [1:0]  u5_col_out_759;
wire  [1:0]  u5_col_out_760;
wire  [1:0]  u5_col_out_761;
wire  [1:0]  u5_col_out_762;
wire  [1:0]  u5_col_out_763;
wire  [1:0]  u5_col_out_764;
wire  [1:0]  u5_col_out_765;
wire  [1:0]  u5_col_out_766;
wire  [1:0]  u5_col_out_767;
wire  [1:0]  u5_col_out_768;
wire  [1:0]  u5_col_out_769;
wire  [1:0]  u5_col_out_770;
wire  [1:0]  u5_col_out_771;
wire  [1:0]  u5_col_out_772;
wire  [1:0]  u5_col_out_773;
wire  [1:0]  u5_col_out_774;
wire  [1:0]  u5_col_out_775;
wire  [1:0]  u5_col_out_776;
wire  [1:0]  u5_col_out_777;
wire  [1:0]  u5_col_out_778;
wire  [1:0]  u5_col_out_779;
wire  [1:0]  u5_col_out_780;
wire  [1:0]  u5_col_out_781;
wire  [1:0]  u5_col_out_782;
wire  [1:0]  u5_col_out_783;
wire  [1:0]  u5_col_out_784;
wire  [1:0]  u5_col_out_785;
wire  [1:0]  u5_col_out_786;
wire  [1:0]  u5_col_out_787;
wire  [1:0]  u5_col_out_788;
wire  [1:0]  u5_col_out_789;
wire  [1:0]  u5_col_out_790;
wire  [1:0]  u5_col_out_791;
wire  [1:0]  u5_col_out_792;
wire  [1:0]  u5_col_out_793;
wire  [1:0]  u5_col_out_794;
wire  [1:0]  u5_col_out_795;
wire  [1:0]  u5_col_out_796;
wire  [1:0]  u5_col_out_797;
wire  [1:0]  u5_col_out_798;
wire  [1:0]  u5_col_out_799;
wire  [1:0]  u5_col_out_800;
wire  [1:0]  u5_col_out_801;
wire  [1:0]  u5_col_out_802;
wire  [1:0]  u5_col_out_803;
wire  [1:0]  u5_col_out_804;
wire  [1:0]  u5_col_out_805;
wire  [1:0]  u5_col_out_806;
wire  [1:0]  u5_col_out_807;
wire  [1:0]  u5_col_out_808;
wire  [1:0]  u5_col_out_809;
wire  [1:0]  u5_col_out_810;
wire  [1:0]  u5_col_out_811;
wire  [1:0]  u5_col_out_812;
wire  [1:0]  u5_col_out_813;
wire  [1:0]  u5_col_out_814;
wire  [1:0]  u5_col_out_815;
wire  [1:0]  u5_col_out_816;
wire  [1:0]  u5_col_out_817;
wire  [1:0]  u5_col_out_818;
wire  [1:0]  u5_col_out_819;
wire  [1:0]  u5_col_out_820;
wire  [1:0]  u5_col_out_821;
wire  [1:0]  u5_col_out_822;
wire  [1:0]  u5_col_out_823;
wire  [1:0]  u5_col_out_824;
wire  [1:0]  u5_col_out_825;
wire  [1:0]  u5_col_out_826;
wire  [1:0]  u5_col_out_827;
wire  [1:0]  u5_col_out_828;
wire  [1:0]  u5_col_out_829;
wire  [1:0]  u5_col_out_830;
wire  [1:0]  u5_col_out_831;
wire  [1:0]  u5_col_out_832;
wire  [1:0]  u5_col_out_833;
wire  [1:0]  u5_col_out_834;
wire  [1:0]  u5_col_out_835;
wire  [1:0]  u5_col_out_836;
wire  [1:0]  u5_col_out_837;
wire  [1:0]  u5_col_out_838;
wire  [1:0]  u5_col_out_839;
wire  [1:0]  u5_col_out_840;
wire  [1:0]  u5_col_out_841;
wire  [1:0]  u5_col_out_842;
wire  [1:0]  u5_col_out_843;
wire  [1:0]  u5_col_out_844;
wire  [1:0]  u5_col_out_845;
wire  [1:0]  u5_col_out_846;
wire  [1:0]  u5_col_out_847;
wire  [1:0]  u5_col_out_848;
wire  [1:0]  u5_col_out_849;
wire  [1:0]  u5_col_out_850;
wire  [1:0]  u5_col_out_851;
wire  [1:0]  u5_col_out_852;
wire  [1:0]  u5_col_out_853;
wire  [1:0]  u5_col_out_854;
wire  [1:0]  u5_col_out_855;
wire  [1:0]  u5_col_out_856;
wire  [1:0]  u5_col_out_857;
wire  [1:0]  u5_col_out_858;
wire  [1:0]  u5_col_out_859;
wire  [1:0]  u5_col_out_860;
wire  [1:0]  u5_col_out_861;
wire  [1:0]  u5_col_out_862;
wire  [1:0]  u5_col_out_863;
wire  [1:0]  u5_col_out_864;
wire  [1:0]  u5_col_out_865;
wire  [1:0]  u5_col_out_866;
wire  [1:0]  u5_col_out_867;
wire  [1:0]  u5_col_out_868;
wire  [1:0]  u5_col_out_869;
wire  [1:0]  u5_col_out_870;
wire  [1:0]  u5_col_out_871;
wire  [1:0]  u5_col_out_872;
wire  [1:0]  u5_col_out_873;
wire  [1:0]  u5_col_out_874;
wire  [1:0]  u5_col_out_875;
wire  [1:0]  u5_col_out_876;
wire  [1:0]  u5_col_out_877;
wire  [1:0]  u5_col_out_878;
wire  [1:0]  u5_col_out_879;
wire  [1:0]  u5_col_out_880;
wire  [1:0]  u5_col_out_881;
wire  [1:0]  u5_col_out_882;
wire  [1:0]  u5_col_out_883;
wire  [1:0]  u5_col_out_884;
wire  [1:0]  u5_col_out_885;
wire  [1:0]  u5_col_out_886;
wire  [1:0]  u5_col_out_887;
wire  [1:0]  u5_col_out_888;
wire  [1:0]  u5_col_out_889;
wire  [1:0]  u5_col_out_890;
wire  [1:0]  u5_col_out_891;
wire  [1:0]  u5_col_out_892;
wire  [1:0]  u5_col_out_893;
wire  [1:0]  u5_col_out_894;
wire  [1:0]  u5_col_out_895;
wire  [1:0]  u5_col_out_896;
wire  [1:0]  u5_col_out_897;
wire  [1:0]  u5_col_out_898;
wire  [1:0]  u5_col_out_899;
wire  [1:0]  u5_col_out_900;
wire  [1:0]  u5_col_out_901;
wire  [1:0]  u5_col_out_902;
wire  [1:0]  u5_col_out_903;
wire  [1:0]  u5_col_out_904;
wire  [1:0]  u5_col_out_905;
wire  [1:0]  u5_col_out_906;
wire  [1:0]  u5_col_out_907;
wire  [1:0]  u5_col_out_908;
wire  [1:0]  u5_col_out_909;
wire  [1:0]  u5_col_out_910;
wire  [1:0]  u5_col_out_911;
wire  [1:0]  u5_col_out_912;
wire  [1:0]  u5_col_out_913;
wire  [1:0]  u5_col_out_914;
wire  [1:0]  u5_col_out_915;
wire  [1:0]  u5_col_out_916;
wire  [1:0]  u5_col_out_917;
wire  [1:0]  u5_col_out_918;
wire  [1:0]  u5_col_out_919;
wire  [1:0]  u5_col_out_920;
wire  [1:0]  u5_col_out_921;
wire  [1:0]  u5_col_out_922;
wire  [1:0]  u5_col_out_923;
wire  [1:0]  u5_col_out_924;
wire  [1:0]  u5_col_out_925;
wire  [1:0]  u5_col_out_926;
wire  [1:0]  u5_col_out_927;
wire  [1:0]  u5_col_out_928;
wire  [1:0]  u5_col_out_929;
wire  [1:0]  u5_col_out_930;
wire  [1:0]  u5_col_out_931;
wire  [1:0]  u5_col_out_932;
wire  [1:0]  u5_col_out_933;
wire  [1:0]  u5_col_out_934;
wire  [1:0]  u5_col_out_935;
wire  [1:0]  u5_col_out_936;
wire  [1:0]  u5_col_out_937;
wire  [1:0]  u5_col_out_938;
wire  [1:0]  u5_col_out_939;
wire  [1:0]  u5_col_out_940;
wire  [1:0]  u5_col_out_941;
wire  [1:0]  u5_col_out_942;
wire  [1:0]  u5_col_out_943;
wire  [1:0]  u5_col_out_944;
wire  [1:0]  u5_col_out_945;
wire  [1:0]  u5_col_out_946;
wire  [1:0]  u5_col_out_947;
wire  [1:0]  u5_col_out_948;
wire  [1:0]  u5_col_out_949;
wire  [1:0]  u5_col_out_950;
wire  [1:0]  u5_col_out_951;
wire  [1:0]  u5_col_out_952;
wire  [1:0]  u5_col_out_953;
wire  [1:0]  u5_col_out_954;
wire  [1:0]  u5_col_out_955;
wire  [1:0]  u5_col_out_956;
wire  [1:0]  u5_col_out_957;
wire  [1:0]  u5_col_out_958;
wire  [1:0]  u5_col_out_959;
wire  [1:0]  u5_col_out_960;
wire  [1:0]  u5_col_out_961;
wire  [1:0]  u5_col_out_962;
wire  [1:0]  u5_col_out_963;
wire  [1:0]  u5_col_out_964;
wire  [1:0]  u5_col_out_965;
wire  [1:0]  u5_col_out_966;
wire  [1:0]  u5_col_out_967;
wire  [1:0]  u5_col_out_968;
wire  [1:0]  u5_col_out_969;
wire  [1:0]  u5_col_out_970;
wire  [1:0]  u5_col_out_971;
wire  [1:0]  u5_col_out_972;
wire  [1:0]  u5_col_out_973;
wire  [1:0]  u5_col_out_974;
wire  [1:0]  u5_col_out_975;
wire  [1:0]  u5_col_out_976;
wire  [1:0]  u5_col_out_977;
wire  [1:0]  u5_col_out_978;
wire  [1:0]  u5_col_out_979;
wire  [1:0]  u5_col_out_980;
wire  [1:0]  u5_col_out_981;
wire  [1:0]  u5_col_out_982;
wire  [1:0]  u5_col_out_983;
wire  [1:0]  u5_col_out_984;
wire  [1:0]  u5_col_out_985;
wire  [1:0]  u5_col_out_986;
wire  [1:0]  u5_col_out_987;
wire  [1:0]  u5_col_out_988;
wire  [1:0]  u5_col_out_989;
wire  [1:0]  u5_col_out_990;
wire  [1:0]  u5_col_out_991;
wire  [1:0]  u5_col_out_992;
wire  [1:0]  u5_col_out_993;
wire  [1:0]  u5_col_out_994;
wire  [1:0]  u5_col_out_995;
wire  [1:0]  u5_col_out_996;
wire  [1:0]  u5_col_out_997;
wire  [1:0]  u5_col_out_998;
wire  [1:0]  u5_col_out_999;
wire  [1:0]  u5_col_out_1000;
wire  [1:0]  u5_col_out_1001;
wire  [1:0]  u5_col_out_1002;
wire  [1:0]  u5_col_out_1003;
wire  [1:0]  u5_col_out_1004;
wire  [1:0]  u5_col_out_1005;
wire  [1:0]  u5_col_out_1006;
wire  [1:0]  u5_col_out_1007;
wire  [1:0]  u5_col_out_1008;
wire  [1:0]  u5_col_out_1009;
wire  [1:0]  u5_col_out_1010;
wire  [1:0]  u5_col_out_1011;
wire  [1:0]  u5_col_out_1012;
wire  [1:0]  u5_col_out_1013;
wire  [1:0]  u5_col_out_1014;
wire  [1:0]  u5_col_out_1015;
wire  [1:0]  u5_col_out_1016;
wire  [1:0]  u5_col_out_1017;
wire  [1:0]  u5_col_out_1018;
wire  [1:0]  u5_col_out_1019;
wire  [1:0]  u5_col_out_1020;
wire  [1:0]  u5_col_out_1021;
wire  [1:0]  u5_col_out_1022;
wire  [1:0]  u5_col_out_1023;
wire  [1:0]  u5_col_out_1024;
wire  [1:0]  u5_col_out_1025;
wire  [1:0]  u5_col_out_1026;
wire  [1:0]  u5_col_out_1027;
wire  [1:0]  u5_col_out_1028;
wire  [1:0]  u5_col_out_1029;
wire  [1:0]  u5_col_out_1030;
wire  [1:0]  u5_col_out_1031;
wire  [1:0]  u5_col_out_1032;
wire  [1:0]  u5_col_out_1033;

compressor_array_3_2_1033  u5_compressor_array_3_2_1033 (
    .col_in_0                ( u4_col_out_0       ),
    .col_in_1                ( u4_col_out_1       ),
    .col_in_2                ( u4_col_out_2       ),
    .col_in_3                ( u4_col_out_3       ),
    .col_in_4                ( u4_col_out_4       ),
    .col_in_5                ( u4_col_out_5       ),
    .col_in_6                ( u4_col_out_6       ),
    .col_in_7                ( u4_col_out_7       ),
    .col_in_8                ( u4_col_out_8       ),
    .col_in_9                ( u4_col_out_9       ),
    .col_in_10               ( u4_col_out_10      ),
    .col_in_11               ( u4_col_out_11      ),
    .col_in_12               ( u4_col_out_12      ),
    .col_in_13               ( u4_col_out_13      ),
    .col_in_14               ( u4_col_out_14      ),
    .col_in_15               ( u4_col_out_15      ),
    .col_in_16               ( u4_col_out_16      ),
    .col_in_17               ( u4_col_out_17      ),
    .col_in_18               ( u4_col_out_18      ),
    .col_in_19               ( u4_col_out_19      ),
    .col_in_20               ( u4_col_out_20      ),
    .col_in_21               ( u4_col_out_21      ),
    .col_in_22               ( u4_col_out_22      ),
    .col_in_23               ( u4_col_out_23      ),
    .col_in_24               ( u4_col_out_24      ),
    .col_in_25               ( u4_col_out_25      ),
    .col_in_26               ( u4_col_out_26      ),
    .col_in_27               ( u4_col_out_27      ),
    .col_in_28               ( u4_col_out_28      ),
    .col_in_29               ( u4_col_out_29      ),
    .col_in_30               ( u4_col_out_30      ),
    .col_in_31               ( u4_col_out_31      ),
    .col_in_32               ( u4_col_out_32      ),
    .col_in_33               ( u4_col_out_33      ),
    .col_in_34               ( u4_col_out_34      ),
    .col_in_35               ( u4_col_out_35      ),
    .col_in_36               ( u4_col_out_36      ),
    .col_in_37               ( u4_col_out_37      ),
    .col_in_38               ( u4_col_out_38      ),
    .col_in_39               ( u4_col_out_39      ),
    .col_in_40               ( u4_col_out_40      ),
    .col_in_41               ( u4_col_out_41      ),
    .col_in_42               ( u4_col_out_42      ),
    .col_in_43               ( u4_col_out_43      ),
    .col_in_44               ( u4_col_out_44      ),
    .col_in_45               ( u4_col_out_45      ),
    .col_in_46               ( u4_col_out_46      ),
    .col_in_47               ( u4_col_out_47      ),
    .col_in_48               ( u4_col_out_48      ),
    .col_in_49               ( u4_col_out_49      ),
    .col_in_50               ( u4_col_out_50      ),
    .col_in_51               ( u4_col_out_51      ),
    .col_in_52               ( u4_col_out_52      ),
    .col_in_53               ( u4_col_out_53      ),
    .col_in_54               ( u4_col_out_54      ),
    .col_in_55               ( u4_col_out_55      ),
    .col_in_56               ( u4_col_out_56      ),
    .col_in_57               ( u4_col_out_57      ),
    .col_in_58               ( u4_col_out_58      ),
    .col_in_59               ( u4_col_out_59      ),
    .col_in_60               ( u4_col_out_60      ),
    .col_in_61               ( u4_col_out_61      ),
    .col_in_62               ( u4_col_out_62      ),
    .col_in_63               ( u4_col_out_63      ),
    .col_in_64               ( u4_col_out_64      ),
    .col_in_65               ( u4_col_out_65      ),
    .col_in_66               ( u4_col_out_66      ),
    .col_in_67               ( u4_col_out_67      ),
    .col_in_68               ( u4_col_out_68      ),
    .col_in_69               ( u4_col_out_69      ),
    .col_in_70               ( u4_col_out_70      ),
    .col_in_71               ( u4_col_out_71      ),
    .col_in_72               ( u4_col_out_72      ),
    .col_in_73               ( u4_col_out_73      ),
    .col_in_74               ( u4_col_out_74      ),
    .col_in_75               ( u4_col_out_75      ),
    .col_in_76               ( u4_col_out_76      ),
    .col_in_77               ( u4_col_out_77      ),
    .col_in_78               ( u4_col_out_78      ),
    .col_in_79               ( u4_col_out_79      ),
    .col_in_80               ( u4_col_out_80      ),
    .col_in_81               ( u4_col_out_81      ),
    .col_in_82               ( u4_col_out_82      ),
    .col_in_83               ( u4_col_out_83      ),
    .col_in_84               ( u4_col_out_84      ),
    .col_in_85               ( u4_col_out_85      ),
    .col_in_86               ( u4_col_out_86      ),
    .col_in_87               ( u4_col_out_87      ),
    .col_in_88               ( u4_col_out_88      ),
    .col_in_89               ( u4_col_out_89      ),
    .col_in_90               ( u4_col_out_90      ),
    .col_in_91               ( u4_col_out_91      ),
    .col_in_92               ( u4_col_out_92      ),
    .col_in_93               ( u4_col_out_93      ),
    .col_in_94               ( u4_col_out_94      ),
    .col_in_95               ( u4_col_out_95      ),
    .col_in_96               ( u4_col_out_96      ),
    .col_in_97               ( u4_col_out_97      ),
    .col_in_98               ( u4_col_out_98      ),
    .col_in_99               ( u4_col_out_99      ),
    .col_in_100              ( u4_col_out_100     ),
    .col_in_101              ( u4_col_out_101     ),
    .col_in_102              ( u4_col_out_102     ),
    .col_in_103              ( u4_col_out_103     ),
    .col_in_104              ( u4_col_out_104     ),
    .col_in_105              ( u4_col_out_105     ),
    .col_in_106              ( u4_col_out_106     ),
    .col_in_107              ( u4_col_out_107     ),
    .col_in_108              ( u4_col_out_108     ),
    .col_in_109              ( u4_col_out_109     ),
    .col_in_110              ( u4_col_out_110     ),
    .col_in_111              ( u4_col_out_111     ),
    .col_in_112              ( u4_col_out_112     ),
    .col_in_113              ( u4_col_out_113     ),
    .col_in_114              ( u4_col_out_114     ),
    .col_in_115              ( u4_col_out_115     ),
    .col_in_116              ( u4_col_out_116     ),
    .col_in_117              ( u4_col_out_117     ),
    .col_in_118              ( u4_col_out_118     ),
    .col_in_119              ( u4_col_out_119     ),
    .col_in_120              ( u4_col_out_120     ),
    .col_in_121              ( u4_col_out_121     ),
    .col_in_122              ( u4_col_out_122     ),
    .col_in_123              ( u4_col_out_123     ),
    .col_in_124              ( u4_col_out_124     ),
    .col_in_125              ( u4_col_out_125     ),
    .col_in_126              ( u4_col_out_126     ),
    .col_in_127              ( u4_col_out_127     ),
    .col_in_128              ( u4_col_out_128     ),
    .col_in_129              ( u4_col_out_129     ),
    .col_in_130              ( u4_col_out_130     ),
    .col_in_131              ( u4_col_out_131     ),
    .col_in_132              ( u4_col_out_132     ),
    .col_in_133              ( u4_col_out_133     ),
    .col_in_134              ( u4_col_out_134     ),
    .col_in_135              ( u4_col_out_135     ),
    .col_in_136              ( u4_col_out_136     ),
    .col_in_137              ( u4_col_out_137     ),
    .col_in_138              ( u4_col_out_138     ),
    .col_in_139              ( u4_col_out_139     ),
    .col_in_140              ( u4_col_out_140     ),
    .col_in_141              ( u4_col_out_141     ),
    .col_in_142              ( u4_col_out_142     ),
    .col_in_143              ( u4_col_out_143     ),
    .col_in_144              ( u4_col_out_144     ),
    .col_in_145              ( u4_col_out_145     ),
    .col_in_146              ( u4_col_out_146     ),
    .col_in_147              ( u4_col_out_147     ),
    .col_in_148              ( u4_col_out_148     ),
    .col_in_149              ( u4_col_out_149     ),
    .col_in_150              ( u4_col_out_150     ),
    .col_in_151              ( u4_col_out_151     ),
    .col_in_152              ( u4_col_out_152     ),
    .col_in_153              ( u4_col_out_153     ),
    .col_in_154              ( u4_col_out_154     ),
    .col_in_155              ( u4_col_out_155     ),
    .col_in_156              ( u4_col_out_156     ),
    .col_in_157              ( u4_col_out_157     ),
    .col_in_158              ( u4_col_out_158     ),
    .col_in_159              ( u4_col_out_159     ),
    .col_in_160              ( u4_col_out_160     ),
    .col_in_161              ( u4_col_out_161     ),
    .col_in_162              ( u4_col_out_162     ),
    .col_in_163              ( u4_col_out_163     ),
    .col_in_164              ( u4_col_out_164     ),
    .col_in_165              ( u4_col_out_165     ),
    .col_in_166              ( u4_col_out_166     ),
    .col_in_167              ( u4_col_out_167     ),
    .col_in_168              ( u4_col_out_168     ),
    .col_in_169              ( u4_col_out_169     ),
    .col_in_170              ( u4_col_out_170     ),
    .col_in_171              ( u4_col_out_171     ),
    .col_in_172              ( u4_col_out_172     ),
    .col_in_173              ( u4_col_out_173     ),
    .col_in_174              ( u4_col_out_174     ),
    .col_in_175              ( u4_col_out_175     ),
    .col_in_176              ( u4_col_out_176     ),
    .col_in_177              ( u4_col_out_177     ),
    .col_in_178              ( u4_col_out_178     ),
    .col_in_179              ( u4_col_out_179     ),
    .col_in_180              ( u4_col_out_180     ),
    .col_in_181              ( u4_col_out_181     ),
    .col_in_182              ( u4_col_out_182     ),
    .col_in_183              ( u4_col_out_183     ),
    .col_in_184              ( u4_col_out_184     ),
    .col_in_185              ( u4_col_out_185     ),
    .col_in_186              ( u4_col_out_186     ),
    .col_in_187              ( u4_col_out_187     ),
    .col_in_188              ( u4_col_out_188     ),
    .col_in_189              ( u4_col_out_189     ),
    .col_in_190              ( u4_col_out_190     ),
    .col_in_191              ( u4_col_out_191     ),
    .col_in_192              ( u4_col_out_192     ),
    .col_in_193              ( u4_col_out_193     ),
    .col_in_194              ( u4_col_out_194     ),
    .col_in_195              ( u4_col_out_195     ),
    .col_in_196              ( u4_col_out_196     ),
    .col_in_197              ( u4_col_out_197     ),
    .col_in_198              ( u4_col_out_198     ),
    .col_in_199              ( u4_col_out_199     ),
    .col_in_200              ( u4_col_out_200     ),
    .col_in_201              ( u4_col_out_201     ),
    .col_in_202              ( u4_col_out_202     ),
    .col_in_203              ( u4_col_out_203     ),
    .col_in_204              ( u4_col_out_204     ),
    .col_in_205              ( u4_col_out_205     ),
    .col_in_206              ( u4_col_out_206     ),
    .col_in_207              ( u4_col_out_207     ),
    .col_in_208              ( u4_col_out_208     ),
    .col_in_209              ( u4_col_out_209     ),
    .col_in_210              ( u4_col_out_210     ),
    .col_in_211              ( u4_col_out_211     ),
    .col_in_212              ( u4_col_out_212     ),
    .col_in_213              ( u4_col_out_213     ),
    .col_in_214              ( u4_col_out_214     ),
    .col_in_215              ( u4_col_out_215     ),
    .col_in_216              ( u4_col_out_216     ),
    .col_in_217              ( u4_col_out_217     ),
    .col_in_218              ( u4_col_out_218     ),
    .col_in_219              ( u4_col_out_219     ),
    .col_in_220              ( u4_col_out_220     ),
    .col_in_221              ( u4_col_out_221     ),
    .col_in_222              ( u4_col_out_222     ),
    .col_in_223              ( u4_col_out_223     ),
    .col_in_224              ( u4_col_out_224     ),
    .col_in_225              ( u4_col_out_225     ),
    .col_in_226              ( u4_col_out_226     ),
    .col_in_227              ( u4_col_out_227     ),
    .col_in_228              ( u4_col_out_228     ),
    .col_in_229              ( u4_col_out_229     ),
    .col_in_230              ( u4_col_out_230     ),
    .col_in_231              ( u4_col_out_231     ),
    .col_in_232              ( u4_col_out_232     ),
    .col_in_233              ( u4_col_out_233     ),
    .col_in_234              ( u4_col_out_234     ),
    .col_in_235              ( u4_col_out_235     ),
    .col_in_236              ( u4_col_out_236     ),
    .col_in_237              ( u4_col_out_237     ),
    .col_in_238              ( u4_col_out_238     ),
    .col_in_239              ( u4_col_out_239     ),
    .col_in_240              ( u4_col_out_240     ),
    .col_in_241              ( u4_col_out_241     ),
    .col_in_242              ( u4_col_out_242     ),
    .col_in_243              ( u4_col_out_243     ),
    .col_in_244              ( u4_col_out_244     ),
    .col_in_245              ( u4_col_out_245     ),
    .col_in_246              ( u4_col_out_246     ),
    .col_in_247              ( u4_col_out_247     ),
    .col_in_248              ( u4_col_out_248     ),
    .col_in_249              ( u4_col_out_249     ),
    .col_in_250              ( u4_col_out_250     ),
    .col_in_251              ( u4_col_out_251     ),
    .col_in_252              ( u4_col_out_252     ),
    .col_in_253              ( u4_col_out_253     ),
    .col_in_254              ( u4_col_out_254     ),
    .col_in_255              ( u4_col_out_255     ),
    .col_in_256              ( u4_col_out_256     ),
    .col_in_257              ( u4_col_out_257     ),
    .col_in_258              ( u4_col_out_258     ),
    .col_in_259              ( u4_col_out_259     ),
    .col_in_260              ( u4_col_out_260     ),
    .col_in_261              ( u4_col_out_261     ),
    .col_in_262              ( u4_col_out_262     ),
    .col_in_263              ( u4_col_out_263     ),
    .col_in_264              ( u4_col_out_264     ),
    .col_in_265              ( u4_col_out_265     ),
    .col_in_266              ( u4_col_out_266     ),
    .col_in_267              ( u4_col_out_267     ),
    .col_in_268              ( u4_col_out_268     ),
    .col_in_269              ( u4_col_out_269     ),
    .col_in_270              ( u4_col_out_270     ),
    .col_in_271              ( u4_col_out_271     ),
    .col_in_272              ( u4_col_out_272     ),
    .col_in_273              ( u4_col_out_273     ),
    .col_in_274              ( u4_col_out_274     ),
    .col_in_275              ( u4_col_out_275     ),
    .col_in_276              ( u4_col_out_276     ),
    .col_in_277              ( u4_col_out_277     ),
    .col_in_278              ( u4_col_out_278     ),
    .col_in_279              ( u4_col_out_279     ),
    .col_in_280              ( u4_col_out_280     ),
    .col_in_281              ( u4_col_out_281     ),
    .col_in_282              ( u4_col_out_282     ),
    .col_in_283              ( u4_col_out_283     ),
    .col_in_284              ( u4_col_out_284     ),
    .col_in_285              ( u4_col_out_285     ),
    .col_in_286              ( u4_col_out_286     ),
    .col_in_287              ( u4_col_out_287     ),
    .col_in_288              ( u4_col_out_288     ),
    .col_in_289              ( u4_col_out_289     ),
    .col_in_290              ( u4_col_out_290     ),
    .col_in_291              ( u4_col_out_291     ),
    .col_in_292              ( u4_col_out_292     ),
    .col_in_293              ( u4_col_out_293     ),
    .col_in_294              ( u4_col_out_294     ),
    .col_in_295              ( u4_col_out_295     ),
    .col_in_296              ( u4_col_out_296     ),
    .col_in_297              ( u4_col_out_297     ),
    .col_in_298              ( u4_col_out_298     ),
    .col_in_299              ( u4_col_out_299     ),
    .col_in_300              ( u4_col_out_300     ),
    .col_in_301              ( u4_col_out_301     ),
    .col_in_302              ( u4_col_out_302     ),
    .col_in_303              ( u4_col_out_303     ),
    .col_in_304              ( u4_col_out_304     ),
    .col_in_305              ( u4_col_out_305     ),
    .col_in_306              ( u4_col_out_306     ),
    .col_in_307              ( u4_col_out_307     ),
    .col_in_308              ( u4_col_out_308     ),
    .col_in_309              ( u4_col_out_309     ),
    .col_in_310              ( u4_col_out_310     ),
    .col_in_311              ( u4_col_out_311     ),
    .col_in_312              ( u4_col_out_312     ),
    .col_in_313              ( u4_col_out_313     ),
    .col_in_314              ( u4_col_out_314     ),
    .col_in_315              ( u4_col_out_315     ),
    .col_in_316              ( u4_col_out_316     ),
    .col_in_317              ( u4_col_out_317     ),
    .col_in_318              ( u4_col_out_318     ),
    .col_in_319              ( u4_col_out_319     ),
    .col_in_320              ( u4_col_out_320     ),
    .col_in_321              ( u4_col_out_321     ),
    .col_in_322              ( u4_col_out_322     ),
    .col_in_323              ( u4_col_out_323     ),
    .col_in_324              ( u4_col_out_324     ),
    .col_in_325              ( u4_col_out_325     ),
    .col_in_326              ( u4_col_out_326     ),
    .col_in_327              ( u4_col_out_327     ),
    .col_in_328              ( u4_col_out_328     ),
    .col_in_329              ( u4_col_out_329     ),
    .col_in_330              ( u4_col_out_330     ),
    .col_in_331              ( u4_col_out_331     ),
    .col_in_332              ( u4_col_out_332     ),
    .col_in_333              ( u4_col_out_333     ),
    .col_in_334              ( u4_col_out_334     ),
    .col_in_335              ( u4_col_out_335     ),
    .col_in_336              ( u4_col_out_336     ),
    .col_in_337              ( u4_col_out_337     ),
    .col_in_338              ( u4_col_out_338     ),
    .col_in_339              ( u4_col_out_339     ),
    .col_in_340              ( u4_col_out_340     ),
    .col_in_341              ( u4_col_out_341     ),
    .col_in_342              ( u4_col_out_342     ),
    .col_in_343              ( u4_col_out_343     ),
    .col_in_344              ( u4_col_out_344     ),
    .col_in_345              ( u4_col_out_345     ),
    .col_in_346              ( u4_col_out_346     ),
    .col_in_347              ( u4_col_out_347     ),
    .col_in_348              ( u4_col_out_348     ),
    .col_in_349              ( u4_col_out_349     ),
    .col_in_350              ( u4_col_out_350     ),
    .col_in_351              ( u4_col_out_351     ),
    .col_in_352              ( u4_col_out_352     ),
    .col_in_353              ( u4_col_out_353     ),
    .col_in_354              ( u4_col_out_354     ),
    .col_in_355              ( u4_col_out_355     ),
    .col_in_356              ( u4_col_out_356     ),
    .col_in_357              ( u4_col_out_357     ),
    .col_in_358              ( u4_col_out_358     ),
    .col_in_359              ( u4_col_out_359     ),
    .col_in_360              ( u4_col_out_360     ),
    .col_in_361              ( u4_col_out_361     ),
    .col_in_362              ( u4_col_out_362     ),
    .col_in_363              ( u4_col_out_363     ),
    .col_in_364              ( u4_col_out_364     ),
    .col_in_365              ( u4_col_out_365     ),
    .col_in_366              ( u4_col_out_366     ),
    .col_in_367              ( u4_col_out_367     ),
    .col_in_368              ( u4_col_out_368     ),
    .col_in_369              ( u4_col_out_369     ),
    .col_in_370              ( u4_col_out_370     ),
    .col_in_371              ( u4_col_out_371     ),
    .col_in_372              ( u4_col_out_372     ),
    .col_in_373              ( u4_col_out_373     ),
    .col_in_374              ( u4_col_out_374     ),
    .col_in_375              ( u4_col_out_375     ),
    .col_in_376              ( u4_col_out_376     ),
    .col_in_377              ( u4_col_out_377     ),
    .col_in_378              ( u4_col_out_378     ),
    .col_in_379              ( u4_col_out_379     ),
    .col_in_380              ( u4_col_out_380     ),
    .col_in_381              ( u4_col_out_381     ),
    .col_in_382              ( u4_col_out_382     ),
    .col_in_383              ( u4_col_out_383     ),
    .col_in_384              ( u4_col_out_384     ),
    .col_in_385              ( u4_col_out_385     ),
    .col_in_386              ( u4_col_out_386     ),
    .col_in_387              ( u4_col_out_387     ),
    .col_in_388              ( u4_col_out_388     ),
    .col_in_389              ( u4_col_out_389     ),
    .col_in_390              ( u4_col_out_390     ),
    .col_in_391              ( u4_col_out_391     ),
    .col_in_392              ( u4_col_out_392     ),
    .col_in_393              ( u4_col_out_393     ),
    .col_in_394              ( u4_col_out_394     ),
    .col_in_395              ( u4_col_out_395     ),
    .col_in_396              ( u4_col_out_396     ),
    .col_in_397              ( u4_col_out_397     ),
    .col_in_398              ( u4_col_out_398     ),
    .col_in_399              ( u4_col_out_399     ),
    .col_in_400              ( u4_col_out_400     ),
    .col_in_401              ( u4_col_out_401     ),
    .col_in_402              ( u4_col_out_402     ),
    .col_in_403              ( u4_col_out_403     ),
    .col_in_404              ( u4_col_out_404     ),
    .col_in_405              ( u4_col_out_405     ),
    .col_in_406              ( u4_col_out_406     ),
    .col_in_407              ( u4_col_out_407     ),
    .col_in_408              ( u4_col_out_408     ),
    .col_in_409              ( u4_col_out_409     ),
    .col_in_410              ( u4_col_out_410     ),
    .col_in_411              ( u4_col_out_411     ),
    .col_in_412              ( u4_col_out_412     ),
    .col_in_413              ( u4_col_out_413     ),
    .col_in_414              ( u4_col_out_414     ),
    .col_in_415              ( u4_col_out_415     ),
    .col_in_416              ( u4_col_out_416     ),
    .col_in_417              ( u4_col_out_417     ),
    .col_in_418              ( u4_col_out_418     ),
    .col_in_419              ( u4_col_out_419     ),
    .col_in_420              ( u4_col_out_420     ),
    .col_in_421              ( u4_col_out_421     ),
    .col_in_422              ( u4_col_out_422     ),
    .col_in_423              ( u4_col_out_423     ),
    .col_in_424              ( u4_col_out_424     ),
    .col_in_425              ( u4_col_out_425     ),
    .col_in_426              ( u4_col_out_426     ),
    .col_in_427              ( u4_col_out_427     ),
    .col_in_428              ( u4_col_out_428     ),
    .col_in_429              ( u4_col_out_429     ),
    .col_in_430              ( u4_col_out_430     ),
    .col_in_431              ( u4_col_out_431     ),
    .col_in_432              ( u4_col_out_432     ),
    .col_in_433              ( u4_col_out_433     ),
    .col_in_434              ( u4_col_out_434     ),
    .col_in_435              ( u4_col_out_435     ),
    .col_in_436              ( u4_col_out_436     ),
    .col_in_437              ( u4_col_out_437     ),
    .col_in_438              ( u4_col_out_438     ),
    .col_in_439              ( u4_col_out_439     ),
    .col_in_440              ( u4_col_out_440     ),
    .col_in_441              ( u4_col_out_441     ),
    .col_in_442              ( u4_col_out_442     ),
    .col_in_443              ( u4_col_out_443     ),
    .col_in_444              ( u4_col_out_444     ),
    .col_in_445              ( u4_col_out_445     ),
    .col_in_446              ( u4_col_out_446     ),
    .col_in_447              ( u4_col_out_447     ),
    .col_in_448              ( u4_col_out_448     ),
    .col_in_449              ( u4_col_out_449     ),
    .col_in_450              ( u4_col_out_450     ),
    .col_in_451              ( u4_col_out_451     ),
    .col_in_452              ( u4_col_out_452     ),
    .col_in_453              ( u4_col_out_453     ),
    .col_in_454              ( u4_col_out_454     ),
    .col_in_455              ( u4_col_out_455     ),
    .col_in_456              ( u4_col_out_456     ),
    .col_in_457              ( u4_col_out_457     ),
    .col_in_458              ( u4_col_out_458     ),
    .col_in_459              ( u4_col_out_459     ),
    .col_in_460              ( u4_col_out_460     ),
    .col_in_461              ( u4_col_out_461     ),
    .col_in_462              ( u4_col_out_462     ),
    .col_in_463              ( u4_col_out_463     ),
    .col_in_464              ( u4_col_out_464     ),
    .col_in_465              ( u4_col_out_465     ),
    .col_in_466              ( u4_col_out_466     ),
    .col_in_467              ( u4_col_out_467     ),
    .col_in_468              ( u4_col_out_468     ),
    .col_in_469              ( u4_col_out_469     ),
    .col_in_470              ( u4_col_out_470     ),
    .col_in_471              ( u4_col_out_471     ),
    .col_in_472              ( u4_col_out_472     ),
    .col_in_473              ( u4_col_out_473     ),
    .col_in_474              ( u4_col_out_474     ),
    .col_in_475              ( u4_col_out_475     ),
    .col_in_476              ( u4_col_out_476     ),
    .col_in_477              ( u4_col_out_477     ),
    .col_in_478              ( u4_col_out_478     ),
    .col_in_479              ( u4_col_out_479     ),
    .col_in_480              ( u4_col_out_480     ),
    .col_in_481              ( u4_col_out_481     ),
    .col_in_482              ( u4_col_out_482     ),
    .col_in_483              ( u4_col_out_483     ),
    .col_in_484              ( u4_col_out_484     ),
    .col_in_485              ( u4_col_out_485     ),
    .col_in_486              ( u4_col_out_486     ),
    .col_in_487              ( u4_col_out_487     ),
    .col_in_488              ( u4_col_out_488     ),
    .col_in_489              ( u4_col_out_489     ),
    .col_in_490              ( u4_col_out_490     ),
    .col_in_491              ( u4_col_out_491     ),
    .col_in_492              ( u4_col_out_492     ),
    .col_in_493              ( u4_col_out_493     ),
    .col_in_494              ( u4_col_out_494     ),
    .col_in_495              ( u4_col_out_495     ),
    .col_in_496              ( u4_col_out_496     ),
    .col_in_497              ( u4_col_out_497     ),
    .col_in_498              ( u4_col_out_498     ),
    .col_in_499              ( u4_col_out_499     ),
    .col_in_500              ( u4_col_out_500     ),
    .col_in_501              ( u4_col_out_501     ),
    .col_in_502              ( u4_col_out_502     ),
    .col_in_503              ( u4_col_out_503     ),
    .col_in_504              ( u4_col_out_504     ),
    .col_in_505              ( u4_col_out_505     ),
    .col_in_506              ( u4_col_out_506     ),
    .col_in_507              ( u4_col_out_507     ),
    .col_in_508              ( u4_col_out_508     ),
    .col_in_509              ( u4_col_out_509     ),
    .col_in_510              ( u4_col_out_510     ),
    .col_in_511              ( u4_col_out_511     ),
    .col_in_512              ( u4_col_out_512     ),
    .col_in_513              ( u4_col_out_513     ),
    .col_in_514              ( u4_col_out_514     ),
    .col_in_515              ( u4_col_out_515     ),
    .col_in_516              ( u4_col_out_516     ),
    .col_in_517              ( u4_col_out_517     ),
    .col_in_518              ( u4_col_out_518     ),
    .col_in_519              ( u4_col_out_519     ),
    .col_in_520              ( u4_col_out_520     ),
    .col_in_521              ( u4_col_out_521     ),
    .col_in_522              ( u4_col_out_522     ),
    .col_in_523              ( u4_col_out_523     ),
    .col_in_524              ( u4_col_out_524     ),
    .col_in_525              ( u4_col_out_525     ),
    .col_in_526              ( u4_col_out_526     ),
    .col_in_527              ( u4_col_out_527     ),
    .col_in_528              ( u4_col_out_528     ),
    .col_in_529              ( u4_col_out_529     ),
    .col_in_530              ( u4_col_out_530     ),
    .col_in_531              ( u4_col_out_531     ),
    .col_in_532              ( u4_col_out_532     ),
    .col_in_533              ( u4_col_out_533     ),
    .col_in_534              ( u4_col_out_534     ),
    .col_in_535              ( u4_col_out_535     ),
    .col_in_536              ( u4_col_out_536     ),
    .col_in_537              ( u4_col_out_537     ),
    .col_in_538              ( u4_col_out_538     ),
    .col_in_539              ( u4_col_out_539     ),
    .col_in_540              ( u4_col_out_540     ),
    .col_in_541              ( u4_col_out_541     ),
    .col_in_542              ( u4_col_out_542     ),
    .col_in_543              ( u4_col_out_543     ),
    .col_in_544              ( u4_col_out_544     ),
    .col_in_545              ( u4_col_out_545     ),
    .col_in_546              ( u4_col_out_546     ),
    .col_in_547              ( u4_col_out_547     ),
    .col_in_548              ( u4_col_out_548     ),
    .col_in_549              ( u4_col_out_549     ),
    .col_in_550              ( u4_col_out_550     ),
    .col_in_551              ( u4_col_out_551     ),
    .col_in_552              ( u4_col_out_552     ),
    .col_in_553              ( u4_col_out_553     ),
    .col_in_554              ( u4_col_out_554     ),
    .col_in_555              ( u4_col_out_555     ),
    .col_in_556              ( u4_col_out_556     ),
    .col_in_557              ( u4_col_out_557     ),
    .col_in_558              ( u4_col_out_558     ),
    .col_in_559              ( u4_col_out_559     ),
    .col_in_560              ( u4_col_out_560     ),
    .col_in_561              ( u4_col_out_561     ),
    .col_in_562              ( u4_col_out_562     ),
    .col_in_563              ( u4_col_out_563     ),
    .col_in_564              ( u4_col_out_564     ),
    .col_in_565              ( u4_col_out_565     ),
    .col_in_566              ( u4_col_out_566     ),
    .col_in_567              ( u4_col_out_567     ),
    .col_in_568              ( u4_col_out_568     ),
    .col_in_569              ( u4_col_out_569     ),
    .col_in_570              ( u4_col_out_570     ),
    .col_in_571              ( u4_col_out_571     ),
    .col_in_572              ( u4_col_out_572     ),
    .col_in_573              ( u4_col_out_573     ),
    .col_in_574              ( u4_col_out_574     ),
    .col_in_575              ( u4_col_out_575     ),
    .col_in_576              ( u4_col_out_576     ),
    .col_in_577              ( u4_col_out_577     ),
    .col_in_578              ( u4_col_out_578     ),
    .col_in_579              ( u4_col_out_579     ),
    .col_in_580              ( u4_col_out_580     ),
    .col_in_581              ( u4_col_out_581     ),
    .col_in_582              ( u4_col_out_582     ),
    .col_in_583              ( u4_col_out_583     ),
    .col_in_584              ( u4_col_out_584     ),
    .col_in_585              ( u4_col_out_585     ),
    .col_in_586              ( u4_col_out_586     ),
    .col_in_587              ( u4_col_out_587     ),
    .col_in_588              ( u4_col_out_588     ),
    .col_in_589              ( u4_col_out_589     ),
    .col_in_590              ( u4_col_out_590     ),
    .col_in_591              ( u4_col_out_591     ),
    .col_in_592              ( u4_col_out_592     ),
    .col_in_593              ( u4_col_out_593     ),
    .col_in_594              ( u4_col_out_594     ),
    .col_in_595              ( u4_col_out_595     ),
    .col_in_596              ( u4_col_out_596     ),
    .col_in_597              ( u4_col_out_597     ),
    .col_in_598              ( u4_col_out_598     ),
    .col_in_599              ( u4_col_out_599     ),
    .col_in_600              ( u4_col_out_600     ),
    .col_in_601              ( u4_col_out_601     ),
    .col_in_602              ( u4_col_out_602     ),
    .col_in_603              ( u4_col_out_603     ),
    .col_in_604              ( u4_col_out_604     ),
    .col_in_605              ( u4_col_out_605     ),
    .col_in_606              ( u4_col_out_606     ),
    .col_in_607              ( u4_col_out_607     ),
    .col_in_608              ( u4_col_out_608     ),
    .col_in_609              ( u4_col_out_609     ),
    .col_in_610              ( u4_col_out_610     ),
    .col_in_611              ( u4_col_out_611     ),
    .col_in_612              ( u4_col_out_612     ),
    .col_in_613              ( u4_col_out_613     ),
    .col_in_614              ( u4_col_out_614     ),
    .col_in_615              ( u4_col_out_615     ),
    .col_in_616              ( u4_col_out_616     ),
    .col_in_617              ( u4_col_out_617     ),
    .col_in_618              ( u4_col_out_618     ),
    .col_in_619              ( u4_col_out_619     ),
    .col_in_620              ( u4_col_out_620     ),
    .col_in_621              ( u4_col_out_621     ),
    .col_in_622              ( u4_col_out_622     ),
    .col_in_623              ( u4_col_out_623     ),
    .col_in_624              ( u4_col_out_624     ),
    .col_in_625              ( u4_col_out_625     ),
    .col_in_626              ( u4_col_out_626     ),
    .col_in_627              ( u4_col_out_627     ),
    .col_in_628              ( u4_col_out_628     ),
    .col_in_629              ( u4_col_out_629     ),
    .col_in_630              ( u4_col_out_630     ),
    .col_in_631              ( u4_col_out_631     ),
    .col_in_632              ( u4_col_out_632     ),
    .col_in_633              ( u4_col_out_633     ),
    .col_in_634              ( u4_col_out_634     ),
    .col_in_635              ( u4_col_out_635     ),
    .col_in_636              ( u4_col_out_636     ),
    .col_in_637              ( u4_col_out_637     ),
    .col_in_638              ( u4_col_out_638     ),
    .col_in_639              ( u4_col_out_639     ),
    .col_in_640              ( u4_col_out_640     ),
    .col_in_641              ( u4_col_out_641     ),
    .col_in_642              ( u4_col_out_642     ),
    .col_in_643              ( u4_col_out_643     ),
    .col_in_644              ( u4_col_out_644     ),
    .col_in_645              ( u4_col_out_645     ),
    .col_in_646              ( u4_col_out_646     ),
    .col_in_647              ( u4_col_out_647     ),
    .col_in_648              ( u4_col_out_648     ),
    .col_in_649              ( u4_col_out_649     ),
    .col_in_650              ( u4_col_out_650     ),
    .col_in_651              ( u4_col_out_651     ),
    .col_in_652              ( u4_col_out_652     ),
    .col_in_653              ( u4_col_out_653     ),
    .col_in_654              ( u4_col_out_654     ),
    .col_in_655              ( u4_col_out_655     ),
    .col_in_656              ( u4_col_out_656     ),
    .col_in_657              ( u4_col_out_657     ),
    .col_in_658              ( u4_col_out_658     ),
    .col_in_659              ( u4_col_out_659     ),
    .col_in_660              ( u4_col_out_660     ),
    .col_in_661              ( u4_col_out_661     ),
    .col_in_662              ( u4_col_out_662     ),
    .col_in_663              ( u4_col_out_663     ),
    .col_in_664              ( u4_col_out_664     ),
    .col_in_665              ( u4_col_out_665     ),
    .col_in_666              ( u4_col_out_666     ),
    .col_in_667              ( u4_col_out_667     ),
    .col_in_668              ( u4_col_out_668     ),
    .col_in_669              ( u4_col_out_669     ),
    .col_in_670              ( u4_col_out_670     ),
    .col_in_671              ( u4_col_out_671     ),
    .col_in_672              ( u4_col_out_672     ),
    .col_in_673              ( u4_col_out_673     ),
    .col_in_674              ( u4_col_out_674     ),
    .col_in_675              ( u4_col_out_675     ),
    .col_in_676              ( u4_col_out_676     ),
    .col_in_677              ( u4_col_out_677     ),
    .col_in_678              ( u4_col_out_678     ),
    .col_in_679              ( u4_col_out_679     ),
    .col_in_680              ( u4_col_out_680     ),
    .col_in_681              ( u4_col_out_681     ),
    .col_in_682              ( u4_col_out_682     ),
    .col_in_683              ( u4_col_out_683     ),
    .col_in_684              ( u4_col_out_684     ),
    .col_in_685              ( u4_col_out_685     ),
    .col_in_686              ( u4_col_out_686     ),
    .col_in_687              ( u4_col_out_687     ),
    .col_in_688              ( u4_col_out_688     ),
    .col_in_689              ( u4_col_out_689     ),
    .col_in_690              ( u4_col_out_690     ),
    .col_in_691              ( u4_col_out_691     ),
    .col_in_692              ( u4_col_out_692     ),
    .col_in_693              ( u4_col_out_693     ),
    .col_in_694              ( u4_col_out_694     ),
    .col_in_695              ( u4_col_out_695     ),
    .col_in_696              ( u4_col_out_696     ),
    .col_in_697              ( u4_col_out_697     ),
    .col_in_698              ( u4_col_out_698     ),
    .col_in_699              ( u4_col_out_699     ),
    .col_in_700              ( u4_col_out_700     ),
    .col_in_701              ( u4_col_out_701     ),
    .col_in_702              ( u4_col_out_702     ),
    .col_in_703              ( u4_col_out_703     ),
    .col_in_704              ( u4_col_out_704     ),
    .col_in_705              ( u4_col_out_705     ),
    .col_in_706              ( u4_col_out_706     ),
    .col_in_707              ( u4_col_out_707     ),
    .col_in_708              ( u4_col_out_708     ),
    .col_in_709              ( u4_col_out_709     ),
    .col_in_710              ( u4_col_out_710     ),
    .col_in_711              ( u4_col_out_711     ),
    .col_in_712              ( u4_col_out_712     ),
    .col_in_713              ( u4_col_out_713     ),
    .col_in_714              ( u4_col_out_714     ),
    .col_in_715              ( u4_col_out_715     ),
    .col_in_716              ( u4_col_out_716     ),
    .col_in_717              ( u4_col_out_717     ),
    .col_in_718              ( u4_col_out_718     ),
    .col_in_719              ( u4_col_out_719     ),
    .col_in_720              ( u4_col_out_720     ),
    .col_in_721              ( u4_col_out_721     ),
    .col_in_722              ( u4_col_out_722     ),
    .col_in_723              ( u4_col_out_723     ),
    .col_in_724              ( u4_col_out_724     ),
    .col_in_725              ( u4_col_out_725     ),
    .col_in_726              ( u4_col_out_726     ),
    .col_in_727              ( u4_col_out_727     ),
    .col_in_728              ( u4_col_out_728     ),
    .col_in_729              ( u4_col_out_729     ),
    .col_in_730              ( u4_col_out_730     ),
    .col_in_731              ( u4_col_out_731     ),
    .col_in_732              ( u4_col_out_732     ),
    .col_in_733              ( u4_col_out_733     ),
    .col_in_734              ( u4_col_out_734     ),
    .col_in_735              ( u4_col_out_735     ),
    .col_in_736              ( u4_col_out_736     ),
    .col_in_737              ( u4_col_out_737     ),
    .col_in_738              ( u4_col_out_738     ),
    .col_in_739              ( u4_col_out_739     ),
    .col_in_740              ( u4_col_out_740     ),
    .col_in_741              ( u4_col_out_741     ),
    .col_in_742              ( u4_col_out_742     ),
    .col_in_743              ( u4_col_out_743     ),
    .col_in_744              ( u4_col_out_744     ),
    .col_in_745              ( u4_col_out_745     ),
    .col_in_746              ( u4_col_out_746     ),
    .col_in_747              ( u4_col_out_747     ),
    .col_in_748              ( u4_col_out_748     ),
    .col_in_749              ( u4_col_out_749     ),
    .col_in_750              ( u4_col_out_750     ),
    .col_in_751              ( u4_col_out_751     ),
    .col_in_752              ( u4_col_out_752     ),
    .col_in_753              ( u4_col_out_753     ),
    .col_in_754              ( u4_col_out_754     ),
    .col_in_755              ( u4_col_out_755     ),
    .col_in_756              ( u4_col_out_756     ),
    .col_in_757              ( u4_col_out_757     ),
    .col_in_758              ( u4_col_out_758     ),
    .col_in_759              ( u4_col_out_759     ),
    .col_in_760              ( u4_col_out_760     ),
    .col_in_761              ( u4_col_out_761     ),
    .col_in_762              ( u4_col_out_762     ),
    .col_in_763              ( u4_col_out_763     ),
    .col_in_764              ( u4_col_out_764     ),
    .col_in_765              ( u4_col_out_765     ),
    .col_in_766              ( u4_col_out_766     ),
    .col_in_767              ( u4_col_out_767     ),
    .col_in_768              ( u4_col_out_768     ),
    .col_in_769              ( u4_col_out_769     ),
    .col_in_770              ( u4_col_out_770     ),
    .col_in_771              ( u4_col_out_771     ),
    .col_in_772              ( u4_col_out_772     ),
    .col_in_773              ( u4_col_out_773     ),
    .col_in_774              ( u4_col_out_774     ),
    .col_in_775              ( u4_col_out_775     ),
    .col_in_776              ( u4_col_out_776     ),
    .col_in_777              ( u4_col_out_777     ),
    .col_in_778              ( u4_col_out_778     ),
    .col_in_779              ( u4_col_out_779     ),
    .col_in_780              ( u4_col_out_780     ),
    .col_in_781              ( u4_col_out_781     ),
    .col_in_782              ( u4_col_out_782     ),
    .col_in_783              ( u4_col_out_783     ),
    .col_in_784              ( u4_col_out_784     ),
    .col_in_785              ( u4_col_out_785     ),
    .col_in_786              ( u4_col_out_786     ),
    .col_in_787              ( u4_col_out_787     ),
    .col_in_788              ( u4_col_out_788     ),
    .col_in_789              ( u4_col_out_789     ),
    .col_in_790              ( u4_col_out_790     ),
    .col_in_791              ( u4_col_out_791     ),
    .col_in_792              ( u4_col_out_792     ),
    .col_in_793              ( u4_col_out_793     ),
    .col_in_794              ( u4_col_out_794     ),
    .col_in_795              ( u4_col_out_795     ),
    .col_in_796              ( u4_col_out_796     ),
    .col_in_797              ( u4_col_out_797     ),
    .col_in_798              ( u4_col_out_798     ),
    .col_in_799              ( u4_col_out_799     ),
    .col_in_800              ( u4_col_out_800     ),
    .col_in_801              ( u4_col_out_801     ),
    .col_in_802              ( u4_col_out_802     ),
    .col_in_803              ( u4_col_out_803     ),
    .col_in_804              ( u4_col_out_804     ),
    .col_in_805              ( u4_col_out_805     ),
    .col_in_806              ( u4_col_out_806     ),
    .col_in_807              ( u4_col_out_807     ),
    .col_in_808              ( u4_col_out_808     ),
    .col_in_809              ( u4_col_out_809     ),
    .col_in_810              ( u4_col_out_810     ),
    .col_in_811              ( u4_col_out_811     ),
    .col_in_812              ( u4_col_out_812     ),
    .col_in_813              ( u4_col_out_813     ),
    .col_in_814              ( u4_col_out_814     ),
    .col_in_815              ( u4_col_out_815     ),
    .col_in_816              ( u4_col_out_816     ),
    .col_in_817              ( u4_col_out_817     ),
    .col_in_818              ( u4_col_out_818     ),
    .col_in_819              ( u4_col_out_819     ),
    .col_in_820              ( u4_col_out_820     ),
    .col_in_821              ( u4_col_out_821     ),
    .col_in_822              ( u4_col_out_822     ),
    .col_in_823              ( u4_col_out_823     ),
    .col_in_824              ( u4_col_out_824     ),
    .col_in_825              ( u4_col_out_825     ),
    .col_in_826              ( u4_col_out_826     ),
    .col_in_827              ( u4_col_out_827     ),
    .col_in_828              ( u4_col_out_828     ),
    .col_in_829              ( u4_col_out_829     ),
    .col_in_830              ( u4_col_out_830     ),
    .col_in_831              ( u4_col_out_831     ),
    .col_in_832              ( u4_col_out_832     ),
    .col_in_833              ( u4_col_out_833     ),
    .col_in_834              ( u4_col_out_834     ),
    .col_in_835              ( u4_col_out_835     ),
    .col_in_836              ( u4_col_out_836     ),
    .col_in_837              ( u4_col_out_837     ),
    .col_in_838              ( u4_col_out_838     ),
    .col_in_839              ( u4_col_out_839     ),
    .col_in_840              ( u4_col_out_840     ),
    .col_in_841              ( u4_col_out_841     ),
    .col_in_842              ( u4_col_out_842     ),
    .col_in_843              ( u4_col_out_843     ),
    .col_in_844              ( u4_col_out_844     ),
    .col_in_845              ( u4_col_out_845     ),
    .col_in_846              ( u4_col_out_846     ),
    .col_in_847              ( u4_col_out_847     ),
    .col_in_848              ( u4_col_out_848     ),
    .col_in_849              ( u4_col_out_849     ),
    .col_in_850              ( u4_col_out_850     ),
    .col_in_851              ( u4_col_out_851     ),
    .col_in_852              ( u4_col_out_852     ),
    .col_in_853              ( u4_col_out_853     ),
    .col_in_854              ( u4_col_out_854     ),
    .col_in_855              ( u4_col_out_855     ),
    .col_in_856              ( u4_col_out_856     ),
    .col_in_857              ( u4_col_out_857     ),
    .col_in_858              ( u4_col_out_858     ),
    .col_in_859              ( u4_col_out_859     ),
    .col_in_860              ( u4_col_out_860     ),
    .col_in_861              ( u4_col_out_861     ),
    .col_in_862              ( u4_col_out_862     ),
    .col_in_863              ( u4_col_out_863     ),
    .col_in_864              ( u4_col_out_864     ),
    .col_in_865              ( u4_col_out_865     ),
    .col_in_866              ( u4_col_out_866     ),
    .col_in_867              ( u4_col_out_867     ),
    .col_in_868              ( u4_col_out_868     ),
    .col_in_869              ( u4_col_out_869     ),
    .col_in_870              ( u4_col_out_870     ),
    .col_in_871              ( u4_col_out_871     ),
    .col_in_872              ( u4_col_out_872     ),
    .col_in_873              ( u4_col_out_873     ),
    .col_in_874              ( u4_col_out_874     ),
    .col_in_875              ( u4_col_out_875     ),
    .col_in_876              ( u4_col_out_876     ),
    .col_in_877              ( u4_col_out_877     ),
    .col_in_878              ( u4_col_out_878     ),
    .col_in_879              ( u4_col_out_879     ),
    .col_in_880              ( u4_col_out_880     ),
    .col_in_881              ( u4_col_out_881     ),
    .col_in_882              ( u4_col_out_882     ),
    .col_in_883              ( u4_col_out_883     ),
    .col_in_884              ( u4_col_out_884     ),
    .col_in_885              ( u4_col_out_885     ),
    .col_in_886              ( u4_col_out_886     ),
    .col_in_887              ( u4_col_out_887     ),
    .col_in_888              ( u4_col_out_888     ),
    .col_in_889              ( u4_col_out_889     ),
    .col_in_890              ( u4_col_out_890     ),
    .col_in_891              ( u4_col_out_891     ),
    .col_in_892              ( u4_col_out_892     ),
    .col_in_893              ( u4_col_out_893     ),
    .col_in_894              ( u4_col_out_894     ),
    .col_in_895              ( u4_col_out_895     ),
    .col_in_896              ( u4_col_out_896     ),
    .col_in_897              ( u4_col_out_897     ),
    .col_in_898              ( u4_col_out_898     ),
    .col_in_899              ( u4_col_out_899     ),
    .col_in_900              ( u4_col_out_900     ),
    .col_in_901              ( u4_col_out_901     ),
    .col_in_902              ( u4_col_out_902     ),
    .col_in_903              ( u4_col_out_903     ),
    .col_in_904              ( u4_col_out_904     ),
    .col_in_905              ( u4_col_out_905     ),
    .col_in_906              ( u4_col_out_906     ),
    .col_in_907              ( u4_col_out_907     ),
    .col_in_908              ( u4_col_out_908     ),
    .col_in_909              ( u4_col_out_909     ),
    .col_in_910              ( u4_col_out_910     ),
    .col_in_911              ( u4_col_out_911     ),
    .col_in_912              ( u4_col_out_912     ),
    .col_in_913              ( u4_col_out_913     ),
    .col_in_914              ( u4_col_out_914     ),
    .col_in_915              ( u4_col_out_915     ),
    .col_in_916              ( u4_col_out_916     ),
    .col_in_917              ( u4_col_out_917     ),
    .col_in_918              ( u4_col_out_918     ),
    .col_in_919              ( u4_col_out_919     ),
    .col_in_920              ( u4_col_out_920     ),
    .col_in_921              ( u4_col_out_921     ),
    .col_in_922              ( u4_col_out_922     ),
    .col_in_923              ( u4_col_out_923     ),
    .col_in_924              ( u4_col_out_924     ),
    .col_in_925              ( u4_col_out_925     ),
    .col_in_926              ( u4_col_out_926     ),
    .col_in_927              ( u4_col_out_927     ),
    .col_in_928              ( u4_col_out_928     ),
    .col_in_929              ( u4_col_out_929     ),
    .col_in_930              ( u4_col_out_930     ),
    .col_in_931              ( u4_col_out_931     ),
    .col_in_932              ( u4_col_out_932     ),
    .col_in_933              ( u4_col_out_933     ),
    .col_in_934              ( u4_col_out_934     ),
    .col_in_935              ( u4_col_out_935     ),
    .col_in_936              ( u4_col_out_936     ),
    .col_in_937              ( u4_col_out_937     ),
    .col_in_938              ( u4_col_out_938     ),
    .col_in_939              ( u4_col_out_939     ),
    .col_in_940              ( u4_col_out_940     ),
    .col_in_941              ( u4_col_out_941     ),
    .col_in_942              ( u4_col_out_942     ),
    .col_in_943              ( u4_col_out_943     ),
    .col_in_944              ( u4_col_out_944     ),
    .col_in_945              ( u4_col_out_945     ),
    .col_in_946              ( u4_col_out_946     ),
    .col_in_947              ( u4_col_out_947     ),
    .col_in_948              ( u4_col_out_948     ),
    .col_in_949              ( u4_col_out_949     ),
    .col_in_950              ( u4_col_out_950     ),
    .col_in_951              ( u4_col_out_951     ),
    .col_in_952              ( u4_col_out_952     ),
    .col_in_953              ( u4_col_out_953     ),
    .col_in_954              ( u4_col_out_954     ),
    .col_in_955              ( u4_col_out_955     ),
    .col_in_956              ( u4_col_out_956     ),
    .col_in_957              ( u4_col_out_957     ),
    .col_in_958              ( u4_col_out_958     ),
    .col_in_959              ( u4_col_out_959     ),
    .col_in_960              ( u4_col_out_960     ),
    .col_in_961              ( u4_col_out_961     ),
    .col_in_962              ( u4_col_out_962     ),
    .col_in_963              ( u4_col_out_963     ),
    .col_in_964              ( u4_col_out_964     ),
    .col_in_965              ( u4_col_out_965     ),
    .col_in_966              ( u4_col_out_966     ),
    .col_in_967              ( u4_col_out_967     ),
    .col_in_968              ( u4_col_out_968     ),
    .col_in_969              ( u4_col_out_969     ),
    .col_in_970              ( u4_col_out_970     ),
    .col_in_971              ( u4_col_out_971     ),
    .col_in_972              ( u4_col_out_972     ),
    .col_in_973              ( u4_col_out_973     ),
    .col_in_974              ( u4_col_out_974     ),
    .col_in_975              ( u4_col_out_975     ),
    .col_in_976              ( u4_col_out_976     ),
    .col_in_977              ( u4_col_out_977     ),
    .col_in_978              ( u4_col_out_978     ),
    .col_in_979              ( u4_col_out_979     ),
    .col_in_980              ( u4_col_out_980     ),
    .col_in_981              ( u4_col_out_981     ),
    .col_in_982              ( u4_col_out_982     ),
    .col_in_983              ( u4_col_out_983     ),
    .col_in_984              ( u4_col_out_984     ),
    .col_in_985              ( u4_col_out_985     ),
    .col_in_986              ( u4_col_out_986     ),
    .col_in_987              ( u4_col_out_987     ),
    .col_in_988              ( u4_col_out_988     ),
    .col_in_989              ( u4_col_out_989     ),
    .col_in_990              ( u4_col_out_990     ),
    .col_in_991              ( u4_col_out_991     ),
    .col_in_992              ( u4_col_out_992     ),
    .col_in_993              ( u4_col_out_993     ),
    .col_in_994              ( u4_col_out_994     ),
    .col_in_995              ( u4_col_out_995     ),
    .col_in_996              ( u4_col_out_996     ),
    .col_in_997              ( u4_col_out_997     ),
    .col_in_998              ( u4_col_out_998     ),
    .col_in_999              ( u4_col_out_999     ),
    .col_in_1000             ( u4_col_out_1000    ),
    .col_in_1001             ( u4_col_out_1001    ),
    .col_in_1002             ( u4_col_out_1002    ),
    .col_in_1003             ( u4_col_out_1003    ),
    .col_in_1004             ( u4_col_out_1004    ),
    .col_in_1005             ( u4_col_out_1005    ),
    .col_in_1006             ( u4_col_out_1006    ),
    .col_in_1007             ( u4_col_out_1007    ),
    .col_in_1008             ( u4_col_out_1008    ),
    .col_in_1009             ( u4_col_out_1009    ),
    .col_in_1010             ( u4_col_out_1010    ),
    .col_in_1011             ( u4_col_out_1011    ),
    .col_in_1012             ( u4_col_out_1012    ),
    .col_in_1013             ( u4_col_out_1013    ),
    .col_in_1014             ( u4_col_out_1014    ),
    .col_in_1015             ( u4_col_out_1015    ),
    .col_in_1016             ( u4_col_out_1016    ),
    .col_in_1017             ( u4_col_out_1017    ),
    .col_in_1018             ( u4_col_out_1018    ),
    .col_in_1019             ( u4_col_out_1019    ),
    .col_in_1020             ( u4_col_out_1020    ),
    .col_in_1021             ( u4_col_out_1021    ),
    .col_in_1022             ( u4_col_out_1022    ),
    .col_in_1023             ( u4_col_out_1023    ),
    .col_in_1024             ( u4_col_out_1024    ),
    .col_in_1025             ( u4_col_out_1025    ),
    .col_in_1026             ( u4_col_out_1026    ),
    .col_in_1027             ( u4_col_out_1027    ),
    .col_in_1028             ( u4_col_out_1028    ),
    .col_in_1029             ( u4_col_out_1029    ),
    .col_in_1030             ( u4_col_out_1030    ),
    .col_in_1031             ( u4_col_out_1031    ),
    .col_in_1032             ( u4_col_out_1032    ),


    .col_out_0               ( u5_col_out_0      ),
    .col_out_1               ( u5_col_out_1      ),
    .col_out_2               ( u5_col_out_2      ),
    .col_out_3               ( u5_col_out_3      ),
    .col_out_4               ( u5_col_out_4      ),
    .col_out_5               ( u5_col_out_5      ),
    .col_out_6               ( u5_col_out_6      ),
    .col_out_7               ( u5_col_out_7      ),
    .col_out_8               ( u5_col_out_8      ),
    .col_out_9               ( u5_col_out_9      ),
    .col_out_10              ( u5_col_out_10     ),
    .col_out_11              ( u5_col_out_11     ),
    .col_out_12              ( u5_col_out_12     ),
    .col_out_13              ( u5_col_out_13     ),
    .col_out_14              ( u5_col_out_14     ),
    .col_out_15              ( u5_col_out_15     ),
    .col_out_16              ( u5_col_out_16     ),
    .col_out_17              ( u5_col_out_17     ),
    .col_out_18              ( u5_col_out_18     ),
    .col_out_19              ( u5_col_out_19     ),
    .col_out_20              ( u5_col_out_20     ),
    .col_out_21              ( u5_col_out_21     ),
    .col_out_22              ( u5_col_out_22     ),
    .col_out_23              ( u5_col_out_23     ),
    .col_out_24              ( u5_col_out_24     ),
    .col_out_25              ( u5_col_out_25     ),
    .col_out_26              ( u5_col_out_26     ),
    .col_out_27              ( u5_col_out_27     ),
    .col_out_28              ( u5_col_out_28     ),
    .col_out_29              ( u5_col_out_29     ),
    .col_out_30              ( u5_col_out_30     ),
    .col_out_31              ( u5_col_out_31     ),
    .col_out_32              ( u5_col_out_32     ),
    .col_out_33              ( u5_col_out_33     ),
    .col_out_34              ( u5_col_out_34     ),
    .col_out_35              ( u5_col_out_35     ),
    .col_out_36              ( u5_col_out_36     ),
    .col_out_37              ( u5_col_out_37     ),
    .col_out_38              ( u5_col_out_38     ),
    .col_out_39              ( u5_col_out_39     ),
    .col_out_40              ( u5_col_out_40     ),
    .col_out_41              ( u5_col_out_41     ),
    .col_out_42              ( u5_col_out_42     ),
    .col_out_43              ( u5_col_out_43     ),
    .col_out_44              ( u5_col_out_44     ),
    .col_out_45              ( u5_col_out_45     ),
    .col_out_46              ( u5_col_out_46     ),
    .col_out_47              ( u5_col_out_47     ),
    .col_out_48              ( u5_col_out_48     ),
    .col_out_49              ( u5_col_out_49     ),
    .col_out_50              ( u5_col_out_50     ),
    .col_out_51              ( u5_col_out_51     ),
    .col_out_52              ( u5_col_out_52     ),
    .col_out_53              ( u5_col_out_53     ),
    .col_out_54              ( u5_col_out_54     ),
    .col_out_55              ( u5_col_out_55     ),
    .col_out_56              ( u5_col_out_56     ),
    .col_out_57              ( u5_col_out_57     ),
    .col_out_58              ( u5_col_out_58     ),
    .col_out_59              ( u5_col_out_59     ),
    .col_out_60              ( u5_col_out_60     ),
    .col_out_61              ( u5_col_out_61     ),
    .col_out_62              ( u5_col_out_62     ),
    .col_out_63              ( u5_col_out_63     ),
    .col_out_64              ( u5_col_out_64     ),
    .col_out_65              ( u5_col_out_65     ),
    .col_out_66              ( u5_col_out_66     ),
    .col_out_67              ( u5_col_out_67     ),
    .col_out_68              ( u5_col_out_68     ),
    .col_out_69              ( u5_col_out_69     ),
    .col_out_70              ( u5_col_out_70     ),
    .col_out_71              ( u5_col_out_71     ),
    .col_out_72              ( u5_col_out_72     ),
    .col_out_73              ( u5_col_out_73     ),
    .col_out_74              ( u5_col_out_74     ),
    .col_out_75              ( u5_col_out_75     ),
    .col_out_76              ( u5_col_out_76     ),
    .col_out_77              ( u5_col_out_77     ),
    .col_out_78              ( u5_col_out_78     ),
    .col_out_79              ( u5_col_out_79     ),
    .col_out_80              ( u5_col_out_80     ),
    .col_out_81              ( u5_col_out_81     ),
    .col_out_82              ( u5_col_out_82     ),
    .col_out_83              ( u5_col_out_83     ),
    .col_out_84              ( u5_col_out_84     ),
    .col_out_85              ( u5_col_out_85     ),
    .col_out_86              ( u5_col_out_86     ),
    .col_out_87              ( u5_col_out_87     ),
    .col_out_88              ( u5_col_out_88     ),
    .col_out_89              ( u5_col_out_89     ),
    .col_out_90              ( u5_col_out_90     ),
    .col_out_91              ( u5_col_out_91     ),
    .col_out_92              ( u5_col_out_92     ),
    .col_out_93              ( u5_col_out_93     ),
    .col_out_94              ( u5_col_out_94     ),
    .col_out_95              ( u5_col_out_95     ),
    .col_out_96              ( u5_col_out_96     ),
    .col_out_97              ( u5_col_out_97     ),
    .col_out_98              ( u5_col_out_98     ),
    .col_out_99              ( u5_col_out_99     ),
    .col_out_100             ( u5_col_out_100    ),
    .col_out_101             ( u5_col_out_101    ),
    .col_out_102             ( u5_col_out_102    ),
    .col_out_103             ( u5_col_out_103    ),
    .col_out_104             ( u5_col_out_104    ),
    .col_out_105             ( u5_col_out_105    ),
    .col_out_106             ( u5_col_out_106    ),
    .col_out_107             ( u5_col_out_107    ),
    .col_out_108             ( u5_col_out_108    ),
    .col_out_109             ( u5_col_out_109    ),
    .col_out_110             ( u5_col_out_110    ),
    .col_out_111             ( u5_col_out_111    ),
    .col_out_112             ( u5_col_out_112    ),
    .col_out_113             ( u5_col_out_113    ),
    .col_out_114             ( u5_col_out_114    ),
    .col_out_115             ( u5_col_out_115    ),
    .col_out_116             ( u5_col_out_116    ),
    .col_out_117             ( u5_col_out_117    ),
    .col_out_118             ( u5_col_out_118    ),
    .col_out_119             ( u5_col_out_119    ),
    .col_out_120             ( u5_col_out_120    ),
    .col_out_121             ( u5_col_out_121    ),
    .col_out_122             ( u5_col_out_122    ),
    .col_out_123             ( u5_col_out_123    ),
    .col_out_124             ( u5_col_out_124    ),
    .col_out_125             ( u5_col_out_125    ),
    .col_out_126             ( u5_col_out_126    ),
    .col_out_127             ( u5_col_out_127    ),
    .col_out_128             ( u5_col_out_128    ),
    .col_out_129             ( u5_col_out_129    ),
    .col_out_130             ( u5_col_out_130    ),
    .col_out_131             ( u5_col_out_131    ),
    .col_out_132             ( u5_col_out_132    ),
    .col_out_133             ( u5_col_out_133    ),
    .col_out_134             ( u5_col_out_134    ),
    .col_out_135             ( u5_col_out_135    ),
    .col_out_136             ( u5_col_out_136    ),
    .col_out_137             ( u5_col_out_137    ),
    .col_out_138             ( u5_col_out_138    ),
    .col_out_139             ( u5_col_out_139    ),
    .col_out_140             ( u5_col_out_140    ),
    .col_out_141             ( u5_col_out_141    ),
    .col_out_142             ( u5_col_out_142    ),
    .col_out_143             ( u5_col_out_143    ),
    .col_out_144             ( u5_col_out_144    ),
    .col_out_145             ( u5_col_out_145    ),
    .col_out_146             ( u5_col_out_146    ),
    .col_out_147             ( u5_col_out_147    ),
    .col_out_148             ( u5_col_out_148    ),
    .col_out_149             ( u5_col_out_149    ),
    .col_out_150             ( u5_col_out_150    ),
    .col_out_151             ( u5_col_out_151    ),
    .col_out_152             ( u5_col_out_152    ),
    .col_out_153             ( u5_col_out_153    ),
    .col_out_154             ( u5_col_out_154    ),
    .col_out_155             ( u5_col_out_155    ),
    .col_out_156             ( u5_col_out_156    ),
    .col_out_157             ( u5_col_out_157    ),
    .col_out_158             ( u5_col_out_158    ),
    .col_out_159             ( u5_col_out_159    ),
    .col_out_160             ( u5_col_out_160    ),
    .col_out_161             ( u5_col_out_161    ),
    .col_out_162             ( u5_col_out_162    ),
    .col_out_163             ( u5_col_out_163    ),
    .col_out_164             ( u5_col_out_164    ),
    .col_out_165             ( u5_col_out_165    ),
    .col_out_166             ( u5_col_out_166    ),
    .col_out_167             ( u5_col_out_167    ),
    .col_out_168             ( u5_col_out_168    ),
    .col_out_169             ( u5_col_out_169    ),
    .col_out_170             ( u5_col_out_170    ),
    .col_out_171             ( u5_col_out_171    ),
    .col_out_172             ( u5_col_out_172    ),
    .col_out_173             ( u5_col_out_173    ),
    .col_out_174             ( u5_col_out_174    ),
    .col_out_175             ( u5_col_out_175    ),
    .col_out_176             ( u5_col_out_176    ),
    .col_out_177             ( u5_col_out_177    ),
    .col_out_178             ( u5_col_out_178    ),
    .col_out_179             ( u5_col_out_179    ),
    .col_out_180             ( u5_col_out_180    ),
    .col_out_181             ( u5_col_out_181    ),
    .col_out_182             ( u5_col_out_182    ),
    .col_out_183             ( u5_col_out_183    ),
    .col_out_184             ( u5_col_out_184    ),
    .col_out_185             ( u5_col_out_185    ),
    .col_out_186             ( u5_col_out_186    ),
    .col_out_187             ( u5_col_out_187    ),
    .col_out_188             ( u5_col_out_188    ),
    .col_out_189             ( u5_col_out_189    ),
    .col_out_190             ( u5_col_out_190    ),
    .col_out_191             ( u5_col_out_191    ),
    .col_out_192             ( u5_col_out_192    ),
    .col_out_193             ( u5_col_out_193    ),
    .col_out_194             ( u5_col_out_194    ),
    .col_out_195             ( u5_col_out_195    ),
    .col_out_196             ( u5_col_out_196    ),
    .col_out_197             ( u5_col_out_197    ),
    .col_out_198             ( u5_col_out_198    ),
    .col_out_199             ( u5_col_out_199    ),
    .col_out_200             ( u5_col_out_200    ),
    .col_out_201             ( u5_col_out_201    ),
    .col_out_202             ( u5_col_out_202    ),
    .col_out_203             ( u5_col_out_203    ),
    .col_out_204             ( u5_col_out_204    ),
    .col_out_205             ( u5_col_out_205    ),
    .col_out_206             ( u5_col_out_206    ),
    .col_out_207             ( u5_col_out_207    ),
    .col_out_208             ( u5_col_out_208    ),
    .col_out_209             ( u5_col_out_209    ),
    .col_out_210             ( u5_col_out_210    ),
    .col_out_211             ( u5_col_out_211    ),
    .col_out_212             ( u5_col_out_212    ),
    .col_out_213             ( u5_col_out_213    ),
    .col_out_214             ( u5_col_out_214    ),
    .col_out_215             ( u5_col_out_215    ),
    .col_out_216             ( u5_col_out_216    ),
    .col_out_217             ( u5_col_out_217    ),
    .col_out_218             ( u5_col_out_218    ),
    .col_out_219             ( u5_col_out_219    ),
    .col_out_220             ( u5_col_out_220    ),
    .col_out_221             ( u5_col_out_221    ),
    .col_out_222             ( u5_col_out_222    ),
    .col_out_223             ( u5_col_out_223    ),
    .col_out_224             ( u5_col_out_224    ),
    .col_out_225             ( u5_col_out_225    ),
    .col_out_226             ( u5_col_out_226    ),
    .col_out_227             ( u5_col_out_227    ),
    .col_out_228             ( u5_col_out_228    ),
    .col_out_229             ( u5_col_out_229    ),
    .col_out_230             ( u5_col_out_230    ),
    .col_out_231             ( u5_col_out_231    ),
    .col_out_232             ( u5_col_out_232    ),
    .col_out_233             ( u5_col_out_233    ),
    .col_out_234             ( u5_col_out_234    ),
    .col_out_235             ( u5_col_out_235    ),
    .col_out_236             ( u5_col_out_236    ),
    .col_out_237             ( u5_col_out_237    ),
    .col_out_238             ( u5_col_out_238    ),
    .col_out_239             ( u5_col_out_239    ),
    .col_out_240             ( u5_col_out_240    ),
    .col_out_241             ( u5_col_out_241    ),
    .col_out_242             ( u5_col_out_242    ),
    .col_out_243             ( u5_col_out_243    ),
    .col_out_244             ( u5_col_out_244    ),
    .col_out_245             ( u5_col_out_245    ),
    .col_out_246             ( u5_col_out_246    ),
    .col_out_247             ( u5_col_out_247    ),
    .col_out_248             ( u5_col_out_248    ),
    .col_out_249             ( u5_col_out_249    ),
    .col_out_250             ( u5_col_out_250    ),
    .col_out_251             ( u5_col_out_251    ),
    .col_out_252             ( u5_col_out_252    ),
    .col_out_253             ( u5_col_out_253    ),
    .col_out_254             ( u5_col_out_254    ),
    .col_out_255             ( u5_col_out_255    ),
    .col_out_256             ( u5_col_out_256    ),
    .col_out_257             ( u5_col_out_257    ),
    .col_out_258             ( u5_col_out_258    ),
    .col_out_259             ( u5_col_out_259    ),
    .col_out_260             ( u5_col_out_260    ),
    .col_out_261             ( u5_col_out_261    ),
    .col_out_262             ( u5_col_out_262    ),
    .col_out_263             ( u5_col_out_263    ),
    .col_out_264             ( u5_col_out_264    ),
    .col_out_265             ( u5_col_out_265    ),
    .col_out_266             ( u5_col_out_266    ),
    .col_out_267             ( u5_col_out_267    ),
    .col_out_268             ( u5_col_out_268    ),
    .col_out_269             ( u5_col_out_269    ),
    .col_out_270             ( u5_col_out_270    ),
    .col_out_271             ( u5_col_out_271    ),
    .col_out_272             ( u5_col_out_272    ),
    .col_out_273             ( u5_col_out_273    ),
    .col_out_274             ( u5_col_out_274    ),
    .col_out_275             ( u5_col_out_275    ),
    .col_out_276             ( u5_col_out_276    ),
    .col_out_277             ( u5_col_out_277    ),
    .col_out_278             ( u5_col_out_278    ),
    .col_out_279             ( u5_col_out_279    ),
    .col_out_280             ( u5_col_out_280    ),
    .col_out_281             ( u5_col_out_281    ),
    .col_out_282             ( u5_col_out_282    ),
    .col_out_283             ( u5_col_out_283    ),
    .col_out_284             ( u5_col_out_284    ),
    .col_out_285             ( u5_col_out_285    ),
    .col_out_286             ( u5_col_out_286    ),
    .col_out_287             ( u5_col_out_287    ),
    .col_out_288             ( u5_col_out_288    ),
    .col_out_289             ( u5_col_out_289    ),
    .col_out_290             ( u5_col_out_290    ),
    .col_out_291             ( u5_col_out_291    ),
    .col_out_292             ( u5_col_out_292    ),
    .col_out_293             ( u5_col_out_293    ),
    .col_out_294             ( u5_col_out_294    ),
    .col_out_295             ( u5_col_out_295    ),
    .col_out_296             ( u5_col_out_296    ),
    .col_out_297             ( u5_col_out_297    ),
    .col_out_298             ( u5_col_out_298    ),
    .col_out_299             ( u5_col_out_299    ),
    .col_out_300             ( u5_col_out_300    ),
    .col_out_301             ( u5_col_out_301    ),
    .col_out_302             ( u5_col_out_302    ),
    .col_out_303             ( u5_col_out_303    ),
    .col_out_304             ( u5_col_out_304    ),
    .col_out_305             ( u5_col_out_305    ),
    .col_out_306             ( u5_col_out_306    ),
    .col_out_307             ( u5_col_out_307    ),
    .col_out_308             ( u5_col_out_308    ),
    .col_out_309             ( u5_col_out_309    ),
    .col_out_310             ( u5_col_out_310    ),
    .col_out_311             ( u5_col_out_311    ),
    .col_out_312             ( u5_col_out_312    ),
    .col_out_313             ( u5_col_out_313    ),
    .col_out_314             ( u5_col_out_314    ),
    .col_out_315             ( u5_col_out_315    ),
    .col_out_316             ( u5_col_out_316    ),
    .col_out_317             ( u5_col_out_317    ),
    .col_out_318             ( u5_col_out_318    ),
    .col_out_319             ( u5_col_out_319    ),
    .col_out_320             ( u5_col_out_320    ),
    .col_out_321             ( u5_col_out_321    ),
    .col_out_322             ( u5_col_out_322    ),
    .col_out_323             ( u5_col_out_323    ),
    .col_out_324             ( u5_col_out_324    ),
    .col_out_325             ( u5_col_out_325    ),
    .col_out_326             ( u5_col_out_326    ),
    .col_out_327             ( u5_col_out_327    ),
    .col_out_328             ( u5_col_out_328    ),
    .col_out_329             ( u5_col_out_329    ),
    .col_out_330             ( u5_col_out_330    ),
    .col_out_331             ( u5_col_out_331    ),
    .col_out_332             ( u5_col_out_332    ),
    .col_out_333             ( u5_col_out_333    ),
    .col_out_334             ( u5_col_out_334    ),
    .col_out_335             ( u5_col_out_335    ),
    .col_out_336             ( u5_col_out_336    ),
    .col_out_337             ( u5_col_out_337    ),
    .col_out_338             ( u5_col_out_338    ),
    .col_out_339             ( u5_col_out_339    ),
    .col_out_340             ( u5_col_out_340    ),
    .col_out_341             ( u5_col_out_341    ),
    .col_out_342             ( u5_col_out_342    ),
    .col_out_343             ( u5_col_out_343    ),
    .col_out_344             ( u5_col_out_344    ),
    .col_out_345             ( u5_col_out_345    ),
    .col_out_346             ( u5_col_out_346    ),
    .col_out_347             ( u5_col_out_347    ),
    .col_out_348             ( u5_col_out_348    ),
    .col_out_349             ( u5_col_out_349    ),
    .col_out_350             ( u5_col_out_350    ),
    .col_out_351             ( u5_col_out_351    ),
    .col_out_352             ( u5_col_out_352    ),
    .col_out_353             ( u5_col_out_353    ),
    .col_out_354             ( u5_col_out_354    ),
    .col_out_355             ( u5_col_out_355    ),
    .col_out_356             ( u5_col_out_356    ),
    .col_out_357             ( u5_col_out_357    ),
    .col_out_358             ( u5_col_out_358    ),
    .col_out_359             ( u5_col_out_359    ),
    .col_out_360             ( u5_col_out_360    ),
    .col_out_361             ( u5_col_out_361    ),
    .col_out_362             ( u5_col_out_362    ),
    .col_out_363             ( u5_col_out_363    ),
    .col_out_364             ( u5_col_out_364    ),
    .col_out_365             ( u5_col_out_365    ),
    .col_out_366             ( u5_col_out_366    ),
    .col_out_367             ( u5_col_out_367    ),
    .col_out_368             ( u5_col_out_368    ),
    .col_out_369             ( u5_col_out_369    ),
    .col_out_370             ( u5_col_out_370    ),
    .col_out_371             ( u5_col_out_371    ),
    .col_out_372             ( u5_col_out_372    ),
    .col_out_373             ( u5_col_out_373    ),
    .col_out_374             ( u5_col_out_374    ),
    .col_out_375             ( u5_col_out_375    ),
    .col_out_376             ( u5_col_out_376    ),
    .col_out_377             ( u5_col_out_377    ),
    .col_out_378             ( u5_col_out_378    ),
    .col_out_379             ( u5_col_out_379    ),
    .col_out_380             ( u5_col_out_380    ),
    .col_out_381             ( u5_col_out_381    ),
    .col_out_382             ( u5_col_out_382    ),
    .col_out_383             ( u5_col_out_383    ),
    .col_out_384             ( u5_col_out_384    ),
    .col_out_385             ( u5_col_out_385    ),
    .col_out_386             ( u5_col_out_386    ),
    .col_out_387             ( u5_col_out_387    ),
    .col_out_388             ( u5_col_out_388    ),
    .col_out_389             ( u5_col_out_389    ),
    .col_out_390             ( u5_col_out_390    ),
    .col_out_391             ( u5_col_out_391    ),
    .col_out_392             ( u5_col_out_392    ),
    .col_out_393             ( u5_col_out_393    ),
    .col_out_394             ( u5_col_out_394    ),
    .col_out_395             ( u5_col_out_395    ),
    .col_out_396             ( u5_col_out_396    ),
    .col_out_397             ( u5_col_out_397    ),
    .col_out_398             ( u5_col_out_398    ),
    .col_out_399             ( u5_col_out_399    ),
    .col_out_400             ( u5_col_out_400    ),
    .col_out_401             ( u5_col_out_401    ),
    .col_out_402             ( u5_col_out_402    ),
    .col_out_403             ( u5_col_out_403    ),
    .col_out_404             ( u5_col_out_404    ),
    .col_out_405             ( u5_col_out_405    ),
    .col_out_406             ( u5_col_out_406    ),
    .col_out_407             ( u5_col_out_407    ),
    .col_out_408             ( u5_col_out_408    ),
    .col_out_409             ( u5_col_out_409    ),
    .col_out_410             ( u5_col_out_410    ),
    .col_out_411             ( u5_col_out_411    ),
    .col_out_412             ( u5_col_out_412    ),
    .col_out_413             ( u5_col_out_413    ),
    .col_out_414             ( u5_col_out_414    ),
    .col_out_415             ( u5_col_out_415    ),
    .col_out_416             ( u5_col_out_416    ),
    .col_out_417             ( u5_col_out_417    ),
    .col_out_418             ( u5_col_out_418    ),
    .col_out_419             ( u5_col_out_419    ),
    .col_out_420             ( u5_col_out_420    ),
    .col_out_421             ( u5_col_out_421    ),
    .col_out_422             ( u5_col_out_422    ),
    .col_out_423             ( u5_col_out_423    ),
    .col_out_424             ( u5_col_out_424    ),
    .col_out_425             ( u5_col_out_425    ),
    .col_out_426             ( u5_col_out_426    ),
    .col_out_427             ( u5_col_out_427    ),
    .col_out_428             ( u5_col_out_428    ),
    .col_out_429             ( u5_col_out_429    ),
    .col_out_430             ( u5_col_out_430    ),
    .col_out_431             ( u5_col_out_431    ),
    .col_out_432             ( u5_col_out_432    ),
    .col_out_433             ( u5_col_out_433    ),
    .col_out_434             ( u5_col_out_434    ),
    .col_out_435             ( u5_col_out_435    ),
    .col_out_436             ( u5_col_out_436    ),
    .col_out_437             ( u5_col_out_437    ),
    .col_out_438             ( u5_col_out_438    ),
    .col_out_439             ( u5_col_out_439    ),
    .col_out_440             ( u5_col_out_440    ),
    .col_out_441             ( u5_col_out_441    ),
    .col_out_442             ( u5_col_out_442    ),
    .col_out_443             ( u5_col_out_443    ),
    .col_out_444             ( u5_col_out_444    ),
    .col_out_445             ( u5_col_out_445    ),
    .col_out_446             ( u5_col_out_446    ),
    .col_out_447             ( u5_col_out_447    ),
    .col_out_448             ( u5_col_out_448    ),
    .col_out_449             ( u5_col_out_449    ),
    .col_out_450             ( u5_col_out_450    ),
    .col_out_451             ( u5_col_out_451    ),
    .col_out_452             ( u5_col_out_452    ),
    .col_out_453             ( u5_col_out_453    ),
    .col_out_454             ( u5_col_out_454    ),
    .col_out_455             ( u5_col_out_455    ),
    .col_out_456             ( u5_col_out_456    ),
    .col_out_457             ( u5_col_out_457    ),
    .col_out_458             ( u5_col_out_458    ),
    .col_out_459             ( u5_col_out_459    ),
    .col_out_460             ( u5_col_out_460    ),
    .col_out_461             ( u5_col_out_461    ),
    .col_out_462             ( u5_col_out_462    ),
    .col_out_463             ( u5_col_out_463    ),
    .col_out_464             ( u5_col_out_464    ),
    .col_out_465             ( u5_col_out_465    ),
    .col_out_466             ( u5_col_out_466    ),
    .col_out_467             ( u5_col_out_467    ),
    .col_out_468             ( u5_col_out_468    ),
    .col_out_469             ( u5_col_out_469    ),
    .col_out_470             ( u5_col_out_470    ),
    .col_out_471             ( u5_col_out_471    ),
    .col_out_472             ( u5_col_out_472    ),
    .col_out_473             ( u5_col_out_473    ),
    .col_out_474             ( u5_col_out_474    ),
    .col_out_475             ( u5_col_out_475    ),
    .col_out_476             ( u5_col_out_476    ),
    .col_out_477             ( u5_col_out_477    ),
    .col_out_478             ( u5_col_out_478    ),
    .col_out_479             ( u5_col_out_479    ),
    .col_out_480             ( u5_col_out_480    ),
    .col_out_481             ( u5_col_out_481    ),
    .col_out_482             ( u5_col_out_482    ),
    .col_out_483             ( u5_col_out_483    ),
    .col_out_484             ( u5_col_out_484    ),
    .col_out_485             ( u5_col_out_485    ),
    .col_out_486             ( u5_col_out_486    ),
    .col_out_487             ( u5_col_out_487    ),
    .col_out_488             ( u5_col_out_488    ),
    .col_out_489             ( u5_col_out_489    ),
    .col_out_490             ( u5_col_out_490    ),
    .col_out_491             ( u5_col_out_491    ),
    .col_out_492             ( u5_col_out_492    ),
    .col_out_493             ( u5_col_out_493    ),
    .col_out_494             ( u5_col_out_494    ),
    .col_out_495             ( u5_col_out_495    ),
    .col_out_496             ( u5_col_out_496    ),
    .col_out_497             ( u5_col_out_497    ),
    .col_out_498             ( u5_col_out_498    ),
    .col_out_499             ( u5_col_out_499    ),
    .col_out_500             ( u5_col_out_500    ),
    .col_out_501             ( u5_col_out_501    ),
    .col_out_502             ( u5_col_out_502    ),
    .col_out_503             ( u5_col_out_503    ),
    .col_out_504             ( u5_col_out_504    ),
    .col_out_505             ( u5_col_out_505    ),
    .col_out_506             ( u5_col_out_506    ),
    .col_out_507             ( u5_col_out_507    ),
    .col_out_508             ( u5_col_out_508    ),
    .col_out_509             ( u5_col_out_509    ),
    .col_out_510             ( u5_col_out_510    ),
    .col_out_511             ( u5_col_out_511    ),
    .col_out_512             ( u5_col_out_512    ),
    .col_out_513             ( u5_col_out_513    ),
    .col_out_514             ( u5_col_out_514    ),
    .col_out_515             ( u5_col_out_515    ),
    .col_out_516             ( u5_col_out_516    ),
    .col_out_517             ( u5_col_out_517    ),
    .col_out_518             ( u5_col_out_518    ),
    .col_out_519             ( u5_col_out_519    ),
    .col_out_520             ( u5_col_out_520    ),
    .col_out_521             ( u5_col_out_521    ),
    .col_out_522             ( u5_col_out_522    ),
    .col_out_523             ( u5_col_out_523    ),
    .col_out_524             ( u5_col_out_524    ),
    .col_out_525             ( u5_col_out_525    ),
    .col_out_526             ( u5_col_out_526    ),
    .col_out_527             ( u5_col_out_527    ),
    .col_out_528             ( u5_col_out_528    ),
    .col_out_529             ( u5_col_out_529    ),
    .col_out_530             ( u5_col_out_530    ),
    .col_out_531             ( u5_col_out_531    ),
    .col_out_532             ( u5_col_out_532    ),
    .col_out_533             ( u5_col_out_533    ),
    .col_out_534             ( u5_col_out_534    ),
    .col_out_535             ( u5_col_out_535    ),
    .col_out_536             ( u5_col_out_536    ),
    .col_out_537             ( u5_col_out_537    ),
    .col_out_538             ( u5_col_out_538    ),
    .col_out_539             ( u5_col_out_539    ),
    .col_out_540             ( u5_col_out_540    ),
    .col_out_541             ( u5_col_out_541    ),
    .col_out_542             ( u5_col_out_542    ),
    .col_out_543             ( u5_col_out_543    ),
    .col_out_544             ( u5_col_out_544    ),
    .col_out_545             ( u5_col_out_545    ),
    .col_out_546             ( u5_col_out_546    ),
    .col_out_547             ( u5_col_out_547    ),
    .col_out_548             ( u5_col_out_548    ),
    .col_out_549             ( u5_col_out_549    ),
    .col_out_550             ( u5_col_out_550    ),
    .col_out_551             ( u5_col_out_551    ),
    .col_out_552             ( u5_col_out_552    ),
    .col_out_553             ( u5_col_out_553    ),
    .col_out_554             ( u5_col_out_554    ),
    .col_out_555             ( u5_col_out_555    ),
    .col_out_556             ( u5_col_out_556    ),
    .col_out_557             ( u5_col_out_557    ),
    .col_out_558             ( u5_col_out_558    ),
    .col_out_559             ( u5_col_out_559    ),
    .col_out_560             ( u5_col_out_560    ),
    .col_out_561             ( u5_col_out_561    ),
    .col_out_562             ( u5_col_out_562    ),
    .col_out_563             ( u5_col_out_563    ),
    .col_out_564             ( u5_col_out_564    ),
    .col_out_565             ( u5_col_out_565    ),
    .col_out_566             ( u5_col_out_566    ),
    .col_out_567             ( u5_col_out_567    ),
    .col_out_568             ( u5_col_out_568    ),
    .col_out_569             ( u5_col_out_569    ),
    .col_out_570             ( u5_col_out_570    ),
    .col_out_571             ( u5_col_out_571    ),
    .col_out_572             ( u5_col_out_572    ),
    .col_out_573             ( u5_col_out_573    ),
    .col_out_574             ( u5_col_out_574    ),
    .col_out_575             ( u5_col_out_575    ),
    .col_out_576             ( u5_col_out_576    ),
    .col_out_577             ( u5_col_out_577    ),
    .col_out_578             ( u5_col_out_578    ),
    .col_out_579             ( u5_col_out_579    ),
    .col_out_580             ( u5_col_out_580    ),
    .col_out_581             ( u5_col_out_581    ),
    .col_out_582             ( u5_col_out_582    ),
    .col_out_583             ( u5_col_out_583    ),
    .col_out_584             ( u5_col_out_584    ),
    .col_out_585             ( u5_col_out_585    ),
    .col_out_586             ( u5_col_out_586    ),
    .col_out_587             ( u5_col_out_587    ),
    .col_out_588             ( u5_col_out_588    ),
    .col_out_589             ( u5_col_out_589    ),
    .col_out_590             ( u5_col_out_590    ),
    .col_out_591             ( u5_col_out_591    ),
    .col_out_592             ( u5_col_out_592    ),
    .col_out_593             ( u5_col_out_593    ),
    .col_out_594             ( u5_col_out_594    ),
    .col_out_595             ( u5_col_out_595    ),
    .col_out_596             ( u5_col_out_596    ),
    .col_out_597             ( u5_col_out_597    ),
    .col_out_598             ( u5_col_out_598    ),
    .col_out_599             ( u5_col_out_599    ),
    .col_out_600             ( u5_col_out_600    ),
    .col_out_601             ( u5_col_out_601    ),
    .col_out_602             ( u5_col_out_602    ),
    .col_out_603             ( u5_col_out_603    ),
    .col_out_604             ( u5_col_out_604    ),
    .col_out_605             ( u5_col_out_605    ),
    .col_out_606             ( u5_col_out_606    ),
    .col_out_607             ( u5_col_out_607    ),
    .col_out_608             ( u5_col_out_608    ),
    .col_out_609             ( u5_col_out_609    ),
    .col_out_610             ( u5_col_out_610    ),
    .col_out_611             ( u5_col_out_611    ),
    .col_out_612             ( u5_col_out_612    ),
    .col_out_613             ( u5_col_out_613    ),
    .col_out_614             ( u5_col_out_614    ),
    .col_out_615             ( u5_col_out_615    ),
    .col_out_616             ( u5_col_out_616    ),
    .col_out_617             ( u5_col_out_617    ),
    .col_out_618             ( u5_col_out_618    ),
    .col_out_619             ( u5_col_out_619    ),
    .col_out_620             ( u5_col_out_620    ),
    .col_out_621             ( u5_col_out_621    ),
    .col_out_622             ( u5_col_out_622    ),
    .col_out_623             ( u5_col_out_623    ),
    .col_out_624             ( u5_col_out_624    ),
    .col_out_625             ( u5_col_out_625    ),
    .col_out_626             ( u5_col_out_626    ),
    .col_out_627             ( u5_col_out_627    ),
    .col_out_628             ( u5_col_out_628    ),
    .col_out_629             ( u5_col_out_629    ),
    .col_out_630             ( u5_col_out_630    ),
    .col_out_631             ( u5_col_out_631    ),
    .col_out_632             ( u5_col_out_632    ),
    .col_out_633             ( u5_col_out_633    ),
    .col_out_634             ( u5_col_out_634    ),
    .col_out_635             ( u5_col_out_635    ),
    .col_out_636             ( u5_col_out_636    ),
    .col_out_637             ( u5_col_out_637    ),
    .col_out_638             ( u5_col_out_638    ),
    .col_out_639             ( u5_col_out_639    ),
    .col_out_640             ( u5_col_out_640    ),
    .col_out_641             ( u5_col_out_641    ),
    .col_out_642             ( u5_col_out_642    ),
    .col_out_643             ( u5_col_out_643    ),
    .col_out_644             ( u5_col_out_644    ),
    .col_out_645             ( u5_col_out_645    ),
    .col_out_646             ( u5_col_out_646    ),
    .col_out_647             ( u5_col_out_647    ),
    .col_out_648             ( u5_col_out_648    ),
    .col_out_649             ( u5_col_out_649    ),
    .col_out_650             ( u5_col_out_650    ),
    .col_out_651             ( u5_col_out_651    ),
    .col_out_652             ( u5_col_out_652    ),
    .col_out_653             ( u5_col_out_653    ),
    .col_out_654             ( u5_col_out_654    ),
    .col_out_655             ( u5_col_out_655    ),
    .col_out_656             ( u5_col_out_656    ),
    .col_out_657             ( u5_col_out_657    ),
    .col_out_658             ( u5_col_out_658    ),
    .col_out_659             ( u5_col_out_659    ),
    .col_out_660             ( u5_col_out_660    ),
    .col_out_661             ( u5_col_out_661    ),
    .col_out_662             ( u5_col_out_662    ),
    .col_out_663             ( u5_col_out_663    ),
    .col_out_664             ( u5_col_out_664    ),
    .col_out_665             ( u5_col_out_665    ),
    .col_out_666             ( u5_col_out_666    ),
    .col_out_667             ( u5_col_out_667    ),
    .col_out_668             ( u5_col_out_668    ),
    .col_out_669             ( u5_col_out_669    ),
    .col_out_670             ( u5_col_out_670    ),
    .col_out_671             ( u5_col_out_671    ),
    .col_out_672             ( u5_col_out_672    ),
    .col_out_673             ( u5_col_out_673    ),
    .col_out_674             ( u5_col_out_674    ),
    .col_out_675             ( u5_col_out_675    ),
    .col_out_676             ( u5_col_out_676    ),
    .col_out_677             ( u5_col_out_677    ),
    .col_out_678             ( u5_col_out_678    ),
    .col_out_679             ( u5_col_out_679    ),
    .col_out_680             ( u5_col_out_680    ),
    .col_out_681             ( u5_col_out_681    ),
    .col_out_682             ( u5_col_out_682    ),
    .col_out_683             ( u5_col_out_683    ),
    .col_out_684             ( u5_col_out_684    ),
    .col_out_685             ( u5_col_out_685    ),
    .col_out_686             ( u5_col_out_686    ),
    .col_out_687             ( u5_col_out_687    ),
    .col_out_688             ( u5_col_out_688    ),
    .col_out_689             ( u5_col_out_689    ),
    .col_out_690             ( u5_col_out_690    ),
    .col_out_691             ( u5_col_out_691    ),
    .col_out_692             ( u5_col_out_692    ),
    .col_out_693             ( u5_col_out_693    ),
    .col_out_694             ( u5_col_out_694    ),
    .col_out_695             ( u5_col_out_695    ),
    .col_out_696             ( u5_col_out_696    ),
    .col_out_697             ( u5_col_out_697    ),
    .col_out_698             ( u5_col_out_698    ),
    .col_out_699             ( u5_col_out_699    ),
    .col_out_700             ( u5_col_out_700    ),
    .col_out_701             ( u5_col_out_701    ),
    .col_out_702             ( u5_col_out_702    ),
    .col_out_703             ( u5_col_out_703    ),
    .col_out_704             ( u5_col_out_704    ),
    .col_out_705             ( u5_col_out_705    ),
    .col_out_706             ( u5_col_out_706    ),
    .col_out_707             ( u5_col_out_707    ),
    .col_out_708             ( u5_col_out_708    ),
    .col_out_709             ( u5_col_out_709    ),
    .col_out_710             ( u5_col_out_710    ),
    .col_out_711             ( u5_col_out_711    ),
    .col_out_712             ( u5_col_out_712    ),
    .col_out_713             ( u5_col_out_713    ),
    .col_out_714             ( u5_col_out_714    ),
    .col_out_715             ( u5_col_out_715    ),
    .col_out_716             ( u5_col_out_716    ),
    .col_out_717             ( u5_col_out_717    ),
    .col_out_718             ( u5_col_out_718    ),
    .col_out_719             ( u5_col_out_719    ),
    .col_out_720             ( u5_col_out_720    ),
    .col_out_721             ( u5_col_out_721    ),
    .col_out_722             ( u5_col_out_722    ),
    .col_out_723             ( u5_col_out_723    ),
    .col_out_724             ( u5_col_out_724    ),
    .col_out_725             ( u5_col_out_725    ),
    .col_out_726             ( u5_col_out_726    ),
    .col_out_727             ( u5_col_out_727    ),
    .col_out_728             ( u5_col_out_728    ),
    .col_out_729             ( u5_col_out_729    ),
    .col_out_730             ( u5_col_out_730    ),
    .col_out_731             ( u5_col_out_731    ),
    .col_out_732             ( u5_col_out_732    ),
    .col_out_733             ( u5_col_out_733    ),
    .col_out_734             ( u5_col_out_734    ),
    .col_out_735             ( u5_col_out_735    ),
    .col_out_736             ( u5_col_out_736    ),
    .col_out_737             ( u5_col_out_737    ),
    .col_out_738             ( u5_col_out_738    ),
    .col_out_739             ( u5_col_out_739    ),
    .col_out_740             ( u5_col_out_740    ),
    .col_out_741             ( u5_col_out_741    ),
    .col_out_742             ( u5_col_out_742    ),
    .col_out_743             ( u5_col_out_743    ),
    .col_out_744             ( u5_col_out_744    ),
    .col_out_745             ( u5_col_out_745    ),
    .col_out_746             ( u5_col_out_746    ),
    .col_out_747             ( u5_col_out_747    ),
    .col_out_748             ( u5_col_out_748    ),
    .col_out_749             ( u5_col_out_749    ),
    .col_out_750             ( u5_col_out_750    ),
    .col_out_751             ( u5_col_out_751    ),
    .col_out_752             ( u5_col_out_752    ),
    .col_out_753             ( u5_col_out_753    ),
    .col_out_754             ( u5_col_out_754    ),
    .col_out_755             ( u5_col_out_755    ),
    .col_out_756             ( u5_col_out_756    ),
    .col_out_757             ( u5_col_out_757    ),
    .col_out_758             ( u5_col_out_758    ),
    .col_out_759             ( u5_col_out_759    ),
    .col_out_760             ( u5_col_out_760    ),
    .col_out_761             ( u5_col_out_761    ),
    .col_out_762             ( u5_col_out_762    ),
    .col_out_763             ( u5_col_out_763    ),
    .col_out_764             ( u5_col_out_764    ),
    .col_out_765             ( u5_col_out_765    ),
    .col_out_766             ( u5_col_out_766    ),
    .col_out_767             ( u5_col_out_767    ),
    .col_out_768             ( u5_col_out_768    ),
    .col_out_769             ( u5_col_out_769    ),
    .col_out_770             ( u5_col_out_770    ),
    .col_out_771             ( u5_col_out_771    ),
    .col_out_772             ( u5_col_out_772    ),
    .col_out_773             ( u5_col_out_773    ),
    .col_out_774             ( u5_col_out_774    ),
    .col_out_775             ( u5_col_out_775    ),
    .col_out_776             ( u5_col_out_776    ),
    .col_out_777             ( u5_col_out_777    ),
    .col_out_778             ( u5_col_out_778    ),
    .col_out_779             ( u5_col_out_779    ),
    .col_out_780             ( u5_col_out_780    ),
    .col_out_781             ( u5_col_out_781    ),
    .col_out_782             ( u5_col_out_782    ),
    .col_out_783             ( u5_col_out_783    ),
    .col_out_784             ( u5_col_out_784    ),
    .col_out_785             ( u5_col_out_785    ),
    .col_out_786             ( u5_col_out_786    ),
    .col_out_787             ( u5_col_out_787    ),
    .col_out_788             ( u5_col_out_788    ),
    .col_out_789             ( u5_col_out_789    ),
    .col_out_790             ( u5_col_out_790    ),
    .col_out_791             ( u5_col_out_791    ),
    .col_out_792             ( u5_col_out_792    ),
    .col_out_793             ( u5_col_out_793    ),
    .col_out_794             ( u5_col_out_794    ),
    .col_out_795             ( u5_col_out_795    ),
    .col_out_796             ( u5_col_out_796    ),
    .col_out_797             ( u5_col_out_797    ),
    .col_out_798             ( u5_col_out_798    ),
    .col_out_799             ( u5_col_out_799    ),
    .col_out_800             ( u5_col_out_800    ),
    .col_out_801             ( u5_col_out_801    ),
    .col_out_802             ( u5_col_out_802    ),
    .col_out_803             ( u5_col_out_803    ),
    .col_out_804             ( u5_col_out_804    ),
    .col_out_805             ( u5_col_out_805    ),
    .col_out_806             ( u5_col_out_806    ),
    .col_out_807             ( u5_col_out_807    ),
    .col_out_808             ( u5_col_out_808    ),
    .col_out_809             ( u5_col_out_809    ),
    .col_out_810             ( u5_col_out_810    ),
    .col_out_811             ( u5_col_out_811    ),
    .col_out_812             ( u5_col_out_812    ),
    .col_out_813             ( u5_col_out_813    ),
    .col_out_814             ( u5_col_out_814    ),
    .col_out_815             ( u5_col_out_815    ),
    .col_out_816             ( u5_col_out_816    ),
    .col_out_817             ( u5_col_out_817    ),
    .col_out_818             ( u5_col_out_818    ),
    .col_out_819             ( u5_col_out_819    ),
    .col_out_820             ( u5_col_out_820    ),
    .col_out_821             ( u5_col_out_821    ),
    .col_out_822             ( u5_col_out_822    ),
    .col_out_823             ( u5_col_out_823    ),
    .col_out_824             ( u5_col_out_824    ),
    .col_out_825             ( u5_col_out_825    ),
    .col_out_826             ( u5_col_out_826    ),
    .col_out_827             ( u5_col_out_827    ),
    .col_out_828             ( u5_col_out_828    ),
    .col_out_829             ( u5_col_out_829    ),
    .col_out_830             ( u5_col_out_830    ),
    .col_out_831             ( u5_col_out_831    ),
    .col_out_832             ( u5_col_out_832    ),
    .col_out_833             ( u5_col_out_833    ),
    .col_out_834             ( u5_col_out_834    ),
    .col_out_835             ( u5_col_out_835    ),
    .col_out_836             ( u5_col_out_836    ),
    .col_out_837             ( u5_col_out_837    ),
    .col_out_838             ( u5_col_out_838    ),
    .col_out_839             ( u5_col_out_839    ),
    .col_out_840             ( u5_col_out_840    ),
    .col_out_841             ( u5_col_out_841    ),
    .col_out_842             ( u5_col_out_842    ),
    .col_out_843             ( u5_col_out_843    ),
    .col_out_844             ( u5_col_out_844    ),
    .col_out_845             ( u5_col_out_845    ),
    .col_out_846             ( u5_col_out_846    ),
    .col_out_847             ( u5_col_out_847    ),
    .col_out_848             ( u5_col_out_848    ),
    .col_out_849             ( u5_col_out_849    ),
    .col_out_850             ( u5_col_out_850    ),
    .col_out_851             ( u5_col_out_851    ),
    .col_out_852             ( u5_col_out_852    ),
    .col_out_853             ( u5_col_out_853    ),
    .col_out_854             ( u5_col_out_854    ),
    .col_out_855             ( u5_col_out_855    ),
    .col_out_856             ( u5_col_out_856    ),
    .col_out_857             ( u5_col_out_857    ),
    .col_out_858             ( u5_col_out_858    ),
    .col_out_859             ( u5_col_out_859    ),
    .col_out_860             ( u5_col_out_860    ),
    .col_out_861             ( u5_col_out_861    ),
    .col_out_862             ( u5_col_out_862    ),
    .col_out_863             ( u5_col_out_863    ),
    .col_out_864             ( u5_col_out_864    ),
    .col_out_865             ( u5_col_out_865    ),
    .col_out_866             ( u5_col_out_866    ),
    .col_out_867             ( u5_col_out_867    ),
    .col_out_868             ( u5_col_out_868    ),
    .col_out_869             ( u5_col_out_869    ),
    .col_out_870             ( u5_col_out_870    ),
    .col_out_871             ( u5_col_out_871    ),
    .col_out_872             ( u5_col_out_872    ),
    .col_out_873             ( u5_col_out_873    ),
    .col_out_874             ( u5_col_out_874    ),
    .col_out_875             ( u5_col_out_875    ),
    .col_out_876             ( u5_col_out_876    ),
    .col_out_877             ( u5_col_out_877    ),
    .col_out_878             ( u5_col_out_878    ),
    .col_out_879             ( u5_col_out_879    ),
    .col_out_880             ( u5_col_out_880    ),
    .col_out_881             ( u5_col_out_881    ),
    .col_out_882             ( u5_col_out_882    ),
    .col_out_883             ( u5_col_out_883    ),
    .col_out_884             ( u5_col_out_884    ),
    .col_out_885             ( u5_col_out_885    ),
    .col_out_886             ( u5_col_out_886    ),
    .col_out_887             ( u5_col_out_887    ),
    .col_out_888             ( u5_col_out_888    ),
    .col_out_889             ( u5_col_out_889    ),
    .col_out_890             ( u5_col_out_890    ),
    .col_out_891             ( u5_col_out_891    ),
    .col_out_892             ( u5_col_out_892    ),
    .col_out_893             ( u5_col_out_893    ),
    .col_out_894             ( u5_col_out_894    ),
    .col_out_895             ( u5_col_out_895    ),
    .col_out_896             ( u5_col_out_896    ),
    .col_out_897             ( u5_col_out_897    ),
    .col_out_898             ( u5_col_out_898    ),
    .col_out_899             ( u5_col_out_899    ),
    .col_out_900             ( u5_col_out_900    ),
    .col_out_901             ( u5_col_out_901    ),
    .col_out_902             ( u5_col_out_902    ),
    .col_out_903             ( u5_col_out_903    ),
    .col_out_904             ( u5_col_out_904    ),
    .col_out_905             ( u5_col_out_905    ),
    .col_out_906             ( u5_col_out_906    ),
    .col_out_907             ( u5_col_out_907    ),
    .col_out_908             ( u5_col_out_908    ),
    .col_out_909             ( u5_col_out_909    ),
    .col_out_910             ( u5_col_out_910    ),
    .col_out_911             ( u5_col_out_911    ),
    .col_out_912             ( u5_col_out_912    ),
    .col_out_913             ( u5_col_out_913    ),
    .col_out_914             ( u5_col_out_914    ),
    .col_out_915             ( u5_col_out_915    ),
    .col_out_916             ( u5_col_out_916    ),
    .col_out_917             ( u5_col_out_917    ),
    .col_out_918             ( u5_col_out_918    ),
    .col_out_919             ( u5_col_out_919    ),
    .col_out_920             ( u5_col_out_920    ),
    .col_out_921             ( u5_col_out_921    ),
    .col_out_922             ( u5_col_out_922    ),
    .col_out_923             ( u5_col_out_923    ),
    .col_out_924             ( u5_col_out_924    ),
    .col_out_925             ( u5_col_out_925    ),
    .col_out_926             ( u5_col_out_926    ),
    .col_out_927             ( u5_col_out_927    ),
    .col_out_928             ( u5_col_out_928    ),
    .col_out_929             ( u5_col_out_929    ),
    .col_out_930             ( u5_col_out_930    ),
    .col_out_931             ( u5_col_out_931    ),
    .col_out_932             ( u5_col_out_932    ),
    .col_out_933             ( u5_col_out_933    ),
    .col_out_934             ( u5_col_out_934    ),
    .col_out_935             ( u5_col_out_935    ),
    .col_out_936             ( u5_col_out_936    ),
    .col_out_937             ( u5_col_out_937    ),
    .col_out_938             ( u5_col_out_938    ),
    .col_out_939             ( u5_col_out_939    ),
    .col_out_940             ( u5_col_out_940    ),
    .col_out_941             ( u5_col_out_941    ),
    .col_out_942             ( u5_col_out_942    ),
    .col_out_943             ( u5_col_out_943    ),
    .col_out_944             ( u5_col_out_944    ),
    .col_out_945             ( u5_col_out_945    ),
    .col_out_946             ( u5_col_out_946    ),
    .col_out_947             ( u5_col_out_947    ),
    .col_out_948             ( u5_col_out_948    ),
    .col_out_949             ( u5_col_out_949    ),
    .col_out_950             ( u5_col_out_950    ),
    .col_out_951             ( u5_col_out_951    ),
    .col_out_952             ( u5_col_out_952    ),
    .col_out_953             ( u5_col_out_953    ),
    .col_out_954             ( u5_col_out_954    ),
    .col_out_955             ( u5_col_out_955    ),
    .col_out_956             ( u5_col_out_956    ),
    .col_out_957             ( u5_col_out_957    ),
    .col_out_958             ( u5_col_out_958    ),
    .col_out_959             ( u5_col_out_959    ),
    .col_out_960             ( u5_col_out_960    ),
    .col_out_961             ( u5_col_out_961    ),
    .col_out_962             ( u5_col_out_962    ),
    .col_out_963             ( u5_col_out_963    ),
    .col_out_964             ( u5_col_out_964    ),
    .col_out_965             ( u5_col_out_965    ),
    .col_out_966             ( u5_col_out_966    ),
    .col_out_967             ( u5_col_out_967    ),
    .col_out_968             ( u5_col_out_968    ),
    .col_out_969             ( u5_col_out_969    ),
    .col_out_970             ( u5_col_out_970    ),
    .col_out_971             ( u5_col_out_971    ),
    .col_out_972             ( u5_col_out_972    ),
    .col_out_973             ( u5_col_out_973    ),
    .col_out_974             ( u5_col_out_974    ),
    .col_out_975             ( u5_col_out_975    ),
    .col_out_976             ( u5_col_out_976    ),
    .col_out_977             ( u5_col_out_977    ),
    .col_out_978             ( u5_col_out_978    ),
    .col_out_979             ( u5_col_out_979    ),
    .col_out_980             ( u5_col_out_980    ),
    .col_out_981             ( u5_col_out_981    ),
    .col_out_982             ( u5_col_out_982    ),
    .col_out_983             ( u5_col_out_983    ),
    .col_out_984             ( u5_col_out_984    ),
    .col_out_985             ( u5_col_out_985    ),
    .col_out_986             ( u5_col_out_986    ),
    .col_out_987             ( u5_col_out_987    ),
    .col_out_988             ( u5_col_out_988    ),
    .col_out_989             ( u5_col_out_989    ),
    .col_out_990             ( u5_col_out_990    ),
    .col_out_991             ( u5_col_out_991    ),
    .col_out_992             ( u5_col_out_992    ),
    .col_out_993             ( u5_col_out_993    ),
    .col_out_994             ( u5_col_out_994    ),
    .col_out_995             ( u5_col_out_995    ),
    .col_out_996             ( u5_col_out_996    ),
    .col_out_997             ( u5_col_out_997    ),
    .col_out_998             ( u5_col_out_998    ),
    .col_out_999             ( u5_col_out_999    ),
    .col_out_1000            ( u5_col_out_1000   ),
    .col_out_1001            ( u5_col_out_1001   ),
    .col_out_1002            ( u5_col_out_1002   ),
    .col_out_1003            ( u5_col_out_1003   ),
    .col_out_1004            ( u5_col_out_1004   ),
    .col_out_1005            ( u5_col_out_1005   ),
    .col_out_1006            ( u5_col_out_1006   ),
    .col_out_1007            ( u5_col_out_1007   ),
    .col_out_1008            ( u5_col_out_1008   ),
    .col_out_1009            ( u5_col_out_1009   ),
    .col_out_1010            ( u5_col_out_1010   ),
    .col_out_1011            ( u5_col_out_1011   ),
    .col_out_1012            ( u5_col_out_1012   ),
    .col_out_1013            ( u5_col_out_1013   ),
    .col_out_1014            ( u5_col_out_1014   ),
    .col_out_1015            ( u5_col_out_1015   ),
    .col_out_1016            ( u5_col_out_1016   ),
    .col_out_1017            ( u5_col_out_1017   ),
    .col_out_1018            ( u5_col_out_1018   ),
    .col_out_1019            ( u5_col_out_1019   ),
    .col_out_1020            ( u5_col_out_1020   ),
    .col_out_1021            ( u5_col_out_1021   ),
    .col_out_1022            ( u5_col_out_1022   ),
    .col_out_1023            ( u5_col_out_1023   ),
    .col_out_1024            ( u5_col_out_1024   ),
    .col_out_1025            ( u5_col_out_1025   ),
    .col_out_1026            ( u5_col_out_1026   ),
    .col_out_1027            ( u5_col_out_1027   ),
    .col_out_1028            ( u5_col_out_1028   ),
    .col_out_1029            ( u5_col_out_1029   ),
    .col_out_1030            ( u5_col_out_1030   ),
    .col_out_1031            ( u5_col_out_1031   ),
    .col_out_1032            ( u5_col_out_1032   ),
    .col_out_1033            ( u5_col_out_1033   )
);






//*****************************************************
//**************输出赋值******************************
//*****************************************************
assign col_out_0 = u5_col_out_0;
assign col_out_1 = u5_col_out_1;
assign col_out_2 = u5_col_out_2;
assign col_out_3 = u5_col_out_3;
assign col_out_4 = u5_col_out_4;
assign col_out_5 = u5_col_out_5;
assign col_out_6 = u5_col_out_6;
assign col_out_7 = u5_col_out_7;
assign col_out_8 = u5_col_out_8;
assign col_out_9 = u5_col_out_9;
assign col_out_10 = u5_col_out_10;
assign col_out_11 = u5_col_out_11;
assign col_out_12 = u5_col_out_12;
assign col_out_13 = u5_col_out_13;
assign col_out_14 = u5_col_out_14;
assign col_out_15 = u5_col_out_15;
assign col_out_16 = u5_col_out_16;
assign col_out_17 = u5_col_out_17;
assign col_out_18 = u5_col_out_18;
assign col_out_19 = u5_col_out_19;
assign col_out_20 = u5_col_out_20;
assign col_out_21 = u5_col_out_21;
assign col_out_22 = u5_col_out_22;
assign col_out_23 = u5_col_out_23;
assign col_out_24 = u5_col_out_24;
assign col_out_25 = u5_col_out_25;
assign col_out_26 = u5_col_out_26;
assign col_out_27 = u5_col_out_27;
assign col_out_28 = u5_col_out_28;
assign col_out_29 = u5_col_out_29;
assign col_out_30 = u5_col_out_30;
assign col_out_31 = u5_col_out_31;
assign col_out_32 = u5_col_out_32;
assign col_out_33 = u5_col_out_33;
assign col_out_34 = u5_col_out_34;
assign col_out_35 = u5_col_out_35;
assign col_out_36 = u5_col_out_36;
assign col_out_37 = u5_col_out_37;
assign col_out_38 = u5_col_out_38;
assign col_out_39 = u5_col_out_39;
assign col_out_40 = u5_col_out_40;
assign col_out_41 = u5_col_out_41;
assign col_out_42 = u5_col_out_42;
assign col_out_43 = u5_col_out_43;
assign col_out_44 = u5_col_out_44;
assign col_out_45 = u5_col_out_45;
assign col_out_46 = u5_col_out_46;
assign col_out_47 = u5_col_out_47;
assign col_out_48 = u5_col_out_48;
assign col_out_49 = u5_col_out_49;
assign col_out_50 = u5_col_out_50;
assign col_out_51 = u5_col_out_51;
assign col_out_52 = u5_col_out_52;
assign col_out_53 = u5_col_out_53;
assign col_out_54 = u5_col_out_54;
assign col_out_55 = u5_col_out_55;
assign col_out_56 = u5_col_out_56;
assign col_out_57 = u5_col_out_57;
assign col_out_58 = u5_col_out_58;
assign col_out_59 = u5_col_out_59;
assign col_out_60 = u5_col_out_60;
assign col_out_61 = u5_col_out_61;
assign col_out_62 = u5_col_out_62;
assign col_out_63 = u5_col_out_63;
assign col_out_64 = u5_col_out_64;
assign col_out_65 = u5_col_out_65;
assign col_out_66 = u5_col_out_66;
assign col_out_67 = u5_col_out_67;
assign col_out_68 = u5_col_out_68;
assign col_out_69 = u5_col_out_69;
assign col_out_70 = u5_col_out_70;
assign col_out_71 = u5_col_out_71;
assign col_out_72 = u5_col_out_72;
assign col_out_73 = u5_col_out_73;
assign col_out_74 = u5_col_out_74;
assign col_out_75 = u5_col_out_75;
assign col_out_76 = u5_col_out_76;
assign col_out_77 = u5_col_out_77;
assign col_out_78 = u5_col_out_78;
assign col_out_79 = u5_col_out_79;
assign col_out_80 = u5_col_out_80;
assign col_out_81 = u5_col_out_81;
assign col_out_82 = u5_col_out_82;
assign col_out_83 = u5_col_out_83;
assign col_out_84 = u5_col_out_84;
assign col_out_85 = u5_col_out_85;
assign col_out_86 = u5_col_out_86;
assign col_out_87 = u5_col_out_87;
assign col_out_88 = u5_col_out_88;
assign col_out_89 = u5_col_out_89;
assign col_out_90 = u5_col_out_90;
assign col_out_91 = u5_col_out_91;
assign col_out_92 = u5_col_out_92;
assign col_out_93 = u5_col_out_93;
assign col_out_94 = u5_col_out_94;
assign col_out_95 = u5_col_out_95;
assign col_out_96 = u5_col_out_96;
assign col_out_97 = u5_col_out_97;
assign col_out_98 = u5_col_out_98;
assign col_out_99 = u5_col_out_99;
assign col_out_100 = u5_col_out_100;
assign col_out_101 = u5_col_out_101;
assign col_out_102 = u5_col_out_102;
assign col_out_103 = u5_col_out_103;
assign col_out_104 = u5_col_out_104;
assign col_out_105 = u5_col_out_105;
assign col_out_106 = u5_col_out_106;
assign col_out_107 = u5_col_out_107;
assign col_out_108 = u5_col_out_108;
assign col_out_109 = u5_col_out_109;
assign col_out_110 = u5_col_out_110;
assign col_out_111 = u5_col_out_111;
assign col_out_112 = u5_col_out_112;
assign col_out_113 = u5_col_out_113;
assign col_out_114 = u5_col_out_114;
assign col_out_115 = u5_col_out_115;
assign col_out_116 = u5_col_out_116;
assign col_out_117 = u5_col_out_117;
assign col_out_118 = u5_col_out_118;
assign col_out_119 = u5_col_out_119;
assign col_out_120 = u5_col_out_120;
assign col_out_121 = u5_col_out_121;
assign col_out_122 = u5_col_out_122;
assign col_out_123 = u5_col_out_123;
assign col_out_124 = u5_col_out_124;
assign col_out_125 = u5_col_out_125;
assign col_out_126 = u5_col_out_126;
assign col_out_127 = u5_col_out_127;
assign col_out_128 = u5_col_out_128;
assign col_out_129 = u5_col_out_129;
assign col_out_130 = u5_col_out_130;
assign col_out_131 = u5_col_out_131;
assign col_out_132 = u5_col_out_132;
assign col_out_133 = u5_col_out_133;
assign col_out_134 = u5_col_out_134;
assign col_out_135 = u5_col_out_135;
assign col_out_136 = u5_col_out_136;
assign col_out_137 = u5_col_out_137;
assign col_out_138 = u5_col_out_138;
assign col_out_139 = u5_col_out_139;
assign col_out_140 = u5_col_out_140;
assign col_out_141 = u5_col_out_141;
assign col_out_142 = u5_col_out_142;
assign col_out_143 = u5_col_out_143;
assign col_out_144 = u5_col_out_144;
assign col_out_145 = u5_col_out_145;
assign col_out_146 = u5_col_out_146;
assign col_out_147 = u5_col_out_147;
assign col_out_148 = u5_col_out_148;
assign col_out_149 = u5_col_out_149;
assign col_out_150 = u5_col_out_150;
assign col_out_151 = u5_col_out_151;
assign col_out_152 = u5_col_out_152;
assign col_out_153 = u5_col_out_153;
assign col_out_154 = u5_col_out_154;
assign col_out_155 = u5_col_out_155;
assign col_out_156 = u5_col_out_156;
assign col_out_157 = u5_col_out_157;
assign col_out_158 = u5_col_out_158;
assign col_out_159 = u5_col_out_159;
assign col_out_160 = u5_col_out_160;
assign col_out_161 = u5_col_out_161;
assign col_out_162 = u5_col_out_162;
assign col_out_163 = u5_col_out_163;
assign col_out_164 = u5_col_out_164;
assign col_out_165 = u5_col_out_165;
assign col_out_166 = u5_col_out_166;
assign col_out_167 = u5_col_out_167;
assign col_out_168 = u5_col_out_168;
assign col_out_169 = u5_col_out_169;
assign col_out_170 = u5_col_out_170;
assign col_out_171 = u5_col_out_171;
assign col_out_172 = u5_col_out_172;
assign col_out_173 = u5_col_out_173;
assign col_out_174 = u5_col_out_174;
assign col_out_175 = u5_col_out_175;
assign col_out_176 = u5_col_out_176;
assign col_out_177 = u5_col_out_177;
assign col_out_178 = u5_col_out_178;
assign col_out_179 = u5_col_out_179;
assign col_out_180 = u5_col_out_180;
assign col_out_181 = u5_col_out_181;
assign col_out_182 = u5_col_out_182;
assign col_out_183 = u5_col_out_183;
assign col_out_184 = u5_col_out_184;
assign col_out_185 = u5_col_out_185;
assign col_out_186 = u5_col_out_186;
assign col_out_187 = u5_col_out_187;
assign col_out_188 = u5_col_out_188;
assign col_out_189 = u5_col_out_189;
assign col_out_190 = u5_col_out_190;
assign col_out_191 = u5_col_out_191;
assign col_out_192 = u5_col_out_192;
assign col_out_193 = u5_col_out_193;
assign col_out_194 = u5_col_out_194;
assign col_out_195 = u5_col_out_195;
assign col_out_196 = u5_col_out_196;
assign col_out_197 = u5_col_out_197;
assign col_out_198 = u5_col_out_198;
assign col_out_199 = u5_col_out_199;
assign col_out_200 = u5_col_out_200;
assign col_out_201 = u5_col_out_201;
assign col_out_202 = u5_col_out_202;
assign col_out_203 = u5_col_out_203;
assign col_out_204 = u5_col_out_204;
assign col_out_205 = u5_col_out_205;
assign col_out_206 = u5_col_out_206;
assign col_out_207 = u5_col_out_207;
assign col_out_208 = u5_col_out_208;
assign col_out_209 = u5_col_out_209;
assign col_out_210 = u5_col_out_210;
assign col_out_211 = u5_col_out_211;
assign col_out_212 = u5_col_out_212;
assign col_out_213 = u5_col_out_213;
assign col_out_214 = u5_col_out_214;
assign col_out_215 = u5_col_out_215;
assign col_out_216 = u5_col_out_216;
assign col_out_217 = u5_col_out_217;
assign col_out_218 = u5_col_out_218;
assign col_out_219 = u5_col_out_219;
assign col_out_220 = u5_col_out_220;
assign col_out_221 = u5_col_out_221;
assign col_out_222 = u5_col_out_222;
assign col_out_223 = u5_col_out_223;
assign col_out_224 = u5_col_out_224;
assign col_out_225 = u5_col_out_225;
assign col_out_226 = u5_col_out_226;
assign col_out_227 = u5_col_out_227;
assign col_out_228 = u5_col_out_228;
assign col_out_229 = u5_col_out_229;
assign col_out_230 = u5_col_out_230;
assign col_out_231 = u5_col_out_231;
assign col_out_232 = u5_col_out_232;
assign col_out_233 = u5_col_out_233;
assign col_out_234 = u5_col_out_234;
assign col_out_235 = u5_col_out_235;
assign col_out_236 = u5_col_out_236;
assign col_out_237 = u5_col_out_237;
assign col_out_238 = u5_col_out_238;
assign col_out_239 = u5_col_out_239;
assign col_out_240 = u5_col_out_240;
assign col_out_241 = u5_col_out_241;
assign col_out_242 = u5_col_out_242;
assign col_out_243 = u5_col_out_243;
assign col_out_244 = u5_col_out_244;
assign col_out_245 = u5_col_out_245;
assign col_out_246 = u5_col_out_246;
assign col_out_247 = u5_col_out_247;
assign col_out_248 = u5_col_out_248;
assign col_out_249 = u5_col_out_249;
assign col_out_250 = u5_col_out_250;
assign col_out_251 = u5_col_out_251;
assign col_out_252 = u5_col_out_252;
assign col_out_253 = u5_col_out_253;
assign col_out_254 = u5_col_out_254;
assign col_out_255 = u5_col_out_255;
assign col_out_256 = u5_col_out_256;
assign col_out_257 = u5_col_out_257;
assign col_out_258 = u5_col_out_258;
assign col_out_259 = u5_col_out_259;
assign col_out_260 = u5_col_out_260;
assign col_out_261 = u5_col_out_261;
assign col_out_262 = u5_col_out_262;
assign col_out_263 = u5_col_out_263;
assign col_out_264 = u5_col_out_264;
assign col_out_265 = u5_col_out_265;
assign col_out_266 = u5_col_out_266;
assign col_out_267 = u5_col_out_267;
assign col_out_268 = u5_col_out_268;
assign col_out_269 = u5_col_out_269;
assign col_out_270 = u5_col_out_270;
assign col_out_271 = u5_col_out_271;
assign col_out_272 = u5_col_out_272;
assign col_out_273 = u5_col_out_273;
assign col_out_274 = u5_col_out_274;
assign col_out_275 = u5_col_out_275;
assign col_out_276 = u5_col_out_276;
assign col_out_277 = u5_col_out_277;
assign col_out_278 = u5_col_out_278;
assign col_out_279 = u5_col_out_279;
assign col_out_280 = u5_col_out_280;
assign col_out_281 = u5_col_out_281;
assign col_out_282 = u5_col_out_282;
assign col_out_283 = u5_col_out_283;
assign col_out_284 = u5_col_out_284;
assign col_out_285 = u5_col_out_285;
assign col_out_286 = u5_col_out_286;
assign col_out_287 = u5_col_out_287;
assign col_out_288 = u5_col_out_288;
assign col_out_289 = u5_col_out_289;
assign col_out_290 = u5_col_out_290;
assign col_out_291 = u5_col_out_291;
assign col_out_292 = u5_col_out_292;
assign col_out_293 = u5_col_out_293;
assign col_out_294 = u5_col_out_294;
assign col_out_295 = u5_col_out_295;
assign col_out_296 = u5_col_out_296;
assign col_out_297 = u5_col_out_297;
assign col_out_298 = u5_col_out_298;
assign col_out_299 = u5_col_out_299;
assign col_out_300 = u5_col_out_300;
assign col_out_301 = u5_col_out_301;
assign col_out_302 = u5_col_out_302;
assign col_out_303 = u5_col_out_303;
assign col_out_304 = u5_col_out_304;
assign col_out_305 = u5_col_out_305;
assign col_out_306 = u5_col_out_306;
assign col_out_307 = u5_col_out_307;
assign col_out_308 = u5_col_out_308;
assign col_out_309 = u5_col_out_309;
assign col_out_310 = u5_col_out_310;
assign col_out_311 = u5_col_out_311;
assign col_out_312 = u5_col_out_312;
assign col_out_313 = u5_col_out_313;
assign col_out_314 = u5_col_out_314;
assign col_out_315 = u5_col_out_315;
assign col_out_316 = u5_col_out_316;
assign col_out_317 = u5_col_out_317;
assign col_out_318 = u5_col_out_318;
assign col_out_319 = u5_col_out_319;
assign col_out_320 = u5_col_out_320;
assign col_out_321 = u5_col_out_321;
assign col_out_322 = u5_col_out_322;
assign col_out_323 = u5_col_out_323;
assign col_out_324 = u5_col_out_324;
assign col_out_325 = u5_col_out_325;
assign col_out_326 = u5_col_out_326;
assign col_out_327 = u5_col_out_327;
assign col_out_328 = u5_col_out_328;
assign col_out_329 = u5_col_out_329;
assign col_out_330 = u5_col_out_330;
assign col_out_331 = u5_col_out_331;
assign col_out_332 = u5_col_out_332;
assign col_out_333 = u5_col_out_333;
assign col_out_334 = u5_col_out_334;
assign col_out_335 = u5_col_out_335;
assign col_out_336 = u5_col_out_336;
assign col_out_337 = u5_col_out_337;
assign col_out_338 = u5_col_out_338;
assign col_out_339 = u5_col_out_339;
assign col_out_340 = u5_col_out_340;
assign col_out_341 = u5_col_out_341;
assign col_out_342 = u5_col_out_342;
assign col_out_343 = u5_col_out_343;
assign col_out_344 = u5_col_out_344;
assign col_out_345 = u5_col_out_345;
assign col_out_346 = u5_col_out_346;
assign col_out_347 = u5_col_out_347;
assign col_out_348 = u5_col_out_348;
assign col_out_349 = u5_col_out_349;
assign col_out_350 = u5_col_out_350;
assign col_out_351 = u5_col_out_351;
assign col_out_352 = u5_col_out_352;
assign col_out_353 = u5_col_out_353;
assign col_out_354 = u5_col_out_354;
assign col_out_355 = u5_col_out_355;
assign col_out_356 = u5_col_out_356;
assign col_out_357 = u5_col_out_357;
assign col_out_358 = u5_col_out_358;
assign col_out_359 = u5_col_out_359;
assign col_out_360 = u5_col_out_360;
assign col_out_361 = u5_col_out_361;
assign col_out_362 = u5_col_out_362;
assign col_out_363 = u5_col_out_363;
assign col_out_364 = u5_col_out_364;
assign col_out_365 = u5_col_out_365;
assign col_out_366 = u5_col_out_366;
assign col_out_367 = u5_col_out_367;
assign col_out_368 = u5_col_out_368;
assign col_out_369 = u5_col_out_369;
assign col_out_370 = u5_col_out_370;
assign col_out_371 = u5_col_out_371;
assign col_out_372 = u5_col_out_372;
assign col_out_373 = u5_col_out_373;
assign col_out_374 = u5_col_out_374;
assign col_out_375 = u5_col_out_375;
assign col_out_376 = u5_col_out_376;
assign col_out_377 = u5_col_out_377;
assign col_out_378 = u5_col_out_378;
assign col_out_379 = u5_col_out_379;
assign col_out_380 = u5_col_out_380;
assign col_out_381 = u5_col_out_381;
assign col_out_382 = u5_col_out_382;
assign col_out_383 = u5_col_out_383;
assign col_out_384 = u5_col_out_384;
assign col_out_385 = u5_col_out_385;
assign col_out_386 = u5_col_out_386;
assign col_out_387 = u5_col_out_387;
assign col_out_388 = u5_col_out_388;
assign col_out_389 = u5_col_out_389;
assign col_out_390 = u5_col_out_390;
assign col_out_391 = u5_col_out_391;
assign col_out_392 = u5_col_out_392;
assign col_out_393 = u5_col_out_393;
assign col_out_394 = u5_col_out_394;
assign col_out_395 = u5_col_out_395;
assign col_out_396 = u5_col_out_396;
assign col_out_397 = u5_col_out_397;
assign col_out_398 = u5_col_out_398;
assign col_out_399 = u5_col_out_399;
assign col_out_400 = u5_col_out_400;
assign col_out_401 = u5_col_out_401;
assign col_out_402 = u5_col_out_402;
assign col_out_403 = u5_col_out_403;
assign col_out_404 = u5_col_out_404;
assign col_out_405 = u5_col_out_405;
assign col_out_406 = u5_col_out_406;
assign col_out_407 = u5_col_out_407;
assign col_out_408 = u5_col_out_408;
assign col_out_409 = u5_col_out_409;
assign col_out_410 = u5_col_out_410;
assign col_out_411 = u5_col_out_411;
assign col_out_412 = u5_col_out_412;
assign col_out_413 = u5_col_out_413;
assign col_out_414 = u5_col_out_414;
assign col_out_415 = u5_col_out_415;
assign col_out_416 = u5_col_out_416;
assign col_out_417 = u5_col_out_417;
assign col_out_418 = u5_col_out_418;
assign col_out_419 = u5_col_out_419;
assign col_out_420 = u5_col_out_420;
assign col_out_421 = u5_col_out_421;
assign col_out_422 = u5_col_out_422;
assign col_out_423 = u5_col_out_423;
assign col_out_424 = u5_col_out_424;
assign col_out_425 = u5_col_out_425;
assign col_out_426 = u5_col_out_426;
assign col_out_427 = u5_col_out_427;
assign col_out_428 = u5_col_out_428;
assign col_out_429 = u5_col_out_429;
assign col_out_430 = u5_col_out_430;
assign col_out_431 = u5_col_out_431;
assign col_out_432 = u5_col_out_432;
assign col_out_433 = u5_col_out_433;
assign col_out_434 = u5_col_out_434;
assign col_out_435 = u5_col_out_435;
assign col_out_436 = u5_col_out_436;
assign col_out_437 = u5_col_out_437;
assign col_out_438 = u5_col_out_438;
assign col_out_439 = u5_col_out_439;
assign col_out_440 = u5_col_out_440;
assign col_out_441 = u5_col_out_441;
assign col_out_442 = u5_col_out_442;
assign col_out_443 = u5_col_out_443;
assign col_out_444 = u5_col_out_444;
assign col_out_445 = u5_col_out_445;
assign col_out_446 = u5_col_out_446;
assign col_out_447 = u5_col_out_447;
assign col_out_448 = u5_col_out_448;
assign col_out_449 = u5_col_out_449;
assign col_out_450 = u5_col_out_450;
assign col_out_451 = u5_col_out_451;
assign col_out_452 = u5_col_out_452;
assign col_out_453 = u5_col_out_453;
assign col_out_454 = u5_col_out_454;
assign col_out_455 = u5_col_out_455;
assign col_out_456 = u5_col_out_456;
assign col_out_457 = u5_col_out_457;
assign col_out_458 = u5_col_out_458;
assign col_out_459 = u5_col_out_459;
assign col_out_460 = u5_col_out_460;
assign col_out_461 = u5_col_out_461;
assign col_out_462 = u5_col_out_462;
assign col_out_463 = u5_col_out_463;
assign col_out_464 = u5_col_out_464;
assign col_out_465 = u5_col_out_465;
assign col_out_466 = u5_col_out_466;
assign col_out_467 = u5_col_out_467;
assign col_out_468 = u5_col_out_468;
assign col_out_469 = u5_col_out_469;
assign col_out_470 = u5_col_out_470;
assign col_out_471 = u5_col_out_471;
assign col_out_472 = u5_col_out_472;
assign col_out_473 = u5_col_out_473;
assign col_out_474 = u5_col_out_474;
assign col_out_475 = u5_col_out_475;
assign col_out_476 = u5_col_out_476;
assign col_out_477 = u5_col_out_477;
assign col_out_478 = u5_col_out_478;
assign col_out_479 = u5_col_out_479;
assign col_out_480 = u5_col_out_480;
assign col_out_481 = u5_col_out_481;
assign col_out_482 = u5_col_out_482;
assign col_out_483 = u5_col_out_483;
assign col_out_484 = u5_col_out_484;
assign col_out_485 = u5_col_out_485;
assign col_out_486 = u5_col_out_486;
assign col_out_487 = u5_col_out_487;
assign col_out_488 = u5_col_out_488;
assign col_out_489 = u5_col_out_489;
assign col_out_490 = u5_col_out_490;
assign col_out_491 = u5_col_out_491;
assign col_out_492 = u5_col_out_492;
assign col_out_493 = u5_col_out_493;
assign col_out_494 = u5_col_out_494;
assign col_out_495 = u5_col_out_495;
assign col_out_496 = u5_col_out_496;
assign col_out_497 = u5_col_out_497;
assign col_out_498 = u5_col_out_498;
assign col_out_499 = u5_col_out_499;
assign col_out_500 = u5_col_out_500;
assign col_out_501 = u5_col_out_501;
assign col_out_502 = u5_col_out_502;
assign col_out_503 = u5_col_out_503;
assign col_out_504 = u5_col_out_504;
assign col_out_505 = u5_col_out_505;
assign col_out_506 = u5_col_out_506;
assign col_out_507 = u5_col_out_507;
assign col_out_508 = u5_col_out_508;
assign col_out_509 = u5_col_out_509;
assign col_out_510 = u5_col_out_510;
assign col_out_511 = u5_col_out_511;
assign col_out_512 = u5_col_out_512;
assign col_out_513 = u5_col_out_513;
assign col_out_514 = u5_col_out_514;
assign col_out_515 = u5_col_out_515;
assign col_out_516 = u5_col_out_516;
assign col_out_517 = u5_col_out_517;
assign col_out_518 = u5_col_out_518;
assign col_out_519 = u5_col_out_519;
assign col_out_520 = u5_col_out_520;
assign col_out_521 = u5_col_out_521;
assign col_out_522 = u5_col_out_522;
assign col_out_523 = u5_col_out_523;
assign col_out_524 = u5_col_out_524;
assign col_out_525 = u5_col_out_525;
assign col_out_526 = u5_col_out_526;
assign col_out_527 = u5_col_out_527;
assign col_out_528 = u5_col_out_528;
assign col_out_529 = u5_col_out_529;
assign col_out_530 = u5_col_out_530;
assign col_out_531 = u5_col_out_531;
assign col_out_532 = u5_col_out_532;
assign col_out_533 = u5_col_out_533;
assign col_out_534 = u5_col_out_534;
assign col_out_535 = u5_col_out_535;
assign col_out_536 = u5_col_out_536;
assign col_out_537 = u5_col_out_537;
assign col_out_538 = u5_col_out_538;
assign col_out_539 = u5_col_out_539;
assign col_out_540 = u5_col_out_540;
assign col_out_541 = u5_col_out_541;
assign col_out_542 = u5_col_out_542;
assign col_out_543 = u5_col_out_543;
assign col_out_544 = u5_col_out_544;
assign col_out_545 = u5_col_out_545;
assign col_out_546 = u5_col_out_546;
assign col_out_547 = u5_col_out_547;
assign col_out_548 = u5_col_out_548;
assign col_out_549 = u5_col_out_549;
assign col_out_550 = u5_col_out_550;
assign col_out_551 = u5_col_out_551;
assign col_out_552 = u5_col_out_552;
assign col_out_553 = u5_col_out_553;
assign col_out_554 = u5_col_out_554;
assign col_out_555 = u5_col_out_555;
assign col_out_556 = u5_col_out_556;
assign col_out_557 = u5_col_out_557;
assign col_out_558 = u5_col_out_558;
assign col_out_559 = u5_col_out_559;
assign col_out_560 = u5_col_out_560;
assign col_out_561 = u5_col_out_561;
assign col_out_562 = u5_col_out_562;
assign col_out_563 = u5_col_out_563;
assign col_out_564 = u5_col_out_564;
assign col_out_565 = u5_col_out_565;
assign col_out_566 = u5_col_out_566;
assign col_out_567 = u5_col_out_567;
assign col_out_568 = u5_col_out_568;
assign col_out_569 = u5_col_out_569;
assign col_out_570 = u5_col_out_570;
assign col_out_571 = u5_col_out_571;
assign col_out_572 = u5_col_out_572;
assign col_out_573 = u5_col_out_573;
assign col_out_574 = u5_col_out_574;
assign col_out_575 = u5_col_out_575;
assign col_out_576 = u5_col_out_576;
assign col_out_577 = u5_col_out_577;
assign col_out_578 = u5_col_out_578;
assign col_out_579 = u5_col_out_579;
assign col_out_580 = u5_col_out_580;
assign col_out_581 = u5_col_out_581;
assign col_out_582 = u5_col_out_582;
assign col_out_583 = u5_col_out_583;
assign col_out_584 = u5_col_out_584;
assign col_out_585 = u5_col_out_585;
assign col_out_586 = u5_col_out_586;
assign col_out_587 = u5_col_out_587;
assign col_out_588 = u5_col_out_588;
assign col_out_589 = u5_col_out_589;
assign col_out_590 = u5_col_out_590;
assign col_out_591 = u5_col_out_591;
assign col_out_592 = u5_col_out_592;
assign col_out_593 = u5_col_out_593;
assign col_out_594 = u5_col_out_594;
assign col_out_595 = u5_col_out_595;
assign col_out_596 = u5_col_out_596;
assign col_out_597 = u5_col_out_597;
assign col_out_598 = u5_col_out_598;
assign col_out_599 = u5_col_out_599;
assign col_out_600 = u5_col_out_600;
assign col_out_601 = u5_col_out_601;
assign col_out_602 = u5_col_out_602;
assign col_out_603 = u5_col_out_603;
assign col_out_604 = u5_col_out_604;
assign col_out_605 = u5_col_out_605;
assign col_out_606 = u5_col_out_606;
assign col_out_607 = u5_col_out_607;
assign col_out_608 = u5_col_out_608;
assign col_out_609 = u5_col_out_609;
assign col_out_610 = u5_col_out_610;
assign col_out_611 = u5_col_out_611;
assign col_out_612 = u5_col_out_612;
assign col_out_613 = u5_col_out_613;
assign col_out_614 = u5_col_out_614;
assign col_out_615 = u5_col_out_615;
assign col_out_616 = u5_col_out_616;
assign col_out_617 = u5_col_out_617;
assign col_out_618 = u5_col_out_618;
assign col_out_619 = u5_col_out_619;
assign col_out_620 = u5_col_out_620;
assign col_out_621 = u5_col_out_621;
assign col_out_622 = u5_col_out_622;
assign col_out_623 = u5_col_out_623;
assign col_out_624 = u5_col_out_624;
assign col_out_625 = u5_col_out_625;
assign col_out_626 = u5_col_out_626;
assign col_out_627 = u5_col_out_627;
assign col_out_628 = u5_col_out_628;
assign col_out_629 = u5_col_out_629;
assign col_out_630 = u5_col_out_630;
assign col_out_631 = u5_col_out_631;
assign col_out_632 = u5_col_out_632;
assign col_out_633 = u5_col_out_633;
assign col_out_634 = u5_col_out_634;
assign col_out_635 = u5_col_out_635;
assign col_out_636 = u5_col_out_636;
assign col_out_637 = u5_col_out_637;
assign col_out_638 = u5_col_out_638;
assign col_out_639 = u5_col_out_639;
assign col_out_640 = u5_col_out_640;
assign col_out_641 = u5_col_out_641;
assign col_out_642 = u5_col_out_642;
assign col_out_643 = u5_col_out_643;
assign col_out_644 = u5_col_out_644;
assign col_out_645 = u5_col_out_645;
assign col_out_646 = u5_col_out_646;
assign col_out_647 = u5_col_out_647;
assign col_out_648 = u5_col_out_648;
assign col_out_649 = u5_col_out_649;
assign col_out_650 = u5_col_out_650;
assign col_out_651 = u5_col_out_651;
assign col_out_652 = u5_col_out_652;
assign col_out_653 = u5_col_out_653;
assign col_out_654 = u5_col_out_654;
assign col_out_655 = u5_col_out_655;
assign col_out_656 = u5_col_out_656;
assign col_out_657 = u5_col_out_657;
assign col_out_658 = u5_col_out_658;
assign col_out_659 = u5_col_out_659;
assign col_out_660 = u5_col_out_660;
assign col_out_661 = u5_col_out_661;
assign col_out_662 = u5_col_out_662;
assign col_out_663 = u5_col_out_663;
assign col_out_664 = u5_col_out_664;
assign col_out_665 = u5_col_out_665;
assign col_out_666 = u5_col_out_666;
assign col_out_667 = u5_col_out_667;
assign col_out_668 = u5_col_out_668;
assign col_out_669 = u5_col_out_669;
assign col_out_670 = u5_col_out_670;
assign col_out_671 = u5_col_out_671;
assign col_out_672 = u5_col_out_672;
assign col_out_673 = u5_col_out_673;
assign col_out_674 = u5_col_out_674;
assign col_out_675 = u5_col_out_675;
assign col_out_676 = u5_col_out_676;
assign col_out_677 = u5_col_out_677;
assign col_out_678 = u5_col_out_678;
assign col_out_679 = u5_col_out_679;
assign col_out_680 = u5_col_out_680;
assign col_out_681 = u5_col_out_681;
assign col_out_682 = u5_col_out_682;
assign col_out_683 = u5_col_out_683;
assign col_out_684 = u5_col_out_684;
assign col_out_685 = u5_col_out_685;
assign col_out_686 = u5_col_out_686;
assign col_out_687 = u5_col_out_687;
assign col_out_688 = u5_col_out_688;
assign col_out_689 = u5_col_out_689;
assign col_out_690 = u5_col_out_690;
assign col_out_691 = u5_col_out_691;
assign col_out_692 = u5_col_out_692;
assign col_out_693 = u5_col_out_693;
assign col_out_694 = u5_col_out_694;
assign col_out_695 = u5_col_out_695;
assign col_out_696 = u5_col_out_696;
assign col_out_697 = u5_col_out_697;
assign col_out_698 = u5_col_out_698;
assign col_out_699 = u5_col_out_699;
assign col_out_700 = u5_col_out_700;
assign col_out_701 = u5_col_out_701;
assign col_out_702 = u5_col_out_702;
assign col_out_703 = u5_col_out_703;
assign col_out_704 = u5_col_out_704;
assign col_out_705 = u5_col_out_705;
assign col_out_706 = u5_col_out_706;
assign col_out_707 = u5_col_out_707;
assign col_out_708 = u5_col_out_708;
assign col_out_709 = u5_col_out_709;
assign col_out_710 = u5_col_out_710;
assign col_out_711 = u5_col_out_711;
assign col_out_712 = u5_col_out_712;
assign col_out_713 = u5_col_out_713;
assign col_out_714 = u5_col_out_714;
assign col_out_715 = u5_col_out_715;
assign col_out_716 = u5_col_out_716;
assign col_out_717 = u5_col_out_717;
assign col_out_718 = u5_col_out_718;
assign col_out_719 = u5_col_out_719;
assign col_out_720 = u5_col_out_720;
assign col_out_721 = u5_col_out_721;
assign col_out_722 = u5_col_out_722;
assign col_out_723 = u5_col_out_723;
assign col_out_724 = u5_col_out_724;
assign col_out_725 = u5_col_out_725;
assign col_out_726 = u5_col_out_726;
assign col_out_727 = u5_col_out_727;
assign col_out_728 = u5_col_out_728;
assign col_out_729 = u5_col_out_729;
assign col_out_730 = u5_col_out_730;
assign col_out_731 = u5_col_out_731;
assign col_out_732 = u5_col_out_732;
assign col_out_733 = u5_col_out_733;
assign col_out_734 = u5_col_out_734;
assign col_out_735 = u5_col_out_735;
assign col_out_736 = u5_col_out_736;
assign col_out_737 = u5_col_out_737;
assign col_out_738 = u5_col_out_738;
assign col_out_739 = u5_col_out_739;
assign col_out_740 = u5_col_out_740;
assign col_out_741 = u5_col_out_741;
assign col_out_742 = u5_col_out_742;
assign col_out_743 = u5_col_out_743;
assign col_out_744 = u5_col_out_744;
assign col_out_745 = u5_col_out_745;
assign col_out_746 = u5_col_out_746;
assign col_out_747 = u5_col_out_747;
assign col_out_748 = u5_col_out_748;
assign col_out_749 = u5_col_out_749;
assign col_out_750 = u5_col_out_750;
assign col_out_751 = u5_col_out_751;
assign col_out_752 = u5_col_out_752;
assign col_out_753 = u5_col_out_753;
assign col_out_754 = u5_col_out_754;
assign col_out_755 = u5_col_out_755;
assign col_out_756 = u5_col_out_756;
assign col_out_757 = u5_col_out_757;
assign col_out_758 = u5_col_out_758;
assign col_out_759 = u5_col_out_759;
assign col_out_760 = u5_col_out_760;
assign col_out_761 = u5_col_out_761;
assign col_out_762 = u5_col_out_762;
assign col_out_763 = u5_col_out_763;
assign col_out_764 = u5_col_out_764;
assign col_out_765 = u5_col_out_765;
assign col_out_766 = u5_col_out_766;
assign col_out_767 = u5_col_out_767;
assign col_out_768 = u5_col_out_768;
assign col_out_769 = u5_col_out_769;
assign col_out_770 = u5_col_out_770;
assign col_out_771 = u5_col_out_771;
assign col_out_772 = u5_col_out_772;
assign col_out_773 = u5_col_out_773;
assign col_out_774 = u5_col_out_774;
assign col_out_775 = u5_col_out_775;
assign col_out_776 = u5_col_out_776;
assign col_out_777 = u5_col_out_777;
assign col_out_778 = u5_col_out_778;
assign col_out_779 = u5_col_out_779;
assign col_out_780 = u5_col_out_780;
assign col_out_781 = u5_col_out_781;
assign col_out_782 = u5_col_out_782;
assign col_out_783 = u5_col_out_783;
assign col_out_784 = u5_col_out_784;
assign col_out_785 = u5_col_out_785;
assign col_out_786 = u5_col_out_786;
assign col_out_787 = u5_col_out_787;
assign col_out_788 = u5_col_out_788;
assign col_out_789 = u5_col_out_789;
assign col_out_790 = u5_col_out_790;
assign col_out_791 = u5_col_out_791;
assign col_out_792 = u5_col_out_792;
assign col_out_793 = u5_col_out_793;
assign col_out_794 = u5_col_out_794;
assign col_out_795 = u5_col_out_795;
assign col_out_796 = u5_col_out_796;
assign col_out_797 = u5_col_out_797;
assign col_out_798 = u5_col_out_798;
assign col_out_799 = u5_col_out_799;
assign col_out_800 = u5_col_out_800;
assign col_out_801 = u5_col_out_801;
assign col_out_802 = u5_col_out_802;
assign col_out_803 = u5_col_out_803;
assign col_out_804 = u5_col_out_804;
assign col_out_805 = u5_col_out_805;
assign col_out_806 = u5_col_out_806;
assign col_out_807 = u5_col_out_807;
assign col_out_808 = u5_col_out_808;
assign col_out_809 = u5_col_out_809;
assign col_out_810 = u5_col_out_810;
assign col_out_811 = u5_col_out_811;
assign col_out_812 = u5_col_out_812;
assign col_out_813 = u5_col_out_813;
assign col_out_814 = u5_col_out_814;
assign col_out_815 = u5_col_out_815;
assign col_out_816 = u5_col_out_816;
assign col_out_817 = u5_col_out_817;
assign col_out_818 = u5_col_out_818;
assign col_out_819 = u5_col_out_819;
assign col_out_820 = u5_col_out_820;
assign col_out_821 = u5_col_out_821;
assign col_out_822 = u5_col_out_822;
assign col_out_823 = u5_col_out_823;
assign col_out_824 = u5_col_out_824;
assign col_out_825 = u5_col_out_825;
assign col_out_826 = u5_col_out_826;
assign col_out_827 = u5_col_out_827;
assign col_out_828 = u5_col_out_828;
assign col_out_829 = u5_col_out_829;
assign col_out_830 = u5_col_out_830;
assign col_out_831 = u5_col_out_831;
assign col_out_832 = u5_col_out_832;
assign col_out_833 = u5_col_out_833;
assign col_out_834 = u5_col_out_834;
assign col_out_835 = u5_col_out_835;
assign col_out_836 = u5_col_out_836;
assign col_out_837 = u5_col_out_837;
assign col_out_838 = u5_col_out_838;
assign col_out_839 = u5_col_out_839;
assign col_out_840 = u5_col_out_840;
assign col_out_841 = u5_col_out_841;
assign col_out_842 = u5_col_out_842;
assign col_out_843 = u5_col_out_843;
assign col_out_844 = u5_col_out_844;
assign col_out_845 = u5_col_out_845;
assign col_out_846 = u5_col_out_846;
assign col_out_847 = u5_col_out_847;
assign col_out_848 = u5_col_out_848;
assign col_out_849 = u5_col_out_849;
assign col_out_850 = u5_col_out_850;
assign col_out_851 = u5_col_out_851;
assign col_out_852 = u5_col_out_852;
assign col_out_853 = u5_col_out_853;
assign col_out_854 = u5_col_out_854;
assign col_out_855 = u5_col_out_855;
assign col_out_856 = u5_col_out_856;
assign col_out_857 = u5_col_out_857;
assign col_out_858 = u5_col_out_858;
assign col_out_859 = u5_col_out_859;
assign col_out_860 = u5_col_out_860;
assign col_out_861 = u5_col_out_861;
assign col_out_862 = u5_col_out_862;
assign col_out_863 = u5_col_out_863;
assign col_out_864 = u5_col_out_864;
assign col_out_865 = u5_col_out_865;
assign col_out_866 = u5_col_out_866;
assign col_out_867 = u5_col_out_867;
assign col_out_868 = u5_col_out_868;
assign col_out_869 = u5_col_out_869;
assign col_out_870 = u5_col_out_870;
assign col_out_871 = u5_col_out_871;
assign col_out_872 = u5_col_out_872;
assign col_out_873 = u5_col_out_873;
assign col_out_874 = u5_col_out_874;
assign col_out_875 = u5_col_out_875;
assign col_out_876 = u5_col_out_876;
assign col_out_877 = u5_col_out_877;
assign col_out_878 = u5_col_out_878;
assign col_out_879 = u5_col_out_879;
assign col_out_880 = u5_col_out_880;
assign col_out_881 = u5_col_out_881;
assign col_out_882 = u5_col_out_882;
assign col_out_883 = u5_col_out_883;
assign col_out_884 = u5_col_out_884;
assign col_out_885 = u5_col_out_885;
assign col_out_886 = u5_col_out_886;
assign col_out_887 = u5_col_out_887;
assign col_out_888 = u5_col_out_888;
assign col_out_889 = u5_col_out_889;
assign col_out_890 = u5_col_out_890;
assign col_out_891 = u5_col_out_891;
assign col_out_892 = u5_col_out_892;
assign col_out_893 = u5_col_out_893;
assign col_out_894 = u5_col_out_894;
assign col_out_895 = u5_col_out_895;
assign col_out_896 = u5_col_out_896;
assign col_out_897 = u5_col_out_897;
assign col_out_898 = u5_col_out_898;
assign col_out_899 = u5_col_out_899;
assign col_out_900 = u5_col_out_900;
assign col_out_901 = u5_col_out_901;
assign col_out_902 = u5_col_out_902;
assign col_out_903 = u5_col_out_903;
assign col_out_904 = u5_col_out_904;
assign col_out_905 = u5_col_out_905;
assign col_out_906 = u5_col_out_906;
assign col_out_907 = u5_col_out_907;
assign col_out_908 = u5_col_out_908;
assign col_out_909 = u5_col_out_909;
assign col_out_910 = u5_col_out_910;
assign col_out_911 = u5_col_out_911;
assign col_out_912 = u5_col_out_912;
assign col_out_913 = u5_col_out_913;
assign col_out_914 = u5_col_out_914;
assign col_out_915 = u5_col_out_915;
assign col_out_916 = u5_col_out_916;
assign col_out_917 = u5_col_out_917;
assign col_out_918 = u5_col_out_918;
assign col_out_919 = u5_col_out_919;
assign col_out_920 = u5_col_out_920;
assign col_out_921 = u5_col_out_921;
assign col_out_922 = u5_col_out_922;
assign col_out_923 = u5_col_out_923;
assign col_out_924 = u5_col_out_924;
assign col_out_925 = u5_col_out_925;
assign col_out_926 = u5_col_out_926;
assign col_out_927 = u5_col_out_927;
assign col_out_928 = u5_col_out_928;
assign col_out_929 = u5_col_out_929;
assign col_out_930 = u5_col_out_930;
assign col_out_931 = u5_col_out_931;
assign col_out_932 = u5_col_out_932;
assign col_out_933 = u5_col_out_933;
assign col_out_934 = u5_col_out_934;
assign col_out_935 = u5_col_out_935;
assign col_out_936 = u5_col_out_936;
assign col_out_937 = u5_col_out_937;
assign col_out_938 = u5_col_out_938;
assign col_out_939 = u5_col_out_939;
assign col_out_940 = u5_col_out_940;
assign col_out_941 = u5_col_out_941;
assign col_out_942 = u5_col_out_942;
assign col_out_943 = u5_col_out_943;
assign col_out_944 = u5_col_out_944;
assign col_out_945 = u5_col_out_945;
assign col_out_946 = u5_col_out_946;
assign col_out_947 = u5_col_out_947;
assign col_out_948 = u5_col_out_948;
assign col_out_949 = u5_col_out_949;
assign col_out_950 = u5_col_out_950;
assign col_out_951 = u5_col_out_951;
assign col_out_952 = u5_col_out_952;
assign col_out_953 = u5_col_out_953;
assign col_out_954 = u5_col_out_954;
assign col_out_955 = u5_col_out_955;
assign col_out_956 = u5_col_out_956;
assign col_out_957 = u5_col_out_957;
assign col_out_958 = u5_col_out_958;
assign col_out_959 = u5_col_out_959;
assign col_out_960 = u5_col_out_960;
assign col_out_961 = u5_col_out_961;
assign col_out_962 = u5_col_out_962;
assign col_out_963 = u5_col_out_963;
assign col_out_964 = u5_col_out_964;
assign col_out_965 = u5_col_out_965;
assign col_out_966 = u5_col_out_966;
assign col_out_967 = u5_col_out_967;
assign col_out_968 = u5_col_out_968;
assign col_out_969 = u5_col_out_969;
assign col_out_970 = u5_col_out_970;
assign col_out_971 = u5_col_out_971;
assign col_out_972 = u5_col_out_972;
assign col_out_973 = u5_col_out_973;
assign col_out_974 = u5_col_out_974;
assign col_out_975 = u5_col_out_975;
assign col_out_976 = u5_col_out_976;
assign col_out_977 = u5_col_out_977;
assign col_out_978 = u5_col_out_978;
assign col_out_979 = u5_col_out_979;
assign col_out_980 = u5_col_out_980;
assign col_out_981 = u5_col_out_981;
assign col_out_982 = u5_col_out_982;
assign col_out_983 = u5_col_out_983;
assign col_out_984 = u5_col_out_984;
assign col_out_985 = u5_col_out_985;
assign col_out_986 = u5_col_out_986;
assign col_out_987 = u5_col_out_987;
assign col_out_988 = u5_col_out_988;
assign col_out_989 = u5_col_out_989;
assign col_out_990 = u5_col_out_990;
assign col_out_991 = u5_col_out_991;
assign col_out_992 = u5_col_out_992;
assign col_out_993 = u5_col_out_993;
assign col_out_994 = u5_col_out_994;
assign col_out_995 = u5_col_out_995;
assign col_out_996 = u5_col_out_996;
assign col_out_997 = u5_col_out_997;
assign col_out_998 = u5_col_out_998;
assign col_out_999 = u5_col_out_999;
assign col_out_1000 = u5_col_out_1000;
assign col_out_1001 = u5_col_out_1001;
assign col_out_1002 = u5_col_out_1002;
assign col_out_1003 = u5_col_out_1003;
assign col_out_1004 = u5_col_out_1004;
assign col_out_1005 = u5_col_out_1005;
assign col_out_1006 = u5_col_out_1006;
assign col_out_1007 = u5_col_out_1007;
assign col_out_1008 = u5_col_out_1008;
assign col_out_1009 = u5_col_out_1009;
assign col_out_1010 = u5_col_out_1010;
assign col_out_1011 = u5_col_out_1011;
assign col_out_1012 = u5_col_out_1012;
assign col_out_1013 = u5_col_out_1013;
assign col_out_1014 = u5_col_out_1014;
assign col_out_1015 = u5_col_out_1015;
assign col_out_1016 = u5_col_out_1016;
assign col_out_1017 = u5_col_out_1017;
assign col_out_1018 = u5_col_out_1018;
assign col_out_1019 = u5_col_out_1019;
assign col_out_1020 = u5_col_out_1020;
assign col_out_1021 = u5_col_out_1021;
assign col_out_1022 = u5_col_out_1022;
assign col_out_1023 = u5_col_out_1023;
assign col_out_1024 = u5_col_out_1024;
assign col_out_1025 = u5_col_out_1025;
assign col_out_1026 = u5_col_out_1026;
assign col_out_1027 = u5_col_out_1027;
assign col_out_1028 = u5_col_out_1028;
assign col_out_1029 = u5_col_out_1029;
assign col_out_1030 = u5_col_out_1030;
assign col_out_1031 = u5_col_out_1031;
assign col_out_1032 = u5_col_out_1032;




endmodule
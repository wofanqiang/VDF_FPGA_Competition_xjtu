module xpb_5_560
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h69e030c962752b49149b89fee6d8afbdf78872dd23a35f30c9641c3f57d9732df18a190f6676dd4055ac19328eaa72c6e66b38ebdd5652c628448376749e8deafc2a00849572291fc9d98a32f09150466070c97fb4af3b78abd7a8a6c8aa610ac4e6c850ebccdc461c022056ab1fb3b09631b0dee2842079dcd530193c2ef08a;
    5'b00010 : xpb = 1024'h23131c3d02fc21c95e319c26bd57182a7d9ae28971cf1dea14eb7f28fcb03953dfcbb4a602c73bf20bf9f31e39f6d4c368bc49f197f9d5409fe9c78eae6aa7248404cc5a7b5354fa811911c34846dc5bccdc9966dcd849e0a222bf52d72a1f835ac5fe7826d0bffeb14459ce5e6f4137dd8982db74bce3c3733ae52def7b7aa9;
    5'b00011 : xpb = 1024'h8cf34d0665714d1272cd2625a42fc7e87523556695727d1ade4f9b685489ac81d155cdb5693e193261a60c50c8a1478a4f2782dd75502806c82e4b052309350f802eccdf10c57e1a4af29bf638d82ca22d4d62e6918785594dfa67f99fd4808e1facc6c9129d9c44cd467a25098ef4e873bb33ba5741043d501015472baa6b33;
    5'b00100 : xpb = 1024'h4626387a05f84392bc63384d7aae3054fb35c512e39e3bd429d6fe51f96072a7bf97694c058e77e417f3e63c73eda986d17893e32ff3aa813fd38f1d5cd54e49080998b4f6a6a9f502322386908db8b799b932cdb9b093c144457ea5ae543f06b58bfcf04da17ffd6288b39cbcde826fbb1305b6e979c786e675ca5bdef6f552;
    5'b00101 : xpb = 1024'hb0066943686d6edbd0fec24c6186e012f2be37f007419b04f33b1a915139e5d5b121825b6c0555246d9fff6f02981c4db7e3cccf0d49fd4768181293d173dc34043399398c18d314cc0badb9811f08fdfa29fc4d6e5fcf39f01d274c76fea0117a72c541396e5c437e8ad3f367fe36205144b695cbfde800c34afa751b25e5dc;
    5'b00110 : xpb = 1024'h693954b708f4655c1a94d4743805487f78d0a79c556d59be3ec27d7af610abfb9f631df20855b3d623edd95aade47e4a3a34ddd4c7ed7fc1dfbd56ac0b3ff56d8c0e650f71f9feef834b3549d8d495136695cc349688dda1e6683df8857e5e8a1051fb6874723ffc13cd0d6b1b4dc3a7989c88925e36ab4a59b0af89ce726ffb;
    5'b00111 : xpb = 1024'h226c402aa97b5bdc642ae69c0e83b0ebfee31748a39918778a49e0649ae772218da4b988a4a61287da3bb3465930e046bc85eeda8291023c57629ac4450c0ea713e930e557db2aca3a8abcda308a2128d3019c1bbeb1ec09dcb354a493fe1d02a631318faf7623b4a90f46e2ce9d512edff45a8ef06f6e93f016649e81befa1a;
    5'b01000 : xpb = 1024'h8c4c70f40bf0872578c6709af55c60a9f66b8a25c73c77a853adfca3f2c0e54f7f2ed2980b1cefc82fe7cc78e7db530da2f127c65fe755027fa71e3ab9aa9c9210133169ed4d53ea0464470d211b716f3372659b73612782888afd4b5ca87e0d6b17f9e09b42fffac511673979bd04df76260b6dd2f38f0dcceb94b7bdedeaa4;
    5'b01001 : xpb = 1024'h457f5c67ac777da5c25c82c2cbdac9167c7df9d2156836619f355f8d9797ab756d706e2ea76d4e79e635a6649327b50a254238cc1a8ad77cf74c6252f376b5cb97edfd3fd32e7fc4bba3ce9d78d0fd849fde35829b8a35ea7ed613f76b283c8600f73007d646e3b35a53a0b12d0c9266bd7ddd6a652c5257635149cc713a74c3;
    5'b01010 : xpb = 1024'haf5f8d310eeca8eed6f80cc1b2b378d474066caf390b959268997bccef711ea35efa873e0de42bba3be1bf9721d227d10bad71b7f7e12a431f90e5c9681543b69417fdc468a0a8e4857d58d069624dcb004eff02503971632aadbc9e33d29d90c5ddf858c213bff97655c107d82c461753af8e4947b072d1402679e5ad69654d;
    5'b01011 : xpb = 1024'h689278a4af739f6f208e1ee98931e140fa18dc5b8737544bb420deb69447e4c94d3c22d4aa348a6bf22f9982cd1e89cd8dfe82bdb284acbd973629e1a1e15cf01bf2c99a4e81d4bf3cbce060c117d9e06cbacee978627fcb20f8d34a42525c095bbd2e7ffd17a3b20b97fa7f8b7bd39e9b076045d9e9361ad68c2efa60b5ef6c;
    5'b01100 : xpb = 1024'h21c564184ffa95ef6a2431115fb049ad802b4c07d5631304ffa841a0391eaaef3b7dbe6b4684e91da87d736e786aebca104f93c36d282f380edb6df9dbad7629a3cd957034630099f3fc67f118cd65f5d9269ed0a08b8e331743e9f650d21a81f19c64a7381b876aa0da33f73ecb6125e25f32426c21f9646cf1e40f1402798b;
    5'b01101 : xpb = 1024'h8ba594e1b26fc1387ebfbb104688f96b77b3bee4f9067235c90c5ddf90f81e1d2d07d77aacfbc65dfe298ca107155e90f6baccaf4a7e81fe371ff170504c04149ff795f4c9d529b9bdd5f224095eb63c39976850553ac9abc31b929d197c7b8cb6832cf823e863b0bcdc544de9eb14d67890e3214ea619de49c7142850316a15;
    5'b01110 : xpb = 1024'h44d8805552f6b7b8c855cd381d0761d7fdc62e91473230ef1493c0c935cee4431b497311494c250fb477668cb261c08d790bddb505220478aec535888a181d4e27d261caafb65594751579b461144251a60338377d63d813b966a94927fc3a054c62631f5eec4769521e8dc59d3aa25dbfe8b51de0dedd27e02cc93d037df434;
    5'b01111 : xpb = 1024'haeb8b11eb56be301dcf1573703e01195f54ea16e6ad5901fddf7dd088da857710cd38c20afc302500a237fbf410c33545f7716a0e278573ed709b8fefeb6ab3923fc624f45287eb43eef03e751a59298067401b73213138c653e51eff0a69b1011492b704ab923af6e20ae1c485a560e561a65fcc362fda1bd01f9563face4be;
    5'b10000 : xpb = 1024'h67eb9c9255f2d9822687695eda5e7a027b61111ab9014ed9297f3ff2327f1d96fb1527b74c136101c07159aaec589550e1c827a69d1bd9b94eaefd173882c472abd72e252b09aa8ef62e8b77a95b1ead72dfd19e5a3c21f45b89689bff265988a728619785bd07680362e793fba9e3959d7237f9559bc0eb5367ae6af2f96edd;
    5'b10001 : xpb = 1024'h211e8805f679d002701d7b86b0dce26f017380c7072d0d927506a2dbd755e3bce956c34de863bfb376bf339697a4f74d641938ac57bf5c33c654412f724eddac33b1f9fb10ead669ad6e13080110aac2df4ba1858265305c51d47f480da618013d0797bec0c0eb2098a5210baef9711ce4ca09f5e7d48434e9cd637fa645f8fc;
    5'b10010 : xpb = 1024'h8afeb8cf58eefb4b84b9058597b5922cf8fbf3a42ad06cc33e6abf1b2f2f56eadae0dc5d4eda9cf3cc6b4cc9264f6a144a8471983515aef9ee98c4a5e6ed6b972fdbfa7fa65cff8977479d3af1a1fb093fbc6b0537146bd4fdac27eed650790c01ee600fac8dc766b4a741625a1924cd7afbbad4ca58a4aec6a29398e274e986;
    5'b10011 : xpb = 1024'h4431a442f975f1cbce4f17ad6e33fa997f0e635078fc2b7c89f22204d4061d10c92277f3eb2afba582b926b4d19bcc10ccd5829defb93174663e08be20b984d0b7b6c6558c3e2b642e8724cb4957871eac283aec5f3d7a3cf3f73e9ae4d0378497cd9636e791ab1f49e97ada0d68b254c2538cd15c9167f85d0848ad95c173a5;
    5'b10100 : xpb = 1024'hae11d50c5beb1d14e2eaa1ac550caa577696d62d9c9f8aad53563e442bdf903ebaac910351a1d8e5d8653fe760463ed7b340bb89cd0f843a8e828c34955812bbb3e0c6da21b05483f860aefe39e8d7650c99046c13ecb5b59fcee741ad7a988f5cb45e87d35e876565eb9b30b888660558853db03f15887239dd78c6d1f0642f;
    5'b10101 : xpb = 1024'h6744c07ffc7213952c80b3d42b8b12c3fca945d9eacb49669edda12dd0b65664a8ee2c99edf237978eb319d30b92a0d43591cc8f87b306b50627d04ccf242bf53bbb92b00791805eafa0368e919e637a7904d4533c15c41d9619fdedbbfa5707f29394af0e626b1dfb2dd4a86bd7f38c9fdd0facd14e4bbbd0432ddb853cee4e;
    5'b10110 : xpb = 1024'h2077abf39cf90a157616c5fc02097b3082bbb58638f7081fea650417758d1c8a972fc8308a4296494500f3beb6df02d0b7e2dd954256892f7dcd146508f0452ec3965e85ed72ac3966dfbe1ee953ef8fe570a43a643ed2858c651499ca7a15808872cad649664ed690700e201f278113e734e1a963870f0566a8e2f03889786d;
    5'b10111 : xpb = 1024'h8a57dcbcff6e355e8ab24ffae8e22aee7a4428635c9a6750b3c92056cd668fb888b9e13ff0b973899aad0cf1458975979e4e16811facdbf5a61197db7d8ed319bfc05f0a82e4d55930b94851d9e53fd645e16dba18ee0dfe383cbd409324768b4d59932735332b1cac722e76ca4734c47d669288460b2f7f437e130974b868f7;
    5'b11000 : xpb = 1024'h438ac8309ff52bded4486222bf60935b0056980faac62609ff508340723d55de76fb7cd68d09d23b50fae6dcf0d5d794209f2786da505e701db6dbf3b75aec53479b2ae068c60133e7f8cfe2319acbebb24d3da141171c662e87d3eca1a43503e338c94e70370ed541b467ee7d96c24bc4be6484d843f2c8d9e3c81e2804f316;
    5'b11001 : xpb = 1024'had6af8fa026a5727e8e3ec21a6394318f7df0aecce69853ac8b49f7fca16c90c688595e5f380af7ba6a7000f7f804a5b070a6072b7a6b13645fb5f6a2bf97a3e43c52b64fe382a53b1d25a15222c1c3212be0720f5c657deda5f7c936a4e960ea81f919f5c03eb1b5db6884528b675fc5af01563bac81342b6b8f8376433e3a0;
    5'b11010 : xpb = 1024'h669de46da2f14da83279fe497cb7ab857df17a991c9543f4143c02696eed8f3256c7317c8fd10e2d5cf4d9fb2accac57895b7178724a33b0bda0a38265c59377cb9ff73ae419562e6911e1a579e1a8477f29d7081def6646d0aa933f78ce54873dfec7c69707ced3f2f8c1bcdc060383a247e7604d00d68c4d1ead4c17806dbf;
    5'b11011 : xpb = 1024'h1fd0cfe1437844287c101071533613f20403ea456ac102ad5fc3655313c455584508cd132c216cdf1342b3e6d6190e540bac827e2cedb62b3545e79a9f91acb1537ac310c9fa820920516935d197345ceb95a6ef461874aec6f5a9eb874e12ffd3ddfdedd20bb28c883afb348f55910ae99fb95cdf3999d5e3846260caccf7de;
    5'b11100 : xpb = 1024'h89b100aaa5ed6f7190ab9a703a0ec3affb8c5d228e6461de292781926b9dc8863692e62292984a1f68eecd1964c3811af217bb6a0a4408f15d8a6b1114303a9c4fa4c3955f6cab28ea2af368c22884a34c06706efac7b02772cd52924ff8740a98c4c63ebdd88ed2a43d1b8b3a7544bb7fd16a3bc1bdba4fc059927a06fbe868;
    5'b11101 : xpb = 1024'h42e3ec1e467465f1da41ac98108d2c1c819ecccedc90209774aee47c10748eac24d481b92ee8a8d11f3ca705100fe3177468cc6fc4e78b6bd52faf294dfc53d5d77f8f6b454dd703a16a7af919de10b8b872405622f0be8f6918693e5e7832832ea3fc65f8dc728b397f5502edc4d242c7293c3853f67d9956bf478eba487287;
    5'b11110 : xpb = 1024'hacc41ce7a8e9913aeedd3696f765dbda79273fac00337fc83e1300bb684e01da165e9ac8955f861174e8c0379eba55de5ad4055ba23dde31fd74329fc29ae1c0d3a98fefdac000236b44052c0a6f60ff18e309d5d79ffa0814f011e52722938df38ac4b6e4a94ed15581755998e485f35d5aed17367a9e13339477a7f6776311;
    5'b11111 : xpb = 1024'h65f7085b497087bb387348becde44446ff39af584e5f3e81899a63a50d24c80004a0365f31afe4c32b369a234a06b7dadd2516615ce160ac751976b7fc66fafa5b845bc5c0a12bfe22838cbc6224ed14854ed9bcffc908700b3b289135a252068969fade1fad3289eac3aed14c34137aa4b2bf13c8b3615cc9fa2cbca9c3ed30;
    endcase
end

endmodule

module compressor_array_512_2_1024_row
(
    input  [511:0] col_in_0,
    input  [511:0] col_in_1,
    input  [511:0] col_in_2,
    input  [511:0] col_in_3,
    input  [511:0] col_in_4,
    input  [511:0] col_in_5,
    input  [511:0] col_in_6,
    input  [511:0] col_in_7,
    input  [511:0] col_in_8,
    input  [511:0] col_in_9,
    input  [511:0] col_in_10,
    input  [511:0] col_in_11,
    input  [511:0] col_in_12,
    input  [511:0] col_in_13,
    input  [511:0] col_in_14,
    input  [511:0] col_in_15,
    input  [511:0] col_in_16,
    input  [511:0] col_in_17,
    input  [511:0] col_in_18,
    input  [511:0] col_in_19,
    input  [511:0] col_in_20,
    input  [511:0] col_in_21,
    input  [511:0] col_in_22,
    input  [511:0] col_in_23,
    input  [511:0] col_in_24,
    input  [511:0] col_in_25,
    input  [511:0] col_in_26,
    input  [511:0] col_in_27,
    input  [511:0] col_in_28,
    input  [511:0] col_in_29,
    input  [511:0] col_in_30,
    input  [511:0] col_in_31,
    input  [511:0] col_in_32,
    input  [511:0] col_in_33,
    input  [511:0] col_in_34,
    input  [511:0] col_in_35,
    input  [511:0] col_in_36,
    input  [511:0] col_in_37,
    input  [511:0] col_in_38,
    input  [511:0] col_in_39,
    input  [511:0] col_in_40,
    input  [511:0] col_in_41,
    input  [511:0] col_in_42,
    input  [511:0] col_in_43,
    input  [511:0] col_in_44,
    input  [511:0] col_in_45,
    input  [511:0] col_in_46,
    input  [511:0] col_in_47,
    input  [511:0] col_in_48,
    input  [511:0] col_in_49,
    input  [511:0] col_in_50,
    input  [511:0] col_in_51,
    input  [511:0] col_in_52,
    input  [511:0] col_in_53,
    input  [511:0] col_in_54,
    input  [511:0] col_in_55,
    input  [511:0] col_in_56,
    input  [511:0] col_in_57,
    input  [511:0] col_in_58,
    input  [511:0] col_in_59,
    input  [511:0] col_in_60,
    input  [511:0] col_in_61,
    input  [511:0] col_in_62,
    input  [511:0] col_in_63,
    input  [511:0] col_in_64,
    input  [511:0] col_in_65,
    input  [511:0] col_in_66,
    input  [511:0] col_in_67,
    input  [511:0] col_in_68,
    input  [511:0] col_in_69,
    input  [511:0] col_in_70,
    input  [511:0] col_in_71,
    input  [511:0] col_in_72,
    input  [511:0] col_in_73,
    input  [511:0] col_in_74,
    input  [511:0] col_in_75,
    input  [511:0] col_in_76,
    input  [511:0] col_in_77,
    input  [511:0] col_in_78,
    input  [511:0] col_in_79,
    input  [511:0] col_in_80,
    input  [511:0] col_in_81,
    input  [511:0] col_in_82,
    input  [511:0] col_in_83,
    input  [511:0] col_in_84,
    input  [511:0] col_in_85,
    input  [511:0] col_in_86,
    input  [511:0] col_in_87,
    input  [511:0] col_in_88,
    input  [511:0] col_in_89,
    input  [511:0] col_in_90,
    input  [511:0] col_in_91,
    input  [511:0] col_in_92,
    input  [511:0] col_in_93,
    input  [511:0] col_in_94,
    input  [511:0] col_in_95,
    input  [511:0] col_in_96,
    input  [511:0] col_in_97,
    input  [511:0] col_in_98,
    input  [511:0] col_in_99,
    input  [511:0] col_in_100,
    input  [511:0] col_in_101,
    input  [511:0] col_in_102,
    input  [511:0] col_in_103,
    input  [511:0] col_in_104,
    input  [511:0] col_in_105,
    input  [511:0] col_in_106,
    input  [511:0] col_in_107,
    input  [511:0] col_in_108,
    input  [511:0] col_in_109,
    input  [511:0] col_in_110,
    input  [511:0] col_in_111,
    input  [511:0] col_in_112,
    input  [511:0] col_in_113,
    input  [511:0] col_in_114,
    input  [511:0] col_in_115,
    input  [511:0] col_in_116,
    input  [511:0] col_in_117,
    input  [511:0] col_in_118,
    input  [511:0] col_in_119,
    input  [511:0] col_in_120,
    input  [511:0] col_in_121,
    input  [511:0] col_in_122,
    input  [511:0] col_in_123,
    input  [511:0] col_in_124,
    input  [511:0] col_in_125,
    input  [511:0] col_in_126,
    input  [511:0] col_in_127,
    input  [511:0] col_in_128,
    input  [511:0] col_in_129,
    input  [511:0] col_in_130,
    input  [511:0] col_in_131,
    input  [511:0] col_in_132,
    input  [511:0] col_in_133,
    input  [511:0] col_in_134,
    input  [511:0] col_in_135,
    input  [511:0] col_in_136,
    input  [511:0] col_in_137,
    input  [511:0] col_in_138,
    input  [511:0] col_in_139,
    input  [511:0] col_in_140,
    input  [511:0] col_in_141,
    input  [511:0] col_in_142,
    input  [511:0] col_in_143,
    input  [511:0] col_in_144,
    input  [511:0] col_in_145,
    input  [511:0] col_in_146,
    input  [511:0] col_in_147,
    input  [511:0] col_in_148,
    input  [511:0] col_in_149,
    input  [511:0] col_in_150,
    input  [511:0] col_in_151,
    input  [511:0] col_in_152,
    input  [511:0] col_in_153,
    input  [511:0] col_in_154,
    input  [511:0] col_in_155,
    input  [511:0] col_in_156,
    input  [511:0] col_in_157,
    input  [511:0] col_in_158,
    input  [511:0] col_in_159,
    input  [511:0] col_in_160,
    input  [511:0] col_in_161,
    input  [511:0] col_in_162,
    input  [511:0] col_in_163,
    input  [511:0] col_in_164,
    input  [511:0] col_in_165,
    input  [511:0] col_in_166,
    input  [511:0] col_in_167,
    input  [511:0] col_in_168,
    input  [511:0] col_in_169,
    input  [511:0] col_in_170,
    input  [511:0] col_in_171,
    input  [511:0] col_in_172,
    input  [511:0] col_in_173,
    input  [511:0] col_in_174,
    input  [511:0] col_in_175,
    input  [511:0] col_in_176,
    input  [511:0] col_in_177,
    input  [511:0] col_in_178,
    input  [511:0] col_in_179,
    input  [511:0] col_in_180,
    input  [511:0] col_in_181,
    input  [511:0] col_in_182,
    input  [511:0] col_in_183,
    input  [511:0] col_in_184,
    input  [511:0] col_in_185,
    input  [511:0] col_in_186,
    input  [511:0] col_in_187,
    input  [511:0] col_in_188,
    input  [511:0] col_in_189,
    input  [511:0] col_in_190,
    input  [511:0] col_in_191,
    input  [511:0] col_in_192,
    input  [511:0] col_in_193,
    input  [511:0] col_in_194,
    input  [511:0] col_in_195,
    input  [511:0] col_in_196,
    input  [511:0] col_in_197,
    input  [511:0] col_in_198,
    input  [511:0] col_in_199,
    input  [511:0] col_in_200,
    input  [511:0] col_in_201,
    input  [511:0] col_in_202,
    input  [511:0] col_in_203,
    input  [511:0] col_in_204,
    input  [511:0] col_in_205,
    input  [511:0] col_in_206,
    input  [511:0] col_in_207,
    input  [511:0] col_in_208,
    input  [511:0] col_in_209,
    input  [511:0] col_in_210,
    input  [511:0] col_in_211,
    input  [511:0] col_in_212,
    input  [511:0] col_in_213,
    input  [511:0] col_in_214,
    input  [511:0] col_in_215,
    input  [511:0] col_in_216,
    input  [511:0] col_in_217,
    input  [511:0] col_in_218,
    input  [511:0] col_in_219,
    input  [511:0] col_in_220,
    input  [511:0] col_in_221,
    input  [511:0] col_in_222,
    input  [511:0] col_in_223,
    input  [511:0] col_in_224,
    input  [511:0] col_in_225,
    input  [511:0] col_in_226,
    input  [511:0] col_in_227,
    input  [511:0] col_in_228,
    input  [511:0] col_in_229,
    input  [511:0] col_in_230,
    input  [511:0] col_in_231,
    input  [511:0] col_in_232,
    input  [511:0] col_in_233,
    input  [511:0] col_in_234,
    input  [511:0] col_in_235,
    input  [511:0] col_in_236,
    input  [511:0] col_in_237,
    input  [511:0] col_in_238,
    input  [511:0] col_in_239,
    input  [511:0] col_in_240,
    input  [511:0] col_in_241,
    input  [511:0] col_in_242,
    input  [511:0] col_in_243,
    input  [511:0] col_in_244,
    input  [511:0] col_in_245,
    input  [511:0] col_in_246,
    input  [511:0] col_in_247,
    input  [511:0] col_in_248,
    input  [511:0] col_in_249,
    input  [511:0] col_in_250,
    input  [511:0] col_in_251,
    input  [511:0] col_in_252,
    input  [511:0] col_in_253,
    input  [511:0] col_in_254,
    input  [511:0] col_in_255,
    input  [511:0] col_in_256,
    input  [511:0] col_in_257,
    input  [511:0] col_in_258,
    input  [511:0] col_in_259,
    input  [511:0] col_in_260,
    input  [511:0] col_in_261,
    input  [511:0] col_in_262,
    input  [511:0] col_in_263,
    input  [511:0] col_in_264,
    input  [511:0] col_in_265,
    input  [511:0] col_in_266,
    input  [511:0] col_in_267,
    input  [511:0] col_in_268,
    input  [511:0] col_in_269,
    input  [511:0] col_in_270,
    input  [511:0] col_in_271,
    input  [511:0] col_in_272,
    input  [511:0] col_in_273,
    input  [511:0] col_in_274,
    input  [511:0] col_in_275,
    input  [511:0] col_in_276,
    input  [511:0] col_in_277,
    input  [511:0] col_in_278,
    input  [511:0] col_in_279,
    input  [511:0] col_in_280,
    input  [511:0] col_in_281,
    input  [511:0] col_in_282,
    input  [511:0] col_in_283,
    input  [511:0] col_in_284,
    input  [511:0] col_in_285,
    input  [511:0] col_in_286,
    input  [511:0] col_in_287,
    input  [511:0] col_in_288,
    input  [511:0] col_in_289,
    input  [511:0] col_in_290,
    input  [511:0] col_in_291,
    input  [511:0] col_in_292,
    input  [511:0] col_in_293,
    input  [511:0] col_in_294,
    input  [511:0] col_in_295,
    input  [511:0] col_in_296,
    input  [511:0] col_in_297,
    input  [511:0] col_in_298,
    input  [511:0] col_in_299,
    input  [511:0] col_in_300,
    input  [511:0] col_in_301,
    input  [511:0] col_in_302,
    input  [511:0] col_in_303,
    input  [511:0] col_in_304,
    input  [511:0] col_in_305,
    input  [511:0] col_in_306,
    input  [511:0] col_in_307,
    input  [511:0] col_in_308,
    input  [511:0] col_in_309,
    input  [511:0] col_in_310,
    input  [511:0] col_in_311,
    input  [511:0] col_in_312,
    input  [511:0] col_in_313,
    input  [511:0] col_in_314,
    input  [511:0] col_in_315,
    input  [511:0] col_in_316,
    input  [511:0] col_in_317,
    input  [511:0] col_in_318,
    input  [511:0] col_in_319,
    input  [511:0] col_in_320,
    input  [511:0] col_in_321,
    input  [511:0] col_in_322,
    input  [511:0] col_in_323,
    input  [511:0] col_in_324,
    input  [511:0] col_in_325,
    input  [511:0] col_in_326,
    input  [511:0] col_in_327,
    input  [511:0] col_in_328,
    input  [511:0] col_in_329,
    input  [511:0] col_in_330,
    input  [511:0] col_in_331,
    input  [511:0] col_in_332,
    input  [511:0] col_in_333,
    input  [511:0] col_in_334,
    input  [511:0] col_in_335,
    input  [511:0] col_in_336,
    input  [511:0] col_in_337,
    input  [511:0] col_in_338,
    input  [511:0] col_in_339,
    input  [511:0] col_in_340,
    input  [511:0] col_in_341,
    input  [511:0] col_in_342,
    input  [511:0] col_in_343,
    input  [511:0] col_in_344,
    input  [511:0] col_in_345,
    input  [511:0] col_in_346,
    input  [511:0] col_in_347,
    input  [511:0] col_in_348,
    input  [511:0] col_in_349,
    input  [511:0] col_in_350,
    input  [511:0] col_in_351,
    input  [511:0] col_in_352,
    input  [511:0] col_in_353,
    input  [511:0] col_in_354,
    input  [511:0] col_in_355,
    input  [511:0] col_in_356,
    input  [511:0] col_in_357,
    input  [511:0] col_in_358,
    input  [511:0] col_in_359,
    input  [511:0] col_in_360,
    input  [511:0] col_in_361,
    input  [511:0] col_in_362,
    input  [511:0] col_in_363,
    input  [511:0] col_in_364,
    input  [511:0] col_in_365,
    input  [511:0] col_in_366,
    input  [511:0] col_in_367,
    input  [511:0] col_in_368,
    input  [511:0] col_in_369,
    input  [511:0] col_in_370,
    input  [511:0] col_in_371,
    input  [511:0] col_in_372,
    input  [511:0] col_in_373,
    input  [511:0] col_in_374,
    input  [511:0] col_in_375,
    input  [511:0] col_in_376,
    input  [511:0] col_in_377,
    input  [511:0] col_in_378,
    input  [511:0] col_in_379,
    input  [511:0] col_in_380,
    input  [511:0] col_in_381,
    input  [511:0] col_in_382,
    input  [511:0] col_in_383,
    input  [511:0] col_in_384,
    input  [511:0] col_in_385,
    input  [511:0] col_in_386,
    input  [511:0] col_in_387,
    input  [511:0] col_in_388,
    input  [511:0] col_in_389,
    input  [511:0] col_in_390,
    input  [511:0] col_in_391,
    input  [511:0] col_in_392,
    input  [511:0] col_in_393,
    input  [511:0] col_in_394,
    input  [511:0] col_in_395,
    input  [511:0] col_in_396,
    input  [511:0] col_in_397,
    input  [511:0] col_in_398,
    input  [511:0] col_in_399,
    input  [511:0] col_in_400,
    input  [511:0] col_in_401,
    input  [511:0] col_in_402,
    input  [511:0] col_in_403,
    input  [511:0] col_in_404,
    input  [511:0] col_in_405,
    input  [511:0] col_in_406,
    input  [511:0] col_in_407,
    input  [511:0] col_in_408,
    input  [511:0] col_in_409,
    input  [511:0] col_in_410,
    input  [511:0] col_in_411,
    input  [511:0] col_in_412,
    input  [511:0] col_in_413,
    input  [511:0] col_in_414,
    input  [511:0] col_in_415,
    input  [511:0] col_in_416,
    input  [511:0] col_in_417,
    input  [511:0] col_in_418,
    input  [511:0] col_in_419,
    input  [511:0] col_in_420,
    input  [511:0] col_in_421,
    input  [511:0] col_in_422,
    input  [511:0] col_in_423,
    input  [511:0] col_in_424,
    input  [511:0] col_in_425,
    input  [511:0] col_in_426,
    input  [511:0] col_in_427,
    input  [511:0] col_in_428,
    input  [511:0] col_in_429,
    input  [511:0] col_in_430,
    input  [511:0] col_in_431,
    input  [511:0] col_in_432,
    input  [511:0] col_in_433,
    input  [511:0] col_in_434,
    input  [511:0] col_in_435,
    input  [511:0] col_in_436,
    input  [511:0] col_in_437,
    input  [511:0] col_in_438,
    input  [511:0] col_in_439,
    input  [511:0] col_in_440,
    input  [511:0] col_in_441,
    input  [511:0] col_in_442,
    input  [511:0] col_in_443,
    input  [511:0] col_in_444,
    input  [511:0] col_in_445,
    input  [511:0] col_in_446,
    input  [511:0] col_in_447,
    input  [511:0] col_in_448,
    input  [511:0] col_in_449,
    input  [511:0] col_in_450,
    input  [511:0] col_in_451,
    input  [511:0] col_in_452,
    input  [511:0] col_in_453,
    input  [511:0] col_in_454,
    input  [511:0] col_in_455,
    input  [511:0] col_in_456,
    input  [511:0] col_in_457,
    input  [511:0] col_in_458,
    input  [511:0] col_in_459,
    input  [511:0] col_in_460,
    input  [511:0] col_in_461,
    input  [511:0] col_in_462,
    input  [511:0] col_in_463,
    input  [511:0] col_in_464,
    input  [511:0] col_in_465,
    input  [511:0] col_in_466,
    input  [511:0] col_in_467,
    input  [511:0] col_in_468,
    input  [511:0] col_in_469,
    input  [511:0] col_in_470,
    input  [511:0] col_in_471,
    input  [511:0] col_in_472,
    input  [511:0] col_in_473,
    input  [511:0] col_in_474,
    input  [511:0] col_in_475,
    input  [511:0] col_in_476,
    input  [511:0] col_in_477,
    input  [511:0] col_in_478,
    input  [511:0] col_in_479,
    input  [511:0] col_in_480,
    input  [511:0] col_in_481,
    input  [511:0] col_in_482,
    input  [511:0] col_in_483,
    input  [511:0] col_in_484,
    input  [511:0] col_in_485,
    input  [511:0] col_in_486,
    input  [511:0] col_in_487,
    input  [511:0] col_in_488,
    input  [511:0] col_in_489,
    input  [511:0] col_in_490,
    input  [511:0] col_in_491,
    input  [511:0] col_in_492,
    input  [511:0] col_in_493,
    input  [511:0] col_in_494,
    input  [511:0] col_in_495,
    input  [511:0] col_in_496,
    input  [511:0] col_in_497,
    input  [511:0] col_in_498,
    input  [511:0] col_in_499,
    input  [511:0] col_in_500,
    input  [511:0] col_in_501,
    input  [511:0] col_in_502,
    input  [511:0] col_in_503,
    input  [511:0] col_in_504,
    input  [511:0] col_in_505,
    input  [511:0] col_in_506,
    input  [511:0] col_in_507,
    input  [511:0] col_in_508,
    input  [511:0] col_in_509,
    input  [511:0] col_in_510,
    input  [511:0] col_in_511,
    input  [511:0] col_in_512,
    input  [511:0] col_in_513,
    input  [511:0] col_in_514,
    input  [511:0] col_in_515,
    input  [511:0] col_in_516,
    input  [511:0] col_in_517,
    input  [511:0] col_in_518,
    input  [511:0] col_in_519,
    input  [511:0] col_in_520,
    input  [511:0] col_in_521,
    input  [511:0] col_in_522,
    input  [511:0] col_in_523,
    input  [511:0] col_in_524,
    input  [511:0] col_in_525,
    input  [511:0] col_in_526,
    input  [511:0] col_in_527,
    input  [511:0] col_in_528,
    input  [511:0] col_in_529,
    input  [511:0] col_in_530,
    input  [511:0] col_in_531,
    input  [511:0] col_in_532,
    input  [511:0] col_in_533,
    input  [511:0] col_in_534,
    input  [511:0] col_in_535,
    input  [511:0] col_in_536,
    input  [511:0] col_in_537,
    input  [511:0] col_in_538,
    input  [511:0] col_in_539,
    input  [511:0] col_in_540,
    input  [511:0] col_in_541,
    input  [511:0] col_in_542,
    input  [511:0] col_in_543,
    input  [511:0] col_in_544,
    input  [511:0] col_in_545,
    input  [511:0] col_in_546,
    input  [511:0] col_in_547,
    input  [511:0] col_in_548,
    input  [511:0] col_in_549,
    input  [511:0] col_in_550,
    input  [511:0] col_in_551,
    input  [511:0] col_in_552,
    input  [511:0] col_in_553,
    input  [511:0] col_in_554,
    input  [511:0] col_in_555,
    input  [511:0] col_in_556,
    input  [511:0] col_in_557,
    input  [511:0] col_in_558,
    input  [511:0] col_in_559,
    input  [511:0] col_in_560,
    input  [511:0] col_in_561,
    input  [511:0] col_in_562,
    input  [511:0] col_in_563,
    input  [511:0] col_in_564,
    input  [511:0] col_in_565,
    input  [511:0] col_in_566,
    input  [511:0] col_in_567,
    input  [511:0] col_in_568,
    input  [511:0] col_in_569,
    input  [511:0] col_in_570,
    input  [511:0] col_in_571,
    input  [511:0] col_in_572,
    input  [511:0] col_in_573,
    input  [511:0] col_in_574,
    input  [511:0] col_in_575,
    input  [511:0] col_in_576,
    input  [511:0] col_in_577,
    input  [511:0] col_in_578,
    input  [511:0] col_in_579,
    input  [511:0] col_in_580,
    input  [511:0] col_in_581,
    input  [511:0] col_in_582,
    input  [511:0] col_in_583,
    input  [511:0] col_in_584,
    input  [511:0] col_in_585,
    input  [511:0] col_in_586,
    input  [511:0] col_in_587,
    input  [511:0] col_in_588,
    input  [511:0] col_in_589,
    input  [511:0] col_in_590,
    input  [511:0] col_in_591,
    input  [511:0] col_in_592,
    input  [511:0] col_in_593,
    input  [511:0] col_in_594,
    input  [511:0] col_in_595,
    input  [511:0] col_in_596,
    input  [511:0] col_in_597,
    input  [511:0] col_in_598,
    input  [511:0] col_in_599,
    input  [511:0] col_in_600,
    input  [511:0] col_in_601,
    input  [511:0] col_in_602,
    input  [511:0] col_in_603,
    input  [511:0] col_in_604,
    input  [511:0] col_in_605,
    input  [511:0] col_in_606,
    input  [511:0] col_in_607,
    input  [511:0] col_in_608,
    input  [511:0] col_in_609,
    input  [511:0] col_in_610,
    input  [511:0] col_in_611,
    input  [511:0] col_in_612,
    input  [511:0] col_in_613,
    input  [511:0] col_in_614,
    input  [511:0] col_in_615,
    input  [511:0] col_in_616,
    input  [511:0] col_in_617,
    input  [511:0] col_in_618,
    input  [511:0] col_in_619,
    input  [511:0] col_in_620,
    input  [511:0] col_in_621,
    input  [511:0] col_in_622,
    input  [511:0] col_in_623,
    input  [511:0] col_in_624,
    input  [511:0] col_in_625,
    input  [511:0] col_in_626,
    input  [511:0] col_in_627,
    input  [511:0] col_in_628,
    input  [511:0] col_in_629,
    input  [511:0] col_in_630,
    input  [511:0] col_in_631,
    input  [511:0] col_in_632,
    input  [511:0] col_in_633,
    input  [511:0] col_in_634,
    input  [511:0] col_in_635,
    input  [511:0] col_in_636,
    input  [511:0] col_in_637,
    input  [511:0] col_in_638,
    input  [511:0] col_in_639,
    input  [511:0] col_in_640,
    input  [511:0] col_in_641,
    input  [511:0] col_in_642,
    input  [511:0] col_in_643,
    input  [511:0] col_in_644,
    input  [511:0] col_in_645,
    input  [511:0] col_in_646,
    input  [511:0] col_in_647,
    input  [511:0] col_in_648,
    input  [511:0] col_in_649,
    input  [511:0] col_in_650,
    input  [511:0] col_in_651,
    input  [511:0] col_in_652,
    input  [511:0] col_in_653,
    input  [511:0] col_in_654,
    input  [511:0] col_in_655,
    input  [511:0] col_in_656,
    input  [511:0] col_in_657,
    input  [511:0] col_in_658,
    input  [511:0] col_in_659,
    input  [511:0] col_in_660,
    input  [511:0] col_in_661,
    input  [511:0] col_in_662,
    input  [511:0] col_in_663,
    input  [511:0] col_in_664,
    input  [511:0] col_in_665,
    input  [511:0] col_in_666,
    input  [511:0] col_in_667,
    input  [511:0] col_in_668,
    input  [511:0] col_in_669,
    input  [511:0] col_in_670,
    input  [511:0] col_in_671,
    input  [511:0] col_in_672,
    input  [511:0] col_in_673,
    input  [511:0] col_in_674,
    input  [511:0] col_in_675,
    input  [511:0] col_in_676,
    input  [511:0] col_in_677,
    input  [511:0] col_in_678,
    input  [511:0] col_in_679,
    input  [511:0] col_in_680,
    input  [511:0] col_in_681,
    input  [511:0] col_in_682,
    input  [511:0] col_in_683,
    input  [511:0] col_in_684,
    input  [511:0] col_in_685,
    input  [511:0] col_in_686,
    input  [511:0] col_in_687,
    input  [511:0] col_in_688,
    input  [511:0] col_in_689,
    input  [511:0] col_in_690,
    input  [511:0] col_in_691,
    input  [511:0] col_in_692,
    input  [511:0] col_in_693,
    input  [511:0] col_in_694,
    input  [511:0] col_in_695,
    input  [511:0] col_in_696,
    input  [511:0] col_in_697,
    input  [511:0] col_in_698,
    input  [511:0] col_in_699,
    input  [511:0] col_in_700,
    input  [511:0] col_in_701,
    input  [511:0] col_in_702,
    input  [511:0] col_in_703,
    input  [511:0] col_in_704,
    input  [511:0] col_in_705,
    input  [511:0] col_in_706,
    input  [511:0] col_in_707,
    input  [511:0] col_in_708,
    input  [511:0] col_in_709,
    input  [511:0] col_in_710,
    input  [511:0] col_in_711,
    input  [511:0] col_in_712,
    input  [511:0] col_in_713,
    input  [511:0] col_in_714,
    input  [511:0] col_in_715,
    input  [511:0] col_in_716,
    input  [511:0] col_in_717,
    input  [511:0] col_in_718,
    input  [511:0] col_in_719,
    input  [511:0] col_in_720,
    input  [511:0] col_in_721,
    input  [511:0] col_in_722,
    input  [511:0] col_in_723,
    input  [511:0] col_in_724,
    input  [511:0] col_in_725,
    input  [511:0] col_in_726,
    input  [511:0] col_in_727,
    input  [511:0] col_in_728,
    input  [511:0] col_in_729,
    input  [511:0] col_in_730,
    input  [511:0] col_in_731,
    input  [511:0] col_in_732,
    input  [511:0] col_in_733,
    input  [511:0] col_in_734,
    input  [511:0] col_in_735,
    input  [511:0] col_in_736,
    input  [511:0] col_in_737,
    input  [511:0] col_in_738,
    input  [511:0] col_in_739,
    input  [511:0] col_in_740,
    input  [511:0] col_in_741,
    input  [511:0] col_in_742,
    input  [511:0] col_in_743,
    input  [511:0] col_in_744,
    input  [511:0] col_in_745,
    input  [511:0] col_in_746,
    input  [511:0] col_in_747,
    input  [511:0] col_in_748,
    input  [511:0] col_in_749,
    input  [511:0] col_in_750,
    input  [511:0] col_in_751,
    input  [511:0] col_in_752,
    input  [511:0] col_in_753,
    input  [511:0] col_in_754,
    input  [511:0] col_in_755,
    input  [511:0] col_in_756,
    input  [511:0] col_in_757,
    input  [511:0] col_in_758,
    input  [511:0] col_in_759,
    input  [511:0] col_in_760,
    input  [511:0] col_in_761,
    input  [511:0] col_in_762,
    input  [511:0] col_in_763,
    input  [511:0] col_in_764,
    input  [511:0] col_in_765,
    input  [511:0] col_in_766,
    input  [511:0] col_in_767,
    input  [511:0] col_in_768,
    input  [511:0] col_in_769,
    input  [511:0] col_in_770,
    input  [511:0] col_in_771,
    input  [511:0] col_in_772,
    input  [511:0] col_in_773,
    input  [511:0] col_in_774,
    input  [511:0] col_in_775,
    input  [511:0] col_in_776,
    input  [511:0] col_in_777,
    input  [511:0] col_in_778,
    input  [511:0] col_in_779,
    input  [511:0] col_in_780,
    input  [511:0] col_in_781,
    input  [511:0] col_in_782,
    input  [511:0] col_in_783,
    input  [511:0] col_in_784,
    input  [511:0] col_in_785,
    input  [511:0] col_in_786,
    input  [511:0] col_in_787,
    input  [511:0] col_in_788,
    input  [511:0] col_in_789,
    input  [511:0] col_in_790,
    input  [511:0] col_in_791,
    input  [511:0] col_in_792,
    input  [511:0] col_in_793,
    input  [511:0] col_in_794,
    input  [511:0] col_in_795,
    input  [511:0] col_in_796,
    input  [511:0] col_in_797,
    input  [511:0] col_in_798,
    input  [511:0] col_in_799,
    input  [511:0] col_in_800,
    input  [511:0] col_in_801,
    input  [511:0] col_in_802,
    input  [511:0] col_in_803,
    input  [511:0] col_in_804,
    input  [511:0] col_in_805,
    input  [511:0] col_in_806,
    input  [511:0] col_in_807,
    input  [511:0] col_in_808,
    input  [511:0] col_in_809,
    input  [511:0] col_in_810,
    input  [511:0] col_in_811,
    input  [511:0] col_in_812,
    input  [511:0] col_in_813,
    input  [511:0] col_in_814,
    input  [511:0] col_in_815,
    input  [511:0] col_in_816,
    input  [511:0] col_in_817,
    input  [511:0] col_in_818,
    input  [511:0] col_in_819,
    input  [511:0] col_in_820,
    input  [511:0] col_in_821,
    input  [511:0] col_in_822,
    input  [511:0] col_in_823,
    input  [511:0] col_in_824,
    input  [511:0] col_in_825,
    input  [511:0] col_in_826,
    input  [511:0] col_in_827,
    input  [511:0] col_in_828,
    input  [511:0] col_in_829,
    input  [511:0] col_in_830,
    input  [511:0] col_in_831,
    input  [511:0] col_in_832,
    input  [511:0] col_in_833,
    input  [511:0] col_in_834,
    input  [511:0] col_in_835,
    input  [511:0] col_in_836,
    input  [511:0] col_in_837,
    input  [511:0] col_in_838,
    input  [511:0] col_in_839,
    input  [511:0] col_in_840,
    input  [511:0] col_in_841,
    input  [511:0] col_in_842,
    input  [511:0] col_in_843,
    input  [511:0] col_in_844,
    input  [511:0] col_in_845,
    input  [511:0] col_in_846,
    input  [511:0] col_in_847,
    input  [511:0] col_in_848,
    input  [511:0] col_in_849,
    input  [511:0] col_in_850,
    input  [511:0] col_in_851,
    input  [511:0] col_in_852,
    input  [511:0] col_in_853,
    input  [511:0] col_in_854,
    input  [511:0] col_in_855,
    input  [511:0] col_in_856,
    input  [511:0] col_in_857,
    input  [511:0] col_in_858,
    input  [511:0] col_in_859,
    input  [511:0] col_in_860,
    input  [511:0] col_in_861,
    input  [511:0] col_in_862,
    input  [511:0] col_in_863,
    input  [511:0] col_in_864,
    input  [511:0] col_in_865,
    input  [511:0] col_in_866,
    input  [511:0] col_in_867,
    input  [511:0] col_in_868,
    input  [511:0] col_in_869,
    input  [511:0] col_in_870,
    input  [511:0] col_in_871,
    input  [511:0] col_in_872,
    input  [511:0] col_in_873,
    input  [511:0] col_in_874,
    input  [511:0] col_in_875,
    input  [511:0] col_in_876,
    input  [511:0] col_in_877,
    input  [511:0] col_in_878,
    input  [511:0] col_in_879,
    input  [511:0] col_in_880,
    input  [511:0] col_in_881,
    input  [511:0] col_in_882,
    input  [511:0] col_in_883,
    input  [511:0] col_in_884,
    input  [511:0] col_in_885,
    input  [511:0] col_in_886,
    input  [511:0] col_in_887,
    input  [511:0] col_in_888,
    input  [511:0] col_in_889,
    input  [511:0] col_in_890,
    input  [511:0] col_in_891,
    input  [511:0] col_in_892,
    input  [511:0] col_in_893,
    input  [511:0] col_in_894,
    input  [511:0] col_in_895,
    input  [511:0] col_in_896,
    input  [511:0] col_in_897,
    input  [511:0] col_in_898,
    input  [511:0] col_in_899,
    input  [511:0] col_in_900,
    input  [511:0] col_in_901,
    input  [511:0] col_in_902,
    input  [511:0] col_in_903,
    input  [511:0] col_in_904,
    input  [511:0] col_in_905,
    input  [511:0] col_in_906,
    input  [511:0] col_in_907,
    input  [511:0] col_in_908,
    input  [511:0] col_in_909,
    input  [511:0] col_in_910,
    input  [511:0] col_in_911,
    input  [511:0] col_in_912,
    input  [511:0] col_in_913,
    input  [511:0] col_in_914,
    input  [511:0] col_in_915,
    input  [511:0] col_in_916,
    input  [511:0] col_in_917,
    input  [511:0] col_in_918,
    input  [511:0] col_in_919,
    input  [511:0] col_in_920,
    input  [511:0] col_in_921,
    input  [511:0] col_in_922,
    input  [511:0] col_in_923,
    input  [511:0] col_in_924,
    input  [511:0] col_in_925,
    input  [511:0] col_in_926,
    input  [511:0] col_in_927,
    input  [511:0] col_in_928,
    input  [511:0] col_in_929,
    input  [511:0] col_in_930,
    input  [511:0] col_in_931,
    input  [511:0] col_in_932,
    input  [511:0] col_in_933,
    input  [511:0] col_in_934,
    input  [511:0] col_in_935,
    input  [511:0] col_in_936,
    input  [511:0] col_in_937,
    input  [511:0] col_in_938,
    input  [511:0] col_in_939,
    input  [511:0] col_in_940,
    input  [511:0] col_in_941,
    input  [511:0] col_in_942,
    input  [511:0] col_in_943,
    input  [511:0] col_in_944,
    input  [511:0] col_in_945,
    input  [511:0] col_in_946,
    input  [511:0] col_in_947,
    input  [511:0] col_in_948,
    input  [511:0] col_in_949,
    input  [511:0] col_in_950,
    input  [511:0] col_in_951,
    input  [511:0] col_in_952,
    input  [511:0] col_in_953,
    input  [511:0] col_in_954,
    input  [511:0] col_in_955,
    input  [511:0] col_in_956,
    input  [511:0] col_in_957,
    input  [511:0] col_in_958,
    input  [511:0] col_in_959,
    input  [511:0] col_in_960,
    input  [511:0] col_in_961,
    input  [511:0] col_in_962,
    input  [511:0] col_in_963,
    input  [511:0] col_in_964,
    input  [511:0] col_in_965,
    input  [511:0] col_in_966,
    input  [511:0] col_in_967,
    input  [511:0] col_in_968,
    input  [511:0] col_in_969,
    input  [511:0] col_in_970,
    input  [511:0] col_in_971,
    input  [511:0] col_in_972,
    input  [511:0] col_in_973,
    input  [511:0] col_in_974,
    input  [511:0] col_in_975,
    input  [511:0] col_in_976,
    input  [511:0] col_in_977,
    input  [511:0] col_in_978,
    input  [511:0] col_in_979,
    input  [511:0] col_in_980,
    input  [511:0] col_in_981,
    input  [511:0] col_in_982,
    input  [511:0] col_in_983,
    input  [511:0] col_in_984,
    input  [511:0] col_in_985,
    input  [511:0] col_in_986,
    input  [511:0] col_in_987,
    input  [511:0] col_in_988,
    input  [511:0] col_in_989,
    input  [511:0] col_in_990,
    input  [511:0] col_in_991,
    input  [511:0] col_in_992,
    input  [511:0] col_in_993,
    input  [511:0] col_in_994,
    input  [511:0] col_in_995,
    input  [511:0] col_in_996,
    input  [511:0] col_in_997,
    input  [511:0] col_in_998,
    input  [511:0] col_in_999,
    input  [511:0] col_in_1000,
    input  [511:0] col_in_1001,
    input  [511:0] col_in_1002,
    input  [511:0] col_in_1003,
    input  [511:0] col_in_1004,
    input  [511:0] col_in_1005,
    input  [511:0] col_in_1006,
    input  [511:0] col_in_1007,
    input  [511:0] col_in_1008,
    input  [511:0] col_in_1009,
    input  [511:0] col_in_1010,
    input  [511:0] col_in_1011,
    input  [511:0] col_in_1012,
    input  [511:0] col_in_1013,
    input  [511:0] col_in_1014,
    input  [511:0] col_in_1015,
    input  [511:0] col_in_1016,
    input  [511:0] col_in_1017,
    input  [511:0] col_in_1018,
    input  [511:0] col_in_1019,
    input  [511:0] col_in_1020,
    input  [511:0] col_in_1021,
    input  [511:0] col_in_1022,
    input  [511:0] col_in_1023,

    output [1032:0] row_out_0,
    output [1032:0] row_out_1
);



// compressor_array_512_2_1024 Outputs
wire  [1:0]  col_out_0;
wire  [1:0]  col_out_1;
wire  [1:0]  col_out_2;
wire  [1:0]  col_out_3;
wire  [1:0]  col_out_4;
wire  [1:0]  col_out_5;
wire  [1:0]  col_out_6;
wire  [1:0]  col_out_7;
wire  [1:0]  col_out_8;
wire  [1:0]  col_out_9;
wire  [1:0]  col_out_10;
wire  [1:0]  col_out_11;
wire  [1:0]  col_out_12;
wire  [1:0]  col_out_13;
wire  [1:0]  col_out_14;
wire  [1:0]  col_out_15;
wire  [1:0]  col_out_16;
wire  [1:0]  col_out_17;
wire  [1:0]  col_out_18;
wire  [1:0]  col_out_19;
wire  [1:0]  col_out_20;
wire  [1:0]  col_out_21;
wire  [1:0]  col_out_22;
wire  [1:0]  col_out_23;
wire  [1:0]  col_out_24;
wire  [1:0]  col_out_25;
wire  [1:0]  col_out_26;
wire  [1:0]  col_out_27;
wire  [1:0]  col_out_28;
wire  [1:0]  col_out_29;
wire  [1:0]  col_out_30;
wire  [1:0]  col_out_31;
wire  [1:0]  col_out_32;
wire  [1:0]  col_out_33;
wire  [1:0]  col_out_34;
wire  [1:0]  col_out_35;
wire  [1:0]  col_out_36;
wire  [1:0]  col_out_37;
wire  [1:0]  col_out_38;
wire  [1:0]  col_out_39;
wire  [1:0]  col_out_40;
wire  [1:0]  col_out_41;
wire  [1:0]  col_out_42;
wire  [1:0]  col_out_43;
wire  [1:0]  col_out_44;
wire  [1:0]  col_out_45;
wire  [1:0]  col_out_46;
wire  [1:0]  col_out_47;
wire  [1:0]  col_out_48;
wire  [1:0]  col_out_49;
wire  [1:0]  col_out_50;
wire  [1:0]  col_out_51;
wire  [1:0]  col_out_52;
wire  [1:0]  col_out_53;
wire  [1:0]  col_out_54;
wire  [1:0]  col_out_55;
wire  [1:0]  col_out_56;
wire  [1:0]  col_out_57;
wire  [1:0]  col_out_58;
wire  [1:0]  col_out_59;
wire  [1:0]  col_out_60;
wire  [1:0]  col_out_61;
wire  [1:0]  col_out_62;
wire  [1:0]  col_out_63;
wire  [1:0]  col_out_64;
wire  [1:0]  col_out_65;
wire  [1:0]  col_out_66;
wire  [1:0]  col_out_67;
wire  [1:0]  col_out_68;
wire  [1:0]  col_out_69;
wire  [1:0]  col_out_70;
wire  [1:0]  col_out_71;
wire  [1:0]  col_out_72;
wire  [1:0]  col_out_73;
wire  [1:0]  col_out_74;
wire  [1:0]  col_out_75;
wire  [1:0]  col_out_76;
wire  [1:0]  col_out_77;
wire  [1:0]  col_out_78;
wire  [1:0]  col_out_79;
wire  [1:0]  col_out_80;
wire  [1:0]  col_out_81;
wire  [1:0]  col_out_82;
wire  [1:0]  col_out_83;
wire  [1:0]  col_out_84;
wire  [1:0]  col_out_85;
wire  [1:0]  col_out_86;
wire  [1:0]  col_out_87;
wire  [1:0]  col_out_88;
wire  [1:0]  col_out_89;
wire  [1:0]  col_out_90;
wire  [1:0]  col_out_91;
wire  [1:0]  col_out_92;
wire  [1:0]  col_out_93;
wire  [1:0]  col_out_94;
wire  [1:0]  col_out_95;
wire  [1:0]  col_out_96;
wire  [1:0]  col_out_97;
wire  [1:0]  col_out_98;
wire  [1:0]  col_out_99;
wire  [1:0]  col_out_100;
wire  [1:0]  col_out_101;
wire  [1:0]  col_out_102;
wire  [1:0]  col_out_103;
wire  [1:0]  col_out_104;
wire  [1:0]  col_out_105;
wire  [1:0]  col_out_106;
wire  [1:0]  col_out_107;
wire  [1:0]  col_out_108;
wire  [1:0]  col_out_109;
wire  [1:0]  col_out_110;
wire  [1:0]  col_out_111;
wire  [1:0]  col_out_112;
wire  [1:0]  col_out_113;
wire  [1:0]  col_out_114;
wire  [1:0]  col_out_115;
wire  [1:0]  col_out_116;
wire  [1:0]  col_out_117;
wire  [1:0]  col_out_118;
wire  [1:0]  col_out_119;
wire  [1:0]  col_out_120;
wire  [1:0]  col_out_121;
wire  [1:0]  col_out_122;
wire  [1:0]  col_out_123;
wire  [1:0]  col_out_124;
wire  [1:0]  col_out_125;
wire  [1:0]  col_out_126;
wire  [1:0]  col_out_127;
wire  [1:0]  col_out_128;
wire  [1:0]  col_out_129;
wire  [1:0]  col_out_130;
wire  [1:0]  col_out_131;
wire  [1:0]  col_out_132;
wire  [1:0]  col_out_133;
wire  [1:0]  col_out_134;
wire  [1:0]  col_out_135;
wire  [1:0]  col_out_136;
wire  [1:0]  col_out_137;
wire  [1:0]  col_out_138;
wire  [1:0]  col_out_139;
wire  [1:0]  col_out_140;
wire  [1:0]  col_out_141;
wire  [1:0]  col_out_142;
wire  [1:0]  col_out_143;
wire  [1:0]  col_out_144;
wire  [1:0]  col_out_145;
wire  [1:0]  col_out_146;
wire  [1:0]  col_out_147;
wire  [1:0]  col_out_148;
wire  [1:0]  col_out_149;
wire  [1:0]  col_out_150;
wire  [1:0]  col_out_151;
wire  [1:0]  col_out_152;
wire  [1:0]  col_out_153;
wire  [1:0]  col_out_154;
wire  [1:0]  col_out_155;
wire  [1:0]  col_out_156;
wire  [1:0]  col_out_157;
wire  [1:0]  col_out_158;
wire  [1:0]  col_out_159;
wire  [1:0]  col_out_160;
wire  [1:0]  col_out_161;
wire  [1:0]  col_out_162;
wire  [1:0]  col_out_163;
wire  [1:0]  col_out_164;
wire  [1:0]  col_out_165;
wire  [1:0]  col_out_166;
wire  [1:0]  col_out_167;
wire  [1:0]  col_out_168;
wire  [1:0]  col_out_169;
wire  [1:0]  col_out_170;
wire  [1:0]  col_out_171;
wire  [1:0]  col_out_172;
wire  [1:0]  col_out_173;
wire  [1:0]  col_out_174;
wire  [1:0]  col_out_175;
wire  [1:0]  col_out_176;
wire  [1:0]  col_out_177;
wire  [1:0]  col_out_178;
wire  [1:0]  col_out_179;
wire  [1:0]  col_out_180;
wire  [1:0]  col_out_181;
wire  [1:0]  col_out_182;
wire  [1:0]  col_out_183;
wire  [1:0]  col_out_184;
wire  [1:0]  col_out_185;
wire  [1:0]  col_out_186;
wire  [1:0]  col_out_187;
wire  [1:0]  col_out_188;
wire  [1:0]  col_out_189;
wire  [1:0]  col_out_190;
wire  [1:0]  col_out_191;
wire  [1:0]  col_out_192;
wire  [1:0]  col_out_193;
wire  [1:0]  col_out_194;
wire  [1:0]  col_out_195;
wire  [1:0]  col_out_196;
wire  [1:0]  col_out_197;
wire  [1:0]  col_out_198;
wire  [1:0]  col_out_199;
wire  [1:0]  col_out_200;
wire  [1:0]  col_out_201;
wire  [1:0]  col_out_202;
wire  [1:0]  col_out_203;
wire  [1:0]  col_out_204;
wire  [1:0]  col_out_205;
wire  [1:0]  col_out_206;
wire  [1:0]  col_out_207;
wire  [1:0]  col_out_208;
wire  [1:0]  col_out_209;
wire  [1:0]  col_out_210;
wire  [1:0]  col_out_211;
wire  [1:0]  col_out_212;
wire  [1:0]  col_out_213;
wire  [1:0]  col_out_214;
wire  [1:0]  col_out_215;
wire  [1:0]  col_out_216;
wire  [1:0]  col_out_217;
wire  [1:0]  col_out_218;
wire  [1:0]  col_out_219;
wire  [1:0]  col_out_220;
wire  [1:0]  col_out_221;
wire  [1:0]  col_out_222;
wire  [1:0]  col_out_223;
wire  [1:0]  col_out_224;
wire  [1:0]  col_out_225;
wire  [1:0]  col_out_226;
wire  [1:0]  col_out_227;
wire  [1:0]  col_out_228;
wire  [1:0]  col_out_229;
wire  [1:0]  col_out_230;
wire  [1:0]  col_out_231;
wire  [1:0]  col_out_232;
wire  [1:0]  col_out_233;
wire  [1:0]  col_out_234;
wire  [1:0]  col_out_235;
wire  [1:0]  col_out_236;
wire  [1:0]  col_out_237;
wire  [1:0]  col_out_238;
wire  [1:0]  col_out_239;
wire  [1:0]  col_out_240;
wire  [1:0]  col_out_241;
wire  [1:0]  col_out_242;
wire  [1:0]  col_out_243;
wire  [1:0]  col_out_244;
wire  [1:0]  col_out_245;
wire  [1:0]  col_out_246;
wire  [1:0]  col_out_247;
wire  [1:0]  col_out_248;
wire  [1:0]  col_out_249;
wire  [1:0]  col_out_250;
wire  [1:0]  col_out_251;
wire  [1:0]  col_out_252;
wire  [1:0]  col_out_253;
wire  [1:0]  col_out_254;
wire  [1:0]  col_out_255;
wire  [1:0]  col_out_256;
wire  [1:0]  col_out_257;
wire  [1:0]  col_out_258;
wire  [1:0]  col_out_259;
wire  [1:0]  col_out_260;
wire  [1:0]  col_out_261;
wire  [1:0]  col_out_262;
wire  [1:0]  col_out_263;
wire  [1:0]  col_out_264;
wire  [1:0]  col_out_265;
wire  [1:0]  col_out_266;
wire  [1:0]  col_out_267;
wire  [1:0]  col_out_268;
wire  [1:0]  col_out_269;
wire  [1:0]  col_out_270;
wire  [1:0]  col_out_271;
wire  [1:0]  col_out_272;
wire  [1:0]  col_out_273;
wire  [1:0]  col_out_274;
wire  [1:0]  col_out_275;
wire  [1:0]  col_out_276;
wire  [1:0]  col_out_277;
wire  [1:0]  col_out_278;
wire  [1:0]  col_out_279;
wire  [1:0]  col_out_280;
wire  [1:0]  col_out_281;
wire  [1:0]  col_out_282;
wire  [1:0]  col_out_283;
wire  [1:0]  col_out_284;
wire  [1:0]  col_out_285;
wire  [1:0]  col_out_286;
wire  [1:0]  col_out_287;
wire  [1:0]  col_out_288;
wire  [1:0]  col_out_289;
wire  [1:0]  col_out_290;
wire  [1:0]  col_out_291;
wire  [1:0]  col_out_292;
wire  [1:0]  col_out_293;
wire  [1:0]  col_out_294;
wire  [1:0]  col_out_295;
wire  [1:0]  col_out_296;
wire  [1:0]  col_out_297;
wire  [1:0]  col_out_298;
wire  [1:0]  col_out_299;
wire  [1:0]  col_out_300;
wire  [1:0]  col_out_301;
wire  [1:0]  col_out_302;
wire  [1:0]  col_out_303;
wire  [1:0]  col_out_304;
wire  [1:0]  col_out_305;
wire  [1:0]  col_out_306;
wire  [1:0]  col_out_307;
wire  [1:0]  col_out_308;
wire  [1:0]  col_out_309;
wire  [1:0]  col_out_310;
wire  [1:0]  col_out_311;
wire  [1:0]  col_out_312;
wire  [1:0]  col_out_313;
wire  [1:0]  col_out_314;
wire  [1:0]  col_out_315;
wire  [1:0]  col_out_316;
wire  [1:0]  col_out_317;
wire  [1:0]  col_out_318;
wire  [1:0]  col_out_319;
wire  [1:0]  col_out_320;
wire  [1:0]  col_out_321;
wire  [1:0]  col_out_322;
wire  [1:0]  col_out_323;
wire  [1:0]  col_out_324;
wire  [1:0]  col_out_325;
wire  [1:0]  col_out_326;
wire  [1:0]  col_out_327;
wire  [1:0]  col_out_328;
wire  [1:0]  col_out_329;
wire  [1:0]  col_out_330;
wire  [1:0]  col_out_331;
wire  [1:0]  col_out_332;
wire  [1:0]  col_out_333;
wire  [1:0]  col_out_334;
wire  [1:0]  col_out_335;
wire  [1:0]  col_out_336;
wire  [1:0]  col_out_337;
wire  [1:0]  col_out_338;
wire  [1:0]  col_out_339;
wire  [1:0]  col_out_340;
wire  [1:0]  col_out_341;
wire  [1:0]  col_out_342;
wire  [1:0]  col_out_343;
wire  [1:0]  col_out_344;
wire  [1:0]  col_out_345;
wire  [1:0]  col_out_346;
wire  [1:0]  col_out_347;
wire  [1:0]  col_out_348;
wire  [1:0]  col_out_349;
wire  [1:0]  col_out_350;
wire  [1:0]  col_out_351;
wire  [1:0]  col_out_352;
wire  [1:0]  col_out_353;
wire  [1:0]  col_out_354;
wire  [1:0]  col_out_355;
wire  [1:0]  col_out_356;
wire  [1:0]  col_out_357;
wire  [1:0]  col_out_358;
wire  [1:0]  col_out_359;
wire  [1:0]  col_out_360;
wire  [1:0]  col_out_361;
wire  [1:0]  col_out_362;
wire  [1:0]  col_out_363;
wire  [1:0]  col_out_364;
wire  [1:0]  col_out_365;
wire  [1:0]  col_out_366;
wire  [1:0]  col_out_367;
wire  [1:0]  col_out_368;
wire  [1:0]  col_out_369;
wire  [1:0]  col_out_370;
wire  [1:0]  col_out_371;
wire  [1:0]  col_out_372;
wire  [1:0]  col_out_373;
wire  [1:0]  col_out_374;
wire  [1:0]  col_out_375;
wire  [1:0]  col_out_376;
wire  [1:0]  col_out_377;
wire  [1:0]  col_out_378;
wire  [1:0]  col_out_379;
wire  [1:0]  col_out_380;
wire  [1:0]  col_out_381;
wire  [1:0]  col_out_382;
wire  [1:0]  col_out_383;
wire  [1:0]  col_out_384;
wire  [1:0]  col_out_385;
wire  [1:0]  col_out_386;
wire  [1:0]  col_out_387;
wire  [1:0]  col_out_388;
wire  [1:0]  col_out_389;
wire  [1:0]  col_out_390;
wire  [1:0]  col_out_391;
wire  [1:0]  col_out_392;
wire  [1:0]  col_out_393;
wire  [1:0]  col_out_394;
wire  [1:0]  col_out_395;
wire  [1:0]  col_out_396;
wire  [1:0]  col_out_397;
wire  [1:0]  col_out_398;
wire  [1:0]  col_out_399;
wire  [1:0]  col_out_400;
wire  [1:0]  col_out_401;
wire  [1:0]  col_out_402;
wire  [1:0]  col_out_403;
wire  [1:0]  col_out_404;
wire  [1:0]  col_out_405;
wire  [1:0]  col_out_406;
wire  [1:0]  col_out_407;
wire  [1:0]  col_out_408;
wire  [1:0]  col_out_409;
wire  [1:0]  col_out_410;
wire  [1:0]  col_out_411;
wire  [1:0]  col_out_412;
wire  [1:0]  col_out_413;
wire  [1:0]  col_out_414;
wire  [1:0]  col_out_415;
wire  [1:0]  col_out_416;
wire  [1:0]  col_out_417;
wire  [1:0]  col_out_418;
wire  [1:0]  col_out_419;
wire  [1:0]  col_out_420;
wire  [1:0]  col_out_421;
wire  [1:0]  col_out_422;
wire  [1:0]  col_out_423;
wire  [1:0]  col_out_424;
wire  [1:0]  col_out_425;
wire  [1:0]  col_out_426;
wire  [1:0]  col_out_427;
wire  [1:0]  col_out_428;
wire  [1:0]  col_out_429;
wire  [1:0]  col_out_430;
wire  [1:0]  col_out_431;
wire  [1:0]  col_out_432;
wire  [1:0]  col_out_433;
wire  [1:0]  col_out_434;
wire  [1:0]  col_out_435;
wire  [1:0]  col_out_436;
wire  [1:0]  col_out_437;
wire  [1:0]  col_out_438;
wire  [1:0]  col_out_439;
wire  [1:0]  col_out_440;
wire  [1:0]  col_out_441;
wire  [1:0]  col_out_442;
wire  [1:0]  col_out_443;
wire  [1:0]  col_out_444;
wire  [1:0]  col_out_445;
wire  [1:0]  col_out_446;
wire  [1:0]  col_out_447;
wire  [1:0]  col_out_448;
wire  [1:0]  col_out_449;
wire  [1:0]  col_out_450;
wire  [1:0]  col_out_451;
wire  [1:0]  col_out_452;
wire  [1:0]  col_out_453;
wire  [1:0]  col_out_454;
wire  [1:0]  col_out_455;
wire  [1:0]  col_out_456;
wire  [1:0]  col_out_457;
wire  [1:0]  col_out_458;
wire  [1:0]  col_out_459;
wire  [1:0]  col_out_460;
wire  [1:0]  col_out_461;
wire  [1:0]  col_out_462;
wire  [1:0]  col_out_463;
wire  [1:0]  col_out_464;
wire  [1:0]  col_out_465;
wire  [1:0]  col_out_466;
wire  [1:0]  col_out_467;
wire  [1:0]  col_out_468;
wire  [1:0]  col_out_469;
wire  [1:0]  col_out_470;
wire  [1:0]  col_out_471;
wire  [1:0]  col_out_472;
wire  [1:0]  col_out_473;
wire  [1:0]  col_out_474;
wire  [1:0]  col_out_475;
wire  [1:0]  col_out_476;
wire  [1:0]  col_out_477;
wire  [1:0]  col_out_478;
wire  [1:0]  col_out_479;
wire  [1:0]  col_out_480;
wire  [1:0]  col_out_481;
wire  [1:0]  col_out_482;
wire  [1:0]  col_out_483;
wire  [1:0]  col_out_484;
wire  [1:0]  col_out_485;
wire  [1:0]  col_out_486;
wire  [1:0]  col_out_487;
wire  [1:0]  col_out_488;
wire  [1:0]  col_out_489;
wire  [1:0]  col_out_490;
wire  [1:0]  col_out_491;
wire  [1:0]  col_out_492;
wire  [1:0]  col_out_493;
wire  [1:0]  col_out_494;
wire  [1:0]  col_out_495;
wire  [1:0]  col_out_496;
wire  [1:0]  col_out_497;
wire  [1:0]  col_out_498;
wire  [1:0]  col_out_499;
wire  [1:0]  col_out_500;
wire  [1:0]  col_out_501;
wire  [1:0]  col_out_502;
wire  [1:0]  col_out_503;
wire  [1:0]  col_out_504;
wire  [1:0]  col_out_505;
wire  [1:0]  col_out_506;
wire  [1:0]  col_out_507;
wire  [1:0]  col_out_508;
wire  [1:0]  col_out_509;
wire  [1:0]  col_out_510;
wire  [1:0]  col_out_511;
wire  [1:0]  col_out_512;
wire  [1:0]  col_out_513;
wire  [1:0]  col_out_514;
wire  [1:0]  col_out_515;
wire  [1:0]  col_out_516;
wire  [1:0]  col_out_517;
wire  [1:0]  col_out_518;
wire  [1:0]  col_out_519;
wire  [1:0]  col_out_520;
wire  [1:0]  col_out_521;
wire  [1:0]  col_out_522;
wire  [1:0]  col_out_523;
wire  [1:0]  col_out_524;
wire  [1:0]  col_out_525;
wire  [1:0]  col_out_526;
wire  [1:0]  col_out_527;
wire  [1:0]  col_out_528;
wire  [1:0]  col_out_529;
wire  [1:0]  col_out_530;
wire  [1:0]  col_out_531;
wire  [1:0]  col_out_532;
wire  [1:0]  col_out_533;
wire  [1:0]  col_out_534;
wire  [1:0]  col_out_535;
wire  [1:0]  col_out_536;
wire  [1:0]  col_out_537;
wire  [1:0]  col_out_538;
wire  [1:0]  col_out_539;
wire  [1:0]  col_out_540;
wire  [1:0]  col_out_541;
wire  [1:0]  col_out_542;
wire  [1:0]  col_out_543;
wire  [1:0]  col_out_544;
wire  [1:0]  col_out_545;
wire  [1:0]  col_out_546;
wire  [1:0]  col_out_547;
wire  [1:0]  col_out_548;
wire  [1:0]  col_out_549;
wire  [1:0]  col_out_550;
wire  [1:0]  col_out_551;
wire  [1:0]  col_out_552;
wire  [1:0]  col_out_553;
wire  [1:0]  col_out_554;
wire  [1:0]  col_out_555;
wire  [1:0]  col_out_556;
wire  [1:0]  col_out_557;
wire  [1:0]  col_out_558;
wire  [1:0]  col_out_559;
wire  [1:0]  col_out_560;
wire  [1:0]  col_out_561;
wire  [1:0]  col_out_562;
wire  [1:0]  col_out_563;
wire  [1:0]  col_out_564;
wire  [1:0]  col_out_565;
wire  [1:0]  col_out_566;
wire  [1:0]  col_out_567;
wire  [1:0]  col_out_568;
wire  [1:0]  col_out_569;
wire  [1:0]  col_out_570;
wire  [1:0]  col_out_571;
wire  [1:0]  col_out_572;
wire  [1:0]  col_out_573;
wire  [1:0]  col_out_574;
wire  [1:0]  col_out_575;
wire  [1:0]  col_out_576;
wire  [1:0]  col_out_577;
wire  [1:0]  col_out_578;
wire  [1:0]  col_out_579;
wire  [1:0]  col_out_580;
wire  [1:0]  col_out_581;
wire  [1:0]  col_out_582;
wire  [1:0]  col_out_583;
wire  [1:0]  col_out_584;
wire  [1:0]  col_out_585;
wire  [1:0]  col_out_586;
wire  [1:0]  col_out_587;
wire  [1:0]  col_out_588;
wire  [1:0]  col_out_589;
wire  [1:0]  col_out_590;
wire  [1:0]  col_out_591;
wire  [1:0]  col_out_592;
wire  [1:0]  col_out_593;
wire  [1:0]  col_out_594;
wire  [1:0]  col_out_595;
wire  [1:0]  col_out_596;
wire  [1:0]  col_out_597;
wire  [1:0]  col_out_598;
wire  [1:0]  col_out_599;
wire  [1:0]  col_out_600;
wire  [1:0]  col_out_601;
wire  [1:0]  col_out_602;
wire  [1:0]  col_out_603;
wire  [1:0]  col_out_604;
wire  [1:0]  col_out_605;
wire  [1:0]  col_out_606;
wire  [1:0]  col_out_607;
wire  [1:0]  col_out_608;
wire  [1:0]  col_out_609;
wire  [1:0]  col_out_610;
wire  [1:0]  col_out_611;
wire  [1:0]  col_out_612;
wire  [1:0]  col_out_613;
wire  [1:0]  col_out_614;
wire  [1:0]  col_out_615;
wire  [1:0]  col_out_616;
wire  [1:0]  col_out_617;
wire  [1:0]  col_out_618;
wire  [1:0]  col_out_619;
wire  [1:0]  col_out_620;
wire  [1:0]  col_out_621;
wire  [1:0]  col_out_622;
wire  [1:0]  col_out_623;
wire  [1:0]  col_out_624;
wire  [1:0]  col_out_625;
wire  [1:0]  col_out_626;
wire  [1:0]  col_out_627;
wire  [1:0]  col_out_628;
wire  [1:0]  col_out_629;
wire  [1:0]  col_out_630;
wire  [1:0]  col_out_631;
wire  [1:0]  col_out_632;
wire  [1:0]  col_out_633;
wire  [1:0]  col_out_634;
wire  [1:0]  col_out_635;
wire  [1:0]  col_out_636;
wire  [1:0]  col_out_637;
wire  [1:0]  col_out_638;
wire  [1:0]  col_out_639;
wire  [1:0]  col_out_640;
wire  [1:0]  col_out_641;
wire  [1:0]  col_out_642;
wire  [1:0]  col_out_643;
wire  [1:0]  col_out_644;
wire  [1:0]  col_out_645;
wire  [1:0]  col_out_646;
wire  [1:0]  col_out_647;
wire  [1:0]  col_out_648;
wire  [1:0]  col_out_649;
wire  [1:0]  col_out_650;
wire  [1:0]  col_out_651;
wire  [1:0]  col_out_652;
wire  [1:0]  col_out_653;
wire  [1:0]  col_out_654;
wire  [1:0]  col_out_655;
wire  [1:0]  col_out_656;
wire  [1:0]  col_out_657;
wire  [1:0]  col_out_658;
wire  [1:0]  col_out_659;
wire  [1:0]  col_out_660;
wire  [1:0]  col_out_661;
wire  [1:0]  col_out_662;
wire  [1:0]  col_out_663;
wire  [1:0]  col_out_664;
wire  [1:0]  col_out_665;
wire  [1:0]  col_out_666;
wire  [1:0]  col_out_667;
wire  [1:0]  col_out_668;
wire  [1:0]  col_out_669;
wire  [1:0]  col_out_670;
wire  [1:0]  col_out_671;
wire  [1:0]  col_out_672;
wire  [1:0]  col_out_673;
wire  [1:0]  col_out_674;
wire  [1:0]  col_out_675;
wire  [1:0]  col_out_676;
wire  [1:0]  col_out_677;
wire  [1:0]  col_out_678;
wire  [1:0]  col_out_679;
wire  [1:0]  col_out_680;
wire  [1:0]  col_out_681;
wire  [1:0]  col_out_682;
wire  [1:0]  col_out_683;
wire  [1:0]  col_out_684;
wire  [1:0]  col_out_685;
wire  [1:0]  col_out_686;
wire  [1:0]  col_out_687;
wire  [1:0]  col_out_688;
wire  [1:0]  col_out_689;
wire  [1:0]  col_out_690;
wire  [1:0]  col_out_691;
wire  [1:0]  col_out_692;
wire  [1:0]  col_out_693;
wire  [1:0]  col_out_694;
wire  [1:0]  col_out_695;
wire  [1:0]  col_out_696;
wire  [1:0]  col_out_697;
wire  [1:0]  col_out_698;
wire  [1:0]  col_out_699;
wire  [1:0]  col_out_700;
wire  [1:0]  col_out_701;
wire  [1:0]  col_out_702;
wire  [1:0]  col_out_703;
wire  [1:0]  col_out_704;
wire  [1:0]  col_out_705;
wire  [1:0]  col_out_706;
wire  [1:0]  col_out_707;
wire  [1:0]  col_out_708;
wire  [1:0]  col_out_709;
wire  [1:0]  col_out_710;
wire  [1:0]  col_out_711;
wire  [1:0]  col_out_712;
wire  [1:0]  col_out_713;
wire  [1:0]  col_out_714;
wire  [1:0]  col_out_715;
wire  [1:0]  col_out_716;
wire  [1:0]  col_out_717;
wire  [1:0]  col_out_718;
wire  [1:0]  col_out_719;
wire  [1:0]  col_out_720;
wire  [1:0]  col_out_721;
wire  [1:0]  col_out_722;
wire  [1:0]  col_out_723;
wire  [1:0]  col_out_724;
wire  [1:0]  col_out_725;
wire  [1:0]  col_out_726;
wire  [1:0]  col_out_727;
wire  [1:0]  col_out_728;
wire  [1:0]  col_out_729;
wire  [1:0]  col_out_730;
wire  [1:0]  col_out_731;
wire  [1:0]  col_out_732;
wire  [1:0]  col_out_733;
wire  [1:0]  col_out_734;
wire  [1:0]  col_out_735;
wire  [1:0]  col_out_736;
wire  [1:0]  col_out_737;
wire  [1:0]  col_out_738;
wire  [1:0]  col_out_739;
wire  [1:0]  col_out_740;
wire  [1:0]  col_out_741;
wire  [1:0]  col_out_742;
wire  [1:0]  col_out_743;
wire  [1:0]  col_out_744;
wire  [1:0]  col_out_745;
wire  [1:0]  col_out_746;
wire  [1:0]  col_out_747;
wire  [1:0]  col_out_748;
wire  [1:0]  col_out_749;
wire  [1:0]  col_out_750;
wire  [1:0]  col_out_751;
wire  [1:0]  col_out_752;
wire  [1:0]  col_out_753;
wire  [1:0]  col_out_754;
wire  [1:0]  col_out_755;
wire  [1:0]  col_out_756;
wire  [1:0]  col_out_757;
wire  [1:0]  col_out_758;
wire  [1:0]  col_out_759;
wire  [1:0]  col_out_760;
wire  [1:0]  col_out_761;
wire  [1:0]  col_out_762;
wire  [1:0]  col_out_763;
wire  [1:0]  col_out_764;
wire  [1:0]  col_out_765;
wire  [1:0]  col_out_766;
wire  [1:0]  col_out_767;
wire  [1:0]  col_out_768;
wire  [1:0]  col_out_769;
wire  [1:0]  col_out_770;
wire  [1:0]  col_out_771;
wire  [1:0]  col_out_772;
wire  [1:0]  col_out_773;
wire  [1:0]  col_out_774;
wire  [1:0]  col_out_775;
wire  [1:0]  col_out_776;
wire  [1:0]  col_out_777;
wire  [1:0]  col_out_778;
wire  [1:0]  col_out_779;
wire  [1:0]  col_out_780;
wire  [1:0]  col_out_781;
wire  [1:0]  col_out_782;
wire  [1:0]  col_out_783;
wire  [1:0]  col_out_784;
wire  [1:0]  col_out_785;
wire  [1:0]  col_out_786;
wire  [1:0]  col_out_787;
wire  [1:0]  col_out_788;
wire  [1:0]  col_out_789;
wire  [1:0]  col_out_790;
wire  [1:0]  col_out_791;
wire  [1:0]  col_out_792;
wire  [1:0]  col_out_793;
wire  [1:0]  col_out_794;
wire  [1:0]  col_out_795;
wire  [1:0]  col_out_796;
wire  [1:0]  col_out_797;
wire  [1:0]  col_out_798;
wire  [1:0]  col_out_799;
wire  [1:0]  col_out_800;
wire  [1:0]  col_out_801;
wire  [1:0]  col_out_802;
wire  [1:0]  col_out_803;
wire  [1:0]  col_out_804;
wire  [1:0]  col_out_805;
wire  [1:0]  col_out_806;
wire  [1:0]  col_out_807;
wire  [1:0]  col_out_808;
wire  [1:0]  col_out_809;
wire  [1:0]  col_out_810;
wire  [1:0]  col_out_811;
wire  [1:0]  col_out_812;
wire  [1:0]  col_out_813;
wire  [1:0]  col_out_814;
wire  [1:0]  col_out_815;
wire  [1:0]  col_out_816;
wire  [1:0]  col_out_817;
wire  [1:0]  col_out_818;
wire  [1:0]  col_out_819;
wire  [1:0]  col_out_820;
wire  [1:0]  col_out_821;
wire  [1:0]  col_out_822;
wire  [1:0]  col_out_823;
wire  [1:0]  col_out_824;
wire  [1:0]  col_out_825;
wire  [1:0]  col_out_826;
wire  [1:0]  col_out_827;
wire  [1:0]  col_out_828;
wire  [1:0]  col_out_829;
wire  [1:0]  col_out_830;
wire  [1:0]  col_out_831;
wire  [1:0]  col_out_832;
wire  [1:0]  col_out_833;
wire  [1:0]  col_out_834;
wire  [1:0]  col_out_835;
wire  [1:0]  col_out_836;
wire  [1:0]  col_out_837;
wire  [1:0]  col_out_838;
wire  [1:0]  col_out_839;
wire  [1:0]  col_out_840;
wire  [1:0]  col_out_841;
wire  [1:0]  col_out_842;
wire  [1:0]  col_out_843;
wire  [1:0]  col_out_844;
wire  [1:0]  col_out_845;
wire  [1:0]  col_out_846;
wire  [1:0]  col_out_847;
wire  [1:0]  col_out_848;
wire  [1:0]  col_out_849;
wire  [1:0]  col_out_850;
wire  [1:0]  col_out_851;
wire  [1:0]  col_out_852;
wire  [1:0]  col_out_853;
wire  [1:0]  col_out_854;
wire  [1:0]  col_out_855;
wire  [1:0]  col_out_856;
wire  [1:0]  col_out_857;
wire  [1:0]  col_out_858;
wire  [1:0]  col_out_859;
wire  [1:0]  col_out_860;
wire  [1:0]  col_out_861;
wire  [1:0]  col_out_862;
wire  [1:0]  col_out_863;
wire  [1:0]  col_out_864;
wire  [1:0]  col_out_865;
wire  [1:0]  col_out_866;
wire  [1:0]  col_out_867;
wire  [1:0]  col_out_868;
wire  [1:0]  col_out_869;
wire  [1:0]  col_out_870;
wire  [1:0]  col_out_871;
wire  [1:0]  col_out_872;
wire  [1:0]  col_out_873;
wire  [1:0]  col_out_874;
wire  [1:0]  col_out_875;
wire  [1:0]  col_out_876;
wire  [1:0]  col_out_877;
wire  [1:0]  col_out_878;
wire  [1:0]  col_out_879;
wire  [1:0]  col_out_880;
wire  [1:0]  col_out_881;
wire  [1:0]  col_out_882;
wire  [1:0]  col_out_883;
wire  [1:0]  col_out_884;
wire  [1:0]  col_out_885;
wire  [1:0]  col_out_886;
wire  [1:0]  col_out_887;
wire  [1:0]  col_out_888;
wire  [1:0]  col_out_889;
wire  [1:0]  col_out_890;
wire  [1:0]  col_out_891;
wire  [1:0]  col_out_892;
wire  [1:0]  col_out_893;
wire  [1:0]  col_out_894;
wire  [1:0]  col_out_895;
wire  [1:0]  col_out_896;
wire  [1:0]  col_out_897;
wire  [1:0]  col_out_898;
wire  [1:0]  col_out_899;
wire  [1:0]  col_out_900;
wire  [1:0]  col_out_901;
wire  [1:0]  col_out_902;
wire  [1:0]  col_out_903;
wire  [1:0]  col_out_904;
wire  [1:0]  col_out_905;
wire  [1:0]  col_out_906;
wire  [1:0]  col_out_907;
wire  [1:0]  col_out_908;
wire  [1:0]  col_out_909;
wire  [1:0]  col_out_910;
wire  [1:0]  col_out_911;
wire  [1:0]  col_out_912;
wire  [1:0]  col_out_913;
wire  [1:0]  col_out_914;
wire  [1:0]  col_out_915;
wire  [1:0]  col_out_916;
wire  [1:0]  col_out_917;
wire  [1:0]  col_out_918;
wire  [1:0]  col_out_919;
wire  [1:0]  col_out_920;
wire  [1:0]  col_out_921;
wire  [1:0]  col_out_922;
wire  [1:0]  col_out_923;
wire  [1:0]  col_out_924;
wire  [1:0]  col_out_925;
wire  [1:0]  col_out_926;
wire  [1:0]  col_out_927;
wire  [1:0]  col_out_928;
wire  [1:0]  col_out_929;
wire  [1:0]  col_out_930;
wire  [1:0]  col_out_931;
wire  [1:0]  col_out_932;
wire  [1:0]  col_out_933;
wire  [1:0]  col_out_934;
wire  [1:0]  col_out_935;
wire  [1:0]  col_out_936;
wire  [1:0]  col_out_937;
wire  [1:0]  col_out_938;
wire  [1:0]  col_out_939;
wire  [1:0]  col_out_940;
wire  [1:0]  col_out_941;
wire  [1:0]  col_out_942;
wire  [1:0]  col_out_943;
wire  [1:0]  col_out_944;
wire  [1:0]  col_out_945;
wire  [1:0]  col_out_946;
wire  [1:0]  col_out_947;
wire  [1:0]  col_out_948;
wire  [1:0]  col_out_949;
wire  [1:0]  col_out_950;
wire  [1:0]  col_out_951;
wire  [1:0]  col_out_952;
wire  [1:0]  col_out_953;
wire  [1:0]  col_out_954;
wire  [1:0]  col_out_955;
wire  [1:0]  col_out_956;
wire  [1:0]  col_out_957;
wire  [1:0]  col_out_958;
wire  [1:0]  col_out_959;
wire  [1:0]  col_out_960;
wire  [1:0]  col_out_961;
wire  [1:0]  col_out_962;
wire  [1:0]  col_out_963;
wire  [1:0]  col_out_964;
wire  [1:0]  col_out_965;
wire  [1:0]  col_out_966;
wire  [1:0]  col_out_967;
wire  [1:0]  col_out_968;
wire  [1:0]  col_out_969;
wire  [1:0]  col_out_970;
wire  [1:0]  col_out_971;
wire  [1:0]  col_out_972;
wire  [1:0]  col_out_973;
wire  [1:0]  col_out_974;
wire  [1:0]  col_out_975;
wire  [1:0]  col_out_976;
wire  [1:0]  col_out_977;
wire  [1:0]  col_out_978;
wire  [1:0]  col_out_979;
wire  [1:0]  col_out_980;
wire  [1:0]  col_out_981;
wire  [1:0]  col_out_982;
wire  [1:0]  col_out_983;
wire  [1:0]  col_out_984;
wire  [1:0]  col_out_985;
wire  [1:0]  col_out_986;
wire  [1:0]  col_out_987;
wire  [1:0]  col_out_988;
wire  [1:0]  col_out_989;
wire  [1:0]  col_out_990;
wire  [1:0]  col_out_991;
wire  [1:0]  col_out_992;
wire  [1:0]  col_out_993;
wire  [1:0]  col_out_994;
wire  [1:0]  col_out_995;
wire  [1:0]  col_out_996;
wire  [1:0]  col_out_997;
wire  [1:0]  col_out_998;
wire  [1:0]  col_out_999;
wire  [1:0]  col_out_1000;
wire  [1:0]  col_out_1001;
wire  [1:0]  col_out_1002;
wire  [1:0]  col_out_1003;
wire  [1:0]  col_out_1004;
wire  [1:0]  col_out_1005;
wire  [1:0]  col_out_1006;
wire  [1:0]  col_out_1007;
wire  [1:0]  col_out_1008;
wire  [1:0]  col_out_1009;
wire  [1:0]  col_out_1010;
wire  [1:0]  col_out_1011;
wire  [1:0]  col_out_1012;
wire  [1:0]  col_out_1013;
wire  [1:0]  col_out_1014;
wire  [1:0]  col_out_1015;
wire  [1:0]  col_out_1016;
wire  [1:0]  col_out_1017;
wire  [1:0]  col_out_1018;
wire  [1:0]  col_out_1019;
wire  [1:0]  col_out_1020;
wire  [1:0]  col_out_1021;
wire  [1:0]  col_out_1022;
wire  [1:0]  col_out_1023;
wire  [1:0]  col_out_1024;
wire  [1:0]  col_out_1025;
wire  [1:0]  col_out_1026;
wire  [1:0]  col_out_1027;
wire  [1:0]  col_out_1028;
wire  [1:0]  col_out_1029;
wire  [1:0]  col_out_1030;
wire  [1:0]  col_out_1031;
wire  [1:0]  col_out_1032;

compressor_array_512_2_1024  u_compressor_array_512_2_1024 (
    .col_in_0                ( col_in_0       ),
    .col_in_1                ( col_in_1       ),
    .col_in_2                ( col_in_2       ),
    .col_in_3                ( col_in_3       ),
    .col_in_4                ( col_in_4       ),
    .col_in_5                ( col_in_5       ),
    .col_in_6                ( col_in_6       ),
    .col_in_7                ( col_in_7       ),
    .col_in_8                ( col_in_8       ),
    .col_in_9                ( col_in_9       ),
    .col_in_10               ( col_in_10      ),
    .col_in_11               ( col_in_11      ),
    .col_in_12               ( col_in_12      ),
    .col_in_13               ( col_in_13      ),
    .col_in_14               ( col_in_14      ),
    .col_in_15               ( col_in_15      ),
    .col_in_16               ( col_in_16      ),
    .col_in_17               ( col_in_17      ),
    .col_in_18               ( col_in_18      ),
    .col_in_19               ( col_in_19      ),
    .col_in_20               ( col_in_20      ),
    .col_in_21               ( col_in_21      ),
    .col_in_22               ( col_in_22      ),
    .col_in_23               ( col_in_23      ),
    .col_in_24               ( col_in_24      ),
    .col_in_25               ( col_in_25      ),
    .col_in_26               ( col_in_26      ),
    .col_in_27               ( col_in_27      ),
    .col_in_28               ( col_in_28      ),
    .col_in_29               ( col_in_29      ),
    .col_in_30               ( col_in_30      ),
    .col_in_31               ( col_in_31      ),
    .col_in_32               ( col_in_32      ),
    .col_in_33               ( col_in_33      ),
    .col_in_34               ( col_in_34      ),
    .col_in_35               ( col_in_35      ),
    .col_in_36               ( col_in_36      ),
    .col_in_37               ( col_in_37      ),
    .col_in_38               ( col_in_38      ),
    .col_in_39               ( col_in_39      ),
    .col_in_40               ( col_in_40      ),
    .col_in_41               ( col_in_41      ),
    .col_in_42               ( col_in_42      ),
    .col_in_43               ( col_in_43      ),
    .col_in_44               ( col_in_44      ),
    .col_in_45               ( col_in_45      ),
    .col_in_46               ( col_in_46      ),
    .col_in_47               ( col_in_47      ),
    .col_in_48               ( col_in_48      ),
    .col_in_49               ( col_in_49      ),
    .col_in_50               ( col_in_50      ),
    .col_in_51               ( col_in_51      ),
    .col_in_52               ( col_in_52      ),
    .col_in_53               ( col_in_53      ),
    .col_in_54               ( col_in_54      ),
    .col_in_55               ( col_in_55      ),
    .col_in_56               ( col_in_56      ),
    .col_in_57               ( col_in_57      ),
    .col_in_58               ( col_in_58      ),
    .col_in_59               ( col_in_59      ),
    .col_in_60               ( col_in_60      ),
    .col_in_61               ( col_in_61      ),
    .col_in_62               ( col_in_62      ),
    .col_in_63               ( col_in_63      ),
    .col_in_64               ( col_in_64      ),
    .col_in_65               ( col_in_65      ),
    .col_in_66               ( col_in_66      ),
    .col_in_67               ( col_in_67      ),
    .col_in_68               ( col_in_68      ),
    .col_in_69               ( col_in_69      ),
    .col_in_70               ( col_in_70      ),
    .col_in_71               ( col_in_71      ),
    .col_in_72               ( col_in_72      ),
    .col_in_73               ( col_in_73      ),
    .col_in_74               ( col_in_74      ),
    .col_in_75               ( col_in_75      ),
    .col_in_76               ( col_in_76      ),
    .col_in_77               ( col_in_77      ),
    .col_in_78               ( col_in_78      ),
    .col_in_79               ( col_in_79      ),
    .col_in_80               ( col_in_80      ),
    .col_in_81               ( col_in_81      ),
    .col_in_82               ( col_in_82      ),
    .col_in_83               ( col_in_83      ),
    .col_in_84               ( col_in_84      ),
    .col_in_85               ( col_in_85      ),
    .col_in_86               ( col_in_86      ),
    .col_in_87               ( col_in_87      ),
    .col_in_88               ( col_in_88      ),
    .col_in_89               ( col_in_89      ),
    .col_in_90               ( col_in_90      ),
    .col_in_91               ( col_in_91      ),
    .col_in_92               ( col_in_92      ),
    .col_in_93               ( col_in_93      ),
    .col_in_94               ( col_in_94      ),
    .col_in_95               ( col_in_95      ),
    .col_in_96               ( col_in_96      ),
    .col_in_97               ( col_in_97      ),
    .col_in_98               ( col_in_98      ),
    .col_in_99               ( col_in_99      ),
    .col_in_100              ( col_in_100     ),
    .col_in_101              ( col_in_101     ),
    .col_in_102              ( col_in_102     ),
    .col_in_103              ( col_in_103     ),
    .col_in_104              ( col_in_104     ),
    .col_in_105              ( col_in_105     ),
    .col_in_106              ( col_in_106     ),
    .col_in_107              ( col_in_107     ),
    .col_in_108              ( col_in_108     ),
    .col_in_109              ( col_in_109     ),
    .col_in_110              ( col_in_110     ),
    .col_in_111              ( col_in_111     ),
    .col_in_112              ( col_in_112     ),
    .col_in_113              ( col_in_113     ),
    .col_in_114              ( col_in_114     ),
    .col_in_115              ( col_in_115     ),
    .col_in_116              ( col_in_116     ),
    .col_in_117              ( col_in_117     ),
    .col_in_118              ( col_in_118     ),
    .col_in_119              ( col_in_119     ),
    .col_in_120              ( col_in_120     ),
    .col_in_121              ( col_in_121     ),
    .col_in_122              ( col_in_122     ),
    .col_in_123              ( col_in_123     ),
    .col_in_124              ( col_in_124     ),
    .col_in_125              ( col_in_125     ),
    .col_in_126              ( col_in_126     ),
    .col_in_127              ( col_in_127     ),
    .col_in_128              ( col_in_128     ),
    .col_in_129              ( col_in_129     ),
    .col_in_130              ( col_in_130     ),
    .col_in_131              ( col_in_131     ),
    .col_in_132              ( col_in_132     ),
    .col_in_133              ( col_in_133     ),
    .col_in_134              ( col_in_134     ),
    .col_in_135              ( col_in_135     ),
    .col_in_136              ( col_in_136     ),
    .col_in_137              ( col_in_137     ),
    .col_in_138              ( col_in_138     ),
    .col_in_139              ( col_in_139     ),
    .col_in_140              ( col_in_140     ),
    .col_in_141              ( col_in_141     ),
    .col_in_142              ( col_in_142     ),
    .col_in_143              ( col_in_143     ),
    .col_in_144              ( col_in_144     ),
    .col_in_145              ( col_in_145     ),
    .col_in_146              ( col_in_146     ),
    .col_in_147              ( col_in_147     ),
    .col_in_148              ( col_in_148     ),
    .col_in_149              ( col_in_149     ),
    .col_in_150              ( col_in_150     ),
    .col_in_151              ( col_in_151     ),
    .col_in_152              ( col_in_152     ),
    .col_in_153              ( col_in_153     ),
    .col_in_154              ( col_in_154     ),
    .col_in_155              ( col_in_155     ),
    .col_in_156              ( col_in_156     ),
    .col_in_157              ( col_in_157     ),
    .col_in_158              ( col_in_158     ),
    .col_in_159              ( col_in_159     ),
    .col_in_160              ( col_in_160     ),
    .col_in_161              ( col_in_161     ),
    .col_in_162              ( col_in_162     ),
    .col_in_163              ( col_in_163     ),
    .col_in_164              ( col_in_164     ),
    .col_in_165              ( col_in_165     ),
    .col_in_166              ( col_in_166     ),
    .col_in_167              ( col_in_167     ),
    .col_in_168              ( col_in_168     ),
    .col_in_169              ( col_in_169     ),
    .col_in_170              ( col_in_170     ),
    .col_in_171              ( col_in_171     ),
    .col_in_172              ( col_in_172     ),
    .col_in_173              ( col_in_173     ),
    .col_in_174              ( col_in_174     ),
    .col_in_175              ( col_in_175     ),
    .col_in_176              ( col_in_176     ),
    .col_in_177              ( col_in_177     ),
    .col_in_178              ( col_in_178     ),
    .col_in_179              ( col_in_179     ),
    .col_in_180              ( col_in_180     ),
    .col_in_181              ( col_in_181     ),
    .col_in_182              ( col_in_182     ),
    .col_in_183              ( col_in_183     ),
    .col_in_184              ( col_in_184     ),
    .col_in_185              ( col_in_185     ),
    .col_in_186              ( col_in_186     ),
    .col_in_187              ( col_in_187     ),
    .col_in_188              ( col_in_188     ),
    .col_in_189              ( col_in_189     ),
    .col_in_190              ( col_in_190     ),
    .col_in_191              ( col_in_191     ),
    .col_in_192              ( col_in_192     ),
    .col_in_193              ( col_in_193     ),
    .col_in_194              ( col_in_194     ),
    .col_in_195              ( col_in_195     ),
    .col_in_196              ( col_in_196     ),
    .col_in_197              ( col_in_197     ),
    .col_in_198              ( col_in_198     ),
    .col_in_199              ( col_in_199     ),
    .col_in_200              ( col_in_200     ),
    .col_in_201              ( col_in_201     ),
    .col_in_202              ( col_in_202     ),
    .col_in_203              ( col_in_203     ),
    .col_in_204              ( col_in_204     ),
    .col_in_205              ( col_in_205     ),
    .col_in_206              ( col_in_206     ),
    .col_in_207              ( col_in_207     ),
    .col_in_208              ( col_in_208     ),
    .col_in_209              ( col_in_209     ),
    .col_in_210              ( col_in_210     ),
    .col_in_211              ( col_in_211     ),
    .col_in_212              ( col_in_212     ),
    .col_in_213              ( col_in_213     ),
    .col_in_214              ( col_in_214     ),
    .col_in_215              ( col_in_215     ),
    .col_in_216              ( col_in_216     ),
    .col_in_217              ( col_in_217     ),
    .col_in_218              ( col_in_218     ),
    .col_in_219              ( col_in_219     ),
    .col_in_220              ( col_in_220     ),
    .col_in_221              ( col_in_221     ),
    .col_in_222              ( col_in_222     ),
    .col_in_223              ( col_in_223     ),
    .col_in_224              ( col_in_224     ),
    .col_in_225              ( col_in_225     ),
    .col_in_226              ( col_in_226     ),
    .col_in_227              ( col_in_227     ),
    .col_in_228              ( col_in_228     ),
    .col_in_229              ( col_in_229     ),
    .col_in_230              ( col_in_230     ),
    .col_in_231              ( col_in_231     ),
    .col_in_232              ( col_in_232     ),
    .col_in_233              ( col_in_233     ),
    .col_in_234              ( col_in_234     ),
    .col_in_235              ( col_in_235     ),
    .col_in_236              ( col_in_236     ),
    .col_in_237              ( col_in_237     ),
    .col_in_238              ( col_in_238     ),
    .col_in_239              ( col_in_239     ),
    .col_in_240              ( col_in_240     ),
    .col_in_241              ( col_in_241     ),
    .col_in_242              ( col_in_242     ),
    .col_in_243              ( col_in_243     ),
    .col_in_244              ( col_in_244     ),
    .col_in_245              ( col_in_245     ),
    .col_in_246              ( col_in_246     ),
    .col_in_247              ( col_in_247     ),
    .col_in_248              ( col_in_248     ),
    .col_in_249              ( col_in_249     ),
    .col_in_250              ( col_in_250     ),
    .col_in_251              ( col_in_251     ),
    .col_in_252              ( col_in_252     ),
    .col_in_253              ( col_in_253     ),
    .col_in_254              ( col_in_254     ),
    .col_in_255              ( col_in_255     ),
    .col_in_256              ( col_in_256     ),
    .col_in_257              ( col_in_257     ),
    .col_in_258              ( col_in_258     ),
    .col_in_259              ( col_in_259     ),
    .col_in_260              ( col_in_260     ),
    .col_in_261              ( col_in_261     ),
    .col_in_262              ( col_in_262     ),
    .col_in_263              ( col_in_263     ),
    .col_in_264              ( col_in_264     ),
    .col_in_265              ( col_in_265     ),
    .col_in_266              ( col_in_266     ),
    .col_in_267              ( col_in_267     ),
    .col_in_268              ( col_in_268     ),
    .col_in_269              ( col_in_269     ),
    .col_in_270              ( col_in_270     ),
    .col_in_271              ( col_in_271     ),
    .col_in_272              ( col_in_272     ),
    .col_in_273              ( col_in_273     ),
    .col_in_274              ( col_in_274     ),
    .col_in_275              ( col_in_275     ),
    .col_in_276              ( col_in_276     ),
    .col_in_277              ( col_in_277     ),
    .col_in_278              ( col_in_278     ),
    .col_in_279              ( col_in_279     ),
    .col_in_280              ( col_in_280     ),
    .col_in_281              ( col_in_281     ),
    .col_in_282              ( col_in_282     ),
    .col_in_283              ( col_in_283     ),
    .col_in_284              ( col_in_284     ),
    .col_in_285              ( col_in_285     ),
    .col_in_286              ( col_in_286     ),
    .col_in_287              ( col_in_287     ),
    .col_in_288              ( col_in_288     ),
    .col_in_289              ( col_in_289     ),
    .col_in_290              ( col_in_290     ),
    .col_in_291              ( col_in_291     ),
    .col_in_292              ( col_in_292     ),
    .col_in_293              ( col_in_293     ),
    .col_in_294              ( col_in_294     ),
    .col_in_295              ( col_in_295     ),
    .col_in_296              ( col_in_296     ),
    .col_in_297              ( col_in_297     ),
    .col_in_298              ( col_in_298     ),
    .col_in_299              ( col_in_299     ),
    .col_in_300              ( col_in_300     ),
    .col_in_301              ( col_in_301     ),
    .col_in_302              ( col_in_302     ),
    .col_in_303              ( col_in_303     ),
    .col_in_304              ( col_in_304     ),
    .col_in_305              ( col_in_305     ),
    .col_in_306              ( col_in_306     ),
    .col_in_307              ( col_in_307     ),
    .col_in_308              ( col_in_308     ),
    .col_in_309              ( col_in_309     ),
    .col_in_310              ( col_in_310     ),
    .col_in_311              ( col_in_311     ),
    .col_in_312              ( col_in_312     ),
    .col_in_313              ( col_in_313     ),
    .col_in_314              ( col_in_314     ),
    .col_in_315              ( col_in_315     ),
    .col_in_316              ( col_in_316     ),
    .col_in_317              ( col_in_317     ),
    .col_in_318              ( col_in_318     ),
    .col_in_319              ( col_in_319     ),
    .col_in_320              ( col_in_320     ),
    .col_in_321              ( col_in_321     ),
    .col_in_322              ( col_in_322     ),
    .col_in_323              ( col_in_323     ),
    .col_in_324              ( col_in_324     ),
    .col_in_325              ( col_in_325     ),
    .col_in_326              ( col_in_326     ),
    .col_in_327              ( col_in_327     ),
    .col_in_328              ( col_in_328     ),
    .col_in_329              ( col_in_329     ),
    .col_in_330              ( col_in_330     ),
    .col_in_331              ( col_in_331     ),
    .col_in_332              ( col_in_332     ),
    .col_in_333              ( col_in_333     ),
    .col_in_334              ( col_in_334     ),
    .col_in_335              ( col_in_335     ),
    .col_in_336              ( col_in_336     ),
    .col_in_337              ( col_in_337     ),
    .col_in_338              ( col_in_338     ),
    .col_in_339              ( col_in_339     ),
    .col_in_340              ( col_in_340     ),
    .col_in_341              ( col_in_341     ),
    .col_in_342              ( col_in_342     ),
    .col_in_343              ( col_in_343     ),
    .col_in_344              ( col_in_344     ),
    .col_in_345              ( col_in_345     ),
    .col_in_346              ( col_in_346     ),
    .col_in_347              ( col_in_347     ),
    .col_in_348              ( col_in_348     ),
    .col_in_349              ( col_in_349     ),
    .col_in_350              ( col_in_350     ),
    .col_in_351              ( col_in_351     ),
    .col_in_352              ( col_in_352     ),
    .col_in_353              ( col_in_353     ),
    .col_in_354              ( col_in_354     ),
    .col_in_355              ( col_in_355     ),
    .col_in_356              ( col_in_356     ),
    .col_in_357              ( col_in_357     ),
    .col_in_358              ( col_in_358     ),
    .col_in_359              ( col_in_359     ),
    .col_in_360              ( col_in_360     ),
    .col_in_361              ( col_in_361     ),
    .col_in_362              ( col_in_362     ),
    .col_in_363              ( col_in_363     ),
    .col_in_364              ( col_in_364     ),
    .col_in_365              ( col_in_365     ),
    .col_in_366              ( col_in_366     ),
    .col_in_367              ( col_in_367     ),
    .col_in_368              ( col_in_368     ),
    .col_in_369              ( col_in_369     ),
    .col_in_370              ( col_in_370     ),
    .col_in_371              ( col_in_371     ),
    .col_in_372              ( col_in_372     ),
    .col_in_373              ( col_in_373     ),
    .col_in_374              ( col_in_374     ),
    .col_in_375              ( col_in_375     ),
    .col_in_376              ( col_in_376     ),
    .col_in_377              ( col_in_377     ),
    .col_in_378              ( col_in_378     ),
    .col_in_379              ( col_in_379     ),
    .col_in_380              ( col_in_380     ),
    .col_in_381              ( col_in_381     ),
    .col_in_382              ( col_in_382     ),
    .col_in_383              ( col_in_383     ),
    .col_in_384              ( col_in_384     ),
    .col_in_385              ( col_in_385     ),
    .col_in_386              ( col_in_386     ),
    .col_in_387              ( col_in_387     ),
    .col_in_388              ( col_in_388     ),
    .col_in_389              ( col_in_389     ),
    .col_in_390              ( col_in_390     ),
    .col_in_391              ( col_in_391     ),
    .col_in_392              ( col_in_392     ),
    .col_in_393              ( col_in_393     ),
    .col_in_394              ( col_in_394     ),
    .col_in_395              ( col_in_395     ),
    .col_in_396              ( col_in_396     ),
    .col_in_397              ( col_in_397     ),
    .col_in_398              ( col_in_398     ),
    .col_in_399              ( col_in_399     ),
    .col_in_400              ( col_in_400     ),
    .col_in_401              ( col_in_401     ),
    .col_in_402              ( col_in_402     ),
    .col_in_403              ( col_in_403     ),
    .col_in_404              ( col_in_404     ),
    .col_in_405              ( col_in_405     ),
    .col_in_406              ( col_in_406     ),
    .col_in_407              ( col_in_407     ),
    .col_in_408              ( col_in_408     ),
    .col_in_409              ( col_in_409     ),
    .col_in_410              ( col_in_410     ),
    .col_in_411              ( col_in_411     ),
    .col_in_412              ( col_in_412     ),
    .col_in_413              ( col_in_413     ),
    .col_in_414              ( col_in_414     ),
    .col_in_415              ( col_in_415     ),
    .col_in_416              ( col_in_416     ),
    .col_in_417              ( col_in_417     ),
    .col_in_418              ( col_in_418     ),
    .col_in_419              ( col_in_419     ),
    .col_in_420              ( col_in_420     ),
    .col_in_421              ( col_in_421     ),
    .col_in_422              ( col_in_422     ),
    .col_in_423              ( col_in_423     ),
    .col_in_424              ( col_in_424     ),
    .col_in_425              ( col_in_425     ),
    .col_in_426              ( col_in_426     ),
    .col_in_427              ( col_in_427     ),
    .col_in_428              ( col_in_428     ),
    .col_in_429              ( col_in_429     ),
    .col_in_430              ( col_in_430     ),
    .col_in_431              ( col_in_431     ),
    .col_in_432              ( col_in_432     ),
    .col_in_433              ( col_in_433     ),
    .col_in_434              ( col_in_434     ),
    .col_in_435              ( col_in_435     ),
    .col_in_436              ( col_in_436     ),
    .col_in_437              ( col_in_437     ),
    .col_in_438              ( col_in_438     ),
    .col_in_439              ( col_in_439     ),
    .col_in_440              ( col_in_440     ),
    .col_in_441              ( col_in_441     ),
    .col_in_442              ( col_in_442     ),
    .col_in_443              ( col_in_443     ),
    .col_in_444              ( col_in_444     ),
    .col_in_445              ( col_in_445     ),
    .col_in_446              ( col_in_446     ),
    .col_in_447              ( col_in_447     ),
    .col_in_448              ( col_in_448     ),
    .col_in_449              ( col_in_449     ),
    .col_in_450              ( col_in_450     ),
    .col_in_451              ( col_in_451     ),
    .col_in_452              ( col_in_452     ),
    .col_in_453              ( col_in_453     ),
    .col_in_454              ( col_in_454     ),
    .col_in_455              ( col_in_455     ),
    .col_in_456              ( col_in_456     ),
    .col_in_457              ( col_in_457     ),
    .col_in_458              ( col_in_458     ),
    .col_in_459              ( col_in_459     ),
    .col_in_460              ( col_in_460     ),
    .col_in_461              ( col_in_461     ),
    .col_in_462              ( col_in_462     ),
    .col_in_463              ( col_in_463     ),
    .col_in_464              ( col_in_464     ),
    .col_in_465              ( col_in_465     ),
    .col_in_466              ( col_in_466     ),
    .col_in_467              ( col_in_467     ),
    .col_in_468              ( col_in_468     ),
    .col_in_469              ( col_in_469     ),
    .col_in_470              ( col_in_470     ),
    .col_in_471              ( col_in_471     ),
    .col_in_472              ( col_in_472     ),
    .col_in_473              ( col_in_473     ),
    .col_in_474              ( col_in_474     ),
    .col_in_475              ( col_in_475     ),
    .col_in_476              ( col_in_476     ),
    .col_in_477              ( col_in_477     ),
    .col_in_478              ( col_in_478     ),
    .col_in_479              ( col_in_479     ),
    .col_in_480              ( col_in_480     ),
    .col_in_481              ( col_in_481     ),
    .col_in_482              ( col_in_482     ),
    .col_in_483              ( col_in_483     ),
    .col_in_484              ( col_in_484     ),
    .col_in_485              ( col_in_485     ),
    .col_in_486              ( col_in_486     ),
    .col_in_487              ( col_in_487     ),
    .col_in_488              ( col_in_488     ),
    .col_in_489              ( col_in_489     ),
    .col_in_490              ( col_in_490     ),
    .col_in_491              ( col_in_491     ),
    .col_in_492              ( col_in_492     ),
    .col_in_493              ( col_in_493     ),
    .col_in_494              ( col_in_494     ),
    .col_in_495              ( col_in_495     ),
    .col_in_496              ( col_in_496     ),
    .col_in_497              ( col_in_497     ),
    .col_in_498              ( col_in_498     ),
    .col_in_499              ( col_in_499     ),
    .col_in_500              ( col_in_500     ),
    .col_in_501              ( col_in_501     ),
    .col_in_502              ( col_in_502     ),
    .col_in_503              ( col_in_503     ),
    .col_in_504              ( col_in_504     ),
    .col_in_505              ( col_in_505     ),
    .col_in_506              ( col_in_506     ),
    .col_in_507              ( col_in_507     ),
    .col_in_508              ( col_in_508     ),
    .col_in_509              ( col_in_509     ),
    .col_in_510              ( col_in_510     ),
    .col_in_511              ( col_in_511     ),
    .col_in_512              ( col_in_512     ),
    .col_in_513              ( col_in_513     ),
    .col_in_514              ( col_in_514     ),
    .col_in_515              ( col_in_515     ),
    .col_in_516              ( col_in_516     ),
    .col_in_517              ( col_in_517     ),
    .col_in_518              ( col_in_518     ),
    .col_in_519              ( col_in_519     ),
    .col_in_520              ( col_in_520     ),
    .col_in_521              ( col_in_521     ),
    .col_in_522              ( col_in_522     ),
    .col_in_523              ( col_in_523     ),
    .col_in_524              ( col_in_524     ),
    .col_in_525              ( col_in_525     ),
    .col_in_526              ( col_in_526     ),
    .col_in_527              ( col_in_527     ),
    .col_in_528              ( col_in_528     ),
    .col_in_529              ( col_in_529     ),
    .col_in_530              ( col_in_530     ),
    .col_in_531              ( col_in_531     ),
    .col_in_532              ( col_in_532     ),
    .col_in_533              ( col_in_533     ),
    .col_in_534              ( col_in_534     ),
    .col_in_535              ( col_in_535     ),
    .col_in_536              ( col_in_536     ),
    .col_in_537              ( col_in_537     ),
    .col_in_538              ( col_in_538     ),
    .col_in_539              ( col_in_539     ),
    .col_in_540              ( col_in_540     ),
    .col_in_541              ( col_in_541     ),
    .col_in_542              ( col_in_542     ),
    .col_in_543              ( col_in_543     ),
    .col_in_544              ( col_in_544     ),
    .col_in_545              ( col_in_545     ),
    .col_in_546              ( col_in_546     ),
    .col_in_547              ( col_in_547     ),
    .col_in_548              ( col_in_548     ),
    .col_in_549              ( col_in_549     ),
    .col_in_550              ( col_in_550     ),
    .col_in_551              ( col_in_551     ),
    .col_in_552              ( col_in_552     ),
    .col_in_553              ( col_in_553     ),
    .col_in_554              ( col_in_554     ),
    .col_in_555              ( col_in_555     ),
    .col_in_556              ( col_in_556     ),
    .col_in_557              ( col_in_557     ),
    .col_in_558              ( col_in_558     ),
    .col_in_559              ( col_in_559     ),
    .col_in_560              ( col_in_560     ),
    .col_in_561              ( col_in_561     ),
    .col_in_562              ( col_in_562     ),
    .col_in_563              ( col_in_563     ),
    .col_in_564              ( col_in_564     ),
    .col_in_565              ( col_in_565     ),
    .col_in_566              ( col_in_566     ),
    .col_in_567              ( col_in_567     ),
    .col_in_568              ( col_in_568     ),
    .col_in_569              ( col_in_569     ),
    .col_in_570              ( col_in_570     ),
    .col_in_571              ( col_in_571     ),
    .col_in_572              ( col_in_572     ),
    .col_in_573              ( col_in_573     ),
    .col_in_574              ( col_in_574     ),
    .col_in_575              ( col_in_575     ),
    .col_in_576              ( col_in_576     ),
    .col_in_577              ( col_in_577     ),
    .col_in_578              ( col_in_578     ),
    .col_in_579              ( col_in_579     ),
    .col_in_580              ( col_in_580     ),
    .col_in_581              ( col_in_581     ),
    .col_in_582              ( col_in_582     ),
    .col_in_583              ( col_in_583     ),
    .col_in_584              ( col_in_584     ),
    .col_in_585              ( col_in_585     ),
    .col_in_586              ( col_in_586     ),
    .col_in_587              ( col_in_587     ),
    .col_in_588              ( col_in_588     ),
    .col_in_589              ( col_in_589     ),
    .col_in_590              ( col_in_590     ),
    .col_in_591              ( col_in_591     ),
    .col_in_592              ( col_in_592     ),
    .col_in_593              ( col_in_593     ),
    .col_in_594              ( col_in_594     ),
    .col_in_595              ( col_in_595     ),
    .col_in_596              ( col_in_596     ),
    .col_in_597              ( col_in_597     ),
    .col_in_598              ( col_in_598     ),
    .col_in_599              ( col_in_599     ),
    .col_in_600              ( col_in_600     ),
    .col_in_601              ( col_in_601     ),
    .col_in_602              ( col_in_602     ),
    .col_in_603              ( col_in_603     ),
    .col_in_604              ( col_in_604     ),
    .col_in_605              ( col_in_605     ),
    .col_in_606              ( col_in_606     ),
    .col_in_607              ( col_in_607     ),
    .col_in_608              ( col_in_608     ),
    .col_in_609              ( col_in_609     ),
    .col_in_610              ( col_in_610     ),
    .col_in_611              ( col_in_611     ),
    .col_in_612              ( col_in_612     ),
    .col_in_613              ( col_in_613     ),
    .col_in_614              ( col_in_614     ),
    .col_in_615              ( col_in_615     ),
    .col_in_616              ( col_in_616     ),
    .col_in_617              ( col_in_617     ),
    .col_in_618              ( col_in_618     ),
    .col_in_619              ( col_in_619     ),
    .col_in_620              ( col_in_620     ),
    .col_in_621              ( col_in_621     ),
    .col_in_622              ( col_in_622     ),
    .col_in_623              ( col_in_623     ),
    .col_in_624              ( col_in_624     ),
    .col_in_625              ( col_in_625     ),
    .col_in_626              ( col_in_626     ),
    .col_in_627              ( col_in_627     ),
    .col_in_628              ( col_in_628     ),
    .col_in_629              ( col_in_629     ),
    .col_in_630              ( col_in_630     ),
    .col_in_631              ( col_in_631     ),
    .col_in_632              ( col_in_632     ),
    .col_in_633              ( col_in_633     ),
    .col_in_634              ( col_in_634     ),
    .col_in_635              ( col_in_635     ),
    .col_in_636              ( col_in_636     ),
    .col_in_637              ( col_in_637     ),
    .col_in_638              ( col_in_638     ),
    .col_in_639              ( col_in_639     ),
    .col_in_640              ( col_in_640     ),
    .col_in_641              ( col_in_641     ),
    .col_in_642              ( col_in_642     ),
    .col_in_643              ( col_in_643     ),
    .col_in_644              ( col_in_644     ),
    .col_in_645              ( col_in_645     ),
    .col_in_646              ( col_in_646     ),
    .col_in_647              ( col_in_647     ),
    .col_in_648              ( col_in_648     ),
    .col_in_649              ( col_in_649     ),
    .col_in_650              ( col_in_650     ),
    .col_in_651              ( col_in_651     ),
    .col_in_652              ( col_in_652     ),
    .col_in_653              ( col_in_653     ),
    .col_in_654              ( col_in_654     ),
    .col_in_655              ( col_in_655     ),
    .col_in_656              ( col_in_656     ),
    .col_in_657              ( col_in_657     ),
    .col_in_658              ( col_in_658     ),
    .col_in_659              ( col_in_659     ),
    .col_in_660              ( col_in_660     ),
    .col_in_661              ( col_in_661     ),
    .col_in_662              ( col_in_662     ),
    .col_in_663              ( col_in_663     ),
    .col_in_664              ( col_in_664     ),
    .col_in_665              ( col_in_665     ),
    .col_in_666              ( col_in_666     ),
    .col_in_667              ( col_in_667     ),
    .col_in_668              ( col_in_668     ),
    .col_in_669              ( col_in_669     ),
    .col_in_670              ( col_in_670     ),
    .col_in_671              ( col_in_671     ),
    .col_in_672              ( col_in_672     ),
    .col_in_673              ( col_in_673     ),
    .col_in_674              ( col_in_674     ),
    .col_in_675              ( col_in_675     ),
    .col_in_676              ( col_in_676     ),
    .col_in_677              ( col_in_677     ),
    .col_in_678              ( col_in_678     ),
    .col_in_679              ( col_in_679     ),
    .col_in_680              ( col_in_680     ),
    .col_in_681              ( col_in_681     ),
    .col_in_682              ( col_in_682     ),
    .col_in_683              ( col_in_683     ),
    .col_in_684              ( col_in_684     ),
    .col_in_685              ( col_in_685     ),
    .col_in_686              ( col_in_686     ),
    .col_in_687              ( col_in_687     ),
    .col_in_688              ( col_in_688     ),
    .col_in_689              ( col_in_689     ),
    .col_in_690              ( col_in_690     ),
    .col_in_691              ( col_in_691     ),
    .col_in_692              ( col_in_692     ),
    .col_in_693              ( col_in_693     ),
    .col_in_694              ( col_in_694     ),
    .col_in_695              ( col_in_695     ),
    .col_in_696              ( col_in_696     ),
    .col_in_697              ( col_in_697     ),
    .col_in_698              ( col_in_698     ),
    .col_in_699              ( col_in_699     ),
    .col_in_700              ( col_in_700     ),
    .col_in_701              ( col_in_701     ),
    .col_in_702              ( col_in_702     ),
    .col_in_703              ( col_in_703     ),
    .col_in_704              ( col_in_704     ),
    .col_in_705              ( col_in_705     ),
    .col_in_706              ( col_in_706     ),
    .col_in_707              ( col_in_707     ),
    .col_in_708              ( col_in_708     ),
    .col_in_709              ( col_in_709     ),
    .col_in_710              ( col_in_710     ),
    .col_in_711              ( col_in_711     ),
    .col_in_712              ( col_in_712     ),
    .col_in_713              ( col_in_713     ),
    .col_in_714              ( col_in_714     ),
    .col_in_715              ( col_in_715     ),
    .col_in_716              ( col_in_716     ),
    .col_in_717              ( col_in_717     ),
    .col_in_718              ( col_in_718     ),
    .col_in_719              ( col_in_719     ),
    .col_in_720              ( col_in_720     ),
    .col_in_721              ( col_in_721     ),
    .col_in_722              ( col_in_722     ),
    .col_in_723              ( col_in_723     ),
    .col_in_724              ( col_in_724     ),
    .col_in_725              ( col_in_725     ),
    .col_in_726              ( col_in_726     ),
    .col_in_727              ( col_in_727     ),
    .col_in_728              ( col_in_728     ),
    .col_in_729              ( col_in_729     ),
    .col_in_730              ( col_in_730     ),
    .col_in_731              ( col_in_731     ),
    .col_in_732              ( col_in_732     ),
    .col_in_733              ( col_in_733     ),
    .col_in_734              ( col_in_734     ),
    .col_in_735              ( col_in_735     ),
    .col_in_736              ( col_in_736     ),
    .col_in_737              ( col_in_737     ),
    .col_in_738              ( col_in_738     ),
    .col_in_739              ( col_in_739     ),
    .col_in_740              ( col_in_740     ),
    .col_in_741              ( col_in_741     ),
    .col_in_742              ( col_in_742     ),
    .col_in_743              ( col_in_743     ),
    .col_in_744              ( col_in_744     ),
    .col_in_745              ( col_in_745     ),
    .col_in_746              ( col_in_746     ),
    .col_in_747              ( col_in_747     ),
    .col_in_748              ( col_in_748     ),
    .col_in_749              ( col_in_749     ),
    .col_in_750              ( col_in_750     ),
    .col_in_751              ( col_in_751     ),
    .col_in_752              ( col_in_752     ),
    .col_in_753              ( col_in_753     ),
    .col_in_754              ( col_in_754     ),
    .col_in_755              ( col_in_755     ),
    .col_in_756              ( col_in_756     ),
    .col_in_757              ( col_in_757     ),
    .col_in_758              ( col_in_758     ),
    .col_in_759              ( col_in_759     ),
    .col_in_760              ( col_in_760     ),
    .col_in_761              ( col_in_761     ),
    .col_in_762              ( col_in_762     ),
    .col_in_763              ( col_in_763     ),
    .col_in_764              ( col_in_764     ),
    .col_in_765              ( col_in_765     ),
    .col_in_766              ( col_in_766     ),
    .col_in_767              ( col_in_767     ),
    .col_in_768              ( col_in_768     ),
    .col_in_769              ( col_in_769     ),
    .col_in_770              ( col_in_770     ),
    .col_in_771              ( col_in_771     ),
    .col_in_772              ( col_in_772     ),
    .col_in_773              ( col_in_773     ),
    .col_in_774              ( col_in_774     ),
    .col_in_775              ( col_in_775     ),
    .col_in_776              ( col_in_776     ),
    .col_in_777              ( col_in_777     ),
    .col_in_778              ( col_in_778     ),
    .col_in_779              ( col_in_779     ),
    .col_in_780              ( col_in_780     ),
    .col_in_781              ( col_in_781     ),
    .col_in_782              ( col_in_782     ),
    .col_in_783              ( col_in_783     ),
    .col_in_784              ( col_in_784     ),
    .col_in_785              ( col_in_785     ),
    .col_in_786              ( col_in_786     ),
    .col_in_787              ( col_in_787     ),
    .col_in_788              ( col_in_788     ),
    .col_in_789              ( col_in_789     ),
    .col_in_790              ( col_in_790     ),
    .col_in_791              ( col_in_791     ),
    .col_in_792              ( col_in_792     ),
    .col_in_793              ( col_in_793     ),
    .col_in_794              ( col_in_794     ),
    .col_in_795              ( col_in_795     ),
    .col_in_796              ( col_in_796     ),
    .col_in_797              ( col_in_797     ),
    .col_in_798              ( col_in_798     ),
    .col_in_799              ( col_in_799     ),
    .col_in_800              ( col_in_800     ),
    .col_in_801              ( col_in_801     ),
    .col_in_802              ( col_in_802     ),
    .col_in_803              ( col_in_803     ),
    .col_in_804              ( col_in_804     ),
    .col_in_805              ( col_in_805     ),
    .col_in_806              ( col_in_806     ),
    .col_in_807              ( col_in_807     ),
    .col_in_808              ( col_in_808     ),
    .col_in_809              ( col_in_809     ),
    .col_in_810              ( col_in_810     ),
    .col_in_811              ( col_in_811     ),
    .col_in_812              ( col_in_812     ),
    .col_in_813              ( col_in_813     ),
    .col_in_814              ( col_in_814     ),
    .col_in_815              ( col_in_815     ),
    .col_in_816              ( col_in_816     ),
    .col_in_817              ( col_in_817     ),
    .col_in_818              ( col_in_818     ),
    .col_in_819              ( col_in_819     ),
    .col_in_820              ( col_in_820     ),
    .col_in_821              ( col_in_821     ),
    .col_in_822              ( col_in_822     ),
    .col_in_823              ( col_in_823     ),
    .col_in_824              ( col_in_824     ),
    .col_in_825              ( col_in_825     ),
    .col_in_826              ( col_in_826     ),
    .col_in_827              ( col_in_827     ),
    .col_in_828              ( col_in_828     ),
    .col_in_829              ( col_in_829     ),
    .col_in_830              ( col_in_830     ),
    .col_in_831              ( col_in_831     ),
    .col_in_832              ( col_in_832     ),
    .col_in_833              ( col_in_833     ),
    .col_in_834              ( col_in_834     ),
    .col_in_835              ( col_in_835     ),
    .col_in_836              ( col_in_836     ),
    .col_in_837              ( col_in_837     ),
    .col_in_838              ( col_in_838     ),
    .col_in_839              ( col_in_839     ),
    .col_in_840              ( col_in_840     ),
    .col_in_841              ( col_in_841     ),
    .col_in_842              ( col_in_842     ),
    .col_in_843              ( col_in_843     ),
    .col_in_844              ( col_in_844     ),
    .col_in_845              ( col_in_845     ),
    .col_in_846              ( col_in_846     ),
    .col_in_847              ( col_in_847     ),
    .col_in_848              ( col_in_848     ),
    .col_in_849              ( col_in_849     ),
    .col_in_850              ( col_in_850     ),
    .col_in_851              ( col_in_851     ),
    .col_in_852              ( col_in_852     ),
    .col_in_853              ( col_in_853     ),
    .col_in_854              ( col_in_854     ),
    .col_in_855              ( col_in_855     ),
    .col_in_856              ( col_in_856     ),
    .col_in_857              ( col_in_857     ),
    .col_in_858              ( col_in_858     ),
    .col_in_859              ( col_in_859     ),
    .col_in_860              ( col_in_860     ),
    .col_in_861              ( col_in_861     ),
    .col_in_862              ( col_in_862     ),
    .col_in_863              ( col_in_863     ),
    .col_in_864              ( col_in_864     ),
    .col_in_865              ( col_in_865     ),
    .col_in_866              ( col_in_866     ),
    .col_in_867              ( col_in_867     ),
    .col_in_868              ( col_in_868     ),
    .col_in_869              ( col_in_869     ),
    .col_in_870              ( col_in_870     ),
    .col_in_871              ( col_in_871     ),
    .col_in_872              ( col_in_872     ),
    .col_in_873              ( col_in_873     ),
    .col_in_874              ( col_in_874     ),
    .col_in_875              ( col_in_875     ),
    .col_in_876              ( col_in_876     ),
    .col_in_877              ( col_in_877     ),
    .col_in_878              ( col_in_878     ),
    .col_in_879              ( col_in_879     ),
    .col_in_880              ( col_in_880     ),
    .col_in_881              ( col_in_881     ),
    .col_in_882              ( col_in_882     ),
    .col_in_883              ( col_in_883     ),
    .col_in_884              ( col_in_884     ),
    .col_in_885              ( col_in_885     ),
    .col_in_886              ( col_in_886     ),
    .col_in_887              ( col_in_887     ),
    .col_in_888              ( col_in_888     ),
    .col_in_889              ( col_in_889     ),
    .col_in_890              ( col_in_890     ),
    .col_in_891              ( col_in_891     ),
    .col_in_892              ( col_in_892     ),
    .col_in_893              ( col_in_893     ),
    .col_in_894              ( col_in_894     ),
    .col_in_895              ( col_in_895     ),
    .col_in_896              ( col_in_896     ),
    .col_in_897              ( col_in_897     ),
    .col_in_898              ( col_in_898     ),
    .col_in_899              ( col_in_899     ),
    .col_in_900              ( col_in_900     ),
    .col_in_901              ( col_in_901     ),
    .col_in_902              ( col_in_902     ),
    .col_in_903              ( col_in_903     ),
    .col_in_904              ( col_in_904     ),
    .col_in_905              ( col_in_905     ),
    .col_in_906              ( col_in_906     ),
    .col_in_907              ( col_in_907     ),
    .col_in_908              ( col_in_908     ),
    .col_in_909              ( col_in_909     ),
    .col_in_910              ( col_in_910     ),
    .col_in_911              ( col_in_911     ),
    .col_in_912              ( col_in_912     ),
    .col_in_913              ( col_in_913     ),
    .col_in_914              ( col_in_914     ),
    .col_in_915              ( col_in_915     ),
    .col_in_916              ( col_in_916     ),
    .col_in_917              ( col_in_917     ),
    .col_in_918              ( col_in_918     ),
    .col_in_919              ( col_in_919     ),
    .col_in_920              ( col_in_920     ),
    .col_in_921              ( col_in_921     ),
    .col_in_922              ( col_in_922     ),
    .col_in_923              ( col_in_923     ),
    .col_in_924              ( col_in_924     ),
    .col_in_925              ( col_in_925     ),
    .col_in_926              ( col_in_926     ),
    .col_in_927              ( col_in_927     ),
    .col_in_928              ( col_in_928     ),
    .col_in_929              ( col_in_929     ),
    .col_in_930              ( col_in_930     ),
    .col_in_931              ( col_in_931     ),
    .col_in_932              ( col_in_932     ),
    .col_in_933              ( col_in_933     ),
    .col_in_934              ( col_in_934     ),
    .col_in_935              ( col_in_935     ),
    .col_in_936              ( col_in_936     ),
    .col_in_937              ( col_in_937     ),
    .col_in_938              ( col_in_938     ),
    .col_in_939              ( col_in_939     ),
    .col_in_940              ( col_in_940     ),
    .col_in_941              ( col_in_941     ),
    .col_in_942              ( col_in_942     ),
    .col_in_943              ( col_in_943     ),
    .col_in_944              ( col_in_944     ),
    .col_in_945              ( col_in_945     ),
    .col_in_946              ( col_in_946     ),
    .col_in_947              ( col_in_947     ),
    .col_in_948              ( col_in_948     ),
    .col_in_949              ( col_in_949     ),
    .col_in_950              ( col_in_950     ),
    .col_in_951              ( col_in_951     ),
    .col_in_952              ( col_in_952     ),
    .col_in_953              ( col_in_953     ),
    .col_in_954              ( col_in_954     ),
    .col_in_955              ( col_in_955     ),
    .col_in_956              ( col_in_956     ),
    .col_in_957              ( col_in_957     ),
    .col_in_958              ( col_in_958     ),
    .col_in_959              ( col_in_959     ),
    .col_in_960              ( col_in_960     ),
    .col_in_961              ( col_in_961     ),
    .col_in_962              ( col_in_962     ),
    .col_in_963              ( col_in_963     ),
    .col_in_964              ( col_in_964     ),
    .col_in_965              ( col_in_965     ),
    .col_in_966              ( col_in_966     ),
    .col_in_967              ( col_in_967     ),
    .col_in_968              ( col_in_968     ),
    .col_in_969              ( col_in_969     ),
    .col_in_970              ( col_in_970     ),
    .col_in_971              ( col_in_971     ),
    .col_in_972              ( col_in_972     ),
    .col_in_973              ( col_in_973     ),
    .col_in_974              ( col_in_974     ),
    .col_in_975              ( col_in_975     ),
    .col_in_976              ( col_in_976     ),
    .col_in_977              ( col_in_977     ),
    .col_in_978              ( col_in_978     ),
    .col_in_979              ( col_in_979     ),
    .col_in_980              ( col_in_980     ),
    .col_in_981              ( col_in_981     ),
    .col_in_982              ( col_in_982     ),
    .col_in_983              ( col_in_983     ),
    .col_in_984              ( col_in_984     ),
    .col_in_985              ( col_in_985     ),
    .col_in_986              ( col_in_986     ),
    .col_in_987              ( col_in_987     ),
    .col_in_988              ( col_in_988     ),
    .col_in_989              ( col_in_989     ),
    .col_in_990              ( col_in_990     ),
    .col_in_991              ( col_in_991     ),
    .col_in_992              ( col_in_992     ),
    .col_in_993              ( col_in_993     ),
    .col_in_994              ( col_in_994     ),
    .col_in_995              ( col_in_995     ),
    .col_in_996              ( col_in_996     ),
    .col_in_997              ( col_in_997     ),
    .col_in_998              ( col_in_998     ),
    .col_in_999              ( col_in_999     ),
    .col_in_1000             ( col_in_1000    ),
    .col_in_1001             ( col_in_1001    ),
    .col_in_1002             ( col_in_1002    ),
    .col_in_1003             ( col_in_1003    ),
    .col_in_1004             ( col_in_1004    ),
    .col_in_1005             ( col_in_1005    ),
    .col_in_1006             ( col_in_1006    ),
    .col_in_1007             ( col_in_1007    ),
    .col_in_1008             ( col_in_1008    ),
    .col_in_1009             ( col_in_1009    ),
    .col_in_1010             ( col_in_1010    ),
    .col_in_1011             ( col_in_1011    ),
    .col_in_1012             ( col_in_1012    ),
    .col_in_1013             ( col_in_1013    ),
    .col_in_1014             ( col_in_1014    ),
    .col_in_1015             ( col_in_1015    ),
    .col_in_1016             ( col_in_1016    ),
    .col_in_1017             ( col_in_1017    ),
    .col_in_1018             ( col_in_1018    ),
    .col_in_1019             ( col_in_1019    ),
    .col_in_1020             ( col_in_1020    ),
    .col_in_1021             ( col_in_1021    ),
    .col_in_1022             ( col_in_1022    ),
    .col_in_1023             ( col_in_1023    ),

    .col_out_0               ( col_out_0      ),
    .col_out_1               ( col_out_1      ),
    .col_out_2               ( col_out_2      ),
    .col_out_3               ( col_out_3      ),
    .col_out_4               ( col_out_4      ),
    .col_out_5               ( col_out_5      ),
    .col_out_6               ( col_out_6      ),
    .col_out_7               ( col_out_7      ),
    .col_out_8               ( col_out_8      ),
    .col_out_9               ( col_out_9      ),
    .col_out_10              ( col_out_10     ),
    .col_out_11              ( col_out_11     ),
    .col_out_12              ( col_out_12     ),
    .col_out_13              ( col_out_13     ),
    .col_out_14              ( col_out_14     ),
    .col_out_15              ( col_out_15     ),
    .col_out_16              ( col_out_16     ),
    .col_out_17              ( col_out_17     ),
    .col_out_18              ( col_out_18     ),
    .col_out_19              ( col_out_19     ),
    .col_out_20              ( col_out_20     ),
    .col_out_21              ( col_out_21     ),
    .col_out_22              ( col_out_22     ),
    .col_out_23              ( col_out_23     ),
    .col_out_24              ( col_out_24     ),
    .col_out_25              ( col_out_25     ),
    .col_out_26              ( col_out_26     ),
    .col_out_27              ( col_out_27     ),
    .col_out_28              ( col_out_28     ),
    .col_out_29              ( col_out_29     ),
    .col_out_30              ( col_out_30     ),
    .col_out_31              ( col_out_31     ),
    .col_out_32              ( col_out_32     ),
    .col_out_33              ( col_out_33     ),
    .col_out_34              ( col_out_34     ),
    .col_out_35              ( col_out_35     ),
    .col_out_36              ( col_out_36     ),
    .col_out_37              ( col_out_37     ),
    .col_out_38              ( col_out_38     ),
    .col_out_39              ( col_out_39     ),
    .col_out_40              ( col_out_40     ),
    .col_out_41              ( col_out_41     ),
    .col_out_42              ( col_out_42     ),
    .col_out_43              ( col_out_43     ),
    .col_out_44              ( col_out_44     ),
    .col_out_45              ( col_out_45     ),
    .col_out_46              ( col_out_46     ),
    .col_out_47              ( col_out_47     ),
    .col_out_48              ( col_out_48     ),
    .col_out_49              ( col_out_49     ),
    .col_out_50              ( col_out_50     ),
    .col_out_51              ( col_out_51     ),
    .col_out_52              ( col_out_52     ),
    .col_out_53              ( col_out_53     ),
    .col_out_54              ( col_out_54     ),
    .col_out_55              ( col_out_55     ),
    .col_out_56              ( col_out_56     ),
    .col_out_57              ( col_out_57     ),
    .col_out_58              ( col_out_58     ),
    .col_out_59              ( col_out_59     ),
    .col_out_60              ( col_out_60     ),
    .col_out_61              ( col_out_61     ),
    .col_out_62              ( col_out_62     ),
    .col_out_63              ( col_out_63     ),
    .col_out_64              ( col_out_64     ),
    .col_out_65              ( col_out_65     ),
    .col_out_66              ( col_out_66     ),
    .col_out_67              ( col_out_67     ),
    .col_out_68              ( col_out_68     ),
    .col_out_69              ( col_out_69     ),
    .col_out_70              ( col_out_70     ),
    .col_out_71              ( col_out_71     ),
    .col_out_72              ( col_out_72     ),
    .col_out_73              ( col_out_73     ),
    .col_out_74              ( col_out_74     ),
    .col_out_75              ( col_out_75     ),
    .col_out_76              ( col_out_76     ),
    .col_out_77              ( col_out_77     ),
    .col_out_78              ( col_out_78     ),
    .col_out_79              ( col_out_79     ),
    .col_out_80              ( col_out_80     ),
    .col_out_81              ( col_out_81     ),
    .col_out_82              ( col_out_82     ),
    .col_out_83              ( col_out_83     ),
    .col_out_84              ( col_out_84     ),
    .col_out_85              ( col_out_85     ),
    .col_out_86              ( col_out_86     ),
    .col_out_87              ( col_out_87     ),
    .col_out_88              ( col_out_88     ),
    .col_out_89              ( col_out_89     ),
    .col_out_90              ( col_out_90     ),
    .col_out_91              ( col_out_91     ),
    .col_out_92              ( col_out_92     ),
    .col_out_93              ( col_out_93     ),
    .col_out_94              ( col_out_94     ),
    .col_out_95              ( col_out_95     ),
    .col_out_96              ( col_out_96     ),
    .col_out_97              ( col_out_97     ),
    .col_out_98              ( col_out_98     ),
    .col_out_99              ( col_out_99     ),
    .col_out_100             ( col_out_100    ),
    .col_out_101             ( col_out_101    ),
    .col_out_102             ( col_out_102    ),
    .col_out_103             ( col_out_103    ),
    .col_out_104             ( col_out_104    ),
    .col_out_105             ( col_out_105    ),
    .col_out_106             ( col_out_106    ),
    .col_out_107             ( col_out_107    ),
    .col_out_108             ( col_out_108    ),
    .col_out_109             ( col_out_109    ),
    .col_out_110             ( col_out_110    ),
    .col_out_111             ( col_out_111    ),
    .col_out_112             ( col_out_112    ),
    .col_out_113             ( col_out_113    ),
    .col_out_114             ( col_out_114    ),
    .col_out_115             ( col_out_115    ),
    .col_out_116             ( col_out_116    ),
    .col_out_117             ( col_out_117    ),
    .col_out_118             ( col_out_118    ),
    .col_out_119             ( col_out_119    ),
    .col_out_120             ( col_out_120    ),
    .col_out_121             ( col_out_121    ),
    .col_out_122             ( col_out_122    ),
    .col_out_123             ( col_out_123    ),
    .col_out_124             ( col_out_124    ),
    .col_out_125             ( col_out_125    ),
    .col_out_126             ( col_out_126    ),
    .col_out_127             ( col_out_127    ),
    .col_out_128             ( col_out_128    ),
    .col_out_129             ( col_out_129    ),
    .col_out_130             ( col_out_130    ),
    .col_out_131             ( col_out_131    ),
    .col_out_132             ( col_out_132    ),
    .col_out_133             ( col_out_133    ),
    .col_out_134             ( col_out_134    ),
    .col_out_135             ( col_out_135    ),
    .col_out_136             ( col_out_136    ),
    .col_out_137             ( col_out_137    ),
    .col_out_138             ( col_out_138    ),
    .col_out_139             ( col_out_139    ),
    .col_out_140             ( col_out_140    ),
    .col_out_141             ( col_out_141    ),
    .col_out_142             ( col_out_142    ),
    .col_out_143             ( col_out_143    ),
    .col_out_144             ( col_out_144    ),
    .col_out_145             ( col_out_145    ),
    .col_out_146             ( col_out_146    ),
    .col_out_147             ( col_out_147    ),
    .col_out_148             ( col_out_148    ),
    .col_out_149             ( col_out_149    ),
    .col_out_150             ( col_out_150    ),
    .col_out_151             ( col_out_151    ),
    .col_out_152             ( col_out_152    ),
    .col_out_153             ( col_out_153    ),
    .col_out_154             ( col_out_154    ),
    .col_out_155             ( col_out_155    ),
    .col_out_156             ( col_out_156    ),
    .col_out_157             ( col_out_157    ),
    .col_out_158             ( col_out_158    ),
    .col_out_159             ( col_out_159    ),
    .col_out_160             ( col_out_160    ),
    .col_out_161             ( col_out_161    ),
    .col_out_162             ( col_out_162    ),
    .col_out_163             ( col_out_163    ),
    .col_out_164             ( col_out_164    ),
    .col_out_165             ( col_out_165    ),
    .col_out_166             ( col_out_166    ),
    .col_out_167             ( col_out_167    ),
    .col_out_168             ( col_out_168    ),
    .col_out_169             ( col_out_169    ),
    .col_out_170             ( col_out_170    ),
    .col_out_171             ( col_out_171    ),
    .col_out_172             ( col_out_172    ),
    .col_out_173             ( col_out_173    ),
    .col_out_174             ( col_out_174    ),
    .col_out_175             ( col_out_175    ),
    .col_out_176             ( col_out_176    ),
    .col_out_177             ( col_out_177    ),
    .col_out_178             ( col_out_178    ),
    .col_out_179             ( col_out_179    ),
    .col_out_180             ( col_out_180    ),
    .col_out_181             ( col_out_181    ),
    .col_out_182             ( col_out_182    ),
    .col_out_183             ( col_out_183    ),
    .col_out_184             ( col_out_184    ),
    .col_out_185             ( col_out_185    ),
    .col_out_186             ( col_out_186    ),
    .col_out_187             ( col_out_187    ),
    .col_out_188             ( col_out_188    ),
    .col_out_189             ( col_out_189    ),
    .col_out_190             ( col_out_190    ),
    .col_out_191             ( col_out_191    ),
    .col_out_192             ( col_out_192    ),
    .col_out_193             ( col_out_193    ),
    .col_out_194             ( col_out_194    ),
    .col_out_195             ( col_out_195    ),
    .col_out_196             ( col_out_196    ),
    .col_out_197             ( col_out_197    ),
    .col_out_198             ( col_out_198    ),
    .col_out_199             ( col_out_199    ),
    .col_out_200             ( col_out_200    ),
    .col_out_201             ( col_out_201    ),
    .col_out_202             ( col_out_202    ),
    .col_out_203             ( col_out_203    ),
    .col_out_204             ( col_out_204    ),
    .col_out_205             ( col_out_205    ),
    .col_out_206             ( col_out_206    ),
    .col_out_207             ( col_out_207    ),
    .col_out_208             ( col_out_208    ),
    .col_out_209             ( col_out_209    ),
    .col_out_210             ( col_out_210    ),
    .col_out_211             ( col_out_211    ),
    .col_out_212             ( col_out_212    ),
    .col_out_213             ( col_out_213    ),
    .col_out_214             ( col_out_214    ),
    .col_out_215             ( col_out_215    ),
    .col_out_216             ( col_out_216    ),
    .col_out_217             ( col_out_217    ),
    .col_out_218             ( col_out_218    ),
    .col_out_219             ( col_out_219    ),
    .col_out_220             ( col_out_220    ),
    .col_out_221             ( col_out_221    ),
    .col_out_222             ( col_out_222    ),
    .col_out_223             ( col_out_223    ),
    .col_out_224             ( col_out_224    ),
    .col_out_225             ( col_out_225    ),
    .col_out_226             ( col_out_226    ),
    .col_out_227             ( col_out_227    ),
    .col_out_228             ( col_out_228    ),
    .col_out_229             ( col_out_229    ),
    .col_out_230             ( col_out_230    ),
    .col_out_231             ( col_out_231    ),
    .col_out_232             ( col_out_232    ),
    .col_out_233             ( col_out_233    ),
    .col_out_234             ( col_out_234    ),
    .col_out_235             ( col_out_235    ),
    .col_out_236             ( col_out_236    ),
    .col_out_237             ( col_out_237    ),
    .col_out_238             ( col_out_238    ),
    .col_out_239             ( col_out_239    ),
    .col_out_240             ( col_out_240    ),
    .col_out_241             ( col_out_241    ),
    .col_out_242             ( col_out_242    ),
    .col_out_243             ( col_out_243    ),
    .col_out_244             ( col_out_244    ),
    .col_out_245             ( col_out_245    ),
    .col_out_246             ( col_out_246    ),
    .col_out_247             ( col_out_247    ),
    .col_out_248             ( col_out_248    ),
    .col_out_249             ( col_out_249    ),
    .col_out_250             ( col_out_250    ),
    .col_out_251             ( col_out_251    ),
    .col_out_252             ( col_out_252    ),
    .col_out_253             ( col_out_253    ),
    .col_out_254             ( col_out_254    ),
    .col_out_255             ( col_out_255    ),
    .col_out_256             ( col_out_256    ),
    .col_out_257             ( col_out_257    ),
    .col_out_258             ( col_out_258    ),
    .col_out_259             ( col_out_259    ),
    .col_out_260             ( col_out_260    ),
    .col_out_261             ( col_out_261    ),
    .col_out_262             ( col_out_262    ),
    .col_out_263             ( col_out_263    ),
    .col_out_264             ( col_out_264    ),
    .col_out_265             ( col_out_265    ),
    .col_out_266             ( col_out_266    ),
    .col_out_267             ( col_out_267    ),
    .col_out_268             ( col_out_268    ),
    .col_out_269             ( col_out_269    ),
    .col_out_270             ( col_out_270    ),
    .col_out_271             ( col_out_271    ),
    .col_out_272             ( col_out_272    ),
    .col_out_273             ( col_out_273    ),
    .col_out_274             ( col_out_274    ),
    .col_out_275             ( col_out_275    ),
    .col_out_276             ( col_out_276    ),
    .col_out_277             ( col_out_277    ),
    .col_out_278             ( col_out_278    ),
    .col_out_279             ( col_out_279    ),
    .col_out_280             ( col_out_280    ),
    .col_out_281             ( col_out_281    ),
    .col_out_282             ( col_out_282    ),
    .col_out_283             ( col_out_283    ),
    .col_out_284             ( col_out_284    ),
    .col_out_285             ( col_out_285    ),
    .col_out_286             ( col_out_286    ),
    .col_out_287             ( col_out_287    ),
    .col_out_288             ( col_out_288    ),
    .col_out_289             ( col_out_289    ),
    .col_out_290             ( col_out_290    ),
    .col_out_291             ( col_out_291    ),
    .col_out_292             ( col_out_292    ),
    .col_out_293             ( col_out_293    ),
    .col_out_294             ( col_out_294    ),
    .col_out_295             ( col_out_295    ),
    .col_out_296             ( col_out_296    ),
    .col_out_297             ( col_out_297    ),
    .col_out_298             ( col_out_298    ),
    .col_out_299             ( col_out_299    ),
    .col_out_300             ( col_out_300    ),
    .col_out_301             ( col_out_301    ),
    .col_out_302             ( col_out_302    ),
    .col_out_303             ( col_out_303    ),
    .col_out_304             ( col_out_304    ),
    .col_out_305             ( col_out_305    ),
    .col_out_306             ( col_out_306    ),
    .col_out_307             ( col_out_307    ),
    .col_out_308             ( col_out_308    ),
    .col_out_309             ( col_out_309    ),
    .col_out_310             ( col_out_310    ),
    .col_out_311             ( col_out_311    ),
    .col_out_312             ( col_out_312    ),
    .col_out_313             ( col_out_313    ),
    .col_out_314             ( col_out_314    ),
    .col_out_315             ( col_out_315    ),
    .col_out_316             ( col_out_316    ),
    .col_out_317             ( col_out_317    ),
    .col_out_318             ( col_out_318    ),
    .col_out_319             ( col_out_319    ),
    .col_out_320             ( col_out_320    ),
    .col_out_321             ( col_out_321    ),
    .col_out_322             ( col_out_322    ),
    .col_out_323             ( col_out_323    ),
    .col_out_324             ( col_out_324    ),
    .col_out_325             ( col_out_325    ),
    .col_out_326             ( col_out_326    ),
    .col_out_327             ( col_out_327    ),
    .col_out_328             ( col_out_328    ),
    .col_out_329             ( col_out_329    ),
    .col_out_330             ( col_out_330    ),
    .col_out_331             ( col_out_331    ),
    .col_out_332             ( col_out_332    ),
    .col_out_333             ( col_out_333    ),
    .col_out_334             ( col_out_334    ),
    .col_out_335             ( col_out_335    ),
    .col_out_336             ( col_out_336    ),
    .col_out_337             ( col_out_337    ),
    .col_out_338             ( col_out_338    ),
    .col_out_339             ( col_out_339    ),
    .col_out_340             ( col_out_340    ),
    .col_out_341             ( col_out_341    ),
    .col_out_342             ( col_out_342    ),
    .col_out_343             ( col_out_343    ),
    .col_out_344             ( col_out_344    ),
    .col_out_345             ( col_out_345    ),
    .col_out_346             ( col_out_346    ),
    .col_out_347             ( col_out_347    ),
    .col_out_348             ( col_out_348    ),
    .col_out_349             ( col_out_349    ),
    .col_out_350             ( col_out_350    ),
    .col_out_351             ( col_out_351    ),
    .col_out_352             ( col_out_352    ),
    .col_out_353             ( col_out_353    ),
    .col_out_354             ( col_out_354    ),
    .col_out_355             ( col_out_355    ),
    .col_out_356             ( col_out_356    ),
    .col_out_357             ( col_out_357    ),
    .col_out_358             ( col_out_358    ),
    .col_out_359             ( col_out_359    ),
    .col_out_360             ( col_out_360    ),
    .col_out_361             ( col_out_361    ),
    .col_out_362             ( col_out_362    ),
    .col_out_363             ( col_out_363    ),
    .col_out_364             ( col_out_364    ),
    .col_out_365             ( col_out_365    ),
    .col_out_366             ( col_out_366    ),
    .col_out_367             ( col_out_367    ),
    .col_out_368             ( col_out_368    ),
    .col_out_369             ( col_out_369    ),
    .col_out_370             ( col_out_370    ),
    .col_out_371             ( col_out_371    ),
    .col_out_372             ( col_out_372    ),
    .col_out_373             ( col_out_373    ),
    .col_out_374             ( col_out_374    ),
    .col_out_375             ( col_out_375    ),
    .col_out_376             ( col_out_376    ),
    .col_out_377             ( col_out_377    ),
    .col_out_378             ( col_out_378    ),
    .col_out_379             ( col_out_379    ),
    .col_out_380             ( col_out_380    ),
    .col_out_381             ( col_out_381    ),
    .col_out_382             ( col_out_382    ),
    .col_out_383             ( col_out_383    ),
    .col_out_384             ( col_out_384    ),
    .col_out_385             ( col_out_385    ),
    .col_out_386             ( col_out_386    ),
    .col_out_387             ( col_out_387    ),
    .col_out_388             ( col_out_388    ),
    .col_out_389             ( col_out_389    ),
    .col_out_390             ( col_out_390    ),
    .col_out_391             ( col_out_391    ),
    .col_out_392             ( col_out_392    ),
    .col_out_393             ( col_out_393    ),
    .col_out_394             ( col_out_394    ),
    .col_out_395             ( col_out_395    ),
    .col_out_396             ( col_out_396    ),
    .col_out_397             ( col_out_397    ),
    .col_out_398             ( col_out_398    ),
    .col_out_399             ( col_out_399    ),
    .col_out_400             ( col_out_400    ),
    .col_out_401             ( col_out_401    ),
    .col_out_402             ( col_out_402    ),
    .col_out_403             ( col_out_403    ),
    .col_out_404             ( col_out_404    ),
    .col_out_405             ( col_out_405    ),
    .col_out_406             ( col_out_406    ),
    .col_out_407             ( col_out_407    ),
    .col_out_408             ( col_out_408    ),
    .col_out_409             ( col_out_409    ),
    .col_out_410             ( col_out_410    ),
    .col_out_411             ( col_out_411    ),
    .col_out_412             ( col_out_412    ),
    .col_out_413             ( col_out_413    ),
    .col_out_414             ( col_out_414    ),
    .col_out_415             ( col_out_415    ),
    .col_out_416             ( col_out_416    ),
    .col_out_417             ( col_out_417    ),
    .col_out_418             ( col_out_418    ),
    .col_out_419             ( col_out_419    ),
    .col_out_420             ( col_out_420    ),
    .col_out_421             ( col_out_421    ),
    .col_out_422             ( col_out_422    ),
    .col_out_423             ( col_out_423    ),
    .col_out_424             ( col_out_424    ),
    .col_out_425             ( col_out_425    ),
    .col_out_426             ( col_out_426    ),
    .col_out_427             ( col_out_427    ),
    .col_out_428             ( col_out_428    ),
    .col_out_429             ( col_out_429    ),
    .col_out_430             ( col_out_430    ),
    .col_out_431             ( col_out_431    ),
    .col_out_432             ( col_out_432    ),
    .col_out_433             ( col_out_433    ),
    .col_out_434             ( col_out_434    ),
    .col_out_435             ( col_out_435    ),
    .col_out_436             ( col_out_436    ),
    .col_out_437             ( col_out_437    ),
    .col_out_438             ( col_out_438    ),
    .col_out_439             ( col_out_439    ),
    .col_out_440             ( col_out_440    ),
    .col_out_441             ( col_out_441    ),
    .col_out_442             ( col_out_442    ),
    .col_out_443             ( col_out_443    ),
    .col_out_444             ( col_out_444    ),
    .col_out_445             ( col_out_445    ),
    .col_out_446             ( col_out_446    ),
    .col_out_447             ( col_out_447    ),
    .col_out_448             ( col_out_448    ),
    .col_out_449             ( col_out_449    ),
    .col_out_450             ( col_out_450    ),
    .col_out_451             ( col_out_451    ),
    .col_out_452             ( col_out_452    ),
    .col_out_453             ( col_out_453    ),
    .col_out_454             ( col_out_454    ),
    .col_out_455             ( col_out_455    ),
    .col_out_456             ( col_out_456    ),
    .col_out_457             ( col_out_457    ),
    .col_out_458             ( col_out_458    ),
    .col_out_459             ( col_out_459    ),
    .col_out_460             ( col_out_460    ),
    .col_out_461             ( col_out_461    ),
    .col_out_462             ( col_out_462    ),
    .col_out_463             ( col_out_463    ),
    .col_out_464             ( col_out_464    ),
    .col_out_465             ( col_out_465    ),
    .col_out_466             ( col_out_466    ),
    .col_out_467             ( col_out_467    ),
    .col_out_468             ( col_out_468    ),
    .col_out_469             ( col_out_469    ),
    .col_out_470             ( col_out_470    ),
    .col_out_471             ( col_out_471    ),
    .col_out_472             ( col_out_472    ),
    .col_out_473             ( col_out_473    ),
    .col_out_474             ( col_out_474    ),
    .col_out_475             ( col_out_475    ),
    .col_out_476             ( col_out_476    ),
    .col_out_477             ( col_out_477    ),
    .col_out_478             ( col_out_478    ),
    .col_out_479             ( col_out_479    ),
    .col_out_480             ( col_out_480    ),
    .col_out_481             ( col_out_481    ),
    .col_out_482             ( col_out_482    ),
    .col_out_483             ( col_out_483    ),
    .col_out_484             ( col_out_484    ),
    .col_out_485             ( col_out_485    ),
    .col_out_486             ( col_out_486    ),
    .col_out_487             ( col_out_487    ),
    .col_out_488             ( col_out_488    ),
    .col_out_489             ( col_out_489    ),
    .col_out_490             ( col_out_490    ),
    .col_out_491             ( col_out_491    ),
    .col_out_492             ( col_out_492    ),
    .col_out_493             ( col_out_493    ),
    .col_out_494             ( col_out_494    ),
    .col_out_495             ( col_out_495    ),
    .col_out_496             ( col_out_496    ),
    .col_out_497             ( col_out_497    ),
    .col_out_498             ( col_out_498    ),
    .col_out_499             ( col_out_499    ),
    .col_out_500             ( col_out_500    ),
    .col_out_501             ( col_out_501    ),
    .col_out_502             ( col_out_502    ),
    .col_out_503             ( col_out_503    ),
    .col_out_504             ( col_out_504    ),
    .col_out_505             ( col_out_505    ),
    .col_out_506             ( col_out_506    ),
    .col_out_507             ( col_out_507    ),
    .col_out_508             ( col_out_508    ),
    .col_out_509             ( col_out_509    ),
    .col_out_510             ( col_out_510    ),
    .col_out_511             ( col_out_511    ),
    .col_out_512             ( col_out_512    ),
    .col_out_513             ( col_out_513    ),
    .col_out_514             ( col_out_514    ),
    .col_out_515             ( col_out_515    ),
    .col_out_516             ( col_out_516    ),
    .col_out_517             ( col_out_517    ),
    .col_out_518             ( col_out_518    ),
    .col_out_519             ( col_out_519    ),
    .col_out_520             ( col_out_520    ),
    .col_out_521             ( col_out_521    ),
    .col_out_522             ( col_out_522    ),
    .col_out_523             ( col_out_523    ),
    .col_out_524             ( col_out_524    ),
    .col_out_525             ( col_out_525    ),
    .col_out_526             ( col_out_526    ),
    .col_out_527             ( col_out_527    ),
    .col_out_528             ( col_out_528    ),
    .col_out_529             ( col_out_529    ),
    .col_out_530             ( col_out_530    ),
    .col_out_531             ( col_out_531    ),
    .col_out_532             ( col_out_532    ),
    .col_out_533             ( col_out_533    ),
    .col_out_534             ( col_out_534    ),
    .col_out_535             ( col_out_535    ),
    .col_out_536             ( col_out_536    ),
    .col_out_537             ( col_out_537    ),
    .col_out_538             ( col_out_538    ),
    .col_out_539             ( col_out_539    ),
    .col_out_540             ( col_out_540    ),
    .col_out_541             ( col_out_541    ),
    .col_out_542             ( col_out_542    ),
    .col_out_543             ( col_out_543    ),
    .col_out_544             ( col_out_544    ),
    .col_out_545             ( col_out_545    ),
    .col_out_546             ( col_out_546    ),
    .col_out_547             ( col_out_547    ),
    .col_out_548             ( col_out_548    ),
    .col_out_549             ( col_out_549    ),
    .col_out_550             ( col_out_550    ),
    .col_out_551             ( col_out_551    ),
    .col_out_552             ( col_out_552    ),
    .col_out_553             ( col_out_553    ),
    .col_out_554             ( col_out_554    ),
    .col_out_555             ( col_out_555    ),
    .col_out_556             ( col_out_556    ),
    .col_out_557             ( col_out_557    ),
    .col_out_558             ( col_out_558    ),
    .col_out_559             ( col_out_559    ),
    .col_out_560             ( col_out_560    ),
    .col_out_561             ( col_out_561    ),
    .col_out_562             ( col_out_562    ),
    .col_out_563             ( col_out_563    ),
    .col_out_564             ( col_out_564    ),
    .col_out_565             ( col_out_565    ),
    .col_out_566             ( col_out_566    ),
    .col_out_567             ( col_out_567    ),
    .col_out_568             ( col_out_568    ),
    .col_out_569             ( col_out_569    ),
    .col_out_570             ( col_out_570    ),
    .col_out_571             ( col_out_571    ),
    .col_out_572             ( col_out_572    ),
    .col_out_573             ( col_out_573    ),
    .col_out_574             ( col_out_574    ),
    .col_out_575             ( col_out_575    ),
    .col_out_576             ( col_out_576    ),
    .col_out_577             ( col_out_577    ),
    .col_out_578             ( col_out_578    ),
    .col_out_579             ( col_out_579    ),
    .col_out_580             ( col_out_580    ),
    .col_out_581             ( col_out_581    ),
    .col_out_582             ( col_out_582    ),
    .col_out_583             ( col_out_583    ),
    .col_out_584             ( col_out_584    ),
    .col_out_585             ( col_out_585    ),
    .col_out_586             ( col_out_586    ),
    .col_out_587             ( col_out_587    ),
    .col_out_588             ( col_out_588    ),
    .col_out_589             ( col_out_589    ),
    .col_out_590             ( col_out_590    ),
    .col_out_591             ( col_out_591    ),
    .col_out_592             ( col_out_592    ),
    .col_out_593             ( col_out_593    ),
    .col_out_594             ( col_out_594    ),
    .col_out_595             ( col_out_595    ),
    .col_out_596             ( col_out_596    ),
    .col_out_597             ( col_out_597    ),
    .col_out_598             ( col_out_598    ),
    .col_out_599             ( col_out_599    ),
    .col_out_600             ( col_out_600    ),
    .col_out_601             ( col_out_601    ),
    .col_out_602             ( col_out_602    ),
    .col_out_603             ( col_out_603    ),
    .col_out_604             ( col_out_604    ),
    .col_out_605             ( col_out_605    ),
    .col_out_606             ( col_out_606    ),
    .col_out_607             ( col_out_607    ),
    .col_out_608             ( col_out_608    ),
    .col_out_609             ( col_out_609    ),
    .col_out_610             ( col_out_610    ),
    .col_out_611             ( col_out_611    ),
    .col_out_612             ( col_out_612    ),
    .col_out_613             ( col_out_613    ),
    .col_out_614             ( col_out_614    ),
    .col_out_615             ( col_out_615    ),
    .col_out_616             ( col_out_616    ),
    .col_out_617             ( col_out_617    ),
    .col_out_618             ( col_out_618    ),
    .col_out_619             ( col_out_619    ),
    .col_out_620             ( col_out_620    ),
    .col_out_621             ( col_out_621    ),
    .col_out_622             ( col_out_622    ),
    .col_out_623             ( col_out_623    ),
    .col_out_624             ( col_out_624    ),
    .col_out_625             ( col_out_625    ),
    .col_out_626             ( col_out_626    ),
    .col_out_627             ( col_out_627    ),
    .col_out_628             ( col_out_628    ),
    .col_out_629             ( col_out_629    ),
    .col_out_630             ( col_out_630    ),
    .col_out_631             ( col_out_631    ),
    .col_out_632             ( col_out_632    ),
    .col_out_633             ( col_out_633    ),
    .col_out_634             ( col_out_634    ),
    .col_out_635             ( col_out_635    ),
    .col_out_636             ( col_out_636    ),
    .col_out_637             ( col_out_637    ),
    .col_out_638             ( col_out_638    ),
    .col_out_639             ( col_out_639    ),
    .col_out_640             ( col_out_640    ),
    .col_out_641             ( col_out_641    ),
    .col_out_642             ( col_out_642    ),
    .col_out_643             ( col_out_643    ),
    .col_out_644             ( col_out_644    ),
    .col_out_645             ( col_out_645    ),
    .col_out_646             ( col_out_646    ),
    .col_out_647             ( col_out_647    ),
    .col_out_648             ( col_out_648    ),
    .col_out_649             ( col_out_649    ),
    .col_out_650             ( col_out_650    ),
    .col_out_651             ( col_out_651    ),
    .col_out_652             ( col_out_652    ),
    .col_out_653             ( col_out_653    ),
    .col_out_654             ( col_out_654    ),
    .col_out_655             ( col_out_655    ),
    .col_out_656             ( col_out_656    ),
    .col_out_657             ( col_out_657    ),
    .col_out_658             ( col_out_658    ),
    .col_out_659             ( col_out_659    ),
    .col_out_660             ( col_out_660    ),
    .col_out_661             ( col_out_661    ),
    .col_out_662             ( col_out_662    ),
    .col_out_663             ( col_out_663    ),
    .col_out_664             ( col_out_664    ),
    .col_out_665             ( col_out_665    ),
    .col_out_666             ( col_out_666    ),
    .col_out_667             ( col_out_667    ),
    .col_out_668             ( col_out_668    ),
    .col_out_669             ( col_out_669    ),
    .col_out_670             ( col_out_670    ),
    .col_out_671             ( col_out_671    ),
    .col_out_672             ( col_out_672    ),
    .col_out_673             ( col_out_673    ),
    .col_out_674             ( col_out_674    ),
    .col_out_675             ( col_out_675    ),
    .col_out_676             ( col_out_676    ),
    .col_out_677             ( col_out_677    ),
    .col_out_678             ( col_out_678    ),
    .col_out_679             ( col_out_679    ),
    .col_out_680             ( col_out_680    ),
    .col_out_681             ( col_out_681    ),
    .col_out_682             ( col_out_682    ),
    .col_out_683             ( col_out_683    ),
    .col_out_684             ( col_out_684    ),
    .col_out_685             ( col_out_685    ),
    .col_out_686             ( col_out_686    ),
    .col_out_687             ( col_out_687    ),
    .col_out_688             ( col_out_688    ),
    .col_out_689             ( col_out_689    ),
    .col_out_690             ( col_out_690    ),
    .col_out_691             ( col_out_691    ),
    .col_out_692             ( col_out_692    ),
    .col_out_693             ( col_out_693    ),
    .col_out_694             ( col_out_694    ),
    .col_out_695             ( col_out_695    ),
    .col_out_696             ( col_out_696    ),
    .col_out_697             ( col_out_697    ),
    .col_out_698             ( col_out_698    ),
    .col_out_699             ( col_out_699    ),
    .col_out_700             ( col_out_700    ),
    .col_out_701             ( col_out_701    ),
    .col_out_702             ( col_out_702    ),
    .col_out_703             ( col_out_703    ),
    .col_out_704             ( col_out_704    ),
    .col_out_705             ( col_out_705    ),
    .col_out_706             ( col_out_706    ),
    .col_out_707             ( col_out_707    ),
    .col_out_708             ( col_out_708    ),
    .col_out_709             ( col_out_709    ),
    .col_out_710             ( col_out_710    ),
    .col_out_711             ( col_out_711    ),
    .col_out_712             ( col_out_712    ),
    .col_out_713             ( col_out_713    ),
    .col_out_714             ( col_out_714    ),
    .col_out_715             ( col_out_715    ),
    .col_out_716             ( col_out_716    ),
    .col_out_717             ( col_out_717    ),
    .col_out_718             ( col_out_718    ),
    .col_out_719             ( col_out_719    ),
    .col_out_720             ( col_out_720    ),
    .col_out_721             ( col_out_721    ),
    .col_out_722             ( col_out_722    ),
    .col_out_723             ( col_out_723    ),
    .col_out_724             ( col_out_724    ),
    .col_out_725             ( col_out_725    ),
    .col_out_726             ( col_out_726    ),
    .col_out_727             ( col_out_727    ),
    .col_out_728             ( col_out_728    ),
    .col_out_729             ( col_out_729    ),
    .col_out_730             ( col_out_730    ),
    .col_out_731             ( col_out_731    ),
    .col_out_732             ( col_out_732    ),
    .col_out_733             ( col_out_733    ),
    .col_out_734             ( col_out_734    ),
    .col_out_735             ( col_out_735    ),
    .col_out_736             ( col_out_736    ),
    .col_out_737             ( col_out_737    ),
    .col_out_738             ( col_out_738    ),
    .col_out_739             ( col_out_739    ),
    .col_out_740             ( col_out_740    ),
    .col_out_741             ( col_out_741    ),
    .col_out_742             ( col_out_742    ),
    .col_out_743             ( col_out_743    ),
    .col_out_744             ( col_out_744    ),
    .col_out_745             ( col_out_745    ),
    .col_out_746             ( col_out_746    ),
    .col_out_747             ( col_out_747    ),
    .col_out_748             ( col_out_748    ),
    .col_out_749             ( col_out_749    ),
    .col_out_750             ( col_out_750    ),
    .col_out_751             ( col_out_751    ),
    .col_out_752             ( col_out_752    ),
    .col_out_753             ( col_out_753    ),
    .col_out_754             ( col_out_754    ),
    .col_out_755             ( col_out_755    ),
    .col_out_756             ( col_out_756    ),
    .col_out_757             ( col_out_757    ),
    .col_out_758             ( col_out_758    ),
    .col_out_759             ( col_out_759    ),
    .col_out_760             ( col_out_760    ),
    .col_out_761             ( col_out_761    ),
    .col_out_762             ( col_out_762    ),
    .col_out_763             ( col_out_763    ),
    .col_out_764             ( col_out_764    ),
    .col_out_765             ( col_out_765    ),
    .col_out_766             ( col_out_766    ),
    .col_out_767             ( col_out_767    ),
    .col_out_768             ( col_out_768    ),
    .col_out_769             ( col_out_769    ),
    .col_out_770             ( col_out_770    ),
    .col_out_771             ( col_out_771    ),
    .col_out_772             ( col_out_772    ),
    .col_out_773             ( col_out_773    ),
    .col_out_774             ( col_out_774    ),
    .col_out_775             ( col_out_775    ),
    .col_out_776             ( col_out_776    ),
    .col_out_777             ( col_out_777    ),
    .col_out_778             ( col_out_778    ),
    .col_out_779             ( col_out_779    ),
    .col_out_780             ( col_out_780    ),
    .col_out_781             ( col_out_781    ),
    .col_out_782             ( col_out_782    ),
    .col_out_783             ( col_out_783    ),
    .col_out_784             ( col_out_784    ),
    .col_out_785             ( col_out_785    ),
    .col_out_786             ( col_out_786    ),
    .col_out_787             ( col_out_787    ),
    .col_out_788             ( col_out_788    ),
    .col_out_789             ( col_out_789    ),
    .col_out_790             ( col_out_790    ),
    .col_out_791             ( col_out_791    ),
    .col_out_792             ( col_out_792    ),
    .col_out_793             ( col_out_793    ),
    .col_out_794             ( col_out_794    ),
    .col_out_795             ( col_out_795    ),
    .col_out_796             ( col_out_796    ),
    .col_out_797             ( col_out_797    ),
    .col_out_798             ( col_out_798    ),
    .col_out_799             ( col_out_799    ),
    .col_out_800             ( col_out_800    ),
    .col_out_801             ( col_out_801    ),
    .col_out_802             ( col_out_802    ),
    .col_out_803             ( col_out_803    ),
    .col_out_804             ( col_out_804    ),
    .col_out_805             ( col_out_805    ),
    .col_out_806             ( col_out_806    ),
    .col_out_807             ( col_out_807    ),
    .col_out_808             ( col_out_808    ),
    .col_out_809             ( col_out_809    ),
    .col_out_810             ( col_out_810    ),
    .col_out_811             ( col_out_811    ),
    .col_out_812             ( col_out_812    ),
    .col_out_813             ( col_out_813    ),
    .col_out_814             ( col_out_814    ),
    .col_out_815             ( col_out_815    ),
    .col_out_816             ( col_out_816    ),
    .col_out_817             ( col_out_817    ),
    .col_out_818             ( col_out_818    ),
    .col_out_819             ( col_out_819    ),
    .col_out_820             ( col_out_820    ),
    .col_out_821             ( col_out_821    ),
    .col_out_822             ( col_out_822    ),
    .col_out_823             ( col_out_823    ),
    .col_out_824             ( col_out_824    ),
    .col_out_825             ( col_out_825    ),
    .col_out_826             ( col_out_826    ),
    .col_out_827             ( col_out_827    ),
    .col_out_828             ( col_out_828    ),
    .col_out_829             ( col_out_829    ),
    .col_out_830             ( col_out_830    ),
    .col_out_831             ( col_out_831    ),
    .col_out_832             ( col_out_832    ),
    .col_out_833             ( col_out_833    ),
    .col_out_834             ( col_out_834    ),
    .col_out_835             ( col_out_835    ),
    .col_out_836             ( col_out_836    ),
    .col_out_837             ( col_out_837    ),
    .col_out_838             ( col_out_838    ),
    .col_out_839             ( col_out_839    ),
    .col_out_840             ( col_out_840    ),
    .col_out_841             ( col_out_841    ),
    .col_out_842             ( col_out_842    ),
    .col_out_843             ( col_out_843    ),
    .col_out_844             ( col_out_844    ),
    .col_out_845             ( col_out_845    ),
    .col_out_846             ( col_out_846    ),
    .col_out_847             ( col_out_847    ),
    .col_out_848             ( col_out_848    ),
    .col_out_849             ( col_out_849    ),
    .col_out_850             ( col_out_850    ),
    .col_out_851             ( col_out_851    ),
    .col_out_852             ( col_out_852    ),
    .col_out_853             ( col_out_853    ),
    .col_out_854             ( col_out_854    ),
    .col_out_855             ( col_out_855    ),
    .col_out_856             ( col_out_856    ),
    .col_out_857             ( col_out_857    ),
    .col_out_858             ( col_out_858    ),
    .col_out_859             ( col_out_859    ),
    .col_out_860             ( col_out_860    ),
    .col_out_861             ( col_out_861    ),
    .col_out_862             ( col_out_862    ),
    .col_out_863             ( col_out_863    ),
    .col_out_864             ( col_out_864    ),
    .col_out_865             ( col_out_865    ),
    .col_out_866             ( col_out_866    ),
    .col_out_867             ( col_out_867    ),
    .col_out_868             ( col_out_868    ),
    .col_out_869             ( col_out_869    ),
    .col_out_870             ( col_out_870    ),
    .col_out_871             ( col_out_871    ),
    .col_out_872             ( col_out_872    ),
    .col_out_873             ( col_out_873    ),
    .col_out_874             ( col_out_874    ),
    .col_out_875             ( col_out_875    ),
    .col_out_876             ( col_out_876    ),
    .col_out_877             ( col_out_877    ),
    .col_out_878             ( col_out_878    ),
    .col_out_879             ( col_out_879    ),
    .col_out_880             ( col_out_880    ),
    .col_out_881             ( col_out_881    ),
    .col_out_882             ( col_out_882    ),
    .col_out_883             ( col_out_883    ),
    .col_out_884             ( col_out_884    ),
    .col_out_885             ( col_out_885    ),
    .col_out_886             ( col_out_886    ),
    .col_out_887             ( col_out_887    ),
    .col_out_888             ( col_out_888    ),
    .col_out_889             ( col_out_889    ),
    .col_out_890             ( col_out_890    ),
    .col_out_891             ( col_out_891    ),
    .col_out_892             ( col_out_892    ),
    .col_out_893             ( col_out_893    ),
    .col_out_894             ( col_out_894    ),
    .col_out_895             ( col_out_895    ),
    .col_out_896             ( col_out_896    ),
    .col_out_897             ( col_out_897    ),
    .col_out_898             ( col_out_898    ),
    .col_out_899             ( col_out_899    ),
    .col_out_900             ( col_out_900    ),
    .col_out_901             ( col_out_901    ),
    .col_out_902             ( col_out_902    ),
    .col_out_903             ( col_out_903    ),
    .col_out_904             ( col_out_904    ),
    .col_out_905             ( col_out_905    ),
    .col_out_906             ( col_out_906    ),
    .col_out_907             ( col_out_907    ),
    .col_out_908             ( col_out_908    ),
    .col_out_909             ( col_out_909    ),
    .col_out_910             ( col_out_910    ),
    .col_out_911             ( col_out_911    ),
    .col_out_912             ( col_out_912    ),
    .col_out_913             ( col_out_913    ),
    .col_out_914             ( col_out_914    ),
    .col_out_915             ( col_out_915    ),
    .col_out_916             ( col_out_916    ),
    .col_out_917             ( col_out_917    ),
    .col_out_918             ( col_out_918    ),
    .col_out_919             ( col_out_919    ),
    .col_out_920             ( col_out_920    ),
    .col_out_921             ( col_out_921    ),
    .col_out_922             ( col_out_922    ),
    .col_out_923             ( col_out_923    ),
    .col_out_924             ( col_out_924    ),
    .col_out_925             ( col_out_925    ),
    .col_out_926             ( col_out_926    ),
    .col_out_927             ( col_out_927    ),
    .col_out_928             ( col_out_928    ),
    .col_out_929             ( col_out_929    ),
    .col_out_930             ( col_out_930    ),
    .col_out_931             ( col_out_931    ),
    .col_out_932             ( col_out_932    ),
    .col_out_933             ( col_out_933    ),
    .col_out_934             ( col_out_934    ),
    .col_out_935             ( col_out_935    ),
    .col_out_936             ( col_out_936    ),
    .col_out_937             ( col_out_937    ),
    .col_out_938             ( col_out_938    ),
    .col_out_939             ( col_out_939    ),
    .col_out_940             ( col_out_940    ),
    .col_out_941             ( col_out_941    ),
    .col_out_942             ( col_out_942    ),
    .col_out_943             ( col_out_943    ),
    .col_out_944             ( col_out_944    ),
    .col_out_945             ( col_out_945    ),
    .col_out_946             ( col_out_946    ),
    .col_out_947             ( col_out_947    ),
    .col_out_948             ( col_out_948    ),
    .col_out_949             ( col_out_949    ),
    .col_out_950             ( col_out_950    ),
    .col_out_951             ( col_out_951    ),
    .col_out_952             ( col_out_952    ),
    .col_out_953             ( col_out_953    ),
    .col_out_954             ( col_out_954    ),
    .col_out_955             ( col_out_955    ),
    .col_out_956             ( col_out_956    ),
    .col_out_957             ( col_out_957    ),
    .col_out_958             ( col_out_958    ),
    .col_out_959             ( col_out_959    ),
    .col_out_960             ( col_out_960    ),
    .col_out_961             ( col_out_961    ),
    .col_out_962             ( col_out_962    ),
    .col_out_963             ( col_out_963    ),
    .col_out_964             ( col_out_964    ),
    .col_out_965             ( col_out_965    ),
    .col_out_966             ( col_out_966    ),
    .col_out_967             ( col_out_967    ),
    .col_out_968             ( col_out_968    ),
    .col_out_969             ( col_out_969    ),
    .col_out_970             ( col_out_970    ),
    .col_out_971             ( col_out_971    ),
    .col_out_972             ( col_out_972    ),
    .col_out_973             ( col_out_973    ),
    .col_out_974             ( col_out_974    ),
    .col_out_975             ( col_out_975    ),
    .col_out_976             ( col_out_976    ),
    .col_out_977             ( col_out_977    ),
    .col_out_978             ( col_out_978    ),
    .col_out_979             ( col_out_979    ),
    .col_out_980             ( col_out_980    ),
    .col_out_981             ( col_out_981    ),
    .col_out_982             ( col_out_982    ),
    .col_out_983             ( col_out_983    ),
    .col_out_984             ( col_out_984    ),
    .col_out_985             ( col_out_985    ),
    .col_out_986             ( col_out_986    ),
    .col_out_987             ( col_out_987    ),
    .col_out_988             ( col_out_988    ),
    .col_out_989             ( col_out_989    ),
    .col_out_990             ( col_out_990    ),
    .col_out_991             ( col_out_991    ),
    .col_out_992             ( col_out_992    ),
    .col_out_993             ( col_out_993    ),
    .col_out_994             ( col_out_994    ),
    .col_out_995             ( col_out_995    ),
    .col_out_996             ( col_out_996    ),
    .col_out_997             ( col_out_997    ),
    .col_out_998             ( col_out_998    ),
    .col_out_999             ( col_out_999    ),
    .col_out_1000            ( col_out_1000   ),
    .col_out_1001            ( col_out_1001   ),
    .col_out_1002            ( col_out_1002   ),
    .col_out_1003            ( col_out_1003   ),
    .col_out_1004            ( col_out_1004   ),
    .col_out_1005            ( col_out_1005   ),
    .col_out_1006            ( col_out_1006   ),
    .col_out_1007            ( col_out_1007   ),
    .col_out_1008            ( col_out_1008   ),
    .col_out_1009            ( col_out_1009   ),
    .col_out_1010            ( col_out_1010   ),
    .col_out_1011            ( col_out_1011   ),
    .col_out_1012            ( col_out_1012   ),
    .col_out_1013            ( col_out_1013   ),
    .col_out_1014            ( col_out_1014   ),
    .col_out_1015            ( col_out_1015   ),
    .col_out_1016            ( col_out_1016   ),
    .col_out_1017            ( col_out_1017   ),
    .col_out_1018            ( col_out_1018   ),
    .col_out_1019            ( col_out_1019   ),
    .col_out_1020            ( col_out_1020   ),
    .col_out_1021            ( col_out_1021   ),
    .col_out_1022            ( col_out_1022   ),
    .col_out_1023            ( col_out_1023   ),
    .col_out_1024            ( col_out_1024   ),
    .col_out_1025            ( col_out_1025   ),
    .col_out_1026            ( col_out_1026   ),
    .col_out_1027            ( col_out_1027   ),
    .col_out_1028            ( col_out_1028   ),
    .col_out_1029            ( col_out_1029   ),
    .col_out_1030            ( col_out_1030   ),
    .col_out_1031            ( col_out_1031   ),
    .col_out_1032            ( col_out_1032   )
);
















//*****************************************************
//**************输出赋值******************************
//*****************************************************
assign row_out_0 = {col_out_1032[0], col_out_1031[0], col_out_1030[0], col_out_1029[0], col_out_1028[0], col_out_1027[0], col_out_1026[0], col_out_1025[0], col_out_1024[0], col_out_1023[0], col_out_1022[0], col_out_1021[0], col_out_1020[0], col_out_1019[0], col_out_1018[0], col_out_1017[0], col_out_1016[0], col_out_1015[0], col_out_1014[0], col_out_1013[0], col_out_1012[0], col_out_1011[0], col_out_1010[0], col_out_1009[0], col_out_1008[0], col_out_1007[0], col_out_1006[0], col_out_1005[0], col_out_1004[0], col_out_1003[0], col_out_1002[0], col_out_1001[0], col_out_1000[0], col_out_999[0], col_out_998[0], col_out_997[0], col_out_996[0], col_out_995[0], col_out_994[0], col_out_993[0], col_out_992[0], col_out_991[0], col_out_990[0], col_out_989[0], col_out_988[0], col_out_987[0], col_out_986[0], col_out_985[0], col_out_984[0], col_out_983[0], col_out_982[0], col_out_981[0], col_out_980[0], col_out_979[0], col_out_978[0], col_out_977[0], col_out_976[0], col_out_975[0], col_out_974[0], col_out_973[0], col_out_972[0], col_out_971[0], col_out_970[0], col_out_969[0], col_out_968[0], col_out_967[0], col_out_966[0], col_out_965[0], col_out_964[0], col_out_963[0], col_out_962[0], col_out_961[0], col_out_960[0], col_out_959[0], col_out_958[0], col_out_957[0], col_out_956[0], col_out_955[0], col_out_954[0], col_out_953[0], col_out_952[0], col_out_951[0], col_out_950[0], col_out_949[0], col_out_948[0], col_out_947[0], col_out_946[0], col_out_945[0], col_out_944[0], col_out_943[0], col_out_942[0], col_out_941[0], col_out_940[0], col_out_939[0], col_out_938[0], col_out_937[0], col_out_936[0], col_out_935[0], col_out_934[0], col_out_933[0], col_out_932[0], col_out_931[0], col_out_930[0], col_out_929[0], col_out_928[0], col_out_927[0], col_out_926[0], col_out_925[0], col_out_924[0], col_out_923[0], col_out_922[0], col_out_921[0], col_out_920[0], col_out_919[0], col_out_918[0], col_out_917[0], col_out_916[0], col_out_915[0], col_out_914[0], col_out_913[0], col_out_912[0], col_out_911[0], col_out_910[0], col_out_909[0], col_out_908[0], col_out_907[0], col_out_906[0], col_out_905[0], col_out_904[0], col_out_903[0], col_out_902[0], col_out_901[0], col_out_900[0], col_out_899[0], col_out_898[0], col_out_897[0], col_out_896[0], col_out_895[0], col_out_894[0], col_out_893[0], col_out_892[0], col_out_891[0], col_out_890[0], col_out_889[0], col_out_888[0], col_out_887[0], col_out_886[0], col_out_885[0], col_out_884[0], col_out_883[0], col_out_882[0], col_out_881[0], col_out_880[0], col_out_879[0], col_out_878[0], col_out_877[0], col_out_876[0], col_out_875[0], col_out_874[0], col_out_873[0], col_out_872[0], col_out_871[0], col_out_870[0], col_out_869[0], col_out_868[0], col_out_867[0], col_out_866[0], col_out_865[0], col_out_864[0], col_out_863[0], col_out_862[0], col_out_861[0], col_out_860[0], col_out_859[0], col_out_858[0], col_out_857[0], col_out_856[0], col_out_855[0], col_out_854[0], col_out_853[0], col_out_852[0], col_out_851[0], col_out_850[0], col_out_849[0], col_out_848[0], col_out_847[0], col_out_846[0], col_out_845[0], col_out_844[0], col_out_843[0], col_out_842[0], col_out_841[0], col_out_840[0], col_out_839[0], col_out_838[0], col_out_837[0], col_out_836[0], col_out_835[0], col_out_834[0], col_out_833[0], col_out_832[0], col_out_831[0], col_out_830[0], col_out_829[0], col_out_828[0], col_out_827[0], col_out_826[0], col_out_825[0], col_out_824[0], col_out_823[0], col_out_822[0], col_out_821[0], col_out_820[0], col_out_819[0], col_out_818[0], col_out_817[0], col_out_816[0], col_out_815[0], col_out_814[0], col_out_813[0], col_out_812[0], col_out_811[0], col_out_810[0], col_out_809[0], col_out_808[0], col_out_807[0], col_out_806[0], col_out_805[0], col_out_804[0], col_out_803[0], col_out_802[0], col_out_801[0], col_out_800[0], col_out_799[0], col_out_798[0], col_out_797[0], col_out_796[0], col_out_795[0], col_out_794[0], col_out_793[0], col_out_792[0], col_out_791[0], col_out_790[0], col_out_789[0], col_out_788[0], col_out_787[0], col_out_786[0], col_out_785[0], col_out_784[0], col_out_783[0], col_out_782[0], col_out_781[0], col_out_780[0], col_out_779[0], col_out_778[0], col_out_777[0], col_out_776[0], col_out_775[0], col_out_774[0], col_out_773[0], col_out_772[0], col_out_771[0], col_out_770[0], col_out_769[0], col_out_768[0], col_out_767[0], col_out_766[0], col_out_765[0], col_out_764[0], col_out_763[0], col_out_762[0], col_out_761[0], col_out_760[0], col_out_759[0], col_out_758[0], col_out_757[0], col_out_756[0], col_out_755[0], col_out_754[0], col_out_753[0], col_out_752[0], col_out_751[0], col_out_750[0], col_out_749[0], col_out_748[0], col_out_747[0], col_out_746[0], col_out_745[0], col_out_744[0], col_out_743[0], col_out_742[0], col_out_741[0], col_out_740[0], col_out_739[0], col_out_738[0], col_out_737[0], col_out_736[0], col_out_735[0], col_out_734[0], col_out_733[0], col_out_732[0], col_out_731[0], col_out_730[0], col_out_729[0], col_out_728[0], col_out_727[0], col_out_726[0], col_out_725[0], col_out_724[0], col_out_723[0], col_out_722[0], col_out_721[0], col_out_720[0], col_out_719[0], col_out_718[0], col_out_717[0], col_out_716[0], col_out_715[0], col_out_714[0], col_out_713[0], col_out_712[0], col_out_711[0], col_out_710[0], col_out_709[0], col_out_708[0], col_out_707[0], col_out_706[0], col_out_705[0], col_out_704[0], col_out_703[0], col_out_702[0], col_out_701[0], col_out_700[0], col_out_699[0], col_out_698[0], col_out_697[0], col_out_696[0], col_out_695[0], col_out_694[0], col_out_693[0], col_out_692[0], col_out_691[0], col_out_690[0], col_out_689[0], col_out_688[0], col_out_687[0], col_out_686[0], col_out_685[0], col_out_684[0], col_out_683[0], col_out_682[0], col_out_681[0], col_out_680[0], col_out_679[0], col_out_678[0], col_out_677[0], col_out_676[0], col_out_675[0], col_out_674[0], col_out_673[0], col_out_672[0], col_out_671[0], col_out_670[0], col_out_669[0], col_out_668[0], col_out_667[0], col_out_666[0], col_out_665[0], col_out_664[0], col_out_663[0], col_out_662[0], col_out_661[0], col_out_660[0], col_out_659[0], col_out_658[0], col_out_657[0], col_out_656[0], col_out_655[0], col_out_654[0], col_out_653[0], col_out_652[0], col_out_651[0], col_out_650[0], col_out_649[0], col_out_648[0], col_out_647[0], col_out_646[0], col_out_645[0], col_out_644[0], col_out_643[0], col_out_642[0], col_out_641[0], col_out_640[0], col_out_639[0], col_out_638[0], col_out_637[0], col_out_636[0], col_out_635[0], col_out_634[0], col_out_633[0], col_out_632[0], col_out_631[0], col_out_630[0], col_out_629[0], col_out_628[0], col_out_627[0], col_out_626[0], col_out_625[0], col_out_624[0], col_out_623[0], col_out_622[0], col_out_621[0], col_out_620[0], col_out_619[0], col_out_618[0], col_out_617[0], col_out_616[0], col_out_615[0], col_out_614[0], col_out_613[0], col_out_612[0], col_out_611[0], col_out_610[0], col_out_609[0], col_out_608[0], col_out_607[0], col_out_606[0], col_out_605[0], col_out_604[0], col_out_603[0], col_out_602[0], col_out_601[0], col_out_600[0], col_out_599[0], col_out_598[0], col_out_597[0], col_out_596[0], col_out_595[0], col_out_594[0], col_out_593[0], col_out_592[0], col_out_591[0], col_out_590[0], col_out_589[0], col_out_588[0], col_out_587[0], col_out_586[0], col_out_585[0], col_out_584[0], col_out_583[0], col_out_582[0], col_out_581[0], col_out_580[0], col_out_579[0], col_out_578[0], col_out_577[0], col_out_576[0], col_out_575[0], col_out_574[0], col_out_573[0], col_out_572[0], col_out_571[0], col_out_570[0], col_out_569[0], col_out_568[0], col_out_567[0], col_out_566[0], col_out_565[0], col_out_564[0], col_out_563[0], col_out_562[0], col_out_561[0], col_out_560[0], col_out_559[0], col_out_558[0], col_out_557[0], col_out_556[0], col_out_555[0], col_out_554[0], col_out_553[0], col_out_552[0], col_out_551[0], col_out_550[0], col_out_549[0], col_out_548[0], col_out_547[0], col_out_546[0], col_out_545[0], col_out_544[0], col_out_543[0], col_out_542[0], col_out_541[0], col_out_540[0], col_out_539[0], col_out_538[0], col_out_537[0], col_out_536[0], col_out_535[0], col_out_534[0], col_out_533[0], col_out_532[0], col_out_531[0], col_out_530[0], col_out_529[0], col_out_528[0], col_out_527[0], col_out_526[0], col_out_525[0], col_out_524[0], col_out_523[0], col_out_522[0], col_out_521[0], col_out_520[0], col_out_519[0], col_out_518[0], col_out_517[0], col_out_516[0], col_out_515[0], col_out_514[0], col_out_513[0], col_out_512[0], col_out_511[0], col_out_510[0], col_out_509[0], col_out_508[0], col_out_507[0], col_out_506[0], col_out_505[0], col_out_504[0], col_out_503[0], col_out_502[0], col_out_501[0], col_out_500[0], col_out_499[0], col_out_498[0], col_out_497[0], col_out_496[0], col_out_495[0], col_out_494[0], col_out_493[0], col_out_492[0], col_out_491[0], col_out_490[0], col_out_489[0], col_out_488[0], col_out_487[0], col_out_486[0], col_out_485[0], col_out_484[0], col_out_483[0], col_out_482[0], col_out_481[0], col_out_480[0], col_out_479[0], col_out_478[0], col_out_477[0], col_out_476[0], col_out_475[0], col_out_474[0], col_out_473[0], col_out_472[0], col_out_471[0], col_out_470[0], col_out_469[0], col_out_468[0], col_out_467[0], col_out_466[0], col_out_465[0], col_out_464[0], col_out_463[0], col_out_462[0], col_out_461[0], col_out_460[0], col_out_459[0], col_out_458[0], col_out_457[0], col_out_456[0], col_out_455[0], col_out_454[0], col_out_453[0], col_out_452[0], col_out_451[0], col_out_450[0], col_out_449[0], col_out_448[0], col_out_447[0], col_out_446[0], col_out_445[0], col_out_444[0], col_out_443[0], col_out_442[0], col_out_441[0], col_out_440[0], col_out_439[0], col_out_438[0], col_out_437[0], col_out_436[0], col_out_435[0], col_out_434[0], col_out_433[0], col_out_432[0], col_out_431[0], col_out_430[0], col_out_429[0], col_out_428[0], col_out_427[0], col_out_426[0], col_out_425[0], col_out_424[0], col_out_423[0], col_out_422[0], col_out_421[0], col_out_420[0], col_out_419[0], col_out_418[0], col_out_417[0], col_out_416[0], col_out_415[0], col_out_414[0], col_out_413[0], col_out_412[0], col_out_411[0], col_out_410[0], col_out_409[0], col_out_408[0], col_out_407[0], col_out_406[0], col_out_405[0], col_out_404[0], col_out_403[0], col_out_402[0], col_out_401[0], col_out_400[0], col_out_399[0], col_out_398[0], col_out_397[0], col_out_396[0], col_out_395[0], col_out_394[0], col_out_393[0], col_out_392[0], col_out_391[0], col_out_390[0], col_out_389[0], col_out_388[0], col_out_387[0], col_out_386[0], col_out_385[0], col_out_384[0], col_out_383[0], col_out_382[0], col_out_381[0], col_out_380[0], col_out_379[0], col_out_378[0], col_out_377[0], col_out_376[0], col_out_375[0], col_out_374[0], col_out_373[0], col_out_372[0], col_out_371[0], col_out_370[0], col_out_369[0], col_out_368[0], col_out_367[0], col_out_366[0], col_out_365[0], col_out_364[0], col_out_363[0], col_out_362[0], col_out_361[0], col_out_360[0], col_out_359[0], col_out_358[0], col_out_357[0], col_out_356[0], col_out_355[0], col_out_354[0], col_out_353[0], col_out_352[0], col_out_351[0], col_out_350[0], col_out_349[0], col_out_348[0], col_out_347[0], col_out_346[0], col_out_345[0], col_out_344[0], col_out_343[0], col_out_342[0], col_out_341[0], col_out_340[0], col_out_339[0], col_out_338[0], col_out_337[0], col_out_336[0], col_out_335[0], col_out_334[0], col_out_333[0], col_out_332[0], col_out_331[0], col_out_330[0], col_out_329[0], col_out_328[0], col_out_327[0], col_out_326[0], col_out_325[0], col_out_324[0], col_out_323[0], col_out_322[0], col_out_321[0], col_out_320[0], col_out_319[0], col_out_318[0], col_out_317[0], col_out_316[0], col_out_315[0], col_out_314[0], col_out_313[0], col_out_312[0], col_out_311[0], col_out_310[0], col_out_309[0], col_out_308[0], col_out_307[0], col_out_306[0], col_out_305[0], col_out_304[0], col_out_303[0], col_out_302[0], col_out_301[0], col_out_300[0], col_out_299[0], col_out_298[0], col_out_297[0], col_out_296[0], col_out_295[0], col_out_294[0], col_out_293[0], col_out_292[0], col_out_291[0], col_out_290[0], col_out_289[0], col_out_288[0], col_out_287[0], col_out_286[0], col_out_285[0], col_out_284[0], col_out_283[0], col_out_282[0], col_out_281[0], col_out_280[0], col_out_279[0], col_out_278[0], col_out_277[0], col_out_276[0], col_out_275[0], col_out_274[0], col_out_273[0], col_out_272[0], col_out_271[0], col_out_270[0], col_out_269[0], col_out_268[0], col_out_267[0], col_out_266[0], col_out_265[0], col_out_264[0], col_out_263[0], col_out_262[0], col_out_261[0], col_out_260[0], col_out_259[0], col_out_258[0], col_out_257[0], col_out_256[0], col_out_255[0], col_out_254[0], col_out_253[0], col_out_252[0], col_out_251[0], col_out_250[0], col_out_249[0], col_out_248[0], col_out_247[0], col_out_246[0], col_out_245[0], col_out_244[0], col_out_243[0], col_out_242[0], col_out_241[0], col_out_240[0], col_out_239[0], col_out_238[0], col_out_237[0], col_out_236[0], col_out_235[0], col_out_234[0], col_out_233[0], col_out_232[0], col_out_231[0], col_out_230[0], col_out_229[0], col_out_228[0], col_out_227[0], col_out_226[0], col_out_225[0], col_out_224[0], col_out_223[0], col_out_222[0], col_out_221[0], col_out_220[0], col_out_219[0], col_out_218[0], col_out_217[0], col_out_216[0], col_out_215[0], col_out_214[0], col_out_213[0], col_out_212[0], col_out_211[0], col_out_210[0], col_out_209[0], col_out_208[0], col_out_207[0], col_out_206[0], col_out_205[0], col_out_204[0], col_out_203[0], col_out_202[0], col_out_201[0], col_out_200[0], col_out_199[0], col_out_198[0], col_out_197[0], col_out_196[0], col_out_195[0], col_out_194[0], col_out_193[0], col_out_192[0], col_out_191[0], col_out_190[0], col_out_189[0], col_out_188[0], col_out_187[0], col_out_186[0], col_out_185[0], col_out_184[0], col_out_183[0], col_out_182[0], col_out_181[0], col_out_180[0], col_out_179[0], col_out_178[0], col_out_177[0], col_out_176[0], col_out_175[0], col_out_174[0], col_out_173[0], col_out_172[0], col_out_171[0], col_out_170[0], col_out_169[0], col_out_168[0], col_out_167[0], col_out_166[0], col_out_165[0], col_out_164[0], col_out_163[0], col_out_162[0], col_out_161[0], col_out_160[0], col_out_159[0], col_out_158[0], col_out_157[0], col_out_156[0], col_out_155[0], col_out_154[0], col_out_153[0], col_out_152[0], col_out_151[0], col_out_150[0], col_out_149[0], col_out_148[0], col_out_147[0], col_out_146[0], col_out_145[0], col_out_144[0], col_out_143[0], col_out_142[0], col_out_141[0], col_out_140[0], col_out_139[0], col_out_138[0], col_out_137[0], col_out_136[0], col_out_135[0], col_out_134[0], col_out_133[0], col_out_132[0], col_out_131[0], col_out_130[0], col_out_129[0], col_out_128[0], col_out_127[0], col_out_126[0], col_out_125[0], col_out_124[0], col_out_123[0], col_out_122[0], col_out_121[0], col_out_120[0], col_out_119[0], col_out_118[0], col_out_117[0], col_out_116[0], col_out_115[0], col_out_114[0], col_out_113[0], col_out_112[0], col_out_111[0], col_out_110[0], col_out_109[0], col_out_108[0], col_out_107[0], col_out_106[0], col_out_105[0], col_out_104[0], col_out_103[0], col_out_102[0], col_out_101[0], col_out_100[0], col_out_99[0], col_out_98[0], col_out_97[0], col_out_96[0], col_out_95[0], col_out_94[0], col_out_93[0], col_out_92[0], col_out_91[0], col_out_90[0], col_out_89[0], col_out_88[0], col_out_87[0], col_out_86[0], col_out_85[0], col_out_84[0], col_out_83[0], col_out_82[0], col_out_81[0], col_out_80[0], col_out_79[0], col_out_78[0], col_out_77[0], col_out_76[0], col_out_75[0], col_out_74[0], col_out_73[0], col_out_72[0], col_out_71[0], col_out_70[0], col_out_69[0], col_out_68[0], col_out_67[0], col_out_66[0], col_out_65[0], col_out_64[0], col_out_63[0], col_out_62[0], col_out_61[0], col_out_60[0], col_out_59[0], col_out_58[0], col_out_57[0], col_out_56[0], col_out_55[0], col_out_54[0], col_out_53[0], col_out_52[0], col_out_51[0], col_out_50[0], col_out_49[0], col_out_48[0], col_out_47[0], col_out_46[0], col_out_45[0], col_out_44[0], col_out_43[0], col_out_42[0], col_out_41[0], col_out_40[0], col_out_39[0], col_out_38[0], col_out_37[0], col_out_36[0], col_out_35[0], col_out_34[0], col_out_33[0], col_out_32[0], col_out_31[0], col_out_30[0], col_out_29[0], col_out_28[0], col_out_27[0], col_out_26[0], col_out_25[0], col_out_24[0], col_out_23[0], col_out_22[0], col_out_21[0], col_out_20[0], col_out_19[0], col_out_18[0], col_out_17[0], col_out_16[0], col_out_15[0], col_out_14[0], col_out_13[0], col_out_12[0], col_out_11[0], col_out_10[0], col_out_9[0], col_out_8[0], col_out_7[0], col_out_6[0], col_out_5[0], col_out_4[0], col_out_3[0], col_out_2[0], col_out_1[0], col_out_0[0]};


assign row_out_1 = {col_out_1032[1], col_out_1031[1], col_out_1030[1], col_out_1029[1], col_out_1028[1], col_out_1027[1], col_out_1026[1], col_out_1025[1], col_out_1024[1], col_out_1023[1], col_out_1022[1], col_out_1021[1], col_out_1020[1], col_out_1019[1], col_out_1018[1], col_out_1017[1], col_out_1016[1], col_out_1015[1], col_out_1014[1], col_out_1013[1], col_out_1012[1], col_out_1011[1], col_out_1010[1], col_out_1009[1], col_out_1008[1], col_out_1007[1], col_out_1006[1], col_out_1005[1], col_out_1004[1], col_out_1003[1], col_out_1002[1], col_out_1001[1], col_out_1000[1], col_out_999[1], col_out_998[1], col_out_997[1], col_out_996[1], col_out_995[1], col_out_994[1], col_out_993[1], col_out_992[1], col_out_991[1], col_out_990[1], col_out_989[1], col_out_988[1], col_out_987[1], col_out_986[1], col_out_985[1], col_out_984[1], col_out_983[1], col_out_982[1], col_out_981[1], col_out_980[1], col_out_979[1], col_out_978[1], col_out_977[1], col_out_976[1], col_out_975[1], col_out_974[1], col_out_973[1], col_out_972[1], col_out_971[1], col_out_970[1], col_out_969[1], col_out_968[1], col_out_967[1], col_out_966[1], col_out_965[1], col_out_964[1], col_out_963[1], col_out_962[1], col_out_961[1], col_out_960[1], col_out_959[1], col_out_958[1], col_out_957[1], col_out_956[1], col_out_955[1], col_out_954[1], col_out_953[1], col_out_952[1], col_out_951[1], col_out_950[1], col_out_949[1], col_out_948[1], col_out_947[1], col_out_946[1], col_out_945[1], col_out_944[1], col_out_943[1], col_out_942[1], col_out_941[1], col_out_940[1], col_out_939[1], col_out_938[1], col_out_937[1], col_out_936[1], col_out_935[1], col_out_934[1], col_out_933[1], col_out_932[1], col_out_931[1], col_out_930[1], col_out_929[1], col_out_928[1], col_out_927[1], col_out_926[1], col_out_925[1], col_out_924[1], col_out_923[1], col_out_922[1], col_out_921[1], col_out_920[1], col_out_919[1], col_out_918[1], col_out_917[1], col_out_916[1], col_out_915[1], col_out_914[1], col_out_913[1], col_out_912[1], col_out_911[1], col_out_910[1], col_out_909[1], col_out_908[1], col_out_907[1], col_out_906[1], col_out_905[1], col_out_904[1], col_out_903[1], col_out_902[1], col_out_901[1], col_out_900[1], col_out_899[1], col_out_898[1], col_out_897[1], col_out_896[1], col_out_895[1], col_out_894[1], col_out_893[1], col_out_892[1], col_out_891[1], col_out_890[1], col_out_889[1], col_out_888[1], col_out_887[1], col_out_886[1], col_out_885[1], col_out_884[1], col_out_883[1], col_out_882[1], col_out_881[1], col_out_880[1], col_out_879[1], col_out_878[1], col_out_877[1], col_out_876[1], col_out_875[1], col_out_874[1], col_out_873[1], col_out_872[1], col_out_871[1], col_out_870[1], col_out_869[1], col_out_868[1], col_out_867[1], col_out_866[1], col_out_865[1], col_out_864[1], col_out_863[1], col_out_862[1], col_out_861[1], col_out_860[1], col_out_859[1], col_out_858[1], col_out_857[1], col_out_856[1], col_out_855[1], col_out_854[1], col_out_853[1], col_out_852[1], col_out_851[1], col_out_850[1], col_out_849[1], col_out_848[1], col_out_847[1], col_out_846[1], col_out_845[1], col_out_844[1], col_out_843[1], col_out_842[1], col_out_841[1], col_out_840[1], col_out_839[1], col_out_838[1], col_out_837[1], col_out_836[1], col_out_835[1], col_out_834[1], col_out_833[1], col_out_832[1], col_out_831[1], col_out_830[1], col_out_829[1], col_out_828[1], col_out_827[1], col_out_826[1], col_out_825[1], col_out_824[1], col_out_823[1], col_out_822[1], col_out_821[1], col_out_820[1], col_out_819[1], col_out_818[1], col_out_817[1], col_out_816[1], col_out_815[1], col_out_814[1], col_out_813[1], col_out_812[1], col_out_811[1], col_out_810[1], col_out_809[1], col_out_808[1], col_out_807[1], col_out_806[1], col_out_805[1], col_out_804[1], col_out_803[1], col_out_802[1], col_out_801[1], col_out_800[1], col_out_799[1], col_out_798[1], col_out_797[1], col_out_796[1], col_out_795[1], col_out_794[1], col_out_793[1], col_out_792[1], col_out_791[1], col_out_790[1], col_out_789[1], col_out_788[1], col_out_787[1], col_out_786[1], col_out_785[1], col_out_784[1], col_out_783[1], col_out_782[1], col_out_781[1], col_out_780[1], col_out_779[1], col_out_778[1], col_out_777[1], col_out_776[1], col_out_775[1], col_out_774[1], col_out_773[1], col_out_772[1], col_out_771[1], col_out_770[1], col_out_769[1], col_out_768[1], col_out_767[1], col_out_766[1], col_out_765[1], col_out_764[1], col_out_763[1], col_out_762[1], col_out_761[1], col_out_760[1], col_out_759[1], col_out_758[1], col_out_757[1], col_out_756[1], col_out_755[1], col_out_754[1], col_out_753[1], col_out_752[1], col_out_751[1], col_out_750[1], col_out_749[1], col_out_748[1], col_out_747[1], col_out_746[1], col_out_745[1], col_out_744[1], col_out_743[1], col_out_742[1], col_out_741[1], col_out_740[1], col_out_739[1], col_out_738[1], col_out_737[1], col_out_736[1], col_out_735[1], col_out_734[1], col_out_733[1], col_out_732[1], col_out_731[1], col_out_730[1], col_out_729[1], col_out_728[1], col_out_727[1], col_out_726[1], col_out_725[1], col_out_724[1], col_out_723[1], col_out_722[1], col_out_721[1], col_out_720[1], col_out_719[1], col_out_718[1], col_out_717[1], col_out_716[1], col_out_715[1], col_out_714[1], col_out_713[1], col_out_712[1], col_out_711[1], col_out_710[1], col_out_709[1], col_out_708[1], col_out_707[1], col_out_706[1], col_out_705[1], col_out_704[1], col_out_703[1], col_out_702[1], col_out_701[1], col_out_700[1], col_out_699[1], col_out_698[1], col_out_697[1], col_out_696[1], col_out_695[1], col_out_694[1], col_out_693[1], col_out_692[1], col_out_691[1], col_out_690[1], col_out_689[1], col_out_688[1], col_out_687[1], col_out_686[1], col_out_685[1], col_out_684[1], col_out_683[1], col_out_682[1], col_out_681[1], col_out_680[1], col_out_679[1], col_out_678[1], col_out_677[1], col_out_676[1], col_out_675[1], col_out_674[1], col_out_673[1], col_out_672[1], col_out_671[1], col_out_670[1], col_out_669[1], col_out_668[1], col_out_667[1], col_out_666[1], col_out_665[1], col_out_664[1], col_out_663[1], col_out_662[1], col_out_661[1], col_out_660[1], col_out_659[1], col_out_658[1], col_out_657[1], col_out_656[1], col_out_655[1], col_out_654[1], col_out_653[1], col_out_652[1], col_out_651[1], col_out_650[1], col_out_649[1], col_out_648[1], col_out_647[1], col_out_646[1], col_out_645[1], col_out_644[1], col_out_643[1], col_out_642[1], col_out_641[1], col_out_640[1], col_out_639[1], col_out_638[1], col_out_637[1], col_out_636[1], col_out_635[1], col_out_634[1], col_out_633[1], col_out_632[1], col_out_631[1], col_out_630[1], col_out_629[1], col_out_628[1], col_out_627[1], col_out_626[1], col_out_625[1], col_out_624[1], col_out_623[1], col_out_622[1], col_out_621[1], col_out_620[1], col_out_619[1], col_out_618[1], col_out_617[1], col_out_616[1], col_out_615[1], col_out_614[1], col_out_613[1], col_out_612[1], col_out_611[1], col_out_610[1], col_out_609[1], col_out_608[1], col_out_607[1], col_out_606[1], col_out_605[1], col_out_604[1], col_out_603[1], col_out_602[1], col_out_601[1], col_out_600[1], col_out_599[1], col_out_598[1], col_out_597[1], col_out_596[1], col_out_595[1], col_out_594[1], col_out_593[1], col_out_592[1], col_out_591[1], col_out_590[1], col_out_589[1], col_out_588[1], col_out_587[1], col_out_586[1], col_out_585[1], col_out_584[1], col_out_583[1], col_out_582[1], col_out_581[1], col_out_580[1], col_out_579[1], col_out_578[1], col_out_577[1], col_out_576[1], col_out_575[1], col_out_574[1], col_out_573[1], col_out_572[1], col_out_571[1], col_out_570[1], col_out_569[1], col_out_568[1], col_out_567[1], col_out_566[1], col_out_565[1], col_out_564[1], col_out_563[1], col_out_562[1], col_out_561[1], col_out_560[1], col_out_559[1], col_out_558[1], col_out_557[1], col_out_556[1], col_out_555[1], col_out_554[1], col_out_553[1], col_out_552[1], col_out_551[1], col_out_550[1], col_out_549[1], col_out_548[1], col_out_547[1], col_out_546[1], col_out_545[1], col_out_544[1], col_out_543[1], col_out_542[1], col_out_541[1], col_out_540[1], col_out_539[1], col_out_538[1], col_out_537[1], col_out_536[1], col_out_535[1], col_out_534[1], col_out_533[1], col_out_532[1], col_out_531[1], col_out_530[1], col_out_529[1], col_out_528[1], col_out_527[1], col_out_526[1], col_out_525[1], col_out_524[1], col_out_523[1], col_out_522[1], col_out_521[1], col_out_520[1], col_out_519[1], col_out_518[1], col_out_517[1], col_out_516[1], col_out_515[1], col_out_514[1], col_out_513[1], col_out_512[1], col_out_511[1], col_out_510[1], col_out_509[1], col_out_508[1], col_out_507[1], col_out_506[1], col_out_505[1], col_out_504[1], col_out_503[1], col_out_502[1], col_out_501[1], col_out_500[1], col_out_499[1], col_out_498[1], col_out_497[1], col_out_496[1], col_out_495[1], col_out_494[1], col_out_493[1], col_out_492[1], col_out_491[1], col_out_490[1], col_out_489[1], col_out_488[1], col_out_487[1], col_out_486[1], col_out_485[1], col_out_484[1], col_out_483[1], col_out_482[1], col_out_481[1], col_out_480[1], col_out_479[1], col_out_478[1], col_out_477[1], col_out_476[1], col_out_475[1], col_out_474[1], col_out_473[1], col_out_472[1], col_out_471[1], col_out_470[1], col_out_469[1], col_out_468[1], col_out_467[1], col_out_466[1], col_out_465[1], col_out_464[1], col_out_463[1], col_out_462[1], col_out_461[1], col_out_460[1], col_out_459[1], col_out_458[1], col_out_457[1], col_out_456[1], col_out_455[1], col_out_454[1], col_out_453[1], col_out_452[1], col_out_451[1], col_out_450[1], col_out_449[1], col_out_448[1], col_out_447[1], col_out_446[1], col_out_445[1], col_out_444[1], col_out_443[1], col_out_442[1], col_out_441[1], col_out_440[1], col_out_439[1], col_out_438[1], col_out_437[1], col_out_436[1], col_out_435[1], col_out_434[1], col_out_433[1], col_out_432[1], col_out_431[1], col_out_430[1], col_out_429[1], col_out_428[1], col_out_427[1], col_out_426[1], col_out_425[1], col_out_424[1], col_out_423[1], col_out_422[1], col_out_421[1], col_out_420[1], col_out_419[1], col_out_418[1], col_out_417[1], col_out_416[1], col_out_415[1], col_out_414[1], col_out_413[1], col_out_412[1], col_out_411[1], col_out_410[1], col_out_409[1], col_out_408[1], col_out_407[1], col_out_406[1], col_out_405[1], col_out_404[1], col_out_403[1], col_out_402[1], col_out_401[1], col_out_400[1], col_out_399[1], col_out_398[1], col_out_397[1], col_out_396[1], col_out_395[1], col_out_394[1], col_out_393[1], col_out_392[1], col_out_391[1], col_out_390[1], col_out_389[1], col_out_388[1], col_out_387[1], col_out_386[1], col_out_385[1], col_out_384[1], col_out_383[1], col_out_382[1], col_out_381[1], col_out_380[1], col_out_379[1], col_out_378[1], col_out_377[1], col_out_376[1], col_out_375[1], col_out_374[1], col_out_373[1], col_out_372[1], col_out_371[1], col_out_370[1], col_out_369[1], col_out_368[1], col_out_367[1], col_out_366[1], col_out_365[1], col_out_364[1], col_out_363[1], col_out_362[1], col_out_361[1], col_out_360[1], col_out_359[1], col_out_358[1], col_out_357[1], col_out_356[1], col_out_355[1], col_out_354[1], col_out_353[1], col_out_352[1], col_out_351[1], col_out_350[1], col_out_349[1], col_out_348[1], col_out_347[1], col_out_346[1], col_out_345[1], col_out_344[1], col_out_343[1], col_out_342[1], col_out_341[1], col_out_340[1], col_out_339[1], col_out_338[1], col_out_337[1], col_out_336[1], col_out_335[1], col_out_334[1], col_out_333[1], col_out_332[1], col_out_331[1], col_out_330[1], col_out_329[1], col_out_328[1], col_out_327[1], col_out_326[1], col_out_325[1], col_out_324[1], col_out_323[1], col_out_322[1], col_out_321[1], col_out_320[1], col_out_319[1], col_out_318[1], col_out_317[1], col_out_316[1], col_out_315[1], col_out_314[1], col_out_313[1], col_out_312[1], col_out_311[1], col_out_310[1], col_out_309[1], col_out_308[1], col_out_307[1], col_out_306[1], col_out_305[1], col_out_304[1], col_out_303[1], col_out_302[1], col_out_301[1], col_out_300[1], col_out_299[1], col_out_298[1], col_out_297[1], col_out_296[1], col_out_295[1], col_out_294[1], col_out_293[1], col_out_292[1], col_out_291[1], col_out_290[1], col_out_289[1], col_out_288[1], col_out_287[1], col_out_286[1], col_out_285[1], col_out_284[1], col_out_283[1], col_out_282[1], col_out_281[1], col_out_280[1], col_out_279[1], col_out_278[1], col_out_277[1], col_out_276[1], col_out_275[1], col_out_274[1], col_out_273[1], col_out_272[1], col_out_271[1], col_out_270[1], col_out_269[1], col_out_268[1], col_out_267[1], col_out_266[1], col_out_265[1], col_out_264[1], col_out_263[1], col_out_262[1], col_out_261[1], col_out_260[1], col_out_259[1], col_out_258[1], col_out_257[1], col_out_256[1], col_out_255[1], col_out_254[1], col_out_253[1], col_out_252[1], col_out_251[1], col_out_250[1], col_out_249[1], col_out_248[1], col_out_247[1], col_out_246[1], col_out_245[1], col_out_244[1], col_out_243[1], col_out_242[1], col_out_241[1], col_out_240[1], col_out_239[1], col_out_238[1], col_out_237[1], col_out_236[1], col_out_235[1], col_out_234[1], col_out_233[1], col_out_232[1], col_out_231[1], col_out_230[1], col_out_229[1], col_out_228[1], col_out_227[1], col_out_226[1], col_out_225[1], col_out_224[1], col_out_223[1], col_out_222[1], col_out_221[1], col_out_220[1], col_out_219[1], col_out_218[1], col_out_217[1], col_out_216[1], col_out_215[1], col_out_214[1], col_out_213[1], col_out_212[1], col_out_211[1], col_out_210[1], col_out_209[1], col_out_208[1], col_out_207[1], col_out_206[1], col_out_205[1], col_out_204[1], col_out_203[1], col_out_202[1], col_out_201[1], col_out_200[1], col_out_199[1], col_out_198[1], col_out_197[1], col_out_196[1], col_out_195[1], col_out_194[1], col_out_193[1], col_out_192[1], col_out_191[1], col_out_190[1], col_out_189[1], col_out_188[1], col_out_187[1], col_out_186[1], col_out_185[1], col_out_184[1], col_out_183[1], col_out_182[1], col_out_181[1], col_out_180[1], col_out_179[1], col_out_178[1], col_out_177[1], col_out_176[1], col_out_175[1], col_out_174[1], col_out_173[1], col_out_172[1], col_out_171[1], col_out_170[1], col_out_169[1], col_out_168[1], col_out_167[1], col_out_166[1], col_out_165[1], col_out_164[1], col_out_163[1], col_out_162[1], col_out_161[1], col_out_160[1], col_out_159[1], col_out_158[1], col_out_157[1], col_out_156[1], col_out_155[1], col_out_154[1], col_out_153[1], col_out_152[1], col_out_151[1], col_out_150[1], col_out_149[1], col_out_148[1], col_out_147[1], col_out_146[1], col_out_145[1], col_out_144[1], col_out_143[1], col_out_142[1], col_out_141[1], col_out_140[1], col_out_139[1], col_out_138[1], col_out_137[1], col_out_136[1], col_out_135[1], col_out_134[1], col_out_133[1], col_out_132[1], col_out_131[1], col_out_130[1], col_out_129[1], col_out_128[1], col_out_127[1], col_out_126[1], col_out_125[1], col_out_124[1], col_out_123[1], col_out_122[1], col_out_121[1], col_out_120[1], col_out_119[1], col_out_118[1], col_out_117[1], col_out_116[1], col_out_115[1], col_out_114[1], col_out_113[1], col_out_112[1], col_out_111[1], col_out_110[1], col_out_109[1], col_out_108[1], col_out_107[1], col_out_106[1], col_out_105[1], col_out_104[1], col_out_103[1], col_out_102[1], col_out_101[1], col_out_100[1], col_out_99[1], col_out_98[1], col_out_97[1], col_out_96[1], col_out_95[1], col_out_94[1], col_out_93[1], col_out_92[1], col_out_91[1], col_out_90[1], col_out_89[1], col_out_88[1], col_out_87[1], col_out_86[1], col_out_85[1], col_out_84[1], col_out_83[1], col_out_82[1], col_out_81[1], col_out_80[1], col_out_79[1], col_out_78[1], col_out_77[1], col_out_76[1], col_out_75[1], col_out_74[1], col_out_73[1], col_out_72[1], col_out_71[1], col_out_70[1], col_out_69[1], col_out_68[1], col_out_67[1], col_out_66[1], col_out_65[1], col_out_64[1], col_out_63[1], col_out_62[1], col_out_61[1], col_out_60[1], col_out_59[1], col_out_58[1], col_out_57[1], col_out_56[1], col_out_55[1], col_out_54[1], col_out_53[1], col_out_52[1], col_out_51[1], col_out_50[1], col_out_49[1], col_out_48[1], col_out_47[1], col_out_46[1], col_out_45[1], col_out_44[1], col_out_43[1], col_out_42[1], col_out_41[1], col_out_40[1], col_out_39[1], col_out_38[1], col_out_37[1], col_out_36[1], col_out_35[1], col_out_34[1], col_out_33[1], col_out_32[1], col_out_31[1], col_out_30[1], col_out_29[1], col_out_28[1], col_out_27[1], col_out_26[1], col_out_25[1], col_out_24[1], col_out_23[1], col_out_22[1], col_out_21[1], col_out_20[1], col_out_19[1], col_out_18[1], col_out_17[1], col_out_16[1], col_out_15[1], col_out_14[1], col_out_13[1], col_out_12[1], col_out_11[1], col_out_10[1], col_out_9[1], col_out_8[1], col_out_7[1], col_out_6[1], col_out_5[1], col_out_4[1], col_out_3[1], col_out_2[1], col_out_1[1], col_out_0[1]};


//---------------------------------------------------------


endmodule
module data_in_mux
(
    input [1023:0] a,
    input sel_hp,

    input   [1023:0]  partial_product_high0,
    input   [1023:0]  partial_product_high1,
    input   [1032:0]  partial_product_low0,
    input   [1032:0]  partial_product_low1,

    input sel_data_in,

    output [511:0] col_out_0,
    output [511:0] col_out_1,
    output [511:0] col_out_2,
    output [511:0] col_out_3,
    output [511:0] col_out_4,
    output [511:0] col_out_5,
    output [511:0] col_out_6,
    output [511:0] col_out_7,
    output [511:0] col_out_8,
    output [511:0] col_out_9,
    output [511:0] col_out_10,
    output [511:0] col_out_11,
    output [511:0] col_out_12,
    output [511:0] col_out_13,
    output [511:0] col_out_14,
    output [511:0] col_out_15,
    output [511:0] col_out_16,
    output [511:0] col_out_17,
    output [511:0] col_out_18,
    output [511:0] col_out_19,
    output [511:0] col_out_20,
    output [511:0] col_out_21,
    output [511:0] col_out_22,
    output [511:0] col_out_23,
    output [511:0] col_out_24,
    output [511:0] col_out_25,
    output [511:0] col_out_26,
    output [511:0] col_out_27,
    output [511:0] col_out_28,
    output [511:0] col_out_29,
    output [511:0] col_out_30,
    output [511:0] col_out_31,
    output [511:0] col_out_32,
    output [511:0] col_out_33,
    output [511:0] col_out_34,
    output [511:0] col_out_35,
    output [511:0] col_out_36,
    output [511:0] col_out_37,
    output [511:0] col_out_38,
    output [511:0] col_out_39,
    output [511:0] col_out_40,
    output [511:0] col_out_41,
    output [511:0] col_out_42,
    output [511:0] col_out_43,
    output [511:0] col_out_44,
    output [511:0] col_out_45,
    output [511:0] col_out_46,
    output [511:0] col_out_47,
    output [511:0] col_out_48,
    output [511:0] col_out_49,
    output [511:0] col_out_50,
    output [511:0] col_out_51,
    output [511:0] col_out_52,
    output [511:0] col_out_53,
    output [511:0] col_out_54,
    output [511:0] col_out_55,
    output [511:0] col_out_56,
    output [511:0] col_out_57,
    output [511:0] col_out_58,
    output [511:0] col_out_59,
    output [511:0] col_out_60,
    output [511:0] col_out_61,
    output [511:0] col_out_62,
    output [511:0] col_out_63,
    output [511:0] col_out_64,
    output [511:0] col_out_65,
    output [511:0] col_out_66,
    output [511:0] col_out_67,
    output [511:0] col_out_68,
    output [511:0] col_out_69,
    output [511:0] col_out_70,
    output [511:0] col_out_71,
    output [511:0] col_out_72,
    output [511:0] col_out_73,
    output [511:0] col_out_74,
    output [511:0] col_out_75,
    output [511:0] col_out_76,
    output [511:0] col_out_77,
    output [511:0] col_out_78,
    output [511:0] col_out_79,
    output [511:0] col_out_80,
    output [511:0] col_out_81,
    output [511:0] col_out_82,
    output [511:0] col_out_83,
    output [511:0] col_out_84,
    output [511:0] col_out_85,
    output [511:0] col_out_86,
    output [511:0] col_out_87,
    output [511:0] col_out_88,
    output [511:0] col_out_89,
    output [511:0] col_out_90,
    output [511:0] col_out_91,
    output [511:0] col_out_92,
    output [511:0] col_out_93,
    output [511:0] col_out_94,
    output [511:0] col_out_95,
    output [511:0] col_out_96,
    output [511:0] col_out_97,
    output [511:0] col_out_98,
    output [511:0] col_out_99,
    output [511:0] col_out_100,
    output [511:0] col_out_101,
    output [511:0] col_out_102,
    output [511:0] col_out_103,
    output [511:0] col_out_104,
    output [511:0] col_out_105,
    output [511:0] col_out_106,
    output [511:0] col_out_107,
    output [511:0] col_out_108,
    output [511:0] col_out_109,
    output [511:0] col_out_110,
    output [511:0] col_out_111,
    output [511:0] col_out_112,
    output [511:0] col_out_113,
    output [511:0] col_out_114,
    output [511:0] col_out_115,
    output [511:0] col_out_116,
    output [511:0] col_out_117,
    output [511:0] col_out_118,
    output [511:0] col_out_119,
    output [511:0] col_out_120,
    output [511:0] col_out_121,
    output [511:0] col_out_122,
    output [511:0] col_out_123,
    output [511:0] col_out_124,
    output [511:0] col_out_125,
    output [511:0] col_out_126,
    output [511:0] col_out_127,
    output [511:0] col_out_128,
    output [511:0] col_out_129,
    output [511:0] col_out_130,
    output [511:0] col_out_131,
    output [511:0] col_out_132,
    output [511:0] col_out_133,
    output [511:0] col_out_134,
    output [511:0] col_out_135,
    output [511:0] col_out_136,
    output [511:0] col_out_137,
    output [511:0] col_out_138,
    output [511:0] col_out_139,
    output [511:0] col_out_140,
    output [511:0] col_out_141,
    output [511:0] col_out_142,
    output [511:0] col_out_143,
    output [511:0] col_out_144,
    output [511:0] col_out_145,
    output [511:0] col_out_146,
    output [511:0] col_out_147,
    output [511:0] col_out_148,
    output [511:0] col_out_149,
    output [511:0] col_out_150,
    output [511:0] col_out_151,
    output [511:0] col_out_152,
    output [511:0] col_out_153,
    output [511:0] col_out_154,
    output [511:0] col_out_155,
    output [511:0] col_out_156,
    output [511:0] col_out_157,
    output [511:0] col_out_158,
    output [511:0] col_out_159,
    output [511:0] col_out_160,
    output [511:0] col_out_161,
    output [511:0] col_out_162,
    output [511:0] col_out_163,
    output [511:0] col_out_164,
    output [511:0] col_out_165,
    output [511:0] col_out_166,
    output [511:0] col_out_167,
    output [511:0] col_out_168,
    output [511:0] col_out_169,
    output [511:0] col_out_170,
    output [511:0] col_out_171,
    output [511:0] col_out_172,
    output [511:0] col_out_173,
    output [511:0] col_out_174,
    output [511:0] col_out_175,
    output [511:0] col_out_176,
    output [511:0] col_out_177,
    output [511:0] col_out_178,
    output [511:0] col_out_179,
    output [511:0] col_out_180,
    output [511:0] col_out_181,
    output [511:0] col_out_182,
    output [511:0] col_out_183,
    output [511:0] col_out_184,
    output [511:0] col_out_185,
    output [511:0] col_out_186,
    output [511:0] col_out_187,
    output [511:0] col_out_188,
    output [511:0] col_out_189,
    output [511:0] col_out_190,
    output [511:0] col_out_191,
    output [511:0] col_out_192,
    output [511:0] col_out_193,
    output [511:0] col_out_194,
    output [511:0] col_out_195,
    output [511:0] col_out_196,
    output [511:0] col_out_197,
    output [511:0] col_out_198,
    output [511:0] col_out_199,
    output [511:0] col_out_200,
    output [511:0] col_out_201,
    output [511:0] col_out_202,
    output [511:0] col_out_203,
    output [511:0] col_out_204,
    output [511:0] col_out_205,
    output [511:0] col_out_206,
    output [511:0] col_out_207,
    output [511:0] col_out_208,
    output [511:0] col_out_209,
    output [511:0] col_out_210,
    output [511:0] col_out_211,
    output [511:0] col_out_212,
    output [511:0] col_out_213,
    output [511:0] col_out_214,
    output [511:0] col_out_215,
    output [511:0] col_out_216,
    output [511:0] col_out_217,
    output [511:0] col_out_218,
    output [511:0] col_out_219,
    output [511:0] col_out_220,
    output [511:0] col_out_221,
    output [511:0] col_out_222,
    output [511:0] col_out_223,
    output [511:0] col_out_224,
    output [511:0] col_out_225,
    output [511:0] col_out_226,
    output [511:0] col_out_227,
    output [511:0] col_out_228,
    output [511:0] col_out_229,
    output [511:0] col_out_230,
    output [511:0] col_out_231,
    output [511:0] col_out_232,
    output [511:0] col_out_233,
    output [511:0] col_out_234,
    output [511:0] col_out_235,
    output [511:0] col_out_236,
    output [511:0] col_out_237,
    output [511:0] col_out_238,
    output [511:0] col_out_239,
    output [511:0] col_out_240,
    output [511:0] col_out_241,
    output [511:0] col_out_242,
    output [511:0] col_out_243,
    output [511:0] col_out_244,
    output [511:0] col_out_245,
    output [511:0] col_out_246,
    output [511:0] col_out_247,
    output [511:0] col_out_248,
    output [511:0] col_out_249,
    output [511:0] col_out_250,
    output [511:0] col_out_251,
    output [511:0] col_out_252,
    output [511:0] col_out_253,
    output [511:0] col_out_254,
    output [511:0] col_out_255,
    output [511:0] col_out_256,
    output [511:0] col_out_257,
    output [511:0] col_out_258,
    output [511:0] col_out_259,
    output [511:0] col_out_260,
    output [511:0] col_out_261,
    output [511:0] col_out_262,
    output [511:0] col_out_263,
    output [511:0] col_out_264,
    output [511:0] col_out_265,
    output [511:0] col_out_266,
    output [511:0] col_out_267,
    output [511:0] col_out_268,
    output [511:0] col_out_269,
    output [511:0] col_out_270,
    output [511:0] col_out_271,
    output [511:0] col_out_272,
    output [511:0] col_out_273,
    output [511:0] col_out_274,
    output [511:0] col_out_275,
    output [511:0] col_out_276,
    output [511:0] col_out_277,
    output [511:0] col_out_278,
    output [511:0] col_out_279,
    output [511:0] col_out_280,
    output [511:0] col_out_281,
    output [511:0] col_out_282,
    output [511:0] col_out_283,
    output [511:0] col_out_284,
    output [511:0] col_out_285,
    output [511:0] col_out_286,
    output [511:0] col_out_287,
    output [511:0] col_out_288,
    output [511:0] col_out_289,
    output [511:0] col_out_290,
    output [511:0] col_out_291,
    output [511:0] col_out_292,
    output [511:0] col_out_293,
    output [511:0] col_out_294,
    output [511:0] col_out_295,
    output [511:0] col_out_296,
    output [511:0] col_out_297,
    output [511:0] col_out_298,
    output [511:0] col_out_299,
    output [511:0] col_out_300,
    output [511:0] col_out_301,
    output [511:0] col_out_302,
    output [511:0] col_out_303,
    output [511:0] col_out_304,
    output [511:0] col_out_305,
    output [511:0] col_out_306,
    output [511:0] col_out_307,
    output [511:0] col_out_308,
    output [511:0] col_out_309,
    output [511:0] col_out_310,
    output [511:0] col_out_311,
    output [511:0] col_out_312,
    output [511:0] col_out_313,
    output [511:0] col_out_314,
    output [511:0] col_out_315,
    output [511:0] col_out_316,
    output [511:0] col_out_317,
    output [511:0] col_out_318,
    output [511:0] col_out_319,
    output [511:0] col_out_320,
    output [511:0] col_out_321,
    output [511:0] col_out_322,
    output [511:0] col_out_323,
    output [511:0] col_out_324,
    output [511:0] col_out_325,
    output [511:0] col_out_326,
    output [511:0] col_out_327,
    output [511:0] col_out_328,
    output [511:0] col_out_329,
    output [511:0] col_out_330,
    output [511:0] col_out_331,
    output [511:0] col_out_332,
    output [511:0] col_out_333,
    output [511:0] col_out_334,
    output [511:0] col_out_335,
    output [511:0] col_out_336,
    output [511:0] col_out_337,
    output [511:0] col_out_338,
    output [511:0] col_out_339,
    output [511:0] col_out_340,
    output [511:0] col_out_341,
    output [511:0] col_out_342,
    output [511:0] col_out_343,
    output [511:0] col_out_344,
    output [511:0] col_out_345,
    output [511:0] col_out_346,
    output [511:0] col_out_347,
    output [511:0] col_out_348,
    output [511:0] col_out_349,
    output [511:0] col_out_350,
    output [511:0] col_out_351,
    output [511:0] col_out_352,
    output [511:0] col_out_353,
    output [511:0] col_out_354,
    output [511:0] col_out_355,
    output [511:0] col_out_356,
    output [511:0] col_out_357,
    output [511:0] col_out_358,
    output [511:0] col_out_359,
    output [511:0] col_out_360,
    output [511:0] col_out_361,
    output [511:0] col_out_362,
    output [511:0] col_out_363,
    output [511:0] col_out_364,
    output [511:0] col_out_365,
    output [511:0] col_out_366,
    output [511:0] col_out_367,
    output [511:0] col_out_368,
    output [511:0] col_out_369,
    output [511:0] col_out_370,
    output [511:0] col_out_371,
    output [511:0] col_out_372,
    output [511:0] col_out_373,
    output [511:0] col_out_374,
    output [511:0] col_out_375,
    output [511:0] col_out_376,
    output [511:0] col_out_377,
    output [511:0] col_out_378,
    output [511:0] col_out_379,
    output [511:0] col_out_380,
    output [511:0] col_out_381,
    output [511:0] col_out_382,
    output [511:0] col_out_383,
    output [511:0] col_out_384,
    output [511:0] col_out_385,
    output [511:0] col_out_386,
    output [511:0] col_out_387,
    output [511:0] col_out_388,
    output [511:0] col_out_389,
    output [511:0] col_out_390,
    output [511:0] col_out_391,
    output [511:0] col_out_392,
    output [511:0] col_out_393,
    output [511:0] col_out_394,
    output [511:0] col_out_395,
    output [511:0] col_out_396,
    output [511:0] col_out_397,
    output [511:0] col_out_398,
    output [511:0] col_out_399,
    output [511:0] col_out_400,
    output [511:0] col_out_401,
    output [511:0] col_out_402,
    output [511:0] col_out_403,
    output [511:0] col_out_404,
    output [511:0] col_out_405,
    output [511:0] col_out_406,
    output [511:0] col_out_407,
    output [511:0] col_out_408,
    output [511:0] col_out_409,
    output [511:0] col_out_410,
    output [511:0] col_out_411,
    output [511:0] col_out_412,
    output [511:0] col_out_413,
    output [511:0] col_out_414,
    output [511:0] col_out_415,
    output [511:0] col_out_416,
    output [511:0] col_out_417,
    output [511:0] col_out_418,
    output [511:0] col_out_419,
    output [511:0] col_out_420,
    output [511:0] col_out_421,
    output [511:0] col_out_422,
    output [511:0] col_out_423,
    output [511:0] col_out_424,
    output [511:0] col_out_425,
    output [511:0] col_out_426,
    output [511:0] col_out_427,
    output [511:0] col_out_428,
    output [511:0] col_out_429,
    output [511:0] col_out_430,
    output [511:0] col_out_431,
    output [511:0] col_out_432,
    output [511:0] col_out_433,
    output [511:0] col_out_434,
    output [511:0] col_out_435,
    output [511:0] col_out_436,
    output [511:0] col_out_437,
    output [511:0] col_out_438,
    output [511:0] col_out_439,
    output [511:0] col_out_440,
    output [511:0] col_out_441,
    output [511:0] col_out_442,
    output [511:0] col_out_443,
    output [511:0] col_out_444,
    output [511:0] col_out_445,
    output [511:0] col_out_446,
    output [511:0] col_out_447,
    output [511:0] col_out_448,
    output [511:0] col_out_449,
    output [511:0] col_out_450,
    output [511:0] col_out_451,
    output [511:0] col_out_452,
    output [511:0] col_out_453,
    output [511:0] col_out_454,
    output [511:0] col_out_455,
    output [511:0] col_out_456,
    output [511:0] col_out_457,
    output [511:0] col_out_458,
    output [511:0] col_out_459,
    output [511:0] col_out_460,
    output [511:0] col_out_461,
    output [511:0] col_out_462,
    output [511:0] col_out_463,
    output [511:0] col_out_464,
    output [511:0] col_out_465,
    output [511:0] col_out_466,
    output [511:0] col_out_467,
    output [511:0] col_out_468,
    output [511:0] col_out_469,
    output [511:0] col_out_470,
    output [511:0] col_out_471,
    output [511:0] col_out_472,
    output [511:0] col_out_473,
    output [511:0] col_out_474,
    output [511:0] col_out_475,
    output [511:0] col_out_476,
    output [511:0] col_out_477,
    output [511:0] col_out_478,
    output [511:0] col_out_479,
    output [511:0] col_out_480,
    output [511:0] col_out_481,
    output [511:0] col_out_482,
    output [511:0] col_out_483,
    output [511:0] col_out_484,
    output [511:0] col_out_485,
    output [511:0] col_out_486,
    output [511:0] col_out_487,
    output [511:0] col_out_488,
    output [511:0] col_out_489,
    output [511:0] col_out_490,
    output [511:0] col_out_491,
    output [511:0] col_out_492,
    output [511:0] col_out_493,
    output [511:0] col_out_494,
    output [511:0] col_out_495,
    output [511:0] col_out_496,
    output [511:0] col_out_497,
    output [511:0] col_out_498,
    output [511:0] col_out_499,
    output [511:0] col_out_500,
    output [511:0] col_out_501,
    output [511:0] col_out_502,
    output [511:0] col_out_503,
    output [511:0] col_out_504,
    output [511:0] col_out_505,
    output [511:0] col_out_506,
    output [511:0] col_out_507,
    output [511:0] col_out_508,
    output [511:0] col_out_509,
    output [511:0] col_out_510,
    output [511:0] col_out_511,
    output [511:0] col_out_512,
    output [511:0] col_out_513,
    output [511:0] col_out_514,
    output [511:0] col_out_515,
    output [511:0] col_out_516,
    output [511:0] col_out_517,
    output [511:0] col_out_518,
    output [511:0] col_out_519,
    output [511:0] col_out_520,
    output [511:0] col_out_521,
    output [511:0] col_out_522,
    output [511:0] col_out_523,
    output [511:0] col_out_524,
    output [511:0] col_out_525,
    output [511:0] col_out_526,
    output [511:0] col_out_527,
    output [511:0] col_out_528,
    output [511:0] col_out_529,
    output [511:0] col_out_530,
    output [511:0] col_out_531,
    output [511:0] col_out_532,
    output [511:0] col_out_533,
    output [511:0] col_out_534,
    output [511:0] col_out_535,
    output [511:0] col_out_536,
    output [511:0] col_out_537,
    output [511:0] col_out_538,
    output [511:0] col_out_539,
    output [511:0] col_out_540,
    output [511:0] col_out_541,
    output [511:0] col_out_542,
    output [511:0] col_out_543,
    output [511:0] col_out_544,
    output [511:0] col_out_545,
    output [511:0] col_out_546,
    output [511:0] col_out_547,
    output [511:0] col_out_548,
    output [511:0] col_out_549,
    output [511:0] col_out_550,
    output [511:0] col_out_551,
    output [511:0] col_out_552,
    output [511:0] col_out_553,
    output [511:0] col_out_554,
    output [511:0] col_out_555,
    output [511:0] col_out_556,
    output [511:0] col_out_557,
    output [511:0] col_out_558,
    output [511:0] col_out_559,
    output [511:0] col_out_560,
    output [511:0] col_out_561,
    output [511:0] col_out_562,
    output [511:0] col_out_563,
    output [511:0] col_out_564,
    output [511:0] col_out_565,
    output [511:0] col_out_566,
    output [511:0] col_out_567,
    output [511:0] col_out_568,
    output [511:0] col_out_569,
    output [511:0] col_out_570,
    output [511:0] col_out_571,
    output [511:0] col_out_572,
    output [511:0] col_out_573,
    output [511:0] col_out_574,
    output [511:0] col_out_575,
    output [511:0] col_out_576,
    output [511:0] col_out_577,
    output [511:0] col_out_578,
    output [511:0] col_out_579,
    output [511:0] col_out_580,
    output [511:0] col_out_581,
    output [511:0] col_out_582,
    output [511:0] col_out_583,
    output [511:0] col_out_584,
    output [511:0] col_out_585,
    output [511:0] col_out_586,
    output [511:0] col_out_587,
    output [511:0] col_out_588,
    output [511:0] col_out_589,
    output [511:0] col_out_590,
    output [511:0] col_out_591,
    output [511:0] col_out_592,
    output [511:0] col_out_593,
    output [511:0] col_out_594,
    output [511:0] col_out_595,
    output [511:0] col_out_596,
    output [511:0] col_out_597,
    output [511:0] col_out_598,
    output [511:0] col_out_599,
    output [511:0] col_out_600,
    output [511:0] col_out_601,
    output [511:0] col_out_602,
    output [511:0] col_out_603,
    output [511:0] col_out_604,
    output [511:0] col_out_605,
    output [511:0] col_out_606,
    output [511:0] col_out_607,
    output [511:0] col_out_608,
    output [511:0] col_out_609,
    output [511:0] col_out_610,
    output [511:0] col_out_611,
    output [511:0] col_out_612,
    output [511:0] col_out_613,
    output [511:0] col_out_614,
    output [511:0] col_out_615,
    output [511:0] col_out_616,
    output [511:0] col_out_617,
    output [511:0] col_out_618,
    output [511:0] col_out_619,
    output [511:0] col_out_620,
    output [511:0] col_out_621,
    output [511:0] col_out_622,
    output [511:0] col_out_623,
    output [511:0] col_out_624,
    output [511:0] col_out_625,
    output [511:0] col_out_626,
    output [511:0] col_out_627,
    output [511:0] col_out_628,
    output [511:0] col_out_629,
    output [511:0] col_out_630,
    output [511:0] col_out_631,
    output [511:0] col_out_632,
    output [511:0] col_out_633,
    output [511:0] col_out_634,
    output [511:0] col_out_635,
    output [511:0] col_out_636,
    output [511:0] col_out_637,
    output [511:0] col_out_638,
    output [511:0] col_out_639,
    output [511:0] col_out_640,
    output [511:0] col_out_641,
    output [511:0] col_out_642,
    output [511:0] col_out_643,
    output [511:0] col_out_644,
    output [511:0] col_out_645,
    output [511:0] col_out_646,
    output [511:0] col_out_647,
    output [511:0] col_out_648,
    output [511:0] col_out_649,
    output [511:0] col_out_650,
    output [511:0] col_out_651,
    output [511:0] col_out_652,
    output [511:0] col_out_653,
    output [511:0] col_out_654,
    output [511:0] col_out_655,
    output [511:0] col_out_656,
    output [511:0] col_out_657,
    output [511:0] col_out_658,
    output [511:0] col_out_659,
    output [511:0] col_out_660,
    output [511:0] col_out_661,
    output [511:0] col_out_662,
    output [511:0] col_out_663,
    output [511:0] col_out_664,
    output [511:0] col_out_665,
    output [511:0] col_out_666,
    output [511:0] col_out_667,
    output [511:0] col_out_668,
    output [511:0] col_out_669,
    output [511:0] col_out_670,
    output [511:0] col_out_671,
    output [511:0] col_out_672,
    output [511:0] col_out_673,
    output [511:0] col_out_674,
    output [511:0] col_out_675,
    output [511:0] col_out_676,
    output [511:0] col_out_677,
    output [511:0] col_out_678,
    output [511:0] col_out_679,
    output [511:0] col_out_680,
    output [511:0] col_out_681,
    output [511:0] col_out_682,
    output [511:0] col_out_683,
    output [511:0] col_out_684,
    output [511:0] col_out_685,
    output [511:0] col_out_686,
    output [511:0] col_out_687,
    output [511:0] col_out_688,
    output [511:0] col_out_689,
    output [511:0] col_out_690,
    output [511:0] col_out_691,
    output [511:0] col_out_692,
    output [511:0] col_out_693,
    output [511:0] col_out_694,
    output [511:0] col_out_695,
    output [511:0] col_out_696,
    output [511:0] col_out_697,
    output [511:0] col_out_698,
    output [511:0] col_out_699,
    output [511:0] col_out_700,
    output [511:0] col_out_701,
    output [511:0] col_out_702,
    output [511:0] col_out_703,
    output [511:0] col_out_704,
    output [511:0] col_out_705,
    output [511:0] col_out_706,
    output [511:0] col_out_707,
    output [511:0] col_out_708,
    output [511:0] col_out_709,
    output [511:0] col_out_710,
    output [511:0] col_out_711,
    output [511:0] col_out_712,
    output [511:0] col_out_713,
    output [511:0] col_out_714,
    output [511:0] col_out_715,
    output [511:0] col_out_716,
    output [511:0] col_out_717,
    output [511:0] col_out_718,
    output [511:0] col_out_719,
    output [511:0] col_out_720,
    output [511:0] col_out_721,
    output [511:0] col_out_722,
    output [511:0] col_out_723,
    output [511:0] col_out_724,
    output [511:0] col_out_725,
    output [511:0] col_out_726,
    output [511:0] col_out_727,
    output [511:0] col_out_728,
    output [511:0] col_out_729,
    output [511:0] col_out_730,
    output [511:0] col_out_731,
    output [511:0] col_out_732,
    output [511:0] col_out_733,
    output [511:0] col_out_734,
    output [511:0] col_out_735,
    output [511:0] col_out_736,
    output [511:0] col_out_737,
    output [511:0] col_out_738,
    output [511:0] col_out_739,
    output [511:0] col_out_740,
    output [511:0] col_out_741,
    output [511:0] col_out_742,
    output [511:0] col_out_743,
    output [511:0] col_out_744,
    output [511:0] col_out_745,
    output [511:0] col_out_746,
    output [511:0] col_out_747,
    output [511:0] col_out_748,
    output [511:0] col_out_749,
    output [511:0] col_out_750,
    output [511:0] col_out_751,
    output [511:0] col_out_752,
    output [511:0] col_out_753,
    output [511:0] col_out_754,
    output [511:0] col_out_755,
    output [511:0] col_out_756,
    output [511:0] col_out_757,
    output [511:0] col_out_758,
    output [511:0] col_out_759,
    output [511:0] col_out_760,
    output [511:0] col_out_761,
    output [511:0] col_out_762,
    output [511:0] col_out_763,
    output [511:0] col_out_764,
    output [511:0] col_out_765,
    output [511:0] col_out_766,
    output [511:0] col_out_767,
    output [511:0] col_out_768,
    output [511:0] col_out_769,
    output [511:0] col_out_770,
    output [511:0] col_out_771,
    output [511:0] col_out_772,
    output [511:0] col_out_773,
    output [511:0] col_out_774,
    output [511:0] col_out_775,
    output [511:0] col_out_776,
    output [511:0] col_out_777,
    output [511:0] col_out_778,
    output [511:0] col_out_779,
    output [511:0] col_out_780,
    output [511:0] col_out_781,
    output [511:0] col_out_782,
    output [511:0] col_out_783,
    output [511:0] col_out_784,
    output [511:0] col_out_785,
    output [511:0] col_out_786,
    output [511:0] col_out_787,
    output [511:0] col_out_788,
    output [511:0] col_out_789,
    output [511:0] col_out_790,
    output [511:0] col_out_791,
    output [511:0] col_out_792,
    output [511:0] col_out_793,
    output [511:0] col_out_794,
    output [511:0] col_out_795,
    output [511:0] col_out_796,
    output [511:0] col_out_797,
    output [511:0] col_out_798,
    output [511:0] col_out_799,
    output [511:0] col_out_800,
    output [511:0] col_out_801,
    output [511:0] col_out_802,
    output [511:0] col_out_803,
    output [511:0] col_out_804,
    output [511:0] col_out_805,
    output [511:0] col_out_806,
    output [511:0] col_out_807,
    output [511:0] col_out_808,
    output [511:0] col_out_809,
    output [511:0] col_out_810,
    output [511:0] col_out_811,
    output [511:0] col_out_812,
    output [511:0] col_out_813,
    output [511:0] col_out_814,
    output [511:0] col_out_815,
    output [511:0] col_out_816,
    output [511:0] col_out_817,
    output [511:0] col_out_818,
    output [511:0] col_out_819,
    output [511:0] col_out_820,
    output [511:0] col_out_821,
    output [511:0] col_out_822,
    output [511:0] col_out_823,
    output [511:0] col_out_824,
    output [511:0] col_out_825,
    output [511:0] col_out_826,
    output [511:0] col_out_827,
    output [511:0] col_out_828,
    output [511:0] col_out_829,
    output [511:0] col_out_830,
    output [511:0] col_out_831,
    output [511:0] col_out_832,
    output [511:0] col_out_833,
    output [511:0] col_out_834,
    output [511:0] col_out_835,
    output [511:0] col_out_836,
    output [511:0] col_out_837,
    output [511:0] col_out_838,
    output [511:0] col_out_839,
    output [511:0] col_out_840,
    output [511:0] col_out_841,
    output [511:0] col_out_842,
    output [511:0] col_out_843,
    output [511:0] col_out_844,
    output [511:0] col_out_845,
    output [511:0] col_out_846,
    output [511:0] col_out_847,
    output [511:0] col_out_848,
    output [511:0] col_out_849,
    output [511:0] col_out_850,
    output [511:0] col_out_851,
    output [511:0] col_out_852,
    output [511:0] col_out_853,
    output [511:0] col_out_854,
    output [511:0] col_out_855,
    output [511:0] col_out_856,
    output [511:0] col_out_857,
    output [511:0] col_out_858,
    output [511:0] col_out_859,
    output [511:0] col_out_860,
    output [511:0] col_out_861,
    output [511:0] col_out_862,
    output [511:0] col_out_863,
    output [511:0] col_out_864,
    output [511:0] col_out_865,
    output [511:0] col_out_866,
    output [511:0] col_out_867,
    output [511:0] col_out_868,
    output [511:0] col_out_869,
    output [511:0] col_out_870,
    output [511:0] col_out_871,
    output [511:0] col_out_872,
    output [511:0] col_out_873,
    output [511:0] col_out_874,
    output [511:0] col_out_875,
    output [511:0] col_out_876,
    output [511:0] col_out_877,
    output [511:0] col_out_878,
    output [511:0] col_out_879,
    output [511:0] col_out_880,
    output [511:0] col_out_881,
    output [511:0] col_out_882,
    output [511:0] col_out_883,
    output [511:0] col_out_884,
    output [511:0] col_out_885,
    output [511:0] col_out_886,
    output [511:0] col_out_887,
    output [511:0] col_out_888,
    output [511:0] col_out_889,
    output [511:0] col_out_890,
    output [511:0] col_out_891,
    output [511:0] col_out_892,
    output [511:0] col_out_893,
    output [511:0] col_out_894,
    output [511:0] col_out_895,
    output [511:0] col_out_896,
    output [511:0] col_out_897,
    output [511:0] col_out_898,
    output [511:0] col_out_899,
    output [511:0] col_out_900,
    output [511:0] col_out_901,
    output [511:0] col_out_902,
    output [511:0] col_out_903,
    output [511:0] col_out_904,
    output [511:0] col_out_905,
    output [511:0] col_out_906,
    output [511:0] col_out_907,
    output [511:0] col_out_908,
    output [511:0] col_out_909,
    output [511:0] col_out_910,
    output [511:0] col_out_911,
    output [511:0] col_out_912,
    output [511:0] col_out_913,
    output [511:0] col_out_914,
    output [511:0] col_out_915,
    output [511:0] col_out_916,
    output [511:0] col_out_917,
    output [511:0] col_out_918,
    output [511:0] col_out_919,
    output [511:0] col_out_920,
    output [511:0] col_out_921,
    output [511:0] col_out_922,
    output [511:0] col_out_923,
    output [511:0] col_out_924,
    output [511:0] col_out_925,
    output [511:0] col_out_926,
    output [511:0] col_out_927,
    output [511:0] col_out_928,
    output [511:0] col_out_929,
    output [511:0] col_out_930,
    output [511:0] col_out_931,
    output [511:0] col_out_932,
    output [511:0] col_out_933,
    output [511:0] col_out_934,
    output [511:0] col_out_935,
    output [511:0] col_out_936,
    output [511:0] col_out_937,
    output [511:0] col_out_938,
    output [511:0] col_out_939,
    output [511:0] col_out_940,
    output [511:0] col_out_941,
    output [511:0] col_out_942,
    output [511:0] col_out_943,
    output [511:0] col_out_944,
    output [511:0] col_out_945,
    output [511:0] col_out_946,
    output [511:0] col_out_947,
    output [511:0] col_out_948,
    output [511:0] col_out_949,
    output [511:0] col_out_950,
    output [511:0] col_out_951,
    output [511:0] col_out_952,
    output [511:0] col_out_953,
    output [511:0] col_out_954,
    output [511:0] col_out_955,
    output [511:0] col_out_956,
    output [511:0] col_out_957,
    output [511:0] col_out_958,
    output [511:0] col_out_959,
    output [511:0] col_out_960,
    output [511:0] col_out_961,
    output [511:0] col_out_962,
    output [511:0] col_out_963,
    output [511:0] col_out_964,
    output [511:0] col_out_965,
    output [511:0] col_out_966,
    output [511:0] col_out_967,
    output [511:0] col_out_968,
    output [511:0] col_out_969,
    output [511:0] col_out_970,
    output [511:0] col_out_971,
    output [511:0] col_out_972,
    output [511:0] col_out_973,
    output [511:0] col_out_974,
    output [511:0] col_out_975,
    output [511:0] col_out_976,
    output [511:0] col_out_977,
    output [511:0] col_out_978,
    output [511:0] col_out_979,
    output [511:0] col_out_980,
    output [511:0] col_out_981,
    output [511:0] col_out_982,
    output [511:0] col_out_983,
    output [511:0] col_out_984,
    output [511:0] col_out_985,
    output [511:0] col_out_986,
    output [511:0] col_out_987,
    output [511:0] col_out_988,
    output [511:0] col_out_989,
    output [511:0] col_out_990,
    output [511:0] col_out_991,
    output [511:0] col_out_992,
    output [511:0] col_out_993,
    output [511:0] col_out_994,
    output [511:0] col_out_995,
    output [511:0] col_out_996,
    output [511:0] col_out_997,
    output [511:0] col_out_998,
    output [511:0] col_out_999,
    output [511:0] col_out_1000,
    output [511:0] col_out_1001,
    output [511:0] col_out_1002,
    output [511:0] col_out_1003,
    output [511:0] col_out_1004,
    output [511:0] col_out_1005,
    output [511:0] col_out_1006,
    output [511:0] col_out_1007,
    output [511:0] col_out_1008,
    output [511:0] col_out_1009,
    output [511:0] col_out_1010,
    output [511:0] col_out_1011,
    output [511:0] col_out_1012,
    output [511:0] col_out_1013,
    output [511:0] col_out_1014,
    output [511:0] col_out_1015,
    output [511:0] col_out_1016,
    output [511:0] col_out_1017,
    output [511:0] col_out_1018,
    output [511:0] col_out_1019,
    output [511:0] col_out_1020,
    output [511:0] col_out_1021,
    output [511:0] col_out_1022,
    output [511:0] col_out_1023
);


// msq_half_product Outputs
wire [511:0] u0_col_out_0;
wire [511:0] u0_col_out_1;
wire [511:0] u0_col_out_2;
wire [511:0] u0_col_out_3;
wire [511:0] u0_col_out_4;
wire [511:0] u0_col_out_5;
wire [511:0] u0_col_out_6;
wire [511:0] u0_col_out_7;
wire [511:0] u0_col_out_8;
wire [511:0] u0_col_out_9;
wire [511:0] u0_col_out_10;
wire [511:0] u0_col_out_11;
wire [511:0] u0_col_out_12;
wire [511:0] u0_col_out_13;
wire [511:0] u0_col_out_14;
wire [511:0] u0_col_out_15;
wire [511:0] u0_col_out_16;
wire [511:0] u0_col_out_17;
wire [511:0] u0_col_out_18;
wire [511:0] u0_col_out_19;
wire [511:0] u0_col_out_20;
wire [511:0] u0_col_out_21;
wire [511:0] u0_col_out_22;
wire [511:0] u0_col_out_23;
wire [511:0] u0_col_out_24;
wire [511:0] u0_col_out_25;
wire [511:0] u0_col_out_26;
wire [511:0] u0_col_out_27;
wire [511:0] u0_col_out_28;
wire [511:0] u0_col_out_29;
wire [511:0] u0_col_out_30;
wire [511:0] u0_col_out_31;
wire [511:0] u0_col_out_32;
wire [511:0] u0_col_out_33;
wire [511:0] u0_col_out_34;
wire [511:0] u0_col_out_35;
wire [511:0] u0_col_out_36;
wire [511:0] u0_col_out_37;
wire [511:0] u0_col_out_38;
wire [511:0] u0_col_out_39;
wire [511:0] u0_col_out_40;
wire [511:0] u0_col_out_41;
wire [511:0] u0_col_out_42;
wire [511:0] u0_col_out_43;
wire [511:0] u0_col_out_44;
wire [511:0] u0_col_out_45;
wire [511:0] u0_col_out_46;
wire [511:0] u0_col_out_47;
wire [511:0] u0_col_out_48;
wire [511:0] u0_col_out_49;
wire [511:0] u0_col_out_50;
wire [511:0] u0_col_out_51;
wire [511:0] u0_col_out_52;
wire [511:0] u0_col_out_53;
wire [511:0] u0_col_out_54;
wire [511:0] u0_col_out_55;
wire [511:0] u0_col_out_56;
wire [511:0] u0_col_out_57;
wire [511:0] u0_col_out_58;
wire [511:0] u0_col_out_59;
wire [511:0] u0_col_out_60;
wire [511:0] u0_col_out_61;
wire [511:0] u0_col_out_62;
wire [511:0] u0_col_out_63;
wire [511:0] u0_col_out_64;
wire [511:0] u0_col_out_65;
wire [511:0] u0_col_out_66;
wire [511:0] u0_col_out_67;
wire [511:0] u0_col_out_68;
wire [511:0] u0_col_out_69;
wire [511:0] u0_col_out_70;
wire [511:0] u0_col_out_71;
wire [511:0] u0_col_out_72;
wire [511:0] u0_col_out_73;
wire [511:0] u0_col_out_74;
wire [511:0] u0_col_out_75;
wire [511:0] u0_col_out_76;
wire [511:0] u0_col_out_77;
wire [511:0] u0_col_out_78;
wire [511:0] u0_col_out_79;
wire [511:0] u0_col_out_80;
wire [511:0] u0_col_out_81;
wire [511:0] u0_col_out_82;
wire [511:0] u0_col_out_83;
wire [511:0] u0_col_out_84;
wire [511:0] u0_col_out_85;
wire [511:0] u0_col_out_86;
wire [511:0] u0_col_out_87;
wire [511:0] u0_col_out_88;
wire [511:0] u0_col_out_89;
wire [511:0] u0_col_out_90;
wire [511:0] u0_col_out_91;
wire [511:0] u0_col_out_92;
wire [511:0] u0_col_out_93;
wire [511:0] u0_col_out_94;
wire [511:0] u0_col_out_95;
wire [511:0] u0_col_out_96;
wire [511:0] u0_col_out_97;
wire [511:0] u0_col_out_98;
wire [511:0] u0_col_out_99;
wire [511:0] u0_col_out_100;
wire [511:0] u0_col_out_101;
wire [511:0] u0_col_out_102;
wire [511:0] u0_col_out_103;
wire [511:0] u0_col_out_104;
wire [511:0] u0_col_out_105;
wire [511:0] u0_col_out_106;
wire [511:0] u0_col_out_107;
wire [511:0] u0_col_out_108;
wire [511:0] u0_col_out_109;
wire [511:0] u0_col_out_110;
wire [511:0] u0_col_out_111;
wire [511:0] u0_col_out_112;
wire [511:0] u0_col_out_113;
wire [511:0] u0_col_out_114;
wire [511:0] u0_col_out_115;
wire [511:0] u0_col_out_116;
wire [511:0] u0_col_out_117;
wire [511:0] u0_col_out_118;
wire [511:0] u0_col_out_119;
wire [511:0] u0_col_out_120;
wire [511:0] u0_col_out_121;
wire [511:0] u0_col_out_122;
wire [511:0] u0_col_out_123;
wire [511:0] u0_col_out_124;
wire [511:0] u0_col_out_125;
wire [511:0] u0_col_out_126;
wire [511:0] u0_col_out_127;
wire [511:0] u0_col_out_128;
wire [511:0] u0_col_out_129;
wire [511:0] u0_col_out_130;
wire [511:0] u0_col_out_131;
wire [511:0] u0_col_out_132;
wire [511:0] u0_col_out_133;
wire [511:0] u0_col_out_134;
wire [511:0] u0_col_out_135;
wire [511:0] u0_col_out_136;
wire [511:0] u0_col_out_137;
wire [511:0] u0_col_out_138;
wire [511:0] u0_col_out_139;
wire [511:0] u0_col_out_140;
wire [511:0] u0_col_out_141;
wire [511:0] u0_col_out_142;
wire [511:0] u0_col_out_143;
wire [511:0] u0_col_out_144;
wire [511:0] u0_col_out_145;
wire [511:0] u0_col_out_146;
wire [511:0] u0_col_out_147;
wire [511:0] u0_col_out_148;
wire [511:0] u0_col_out_149;
wire [511:0] u0_col_out_150;
wire [511:0] u0_col_out_151;
wire [511:0] u0_col_out_152;
wire [511:0] u0_col_out_153;
wire [511:0] u0_col_out_154;
wire [511:0] u0_col_out_155;
wire [511:0] u0_col_out_156;
wire [511:0] u0_col_out_157;
wire [511:0] u0_col_out_158;
wire [511:0] u0_col_out_159;
wire [511:0] u0_col_out_160;
wire [511:0] u0_col_out_161;
wire [511:0] u0_col_out_162;
wire [511:0] u0_col_out_163;
wire [511:0] u0_col_out_164;
wire [511:0] u0_col_out_165;
wire [511:0] u0_col_out_166;
wire [511:0] u0_col_out_167;
wire [511:0] u0_col_out_168;
wire [511:0] u0_col_out_169;
wire [511:0] u0_col_out_170;
wire [511:0] u0_col_out_171;
wire [511:0] u0_col_out_172;
wire [511:0] u0_col_out_173;
wire [511:0] u0_col_out_174;
wire [511:0] u0_col_out_175;
wire [511:0] u0_col_out_176;
wire [511:0] u0_col_out_177;
wire [511:0] u0_col_out_178;
wire [511:0] u0_col_out_179;
wire [511:0] u0_col_out_180;
wire [511:0] u0_col_out_181;
wire [511:0] u0_col_out_182;
wire [511:0] u0_col_out_183;
wire [511:0] u0_col_out_184;
wire [511:0] u0_col_out_185;
wire [511:0] u0_col_out_186;
wire [511:0] u0_col_out_187;
wire [511:0] u0_col_out_188;
wire [511:0] u0_col_out_189;
wire [511:0] u0_col_out_190;
wire [511:0] u0_col_out_191;
wire [511:0] u0_col_out_192;
wire [511:0] u0_col_out_193;
wire [511:0] u0_col_out_194;
wire [511:0] u0_col_out_195;
wire [511:0] u0_col_out_196;
wire [511:0] u0_col_out_197;
wire [511:0] u0_col_out_198;
wire [511:0] u0_col_out_199;
wire [511:0] u0_col_out_200;
wire [511:0] u0_col_out_201;
wire [511:0] u0_col_out_202;
wire [511:0] u0_col_out_203;
wire [511:0] u0_col_out_204;
wire [511:0] u0_col_out_205;
wire [511:0] u0_col_out_206;
wire [511:0] u0_col_out_207;
wire [511:0] u0_col_out_208;
wire [511:0] u0_col_out_209;
wire [511:0] u0_col_out_210;
wire [511:0] u0_col_out_211;
wire [511:0] u0_col_out_212;
wire [511:0] u0_col_out_213;
wire [511:0] u0_col_out_214;
wire [511:0] u0_col_out_215;
wire [511:0] u0_col_out_216;
wire [511:0] u0_col_out_217;
wire [511:0] u0_col_out_218;
wire [511:0] u0_col_out_219;
wire [511:0] u0_col_out_220;
wire [511:0] u0_col_out_221;
wire [511:0] u0_col_out_222;
wire [511:0] u0_col_out_223;
wire [511:0] u0_col_out_224;
wire [511:0] u0_col_out_225;
wire [511:0] u0_col_out_226;
wire [511:0] u0_col_out_227;
wire [511:0] u0_col_out_228;
wire [511:0] u0_col_out_229;
wire [511:0] u0_col_out_230;
wire [511:0] u0_col_out_231;
wire [511:0] u0_col_out_232;
wire [511:0] u0_col_out_233;
wire [511:0] u0_col_out_234;
wire [511:0] u0_col_out_235;
wire [511:0] u0_col_out_236;
wire [511:0] u0_col_out_237;
wire [511:0] u0_col_out_238;
wire [511:0] u0_col_out_239;
wire [511:0] u0_col_out_240;
wire [511:0] u0_col_out_241;
wire [511:0] u0_col_out_242;
wire [511:0] u0_col_out_243;
wire [511:0] u0_col_out_244;
wire [511:0] u0_col_out_245;
wire [511:0] u0_col_out_246;
wire [511:0] u0_col_out_247;
wire [511:0] u0_col_out_248;
wire [511:0] u0_col_out_249;
wire [511:0] u0_col_out_250;
wire [511:0] u0_col_out_251;
wire [511:0] u0_col_out_252;
wire [511:0] u0_col_out_253;
wire [511:0] u0_col_out_254;
wire [511:0] u0_col_out_255;
wire [511:0] u0_col_out_256;
wire [511:0] u0_col_out_257;
wire [511:0] u0_col_out_258;
wire [511:0] u0_col_out_259;
wire [511:0] u0_col_out_260;
wire [511:0] u0_col_out_261;
wire [511:0] u0_col_out_262;
wire [511:0] u0_col_out_263;
wire [511:0] u0_col_out_264;
wire [511:0] u0_col_out_265;
wire [511:0] u0_col_out_266;
wire [511:0] u0_col_out_267;
wire [511:0] u0_col_out_268;
wire [511:0] u0_col_out_269;
wire [511:0] u0_col_out_270;
wire [511:0] u0_col_out_271;
wire [511:0] u0_col_out_272;
wire [511:0] u0_col_out_273;
wire [511:0] u0_col_out_274;
wire [511:0] u0_col_out_275;
wire [511:0] u0_col_out_276;
wire [511:0] u0_col_out_277;
wire [511:0] u0_col_out_278;
wire [511:0] u0_col_out_279;
wire [511:0] u0_col_out_280;
wire [511:0] u0_col_out_281;
wire [511:0] u0_col_out_282;
wire [511:0] u0_col_out_283;
wire [511:0] u0_col_out_284;
wire [511:0] u0_col_out_285;
wire [511:0] u0_col_out_286;
wire [511:0] u0_col_out_287;
wire [511:0] u0_col_out_288;
wire [511:0] u0_col_out_289;
wire [511:0] u0_col_out_290;
wire [511:0] u0_col_out_291;
wire [511:0] u0_col_out_292;
wire [511:0] u0_col_out_293;
wire [511:0] u0_col_out_294;
wire [511:0] u0_col_out_295;
wire [511:0] u0_col_out_296;
wire [511:0] u0_col_out_297;
wire [511:0] u0_col_out_298;
wire [511:0] u0_col_out_299;
wire [511:0] u0_col_out_300;
wire [511:0] u0_col_out_301;
wire [511:0] u0_col_out_302;
wire [511:0] u0_col_out_303;
wire [511:0] u0_col_out_304;
wire [511:0] u0_col_out_305;
wire [511:0] u0_col_out_306;
wire [511:0] u0_col_out_307;
wire [511:0] u0_col_out_308;
wire [511:0] u0_col_out_309;
wire [511:0] u0_col_out_310;
wire [511:0] u0_col_out_311;
wire [511:0] u0_col_out_312;
wire [511:0] u0_col_out_313;
wire [511:0] u0_col_out_314;
wire [511:0] u0_col_out_315;
wire [511:0] u0_col_out_316;
wire [511:0] u0_col_out_317;
wire [511:0] u0_col_out_318;
wire [511:0] u0_col_out_319;
wire [511:0] u0_col_out_320;
wire [511:0] u0_col_out_321;
wire [511:0] u0_col_out_322;
wire [511:0] u0_col_out_323;
wire [511:0] u0_col_out_324;
wire [511:0] u0_col_out_325;
wire [511:0] u0_col_out_326;
wire [511:0] u0_col_out_327;
wire [511:0] u0_col_out_328;
wire [511:0] u0_col_out_329;
wire [511:0] u0_col_out_330;
wire [511:0] u0_col_out_331;
wire [511:0] u0_col_out_332;
wire [511:0] u0_col_out_333;
wire [511:0] u0_col_out_334;
wire [511:0] u0_col_out_335;
wire [511:0] u0_col_out_336;
wire [511:0] u0_col_out_337;
wire [511:0] u0_col_out_338;
wire [511:0] u0_col_out_339;
wire [511:0] u0_col_out_340;
wire [511:0] u0_col_out_341;
wire [511:0] u0_col_out_342;
wire [511:0] u0_col_out_343;
wire [511:0] u0_col_out_344;
wire [511:0] u0_col_out_345;
wire [511:0] u0_col_out_346;
wire [511:0] u0_col_out_347;
wire [511:0] u0_col_out_348;
wire [511:0] u0_col_out_349;
wire [511:0] u0_col_out_350;
wire [511:0] u0_col_out_351;
wire [511:0] u0_col_out_352;
wire [511:0] u0_col_out_353;
wire [511:0] u0_col_out_354;
wire [511:0] u0_col_out_355;
wire [511:0] u0_col_out_356;
wire [511:0] u0_col_out_357;
wire [511:0] u0_col_out_358;
wire [511:0] u0_col_out_359;
wire [511:0] u0_col_out_360;
wire [511:0] u0_col_out_361;
wire [511:0] u0_col_out_362;
wire [511:0] u0_col_out_363;
wire [511:0] u0_col_out_364;
wire [511:0] u0_col_out_365;
wire [511:0] u0_col_out_366;
wire [511:0] u0_col_out_367;
wire [511:0] u0_col_out_368;
wire [511:0] u0_col_out_369;
wire [511:0] u0_col_out_370;
wire [511:0] u0_col_out_371;
wire [511:0] u0_col_out_372;
wire [511:0] u0_col_out_373;
wire [511:0] u0_col_out_374;
wire [511:0] u0_col_out_375;
wire [511:0] u0_col_out_376;
wire [511:0] u0_col_out_377;
wire [511:0] u0_col_out_378;
wire [511:0] u0_col_out_379;
wire [511:0] u0_col_out_380;
wire [511:0] u0_col_out_381;
wire [511:0] u0_col_out_382;
wire [511:0] u0_col_out_383;
wire [511:0] u0_col_out_384;
wire [511:0] u0_col_out_385;
wire [511:0] u0_col_out_386;
wire [511:0] u0_col_out_387;
wire [511:0] u0_col_out_388;
wire [511:0] u0_col_out_389;
wire [511:0] u0_col_out_390;
wire [511:0] u0_col_out_391;
wire [511:0] u0_col_out_392;
wire [511:0] u0_col_out_393;
wire [511:0] u0_col_out_394;
wire [511:0] u0_col_out_395;
wire [511:0] u0_col_out_396;
wire [511:0] u0_col_out_397;
wire [511:0] u0_col_out_398;
wire [511:0] u0_col_out_399;
wire [511:0] u0_col_out_400;
wire [511:0] u0_col_out_401;
wire [511:0] u0_col_out_402;
wire [511:0] u0_col_out_403;
wire [511:0] u0_col_out_404;
wire [511:0] u0_col_out_405;
wire [511:0] u0_col_out_406;
wire [511:0] u0_col_out_407;
wire [511:0] u0_col_out_408;
wire [511:0] u0_col_out_409;
wire [511:0] u0_col_out_410;
wire [511:0] u0_col_out_411;
wire [511:0] u0_col_out_412;
wire [511:0] u0_col_out_413;
wire [511:0] u0_col_out_414;
wire [511:0] u0_col_out_415;
wire [511:0] u0_col_out_416;
wire [511:0] u0_col_out_417;
wire [511:0] u0_col_out_418;
wire [511:0] u0_col_out_419;
wire [511:0] u0_col_out_420;
wire [511:0] u0_col_out_421;
wire [511:0] u0_col_out_422;
wire [511:0] u0_col_out_423;
wire [511:0] u0_col_out_424;
wire [511:0] u0_col_out_425;
wire [511:0] u0_col_out_426;
wire [511:0] u0_col_out_427;
wire [511:0] u0_col_out_428;
wire [511:0] u0_col_out_429;
wire [511:0] u0_col_out_430;
wire [511:0] u0_col_out_431;
wire [511:0] u0_col_out_432;
wire [511:0] u0_col_out_433;
wire [511:0] u0_col_out_434;
wire [511:0] u0_col_out_435;
wire [511:0] u0_col_out_436;
wire [511:0] u0_col_out_437;
wire [511:0] u0_col_out_438;
wire [511:0] u0_col_out_439;
wire [511:0] u0_col_out_440;
wire [511:0] u0_col_out_441;
wire [511:0] u0_col_out_442;
wire [511:0] u0_col_out_443;
wire [511:0] u0_col_out_444;
wire [511:0] u0_col_out_445;
wire [511:0] u0_col_out_446;
wire [511:0] u0_col_out_447;
wire [511:0] u0_col_out_448;
wire [511:0] u0_col_out_449;
wire [511:0] u0_col_out_450;
wire [511:0] u0_col_out_451;
wire [511:0] u0_col_out_452;
wire [511:0] u0_col_out_453;
wire [511:0] u0_col_out_454;
wire [511:0] u0_col_out_455;
wire [511:0] u0_col_out_456;
wire [511:0] u0_col_out_457;
wire [511:0] u0_col_out_458;
wire [511:0] u0_col_out_459;
wire [511:0] u0_col_out_460;
wire [511:0] u0_col_out_461;
wire [511:0] u0_col_out_462;
wire [511:0] u0_col_out_463;
wire [511:0] u0_col_out_464;
wire [511:0] u0_col_out_465;
wire [511:0] u0_col_out_466;
wire [511:0] u0_col_out_467;
wire [511:0] u0_col_out_468;
wire [511:0] u0_col_out_469;
wire [511:0] u0_col_out_470;
wire [511:0] u0_col_out_471;
wire [511:0] u0_col_out_472;
wire [511:0] u0_col_out_473;
wire [511:0] u0_col_out_474;
wire [511:0] u0_col_out_475;
wire [511:0] u0_col_out_476;
wire [511:0] u0_col_out_477;
wire [511:0] u0_col_out_478;
wire [511:0] u0_col_out_479;
wire [511:0] u0_col_out_480;
wire [511:0] u0_col_out_481;
wire [511:0] u0_col_out_482;
wire [511:0] u0_col_out_483;
wire [511:0] u0_col_out_484;
wire [511:0] u0_col_out_485;
wire [511:0] u0_col_out_486;
wire [511:0] u0_col_out_487;
wire [511:0] u0_col_out_488;
wire [511:0] u0_col_out_489;
wire [511:0] u0_col_out_490;
wire [511:0] u0_col_out_491;
wire [511:0] u0_col_out_492;
wire [511:0] u0_col_out_493;
wire [511:0] u0_col_out_494;
wire [511:0] u0_col_out_495;
wire [511:0] u0_col_out_496;
wire [511:0] u0_col_out_497;
wire [511:0] u0_col_out_498;
wire [511:0] u0_col_out_499;
wire [511:0] u0_col_out_500;
wire [511:0] u0_col_out_501;
wire [511:0] u0_col_out_502;
wire [511:0] u0_col_out_503;
wire [511:0] u0_col_out_504;
wire [511:0] u0_col_out_505;
wire [511:0] u0_col_out_506;
wire [511:0] u0_col_out_507;
wire [511:0] u0_col_out_508;
wire [511:0] u0_col_out_509;
wire [511:0] u0_col_out_510;
wire [511:0] u0_col_out_511;
wire [511:0] u0_col_out_512;
wire [511:0] u0_col_out_513;
wire [511:0] u0_col_out_514;
wire [511:0] u0_col_out_515;
wire [511:0] u0_col_out_516;
wire [511:0] u0_col_out_517;
wire [511:0] u0_col_out_518;
wire [511:0] u0_col_out_519;
wire [511:0] u0_col_out_520;
wire [511:0] u0_col_out_521;
wire [511:0] u0_col_out_522;
wire [511:0] u0_col_out_523;
wire [511:0] u0_col_out_524;
wire [511:0] u0_col_out_525;
wire [511:0] u0_col_out_526;
wire [511:0] u0_col_out_527;
wire [511:0] u0_col_out_528;
wire [511:0] u0_col_out_529;
wire [511:0] u0_col_out_530;
wire [511:0] u0_col_out_531;
wire [511:0] u0_col_out_532;
wire [511:0] u0_col_out_533;
wire [511:0] u0_col_out_534;
wire [511:0] u0_col_out_535;
wire [511:0] u0_col_out_536;
wire [511:0] u0_col_out_537;
wire [511:0] u0_col_out_538;
wire [511:0] u0_col_out_539;
wire [511:0] u0_col_out_540;
wire [511:0] u0_col_out_541;
wire [511:0] u0_col_out_542;
wire [511:0] u0_col_out_543;
wire [511:0] u0_col_out_544;
wire [511:0] u0_col_out_545;
wire [511:0] u0_col_out_546;
wire [511:0] u0_col_out_547;
wire [511:0] u0_col_out_548;
wire [511:0] u0_col_out_549;
wire [511:0] u0_col_out_550;
wire [511:0] u0_col_out_551;
wire [511:0] u0_col_out_552;
wire [511:0] u0_col_out_553;
wire [511:0] u0_col_out_554;
wire [511:0] u0_col_out_555;
wire [511:0] u0_col_out_556;
wire [511:0] u0_col_out_557;
wire [511:0] u0_col_out_558;
wire [511:0] u0_col_out_559;
wire [511:0] u0_col_out_560;
wire [511:0] u0_col_out_561;
wire [511:0] u0_col_out_562;
wire [511:0] u0_col_out_563;
wire [511:0] u0_col_out_564;
wire [511:0] u0_col_out_565;
wire [511:0] u0_col_out_566;
wire [511:0] u0_col_out_567;
wire [511:0] u0_col_out_568;
wire [511:0] u0_col_out_569;
wire [511:0] u0_col_out_570;
wire [511:0] u0_col_out_571;
wire [511:0] u0_col_out_572;
wire [511:0] u0_col_out_573;
wire [511:0] u0_col_out_574;
wire [511:0] u0_col_out_575;
wire [511:0] u0_col_out_576;
wire [511:0] u0_col_out_577;
wire [511:0] u0_col_out_578;
wire [511:0] u0_col_out_579;
wire [511:0] u0_col_out_580;
wire [511:0] u0_col_out_581;
wire [511:0] u0_col_out_582;
wire [511:0] u0_col_out_583;
wire [511:0] u0_col_out_584;
wire [511:0] u0_col_out_585;
wire [511:0] u0_col_out_586;
wire [511:0] u0_col_out_587;
wire [511:0] u0_col_out_588;
wire [511:0] u0_col_out_589;
wire [511:0] u0_col_out_590;
wire [511:0] u0_col_out_591;
wire [511:0] u0_col_out_592;
wire [511:0] u0_col_out_593;
wire [511:0] u0_col_out_594;
wire [511:0] u0_col_out_595;
wire [511:0] u0_col_out_596;
wire [511:0] u0_col_out_597;
wire [511:0] u0_col_out_598;
wire [511:0] u0_col_out_599;
wire [511:0] u0_col_out_600;
wire [511:0] u0_col_out_601;
wire [511:0] u0_col_out_602;
wire [511:0] u0_col_out_603;
wire [511:0] u0_col_out_604;
wire [511:0] u0_col_out_605;
wire [511:0] u0_col_out_606;
wire [511:0] u0_col_out_607;
wire [511:0] u0_col_out_608;
wire [511:0] u0_col_out_609;
wire [511:0] u0_col_out_610;
wire [511:0] u0_col_out_611;
wire [511:0] u0_col_out_612;
wire [511:0] u0_col_out_613;
wire [511:0] u0_col_out_614;
wire [511:0] u0_col_out_615;
wire [511:0] u0_col_out_616;
wire [511:0] u0_col_out_617;
wire [511:0] u0_col_out_618;
wire [511:0] u0_col_out_619;
wire [511:0] u0_col_out_620;
wire [511:0] u0_col_out_621;
wire [511:0] u0_col_out_622;
wire [511:0] u0_col_out_623;
wire [511:0] u0_col_out_624;
wire [511:0] u0_col_out_625;
wire [511:0] u0_col_out_626;
wire [511:0] u0_col_out_627;
wire [511:0] u0_col_out_628;
wire [511:0] u0_col_out_629;
wire [511:0] u0_col_out_630;
wire [511:0] u0_col_out_631;
wire [511:0] u0_col_out_632;
wire [511:0] u0_col_out_633;
wire [511:0] u0_col_out_634;
wire [511:0] u0_col_out_635;
wire [511:0] u0_col_out_636;
wire [511:0] u0_col_out_637;
wire [511:0] u0_col_out_638;
wire [511:0] u0_col_out_639;
wire [511:0] u0_col_out_640;
wire [511:0] u0_col_out_641;
wire [511:0] u0_col_out_642;
wire [511:0] u0_col_out_643;
wire [511:0] u0_col_out_644;
wire [511:0] u0_col_out_645;
wire [511:0] u0_col_out_646;
wire [511:0] u0_col_out_647;
wire [511:0] u0_col_out_648;
wire [511:0] u0_col_out_649;
wire [511:0] u0_col_out_650;
wire [511:0] u0_col_out_651;
wire [511:0] u0_col_out_652;
wire [511:0] u0_col_out_653;
wire [511:0] u0_col_out_654;
wire [511:0] u0_col_out_655;
wire [511:0] u0_col_out_656;
wire [511:0] u0_col_out_657;
wire [511:0] u0_col_out_658;
wire [511:0] u0_col_out_659;
wire [511:0] u0_col_out_660;
wire [511:0] u0_col_out_661;
wire [511:0] u0_col_out_662;
wire [511:0] u0_col_out_663;
wire [511:0] u0_col_out_664;
wire [511:0] u0_col_out_665;
wire [511:0] u0_col_out_666;
wire [511:0] u0_col_out_667;
wire [511:0] u0_col_out_668;
wire [511:0] u0_col_out_669;
wire [511:0] u0_col_out_670;
wire [511:0] u0_col_out_671;
wire [511:0] u0_col_out_672;
wire [511:0] u0_col_out_673;
wire [511:0] u0_col_out_674;
wire [511:0] u0_col_out_675;
wire [511:0] u0_col_out_676;
wire [511:0] u0_col_out_677;
wire [511:0] u0_col_out_678;
wire [511:0] u0_col_out_679;
wire [511:0] u0_col_out_680;
wire [511:0] u0_col_out_681;
wire [511:0] u0_col_out_682;
wire [511:0] u0_col_out_683;
wire [511:0] u0_col_out_684;
wire [511:0] u0_col_out_685;
wire [511:0] u0_col_out_686;
wire [511:0] u0_col_out_687;
wire [511:0] u0_col_out_688;
wire [511:0] u0_col_out_689;
wire [511:0] u0_col_out_690;
wire [511:0] u0_col_out_691;
wire [511:0] u0_col_out_692;
wire [511:0] u0_col_out_693;
wire [511:0] u0_col_out_694;
wire [511:0] u0_col_out_695;
wire [511:0] u0_col_out_696;
wire [511:0] u0_col_out_697;
wire [511:0] u0_col_out_698;
wire [511:0] u0_col_out_699;
wire [511:0] u0_col_out_700;
wire [511:0] u0_col_out_701;
wire [511:0] u0_col_out_702;
wire [511:0] u0_col_out_703;
wire [511:0] u0_col_out_704;
wire [511:0] u0_col_out_705;
wire [511:0] u0_col_out_706;
wire [511:0] u0_col_out_707;
wire [511:0] u0_col_out_708;
wire [511:0] u0_col_out_709;
wire [511:0] u0_col_out_710;
wire [511:0] u0_col_out_711;
wire [511:0] u0_col_out_712;
wire [511:0] u0_col_out_713;
wire [511:0] u0_col_out_714;
wire [511:0] u0_col_out_715;
wire [511:0] u0_col_out_716;
wire [511:0] u0_col_out_717;
wire [511:0] u0_col_out_718;
wire [511:0] u0_col_out_719;
wire [511:0] u0_col_out_720;
wire [511:0] u0_col_out_721;
wire [511:0] u0_col_out_722;
wire [511:0] u0_col_out_723;
wire [511:0] u0_col_out_724;
wire [511:0] u0_col_out_725;
wire [511:0] u0_col_out_726;
wire [511:0] u0_col_out_727;
wire [511:0] u0_col_out_728;
wire [511:0] u0_col_out_729;
wire [511:0] u0_col_out_730;
wire [511:0] u0_col_out_731;
wire [511:0] u0_col_out_732;
wire [511:0] u0_col_out_733;
wire [511:0] u0_col_out_734;
wire [511:0] u0_col_out_735;
wire [511:0] u0_col_out_736;
wire [511:0] u0_col_out_737;
wire [511:0] u0_col_out_738;
wire [511:0] u0_col_out_739;
wire [511:0] u0_col_out_740;
wire [511:0] u0_col_out_741;
wire [511:0] u0_col_out_742;
wire [511:0] u0_col_out_743;
wire [511:0] u0_col_out_744;
wire [511:0] u0_col_out_745;
wire [511:0] u0_col_out_746;
wire [511:0] u0_col_out_747;
wire [511:0] u0_col_out_748;
wire [511:0] u0_col_out_749;
wire [511:0] u0_col_out_750;
wire [511:0] u0_col_out_751;
wire [511:0] u0_col_out_752;
wire [511:0] u0_col_out_753;
wire [511:0] u0_col_out_754;
wire [511:0] u0_col_out_755;
wire [511:0] u0_col_out_756;
wire [511:0] u0_col_out_757;
wire [511:0] u0_col_out_758;
wire [511:0] u0_col_out_759;
wire [511:0] u0_col_out_760;
wire [511:0] u0_col_out_761;
wire [511:0] u0_col_out_762;
wire [511:0] u0_col_out_763;
wire [511:0] u0_col_out_764;
wire [511:0] u0_col_out_765;
wire [511:0] u0_col_out_766;
wire [511:0] u0_col_out_767;
wire [511:0] u0_col_out_768;
wire [511:0] u0_col_out_769;
wire [511:0] u0_col_out_770;
wire [511:0] u0_col_out_771;
wire [511:0] u0_col_out_772;
wire [511:0] u0_col_out_773;
wire [511:0] u0_col_out_774;
wire [511:0] u0_col_out_775;
wire [511:0] u0_col_out_776;
wire [511:0] u0_col_out_777;
wire [511:0] u0_col_out_778;
wire [511:0] u0_col_out_779;
wire [511:0] u0_col_out_780;
wire [511:0] u0_col_out_781;
wire [511:0] u0_col_out_782;
wire [511:0] u0_col_out_783;
wire [511:0] u0_col_out_784;
wire [511:0] u0_col_out_785;
wire [511:0] u0_col_out_786;
wire [511:0] u0_col_out_787;
wire [511:0] u0_col_out_788;
wire [511:0] u0_col_out_789;
wire [511:0] u0_col_out_790;
wire [511:0] u0_col_out_791;
wire [511:0] u0_col_out_792;
wire [511:0] u0_col_out_793;
wire [511:0] u0_col_out_794;
wire [511:0] u0_col_out_795;
wire [511:0] u0_col_out_796;
wire [511:0] u0_col_out_797;
wire [511:0] u0_col_out_798;
wire [511:0] u0_col_out_799;
wire [511:0] u0_col_out_800;
wire [511:0] u0_col_out_801;
wire [511:0] u0_col_out_802;
wire [511:0] u0_col_out_803;
wire [511:0] u0_col_out_804;
wire [511:0] u0_col_out_805;
wire [511:0] u0_col_out_806;
wire [511:0] u0_col_out_807;
wire [511:0] u0_col_out_808;
wire [511:0] u0_col_out_809;
wire [511:0] u0_col_out_810;
wire [511:0] u0_col_out_811;
wire [511:0] u0_col_out_812;
wire [511:0] u0_col_out_813;
wire [511:0] u0_col_out_814;
wire [511:0] u0_col_out_815;
wire [511:0] u0_col_out_816;
wire [511:0] u0_col_out_817;
wire [511:0] u0_col_out_818;
wire [511:0] u0_col_out_819;
wire [511:0] u0_col_out_820;
wire [511:0] u0_col_out_821;
wire [511:0] u0_col_out_822;
wire [511:0] u0_col_out_823;
wire [511:0] u0_col_out_824;
wire [511:0] u0_col_out_825;
wire [511:0] u0_col_out_826;
wire [511:0] u0_col_out_827;
wire [511:0] u0_col_out_828;
wire [511:0] u0_col_out_829;
wire [511:0] u0_col_out_830;
wire [511:0] u0_col_out_831;
wire [511:0] u0_col_out_832;
wire [511:0] u0_col_out_833;
wire [511:0] u0_col_out_834;
wire [511:0] u0_col_out_835;
wire [511:0] u0_col_out_836;
wire [511:0] u0_col_out_837;
wire [511:0] u0_col_out_838;
wire [511:0] u0_col_out_839;
wire [511:0] u0_col_out_840;
wire [511:0] u0_col_out_841;
wire [511:0] u0_col_out_842;
wire [511:0] u0_col_out_843;
wire [511:0] u0_col_out_844;
wire [511:0] u0_col_out_845;
wire [511:0] u0_col_out_846;
wire [511:0] u0_col_out_847;
wire [511:0] u0_col_out_848;
wire [511:0] u0_col_out_849;
wire [511:0] u0_col_out_850;
wire [511:0] u0_col_out_851;
wire [511:0] u0_col_out_852;
wire [511:0] u0_col_out_853;
wire [511:0] u0_col_out_854;
wire [511:0] u0_col_out_855;
wire [511:0] u0_col_out_856;
wire [511:0] u0_col_out_857;
wire [511:0] u0_col_out_858;
wire [511:0] u0_col_out_859;
wire [511:0] u0_col_out_860;
wire [511:0] u0_col_out_861;
wire [511:0] u0_col_out_862;
wire [511:0] u0_col_out_863;
wire [511:0] u0_col_out_864;
wire [511:0] u0_col_out_865;
wire [511:0] u0_col_out_866;
wire [511:0] u0_col_out_867;
wire [511:0] u0_col_out_868;
wire [511:0] u0_col_out_869;
wire [511:0] u0_col_out_870;
wire [511:0] u0_col_out_871;
wire [511:0] u0_col_out_872;
wire [511:0] u0_col_out_873;
wire [511:0] u0_col_out_874;
wire [511:0] u0_col_out_875;
wire [511:0] u0_col_out_876;
wire [511:0] u0_col_out_877;
wire [511:0] u0_col_out_878;
wire [511:0] u0_col_out_879;
wire [511:0] u0_col_out_880;
wire [511:0] u0_col_out_881;
wire [511:0] u0_col_out_882;
wire [511:0] u0_col_out_883;
wire [511:0] u0_col_out_884;
wire [511:0] u0_col_out_885;
wire [511:0] u0_col_out_886;
wire [511:0] u0_col_out_887;
wire [511:0] u0_col_out_888;
wire [511:0] u0_col_out_889;
wire [511:0] u0_col_out_890;
wire [511:0] u0_col_out_891;
wire [511:0] u0_col_out_892;
wire [511:0] u0_col_out_893;
wire [511:0] u0_col_out_894;
wire [511:0] u0_col_out_895;
wire [511:0] u0_col_out_896;
wire [511:0] u0_col_out_897;
wire [511:0] u0_col_out_898;
wire [511:0] u0_col_out_899;
wire [511:0] u0_col_out_900;
wire [511:0] u0_col_out_901;
wire [511:0] u0_col_out_902;
wire [511:0] u0_col_out_903;
wire [511:0] u0_col_out_904;
wire [511:0] u0_col_out_905;
wire [511:0] u0_col_out_906;
wire [511:0] u0_col_out_907;
wire [511:0] u0_col_out_908;
wire [511:0] u0_col_out_909;
wire [511:0] u0_col_out_910;
wire [511:0] u0_col_out_911;
wire [511:0] u0_col_out_912;
wire [511:0] u0_col_out_913;
wire [511:0] u0_col_out_914;
wire [511:0] u0_col_out_915;
wire [511:0] u0_col_out_916;
wire [511:0] u0_col_out_917;
wire [511:0] u0_col_out_918;
wire [511:0] u0_col_out_919;
wire [511:0] u0_col_out_920;
wire [511:0] u0_col_out_921;
wire [511:0] u0_col_out_922;
wire [511:0] u0_col_out_923;
wire [511:0] u0_col_out_924;
wire [511:0] u0_col_out_925;
wire [511:0] u0_col_out_926;
wire [511:0] u0_col_out_927;
wire [511:0] u0_col_out_928;
wire [511:0] u0_col_out_929;
wire [511:0] u0_col_out_930;
wire [511:0] u0_col_out_931;
wire [511:0] u0_col_out_932;
wire [511:0] u0_col_out_933;
wire [511:0] u0_col_out_934;
wire [511:0] u0_col_out_935;
wire [511:0] u0_col_out_936;
wire [511:0] u0_col_out_937;
wire [511:0] u0_col_out_938;
wire [511:0] u0_col_out_939;
wire [511:0] u0_col_out_940;
wire [511:0] u0_col_out_941;
wire [511:0] u0_col_out_942;
wire [511:0] u0_col_out_943;
wire [511:0] u0_col_out_944;
wire [511:0] u0_col_out_945;
wire [511:0] u0_col_out_946;
wire [511:0] u0_col_out_947;
wire [511:0] u0_col_out_948;
wire [511:0] u0_col_out_949;
wire [511:0] u0_col_out_950;
wire [511:0] u0_col_out_951;
wire [511:0] u0_col_out_952;
wire [511:0] u0_col_out_953;
wire [511:0] u0_col_out_954;
wire [511:0] u0_col_out_955;
wire [511:0] u0_col_out_956;
wire [511:0] u0_col_out_957;
wire [511:0] u0_col_out_958;
wire [511:0] u0_col_out_959;
wire [511:0] u0_col_out_960;
wire [511:0] u0_col_out_961;
wire [511:0] u0_col_out_962;
wire [511:0] u0_col_out_963;
wire [511:0] u0_col_out_964;
wire [511:0] u0_col_out_965;
wire [511:0] u0_col_out_966;
wire [511:0] u0_col_out_967;
wire [511:0] u0_col_out_968;
wire [511:0] u0_col_out_969;
wire [511:0] u0_col_out_970;
wire [511:0] u0_col_out_971;
wire [511:0] u0_col_out_972;
wire [511:0] u0_col_out_973;
wire [511:0] u0_col_out_974;
wire [511:0] u0_col_out_975;
wire [511:0] u0_col_out_976;
wire [511:0] u0_col_out_977;
wire [511:0] u0_col_out_978;
wire [511:0] u0_col_out_979;
wire [511:0] u0_col_out_980;
wire [511:0] u0_col_out_981;
wire [511:0] u0_col_out_982;
wire [511:0] u0_col_out_983;
wire [511:0] u0_col_out_984;
wire [511:0] u0_col_out_985;
wire [511:0] u0_col_out_986;
wire [511:0] u0_col_out_987;
wire [511:0] u0_col_out_988;
wire [511:0] u0_col_out_989;
wire [511:0] u0_col_out_990;
wire [511:0] u0_col_out_991;
wire [511:0] u0_col_out_992;
wire [511:0] u0_col_out_993;
wire [511:0] u0_col_out_994;
wire [511:0] u0_col_out_995;
wire [511:0] u0_col_out_996;
wire [511:0] u0_col_out_997;
wire [511:0] u0_col_out_998;
wire [511:0] u0_col_out_999;
wire [511:0] u0_col_out_1000;
wire [511:0] u0_col_out_1001;
wire [511:0] u0_col_out_1002;
wire [511:0] u0_col_out_1003;
wire [511:0] u0_col_out_1004;
wire [511:0] u0_col_out_1005;
wire [511:0] u0_col_out_1006;
wire [511:0] u0_col_out_1007;
wire [511:0] u0_col_out_1008;
wire [511:0] u0_col_out_1009;
wire [511:0] u0_col_out_1010;
wire [511:0] u0_col_out_1011;
wire [511:0] u0_col_out_1012;
wire [511:0] u0_col_out_1013;
wire [511:0] u0_col_out_1014;
wire [511:0] u0_col_out_1015;
wire [511:0] u0_col_out_1016;
wire [511:0] u0_col_out_1017;
wire [511:0] u0_col_out_1018;
wire [511:0] u0_col_out_1019;
wire [511:0] u0_col_out_1020;
wire [511:0] u0_col_out_1021;
wire [511:0] u0_col_out_1022;
wire [511:0] u0_col_out_1023;


msq_half_product_gene u0_msq_half_product_gene
(
    .a(a),
    .sel(sel_hp),

    .col_0(u0_col_out_0),
    .col_1(u0_col_out_1),
    .col_2(u0_col_out_2),
    .col_3(u0_col_out_3),
    .col_4(u0_col_out_4),
    .col_5(u0_col_out_5),
    .col_6(u0_col_out_6),
    .col_7(u0_col_out_7),
    .col_8(u0_col_out_8),
    .col_9(u0_col_out_9),
    .col_10(u0_col_out_10),
    .col_11(u0_col_out_11),
    .col_12(u0_col_out_12),
    .col_13(u0_col_out_13),
    .col_14(u0_col_out_14),
    .col_15(u0_col_out_15),
    .col_16(u0_col_out_16),
    .col_17(u0_col_out_17),
    .col_18(u0_col_out_18),
    .col_19(u0_col_out_19),
    .col_20(u0_col_out_20),
    .col_21(u0_col_out_21),
    .col_22(u0_col_out_22),
    .col_23(u0_col_out_23),
    .col_24(u0_col_out_24),
    .col_25(u0_col_out_25),
    .col_26(u0_col_out_26),
    .col_27(u0_col_out_27),
    .col_28(u0_col_out_28),
    .col_29(u0_col_out_29),
    .col_30(u0_col_out_30),
    .col_31(u0_col_out_31),
    .col_32(u0_col_out_32),
    .col_33(u0_col_out_33),
    .col_34(u0_col_out_34),
    .col_35(u0_col_out_35),
    .col_36(u0_col_out_36),
    .col_37(u0_col_out_37),
    .col_38(u0_col_out_38),
    .col_39(u0_col_out_39),
    .col_40(u0_col_out_40),
    .col_41(u0_col_out_41),
    .col_42(u0_col_out_42),
    .col_43(u0_col_out_43),
    .col_44(u0_col_out_44),
    .col_45(u0_col_out_45),
    .col_46(u0_col_out_46),
    .col_47(u0_col_out_47),
    .col_48(u0_col_out_48),
    .col_49(u0_col_out_49),
    .col_50(u0_col_out_50),
    .col_51(u0_col_out_51),
    .col_52(u0_col_out_52),
    .col_53(u0_col_out_53),
    .col_54(u0_col_out_54),
    .col_55(u0_col_out_55),
    .col_56(u0_col_out_56),
    .col_57(u0_col_out_57),
    .col_58(u0_col_out_58),
    .col_59(u0_col_out_59),
    .col_60(u0_col_out_60),
    .col_61(u0_col_out_61),
    .col_62(u0_col_out_62),
    .col_63(u0_col_out_63),
    .col_64(u0_col_out_64),
    .col_65(u0_col_out_65),
    .col_66(u0_col_out_66),
    .col_67(u0_col_out_67),
    .col_68(u0_col_out_68),
    .col_69(u0_col_out_69),
    .col_70(u0_col_out_70),
    .col_71(u0_col_out_71),
    .col_72(u0_col_out_72),
    .col_73(u0_col_out_73),
    .col_74(u0_col_out_74),
    .col_75(u0_col_out_75),
    .col_76(u0_col_out_76),
    .col_77(u0_col_out_77),
    .col_78(u0_col_out_78),
    .col_79(u0_col_out_79),
    .col_80(u0_col_out_80),
    .col_81(u0_col_out_81),
    .col_82(u0_col_out_82),
    .col_83(u0_col_out_83),
    .col_84(u0_col_out_84),
    .col_85(u0_col_out_85),
    .col_86(u0_col_out_86),
    .col_87(u0_col_out_87),
    .col_88(u0_col_out_88),
    .col_89(u0_col_out_89),
    .col_90(u0_col_out_90),
    .col_91(u0_col_out_91),
    .col_92(u0_col_out_92),
    .col_93(u0_col_out_93),
    .col_94(u0_col_out_94),
    .col_95(u0_col_out_95),
    .col_96(u0_col_out_96),
    .col_97(u0_col_out_97),
    .col_98(u0_col_out_98),
    .col_99(u0_col_out_99),
    .col_100(u0_col_out_100),
    .col_101(u0_col_out_101),
    .col_102(u0_col_out_102),
    .col_103(u0_col_out_103),
    .col_104(u0_col_out_104),
    .col_105(u0_col_out_105),
    .col_106(u0_col_out_106),
    .col_107(u0_col_out_107),
    .col_108(u0_col_out_108),
    .col_109(u0_col_out_109),
    .col_110(u0_col_out_110),
    .col_111(u0_col_out_111),
    .col_112(u0_col_out_112),
    .col_113(u0_col_out_113),
    .col_114(u0_col_out_114),
    .col_115(u0_col_out_115),
    .col_116(u0_col_out_116),
    .col_117(u0_col_out_117),
    .col_118(u0_col_out_118),
    .col_119(u0_col_out_119),
    .col_120(u0_col_out_120),
    .col_121(u0_col_out_121),
    .col_122(u0_col_out_122),
    .col_123(u0_col_out_123),
    .col_124(u0_col_out_124),
    .col_125(u0_col_out_125),
    .col_126(u0_col_out_126),
    .col_127(u0_col_out_127),
    .col_128(u0_col_out_128),
    .col_129(u0_col_out_129),
    .col_130(u0_col_out_130),
    .col_131(u0_col_out_131),
    .col_132(u0_col_out_132),
    .col_133(u0_col_out_133),
    .col_134(u0_col_out_134),
    .col_135(u0_col_out_135),
    .col_136(u0_col_out_136),
    .col_137(u0_col_out_137),
    .col_138(u0_col_out_138),
    .col_139(u0_col_out_139),
    .col_140(u0_col_out_140),
    .col_141(u0_col_out_141),
    .col_142(u0_col_out_142),
    .col_143(u0_col_out_143),
    .col_144(u0_col_out_144),
    .col_145(u0_col_out_145),
    .col_146(u0_col_out_146),
    .col_147(u0_col_out_147),
    .col_148(u0_col_out_148),
    .col_149(u0_col_out_149),
    .col_150(u0_col_out_150),
    .col_151(u0_col_out_151),
    .col_152(u0_col_out_152),
    .col_153(u0_col_out_153),
    .col_154(u0_col_out_154),
    .col_155(u0_col_out_155),
    .col_156(u0_col_out_156),
    .col_157(u0_col_out_157),
    .col_158(u0_col_out_158),
    .col_159(u0_col_out_159),
    .col_160(u0_col_out_160),
    .col_161(u0_col_out_161),
    .col_162(u0_col_out_162),
    .col_163(u0_col_out_163),
    .col_164(u0_col_out_164),
    .col_165(u0_col_out_165),
    .col_166(u0_col_out_166),
    .col_167(u0_col_out_167),
    .col_168(u0_col_out_168),
    .col_169(u0_col_out_169),
    .col_170(u0_col_out_170),
    .col_171(u0_col_out_171),
    .col_172(u0_col_out_172),
    .col_173(u0_col_out_173),
    .col_174(u0_col_out_174),
    .col_175(u0_col_out_175),
    .col_176(u0_col_out_176),
    .col_177(u0_col_out_177),
    .col_178(u0_col_out_178),
    .col_179(u0_col_out_179),
    .col_180(u0_col_out_180),
    .col_181(u0_col_out_181),
    .col_182(u0_col_out_182),
    .col_183(u0_col_out_183),
    .col_184(u0_col_out_184),
    .col_185(u0_col_out_185),
    .col_186(u0_col_out_186),
    .col_187(u0_col_out_187),
    .col_188(u0_col_out_188),
    .col_189(u0_col_out_189),
    .col_190(u0_col_out_190),
    .col_191(u0_col_out_191),
    .col_192(u0_col_out_192),
    .col_193(u0_col_out_193),
    .col_194(u0_col_out_194),
    .col_195(u0_col_out_195),
    .col_196(u0_col_out_196),
    .col_197(u0_col_out_197),
    .col_198(u0_col_out_198),
    .col_199(u0_col_out_199),
    .col_200(u0_col_out_200),
    .col_201(u0_col_out_201),
    .col_202(u0_col_out_202),
    .col_203(u0_col_out_203),
    .col_204(u0_col_out_204),
    .col_205(u0_col_out_205),
    .col_206(u0_col_out_206),
    .col_207(u0_col_out_207),
    .col_208(u0_col_out_208),
    .col_209(u0_col_out_209),
    .col_210(u0_col_out_210),
    .col_211(u0_col_out_211),
    .col_212(u0_col_out_212),
    .col_213(u0_col_out_213),
    .col_214(u0_col_out_214),
    .col_215(u0_col_out_215),
    .col_216(u0_col_out_216),
    .col_217(u0_col_out_217),
    .col_218(u0_col_out_218),
    .col_219(u0_col_out_219),
    .col_220(u0_col_out_220),
    .col_221(u0_col_out_221),
    .col_222(u0_col_out_222),
    .col_223(u0_col_out_223),
    .col_224(u0_col_out_224),
    .col_225(u0_col_out_225),
    .col_226(u0_col_out_226),
    .col_227(u0_col_out_227),
    .col_228(u0_col_out_228),
    .col_229(u0_col_out_229),
    .col_230(u0_col_out_230),
    .col_231(u0_col_out_231),
    .col_232(u0_col_out_232),
    .col_233(u0_col_out_233),
    .col_234(u0_col_out_234),
    .col_235(u0_col_out_235),
    .col_236(u0_col_out_236),
    .col_237(u0_col_out_237),
    .col_238(u0_col_out_238),
    .col_239(u0_col_out_239),
    .col_240(u0_col_out_240),
    .col_241(u0_col_out_241),
    .col_242(u0_col_out_242),
    .col_243(u0_col_out_243),
    .col_244(u0_col_out_244),
    .col_245(u0_col_out_245),
    .col_246(u0_col_out_246),
    .col_247(u0_col_out_247),
    .col_248(u0_col_out_248),
    .col_249(u0_col_out_249),
    .col_250(u0_col_out_250),
    .col_251(u0_col_out_251),
    .col_252(u0_col_out_252),
    .col_253(u0_col_out_253),
    .col_254(u0_col_out_254),
    .col_255(u0_col_out_255),
    .col_256(u0_col_out_256),
    .col_257(u0_col_out_257),
    .col_258(u0_col_out_258),
    .col_259(u0_col_out_259),
    .col_260(u0_col_out_260),
    .col_261(u0_col_out_261),
    .col_262(u0_col_out_262),
    .col_263(u0_col_out_263),
    .col_264(u0_col_out_264),
    .col_265(u0_col_out_265),
    .col_266(u0_col_out_266),
    .col_267(u0_col_out_267),
    .col_268(u0_col_out_268),
    .col_269(u0_col_out_269),
    .col_270(u0_col_out_270),
    .col_271(u0_col_out_271),
    .col_272(u0_col_out_272),
    .col_273(u0_col_out_273),
    .col_274(u0_col_out_274),
    .col_275(u0_col_out_275),
    .col_276(u0_col_out_276),
    .col_277(u0_col_out_277),
    .col_278(u0_col_out_278),
    .col_279(u0_col_out_279),
    .col_280(u0_col_out_280),
    .col_281(u0_col_out_281),
    .col_282(u0_col_out_282),
    .col_283(u0_col_out_283),
    .col_284(u0_col_out_284),
    .col_285(u0_col_out_285),
    .col_286(u0_col_out_286),
    .col_287(u0_col_out_287),
    .col_288(u0_col_out_288),
    .col_289(u0_col_out_289),
    .col_290(u0_col_out_290),
    .col_291(u0_col_out_291),
    .col_292(u0_col_out_292),
    .col_293(u0_col_out_293),
    .col_294(u0_col_out_294),
    .col_295(u0_col_out_295),
    .col_296(u0_col_out_296),
    .col_297(u0_col_out_297),
    .col_298(u0_col_out_298),
    .col_299(u0_col_out_299),
    .col_300(u0_col_out_300),
    .col_301(u0_col_out_301),
    .col_302(u0_col_out_302),
    .col_303(u0_col_out_303),
    .col_304(u0_col_out_304),
    .col_305(u0_col_out_305),
    .col_306(u0_col_out_306),
    .col_307(u0_col_out_307),
    .col_308(u0_col_out_308),
    .col_309(u0_col_out_309),
    .col_310(u0_col_out_310),
    .col_311(u0_col_out_311),
    .col_312(u0_col_out_312),
    .col_313(u0_col_out_313),
    .col_314(u0_col_out_314),
    .col_315(u0_col_out_315),
    .col_316(u0_col_out_316),
    .col_317(u0_col_out_317),
    .col_318(u0_col_out_318),
    .col_319(u0_col_out_319),
    .col_320(u0_col_out_320),
    .col_321(u0_col_out_321),
    .col_322(u0_col_out_322),
    .col_323(u0_col_out_323),
    .col_324(u0_col_out_324),
    .col_325(u0_col_out_325),
    .col_326(u0_col_out_326),
    .col_327(u0_col_out_327),
    .col_328(u0_col_out_328),
    .col_329(u0_col_out_329),
    .col_330(u0_col_out_330),
    .col_331(u0_col_out_331),
    .col_332(u0_col_out_332),
    .col_333(u0_col_out_333),
    .col_334(u0_col_out_334),
    .col_335(u0_col_out_335),
    .col_336(u0_col_out_336),
    .col_337(u0_col_out_337),
    .col_338(u0_col_out_338),
    .col_339(u0_col_out_339),
    .col_340(u0_col_out_340),
    .col_341(u0_col_out_341),
    .col_342(u0_col_out_342),
    .col_343(u0_col_out_343),
    .col_344(u0_col_out_344),
    .col_345(u0_col_out_345),
    .col_346(u0_col_out_346),
    .col_347(u0_col_out_347),
    .col_348(u0_col_out_348),
    .col_349(u0_col_out_349),
    .col_350(u0_col_out_350),
    .col_351(u0_col_out_351),
    .col_352(u0_col_out_352),
    .col_353(u0_col_out_353),
    .col_354(u0_col_out_354),
    .col_355(u0_col_out_355),
    .col_356(u0_col_out_356),
    .col_357(u0_col_out_357),
    .col_358(u0_col_out_358),
    .col_359(u0_col_out_359),
    .col_360(u0_col_out_360),
    .col_361(u0_col_out_361),
    .col_362(u0_col_out_362),
    .col_363(u0_col_out_363),
    .col_364(u0_col_out_364),
    .col_365(u0_col_out_365),
    .col_366(u0_col_out_366),
    .col_367(u0_col_out_367),
    .col_368(u0_col_out_368),
    .col_369(u0_col_out_369),
    .col_370(u0_col_out_370),
    .col_371(u0_col_out_371),
    .col_372(u0_col_out_372),
    .col_373(u0_col_out_373),
    .col_374(u0_col_out_374),
    .col_375(u0_col_out_375),
    .col_376(u0_col_out_376),
    .col_377(u0_col_out_377),
    .col_378(u0_col_out_378),
    .col_379(u0_col_out_379),
    .col_380(u0_col_out_380),
    .col_381(u0_col_out_381),
    .col_382(u0_col_out_382),
    .col_383(u0_col_out_383),
    .col_384(u0_col_out_384),
    .col_385(u0_col_out_385),
    .col_386(u0_col_out_386),
    .col_387(u0_col_out_387),
    .col_388(u0_col_out_388),
    .col_389(u0_col_out_389),
    .col_390(u0_col_out_390),
    .col_391(u0_col_out_391),
    .col_392(u0_col_out_392),
    .col_393(u0_col_out_393),
    .col_394(u0_col_out_394),
    .col_395(u0_col_out_395),
    .col_396(u0_col_out_396),
    .col_397(u0_col_out_397),
    .col_398(u0_col_out_398),
    .col_399(u0_col_out_399),
    .col_400(u0_col_out_400),
    .col_401(u0_col_out_401),
    .col_402(u0_col_out_402),
    .col_403(u0_col_out_403),
    .col_404(u0_col_out_404),
    .col_405(u0_col_out_405),
    .col_406(u0_col_out_406),
    .col_407(u0_col_out_407),
    .col_408(u0_col_out_408),
    .col_409(u0_col_out_409),
    .col_410(u0_col_out_410),
    .col_411(u0_col_out_411),
    .col_412(u0_col_out_412),
    .col_413(u0_col_out_413),
    .col_414(u0_col_out_414),
    .col_415(u0_col_out_415),
    .col_416(u0_col_out_416),
    .col_417(u0_col_out_417),
    .col_418(u0_col_out_418),
    .col_419(u0_col_out_419),
    .col_420(u0_col_out_420),
    .col_421(u0_col_out_421),
    .col_422(u0_col_out_422),
    .col_423(u0_col_out_423),
    .col_424(u0_col_out_424),
    .col_425(u0_col_out_425),
    .col_426(u0_col_out_426),
    .col_427(u0_col_out_427),
    .col_428(u0_col_out_428),
    .col_429(u0_col_out_429),
    .col_430(u0_col_out_430),
    .col_431(u0_col_out_431),
    .col_432(u0_col_out_432),
    .col_433(u0_col_out_433),
    .col_434(u0_col_out_434),
    .col_435(u0_col_out_435),
    .col_436(u0_col_out_436),
    .col_437(u0_col_out_437),
    .col_438(u0_col_out_438),
    .col_439(u0_col_out_439),
    .col_440(u0_col_out_440),
    .col_441(u0_col_out_441),
    .col_442(u0_col_out_442),
    .col_443(u0_col_out_443),
    .col_444(u0_col_out_444),
    .col_445(u0_col_out_445),
    .col_446(u0_col_out_446),
    .col_447(u0_col_out_447),
    .col_448(u0_col_out_448),
    .col_449(u0_col_out_449),
    .col_450(u0_col_out_450),
    .col_451(u0_col_out_451),
    .col_452(u0_col_out_452),
    .col_453(u0_col_out_453),
    .col_454(u0_col_out_454),
    .col_455(u0_col_out_455),
    .col_456(u0_col_out_456),
    .col_457(u0_col_out_457),
    .col_458(u0_col_out_458),
    .col_459(u0_col_out_459),
    .col_460(u0_col_out_460),
    .col_461(u0_col_out_461),
    .col_462(u0_col_out_462),
    .col_463(u0_col_out_463),
    .col_464(u0_col_out_464),
    .col_465(u0_col_out_465),
    .col_466(u0_col_out_466),
    .col_467(u0_col_out_467),
    .col_468(u0_col_out_468),
    .col_469(u0_col_out_469),
    .col_470(u0_col_out_470),
    .col_471(u0_col_out_471),
    .col_472(u0_col_out_472),
    .col_473(u0_col_out_473),
    .col_474(u0_col_out_474),
    .col_475(u0_col_out_475),
    .col_476(u0_col_out_476),
    .col_477(u0_col_out_477),
    .col_478(u0_col_out_478),
    .col_479(u0_col_out_479),
    .col_480(u0_col_out_480),
    .col_481(u0_col_out_481),
    .col_482(u0_col_out_482),
    .col_483(u0_col_out_483),
    .col_484(u0_col_out_484),
    .col_485(u0_col_out_485),
    .col_486(u0_col_out_486),
    .col_487(u0_col_out_487),
    .col_488(u0_col_out_488),
    .col_489(u0_col_out_489),
    .col_490(u0_col_out_490),
    .col_491(u0_col_out_491),
    .col_492(u0_col_out_492),
    .col_493(u0_col_out_493),
    .col_494(u0_col_out_494),
    .col_495(u0_col_out_495),
    .col_496(u0_col_out_496),
    .col_497(u0_col_out_497),
    .col_498(u0_col_out_498),
    .col_499(u0_col_out_499),
    .col_500(u0_col_out_500),
    .col_501(u0_col_out_501),
    .col_502(u0_col_out_502),
    .col_503(u0_col_out_503),
    .col_504(u0_col_out_504),
    .col_505(u0_col_out_505),
    .col_506(u0_col_out_506),
    .col_507(u0_col_out_507),
    .col_508(u0_col_out_508),
    .col_509(u0_col_out_509),
    .col_510(u0_col_out_510),
    .col_511(u0_col_out_511),
    .col_512(u0_col_out_512),
    .col_513(u0_col_out_513),
    .col_514(u0_col_out_514),
    .col_515(u0_col_out_515),
    .col_516(u0_col_out_516),
    .col_517(u0_col_out_517),
    .col_518(u0_col_out_518),
    .col_519(u0_col_out_519),
    .col_520(u0_col_out_520),
    .col_521(u0_col_out_521),
    .col_522(u0_col_out_522),
    .col_523(u0_col_out_523),
    .col_524(u0_col_out_524),
    .col_525(u0_col_out_525),
    .col_526(u0_col_out_526),
    .col_527(u0_col_out_527),
    .col_528(u0_col_out_528),
    .col_529(u0_col_out_529),
    .col_530(u0_col_out_530),
    .col_531(u0_col_out_531),
    .col_532(u0_col_out_532),
    .col_533(u0_col_out_533),
    .col_534(u0_col_out_534),
    .col_535(u0_col_out_535),
    .col_536(u0_col_out_536),
    .col_537(u0_col_out_537),
    .col_538(u0_col_out_538),
    .col_539(u0_col_out_539),
    .col_540(u0_col_out_540),
    .col_541(u0_col_out_541),
    .col_542(u0_col_out_542),
    .col_543(u0_col_out_543),
    .col_544(u0_col_out_544),
    .col_545(u0_col_out_545),
    .col_546(u0_col_out_546),
    .col_547(u0_col_out_547),
    .col_548(u0_col_out_548),
    .col_549(u0_col_out_549),
    .col_550(u0_col_out_550),
    .col_551(u0_col_out_551),
    .col_552(u0_col_out_552),
    .col_553(u0_col_out_553),
    .col_554(u0_col_out_554),
    .col_555(u0_col_out_555),
    .col_556(u0_col_out_556),
    .col_557(u0_col_out_557),
    .col_558(u0_col_out_558),
    .col_559(u0_col_out_559),
    .col_560(u0_col_out_560),
    .col_561(u0_col_out_561),
    .col_562(u0_col_out_562),
    .col_563(u0_col_out_563),
    .col_564(u0_col_out_564),
    .col_565(u0_col_out_565),
    .col_566(u0_col_out_566),
    .col_567(u0_col_out_567),
    .col_568(u0_col_out_568),
    .col_569(u0_col_out_569),
    .col_570(u0_col_out_570),
    .col_571(u0_col_out_571),
    .col_572(u0_col_out_572),
    .col_573(u0_col_out_573),
    .col_574(u0_col_out_574),
    .col_575(u0_col_out_575),
    .col_576(u0_col_out_576),
    .col_577(u0_col_out_577),
    .col_578(u0_col_out_578),
    .col_579(u0_col_out_579),
    .col_580(u0_col_out_580),
    .col_581(u0_col_out_581),
    .col_582(u0_col_out_582),
    .col_583(u0_col_out_583),
    .col_584(u0_col_out_584),
    .col_585(u0_col_out_585),
    .col_586(u0_col_out_586),
    .col_587(u0_col_out_587),
    .col_588(u0_col_out_588),
    .col_589(u0_col_out_589),
    .col_590(u0_col_out_590),
    .col_591(u0_col_out_591),
    .col_592(u0_col_out_592),
    .col_593(u0_col_out_593),
    .col_594(u0_col_out_594),
    .col_595(u0_col_out_595),
    .col_596(u0_col_out_596),
    .col_597(u0_col_out_597),
    .col_598(u0_col_out_598),
    .col_599(u0_col_out_599),
    .col_600(u0_col_out_600),
    .col_601(u0_col_out_601),
    .col_602(u0_col_out_602),
    .col_603(u0_col_out_603),
    .col_604(u0_col_out_604),
    .col_605(u0_col_out_605),
    .col_606(u0_col_out_606),
    .col_607(u0_col_out_607),
    .col_608(u0_col_out_608),
    .col_609(u0_col_out_609),
    .col_610(u0_col_out_610),
    .col_611(u0_col_out_611),
    .col_612(u0_col_out_612),
    .col_613(u0_col_out_613),
    .col_614(u0_col_out_614),
    .col_615(u0_col_out_615),
    .col_616(u0_col_out_616),
    .col_617(u0_col_out_617),
    .col_618(u0_col_out_618),
    .col_619(u0_col_out_619),
    .col_620(u0_col_out_620),
    .col_621(u0_col_out_621),
    .col_622(u0_col_out_622),
    .col_623(u0_col_out_623),
    .col_624(u0_col_out_624),
    .col_625(u0_col_out_625),
    .col_626(u0_col_out_626),
    .col_627(u0_col_out_627),
    .col_628(u0_col_out_628),
    .col_629(u0_col_out_629),
    .col_630(u0_col_out_630),
    .col_631(u0_col_out_631),
    .col_632(u0_col_out_632),
    .col_633(u0_col_out_633),
    .col_634(u0_col_out_634),
    .col_635(u0_col_out_635),
    .col_636(u0_col_out_636),
    .col_637(u0_col_out_637),
    .col_638(u0_col_out_638),
    .col_639(u0_col_out_639),
    .col_640(u0_col_out_640),
    .col_641(u0_col_out_641),
    .col_642(u0_col_out_642),
    .col_643(u0_col_out_643),
    .col_644(u0_col_out_644),
    .col_645(u0_col_out_645),
    .col_646(u0_col_out_646),
    .col_647(u0_col_out_647),
    .col_648(u0_col_out_648),
    .col_649(u0_col_out_649),
    .col_650(u0_col_out_650),
    .col_651(u0_col_out_651),
    .col_652(u0_col_out_652),
    .col_653(u0_col_out_653),
    .col_654(u0_col_out_654),
    .col_655(u0_col_out_655),
    .col_656(u0_col_out_656),
    .col_657(u0_col_out_657),
    .col_658(u0_col_out_658),
    .col_659(u0_col_out_659),
    .col_660(u0_col_out_660),
    .col_661(u0_col_out_661),
    .col_662(u0_col_out_662),
    .col_663(u0_col_out_663),
    .col_664(u0_col_out_664),
    .col_665(u0_col_out_665),
    .col_666(u0_col_out_666),
    .col_667(u0_col_out_667),
    .col_668(u0_col_out_668),
    .col_669(u0_col_out_669),
    .col_670(u0_col_out_670),
    .col_671(u0_col_out_671),
    .col_672(u0_col_out_672),
    .col_673(u0_col_out_673),
    .col_674(u0_col_out_674),
    .col_675(u0_col_out_675),
    .col_676(u0_col_out_676),
    .col_677(u0_col_out_677),
    .col_678(u0_col_out_678),
    .col_679(u0_col_out_679),
    .col_680(u0_col_out_680),
    .col_681(u0_col_out_681),
    .col_682(u0_col_out_682),
    .col_683(u0_col_out_683),
    .col_684(u0_col_out_684),
    .col_685(u0_col_out_685),
    .col_686(u0_col_out_686),
    .col_687(u0_col_out_687),
    .col_688(u0_col_out_688),
    .col_689(u0_col_out_689),
    .col_690(u0_col_out_690),
    .col_691(u0_col_out_691),
    .col_692(u0_col_out_692),
    .col_693(u0_col_out_693),
    .col_694(u0_col_out_694),
    .col_695(u0_col_out_695),
    .col_696(u0_col_out_696),
    .col_697(u0_col_out_697),
    .col_698(u0_col_out_698),
    .col_699(u0_col_out_699),
    .col_700(u0_col_out_700),
    .col_701(u0_col_out_701),
    .col_702(u0_col_out_702),
    .col_703(u0_col_out_703),
    .col_704(u0_col_out_704),
    .col_705(u0_col_out_705),
    .col_706(u0_col_out_706),
    .col_707(u0_col_out_707),
    .col_708(u0_col_out_708),
    .col_709(u0_col_out_709),
    .col_710(u0_col_out_710),
    .col_711(u0_col_out_711),
    .col_712(u0_col_out_712),
    .col_713(u0_col_out_713),
    .col_714(u0_col_out_714),
    .col_715(u0_col_out_715),
    .col_716(u0_col_out_716),
    .col_717(u0_col_out_717),
    .col_718(u0_col_out_718),
    .col_719(u0_col_out_719),
    .col_720(u0_col_out_720),
    .col_721(u0_col_out_721),
    .col_722(u0_col_out_722),
    .col_723(u0_col_out_723),
    .col_724(u0_col_out_724),
    .col_725(u0_col_out_725),
    .col_726(u0_col_out_726),
    .col_727(u0_col_out_727),
    .col_728(u0_col_out_728),
    .col_729(u0_col_out_729),
    .col_730(u0_col_out_730),
    .col_731(u0_col_out_731),
    .col_732(u0_col_out_732),
    .col_733(u0_col_out_733),
    .col_734(u0_col_out_734),
    .col_735(u0_col_out_735),
    .col_736(u0_col_out_736),
    .col_737(u0_col_out_737),
    .col_738(u0_col_out_738),
    .col_739(u0_col_out_739),
    .col_740(u0_col_out_740),
    .col_741(u0_col_out_741),
    .col_742(u0_col_out_742),
    .col_743(u0_col_out_743),
    .col_744(u0_col_out_744),
    .col_745(u0_col_out_745),
    .col_746(u0_col_out_746),
    .col_747(u0_col_out_747),
    .col_748(u0_col_out_748),
    .col_749(u0_col_out_749),
    .col_750(u0_col_out_750),
    .col_751(u0_col_out_751),
    .col_752(u0_col_out_752),
    .col_753(u0_col_out_753),
    .col_754(u0_col_out_754),
    .col_755(u0_col_out_755),
    .col_756(u0_col_out_756),
    .col_757(u0_col_out_757),
    .col_758(u0_col_out_758),
    .col_759(u0_col_out_759),
    .col_760(u0_col_out_760),
    .col_761(u0_col_out_761),
    .col_762(u0_col_out_762),
    .col_763(u0_col_out_763),
    .col_764(u0_col_out_764),
    .col_765(u0_col_out_765),
    .col_766(u0_col_out_766),
    .col_767(u0_col_out_767),
    .col_768(u0_col_out_768),
    .col_769(u0_col_out_769),
    .col_770(u0_col_out_770),
    .col_771(u0_col_out_771),
    .col_772(u0_col_out_772),
    .col_773(u0_col_out_773),
    .col_774(u0_col_out_774),
    .col_775(u0_col_out_775),
    .col_776(u0_col_out_776),
    .col_777(u0_col_out_777),
    .col_778(u0_col_out_778),
    .col_779(u0_col_out_779),
    .col_780(u0_col_out_780),
    .col_781(u0_col_out_781),
    .col_782(u0_col_out_782),
    .col_783(u0_col_out_783),
    .col_784(u0_col_out_784),
    .col_785(u0_col_out_785),
    .col_786(u0_col_out_786),
    .col_787(u0_col_out_787),
    .col_788(u0_col_out_788),
    .col_789(u0_col_out_789),
    .col_790(u0_col_out_790),
    .col_791(u0_col_out_791),
    .col_792(u0_col_out_792),
    .col_793(u0_col_out_793),
    .col_794(u0_col_out_794),
    .col_795(u0_col_out_795),
    .col_796(u0_col_out_796),
    .col_797(u0_col_out_797),
    .col_798(u0_col_out_798),
    .col_799(u0_col_out_799),
    .col_800(u0_col_out_800),
    .col_801(u0_col_out_801),
    .col_802(u0_col_out_802),
    .col_803(u0_col_out_803),
    .col_804(u0_col_out_804),
    .col_805(u0_col_out_805),
    .col_806(u0_col_out_806),
    .col_807(u0_col_out_807),
    .col_808(u0_col_out_808),
    .col_809(u0_col_out_809),
    .col_810(u0_col_out_810),
    .col_811(u0_col_out_811),
    .col_812(u0_col_out_812),
    .col_813(u0_col_out_813),
    .col_814(u0_col_out_814),
    .col_815(u0_col_out_815),
    .col_816(u0_col_out_816),
    .col_817(u0_col_out_817),
    .col_818(u0_col_out_818),
    .col_819(u0_col_out_819),
    .col_820(u0_col_out_820),
    .col_821(u0_col_out_821),
    .col_822(u0_col_out_822),
    .col_823(u0_col_out_823),
    .col_824(u0_col_out_824),
    .col_825(u0_col_out_825),
    .col_826(u0_col_out_826),
    .col_827(u0_col_out_827),
    .col_828(u0_col_out_828),
    .col_829(u0_col_out_829),
    .col_830(u0_col_out_830),
    .col_831(u0_col_out_831),
    .col_832(u0_col_out_832),
    .col_833(u0_col_out_833),
    .col_834(u0_col_out_834),
    .col_835(u0_col_out_835),
    .col_836(u0_col_out_836),
    .col_837(u0_col_out_837),
    .col_838(u0_col_out_838),
    .col_839(u0_col_out_839),
    .col_840(u0_col_out_840),
    .col_841(u0_col_out_841),
    .col_842(u0_col_out_842),
    .col_843(u0_col_out_843),
    .col_844(u0_col_out_844),
    .col_845(u0_col_out_845),
    .col_846(u0_col_out_846),
    .col_847(u0_col_out_847),
    .col_848(u0_col_out_848),
    .col_849(u0_col_out_849),
    .col_850(u0_col_out_850),
    .col_851(u0_col_out_851),
    .col_852(u0_col_out_852),
    .col_853(u0_col_out_853),
    .col_854(u0_col_out_854),
    .col_855(u0_col_out_855),
    .col_856(u0_col_out_856),
    .col_857(u0_col_out_857),
    .col_858(u0_col_out_858),
    .col_859(u0_col_out_859),
    .col_860(u0_col_out_860),
    .col_861(u0_col_out_861),
    .col_862(u0_col_out_862),
    .col_863(u0_col_out_863),
    .col_864(u0_col_out_864),
    .col_865(u0_col_out_865),
    .col_866(u0_col_out_866),
    .col_867(u0_col_out_867),
    .col_868(u0_col_out_868),
    .col_869(u0_col_out_869),
    .col_870(u0_col_out_870),
    .col_871(u0_col_out_871),
    .col_872(u0_col_out_872),
    .col_873(u0_col_out_873),
    .col_874(u0_col_out_874),
    .col_875(u0_col_out_875),
    .col_876(u0_col_out_876),
    .col_877(u0_col_out_877),
    .col_878(u0_col_out_878),
    .col_879(u0_col_out_879),
    .col_880(u0_col_out_880),
    .col_881(u0_col_out_881),
    .col_882(u0_col_out_882),
    .col_883(u0_col_out_883),
    .col_884(u0_col_out_884),
    .col_885(u0_col_out_885),
    .col_886(u0_col_out_886),
    .col_887(u0_col_out_887),
    .col_888(u0_col_out_888),
    .col_889(u0_col_out_889),
    .col_890(u0_col_out_890),
    .col_891(u0_col_out_891),
    .col_892(u0_col_out_892),
    .col_893(u0_col_out_893),
    .col_894(u0_col_out_894),
    .col_895(u0_col_out_895),
    .col_896(u0_col_out_896),
    .col_897(u0_col_out_897),
    .col_898(u0_col_out_898),
    .col_899(u0_col_out_899),
    .col_900(u0_col_out_900),
    .col_901(u0_col_out_901),
    .col_902(u0_col_out_902),
    .col_903(u0_col_out_903),
    .col_904(u0_col_out_904),
    .col_905(u0_col_out_905),
    .col_906(u0_col_out_906),
    .col_907(u0_col_out_907),
    .col_908(u0_col_out_908),
    .col_909(u0_col_out_909),
    .col_910(u0_col_out_910),
    .col_911(u0_col_out_911),
    .col_912(u0_col_out_912),
    .col_913(u0_col_out_913),
    .col_914(u0_col_out_914),
    .col_915(u0_col_out_915),
    .col_916(u0_col_out_916),
    .col_917(u0_col_out_917),
    .col_918(u0_col_out_918),
    .col_919(u0_col_out_919),
    .col_920(u0_col_out_920),
    .col_921(u0_col_out_921),
    .col_922(u0_col_out_922),
    .col_923(u0_col_out_923),
    .col_924(u0_col_out_924),
    .col_925(u0_col_out_925),
    .col_926(u0_col_out_926),
    .col_927(u0_col_out_927),
    .col_928(u0_col_out_928),
    .col_929(u0_col_out_929),
    .col_930(u0_col_out_930),
    .col_931(u0_col_out_931),
    .col_932(u0_col_out_932),
    .col_933(u0_col_out_933),
    .col_934(u0_col_out_934),
    .col_935(u0_col_out_935),
    .col_936(u0_col_out_936),
    .col_937(u0_col_out_937),
    .col_938(u0_col_out_938),
    .col_939(u0_col_out_939),
    .col_940(u0_col_out_940),
    .col_941(u0_col_out_941),
    .col_942(u0_col_out_942),
    .col_943(u0_col_out_943),
    .col_944(u0_col_out_944),
    .col_945(u0_col_out_945),
    .col_946(u0_col_out_946),
    .col_947(u0_col_out_947),
    .col_948(u0_col_out_948),
    .col_949(u0_col_out_949),
    .col_950(u0_col_out_950),
    .col_951(u0_col_out_951),
    .col_952(u0_col_out_952),
    .col_953(u0_col_out_953),
    .col_954(u0_col_out_954),
    .col_955(u0_col_out_955),
    .col_956(u0_col_out_956),
    .col_957(u0_col_out_957),
    .col_958(u0_col_out_958),
    .col_959(u0_col_out_959),
    .col_960(u0_col_out_960),
    .col_961(u0_col_out_961),
    .col_962(u0_col_out_962),
    .col_963(u0_col_out_963),
    .col_964(u0_col_out_964),
    .col_965(u0_col_out_965),
    .col_966(u0_col_out_966),
    .col_967(u0_col_out_967),
    .col_968(u0_col_out_968),
    .col_969(u0_col_out_969),
    .col_970(u0_col_out_970),
    .col_971(u0_col_out_971),
    .col_972(u0_col_out_972),
    .col_973(u0_col_out_973),
    .col_974(u0_col_out_974),
    .col_975(u0_col_out_975),
    .col_976(u0_col_out_976),
    .col_977(u0_col_out_977),
    .col_978(u0_col_out_978),
    .col_979(u0_col_out_979),
    .col_980(u0_col_out_980),
    .col_981(u0_col_out_981),
    .col_982(u0_col_out_982),
    .col_983(u0_col_out_983),
    .col_984(u0_col_out_984),
    .col_985(u0_col_out_985),
    .col_986(u0_col_out_986),
    .col_987(u0_col_out_987),
    .col_988(u0_col_out_988),
    .col_989(u0_col_out_989),
    .col_990(u0_col_out_990),
    .col_991(u0_col_out_991),
    .col_992(u0_col_out_992),
    .col_993(u0_col_out_993),
    .col_994(u0_col_out_994),
    .col_995(u0_col_out_995),
    .col_996(u0_col_out_996),
    .col_997(u0_col_out_997),
    .col_998(u0_col_out_998),
    .col_999(u0_col_out_999),
    .col_1000(u0_col_out_1000),
    .col_1001(u0_col_out_1001),
    .col_1002(u0_col_out_1002),
    .col_1003(u0_col_out_1003),
    .col_1004(u0_col_out_1004),
    .col_1005(u0_col_out_1005),
    .col_1006(u0_col_out_1006),
    .col_1007(u0_col_out_1007),
    .col_1008(u0_col_out_1008),
    .col_1009(u0_col_out_1009),
    .col_1010(u0_col_out_1010),
    .col_1011(u0_col_out_1011),
    .col_1012(u0_col_out_1012),
    .col_1013(u0_col_out_1013),
    .col_1014(u0_col_out_1014),
    .col_1015(u0_col_out_1015),
    .col_1016(u0_col_out_1016),
    .col_1017(u0_col_out_1017),
    .col_1018(u0_col_out_1018),
    .col_1019(u0_col_out_1019),
    .col_1020(u0_col_out_1020),
    .col_1021(u0_col_out_1021),
    .col_1022(u0_col_out_1022),
    .col_1023(u0_col_out_1023)
);




// first_reduction_data Outputs
wire  [511:0]  u1_col_out_0;
wire  [511:0]  u1_col_out_1;
wire  [511:0]  u1_col_out_2;
wire  [511:0]  u1_col_out_3;
wire  [511:0]  u1_col_out_4;
wire  [511:0]  u1_col_out_5;
wire  [511:0]  u1_col_out_6;
wire  [511:0]  u1_col_out_7;
wire  [511:0]  u1_col_out_8;
wire  [511:0]  u1_col_out_9;
wire  [511:0]  u1_col_out_10;
wire  [511:0]  u1_col_out_11;
wire  [511:0]  u1_col_out_12;
wire  [511:0]  u1_col_out_13;
wire  [511:0]  u1_col_out_14;
wire  [511:0]  u1_col_out_15;
wire  [511:0]  u1_col_out_16;
wire  [511:0]  u1_col_out_17;
wire  [511:0]  u1_col_out_18;
wire  [511:0]  u1_col_out_19;
wire  [511:0]  u1_col_out_20;
wire  [511:0]  u1_col_out_21;
wire  [511:0]  u1_col_out_22;
wire  [511:0]  u1_col_out_23;
wire  [511:0]  u1_col_out_24;
wire  [511:0]  u1_col_out_25;
wire  [511:0]  u1_col_out_26;
wire  [511:0]  u1_col_out_27;
wire  [511:0]  u1_col_out_28;
wire  [511:0]  u1_col_out_29;
wire  [511:0]  u1_col_out_30;
wire  [511:0]  u1_col_out_31;
wire  [511:0]  u1_col_out_32;
wire  [511:0]  u1_col_out_33;
wire  [511:0]  u1_col_out_34;
wire  [511:0]  u1_col_out_35;
wire  [511:0]  u1_col_out_36;
wire  [511:0]  u1_col_out_37;
wire  [511:0]  u1_col_out_38;
wire  [511:0]  u1_col_out_39;
wire  [511:0]  u1_col_out_40;
wire  [511:0]  u1_col_out_41;
wire  [511:0]  u1_col_out_42;
wire  [511:0]  u1_col_out_43;
wire  [511:0]  u1_col_out_44;
wire  [511:0]  u1_col_out_45;
wire  [511:0]  u1_col_out_46;
wire  [511:0]  u1_col_out_47;
wire  [511:0]  u1_col_out_48;
wire  [511:0]  u1_col_out_49;
wire  [511:0]  u1_col_out_50;
wire  [511:0]  u1_col_out_51;
wire  [511:0]  u1_col_out_52;
wire  [511:0]  u1_col_out_53;
wire  [511:0]  u1_col_out_54;
wire  [511:0]  u1_col_out_55;
wire  [511:0]  u1_col_out_56;
wire  [511:0]  u1_col_out_57;
wire  [511:0]  u1_col_out_58;
wire  [511:0]  u1_col_out_59;
wire  [511:0]  u1_col_out_60;
wire  [511:0]  u1_col_out_61;
wire  [511:0]  u1_col_out_62;
wire  [511:0]  u1_col_out_63;
wire  [511:0]  u1_col_out_64;
wire  [511:0]  u1_col_out_65;
wire  [511:0]  u1_col_out_66;
wire  [511:0]  u1_col_out_67;
wire  [511:0]  u1_col_out_68;
wire  [511:0]  u1_col_out_69;
wire  [511:0]  u1_col_out_70;
wire  [511:0]  u1_col_out_71;
wire  [511:0]  u1_col_out_72;
wire  [511:0]  u1_col_out_73;
wire  [511:0]  u1_col_out_74;
wire  [511:0]  u1_col_out_75;
wire  [511:0]  u1_col_out_76;
wire  [511:0]  u1_col_out_77;
wire  [511:0]  u1_col_out_78;
wire  [511:0]  u1_col_out_79;
wire  [511:0]  u1_col_out_80;
wire  [511:0]  u1_col_out_81;
wire  [511:0]  u1_col_out_82;
wire  [511:0]  u1_col_out_83;
wire  [511:0]  u1_col_out_84;
wire  [511:0]  u1_col_out_85;
wire  [511:0]  u1_col_out_86;
wire  [511:0]  u1_col_out_87;
wire  [511:0]  u1_col_out_88;
wire  [511:0]  u1_col_out_89;
wire  [511:0]  u1_col_out_90;
wire  [511:0]  u1_col_out_91;
wire  [511:0]  u1_col_out_92;
wire  [511:0]  u1_col_out_93;
wire  [511:0]  u1_col_out_94;
wire  [511:0]  u1_col_out_95;
wire  [511:0]  u1_col_out_96;
wire  [511:0]  u1_col_out_97;
wire  [511:0]  u1_col_out_98;
wire  [511:0]  u1_col_out_99;
wire  [511:0]  u1_col_out_100;
wire  [511:0]  u1_col_out_101;
wire  [511:0]  u1_col_out_102;
wire  [511:0]  u1_col_out_103;
wire  [511:0]  u1_col_out_104;
wire  [511:0]  u1_col_out_105;
wire  [511:0]  u1_col_out_106;
wire  [511:0]  u1_col_out_107;
wire  [511:0]  u1_col_out_108;
wire  [511:0]  u1_col_out_109;
wire  [511:0]  u1_col_out_110;
wire  [511:0]  u1_col_out_111;
wire  [511:0]  u1_col_out_112;
wire  [511:0]  u1_col_out_113;
wire  [511:0]  u1_col_out_114;
wire  [511:0]  u1_col_out_115;
wire  [511:0]  u1_col_out_116;
wire  [511:0]  u1_col_out_117;
wire  [511:0]  u1_col_out_118;
wire  [511:0]  u1_col_out_119;
wire  [511:0]  u1_col_out_120;
wire  [511:0]  u1_col_out_121;
wire  [511:0]  u1_col_out_122;
wire  [511:0]  u1_col_out_123;
wire  [511:0]  u1_col_out_124;
wire  [511:0]  u1_col_out_125;
wire  [511:0]  u1_col_out_126;
wire  [511:0]  u1_col_out_127;
wire  [511:0]  u1_col_out_128;
wire  [511:0]  u1_col_out_129;
wire  [511:0]  u1_col_out_130;
wire  [511:0]  u1_col_out_131;
wire  [511:0]  u1_col_out_132;
wire  [511:0]  u1_col_out_133;
wire  [511:0]  u1_col_out_134;
wire  [511:0]  u1_col_out_135;
wire  [511:0]  u1_col_out_136;
wire  [511:0]  u1_col_out_137;
wire  [511:0]  u1_col_out_138;
wire  [511:0]  u1_col_out_139;
wire  [511:0]  u1_col_out_140;
wire  [511:0]  u1_col_out_141;
wire  [511:0]  u1_col_out_142;
wire  [511:0]  u1_col_out_143;
wire  [511:0]  u1_col_out_144;
wire  [511:0]  u1_col_out_145;
wire  [511:0]  u1_col_out_146;
wire  [511:0]  u1_col_out_147;
wire  [511:0]  u1_col_out_148;
wire  [511:0]  u1_col_out_149;
wire  [511:0]  u1_col_out_150;
wire  [511:0]  u1_col_out_151;
wire  [511:0]  u1_col_out_152;
wire  [511:0]  u1_col_out_153;
wire  [511:0]  u1_col_out_154;
wire  [511:0]  u1_col_out_155;
wire  [511:0]  u1_col_out_156;
wire  [511:0]  u1_col_out_157;
wire  [511:0]  u1_col_out_158;
wire  [511:0]  u1_col_out_159;
wire  [511:0]  u1_col_out_160;
wire  [511:0]  u1_col_out_161;
wire  [511:0]  u1_col_out_162;
wire  [511:0]  u1_col_out_163;
wire  [511:0]  u1_col_out_164;
wire  [511:0]  u1_col_out_165;
wire  [511:0]  u1_col_out_166;
wire  [511:0]  u1_col_out_167;
wire  [511:0]  u1_col_out_168;
wire  [511:0]  u1_col_out_169;
wire  [511:0]  u1_col_out_170;
wire  [511:0]  u1_col_out_171;
wire  [511:0]  u1_col_out_172;
wire  [511:0]  u1_col_out_173;
wire  [511:0]  u1_col_out_174;
wire  [511:0]  u1_col_out_175;
wire  [511:0]  u1_col_out_176;
wire  [511:0]  u1_col_out_177;
wire  [511:0]  u1_col_out_178;
wire  [511:0]  u1_col_out_179;
wire  [511:0]  u1_col_out_180;
wire  [511:0]  u1_col_out_181;
wire  [511:0]  u1_col_out_182;
wire  [511:0]  u1_col_out_183;
wire  [511:0]  u1_col_out_184;
wire  [511:0]  u1_col_out_185;
wire  [511:0]  u1_col_out_186;
wire  [511:0]  u1_col_out_187;
wire  [511:0]  u1_col_out_188;
wire  [511:0]  u1_col_out_189;
wire  [511:0]  u1_col_out_190;
wire  [511:0]  u1_col_out_191;
wire  [511:0]  u1_col_out_192;
wire  [511:0]  u1_col_out_193;
wire  [511:0]  u1_col_out_194;
wire  [511:0]  u1_col_out_195;
wire  [511:0]  u1_col_out_196;
wire  [511:0]  u1_col_out_197;
wire  [511:0]  u1_col_out_198;
wire  [511:0]  u1_col_out_199;
wire  [511:0]  u1_col_out_200;
wire  [511:0]  u1_col_out_201;
wire  [511:0]  u1_col_out_202;
wire  [511:0]  u1_col_out_203;
wire  [511:0]  u1_col_out_204;
wire  [511:0]  u1_col_out_205;
wire  [511:0]  u1_col_out_206;
wire  [511:0]  u1_col_out_207;
wire  [511:0]  u1_col_out_208;
wire  [511:0]  u1_col_out_209;
wire  [511:0]  u1_col_out_210;
wire  [511:0]  u1_col_out_211;
wire  [511:0]  u1_col_out_212;
wire  [511:0]  u1_col_out_213;
wire  [511:0]  u1_col_out_214;
wire  [511:0]  u1_col_out_215;
wire  [511:0]  u1_col_out_216;
wire  [511:0]  u1_col_out_217;
wire  [511:0]  u1_col_out_218;
wire  [511:0]  u1_col_out_219;
wire  [511:0]  u1_col_out_220;
wire  [511:0]  u1_col_out_221;
wire  [511:0]  u1_col_out_222;
wire  [511:0]  u1_col_out_223;
wire  [511:0]  u1_col_out_224;
wire  [511:0]  u1_col_out_225;
wire  [511:0]  u1_col_out_226;
wire  [511:0]  u1_col_out_227;
wire  [511:0]  u1_col_out_228;
wire  [511:0]  u1_col_out_229;
wire  [511:0]  u1_col_out_230;
wire  [511:0]  u1_col_out_231;
wire  [511:0]  u1_col_out_232;
wire  [511:0]  u1_col_out_233;
wire  [511:0]  u1_col_out_234;
wire  [511:0]  u1_col_out_235;
wire  [511:0]  u1_col_out_236;
wire  [511:0]  u1_col_out_237;
wire  [511:0]  u1_col_out_238;
wire  [511:0]  u1_col_out_239;
wire  [511:0]  u1_col_out_240;
wire  [511:0]  u1_col_out_241;
wire  [511:0]  u1_col_out_242;
wire  [511:0]  u1_col_out_243;
wire  [511:0]  u1_col_out_244;
wire  [511:0]  u1_col_out_245;
wire  [511:0]  u1_col_out_246;
wire  [511:0]  u1_col_out_247;
wire  [511:0]  u1_col_out_248;
wire  [511:0]  u1_col_out_249;
wire  [511:0]  u1_col_out_250;
wire  [511:0]  u1_col_out_251;
wire  [511:0]  u1_col_out_252;
wire  [511:0]  u1_col_out_253;
wire  [511:0]  u1_col_out_254;
wire  [511:0]  u1_col_out_255;
wire  [511:0]  u1_col_out_256;
wire  [511:0]  u1_col_out_257;
wire  [511:0]  u1_col_out_258;
wire  [511:0]  u1_col_out_259;
wire  [511:0]  u1_col_out_260;
wire  [511:0]  u1_col_out_261;
wire  [511:0]  u1_col_out_262;
wire  [511:0]  u1_col_out_263;
wire  [511:0]  u1_col_out_264;
wire  [511:0]  u1_col_out_265;
wire  [511:0]  u1_col_out_266;
wire  [511:0]  u1_col_out_267;
wire  [511:0]  u1_col_out_268;
wire  [511:0]  u1_col_out_269;
wire  [511:0]  u1_col_out_270;
wire  [511:0]  u1_col_out_271;
wire  [511:0]  u1_col_out_272;
wire  [511:0]  u1_col_out_273;
wire  [511:0]  u1_col_out_274;
wire  [511:0]  u1_col_out_275;
wire  [511:0]  u1_col_out_276;
wire  [511:0]  u1_col_out_277;
wire  [511:0]  u1_col_out_278;
wire  [511:0]  u1_col_out_279;
wire  [511:0]  u1_col_out_280;
wire  [511:0]  u1_col_out_281;
wire  [511:0]  u1_col_out_282;
wire  [511:0]  u1_col_out_283;
wire  [511:0]  u1_col_out_284;
wire  [511:0]  u1_col_out_285;
wire  [511:0]  u1_col_out_286;
wire  [511:0]  u1_col_out_287;
wire  [511:0]  u1_col_out_288;
wire  [511:0]  u1_col_out_289;
wire  [511:0]  u1_col_out_290;
wire  [511:0]  u1_col_out_291;
wire  [511:0]  u1_col_out_292;
wire  [511:0]  u1_col_out_293;
wire  [511:0]  u1_col_out_294;
wire  [511:0]  u1_col_out_295;
wire  [511:0]  u1_col_out_296;
wire  [511:0]  u1_col_out_297;
wire  [511:0]  u1_col_out_298;
wire  [511:0]  u1_col_out_299;
wire  [511:0]  u1_col_out_300;
wire  [511:0]  u1_col_out_301;
wire  [511:0]  u1_col_out_302;
wire  [511:0]  u1_col_out_303;
wire  [511:0]  u1_col_out_304;
wire  [511:0]  u1_col_out_305;
wire  [511:0]  u1_col_out_306;
wire  [511:0]  u1_col_out_307;
wire  [511:0]  u1_col_out_308;
wire  [511:0]  u1_col_out_309;
wire  [511:0]  u1_col_out_310;
wire  [511:0]  u1_col_out_311;
wire  [511:0]  u1_col_out_312;
wire  [511:0]  u1_col_out_313;
wire  [511:0]  u1_col_out_314;
wire  [511:0]  u1_col_out_315;
wire  [511:0]  u1_col_out_316;
wire  [511:0]  u1_col_out_317;
wire  [511:0]  u1_col_out_318;
wire  [511:0]  u1_col_out_319;
wire  [511:0]  u1_col_out_320;
wire  [511:0]  u1_col_out_321;
wire  [511:0]  u1_col_out_322;
wire  [511:0]  u1_col_out_323;
wire  [511:0]  u1_col_out_324;
wire  [511:0]  u1_col_out_325;
wire  [511:0]  u1_col_out_326;
wire  [511:0]  u1_col_out_327;
wire  [511:0]  u1_col_out_328;
wire  [511:0]  u1_col_out_329;
wire  [511:0]  u1_col_out_330;
wire  [511:0]  u1_col_out_331;
wire  [511:0]  u1_col_out_332;
wire  [511:0]  u1_col_out_333;
wire  [511:0]  u1_col_out_334;
wire  [511:0]  u1_col_out_335;
wire  [511:0]  u1_col_out_336;
wire  [511:0]  u1_col_out_337;
wire  [511:0]  u1_col_out_338;
wire  [511:0]  u1_col_out_339;
wire  [511:0]  u1_col_out_340;
wire  [511:0]  u1_col_out_341;
wire  [511:0]  u1_col_out_342;
wire  [511:0]  u1_col_out_343;
wire  [511:0]  u1_col_out_344;
wire  [511:0]  u1_col_out_345;
wire  [511:0]  u1_col_out_346;
wire  [511:0]  u1_col_out_347;
wire  [511:0]  u1_col_out_348;
wire  [511:0]  u1_col_out_349;
wire  [511:0]  u1_col_out_350;
wire  [511:0]  u1_col_out_351;
wire  [511:0]  u1_col_out_352;
wire  [511:0]  u1_col_out_353;
wire  [511:0]  u1_col_out_354;
wire  [511:0]  u1_col_out_355;
wire  [511:0]  u1_col_out_356;
wire  [511:0]  u1_col_out_357;
wire  [511:0]  u1_col_out_358;
wire  [511:0]  u1_col_out_359;
wire  [511:0]  u1_col_out_360;
wire  [511:0]  u1_col_out_361;
wire  [511:0]  u1_col_out_362;
wire  [511:0]  u1_col_out_363;
wire  [511:0]  u1_col_out_364;
wire  [511:0]  u1_col_out_365;
wire  [511:0]  u1_col_out_366;
wire  [511:0]  u1_col_out_367;
wire  [511:0]  u1_col_out_368;
wire  [511:0]  u1_col_out_369;
wire  [511:0]  u1_col_out_370;
wire  [511:0]  u1_col_out_371;
wire  [511:0]  u1_col_out_372;
wire  [511:0]  u1_col_out_373;
wire  [511:0]  u1_col_out_374;
wire  [511:0]  u1_col_out_375;
wire  [511:0]  u1_col_out_376;
wire  [511:0]  u1_col_out_377;
wire  [511:0]  u1_col_out_378;
wire  [511:0]  u1_col_out_379;
wire  [511:0]  u1_col_out_380;
wire  [511:0]  u1_col_out_381;
wire  [511:0]  u1_col_out_382;
wire  [511:0]  u1_col_out_383;
wire  [511:0]  u1_col_out_384;
wire  [511:0]  u1_col_out_385;
wire  [511:0]  u1_col_out_386;
wire  [511:0]  u1_col_out_387;
wire  [511:0]  u1_col_out_388;
wire  [511:0]  u1_col_out_389;
wire  [511:0]  u1_col_out_390;
wire  [511:0]  u1_col_out_391;
wire  [511:0]  u1_col_out_392;
wire  [511:0]  u1_col_out_393;
wire  [511:0]  u1_col_out_394;
wire  [511:0]  u1_col_out_395;
wire  [511:0]  u1_col_out_396;
wire  [511:0]  u1_col_out_397;
wire  [511:0]  u1_col_out_398;
wire  [511:0]  u1_col_out_399;
wire  [511:0]  u1_col_out_400;
wire  [511:0]  u1_col_out_401;
wire  [511:0]  u1_col_out_402;
wire  [511:0]  u1_col_out_403;
wire  [511:0]  u1_col_out_404;
wire  [511:0]  u1_col_out_405;
wire  [511:0]  u1_col_out_406;
wire  [511:0]  u1_col_out_407;
wire  [511:0]  u1_col_out_408;
wire  [511:0]  u1_col_out_409;
wire  [511:0]  u1_col_out_410;
wire  [511:0]  u1_col_out_411;
wire  [511:0]  u1_col_out_412;
wire  [511:0]  u1_col_out_413;
wire  [511:0]  u1_col_out_414;
wire  [511:0]  u1_col_out_415;
wire  [511:0]  u1_col_out_416;
wire  [511:0]  u1_col_out_417;
wire  [511:0]  u1_col_out_418;
wire  [511:0]  u1_col_out_419;
wire  [511:0]  u1_col_out_420;
wire  [511:0]  u1_col_out_421;
wire  [511:0]  u1_col_out_422;
wire  [511:0]  u1_col_out_423;
wire  [511:0]  u1_col_out_424;
wire  [511:0]  u1_col_out_425;
wire  [511:0]  u1_col_out_426;
wire  [511:0]  u1_col_out_427;
wire  [511:0]  u1_col_out_428;
wire  [511:0]  u1_col_out_429;
wire  [511:0]  u1_col_out_430;
wire  [511:0]  u1_col_out_431;
wire  [511:0]  u1_col_out_432;
wire  [511:0]  u1_col_out_433;
wire  [511:0]  u1_col_out_434;
wire  [511:0]  u1_col_out_435;
wire  [511:0]  u1_col_out_436;
wire  [511:0]  u1_col_out_437;
wire  [511:0]  u1_col_out_438;
wire  [511:0]  u1_col_out_439;
wire  [511:0]  u1_col_out_440;
wire  [511:0]  u1_col_out_441;
wire  [511:0]  u1_col_out_442;
wire  [511:0]  u1_col_out_443;
wire  [511:0]  u1_col_out_444;
wire  [511:0]  u1_col_out_445;
wire  [511:0]  u1_col_out_446;
wire  [511:0]  u1_col_out_447;
wire  [511:0]  u1_col_out_448;
wire  [511:0]  u1_col_out_449;
wire  [511:0]  u1_col_out_450;
wire  [511:0]  u1_col_out_451;
wire  [511:0]  u1_col_out_452;
wire  [511:0]  u1_col_out_453;
wire  [511:0]  u1_col_out_454;
wire  [511:0]  u1_col_out_455;
wire  [511:0]  u1_col_out_456;
wire  [511:0]  u1_col_out_457;
wire  [511:0]  u1_col_out_458;
wire  [511:0]  u1_col_out_459;
wire  [511:0]  u1_col_out_460;
wire  [511:0]  u1_col_out_461;
wire  [511:0]  u1_col_out_462;
wire  [511:0]  u1_col_out_463;
wire  [511:0]  u1_col_out_464;
wire  [511:0]  u1_col_out_465;
wire  [511:0]  u1_col_out_466;
wire  [511:0]  u1_col_out_467;
wire  [511:0]  u1_col_out_468;
wire  [511:0]  u1_col_out_469;
wire  [511:0]  u1_col_out_470;
wire  [511:0]  u1_col_out_471;
wire  [511:0]  u1_col_out_472;
wire  [511:0]  u1_col_out_473;
wire  [511:0]  u1_col_out_474;
wire  [511:0]  u1_col_out_475;
wire  [511:0]  u1_col_out_476;
wire  [511:0]  u1_col_out_477;
wire  [511:0]  u1_col_out_478;
wire  [511:0]  u1_col_out_479;
wire  [511:0]  u1_col_out_480;
wire  [511:0]  u1_col_out_481;
wire  [511:0]  u1_col_out_482;
wire  [511:0]  u1_col_out_483;
wire  [511:0]  u1_col_out_484;
wire  [511:0]  u1_col_out_485;
wire  [511:0]  u1_col_out_486;
wire  [511:0]  u1_col_out_487;
wire  [511:0]  u1_col_out_488;
wire  [511:0]  u1_col_out_489;
wire  [511:0]  u1_col_out_490;
wire  [511:0]  u1_col_out_491;
wire  [511:0]  u1_col_out_492;
wire  [511:0]  u1_col_out_493;
wire  [511:0]  u1_col_out_494;
wire  [511:0]  u1_col_out_495;
wire  [511:0]  u1_col_out_496;
wire  [511:0]  u1_col_out_497;
wire  [511:0]  u1_col_out_498;
wire  [511:0]  u1_col_out_499;
wire  [511:0]  u1_col_out_500;
wire  [511:0]  u1_col_out_501;
wire  [511:0]  u1_col_out_502;
wire  [511:0]  u1_col_out_503;
wire  [511:0]  u1_col_out_504;
wire  [511:0]  u1_col_out_505;
wire  [511:0]  u1_col_out_506;
wire  [511:0]  u1_col_out_507;
wire  [511:0]  u1_col_out_508;
wire  [511:0]  u1_col_out_509;
wire  [511:0]  u1_col_out_510;
wire  [511:0]  u1_col_out_511;
wire  [511:0]  u1_col_out_512;
wire  [511:0]  u1_col_out_513;
wire  [511:0]  u1_col_out_514;
wire  [511:0]  u1_col_out_515;
wire  [511:0]  u1_col_out_516;
wire  [511:0]  u1_col_out_517;
wire  [511:0]  u1_col_out_518;
wire  [511:0]  u1_col_out_519;
wire  [511:0]  u1_col_out_520;
wire  [511:0]  u1_col_out_521;
wire  [511:0]  u1_col_out_522;
wire  [511:0]  u1_col_out_523;
wire  [511:0]  u1_col_out_524;
wire  [511:0]  u1_col_out_525;
wire  [511:0]  u1_col_out_526;
wire  [511:0]  u1_col_out_527;
wire  [511:0]  u1_col_out_528;
wire  [511:0]  u1_col_out_529;
wire  [511:0]  u1_col_out_530;
wire  [511:0]  u1_col_out_531;
wire  [511:0]  u1_col_out_532;
wire  [511:0]  u1_col_out_533;
wire  [511:0]  u1_col_out_534;
wire  [511:0]  u1_col_out_535;
wire  [511:0]  u1_col_out_536;
wire  [511:0]  u1_col_out_537;
wire  [511:0]  u1_col_out_538;
wire  [511:0]  u1_col_out_539;
wire  [511:0]  u1_col_out_540;
wire  [511:0]  u1_col_out_541;
wire  [511:0]  u1_col_out_542;
wire  [511:0]  u1_col_out_543;
wire  [511:0]  u1_col_out_544;
wire  [511:0]  u1_col_out_545;
wire  [511:0]  u1_col_out_546;
wire  [511:0]  u1_col_out_547;
wire  [511:0]  u1_col_out_548;
wire  [511:0]  u1_col_out_549;
wire  [511:0]  u1_col_out_550;
wire  [511:0]  u1_col_out_551;
wire  [511:0]  u1_col_out_552;
wire  [511:0]  u1_col_out_553;
wire  [511:0]  u1_col_out_554;
wire  [511:0]  u1_col_out_555;
wire  [511:0]  u1_col_out_556;
wire  [511:0]  u1_col_out_557;
wire  [511:0]  u1_col_out_558;
wire  [511:0]  u1_col_out_559;
wire  [511:0]  u1_col_out_560;
wire  [511:0]  u1_col_out_561;
wire  [511:0]  u1_col_out_562;
wire  [511:0]  u1_col_out_563;
wire  [511:0]  u1_col_out_564;
wire  [511:0]  u1_col_out_565;
wire  [511:0]  u1_col_out_566;
wire  [511:0]  u1_col_out_567;
wire  [511:0]  u1_col_out_568;
wire  [511:0]  u1_col_out_569;
wire  [511:0]  u1_col_out_570;
wire  [511:0]  u1_col_out_571;
wire  [511:0]  u1_col_out_572;
wire  [511:0]  u1_col_out_573;
wire  [511:0]  u1_col_out_574;
wire  [511:0]  u1_col_out_575;
wire  [511:0]  u1_col_out_576;
wire  [511:0]  u1_col_out_577;
wire  [511:0]  u1_col_out_578;
wire  [511:0]  u1_col_out_579;
wire  [511:0]  u1_col_out_580;
wire  [511:0]  u1_col_out_581;
wire  [511:0]  u1_col_out_582;
wire  [511:0]  u1_col_out_583;
wire  [511:0]  u1_col_out_584;
wire  [511:0]  u1_col_out_585;
wire  [511:0]  u1_col_out_586;
wire  [511:0]  u1_col_out_587;
wire  [511:0]  u1_col_out_588;
wire  [511:0]  u1_col_out_589;
wire  [511:0]  u1_col_out_590;
wire  [511:0]  u1_col_out_591;
wire  [511:0]  u1_col_out_592;
wire  [511:0]  u1_col_out_593;
wire  [511:0]  u1_col_out_594;
wire  [511:0]  u1_col_out_595;
wire  [511:0]  u1_col_out_596;
wire  [511:0]  u1_col_out_597;
wire  [511:0]  u1_col_out_598;
wire  [511:0]  u1_col_out_599;
wire  [511:0]  u1_col_out_600;
wire  [511:0]  u1_col_out_601;
wire  [511:0]  u1_col_out_602;
wire  [511:0]  u1_col_out_603;
wire  [511:0]  u1_col_out_604;
wire  [511:0]  u1_col_out_605;
wire  [511:0]  u1_col_out_606;
wire  [511:0]  u1_col_out_607;
wire  [511:0]  u1_col_out_608;
wire  [511:0]  u1_col_out_609;
wire  [511:0]  u1_col_out_610;
wire  [511:0]  u1_col_out_611;
wire  [511:0]  u1_col_out_612;
wire  [511:0]  u1_col_out_613;
wire  [511:0]  u1_col_out_614;
wire  [511:0]  u1_col_out_615;
wire  [511:0]  u1_col_out_616;
wire  [511:0]  u1_col_out_617;
wire  [511:0]  u1_col_out_618;
wire  [511:0]  u1_col_out_619;
wire  [511:0]  u1_col_out_620;
wire  [511:0]  u1_col_out_621;
wire  [511:0]  u1_col_out_622;
wire  [511:0]  u1_col_out_623;
wire  [511:0]  u1_col_out_624;
wire  [511:0]  u1_col_out_625;
wire  [511:0]  u1_col_out_626;
wire  [511:0]  u1_col_out_627;
wire  [511:0]  u1_col_out_628;
wire  [511:0]  u1_col_out_629;
wire  [511:0]  u1_col_out_630;
wire  [511:0]  u1_col_out_631;
wire  [511:0]  u1_col_out_632;
wire  [511:0]  u1_col_out_633;
wire  [511:0]  u1_col_out_634;
wire  [511:0]  u1_col_out_635;
wire  [511:0]  u1_col_out_636;
wire  [511:0]  u1_col_out_637;
wire  [511:0]  u1_col_out_638;
wire  [511:0]  u1_col_out_639;
wire  [511:0]  u1_col_out_640;
wire  [511:0]  u1_col_out_641;
wire  [511:0]  u1_col_out_642;
wire  [511:0]  u1_col_out_643;
wire  [511:0]  u1_col_out_644;
wire  [511:0]  u1_col_out_645;
wire  [511:0]  u1_col_out_646;
wire  [511:0]  u1_col_out_647;
wire  [511:0]  u1_col_out_648;
wire  [511:0]  u1_col_out_649;
wire  [511:0]  u1_col_out_650;
wire  [511:0]  u1_col_out_651;
wire  [511:0]  u1_col_out_652;
wire  [511:0]  u1_col_out_653;
wire  [511:0]  u1_col_out_654;
wire  [511:0]  u1_col_out_655;
wire  [511:0]  u1_col_out_656;
wire  [511:0]  u1_col_out_657;
wire  [511:0]  u1_col_out_658;
wire  [511:0]  u1_col_out_659;
wire  [511:0]  u1_col_out_660;
wire  [511:0]  u1_col_out_661;
wire  [511:0]  u1_col_out_662;
wire  [511:0]  u1_col_out_663;
wire  [511:0]  u1_col_out_664;
wire  [511:0]  u1_col_out_665;
wire  [511:0]  u1_col_out_666;
wire  [511:0]  u1_col_out_667;
wire  [511:0]  u1_col_out_668;
wire  [511:0]  u1_col_out_669;
wire  [511:0]  u1_col_out_670;
wire  [511:0]  u1_col_out_671;
wire  [511:0]  u1_col_out_672;
wire  [511:0]  u1_col_out_673;
wire  [511:0]  u1_col_out_674;
wire  [511:0]  u1_col_out_675;
wire  [511:0]  u1_col_out_676;
wire  [511:0]  u1_col_out_677;
wire  [511:0]  u1_col_out_678;
wire  [511:0]  u1_col_out_679;
wire  [511:0]  u1_col_out_680;
wire  [511:0]  u1_col_out_681;
wire  [511:0]  u1_col_out_682;
wire  [511:0]  u1_col_out_683;
wire  [511:0]  u1_col_out_684;
wire  [511:0]  u1_col_out_685;
wire  [511:0]  u1_col_out_686;
wire  [511:0]  u1_col_out_687;
wire  [511:0]  u1_col_out_688;
wire  [511:0]  u1_col_out_689;
wire  [511:0]  u1_col_out_690;
wire  [511:0]  u1_col_out_691;
wire  [511:0]  u1_col_out_692;
wire  [511:0]  u1_col_out_693;
wire  [511:0]  u1_col_out_694;
wire  [511:0]  u1_col_out_695;
wire  [511:0]  u1_col_out_696;
wire  [511:0]  u1_col_out_697;
wire  [511:0]  u1_col_out_698;
wire  [511:0]  u1_col_out_699;
wire  [511:0]  u1_col_out_700;
wire  [511:0]  u1_col_out_701;
wire  [511:0]  u1_col_out_702;
wire  [511:0]  u1_col_out_703;
wire  [511:0]  u1_col_out_704;
wire  [511:0]  u1_col_out_705;
wire  [511:0]  u1_col_out_706;
wire  [511:0]  u1_col_out_707;
wire  [511:0]  u1_col_out_708;
wire  [511:0]  u1_col_out_709;
wire  [511:0]  u1_col_out_710;
wire  [511:0]  u1_col_out_711;
wire  [511:0]  u1_col_out_712;
wire  [511:0]  u1_col_out_713;
wire  [511:0]  u1_col_out_714;
wire  [511:0]  u1_col_out_715;
wire  [511:0]  u1_col_out_716;
wire  [511:0]  u1_col_out_717;
wire  [511:0]  u1_col_out_718;
wire  [511:0]  u1_col_out_719;
wire  [511:0]  u1_col_out_720;
wire  [511:0]  u1_col_out_721;
wire  [511:0]  u1_col_out_722;
wire  [511:0]  u1_col_out_723;
wire  [511:0]  u1_col_out_724;
wire  [511:0]  u1_col_out_725;
wire  [511:0]  u1_col_out_726;
wire  [511:0]  u1_col_out_727;
wire  [511:0]  u1_col_out_728;
wire  [511:0]  u1_col_out_729;
wire  [511:0]  u1_col_out_730;
wire  [511:0]  u1_col_out_731;
wire  [511:0]  u1_col_out_732;
wire  [511:0]  u1_col_out_733;
wire  [511:0]  u1_col_out_734;
wire  [511:0]  u1_col_out_735;
wire  [511:0]  u1_col_out_736;
wire  [511:0]  u1_col_out_737;
wire  [511:0]  u1_col_out_738;
wire  [511:0]  u1_col_out_739;
wire  [511:0]  u1_col_out_740;
wire  [511:0]  u1_col_out_741;
wire  [511:0]  u1_col_out_742;
wire  [511:0]  u1_col_out_743;
wire  [511:0]  u1_col_out_744;
wire  [511:0]  u1_col_out_745;
wire  [511:0]  u1_col_out_746;
wire  [511:0]  u1_col_out_747;
wire  [511:0]  u1_col_out_748;
wire  [511:0]  u1_col_out_749;
wire  [511:0]  u1_col_out_750;
wire  [511:0]  u1_col_out_751;
wire  [511:0]  u1_col_out_752;
wire  [511:0]  u1_col_out_753;
wire  [511:0]  u1_col_out_754;
wire  [511:0]  u1_col_out_755;
wire  [511:0]  u1_col_out_756;
wire  [511:0]  u1_col_out_757;
wire  [511:0]  u1_col_out_758;
wire  [511:0]  u1_col_out_759;
wire  [511:0]  u1_col_out_760;
wire  [511:0]  u1_col_out_761;
wire  [511:0]  u1_col_out_762;
wire  [511:0]  u1_col_out_763;
wire  [511:0]  u1_col_out_764;
wire  [511:0]  u1_col_out_765;
wire  [511:0]  u1_col_out_766;
wire  [511:0]  u1_col_out_767;
wire  [511:0]  u1_col_out_768;
wire  [511:0]  u1_col_out_769;
wire  [511:0]  u1_col_out_770;
wire  [511:0]  u1_col_out_771;
wire  [511:0]  u1_col_out_772;
wire  [511:0]  u1_col_out_773;
wire  [511:0]  u1_col_out_774;
wire  [511:0]  u1_col_out_775;
wire  [511:0]  u1_col_out_776;
wire  [511:0]  u1_col_out_777;
wire  [511:0]  u1_col_out_778;
wire  [511:0]  u1_col_out_779;
wire  [511:0]  u1_col_out_780;
wire  [511:0]  u1_col_out_781;
wire  [511:0]  u1_col_out_782;
wire  [511:0]  u1_col_out_783;
wire  [511:0]  u1_col_out_784;
wire  [511:0]  u1_col_out_785;
wire  [511:0]  u1_col_out_786;
wire  [511:0]  u1_col_out_787;
wire  [511:0]  u1_col_out_788;
wire  [511:0]  u1_col_out_789;
wire  [511:0]  u1_col_out_790;
wire  [511:0]  u1_col_out_791;
wire  [511:0]  u1_col_out_792;
wire  [511:0]  u1_col_out_793;
wire  [511:0]  u1_col_out_794;
wire  [511:0]  u1_col_out_795;
wire  [511:0]  u1_col_out_796;
wire  [511:0]  u1_col_out_797;
wire  [511:0]  u1_col_out_798;
wire  [511:0]  u1_col_out_799;
wire  [511:0]  u1_col_out_800;
wire  [511:0]  u1_col_out_801;
wire  [511:0]  u1_col_out_802;
wire  [511:0]  u1_col_out_803;
wire  [511:0]  u1_col_out_804;
wire  [511:0]  u1_col_out_805;
wire  [511:0]  u1_col_out_806;
wire  [511:0]  u1_col_out_807;
wire  [511:0]  u1_col_out_808;
wire  [511:0]  u1_col_out_809;
wire  [511:0]  u1_col_out_810;
wire  [511:0]  u1_col_out_811;
wire  [511:0]  u1_col_out_812;
wire  [511:0]  u1_col_out_813;
wire  [511:0]  u1_col_out_814;
wire  [511:0]  u1_col_out_815;
wire  [511:0]  u1_col_out_816;
wire  [511:0]  u1_col_out_817;
wire  [511:0]  u1_col_out_818;
wire  [511:0]  u1_col_out_819;
wire  [511:0]  u1_col_out_820;
wire  [511:0]  u1_col_out_821;
wire  [511:0]  u1_col_out_822;
wire  [511:0]  u1_col_out_823;
wire  [511:0]  u1_col_out_824;
wire  [511:0]  u1_col_out_825;
wire  [511:0]  u1_col_out_826;
wire  [511:0]  u1_col_out_827;
wire  [511:0]  u1_col_out_828;
wire  [511:0]  u1_col_out_829;
wire  [511:0]  u1_col_out_830;
wire  [511:0]  u1_col_out_831;
wire  [511:0]  u1_col_out_832;
wire  [511:0]  u1_col_out_833;
wire  [511:0]  u1_col_out_834;
wire  [511:0]  u1_col_out_835;
wire  [511:0]  u1_col_out_836;
wire  [511:0]  u1_col_out_837;
wire  [511:0]  u1_col_out_838;
wire  [511:0]  u1_col_out_839;
wire  [511:0]  u1_col_out_840;
wire  [511:0]  u1_col_out_841;
wire  [511:0]  u1_col_out_842;
wire  [511:0]  u1_col_out_843;
wire  [511:0]  u1_col_out_844;
wire  [511:0]  u1_col_out_845;
wire  [511:0]  u1_col_out_846;
wire  [511:0]  u1_col_out_847;
wire  [511:0]  u1_col_out_848;
wire  [511:0]  u1_col_out_849;
wire  [511:0]  u1_col_out_850;
wire  [511:0]  u1_col_out_851;
wire  [511:0]  u1_col_out_852;
wire  [511:0]  u1_col_out_853;
wire  [511:0]  u1_col_out_854;
wire  [511:0]  u1_col_out_855;
wire  [511:0]  u1_col_out_856;
wire  [511:0]  u1_col_out_857;
wire  [511:0]  u1_col_out_858;
wire  [511:0]  u1_col_out_859;
wire  [511:0]  u1_col_out_860;
wire  [511:0]  u1_col_out_861;
wire  [511:0]  u1_col_out_862;
wire  [511:0]  u1_col_out_863;
wire  [511:0]  u1_col_out_864;
wire  [511:0]  u1_col_out_865;
wire  [511:0]  u1_col_out_866;
wire  [511:0]  u1_col_out_867;
wire  [511:0]  u1_col_out_868;
wire  [511:0]  u1_col_out_869;
wire  [511:0]  u1_col_out_870;
wire  [511:0]  u1_col_out_871;
wire  [511:0]  u1_col_out_872;
wire  [511:0]  u1_col_out_873;
wire  [511:0]  u1_col_out_874;
wire  [511:0]  u1_col_out_875;
wire  [511:0]  u1_col_out_876;
wire  [511:0]  u1_col_out_877;
wire  [511:0]  u1_col_out_878;
wire  [511:0]  u1_col_out_879;
wire  [511:0]  u1_col_out_880;
wire  [511:0]  u1_col_out_881;
wire  [511:0]  u1_col_out_882;
wire  [511:0]  u1_col_out_883;
wire  [511:0]  u1_col_out_884;
wire  [511:0]  u1_col_out_885;
wire  [511:0]  u1_col_out_886;
wire  [511:0]  u1_col_out_887;
wire  [511:0]  u1_col_out_888;
wire  [511:0]  u1_col_out_889;
wire  [511:0]  u1_col_out_890;
wire  [511:0]  u1_col_out_891;
wire  [511:0]  u1_col_out_892;
wire  [511:0]  u1_col_out_893;
wire  [511:0]  u1_col_out_894;
wire  [511:0]  u1_col_out_895;
wire  [511:0]  u1_col_out_896;
wire  [511:0]  u1_col_out_897;
wire  [511:0]  u1_col_out_898;
wire  [511:0]  u1_col_out_899;
wire  [511:0]  u1_col_out_900;
wire  [511:0]  u1_col_out_901;
wire  [511:0]  u1_col_out_902;
wire  [511:0]  u1_col_out_903;
wire  [511:0]  u1_col_out_904;
wire  [511:0]  u1_col_out_905;
wire  [511:0]  u1_col_out_906;
wire  [511:0]  u1_col_out_907;
wire  [511:0]  u1_col_out_908;
wire  [511:0]  u1_col_out_909;
wire  [511:0]  u1_col_out_910;
wire  [511:0]  u1_col_out_911;
wire  [511:0]  u1_col_out_912;
wire  [511:0]  u1_col_out_913;
wire  [511:0]  u1_col_out_914;
wire  [511:0]  u1_col_out_915;
wire  [511:0]  u1_col_out_916;
wire  [511:0]  u1_col_out_917;
wire  [511:0]  u1_col_out_918;
wire  [511:0]  u1_col_out_919;
wire  [511:0]  u1_col_out_920;
wire  [511:0]  u1_col_out_921;
wire  [511:0]  u1_col_out_922;
wire  [511:0]  u1_col_out_923;
wire  [511:0]  u1_col_out_924;
wire  [511:0]  u1_col_out_925;
wire  [511:0]  u1_col_out_926;
wire  [511:0]  u1_col_out_927;
wire  [511:0]  u1_col_out_928;
wire  [511:0]  u1_col_out_929;
wire  [511:0]  u1_col_out_930;
wire  [511:0]  u1_col_out_931;
wire  [511:0]  u1_col_out_932;
wire  [511:0]  u1_col_out_933;
wire  [511:0]  u1_col_out_934;
wire  [511:0]  u1_col_out_935;
wire  [511:0]  u1_col_out_936;
wire  [511:0]  u1_col_out_937;
wire  [511:0]  u1_col_out_938;
wire  [511:0]  u1_col_out_939;
wire  [511:0]  u1_col_out_940;
wire  [511:0]  u1_col_out_941;
wire  [511:0]  u1_col_out_942;
wire  [511:0]  u1_col_out_943;
wire  [511:0]  u1_col_out_944;
wire  [511:0]  u1_col_out_945;
wire  [511:0]  u1_col_out_946;
wire  [511:0]  u1_col_out_947;
wire  [511:0]  u1_col_out_948;
wire  [511:0]  u1_col_out_949;
wire  [511:0]  u1_col_out_950;
wire  [511:0]  u1_col_out_951;
wire  [511:0]  u1_col_out_952;
wire  [511:0]  u1_col_out_953;
wire  [511:0]  u1_col_out_954;
wire  [511:0]  u1_col_out_955;
wire  [511:0]  u1_col_out_956;
wire  [511:0]  u1_col_out_957;
wire  [511:0]  u1_col_out_958;
wire  [511:0]  u1_col_out_959;
wire  [511:0]  u1_col_out_960;
wire  [511:0]  u1_col_out_961;
wire  [511:0]  u1_col_out_962;
wire  [511:0]  u1_col_out_963;
wire  [511:0]  u1_col_out_964;
wire  [511:0]  u1_col_out_965;
wire  [511:0]  u1_col_out_966;
wire  [511:0]  u1_col_out_967;
wire  [511:0]  u1_col_out_968;
wire  [511:0]  u1_col_out_969;
wire  [511:0]  u1_col_out_970;
wire  [511:0]  u1_col_out_971;
wire  [511:0]  u1_col_out_972;
wire  [511:0]  u1_col_out_973;
wire  [511:0]  u1_col_out_974;
wire  [511:0]  u1_col_out_975;
wire  [511:0]  u1_col_out_976;
wire  [511:0]  u1_col_out_977;
wire  [511:0]  u1_col_out_978;
wire  [511:0]  u1_col_out_979;
wire  [511:0]  u1_col_out_980;
wire  [511:0]  u1_col_out_981;
wire  [511:0]  u1_col_out_982;
wire  [511:0]  u1_col_out_983;
wire  [511:0]  u1_col_out_984;
wire  [511:0]  u1_col_out_985;
wire  [511:0]  u1_col_out_986;
wire  [511:0]  u1_col_out_987;
wire  [511:0]  u1_col_out_988;
wire  [511:0]  u1_col_out_989;
wire  [511:0]  u1_col_out_990;
wire  [511:0]  u1_col_out_991;
wire  [511:0]  u1_col_out_992;
wire  [511:0]  u1_col_out_993;
wire  [511:0]  u1_col_out_994;
wire  [511:0]  u1_col_out_995;
wire  [511:0]  u1_col_out_996;
wire  [511:0]  u1_col_out_997;
wire  [511:0]  u1_col_out_998;
wire  [511:0]  u1_col_out_999;
wire  [511:0]  u1_col_out_1000;
wire  [511:0]  u1_col_out_1001;
wire  [511:0]  u1_col_out_1002;
wire  [511:0]  u1_col_out_1003;
wire  [511:0]  u1_col_out_1004;
wire  [511:0]  u1_col_out_1005;
wire  [511:0]  u1_col_out_1006;
wire  [511:0]  u1_col_out_1007;
wire  [511:0]  u1_col_out_1008;
wire  [511:0]  u1_col_out_1009;
wire  [511:0]  u1_col_out_1010;
wire  [511:0]  u1_col_out_1011;
wire  [511:0]  u1_col_out_1012;
wire  [511:0]  u1_col_out_1013;
wire  [511:0]  u1_col_out_1014;
wire  [511:0]  u1_col_out_1015;
wire  [511:0]  u1_col_out_1016;
wire  [511:0]  u1_col_out_1017;
wire  [511:0]  u1_col_out_1018;
wire  [511:0]  u1_col_out_1019;
wire  [511:0]  u1_col_out_1020;
wire  [511:0]  u1_col_out_1021;
wire  [511:0]  u1_col_out_1022;
wire  [511:0]  u1_col_out_1023;

first_reduction_data  u1_first_reduction_data (
    .partial_product_high0   ( partial_product_high0   ),
    .partial_product_high1   ( partial_product_high1   ),
    .partial_product_low0    ( partial_product_low0    ),
    .partial_product_low1    ( partial_product_low1    ),

    .col_out_0               ( u1_col_out_0               ),
    .col_out_1               ( u1_col_out_1               ),
    .col_out_2               ( u1_col_out_2               ),
    .col_out_3               ( u1_col_out_3               ),
    .col_out_4               ( u1_col_out_4               ),
    .col_out_5               ( u1_col_out_5               ),
    .col_out_6               ( u1_col_out_6               ),
    .col_out_7               ( u1_col_out_7               ),
    .col_out_8               ( u1_col_out_8               ),
    .col_out_9               ( u1_col_out_9               ),
    .col_out_10              ( u1_col_out_10              ),
    .col_out_11              ( u1_col_out_11              ),
    .col_out_12              ( u1_col_out_12              ),
    .col_out_13              ( u1_col_out_13              ),
    .col_out_14              ( u1_col_out_14              ),
    .col_out_15              ( u1_col_out_15              ),
    .col_out_16              ( u1_col_out_16              ),
    .col_out_17              ( u1_col_out_17              ),
    .col_out_18              ( u1_col_out_18              ),
    .col_out_19              ( u1_col_out_19              ),
    .col_out_20              ( u1_col_out_20              ),
    .col_out_21              ( u1_col_out_21              ),
    .col_out_22              ( u1_col_out_22              ),
    .col_out_23              ( u1_col_out_23              ),
    .col_out_24              ( u1_col_out_24              ),
    .col_out_25              ( u1_col_out_25              ),
    .col_out_26              ( u1_col_out_26              ),
    .col_out_27              ( u1_col_out_27              ),
    .col_out_28              ( u1_col_out_28              ),
    .col_out_29              ( u1_col_out_29              ),
    .col_out_30              ( u1_col_out_30              ),
    .col_out_31              ( u1_col_out_31              ),
    .col_out_32              ( u1_col_out_32              ),
    .col_out_33              ( u1_col_out_33              ),
    .col_out_34              ( u1_col_out_34              ),
    .col_out_35              ( u1_col_out_35              ),
    .col_out_36              ( u1_col_out_36              ),
    .col_out_37              ( u1_col_out_37              ),
    .col_out_38              ( u1_col_out_38              ),
    .col_out_39              ( u1_col_out_39              ),
    .col_out_40              ( u1_col_out_40              ),
    .col_out_41              ( u1_col_out_41              ),
    .col_out_42              ( u1_col_out_42              ),
    .col_out_43              ( u1_col_out_43              ),
    .col_out_44              ( u1_col_out_44              ),
    .col_out_45              ( u1_col_out_45              ),
    .col_out_46              ( u1_col_out_46              ),
    .col_out_47              ( u1_col_out_47              ),
    .col_out_48              ( u1_col_out_48              ),
    .col_out_49              ( u1_col_out_49              ),
    .col_out_50              ( u1_col_out_50              ),
    .col_out_51              ( u1_col_out_51              ),
    .col_out_52              ( u1_col_out_52              ),
    .col_out_53              ( u1_col_out_53              ),
    .col_out_54              ( u1_col_out_54              ),
    .col_out_55              ( u1_col_out_55              ),
    .col_out_56              ( u1_col_out_56              ),
    .col_out_57              ( u1_col_out_57              ),
    .col_out_58              ( u1_col_out_58              ),
    .col_out_59              ( u1_col_out_59              ),
    .col_out_60              ( u1_col_out_60              ),
    .col_out_61              ( u1_col_out_61              ),
    .col_out_62              ( u1_col_out_62              ),
    .col_out_63              ( u1_col_out_63              ),
    .col_out_64              ( u1_col_out_64              ),
    .col_out_65              ( u1_col_out_65              ),
    .col_out_66              ( u1_col_out_66              ),
    .col_out_67              ( u1_col_out_67              ),
    .col_out_68              ( u1_col_out_68              ),
    .col_out_69              ( u1_col_out_69              ),
    .col_out_70              ( u1_col_out_70              ),
    .col_out_71              ( u1_col_out_71              ),
    .col_out_72              ( u1_col_out_72              ),
    .col_out_73              ( u1_col_out_73              ),
    .col_out_74              ( u1_col_out_74              ),
    .col_out_75              ( u1_col_out_75              ),
    .col_out_76              ( u1_col_out_76              ),
    .col_out_77              ( u1_col_out_77              ),
    .col_out_78              ( u1_col_out_78              ),
    .col_out_79              ( u1_col_out_79              ),
    .col_out_80              ( u1_col_out_80              ),
    .col_out_81              ( u1_col_out_81              ),
    .col_out_82              ( u1_col_out_82              ),
    .col_out_83              ( u1_col_out_83              ),
    .col_out_84              ( u1_col_out_84              ),
    .col_out_85              ( u1_col_out_85              ),
    .col_out_86              ( u1_col_out_86              ),
    .col_out_87              ( u1_col_out_87              ),
    .col_out_88              ( u1_col_out_88              ),
    .col_out_89              ( u1_col_out_89              ),
    .col_out_90              ( u1_col_out_90              ),
    .col_out_91              ( u1_col_out_91              ),
    .col_out_92              ( u1_col_out_92              ),
    .col_out_93              ( u1_col_out_93              ),
    .col_out_94              ( u1_col_out_94              ),
    .col_out_95              ( u1_col_out_95              ),
    .col_out_96              ( u1_col_out_96              ),
    .col_out_97              ( u1_col_out_97              ),
    .col_out_98              ( u1_col_out_98              ),
    .col_out_99              ( u1_col_out_99              ),
    .col_out_100             ( u1_col_out_100             ),
    .col_out_101             ( u1_col_out_101             ),
    .col_out_102             ( u1_col_out_102             ),
    .col_out_103             ( u1_col_out_103             ),
    .col_out_104             ( u1_col_out_104             ),
    .col_out_105             ( u1_col_out_105             ),
    .col_out_106             ( u1_col_out_106             ),
    .col_out_107             ( u1_col_out_107             ),
    .col_out_108             ( u1_col_out_108             ),
    .col_out_109             ( u1_col_out_109             ),
    .col_out_110             ( u1_col_out_110             ),
    .col_out_111             ( u1_col_out_111             ),
    .col_out_112             ( u1_col_out_112             ),
    .col_out_113             ( u1_col_out_113             ),
    .col_out_114             ( u1_col_out_114             ),
    .col_out_115             ( u1_col_out_115             ),
    .col_out_116             ( u1_col_out_116             ),
    .col_out_117             ( u1_col_out_117             ),
    .col_out_118             ( u1_col_out_118             ),
    .col_out_119             ( u1_col_out_119             ),
    .col_out_120             ( u1_col_out_120             ),
    .col_out_121             ( u1_col_out_121             ),
    .col_out_122             ( u1_col_out_122             ),
    .col_out_123             ( u1_col_out_123             ),
    .col_out_124             ( u1_col_out_124             ),
    .col_out_125             ( u1_col_out_125             ),
    .col_out_126             ( u1_col_out_126             ),
    .col_out_127             ( u1_col_out_127             ),
    .col_out_128             ( u1_col_out_128             ),
    .col_out_129             ( u1_col_out_129             ),
    .col_out_130             ( u1_col_out_130             ),
    .col_out_131             ( u1_col_out_131             ),
    .col_out_132             ( u1_col_out_132             ),
    .col_out_133             ( u1_col_out_133             ),
    .col_out_134             ( u1_col_out_134             ),
    .col_out_135             ( u1_col_out_135             ),
    .col_out_136             ( u1_col_out_136             ),
    .col_out_137             ( u1_col_out_137             ),
    .col_out_138             ( u1_col_out_138             ),
    .col_out_139             ( u1_col_out_139             ),
    .col_out_140             ( u1_col_out_140             ),
    .col_out_141             ( u1_col_out_141             ),
    .col_out_142             ( u1_col_out_142             ),
    .col_out_143             ( u1_col_out_143             ),
    .col_out_144             ( u1_col_out_144             ),
    .col_out_145             ( u1_col_out_145             ),
    .col_out_146             ( u1_col_out_146             ),
    .col_out_147             ( u1_col_out_147             ),
    .col_out_148             ( u1_col_out_148             ),
    .col_out_149             ( u1_col_out_149             ),
    .col_out_150             ( u1_col_out_150             ),
    .col_out_151             ( u1_col_out_151             ),
    .col_out_152             ( u1_col_out_152             ),
    .col_out_153             ( u1_col_out_153             ),
    .col_out_154             ( u1_col_out_154             ),
    .col_out_155             ( u1_col_out_155             ),
    .col_out_156             ( u1_col_out_156             ),
    .col_out_157             ( u1_col_out_157             ),
    .col_out_158             ( u1_col_out_158             ),
    .col_out_159             ( u1_col_out_159             ),
    .col_out_160             ( u1_col_out_160             ),
    .col_out_161             ( u1_col_out_161             ),
    .col_out_162             ( u1_col_out_162             ),
    .col_out_163             ( u1_col_out_163             ),
    .col_out_164             ( u1_col_out_164             ),
    .col_out_165             ( u1_col_out_165             ),
    .col_out_166             ( u1_col_out_166             ),
    .col_out_167             ( u1_col_out_167             ),
    .col_out_168             ( u1_col_out_168             ),
    .col_out_169             ( u1_col_out_169             ),
    .col_out_170             ( u1_col_out_170             ),
    .col_out_171             ( u1_col_out_171             ),
    .col_out_172             ( u1_col_out_172             ),
    .col_out_173             ( u1_col_out_173             ),
    .col_out_174             ( u1_col_out_174             ),
    .col_out_175             ( u1_col_out_175             ),
    .col_out_176             ( u1_col_out_176             ),
    .col_out_177             ( u1_col_out_177             ),
    .col_out_178             ( u1_col_out_178             ),
    .col_out_179             ( u1_col_out_179             ),
    .col_out_180             ( u1_col_out_180             ),
    .col_out_181             ( u1_col_out_181             ),
    .col_out_182             ( u1_col_out_182             ),
    .col_out_183             ( u1_col_out_183             ),
    .col_out_184             ( u1_col_out_184             ),
    .col_out_185             ( u1_col_out_185             ),
    .col_out_186             ( u1_col_out_186             ),
    .col_out_187             ( u1_col_out_187             ),
    .col_out_188             ( u1_col_out_188             ),
    .col_out_189             ( u1_col_out_189             ),
    .col_out_190             ( u1_col_out_190             ),
    .col_out_191             ( u1_col_out_191             ),
    .col_out_192             ( u1_col_out_192             ),
    .col_out_193             ( u1_col_out_193             ),
    .col_out_194             ( u1_col_out_194             ),
    .col_out_195             ( u1_col_out_195             ),
    .col_out_196             ( u1_col_out_196             ),
    .col_out_197             ( u1_col_out_197             ),
    .col_out_198             ( u1_col_out_198             ),
    .col_out_199             ( u1_col_out_199             ),
    .col_out_200             ( u1_col_out_200             ),
    .col_out_201             ( u1_col_out_201             ),
    .col_out_202             ( u1_col_out_202             ),
    .col_out_203             ( u1_col_out_203             ),
    .col_out_204             ( u1_col_out_204             ),
    .col_out_205             ( u1_col_out_205             ),
    .col_out_206             ( u1_col_out_206             ),
    .col_out_207             ( u1_col_out_207             ),
    .col_out_208             ( u1_col_out_208             ),
    .col_out_209             ( u1_col_out_209             ),
    .col_out_210             ( u1_col_out_210             ),
    .col_out_211             ( u1_col_out_211             ),
    .col_out_212             ( u1_col_out_212             ),
    .col_out_213             ( u1_col_out_213             ),
    .col_out_214             ( u1_col_out_214             ),
    .col_out_215             ( u1_col_out_215             ),
    .col_out_216             ( u1_col_out_216             ),
    .col_out_217             ( u1_col_out_217             ),
    .col_out_218             ( u1_col_out_218             ),
    .col_out_219             ( u1_col_out_219             ),
    .col_out_220             ( u1_col_out_220             ),
    .col_out_221             ( u1_col_out_221             ),
    .col_out_222             ( u1_col_out_222             ),
    .col_out_223             ( u1_col_out_223             ),
    .col_out_224             ( u1_col_out_224             ),
    .col_out_225             ( u1_col_out_225             ),
    .col_out_226             ( u1_col_out_226             ),
    .col_out_227             ( u1_col_out_227             ),
    .col_out_228             ( u1_col_out_228             ),
    .col_out_229             ( u1_col_out_229             ),
    .col_out_230             ( u1_col_out_230             ),
    .col_out_231             ( u1_col_out_231             ),
    .col_out_232             ( u1_col_out_232             ),
    .col_out_233             ( u1_col_out_233             ),
    .col_out_234             ( u1_col_out_234             ),
    .col_out_235             ( u1_col_out_235             ),
    .col_out_236             ( u1_col_out_236             ),
    .col_out_237             ( u1_col_out_237             ),
    .col_out_238             ( u1_col_out_238             ),
    .col_out_239             ( u1_col_out_239             ),
    .col_out_240             ( u1_col_out_240             ),
    .col_out_241             ( u1_col_out_241             ),
    .col_out_242             ( u1_col_out_242             ),
    .col_out_243             ( u1_col_out_243             ),
    .col_out_244             ( u1_col_out_244             ),
    .col_out_245             ( u1_col_out_245             ),
    .col_out_246             ( u1_col_out_246             ),
    .col_out_247             ( u1_col_out_247             ),
    .col_out_248             ( u1_col_out_248             ),
    .col_out_249             ( u1_col_out_249             ),
    .col_out_250             ( u1_col_out_250             ),
    .col_out_251             ( u1_col_out_251             ),
    .col_out_252             ( u1_col_out_252             ),
    .col_out_253             ( u1_col_out_253             ),
    .col_out_254             ( u1_col_out_254             ),
    .col_out_255             ( u1_col_out_255             ),
    .col_out_256             ( u1_col_out_256             ),
    .col_out_257             ( u1_col_out_257             ),
    .col_out_258             ( u1_col_out_258             ),
    .col_out_259             ( u1_col_out_259             ),
    .col_out_260             ( u1_col_out_260             ),
    .col_out_261             ( u1_col_out_261             ),
    .col_out_262             ( u1_col_out_262             ),
    .col_out_263             ( u1_col_out_263             ),
    .col_out_264             ( u1_col_out_264             ),
    .col_out_265             ( u1_col_out_265             ),
    .col_out_266             ( u1_col_out_266             ),
    .col_out_267             ( u1_col_out_267             ),
    .col_out_268             ( u1_col_out_268             ),
    .col_out_269             ( u1_col_out_269             ),
    .col_out_270             ( u1_col_out_270             ),
    .col_out_271             ( u1_col_out_271             ),
    .col_out_272             ( u1_col_out_272             ),
    .col_out_273             ( u1_col_out_273             ),
    .col_out_274             ( u1_col_out_274             ),
    .col_out_275             ( u1_col_out_275             ),
    .col_out_276             ( u1_col_out_276             ),
    .col_out_277             ( u1_col_out_277             ),
    .col_out_278             ( u1_col_out_278             ),
    .col_out_279             ( u1_col_out_279             ),
    .col_out_280             ( u1_col_out_280             ),
    .col_out_281             ( u1_col_out_281             ),
    .col_out_282             ( u1_col_out_282             ),
    .col_out_283             ( u1_col_out_283             ),
    .col_out_284             ( u1_col_out_284             ),
    .col_out_285             ( u1_col_out_285             ),
    .col_out_286             ( u1_col_out_286             ),
    .col_out_287             ( u1_col_out_287             ),
    .col_out_288             ( u1_col_out_288             ),
    .col_out_289             ( u1_col_out_289             ),
    .col_out_290             ( u1_col_out_290             ),
    .col_out_291             ( u1_col_out_291             ),
    .col_out_292             ( u1_col_out_292             ),
    .col_out_293             ( u1_col_out_293             ),
    .col_out_294             ( u1_col_out_294             ),
    .col_out_295             ( u1_col_out_295             ),
    .col_out_296             ( u1_col_out_296             ),
    .col_out_297             ( u1_col_out_297             ),
    .col_out_298             ( u1_col_out_298             ),
    .col_out_299             ( u1_col_out_299             ),
    .col_out_300             ( u1_col_out_300             ),
    .col_out_301             ( u1_col_out_301             ),
    .col_out_302             ( u1_col_out_302             ),
    .col_out_303             ( u1_col_out_303             ),
    .col_out_304             ( u1_col_out_304             ),
    .col_out_305             ( u1_col_out_305             ),
    .col_out_306             ( u1_col_out_306             ),
    .col_out_307             ( u1_col_out_307             ),
    .col_out_308             ( u1_col_out_308             ),
    .col_out_309             ( u1_col_out_309             ),
    .col_out_310             ( u1_col_out_310             ),
    .col_out_311             ( u1_col_out_311             ),
    .col_out_312             ( u1_col_out_312             ),
    .col_out_313             ( u1_col_out_313             ),
    .col_out_314             ( u1_col_out_314             ),
    .col_out_315             ( u1_col_out_315             ),
    .col_out_316             ( u1_col_out_316             ),
    .col_out_317             ( u1_col_out_317             ),
    .col_out_318             ( u1_col_out_318             ),
    .col_out_319             ( u1_col_out_319             ),
    .col_out_320             ( u1_col_out_320             ),
    .col_out_321             ( u1_col_out_321             ),
    .col_out_322             ( u1_col_out_322             ),
    .col_out_323             ( u1_col_out_323             ),
    .col_out_324             ( u1_col_out_324             ),
    .col_out_325             ( u1_col_out_325             ),
    .col_out_326             ( u1_col_out_326             ),
    .col_out_327             ( u1_col_out_327             ),
    .col_out_328             ( u1_col_out_328             ),
    .col_out_329             ( u1_col_out_329             ),
    .col_out_330             ( u1_col_out_330             ),
    .col_out_331             ( u1_col_out_331             ),
    .col_out_332             ( u1_col_out_332             ),
    .col_out_333             ( u1_col_out_333             ),
    .col_out_334             ( u1_col_out_334             ),
    .col_out_335             ( u1_col_out_335             ),
    .col_out_336             ( u1_col_out_336             ),
    .col_out_337             ( u1_col_out_337             ),
    .col_out_338             ( u1_col_out_338             ),
    .col_out_339             ( u1_col_out_339             ),
    .col_out_340             ( u1_col_out_340             ),
    .col_out_341             ( u1_col_out_341             ),
    .col_out_342             ( u1_col_out_342             ),
    .col_out_343             ( u1_col_out_343             ),
    .col_out_344             ( u1_col_out_344             ),
    .col_out_345             ( u1_col_out_345             ),
    .col_out_346             ( u1_col_out_346             ),
    .col_out_347             ( u1_col_out_347             ),
    .col_out_348             ( u1_col_out_348             ),
    .col_out_349             ( u1_col_out_349             ),
    .col_out_350             ( u1_col_out_350             ),
    .col_out_351             ( u1_col_out_351             ),
    .col_out_352             ( u1_col_out_352             ),
    .col_out_353             ( u1_col_out_353             ),
    .col_out_354             ( u1_col_out_354             ),
    .col_out_355             ( u1_col_out_355             ),
    .col_out_356             ( u1_col_out_356             ),
    .col_out_357             ( u1_col_out_357             ),
    .col_out_358             ( u1_col_out_358             ),
    .col_out_359             ( u1_col_out_359             ),
    .col_out_360             ( u1_col_out_360             ),
    .col_out_361             ( u1_col_out_361             ),
    .col_out_362             ( u1_col_out_362             ),
    .col_out_363             ( u1_col_out_363             ),
    .col_out_364             ( u1_col_out_364             ),
    .col_out_365             ( u1_col_out_365             ),
    .col_out_366             ( u1_col_out_366             ),
    .col_out_367             ( u1_col_out_367             ),
    .col_out_368             ( u1_col_out_368             ),
    .col_out_369             ( u1_col_out_369             ),
    .col_out_370             ( u1_col_out_370             ),
    .col_out_371             ( u1_col_out_371             ),
    .col_out_372             ( u1_col_out_372             ),
    .col_out_373             ( u1_col_out_373             ),
    .col_out_374             ( u1_col_out_374             ),
    .col_out_375             ( u1_col_out_375             ),
    .col_out_376             ( u1_col_out_376             ),
    .col_out_377             ( u1_col_out_377             ),
    .col_out_378             ( u1_col_out_378             ),
    .col_out_379             ( u1_col_out_379             ),
    .col_out_380             ( u1_col_out_380             ),
    .col_out_381             ( u1_col_out_381             ),
    .col_out_382             ( u1_col_out_382             ),
    .col_out_383             ( u1_col_out_383             ),
    .col_out_384             ( u1_col_out_384             ),
    .col_out_385             ( u1_col_out_385             ),
    .col_out_386             ( u1_col_out_386             ),
    .col_out_387             ( u1_col_out_387             ),
    .col_out_388             ( u1_col_out_388             ),
    .col_out_389             ( u1_col_out_389             ),
    .col_out_390             ( u1_col_out_390             ),
    .col_out_391             ( u1_col_out_391             ),
    .col_out_392             ( u1_col_out_392             ),
    .col_out_393             ( u1_col_out_393             ),
    .col_out_394             ( u1_col_out_394             ),
    .col_out_395             ( u1_col_out_395             ),
    .col_out_396             ( u1_col_out_396             ),
    .col_out_397             ( u1_col_out_397             ),
    .col_out_398             ( u1_col_out_398             ),
    .col_out_399             ( u1_col_out_399             ),
    .col_out_400             ( u1_col_out_400             ),
    .col_out_401             ( u1_col_out_401             ),
    .col_out_402             ( u1_col_out_402             ),
    .col_out_403             ( u1_col_out_403             ),
    .col_out_404             ( u1_col_out_404             ),
    .col_out_405             ( u1_col_out_405             ),
    .col_out_406             ( u1_col_out_406             ),
    .col_out_407             ( u1_col_out_407             ),
    .col_out_408             ( u1_col_out_408             ),
    .col_out_409             ( u1_col_out_409             ),
    .col_out_410             ( u1_col_out_410             ),
    .col_out_411             ( u1_col_out_411             ),
    .col_out_412             ( u1_col_out_412             ),
    .col_out_413             ( u1_col_out_413             ),
    .col_out_414             ( u1_col_out_414             ),
    .col_out_415             ( u1_col_out_415             ),
    .col_out_416             ( u1_col_out_416             ),
    .col_out_417             ( u1_col_out_417             ),
    .col_out_418             ( u1_col_out_418             ),
    .col_out_419             ( u1_col_out_419             ),
    .col_out_420             ( u1_col_out_420             ),
    .col_out_421             ( u1_col_out_421             ),
    .col_out_422             ( u1_col_out_422             ),
    .col_out_423             ( u1_col_out_423             ),
    .col_out_424             ( u1_col_out_424             ),
    .col_out_425             ( u1_col_out_425             ),
    .col_out_426             ( u1_col_out_426             ),
    .col_out_427             ( u1_col_out_427             ),
    .col_out_428             ( u1_col_out_428             ),
    .col_out_429             ( u1_col_out_429             ),
    .col_out_430             ( u1_col_out_430             ),
    .col_out_431             ( u1_col_out_431             ),
    .col_out_432             ( u1_col_out_432             ),
    .col_out_433             ( u1_col_out_433             ),
    .col_out_434             ( u1_col_out_434             ),
    .col_out_435             ( u1_col_out_435             ),
    .col_out_436             ( u1_col_out_436             ),
    .col_out_437             ( u1_col_out_437             ),
    .col_out_438             ( u1_col_out_438             ),
    .col_out_439             ( u1_col_out_439             ),
    .col_out_440             ( u1_col_out_440             ),
    .col_out_441             ( u1_col_out_441             ),
    .col_out_442             ( u1_col_out_442             ),
    .col_out_443             ( u1_col_out_443             ),
    .col_out_444             ( u1_col_out_444             ),
    .col_out_445             ( u1_col_out_445             ),
    .col_out_446             ( u1_col_out_446             ),
    .col_out_447             ( u1_col_out_447             ),
    .col_out_448             ( u1_col_out_448             ),
    .col_out_449             ( u1_col_out_449             ),
    .col_out_450             ( u1_col_out_450             ),
    .col_out_451             ( u1_col_out_451             ),
    .col_out_452             ( u1_col_out_452             ),
    .col_out_453             ( u1_col_out_453             ),
    .col_out_454             ( u1_col_out_454             ),
    .col_out_455             ( u1_col_out_455             ),
    .col_out_456             ( u1_col_out_456             ),
    .col_out_457             ( u1_col_out_457             ),
    .col_out_458             ( u1_col_out_458             ),
    .col_out_459             ( u1_col_out_459             ),
    .col_out_460             ( u1_col_out_460             ),
    .col_out_461             ( u1_col_out_461             ),
    .col_out_462             ( u1_col_out_462             ),
    .col_out_463             ( u1_col_out_463             ),
    .col_out_464             ( u1_col_out_464             ),
    .col_out_465             ( u1_col_out_465             ),
    .col_out_466             ( u1_col_out_466             ),
    .col_out_467             ( u1_col_out_467             ),
    .col_out_468             ( u1_col_out_468             ),
    .col_out_469             ( u1_col_out_469             ),
    .col_out_470             ( u1_col_out_470             ),
    .col_out_471             ( u1_col_out_471             ),
    .col_out_472             ( u1_col_out_472             ),
    .col_out_473             ( u1_col_out_473             ),
    .col_out_474             ( u1_col_out_474             ),
    .col_out_475             ( u1_col_out_475             ),
    .col_out_476             ( u1_col_out_476             ),
    .col_out_477             ( u1_col_out_477             ),
    .col_out_478             ( u1_col_out_478             ),
    .col_out_479             ( u1_col_out_479             ),
    .col_out_480             ( u1_col_out_480             ),
    .col_out_481             ( u1_col_out_481             ),
    .col_out_482             ( u1_col_out_482             ),
    .col_out_483             ( u1_col_out_483             ),
    .col_out_484             ( u1_col_out_484             ),
    .col_out_485             ( u1_col_out_485             ),
    .col_out_486             ( u1_col_out_486             ),
    .col_out_487             ( u1_col_out_487             ),
    .col_out_488             ( u1_col_out_488             ),
    .col_out_489             ( u1_col_out_489             ),
    .col_out_490             ( u1_col_out_490             ),
    .col_out_491             ( u1_col_out_491             ),
    .col_out_492             ( u1_col_out_492             ),
    .col_out_493             ( u1_col_out_493             ),
    .col_out_494             ( u1_col_out_494             ),
    .col_out_495             ( u1_col_out_495             ),
    .col_out_496             ( u1_col_out_496             ),
    .col_out_497             ( u1_col_out_497             ),
    .col_out_498             ( u1_col_out_498             ),
    .col_out_499             ( u1_col_out_499             ),
    .col_out_500             ( u1_col_out_500             ),
    .col_out_501             ( u1_col_out_501             ),
    .col_out_502             ( u1_col_out_502             ),
    .col_out_503             ( u1_col_out_503             ),
    .col_out_504             ( u1_col_out_504             ),
    .col_out_505             ( u1_col_out_505             ),
    .col_out_506             ( u1_col_out_506             ),
    .col_out_507             ( u1_col_out_507             ),
    .col_out_508             ( u1_col_out_508             ),
    .col_out_509             ( u1_col_out_509             ),
    .col_out_510             ( u1_col_out_510             ),
    .col_out_511             ( u1_col_out_511             ),
    .col_out_512             ( u1_col_out_512             ),
    .col_out_513             ( u1_col_out_513             ),
    .col_out_514             ( u1_col_out_514             ),
    .col_out_515             ( u1_col_out_515             ),
    .col_out_516             ( u1_col_out_516             ),
    .col_out_517             ( u1_col_out_517             ),
    .col_out_518             ( u1_col_out_518             ),
    .col_out_519             ( u1_col_out_519             ),
    .col_out_520             ( u1_col_out_520             ),
    .col_out_521             ( u1_col_out_521             ),
    .col_out_522             ( u1_col_out_522             ),
    .col_out_523             ( u1_col_out_523             ),
    .col_out_524             ( u1_col_out_524             ),
    .col_out_525             ( u1_col_out_525             ),
    .col_out_526             ( u1_col_out_526             ),
    .col_out_527             ( u1_col_out_527             ),
    .col_out_528             ( u1_col_out_528             ),
    .col_out_529             ( u1_col_out_529             ),
    .col_out_530             ( u1_col_out_530             ),
    .col_out_531             ( u1_col_out_531             ),
    .col_out_532             ( u1_col_out_532             ),
    .col_out_533             ( u1_col_out_533             ),
    .col_out_534             ( u1_col_out_534             ),
    .col_out_535             ( u1_col_out_535             ),
    .col_out_536             ( u1_col_out_536             ),
    .col_out_537             ( u1_col_out_537             ),
    .col_out_538             ( u1_col_out_538             ),
    .col_out_539             ( u1_col_out_539             ),
    .col_out_540             ( u1_col_out_540             ),
    .col_out_541             ( u1_col_out_541             ),
    .col_out_542             ( u1_col_out_542             ),
    .col_out_543             ( u1_col_out_543             ),
    .col_out_544             ( u1_col_out_544             ),
    .col_out_545             ( u1_col_out_545             ),
    .col_out_546             ( u1_col_out_546             ),
    .col_out_547             ( u1_col_out_547             ),
    .col_out_548             ( u1_col_out_548             ),
    .col_out_549             ( u1_col_out_549             ),
    .col_out_550             ( u1_col_out_550             ),
    .col_out_551             ( u1_col_out_551             ),
    .col_out_552             ( u1_col_out_552             ),
    .col_out_553             ( u1_col_out_553             ),
    .col_out_554             ( u1_col_out_554             ),
    .col_out_555             ( u1_col_out_555             ),
    .col_out_556             ( u1_col_out_556             ),
    .col_out_557             ( u1_col_out_557             ),
    .col_out_558             ( u1_col_out_558             ),
    .col_out_559             ( u1_col_out_559             ),
    .col_out_560             ( u1_col_out_560             ),
    .col_out_561             ( u1_col_out_561             ),
    .col_out_562             ( u1_col_out_562             ),
    .col_out_563             ( u1_col_out_563             ),
    .col_out_564             ( u1_col_out_564             ),
    .col_out_565             ( u1_col_out_565             ),
    .col_out_566             ( u1_col_out_566             ),
    .col_out_567             ( u1_col_out_567             ),
    .col_out_568             ( u1_col_out_568             ),
    .col_out_569             ( u1_col_out_569             ),
    .col_out_570             ( u1_col_out_570             ),
    .col_out_571             ( u1_col_out_571             ),
    .col_out_572             ( u1_col_out_572             ),
    .col_out_573             ( u1_col_out_573             ),
    .col_out_574             ( u1_col_out_574             ),
    .col_out_575             ( u1_col_out_575             ),
    .col_out_576             ( u1_col_out_576             ),
    .col_out_577             ( u1_col_out_577             ),
    .col_out_578             ( u1_col_out_578             ),
    .col_out_579             ( u1_col_out_579             ),
    .col_out_580             ( u1_col_out_580             ),
    .col_out_581             ( u1_col_out_581             ),
    .col_out_582             ( u1_col_out_582             ),
    .col_out_583             ( u1_col_out_583             ),
    .col_out_584             ( u1_col_out_584             ),
    .col_out_585             ( u1_col_out_585             ),
    .col_out_586             ( u1_col_out_586             ),
    .col_out_587             ( u1_col_out_587             ),
    .col_out_588             ( u1_col_out_588             ),
    .col_out_589             ( u1_col_out_589             ),
    .col_out_590             ( u1_col_out_590             ),
    .col_out_591             ( u1_col_out_591             ),
    .col_out_592             ( u1_col_out_592             ),
    .col_out_593             ( u1_col_out_593             ),
    .col_out_594             ( u1_col_out_594             ),
    .col_out_595             ( u1_col_out_595             ),
    .col_out_596             ( u1_col_out_596             ),
    .col_out_597             ( u1_col_out_597             ),
    .col_out_598             ( u1_col_out_598             ),
    .col_out_599             ( u1_col_out_599             ),
    .col_out_600             ( u1_col_out_600             ),
    .col_out_601             ( u1_col_out_601             ),
    .col_out_602             ( u1_col_out_602             ),
    .col_out_603             ( u1_col_out_603             ),
    .col_out_604             ( u1_col_out_604             ),
    .col_out_605             ( u1_col_out_605             ),
    .col_out_606             ( u1_col_out_606             ),
    .col_out_607             ( u1_col_out_607             ),
    .col_out_608             ( u1_col_out_608             ),
    .col_out_609             ( u1_col_out_609             ),
    .col_out_610             ( u1_col_out_610             ),
    .col_out_611             ( u1_col_out_611             ),
    .col_out_612             ( u1_col_out_612             ),
    .col_out_613             ( u1_col_out_613             ),
    .col_out_614             ( u1_col_out_614             ),
    .col_out_615             ( u1_col_out_615             ),
    .col_out_616             ( u1_col_out_616             ),
    .col_out_617             ( u1_col_out_617             ),
    .col_out_618             ( u1_col_out_618             ),
    .col_out_619             ( u1_col_out_619             ),
    .col_out_620             ( u1_col_out_620             ),
    .col_out_621             ( u1_col_out_621             ),
    .col_out_622             ( u1_col_out_622             ),
    .col_out_623             ( u1_col_out_623             ),
    .col_out_624             ( u1_col_out_624             ),
    .col_out_625             ( u1_col_out_625             ),
    .col_out_626             ( u1_col_out_626             ),
    .col_out_627             ( u1_col_out_627             ),
    .col_out_628             ( u1_col_out_628             ),
    .col_out_629             ( u1_col_out_629             ),
    .col_out_630             ( u1_col_out_630             ),
    .col_out_631             ( u1_col_out_631             ),
    .col_out_632             ( u1_col_out_632             ),
    .col_out_633             ( u1_col_out_633             ),
    .col_out_634             ( u1_col_out_634             ),
    .col_out_635             ( u1_col_out_635             ),
    .col_out_636             ( u1_col_out_636             ),
    .col_out_637             ( u1_col_out_637             ),
    .col_out_638             ( u1_col_out_638             ),
    .col_out_639             ( u1_col_out_639             ),
    .col_out_640             ( u1_col_out_640             ),
    .col_out_641             ( u1_col_out_641             ),
    .col_out_642             ( u1_col_out_642             ),
    .col_out_643             ( u1_col_out_643             ),
    .col_out_644             ( u1_col_out_644             ),
    .col_out_645             ( u1_col_out_645             ),
    .col_out_646             ( u1_col_out_646             ),
    .col_out_647             ( u1_col_out_647             ),
    .col_out_648             ( u1_col_out_648             ),
    .col_out_649             ( u1_col_out_649             ),
    .col_out_650             ( u1_col_out_650             ),
    .col_out_651             ( u1_col_out_651             ),
    .col_out_652             ( u1_col_out_652             ),
    .col_out_653             ( u1_col_out_653             ),
    .col_out_654             ( u1_col_out_654             ),
    .col_out_655             ( u1_col_out_655             ),
    .col_out_656             ( u1_col_out_656             ),
    .col_out_657             ( u1_col_out_657             ),
    .col_out_658             ( u1_col_out_658             ),
    .col_out_659             ( u1_col_out_659             ),
    .col_out_660             ( u1_col_out_660             ),
    .col_out_661             ( u1_col_out_661             ),
    .col_out_662             ( u1_col_out_662             ),
    .col_out_663             ( u1_col_out_663             ),
    .col_out_664             ( u1_col_out_664             ),
    .col_out_665             ( u1_col_out_665             ),
    .col_out_666             ( u1_col_out_666             ),
    .col_out_667             ( u1_col_out_667             ),
    .col_out_668             ( u1_col_out_668             ),
    .col_out_669             ( u1_col_out_669             ),
    .col_out_670             ( u1_col_out_670             ),
    .col_out_671             ( u1_col_out_671             ),
    .col_out_672             ( u1_col_out_672             ),
    .col_out_673             ( u1_col_out_673             ),
    .col_out_674             ( u1_col_out_674             ),
    .col_out_675             ( u1_col_out_675             ),
    .col_out_676             ( u1_col_out_676             ),
    .col_out_677             ( u1_col_out_677             ),
    .col_out_678             ( u1_col_out_678             ),
    .col_out_679             ( u1_col_out_679             ),
    .col_out_680             ( u1_col_out_680             ),
    .col_out_681             ( u1_col_out_681             ),
    .col_out_682             ( u1_col_out_682             ),
    .col_out_683             ( u1_col_out_683             ),
    .col_out_684             ( u1_col_out_684             ),
    .col_out_685             ( u1_col_out_685             ),
    .col_out_686             ( u1_col_out_686             ),
    .col_out_687             ( u1_col_out_687             ),
    .col_out_688             ( u1_col_out_688             ),
    .col_out_689             ( u1_col_out_689             ),
    .col_out_690             ( u1_col_out_690             ),
    .col_out_691             ( u1_col_out_691             ),
    .col_out_692             ( u1_col_out_692             ),
    .col_out_693             ( u1_col_out_693             ),
    .col_out_694             ( u1_col_out_694             ),
    .col_out_695             ( u1_col_out_695             ),
    .col_out_696             ( u1_col_out_696             ),
    .col_out_697             ( u1_col_out_697             ),
    .col_out_698             ( u1_col_out_698             ),
    .col_out_699             ( u1_col_out_699             ),
    .col_out_700             ( u1_col_out_700             ),
    .col_out_701             ( u1_col_out_701             ),
    .col_out_702             ( u1_col_out_702             ),
    .col_out_703             ( u1_col_out_703             ),
    .col_out_704             ( u1_col_out_704             ),
    .col_out_705             ( u1_col_out_705             ),
    .col_out_706             ( u1_col_out_706             ),
    .col_out_707             ( u1_col_out_707             ),
    .col_out_708             ( u1_col_out_708             ),
    .col_out_709             ( u1_col_out_709             ),
    .col_out_710             ( u1_col_out_710             ),
    .col_out_711             ( u1_col_out_711             ),
    .col_out_712             ( u1_col_out_712             ),
    .col_out_713             ( u1_col_out_713             ),
    .col_out_714             ( u1_col_out_714             ),
    .col_out_715             ( u1_col_out_715             ),
    .col_out_716             ( u1_col_out_716             ),
    .col_out_717             ( u1_col_out_717             ),
    .col_out_718             ( u1_col_out_718             ),
    .col_out_719             ( u1_col_out_719             ),
    .col_out_720             ( u1_col_out_720             ),
    .col_out_721             ( u1_col_out_721             ),
    .col_out_722             ( u1_col_out_722             ),
    .col_out_723             ( u1_col_out_723             ),
    .col_out_724             ( u1_col_out_724             ),
    .col_out_725             ( u1_col_out_725             ),
    .col_out_726             ( u1_col_out_726             ),
    .col_out_727             ( u1_col_out_727             ),
    .col_out_728             ( u1_col_out_728             ),
    .col_out_729             ( u1_col_out_729             ),
    .col_out_730             ( u1_col_out_730             ),
    .col_out_731             ( u1_col_out_731             ),
    .col_out_732             ( u1_col_out_732             ),
    .col_out_733             ( u1_col_out_733             ),
    .col_out_734             ( u1_col_out_734             ),
    .col_out_735             ( u1_col_out_735             ),
    .col_out_736             ( u1_col_out_736             ),
    .col_out_737             ( u1_col_out_737             ),
    .col_out_738             ( u1_col_out_738             ),
    .col_out_739             ( u1_col_out_739             ),
    .col_out_740             ( u1_col_out_740             ),
    .col_out_741             ( u1_col_out_741             ),
    .col_out_742             ( u1_col_out_742             ),
    .col_out_743             ( u1_col_out_743             ),
    .col_out_744             ( u1_col_out_744             ),
    .col_out_745             ( u1_col_out_745             ),
    .col_out_746             ( u1_col_out_746             ),
    .col_out_747             ( u1_col_out_747             ),
    .col_out_748             ( u1_col_out_748             ),
    .col_out_749             ( u1_col_out_749             ),
    .col_out_750             ( u1_col_out_750             ),
    .col_out_751             ( u1_col_out_751             ),
    .col_out_752             ( u1_col_out_752             ),
    .col_out_753             ( u1_col_out_753             ),
    .col_out_754             ( u1_col_out_754             ),
    .col_out_755             ( u1_col_out_755             ),
    .col_out_756             ( u1_col_out_756             ),
    .col_out_757             ( u1_col_out_757             ),
    .col_out_758             ( u1_col_out_758             ),
    .col_out_759             ( u1_col_out_759             ),
    .col_out_760             ( u1_col_out_760             ),
    .col_out_761             ( u1_col_out_761             ),
    .col_out_762             ( u1_col_out_762             ),
    .col_out_763             ( u1_col_out_763             ),
    .col_out_764             ( u1_col_out_764             ),
    .col_out_765             ( u1_col_out_765             ),
    .col_out_766             ( u1_col_out_766             ),
    .col_out_767             ( u1_col_out_767             ),
    .col_out_768             ( u1_col_out_768             ),
    .col_out_769             ( u1_col_out_769             ),
    .col_out_770             ( u1_col_out_770             ),
    .col_out_771             ( u1_col_out_771             ),
    .col_out_772             ( u1_col_out_772             ),
    .col_out_773             ( u1_col_out_773             ),
    .col_out_774             ( u1_col_out_774             ),
    .col_out_775             ( u1_col_out_775             ),
    .col_out_776             ( u1_col_out_776             ),
    .col_out_777             ( u1_col_out_777             ),
    .col_out_778             ( u1_col_out_778             ),
    .col_out_779             ( u1_col_out_779             ),
    .col_out_780             ( u1_col_out_780             ),
    .col_out_781             ( u1_col_out_781             ),
    .col_out_782             ( u1_col_out_782             ),
    .col_out_783             ( u1_col_out_783             ),
    .col_out_784             ( u1_col_out_784             ),
    .col_out_785             ( u1_col_out_785             ),
    .col_out_786             ( u1_col_out_786             ),
    .col_out_787             ( u1_col_out_787             ),
    .col_out_788             ( u1_col_out_788             ),
    .col_out_789             ( u1_col_out_789             ),
    .col_out_790             ( u1_col_out_790             ),
    .col_out_791             ( u1_col_out_791             ),
    .col_out_792             ( u1_col_out_792             ),
    .col_out_793             ( u1_col_out_793             ),
    .col_out_794             ( u1_col_out_794             ),
    .col_out_795             ( u1_col_out_795             ),
    .col_out_796             ( u1_col_out_796             ),
    .col_out_797             ( u1_col_out_797             ),
    .col_out_798             ( u1_col_out_798             ),
    .col_out_799             ( u1_col_out_799             ),
    .col_out_800             ( u1_col_out_800             ),
    .col_out_801             ( u1_col_out_801             ),
    .col_out_802             ( u1_col_out_802             ),
    .col_out_803             ( u1_col_out_803             ),
    .col_out_804             ( u1_col_out_804             ),
    .col_out_805             ( u1_col_out_805             ),
    .col_out_806             ( u1_col_out_806             ),
    .col_out_807             ( u1_col_out_807             ),
    .col_out_808             ( u1_col_out_808             ),
    .col_out_809             ( u1_col_out_809             ),
    .col_out_810             ( u1_col_out_810             ),
    .col_out_811             ( u1_col_out_811             ),
    .col_out_812             ( u1_col_out_812             ),
    .col_out_813             ( u1_col_out_813             ),
    .col_out_814             ( u1_col_out_814             ),
    .col_out_815             ( u1_col_out_815             ),
    .col_out_816             ( u1_col_out_816             ),
    .col_out_817             ( u1_col_out_817             ),
    .col_out_818             ( u1_col_out_818             ),
    .col_out_819             ( u1_col_out_819             ),
    .col_out_820             ( u1_col_out_820             ),
    .col_out_821             ( u1_col_out_821             ),
    .col_out_822             ( u1_col_out_822             ),
    .col_out_823             ( u1_col_out_823             ),
    .col_out_824             ( u1_col_out_824             ),
    .col_out_825             ( u1_col_out_825             ),
    .col_out_826             ( u1_col_out_826             ),
    .col_out_827             ( u1_col_out_827             ),
    .col_out_828             ( u1_col_out_828             ),
    .col_out_829             ( u1_col_out_829             ),
    .col_out_830             ( u1_col_out_830             ),
    .col_out_831             ( u1_col_out_831             ),
    .col_out_832             ( u1_col_out_832             ),
    .col_out_833             ( u1_col_out_833             ),
    .col_out_834             ( u1_col_out_834             ),
    .col_out_835             ( u1_col_out_835             ),
    .col_out_836             ( u1_col_out_836             ),
    .col_out_837             ( u1_col_out_837             ),
    .col_out_838             ( u1_col_out_838             ),
    .col_out_839             ( u1_col_out_839             ),
    .col_out_840             ( u1_col_out_840             ),
    .col_out_841             ( u1_col_out_841             ),
    .col_out_842             ( u1_col_out_842             ),
    .col_out_843             ( u1_col_out_843             ),
    .col_out_844             ( u1_col_out_844             ),
    .col_out_845             ( u1_col_out_845             ),
    .col_out_846             ( u1_col_out_846             ),
    .col_out_847             ( u1_col_out_847             ),
    .col_out_848             ( u1_col_out_848             ),
    .col_out_849             ( u1_col_out_849             ),
    .col_out_850             ( u1_col_out_850             ),
    .col_out_851             ( u1_col_out_851             ),
    .col_out_852             ( u1_col_out_852             ),
    .col_out_853             ( u1_col_out_853             ),
    .col_out_854             ( u1_col_out_854             ),
    .col_out_855             ( u1_col_out_855             ),
    .col_out_856             ( u1_col_out_856             ),
    .col_out_857             ( u1_col_out_857             ),
    .col_out_858             ( u1_col_out_858             ),
    .col_out_859             ( u1_col_out_859             ),
    .col_out_860             ( u1_col_out_860             ),
    .col_out_861             ( u1_col_out_861             ),
    .col_out_862             ( u1_col_out_862             ),
    .col_out_863             ( u1_col_out_863             ),
    .col_out_864             ( u1_col_out_864             ),
    .col_out_865             ( u1_col_out_865             ),
    .col_out_866             ( u1_col_out_866             ),
    .col_out_867             ( u1_col_out_867             ),
    .col_out_868             ( u1_col_out_868             ),
    .col_out_869             ( u1_col_out_869             ),
    .col_out_870             ( u1_col_out_870             ),
    .col_out_871             ( u1_col_out_871             ),
    .col_out_872             ( u1_col_out_872             ),
    .col_out_873             ( u1_col_out_873             ),
    .col_out_874             ( u1_col_out_874             ),
    .col_out_875             ( u1_col_out_875             ),
    .col_out_876             ( u1_col_out_876             ),
    .col_out_877             ( u1_col_out_877             ),
    .col_out_878             ( u1_col_out_878             ),
    .col_out_879             ( u1_col_out_879             ),
    .col_out_880             ( u1_col_out_880             ),
    .col_out_881             ( u1_col_out_881             ),
    .col_out_882             ( u1_col_out_882             ),
    .col_out_883             ( u1_col_out_883             ),
    .col_out_884             ( u1_col_out_884             ),
    .col_out_885             ( u1_col_out_885             ),
    .col_out_886             ( u1_col_out_886             ),
    .col_out_887             ( u1_col_out_887             ),
    .col_out_888             ( u1_col_out_888             ),
    .col_out_889             ( u1_col_out_889             ),
    .col_out_890             ( u1_col_out_890             ),
    .col_out_891             ( u1_col_out_891             ),
    .col_out_892             ( u1_col_out_892             ),
    .col_out_893             ( u1_col_out_893             ),
    .col_out_894             ( u1_col_out_894             ),
    .col_out_895             ( u1_col_out_895             ),
    .col_out_896             ( u1_col_out_896             ),
    .col_out_897             ( u1_col_out_897             ),
    .col_out_898             ( u1_col_out_898             ),
    .col_out_899             ( u1_col_out_899             ),
    .col_out_900             ( u1_col_out_900             ),
    .col_out_901             ( u1_col_out_901             ),
    .col_out_902             ( u1_col_out_902             ),
    .col_out_903             ( u1_col_out_903             ),
    .col_out_904             ( u1_col_out_904             ),
    .col_out_905             ( u1_col_out_905             ),
    .col_out_906             ( u1_col_out_906             ),
    .col_out_907             ( u1_col_out_907             ),
    .col_out_908             ( u1_col_out_908             ),
    .col_out_909             ( u1_col_out_909             ),
    .col_out_910             ( u1_col_out_910             ),
    .col_out_911             ( u1_col_out_911             ),
    .col_out_912             ( u1_col_out_912             ),
    .col_out_913             ( u1_col_out_913             ),
    .col_out_914             ( u1_col_out_914             ),
    .col_out_915             ( u1_col_out_915             ),
    .col_out_916             ( u1_col_out_916             ),
    .col_out_917             ( u1_col_out_917             ),
    .col_out_918             ( u1_col_out_918             ),
    .col_out_919             ( u1_col_out_919             ),
    .col_out_920             ( u1_col_out_920             ),
    .col_out_921             ( u1_col_out_921             ),
    .col_out_922             ( u1_col_out_922             ),
    .col_out_923             ( u1_col_out_923             ),
    .col_out_924             ( u1_col_out_924             ),
    .col_out_925             ( u1_col_out_925             ),
    .col_out_926             ( u1_col_out_926             ),
    .col_out_927             ( u1_col_out_927             ),
    .col_out_928             ( u1_col_out_928             ),
    .col_out_929             ( u1_col_out_929             ),
    .col_out_930             ( u1_col_out_930             ),
    .col_out_931             ( u1_col_out_931             ),
    .col_out_932             ( u1_col_out_932             ),
    .col_out_933             ( u1_col_out_933             ),
    .col_out_934             ( u1_col_out_934             ),
    .col_out_935             ( u1_col_out_935             ),
    .col_out_936             ( u1_col_out_936             ),
    .col_out_937             ( u1_col_out_937             ),
    .col_out_938             ( u1_col_out_938             ),
    .col_out_939             ( u1_col_out_939             ),
    .col_out_940             ( u1_col_out_940             ),
    .col_out_941             ( u1_col_out_941             ),
    .col_out_942             ( u1_col_out_942             ),
    .col_out_943             ( u1_col_out_943             ),
    .col_out_944             ( u1_col_out_944             ),
    .col_out_945             ( u1_col_out_945             ),
    .col_out_946             ( u1_col_out_946             ),
    .col_out_947             ( u1_col_out_947             ),
    .col_out_948             ( u1_col_out_948             ),
    .col_out_949             ( u1_col_out_949             ),
    .col_out_950             ( u1_col_out_950             ),
    .col_out_951             ( u1_col_out_951             ),
    .col_out_952             ( u1_col_out_952             ),
    .col_out_953             ( u1_col_out_953             ),
    .col_out_954             ( u1_col_out_954             ),
    .col_out_955             ( u1_col_out_955             ),
    .col_out_956             ( u1_col_out_956             ),
    .col_out_957             ( u1_col_out_957             ),
    .col_out_958             ( u1_col_out_958             ),
    .col_out_959             ( u1_col_out_959             ),
    .col_out_960             ( u1_col_out_960             ),
    .col_out_961             ( u1_col_out_961             ),
    .col_out_962             ( u1_col_out_962             ),
    .col_out_963             ( u1_col_out_963             ),
    .col_out_964             ( u1_col_out_964             ),
    .col_out_965             ( u1_col_out_965             ),
    .col_out_966             ( u1_col_out_966             ),
    .col_out_967             ( u1_col_out_967             ),
    .col_out_968             ( u1_col_out_968             ),
    .col_out_969             ( u1_col_out_969             ),
    .col_out_970             ( u1_col_out_970             ),
    .col_out_971             ( u1_col_out_971             ),
    .col_out_972             ( u1_col_out_972             ),
    .col_out_973             ( u1_col_out_973             ),
    .col_out_974             ( u1_col_out_974             ),
    .col_out_975             ( u1_col_out_975             ),
    .col_out_976             ( u1_col_out_976             ),
    .col_out_977             ( u1_col_out_977             ),
    .col_out_978             ( u1_col_out_978             ),
    .col_out_979             ( u1_col_out_979             ),
    .col_out_980             ( u1_col_out_980             ),
    .col_out_981             ( u1_col_out_981             ),
    .col_out_982             ( u1_col_out_982             ),
    .col_out_983             ( u1_col_out_983             ),
    .col_out_984             ( u1_col_out_984             ),
    .col_out_985             ( u1_col_out_985             ),
    .col_out_986             ( u1_col_out_986             ),
    .col_out_987             ( u1_col_out_987             ),
    .col_out_988             ( u1_col_out_988             ),
    .col_out_989             ( u1_col_out_989             ),
    .col_out_990             ( u1_col_out_990             ),
    .col_out_991             ( u1_col_out_991             ),
    .col_out_992             ( u1_col_out_992             ),
    .col_out_993             ( u1_col_out_993             ),
    .col_out_994             ( u1_col_out_994             ),
    .col_out_995             ( u1_col_out_995             ),
    .col_out_996             ( u1_col_out_996             ),
    .col_out_997             ( u1_col_out_997             ),
    .col_out_998             ( u1_col_out_998             ),
    .col_out_999             ( u1_col_out_999             ),
    .col_out_1000            ( u1_col_out_1000            ),
    .col_out_1001            ( u1_col_out_1001            ),
    .col_out_1002            ( u1_col_out_1002            ),
    .col_out_1003            ( u1_col_out_1003            ),
    .col_out_1004            ( u1_col_out_1004            ),
    .col_out_1005            ( u1_col_out_1005            ),
    .col_out_1006            ( u1_col_out_1006            ),
    .col_out_1007            ( u1_col_out_1007            ),
    .col_out_1008            ( u1_col_out_1008            ),
    .col_out_1009            ( u1_col_out_1009            ),
    .col_out_1010            ( u1_col_out_1010            ),
    .col_out_1011            ( u1_col_out_1011            ),
    .col_out_1012            ( u1_col_out_1012            ),
    .col_out_1013            ( u1_col_out_1013            ),
    .col_out_1014            ( u1_col_out_1014            ),
    .col_out_1015            ( u1_col_out_1015            ),
    .col_out_1016            ( u1_col_out_1016            ),
    .col_out_1017            ( u1_col_out_1017            ),
    .col_out_1018            ( u1_col_out_1018            ),
    .col_out_1019            ( u1_col_out_1019            ),
    .col_out_1020            ( u1_col_out_1020            ),
    .col_out_1021            ( u1_col_out_1021            ),
    .col_out_1022            ( u1_col_out_1022            ),
    .col_out_1023            ( u1_col_out_1023            )
);






assign col_out_0 = (sel_data_in)? u0_col_out_0 : u1_col_out_0;
assign col_out_1 = (sel_data_in)? u0_col_out_1 : u1_col_out_1;
assign col_out_2 = (sel_data_in)? u0_col_out_2 : u1_col_out_2;
assign col_out_3 = (sel_data_in)? u0_col_out_3 : u1_col_out_3;
assign col_out_4 = (sel_data_in)? u0_col_out_4 : u1_col_out_4;
assign col_out_5 = (sel_data_in)? u0_col_out_5 : u1_col_out_5;
assign col_out_6 = (sel_data_in)? u0_col_out_6 : u1_col_out_6;
assign col_out_7 = (sel_data_in)? u0_col_out_7 : u1_col_out_7;
assign col_out_8 = (sel_data_in)? u0_col_out_8 : u1_col_out_8;
assign col_out_9 = (sel_data_in)? u0_col_out_9 : u1_col_out_9;
assign col_out_10 = (sel_data_in)? u0_col_out_10 : u1_col_out_10;
assign col_out_11 = (sel_data_in)? u0_col_out_11 : u1_col_out_11;
assign col_out_12 = (sel_data_in)? u0_col_out_12 : u1_col_out_12;
assign col_out_13 = (sel_data_in)? u0_col_out_13 : u1_col_out_13;
assign col_out_14 = (sel_data_in)? u0_col_out_14 : u1_col_out_14;
assign col_out_15 = (sel_data_in)? u0_col_out_15 : u1_col_out_15;
assign col_out_16 = (sel_data_in)? u0_col_out_16 : u1_col_out_16;
assign col_out_17 = (sel_data_in)? u0_col_out_17 : u1_col_out_17;
assign col_out_18 = (sel_data_in)? u0_col_out_18 : u1_col_out_18;
assign col_out_19 = (sel_data_in)? u0_col_out_19 : u1_col_out_19;
assign col_out_20 = (sel_data_in)? u0_col_out_20 : u1_col_out_20;
assign col_out_21 = (sel_data_in)? u0_col_out_21 : u1_col_out_21;
assign col_out_22 = (sel_data_in)? u0_col_out_22 : u1_col_out_22;
assign col_out_23 = (sel_data_in)? u0_col_out_23 : u1_col_out_23;
assign col_out_24 = (sel_data_in)? u0_col_out_24 : u1_col_out_24;
assign col_out_25 = (sel_data_in)? u0_col_out_25 : u1_col_out_25;
assign col_out_26 = (sel_data_in)? u0_col_out_26 : u1_col_out_26;
assign col_out_27 = (sel_data_in)? u0_col_out_27 : u1_col_out_27;
assign col_out_28 = (sel_data_in)? u0_col_out_28 : u1_col_out_28;
assign col_out_29 = (sel_data_in)? u0_col_out_29 : u1_col_out_29;
assign col_out_30 = (sel_data_in)? u0_col_out_30 : u1_col_out_30;
assign col_out_31 = (sel_data_in)? u0_col_out_31 : u1_col_out_31;
assign col_out_32 = (sel_data_in)? u0_col_out_32 : u1_col_out_32;
assign col_out_33 = (sel_data_in)? u0_col_out_33 : u1_col_out_33;
assign col_out_34 = (sel_data_in)? u0_col_out_34 : u1_col_out_34;
assign col_out_35 = (sel_data_in)? u0_col_out_35 : u1_col_out_35;
assign col_out_36 = (sel_data_in)? u0_col_out_36 : u1_col_out_36;
assign col_out_37 = (sel_data_in)? u0_col_out_37 : u1_col_out_37;
assign col_out_38 = (sel_data_in)? u0_col_out_38 : u1_col_out_38;
assign col_out_39 = (sel_data_in)? u0_col_out_39 : u1_col_out_39;
assign col_out_40 = (sel_data_in)? u0_col_out_40 : u1_col_out_40;
assign col_out_41 = (sel_data_in)? u0_col_out_41 : u1_col_out_41;
assign col_out_42 = (sel_data_in)? u0_col_out_42 : u1_col_out_42;
assign col_out_43 = (sel_data_in)? u0_col_out_43 : u1_col_out_43;
assign col_out_44 = (sel_data_in)? u0_col_out_44 : u1_col_out_44;
assign col_out_45 = (sel_data_in)? u0_col_out_45 : u1_col_out_45;
assign col_out_46 = (sel_data_in)? u0_col_out_46 : u1_col_out_46;
assign col_out_47 = (sel_data_in)? u0_col_out_47 : u1_col_out_47;
assign col_out_48 = (sel_data_in)? u0_col_out_48 : u1_col_out_48;
assign col_out_49 = (sel_data_in)? u0_col_out_49 : u1_col_out_49;
assign col_out_50 = (sel_data_in)? u0_col_out_50 : u1_col_out_50;
assign col_out_51 = (sel_data_in)? u0_col_out_51 : u1_col_out_51;
assign col_out_52 = (sel_data_in)? u0_col_out_52 : u1_col_out_52;
assign col_out_53 = (sel_data_in)? u0_col_out_53 : u1_col_out_53;
assign col_out_54 = (sel_data_in)? u0_col_out_54 : u1_col_out_54;
assign col_out_55 = (sel_data_in)? u0_col_out_55 : u1_col_out_55;
assign col_out_56 = (sel_data_in)? u0_col_out_56 : u1_col_out_56;
assign col_out_57 = (sel_data_in)? u0_col_out_57 : u1_col_out_57;
assign col_out_58 = (sel_data_in)? u0_col_out_58 : u1_col_out_58;
assign col_out_59 = (sel_data_in)? u0_col_out_59 : u1_col_out_59;
assign col_out_60 = (sel_data_in)? u0_col_out_60 : u1_col_out_60;
assign col_out_61 = (sel_data_in)? u0_col_out_61 : u1_col_out_61;
assign col_out_62 = (sel_data_in)? u0_col_out_62 : u1_col_out_62;
assign col_out_63 = (sel_data_in)? u0_col_out_63 : u1_col_out_63;
assign col_out_64 = (sel_data_in)? u0_col_out_64 : u1_col_out_64;
assign col_out_65 = (sel_data_in)? u0_col_out_65 : u1_col_out_65;
assign col_out_66 = (sel_data_in)? u0_col_out_66 : u1_col_out_66;
assign col_out_67 = (sel_data_in)? u0_col_out_67 : u1_col_out_67;
assign col_out_68 = (sel_data_in)? u0_col_out_68 : u1_col_out_68;
assign col_out_69 = (sel_data_in)? u0_col_out_69 : u1_col_out_69;
assign col_out_70 = (sel_data_in)? u0_col_out_70 : u1_col_out_70;
assign col_out_71 = (sel_data_in)? u0_col_out_71 : u1_col_out_71;
assign col_out_72 = (sel_data_in)? u0_col_out_72 : u1_col_out_72;
assign col_out_73 = (sel_data_in)? u0_col_out_73 : u1_col_out_73;
assign col_out_74 = (sel_data_in)? u0_col_out_74 : u1_col_out_74;
assign col_out_75 = (sel_data_in)? u0_col_out_75 : u1_col_out_75;
assign col_out_76 = (sel_data_in)? u0_col_out_76 : u1_col_out_76;
assign col_out_77 = (sel_data_in)? u0_col_out_77 : u1_col_out_77;
assign col_out_78 = (sel_data_in)? u0_col_out_78 : u1_col_out_78;
assign col_out_79 = (sel_data_in)? u0_col_out_79 : u1_col_out_79;
assign col_out_80 = (sel_data_in)? u0_col_out_80 : u1_col_out_80;
assign col_out_81 = (sel_data_in)? u0_col_out_81 : u1_col_out_81;
assign col_out_82 = (sel_data_in)? u0_col_out_82 : u1_col_out_82;
assign col_out_83 = (sel_data_in)? u0_col_out_83 : u1_col_out_83;
assign col_out_84 = (sel_data_in)? u0_col_out_84 : u1_col_out_84;
assign col_out_85 = (sel_data_in)? u0_col_out_85 : u1_col_out_85;
assign col_out_86 = (sel_data_in)? u0_col_out_86 : u1_col_out_86;
assign col_out_87 = (sel_data_in)? u0_col_out_87 : u1_col_out_87;
assign col_out_88 = (sel_data_in)? u0_col_out_88 : u1_col_out_88;
assign col_out_89 = (sel_data_in)? u0_col_out_89 : u1_col_out_89;
assign col_out_90 = (sel_data_in)? u0_col_out_90 : u1_col_out_90;
assign col_out_91 = (sel_data_in)? u0_col_out_91 : u1_col_out_91;
assign col_out_92 = (sel_data_in)? u0_col_out_92 : u1_col_out_92;
assign col_out_93 = (sel_data_in)? u0_col_out_93 : u1_col_out_93;
assign col_out_94 = (sel_data_in)? u0_col_out_94 : u1_col_out_94;
assign col_out_95 = (sel_data_in)? u0_col_out_95 : u1_col_out_95;
assign col_out_96 = (sel_data_in)? u0_col_out_96 : u1_col_out_96;
assign col_out_97 = (sel_data_in)? u0_col_out_97 : u1_col_out_97;
assign col_out_98 = (sel_data_in)? u0_col_out_98 : u1_col_out_98;
assign col_out_99 = (sel_data_in)? u0_col_out_99 : u1_col_out_99;
assign col_out_100 = (sel_data_in)? u0_col_out_100 : u1_col_out_100;
assign col_out_101 = (sel_data_in)? u0_col_out_101 : u1_col_out_101;
assign col_out_102 = (sel_data_in)? u0_col_out_102 : u1_col_out_102;
assign col_out_103 = (sel_data_in)? u0_col_out_103 : u1_col_out_103;
assign col_out_104 = (sel_data_in)? u0_col_out_104 : u1_col_out_104;
assign col_out_105 = (sel_data_in)? u0_col_out_105 : u1_col_out_105;
assign col_out_106 = (sel_data_in)? u0_col_out_106 : u1_col_out_106;
assign col_out_107 = (sel_data_in)? u0_col_out_107 : u1_col_out_107;
assign col_out_108 = (sel_data_in)? u0_col_out_108 : u1_col_out_108;
assign col_out_109 = (sel_data_in)? u0_col_out_109 : u1_col_out_109;
assign col_out_110 = (sel_data_in)? u0_col_out_110 : u1_col_out_110;
assign col_out_111 = (sel_data_in)? u0_col_out_111 : u1_col_out_111;
assign col_out_112 = (sel_data_in)? u0_col_out_112 : u1_col_out_112;
assign col_out_113 = (sel_data_in)? u0_col_out_113 : u1_col_out_113;
assign col_out_114 = (sel_data_in)? u0_col_out_114 : u1_col_out_114;
assign col_out_115 = (sel_data_in)? u0_col_out_115 : u1_col_out_115;
assign col_out_116 = (sel_data_in)? u0_col_out_116 : u1_col_out_116;
assign col_out_117 = (sel_data_in)? u0_col_out_117 : u1_col_out_117;
assign col_out_118 = (sel_data_in)? u0_col_out_118 : u1_col_out_118;
assign col_out_119 = (sel_data_in)? u0_col_out_119 : u1_col_out_119;
assign col_out_120 = (sel_data_in)? u0_col_out_120 : u1_col_out_120;
assign col_out_121 = (sel_data_in)? u0_col_out_121 : u1_col_out_121;
assign col_out_122 = (sel_data_in)? u0_col_out_122 : u1_col_out_122;
assign col_out_123 = (sel_data_in)? u0_col_out_123 : u1_col_out_123;
assign col_out_124 = (sel_data_in)? u0_col_out_124 : u1_col_out_124;
assign col_out_125 = (sel_data_in)? u0_col_out_125 : u1_col_out_125;
assign col_out_126 = (sel_data_in)? u0_col_out_126 : u1_col_out_126;
assign col_out_127 = (sel_data_in)? u0_col_out_127 : u1_col_out_127;
assign col_out_128 = (sel_data_in)? u0_col_out_128 : u1_col_out_128;
assign col_out_129 = (sel_data_in)? u0_col_out_129 : u1_col_out_129;
assign col_out_130 = (sel_data_in)? u0_col_out_130 : u1_col_out_130;
assign col_out_131 = (sel_data_in)? u0_col_out_131 : u1_col_out_131;
assign col_out_132 = (sel_data_in)? u0_col_out_132 : u1_col_out_132;
assign col_out_133 = (sel_data_in)? u0_col_out_133 : u1_col_out_133;
assign col_out_134 = (sel_data_in)? u0_col_out_134 : u1_col_out_134;
assign col_out_135 = (sel_data_in)? u0_col_out_135 : u1_col_out_135;
assign col_out_136 = (sel_data_in)? u0_col_out_136 : u1_col_out_136;
assign col_out_137 = (sel_data_in)? u0_col_out_137 : u1_col_out_137;
assign col_out_138 = (sel_data_in)? u0_col_out_138 : u1_col_out_138;
assign col_out_139 = (sel_data_in)? u0_col_out_139 : u1_col_out_139;
assign col_out_140 = (sel_data_in)? u0_col_out_140 : u1_col_out_140;
assign col_out_141 = (sel_data_in)? u0_col_out_141 : u1_col_out_141;
assign col_out_142 = (sel_data_in)? u0_col_out_142 : u1_col_out_142;
assign col_out_143 = (sel_data_in)? u0_col_out_143 : u1_col_out_143;
assign col_out_144 = (sel_data_in)? u0_col_out_144 : u1_col_out_144;
assign col_out_145 = (sel_data_in)? u0_col_out_145 : u1_col_out_145;
assign col_out_146 = (sel_data_in)? u0_col_out_146 : u1_col_out_146;
assign col_out_147 = (sel_data_in)? u0_col_out_147 : u1_col_out_147;
assign col_out_148 = (sel_data_in)? u0_col_out_148 : u1_col_out_148;
assign col_out_149 = (sel_data_in)? u0_col_out_149 : u1_col_out_149;
assign col_out_150 = (sel_data_in)? u0_col_out_150 : u1_col_out_150;
assign col_out_151 = (sel_data_in)? u0_col_out_151 : u1_col_out_151;
assign col_out_152 = (sel_data_in)? u0_col_out_152 : u1_col_out_152;
assign col_out_153 = (sel_data_in)? u0_col_out_153 : u1_col_out_153;
assign col_out_154 = (sel_data_in)? u0_col_out_154 : u1_col_out_154;
assign col_out_155 = (sel_data_in)? u0_col_out_155 : u1_col_out_155;
assign col_out_156 = (sel_data_in)? u0_col_out_156 : u1_col_out_156;
assign col_out_157 = (sel_data_in)? u0_col_out_157 : u1_col_out_157;
assign col_out_158 = (sel_data_in)? u0_col_out_158 : u1_col_out_158;
assign col_out_159 = (sel_data_in)? u0_col_out_159 : u1_col_out_159;
assign col_out_160 = (sel_data_in)? u0_col_out_160 : u1_col_out_160;
assign col_out_161 = (sel_data_in)? u0_col_out_161 : u1_col_out_161;
assign col_out_162 = (sel_data_in)? u0_col_out_162 : u1_col_out_162;
assign col_out_163 = (sel_data_in)? u0_col_out_163 : u1_col_out_163;
assign col_out_164 = (sel_data_in)? u0_col_out_164 : u1_col_out_164;
assign col_out_165 = (sel_data_in)? u0_col_out_165 : u1_col_out_165;
assign col_out_166 = (sel_data_in)? u0_col_out_166 : u1_col_out_166;
assign col_out_167 = (sel_data_in)? u0_col_out_167 : u1_col_out_167;
assign col_out_168 = (sel_data_in)? u0_col_out_168 : u1_col_out_168;
assign col_out_169 = (sel_data_in)? u0_col_out_169 : u1_col_out_169;
assign col_out_170 = (sel_data_in)? u0_col_out_170 : u1_col_out_170;
assign col_out_171 = (sel_data_in)? u0_col_out_171 : u1_col_out_171;
assign col_out_172 = (sel_data_in)? u0_col_out_172 : u1_col_out_172;
assign col_out_173 = (sel_data_in)? u0_col_out_173 : u1_col_out_173;
assign col_out_174 = (sel_data_in)? u0_col_out_174 : u1_col_out_174;
assign col_out_175 = (sel_data_in)? u0_col_out_175 : u1_col_out_175;
assign col_out_176 = (sel_data_in)? u0_col_out_176 : u1_col_out_176;
assign col_out_177 = (sel_data_in)? u0_col_out_177 : u1_col_out_177;
assign col_out_178 = (sel_data_in)? u0_col_out_178 : u1_col_out_178;
assign col_out_179 = (sel_data_in)? u0_col_out_179 : u1_col_out_179;
assign col_out_180 = (sel_data_in)? u0_col_out_180 : u1_col_out_180;
assign col_out_181 = (sel_data_in)? u0_col_out_181 : u1_col_out_181;
assign col_out_182 = (sel_data_in)? u0_col_out_182 : u1_col_out_182;
assign col_out_183 = (sel_data_in)? u0_col_out_183 : u1_col_out_183;
assign col_out_184 = (sel_data_in)? u0_col_out_184 : u1_col_out_184;
assign col_out_185 = (sel_data_in)? u0_col_out_185 : u1_col_out_185;
assign col_out_186 = (sel_data_in)? u0_col_out_186 : u1_col_out_186;
assign col_out_187 = (sel_data_in)? u0_col_out_187 : u1_col_out_187;
assign col_out_188 = (sel_data_in)? u0_col_out_188 : u1_col_out_188;
assign col_out_189 = (sel_data_in)? u0_col_out_189 : u1_col_out_189;
assign col_out_190 = (sel_data_in)? u0_col_out_190 : u1_col_out_190;
assign col_out_191 = (sel_data_in)? u0_col_out_191 : u1_col_out_191;
assign col_out_192 = (sel_data_in)? u0_col_out_192 : u1_col_out_192;
assign col_out_193 = (sel_data_in)? u0_col_out_193 : u1_col_out_193;
assign col_out_194 = (sel_data_in)? u0_col_out_194 : u1_col_out_194;
assign col_out_195 = (sel_data_in)? u0_col_out_195 : u1_col_out_195;
assign col_out_196 = (sel_data_in)? u0_col_out_196 : u1_col_out_196;
assign col_out_197 = (sel_data_in)? u0_col_out_197 : u1_col_out_197;
assign col_out_198 = (sel_data_in)? u0_col_out_198 : u1_col_out_198;
assign col_out_199 = (sel_data_in)? u0_col_out_199 : u1_col_out_199;
assign col_out_200 = (sel_data_in)? u0_col_out_200 : u1_col_out_200;
assign col_out_201 = (sel_data_in)? u0_col_out_201 : u1_col_out_201;
assign col_out_202 = (sel_data_in)? u0_col_out_202 : u1_col_out_202;
assign col_out_203 = (sel_data_in)? u0_col_out_203 : u1_col_out_203;
assign col_out_204 = (sel_data_in)? u0_col_out_204 : u1_col_out_204;
assign col_out_205 = (sel_data_in)? u0_col_out_205 : u1_col_out_205;
assign col_out_206 = (sel_data_in)? u0_col_out_206 : u1_col_out_206;
assign col_out_207 = (sel_data_in)? u0_col_out_207 : u1_col_out_207;
assign col_out_208 = (sel_data_in)? u0_col_out_208 : u1_col_out_208;
assign col_out_209 = (sel_data_in)? u0_col_out_209 : u1_col_out_209;
assign col_out_210 = (sel_data_in)? u0_col_out_210 : u1_col_out_210;
assign col_out_211 = (sel_data_in)? u0_col_out_211 : u1_col_out_211;
assign col_out_212 = (sel_data_in)? u0_col_out_212 : u1_col_out_212;
assign col_out_213 = (sel_data_in)? u0_col_out_213 : u1_col_out_213;
assign col_out_214 = (sel_data_in)? u0_col_out_214 : u1_col_out_214;
assign col_out_215 = (sel_data_in)? u0_col_out_215 : u1_col_out_215;
assign col_out_216 = (sel_data_in)? u0_col_out_216 : u1_col_out_216;
assign col_out_217 = (sel_data_in)? u0_col_out_217 : u1_col_out_217;
assign col_out_218 = (sel_data_in)? u0_col_out_218 : u1_col_out_218;
assign col_out_219 = (sel_data_in)? u0_col_out_219 : u1_col_out_219;
assign col_out_220 = (sel_data_in)? u0_col_out_220 : u1_col_out_220;
assign col_out_221 = (sel_data_in)? u0_col_out_221 : u1_col_out_221;
assign col_out_222 = (sel_data_in)? u0_col_out_222 : u1_col_out_222;
assign col_out_223 = (sel_data_in)? u0_col_out_223 : u1_col_out_223;
assign col_out_224 = (sel_data_in)? u0_col_out_224 : u1_col_out_224;
assign col_out_225 = (sel_data_in)? u0_col_out_225 : u1_col_out_225;
assign col_out_226 = (sel_data_in)? u0_col_out_226 : u1_col_out_226;
assign col_out_227 = (sel_data_in)? u0_col_out_227 : u1_col_out_227;
assign col_out_228 = (sel_data_in)? u0_col_out_228 : u1_col_out_228;
assign col_out_229 = (sel_data_in)? u0_col_out_229 : u1_col_out_229;
assign col_out_230 = (sel_data_in)? u0_col_out_230 : u1_col_out_230;
assign col_out_231 = (sel_data_in)? u0_col_out_231 : u1_col_out_231;
assign col_out_232 = (sel_data_in)? u0_col_out_232 : u1_col_out_232;
assign col_out_233 = (sel_data_in)? u0_col_out_233 : u1_col_out_233;
assign col_out_234 = (sel_data_in)? u0_col_out_234 : u1_col_out_234;
assign col_out_235 = (sel_data_in)? u0_col_out_235 : u1_col_out_235;
assign col_out_236 = (sel_data_in)? u0_col_out_236 : u1_col_out_236;
assign col_out_237 = (sel_data_in)? u0_col_out_237 : u1_col_out_237;
assign col_out_238 = (sel_data_in)? u0_col_out_238 : u1_col_out_238;
assign col_out_239 = (sel_data_in)? u0_col_out_239 : u1_col_out_239;
assign col_out_240 = (sel_data_in)? u0_col_out_240 : u1_col_out_240;
assign col_out_241 = (sel_data_in)? u0_col_out_241 : u1_col_out_241;
assign col_out_242 = (sel_data_in)? u0_col_out_242 : u1_col_out_242;
assign col_out_243 = (sel_data_in)? u0_col_out_243 : u1_col_out_243;
assign col_out_244 = (sel_data_in)? u0_col_out_244 : u1_col_out_244;
assign col_out_245 = (sel_data_in)? u0_col_out_245 : u1_col_out_245;
assign col_out_246 = (sel_data_in)? u0_col_out_246 : u1_col_out_246;
assign col_out_247 = (sel_data_in)? u0_col_out_247 : u1_col_out_247;
assign col_out_248 = (sel_data_in)? u0_col_out_248 : u1_col_out_248;
assign col_out_249 = (sel_data_in)? u0_col_out_249 : u1_col_out_249;
assign col_out_250 = (sel_data_in)? u0_col_out_250 : u1_col_out_250;
assign col_out_251 = (sel_data_in)? u0_col_out_251 : u1_col_out_251;
assign col_out_252 = (sel_data_in)? u0_col_out_252 : u1_col_out_252;
assign col_out_253 = (sel_data_in)? u0_col_out_253 : u1_col_out_253;
assign col_out_254 = (sel_data_in)? u0_col_out_254 : u1_col_out_254;
assign col_out_255 = (sel_data_in)? u0_col_out_255 : u1_col_out_255;
assign col_out_256 = (sel_data_in)? u0_col_out_256 : u1_col_out_256;
assign col_out_257 = (sel_data_in)? u0_col_out_257 : u1_col_out_257;
assign col_out_258 = (sel_data_in)? u0_col_out_258 : u1_col_out_258;
assign col_out_259 = (sel_data_in)? u0_col_out_259 : u1_col_out_259;
assign col_out_260 = (sel_data_in)? u0_col_out_260 : u1_col_out_260;
assign col_out_261 = (sel_data_in)? u0_col_out_261 : u1_col_out_261;
assign col_out_262 = (sel_data_in)? u0_col_out_262 : u1_col_out_262;
assign col_out_263 = (sel_data_in)? u0_col_out_263 : u1_col_out_263;
assign col_out_264 = (sel_data_in)? u0_col_out_264 : u1_col_out_264;
assign col_out_265 = (sel_data_in)? u0_col_out_265 : u1_col_out_265;
assign col_out_266 = (sel_data_in)? u0_col_out_266 : u1_col_out_266;
assign col_out_267 = (sel_data_in)? u0_col_out_267 : u1_col_out_267;
assign col_out_268 = (sel_data_in)? u0_col_out_268 : u1_col_out_268;
assign col_out_269 = (sel_data_in)? u0_col_out_269 : u1_col_out_269;
assign col_out_270 = (sel_data_in)? u0_col_out_270 : u1_col_out_270;
assign col_out_271 = (sel_data_in)? u0_col_out_271 : u1_col_out_271;
assign col_out_272 = (sel_data_in)? u0_col_out_272 : u1_col_out_272;
assign col_out_273 = (sel_data_in)? u0_col_out_273 : u1_col_out_273;
assign col_out_274 = (sel_data_in)? u0_col_out_274 : u1_col_out_274;
assign col_out_275 = (sel_data_in)? u0_col_out_275 : u1_col_out_275;
assign col_out_276 = (sel_data_in)? u0_col_out_276 : u1_col_out_276;
assign col_out_277 = (sel_data_in)? u0_col_out_277 : u1_col_out_277;
assign col_out_278 = (sel_data_in)? u0_col_out_278 : u1_col_out_278;
assign col_out_279 = (sel_data_in)? u0_col_out_279 : u1_col_out_279;
assign col_out_280 = (sel_data_in)? u0_col_out_280 : u1_col_out_280;
assign col_out_281 = (sel_data_in)? u0_col_out_281 : u1_col_out_281;
assign col_out_282 = (sel_data_in)? u0_col_out_282 : u1_col_out_282;
assign col_out_283 = (sel_data_in)? u0_col_out_283 : u1_col_out_283;
assign col_out_284 = (sel_data_in)? u0_col_out_284 : u1_col_out_284;
assign col_out_285 = (sel_data_in)? u0_col_out_285 : u1_col_out_285;
assign col_out_286 = (sel_data_in)? u0_col_out_286 : u1_col_out_286;
assign col_out_287 = (sel_data_in)? u0_col_out_287 : u1_col_out_287;
assign col_out_288 = (sel_data_in)? u0_col_out_288 : u1_col_out_288;
assign col_out_289 = (sel_data_in)? u0_col_out_289 : u1_col_out_289;
assign col_out_290 = (sel_data_in)? u0_col_out_290 : u1_col_out_290;
assign col_out_291 = (sel_data_in)? u0_col_out_291 : u1_col_out_291;
assign col_out_292 = (sel_data_in)? u0_col_out_292 : u1_col_out_292;
assign col_out_293 = (sel_data_in)? u0_col_out_293 : u1_col_out_293;
assign col_out_294 = (sel_data_in)? u0_col_out_294 : u1_col_out_294;
assign col_out_295 = (sel_data_in)? u0_col_out_295 : u1_col_out_295;
assign col_out_296 = (sel_data_in)? u0_col_out_296 : u1_col_out_296;
assign col_out_297 = (sel_data_in)? u0_col_out_297 : u1_col_out_297;
assign col_out_298 = (sel_data_in)? u0_col_out_298 : u1_col_out_298;
assign col_out_299 = (sel_data_in)? u0_col_out_299 : u1_col_out_299;
assign col_out_300 = (sel_data_in)? u0_col_out_300 : u1_col_out_300;
assign col_out_301 = (sel_data_in)? u0_col_out_301 : u1_col_out_301;
assign col_out_302 = (sel_data_in)? u0_col_out_302 : u1_col_out_302;
assign col_out_303 = (sel_data_in)? u0_col_out_303 : u1_col_out_303;
assign col_out_304 = (sel_data_in)? u0_col_out_304 : u1_col_out_304;
assign col_out_305 = (sel_data_in)? u0_col_out_305 : u1_col_out_305;
assign col_out_306 = (sel_data_in)? u0_col_out_306 : u1_col_out_306;
assign col_out_307 = (sel_data_in)? u0_col_out_307 : u1_col_out_307;
assign col_out_308 = (sel_data_in)? u0_col_out_308 : u1_col_out_308;
assign col_out_309 = (sel_data_in)? u0_col_out_309 : u1_col_out_309;
assign col_out_310 = (sel_data_in)? u0_col_out_310 : u1_col_out_310;
assign col_out_311 = (sel_data_in)? u0_col_out_311 : u1_col_out_311;
assign col_out_312 = (sel_data_in)? u0_col_out_312 : u1_col_out_312;
assign col_out_313 = (sel_data_in)? u0_col_out_313 : u1_col_out_313;
assign col_out_314 = (sel_data_in)? u0_col_out_314 : u1_col_out_314;
assign col_out_315 = (sel_data_in)? u0_col_out_315 : u1_col_out_315;
assign col_out_316 = (sel_data_in)? u0_col_out_316 : u1_col_out_316;
assign col_out_317 = (sel_data_in)? u0_col_out_317 : u1_col_out_317;
assign col_out_318 = (sel_data_in)? u0_col_out_318 : u1_col_out_318;
assign col_out_319 = (sel_data_in)? u0_col_out_319 : u1_col_out_319;
assign col_out_320 = (sel_data_in)? u0_col_out_320 : u1_col_out_320;
assign col_out_321 = (sel_data_in)? u0_col_out_321 : u1_col_out_321;
assign col_out_322 = (sel_data_in)? u0_col_out_322 : u1_col_out_322;
assign col_out_323 = (sel_data_in)? u0_col_out_323 : u1_col_out_323;
assign col_out_324 = (sel_data_in)? u0_col_out_324 : u1_col_out_324;
assign col_out_325 = (sel_data_in)? u0_col_out_325 : u1_col_out_325;
assign col_out_326 = (sel_data_in)? u0_col_out_326 : u1_col_out_326;
assign col_out_327 = (sel_data_in)? u0_col_out_327 : u1_col_out_327;
assign col_out_328 = (sel_data_in)? u0_col_out_328 : u1_col_out_328;
assign col_out_329 = (sel_data_in)? u0_col_out_329 : u1_col_out_329;
assign col_out_330 = (sel_data_in)? u0_col_out_330 : u1_col_out_330;
assign col_out_331 = (sel_data_in)? u0_col_out_331 : u1_col_out_331;
assign col_out_332 = (sel_data_in)? u0_col_out_332 : u1_col_out_332;
assign col_out_333 = (sel_data_in)? u0_col_out_333 : u1_col_out_333;
assign col_out_334 = (sel_data_in)? u0_col_out_334 : u1_col_out_334;
assign col_out_335 = (sel_data_in)? u0_col_out_335 : u1_col_out_335;
assign col_out_336 = (sel_data_in)? u0_col_out_336 : u1_col_out_336;
assign col_out_337 = (sel_data_in)? u0_col_out_337 : u1_col_out_337;
assign col_out_338 = (sel_data_in)? u0_col_out_338 : u1_col_out_338;
assign col_out_339 = (sel_data_in)? u0_col_out_339 : u1_col_out_339;
assign col_out_340 = (sel_data_in)? u0_col_out_340 : u1_col_out_340;
assign col_out_341 = (sel_data_in)? u0_col_out_341 : u1_col_out_341;
assign col_out_342 = (sel_data_in)? u0_col_out_342 : u1_col_out_342;
assign col_out_343 = (sel_data_in)? u0_col_out_343 : u1_col_out_343;
assign col_out_344 = (sel_data_in)? u0_col_out_344 : u1_col_out_344;
assign col_out_345 = (sel_data_in)? u0_col_out_345 : u1_col_out_345;
assign col_out_346 = (sel_data_in)? u0_col_out_346 : u1_col_out_346;
assign col_out_347 = (sel_data_in)? u0_col_out_347 : u1_col_out_347;
assign col_out_348 = (sel_data_in)? u0_col_out_348 : u1_col_out_348;
assign col_out_349 = (sel_data_in)? u0_col_out_349 : u1_col_out_349;
assign col_out_350 = (sel_data_in)? u0_col_out_350 : u1_col_out_350;
assign col_out_351 = (sel_data_in)? u0_col_out_351 : u1_col_out_351;
assign col_out_352 = (sel_data_in)? u0_col_out_352 : u1_col_out_352;
assign col_out_353 = (sel_data_in)? u0_col_out_353 : u1_col_out_353;
assign col_out_354 = (sel_data_in)? u0_col_out_354 : u1_col_out_354;
assign col_out_355 = (sel_data_in)? u0_col_out_355 : u1_col_out_355;
assign col_out_356 = (sel_data_in)? u0_col_out_356 : u1_col_out_356;
assign col_out_357 = (sel_data_in)? u0_col_out_357 : u1_col_out_357;
assign col_out_358 = (sel_data_in)? u0_col_out_358 : u1_col_out_358;
assign col_out_359 = (sel_data_in)? u0_col_out_359 : u1_col_out_359;
assign col_out_360 = (sel_data_in)? u0_col_out_360 : u1_col_out_360;
assign col_out_361 = (sel_data_in)? u0_col_out_361 : u1_col_out_361;
assign col_out_362 = (sel_data_in)? u0_col_out_362 : u1_col_out_362;
assign col_out_363 = (sel_data_in)? u0_col_out_363 : u1_col_out_363;
assign col_out_364 = (sel_data_in)? u0_col_out_364 : u1_col_out_364;
assign col_out_365 = (sel_data_in)? u0_col_out_365 : u1_col_out_365;
assign col_out_366 = (sel_data_in)? u0_col_out_366 : u1_col_out_366;
assign col_out_367 = (sel_data_in)? u0_col_out_367 : u1_col_out_367;
assign col_out_368 = (sel_data_in)? u0_col_out_368 : u1_col_out_368;
assign col_out_369 = (sel_data_in)? u0_col_out_369 : u1_col_out_369;
assign col_out_370 = (sel_data_in)? u0_col_out_370 : u1_col_out_370;
assign col_out_371 = (sel_data_in)? u0_col_out_371 : u1_col_out_371;
assign col_out_372 = (sel_data_in)? u0_col_out_372 : u1_col_out_372;
assign col_out_373 = (sel_data_in)? u0_col_out_373 : u1_col_out_373;
assign col_out_374 = (sel_data_in)? u0_col_out_374 : u1_col_out_374;
assign col_out_375 = (sel_data_in)? u0_col_out_375 : u1_col_out_375;
assign col_out_376 = (sel_data_in)? u0_col_out_376 : u1_col_out_376;
assign col_out_377 = (sel_data_in)? u0_col_out_377 : u1_col_out_377;
assign col_out_378 = (sel_data_in)? u0_col_out_378 : u1_col_out_378;
assign col_out_379 = (sel_data_in)? u0_col_out_379 : u1_col_out_379;
assign col_out_380 = (sel_data_in)? u0_col_out_380 : u1_col_out_380;
assign col_out_381 = (sel_data_in)? u0_col_out_381 : u1_col_out_381;
assign col_out_382 = (sel_data_in)? u0_col_out_382 : u1_col_out_382;
assign col_out_383 = (sel_data_in)? u0_col_out_383 : u1_col_out_383;
assign col_out_384 = (sel_data_in)? u0_col_out_384 : u1_col_out_384;
assign col_out_385 = (sel_data_in)? u0_col_out_385 : u1_col_out_385;
assign col_out_386 = (sel_data_in)? u0_col_out_386 : u1_col_out_386;
assign col_out_387 = (sel_data_in)? u0_col_out_387 : u1_col_out_387;
assign col_out_388 = (sel_data_in)? u0_col_out_388 : u1_col_out_388;
assign col_out_389 = (sel_data_in)? u0_col_out_389 : u1_col_out_389;
assign col_out_390 = (sel_data_in)? u0_col_out_390 : u1_col_out_390;
assign col_out_391 = (sel_data_in)? u0_col_out_391 : u1_col_out_391;
assign col_out_392 = (sel_data_in)? u0_col_out_392 : u1_col_out_392;
assign col_out_393 = (sel_data_in)? u0_col_out_393 : u1_col_out_393;
assign col_out_394 = (sel_data_in)? u0_col_out_394 : u1_col_out_394;
assign col_out_395 = (sel_data_in)? u0_col_out_395 : u1_col_out_395;
assign col_out_396 = (sel_data_in)? u0_col_out_396 : u1_col_out_396;
assign col_out_397 = (sel_data_in)? u0_col_out_397 : u1_col_out_397;
assign col_out_398 = (sel_data_in)? u0_col_out_398 : u1_col_out_398;
assign col_out_399 = (sel_data_in)? u0_col_out_399 : u1_col_out_399;
assign col_out_400 = (sel_data_in)? u0_col_out_400 : u1_col_out_400;
assign col_out_401 = (sel_data_in)? u0_col_out_401 : u1_col_out_401;
assign col_out_402 = (sel_data_in)? u0_col_out_402 : u1_col_out_402;
assign col_out_403 = (sel_data_in)? u0_col_out_403 : u1_col_out_403;
assign col_out_404 = (sel_data_in)? u0_col_out_404 : u1_col_out_404;
assign col_out_405 = (sel_data_in)? u0_col_out_405 : u1_col_out_405;
assign col_out_406 = (sel_data_in)? u0_col_out_406 : u1_col_out_406;
assign col_out_407 = (sel_data_in)? u0_col_out_407 : u1_col_out_407;
assign col_out_408 = (sel_data_in)? u0_col_out_408 : u1_col_out_408;
assign col_out_409 = (sel_data_in)? u0_col_out_409 : u1_col_out_409;
assign col_out_410 = (sel_data_in)? u0_col_out_410 : u1_col_out_410;
assign col_out_411 = (sel_data_in)? u0_col_out_411 : u1_col_out_411;
assign col_out_412 = (sel_data_in)? u0_col_out_412 : u1_col_out_412;
assign col_out_413 = (sel_data_in)? u0_col_out_413 : u1_col_out_413;
assign col_out_414 = (sel_data_in)? u0_col_out_414 : u1_col_out_414;
assign col_out_415 = (sel_data_in)? u0_col_out_415 : u1_col_out_415;
assign col_out_416 = (sel_data_in)? u0_col_out_416 : u1_col_out_416;
assign col_out_417 = (sel_data_in)? u0_col_out_417 : u1_col_out_417;
assign col_out_418 = (sel_data_in)? u0_col_out_418 : u1_col_out_418;
assign col_out_419 = (sel_data_in)? u0_col_out_419 : u1_col_out_419;
assign col_out_420 = (sel_data_in)? u0_col_out_420 : u1_col_out_420;
assign col_out_421 = (sel_data_in)? u0_col_out_421 : u1_col_out_421;
assign col_out_422 = (sel_data_in)? u0_col_out_422 : u1_col_out_422;
assign col_out_423 = (sel_data_in)? u0_col_out_423 : u1_col_out_423;
assign col_out_424 = (sel_data_in)? u0_col_out_424 : u1_col_out_424;
assign col_out_425 = (sel_data_in)? u0_col_out_425 : u1_col_out_425;
assign col_out_426 = (sel_data_in)? u0_col_out_426 : u1_col_out_426;
assign col_out_427 = (sel_data_in)? u0_col_out_427 : u1_col_out_427;
assign col_out_428 = (sel_data_in)? u0_col_out_428 : u1_col_out_428;
assign col_out_429 = (sel_data_in)? u0_col_out_429 : u1_col_out_429;
assign col_out_430 = (sel_data_in)? u0_col_out_430 : u1_col_out_430;
assign col_out_431 = (sel_data_in)? u0_col_out_431 : u1_col_out_431;
assign col_out_432 = (sel_data_in)? u0_col_out_432 : u1_col_out_432;
assign col_out_433 = (sel_data_in)? u0_col_out_433 : u1_col_out_433;
assign col_out_434 = (sel_data_in)? u0_col_out_434 : u1_col_out_434;
assign col_out_435 = (sel_data_in)? u0_col_out_435 : u1_col_out_435;
assign col_out_436 = (sel_data_in)? u0_col_out_436 : u1_col_out_436;
assign col_out_437 = (sel_data_in)? u0_col_out_437 : u1_col_out_437;
assign col_out_438 = (sel_data_in)? u0_col_out_438 : u1_col_out_438;
assign col_out_439 = (sel_data_in)? u0_col_out_439 : u1_col_out_439;
assign col_out_440 = (sel_data_in)? u0_col_out_440 : u1_col_out_440;
assign col_out_441 = (sel_data_in)? u0_col_out_441 : u1_col_out_441;
assign col_out_442 = (sel_data_in)? u0_col_out_442 : u1_col_out_442;
assign col_out_443 = (sel_data_in)? u0_col_out_443 : u1_col_out_443;
assign col_out_444 = (sel_data_in)? u0_col_out_444 : u1_col_out_444;
assign col_out_445 = (sel_data_in)? u0_col_out_445 : u1_col_out_445;
assign col_out_446 = (sel_data_in)? u0_col_out_446 : u1_col_out_446;
assign col_out_447 = (sel_data_in)? u0_col_out_447 : u1_col_out_447;
assign col_out_448 = (sel_data_in)? u0_col_out_448 : u1_col_out_448;
assign col_out_449 = (sel_data_in)? u0_col_out_449 : u1_col_out_449;
assign col_out_450 = (sel_data_in)? u0_col_out_450 : u1_col_out_450;
assign col_out_451 = (sel_data_in)? u0_col_out_451 : u1_col_out_451;
assign col_out_452 = (sel_data_in)? u0_col_out_452 : u1_col_out_452;
assign col_out_453 = (sel_data_in)? u0_col_out_453 : u1_col_out_453;
assign col_out_454 = (sel_data_in)? u0_col_out_454 : u1_col_out_454;
assign col_out_455 = (sel_data_in)? u0_col_out_455 : u1_col_out_455;
assign col_out_456 = (sel_data_in)? u0_col_out_456 : u1_col_out_456;
assign col_out_457 = (sel_data_in)? u0_col_out_457 : u1_col_out_457;
assign col_out_458 = (sel_data_in)? u0_col_out_458 : u1_col_out_458;
assign col_out_459 = (sel_data_in)? u0_col_out_459 : u1_col_out_459;
assign col_out_460 = (sel_data_in)? u0_col_out_460 : u1_col_out_460;
assign col_out_461 = (sel_data_in)? u0_col_out_461 : u1_col_out_461;
assign col_out_462 = (sel_data_in)? u0_col_out_462 : u1_col_out_462;
assign col_out_463 = (sel_data_in)? u0_col_out_463 : u1_col_out_463;
assign col_out_464 = (sel_data_in)? u0_col_out_464 : u1_col_out_464;
assign col_out_465 = (sel_data_in)? u0_col_out_465 : u1_col_out_465;
assign col_out_466 = (sel_data_in)? u0_col_out_466 : u1_col_out_466;
assign col_out_467 = (sel_data_in)? u0_col_out_467 : u1_col_out_467;
assign col_out_468 = (sel_data_in)? u0_col_out_468 : u1_col_out_468;
assign col_out_469 = (sel_data_in)? u0_col_out_469 : u1_col_out_469;
assign col_out_470 = (sel_data_in)? u0_col_out_470 : u1_col_out_470;
assign col_out_471 = (sel_data_in)? u0_col_out_471 : u1_col_out_471;
assign col_out_472 = (sel_data_in)? u0_col_out_472 : u1_col_out_472;
assign col_out_473 = (sel_data_in)? u0_col_out_473 : u1_col_out_473;
assign col_out_474 = (sel_data_in)? u0_col_out_474 : u1_col_out_474;
assign col_out_475 = (sel_data_in)? u0_col_out_475 : u1_col_out_475;
assign col_out_476 = (sel_data_in)? u0_col_out_476 : u1_col_out_476;
assign col_out_477 = (sel_data_in)? u0_col_out_477 : u1_col_out_477;
assign col_out_478 = (sel_data_in)? u0_col_out_478 : u1_col_out_478;
assign col_out_479 = (sel_data_in)? u0_col_out_479 : u1_col_out_479;
assign col_out_480 = (sel_data_in)? u0_col_out_480 : u1_col_out_480;
assign col_out_481 = (sel_data_in)? u0_col_out_481 : u1_col_out_481;
assign col_out_482 = (sel_data_in)? u0_col_out_482 : u1_col_out_482;
assign col_out_483 = (sel_data_in)? u0_col_out_483 : u1_col_out_483;
assign col_out_484 = (sel_data_in)? u0_col_out_484 : u1_col_out_484;
assign col_out_485 = (sel_data_in)? u0_col_out_485 : u1_col_out_485;
assign col_out_486 = (sel_data_in)? u0_col_out_486 : u1_col_out_486;
assign col_out_487 = (sel_data_in)? u0_col_out_487 : u1_col_out_487;
assign col_out_488 = (sel_data_in)? u0_col_out_488 : u1_col_out_488;
assign col_out_489 = (sel_data_in)? u0_col_out_489 : u1_col_out_489;
assign col_out_490 = (sel_data_in)? u0_col_out_490 : u1_col_out_490;
assign col_out_491 = (sel_data_in)? u0_col_out_491 : u1_col_out_491;
assign col_out_492 = (sel_data_in)? u0_col_out_492 : u1_col_out_492;
assign col_out_493 = (sel_data_in)? u0_col_out_493 : u1_col_out_493;
assign col_out_494 = (sel_data_in)? u0_col_out_494 : u1_col_out_494;
assign col_out_495 = (sel_data_in)? u0_col_out_495 : u1_col_out_495;
assign col_out_496 = (sel_data_in)? u0_col_out_496 : u1_col_out_496;
assign col_out_497 = (sel_data_in)? u0_col_out_497 : u1_col_out_497;
assign col_out_498 = (sel_data_in)? u0_col_out_498 : u1_col_out_498;
assign col_out_499 = (sel_data_in)? u0_col_out_499 : u1_col_out_499;
assign col_out_500 = (sel_data_in)? u0_col_out_500 : u1_col_out_500;
assign col_out_501 = (sel_data_in)? u0_col_out_501 : u1_col_out_501;
assign col_out_502 = (sel_data_in)? u0_col_out_502 : u1_col_out_502;
assign col_out_503 = (sel_data_in)? u0_col_out_503 : u1_col_out_503;
assign col_out_504 = (sel_data_in)? u0_col_out_504 : u1_col_out_504;
assign col_out_505 = (sel_data_in)? u0_col_out_505 : u1_col_out_505;
assign col_out_506 = (sel_data_in)? u0_col_out_506 : u1_col_out_506;
assign col_out_507 = (sel_data_in)? u0_col_out_507 : u1_col_out_507;
assign col_out_508 = (sel_data_in)? u0_col_out_508 : u1_col_out_508;
assign col_out_509 = (sel_data_in)? u0_col_out_509 : u1_col_out_509;
assign col_out_510 = (sel_data_in)? u0_col_out_510 : u1_col_out_510;
assign col_out_511 = (sel_data_in)? u0_col_out_511 : u1_col_out_511;
assign col_out_512 = (sel_data_in)? u0_col_out_512 : u1_col_out_512;
assign col_out_513 = (sel_data_in)? u0_col_out_513 : u1_col_out_513;
assign col_out_514 = (sel_data_in)? u0_col_out_514 : u1_col_out_514;
assign col_out_515 = (sel_data_in)? u0_col_out_515 : u1_col_out_515;
assign col_out_516 = (sel_data_in)? u0_col_out_516 : u1_col_out_516;
assign col_out_517 = (sel_data_in)? u0_col_out_517 : u1_col_out_517;
assign col_out_518 = (sel_data_in)? u0_col_out_518 : u1_col_out_518;
assign col_out_519 = (sel_data_in)? u0_col_out_519 : u1_col_out_519;
assign col_out_520 = (sel_data_in)? u0_col_out_520 : u1_col_out_520;
assign col_out_521 = (sel_data_in)? u0_col_out_521 : u1_col_out_521;
assign col_out_522 = (sel_data_in)? u0_col_out_522 : u1_col_out_522;
assign col_out_523 = (sel_data_in)? u0_col_out_523 : u1_col_out_523;
assign col_out_524 = (sel_data_in)? u0_col_out_524 : u1_col_out_524;
assign col_out_525 = (sel_data_in)? u0_col_out_525 : u1_col_out_525;
assign col_out_526 = (sel_data_in)? u0_col_out_526 : u1_col_out_526;
assign col_out_527 = (sel_data_in)? u0_col_out_527 : u1_col_out_527;
assign col_out_528 = (sel_data_in)? u0_col_out_528 : u1_col_out_528;
assign col_out_529 = (sel_data_in)? u0_col_out_529 : u1_col_out_529;
assign col_out_530 = (sel_data_in)? u0_col_out_530 : u1_col_out_530;
assign col_out_531 = (sel_data_in)? u0_col_out_531 : u1_col_out_531;
assign col_out_532 = (sel_data_in)? u0_col_out_532 : u1_col_out_532;
assign col_out_533 = (sel_data_in)? u0_col_out_533 : u1_col_out_533;
assign col_out_534 = (sel_data_in)? u0_col_out_534 : u1_col_out_534;
assign col_out_535 = (sel_data_in)? u0_col_out_535 : u1_col_out_535;
assign col_out_536 = (sel_data_in)? u0_col_out_536 : u1_col_out_536;
assign col_out_537 = (sel_data_in)? u0_col_out_537 : u1_col_out_537;
assign col_out_538 = (sel_data_in)? u0_col_out_538 : u1_col_out_538;
assign col_out_539 = (sel_data_in)? u0_col_out_539 : u1_col_out_539;
assign col_out_540 = (sel_data_in)? u0_col_out_540 : u1_col_out_540;
assign col_out_541 = (sel_data_in)? u0_col_out_541 : u1_col_out_541;
assign col_out_542 = (sel_data_in)? u0_col_out_542 : u1_col_out_542;
assign col_out_543 = (sel_data_in)? u0_col_out_543 : u1_col_out_543;
assign col_out_544 = (sel_data_in)? u0_col_out_544 : u1_col_out_544;
assign col_out_545 = (sel_data_in)? u0_col_out_545 : u1_col_out_545;
assign col_out_546 = (sel_data_in)? u0_col_out_546 : u1_col_out_546;
assign col_out_547 = (sel_data_in)? u0_col_out_547 : u1_col_out_547;
assign col_out_548 = (sel_data_in)? u0_col_out_548 : u1_col_out_548;
assign col_out_549 = (sel_data_in)? u0_col_out_549 : u1_col_out_549;
assign col_out_550 = (sel_data_in)? u0_col_out_550 : u1_col_out_550;
assign col_out_551 = (sel_data_in)? u0_col_out_551 : u1_col_out_551;
assign col_out_552 = (sel_data_in)? u0_col_out_552 : u1_col_out_552;
assign col_out_553 = (sel_data_in)? u0_col_out_553 : u1_col_out_553;
assign col_out_554 = (sel_data_in)? u0_col_out_554 : u1_col_out_554;
assign col_out_555 = (sel_data_in)? u0_col_out_555 : u1_col_out_555;
assign col_out_556 = (sel_data_in)? u0_col_out_556 : u1_col_out_556;
assign col_out_557 = (sel_data_in)? u0_col_out_557 : u1_col_out_557;
assign col_out_558 = (sel_data_in)? u0_col_out_558 : u1_col_out_558;
assign col_out_559 = (sel_data_in)? u0_col_out_559 : u1_col_out_559;
assign col_out_560 = (sel_data_in)? u0_col_out_560 : u1_col_out_560;
assign col_out_561 = (sel_data_in)? u0_col_out_561 : u1_col_out_561;
assign col_out_562 = (sel_data_in)? u0_col_out_562 : u1_col_out_562;
assign col_out_563 = (sel_data_in)? u0_col_out_563 : u1_col_out_563;
assign col_out_564 = (sel_data_in)? u0_col_out_564 : u1_col_out_564;
assign col_out_565 = (sel_data_in)? u0_col_out_565 : u1_col_out_565;
assign col_out_566 = (sel_data_in)? u0_col_out_566 : u1_col_out_566;
assign col_out_567 = (sel_data_in)? u0_col_out_567 : u1_col_out_567;
assign col_out_568 = (sel_data_in)? u0_col_out_568 : u1_col_out_568;
assign col_out_569 = (sel_data_in)? u0_col_out_569 : u1_col_out_569;
assign col_out_570 = (sel_data_in)? u0_col_out_570 : u1_col_out_570;
assign col_out_571 = (sel_data_in)? u0_col_out_571 : u1_col_out_571;
assign col_out_572 = (sel_data_in)? u0_col_out_572 : u1_col_out_572;
assign col_out_573 = (sel_data_in)? u0_col_out_573 : u1_col_out_573;
assign col_out_574 = (sel_data_in)? u0_col_out_574 : u1_col_out_574;
assign col_out_575 = (sel_data_in)? u0_col_out_575 : u1_col_out_575;
assign col_out_576 = (sel_data_in)? u0_col_out_576 : u1_col_out_576;
assign col_out_577 = (sel_data_in)? u0_col_out_577 : u1_col_out_577;
assign col_out_578 = (sel_data_in)? u0_col_out_578 : u1_col_out_578;
assign col_out_579 = (sel_data_in)? u0_col_out_579 : u1_col_out_579;
assign col_out_580 = (sel_data_in)? u0_col_out_580 : u1_col_out_580;
assign col_out_581 = (sel_data_in)? u0_col_out_581 : u1_col_out_581;
assign col_out_582 = (sel_data_in)? u0_col_out_582 : u1_col_out_582;
assign col_out_583 = (sel_data_in)? u0_col_out_583 : u1_col_out_583;
assign col_out_584 = (sel_data_in)? u0_col_out_584 : u1_col_out_584;
assign col_out_585 = (sel_data_in)? u0_col_out_585 : u1_col_out_585;
assign col_out_586 = (sel_data_in)? u0_col_out_586 : u1_col_out_586;
assign col_out_587 = (sel_data_in)? u0_col_out_587 : u1_col_out_587;
assign col_out_588 = (sel_data_in)? u0_col_out_588 : u1_col_out_588;
assign col_out_589 = (sel_data_in)? u0_col_out_589 : u1_col_out_589;
assign col_out_590 = (sel_data_in)? u0_col_out_590 : u1_col_out_590;
assign col_out_591 = (sel_data_in)? u0_col_out_591 : u1_col_out_591;
assign col_out_592 = (sel_data_in)? u0_col_out_592 : u1_col_out_592;
assign col_out_593 = (sel_data_in)? u0_col_out_593 : u1_col_out_593;
assign col_out_594 = (sel_data_in)? u0_col_out_594 : u1_col_out_594;
assign col_out_595 = (sel_data_in)? u0_col_out_595 : u1_col_out_595;
assign col_out_596 = (sel_data_in)? u0_col_out_596 : u1_col_out_596;
assign col_out_597 = (sel_data_in)? u0_col_out_597 : u1_col_out_597;
assign col_out_598 = (sel_data_in)? u0_col_out_598 : u1_col_out_598;
assign col_out_599 = (sel_data_in)? u0_col_out_599 : u1_col_out_599;
assign col_out_600 = (sel_data_in)? u0_col_out_600 : u1_col_out_600;
assign col_out_601 = (sel_data_in)? u0_col_out_601 : u1_col_out_601;
assign col_out_602 = (sel_data_in)? u0_col_out_602 : u1_col_out_602;
assign col_out_603 = (sel_data_in)? u0_col_out_603 : u1_col_out_603;
assign col_out_604 = (sel_data_in)? u0_col_out_604 : u1_col_out_604;
assign col_out_605 = (sel_data_in)? u0_col_out_605 : u1_col_out_605;
assign col_out_606 = (sel_data_in)? u0_col_out_606 : u1_col_out_606;
assign col_out_607 = (sel_data_in)? u0_col_out_607 : u1_col_out_607;
assign col_out_608 = (sel_data_in)? u0_col_out_608 : u1_col_out_608;
assign col_out_609 = (sel_data_in)? u0_col_out_609 : u1_col_out_609;
assign col_out_610 = (sel_data_in)? u0_col_out_610 : u1_col_out_610;
assign col_out_611 = (sel_data_in)? u0_col_out_611 : u1_col_out_611;
assign col_out_612 = (sel_data_in)? u0_col_out_612 : u1_col_out_612;
assign col_out_613 = (sel_data_in)? u0_col_out_613 : u1_col_out_613;
assign col_out_614 = (sel_data_in)? u0_col_out_614 : u1_col_out_614;
assign col_out_615 = (sel_data_in)? u0_col_out_615 : u1_col_out_615;
assign col_out_616 = (sel_data_in)? u0_col_out_616 : u1_col_out_616;
assign col_out_617 = (sel_data_in)? u0_col_out_617 : u1_col_out_617;
assign col_out_618 = (sel_data_in)? u0_col_out_618 : u1_col_out_618;
assign col_out_619 = (sel_data_in)? u0_col_out_619 : u1_col_out_619;
assign col_out_620 = (sel_data_in)? u0_col_out_620 : u1_col_out_620;
assign col_out_621 = (sel_data_in)? u0_col_out_621 : u1_col_out_621;
assign col_out_622 = (sel_data_in)? u0_col_out_622 : u1_col_out_622;
assign col_out_623 = (sel_data_in)? u0_col_out_623 : u1_col_out_623;
assign col_out_624 = (sel_data_in)? u0_col_out_624 : u1_col_out_624;
assign col_out_625 = (sel_data_in)? u0_col_out_625 : u1_col_out_625;
assign col_out_626 = (sel_data_in)? u0_col_out_626 : u1_col_out_626;
assign col_out_627 = (sel_data_in)? u0_col_out_627 : u1_col_out_627;
assign col_out_628 = (sel_data_in)? u0_col_out_628 : u1_col_out_628;
assign col_out_629 = (sel_data_in)? u0_col_out_629 : u1_col_out_629;
assign col_out_630 = (sel_data_in)? u0_col_out_630 : u1_col_out_630;
assign col_out_631 = (sel_data_in)? u0_col_out_631 : u1_col_out_631;
assign col_out_632 = (sel_data_in)? u0_col_out_632 : u1_col_out_632;
assign col_out_633 = (sel_data_in)? u0_col_out_633 : u1_col_out_633;
assign col_out_634 = (sel_data_in)? u0_col_out_634 : u1_col_out_634;
assign col_out_635 = (sel_data_in)? u0_col_out_635 : u1_col_out_635;
assign col_out_636 = (sel_data_in)? u0_col_out_636 : u1_col_out_636;
assign col_out_637 = (sel_data_in)? u0_col_out_637 : u1_col_out_637;
assign col_out_638 = (sel_data_in)? u0_col_out_638 : u1_col_out_638;
assign col_out_639 = (sel_data_in)? u0_col_out_639 : u1_col_out_639;
assign col_out_640 = (sel_data_in)? u0_col_out_640 : u1_col_out_640;
assign col_out_641 = (sel_data_in)? u0_col_out_641 : u1_col_out_641;
assign col_out_642 = (sel_data_in)? u0_col_out_642 : u1_col_out_642;
assign col_out_643 = (sel_data_in)? u0_col_out_643 : u1_col_out_643;
assign col_out_644 = (sel_data_in)? u0_col_out_644 : u1_col_out_644;
assign col_out_645 = (sel_data_in)? u0_col_out_645 : u1_col_out_645;
assign col_out_646 = (sel_data_in)? u0_col_out_646 : u1_col_out_646;
assign col_out_647 = (sel_data_in)? u0_col_out_647 : u1_col_out_647;
assign col_out_648 = (sel_data_in)? u0_col_out_648 : u1_col_out_648;
assign col_out_649 = (sel_data_in)? u0_col_out_649 : u1_col_out_649;
assign col_out_650 = (sel_data_in)? u0_col_out_650 : u1_col_out_650;
assign col_out_651 = (sel_data_in)? u0_col_out_651 : u1_col_out_651;
assign col_out_652 = (sel_data_in)? u0_col_out_652 : u1_col_out_652;
assign col_out_653 = (sel_data_in)? u0_col_out_653 : u1_col_out_653;
assign col_out_654 = (sel_data_in)? u0_col_out_654 : u1_col_out_654;
assign col_out_655 = (sel_data_in)? u0_col_out_655 : u1_col_out_655;
assign col_out_656 = (sel_data_in)? u0_col_out_656 : u1_col_out_656;
assign col_out_657 = (sel_data_in)? u0_col_out_657 : u1_col_out_657;
assign col_out_658 = (sel_data_in)? u0_col_out_658 : u1_col_out_658;
assign col_out_659 = (sel_data_in)? u0_col_out_659 : u1_col_out_659;
assign col_out_660 = (sel_data_in)? u0_col_out_660 : u1_col_out_660;
assign col_out_661 = (sel_data_in)? u0_col_out_661 : u1_col_out_661;
assign col_out_662 = (sel_data_in)? u0_col_out_662 : u1_col_out_662;
assign col_out_663 = (sel_data_in)? u0_col_out_663 : u1_col_out_663;
assign col_out_664 = (sel_data_in)? u0_col_out_664 : u1_col_out_664;
assign col_out_665 = (sel_data_in)? u0_col_out_665 : u1_col_out_665;
assign col_out_666 = (sel_data_in)? u0_col_out_666 : u1_col_out_666;
assign col_out_667 = (sel_data_in)? u0_col_out_667 : u1_col_out_667;
assign col_out_668 = (sel_data_in)? u0_col_out_668 : u1_col_out_668;
assign col_out_669 = (sel_data_in)? u0_col_out_669 : u1_col_out_669;
assign col_out_670 = (sel_data_in)? u0_col_out_670 : u1_col_out_670;
assign col_out_671 = (sel_data_in)? u0_col_out_671 : u1_col_out_671;
assign col_out_672 = (sel_data_in)? u0_col_out_672 : u1_col_out_672;
assign col_out_673 = (sel_data_in)? u0_col_out_673 : u1_col_out_673;
assign col_out_674 = (sel_data_in)? u0_col_out_674 : u1_col_out_674;
assign col_out_675 = (sel_data_in)? u0_col_out_675 : u1_col_out_675;
assign col_out_676 = (sel_data_in)? u0_col_out_676 : u1_col_out_676;
assign col_out_677 = (sel_data_in)? u0_col_out_677 : u1_col_out_677;
assign col_out_678 = (sel_data_in)? u0_col_out_678 : u1_col_out_678;
assign col_out_679 = (sel_data_in)? u0_col_out_679 : u1_col_out_679;
assign col_out_680 = (sel_data_in)? u0_col_out_680 : u1_col_out_680;
assign col_out_681 = (sel_data_in)? u0_col_out_681 : u1_col_out_681;
assign col_out_682 = (sel_data_in)? u0_col_out_682 : u1_col_out_682;
assign col_out_683 = (sel_data_in)? u0_col_out_683 : u1_col_out_683;
assign col_out_684 = (sel_data_in)? u0_col_out_684 : u1_col_out_684;
assign col_out_685 = (sel_data_in)? u0_col_out_685 : u1_col_out_685;
assign col_out_686 = (sel_data_in)? u0_col_out_686 : u1_col_out_686;
assign col_out_687 = (sel_data_in)? u0_col_out_687 : u1_col_out_687;
assign col_out_688 = (sel_data_in)? u0_col_out_688 : u1_col_out_688;
assign col_out_689 = (sel_data_in)? u0_col_out_689 : u1_col_out_689;
assign col_out_690 = (sel_data_in)? u0_col_out_690 : u1_col_out_690;
assign col_out_691 = (sel_data_in)? u0_col_out_691 : u1_col_out_691;
assign col_out_692 = (sel_data_in)? u0_col_out_692 : u1_col_out_692;
assign col_out_693 = (sel_data_in)? u0_col_out_693 : u1_col_out_693;
assign col_out_694 = (sel_data_in)? u0_col_out_694 : u1_col_out_694;
assign col_out_695 = (sel_data_in)? u0_col_out_695 : u1_col_out_695;
assign col_out_696 = (sel_data_in)? u0_col_out_696 : u1_col_out_696;
assign col_out_697 = (sel_data_in)? u0_col_out_697 : u1_col_out_697;
assign col_out_698 = (sel_data_in)? u0_col_out_698 : u1_col_out_698;
assign col_out_699 = (sel_data_in)? u0_col_out_699 : u1_col_out_699;
assign col_out_700 = (sel_data_in)? u0_col_out_700 : u1_col_out_700;
assign col_out_701 = (sel_data_in)? u0_col_out_701 : u1_col_out_701;
assign col_out_702 = (sel_data_in)? u0_col_out_702 : u1_col_out_702;
assign col_out_703 = (sel_data_in)? u0_col_out_703 : u1_col_out_703;
assign col_out_704 = (sel_data_in)? u0_col_out_704 : u1_col_out_704;
assign col_out_705 = (sel_data_in)? u0_col_out_705 : u1_col_out_705;
assign col_out_706 = (sel_data_in)? u0_col_out_706 : u1_col_out_706;
assign col_out_707 = (sel_data_in)? u0_col_out_707 : u1_col_out_707;
assign col_out_708 = (sel_data_in)? u0_col_out_708 : u1_col_out_708;
assign col_out_709 = (sel_data_in)? u0_col_out_709 : u1_col_out_709;
assign col_out_710 = (sel_data_in)? u0_col_out_710 : u1_col_out_710;
assign col_out_711 = (sel_data_in)? u0_col_out_711 : u1_col_out_711;
assign col_out_712 = (sel_data_in)? u0_col_out_712 : u1_col_out_712;
assign col_out_713 = (sel_data_in)? u0_col_out_713 : u1_col_out_713;
assign col_out_714 = (sel_data_in)? u0_col_out_714 : u1_col_out_714;
assign col_out_715 = (sel_data_in)? u0_col_out_715 : u1_col_out_715;
assign col_out_716 = (sel_data_in)? u0_col_out_716 : u1_col_out_716;
assign col_out_717 = (sel_data_in)? u0_col_out_717 : u1_col_out_717;
assign col_out_718 = (sel_data_in)? u0_col_out_718 : u1_col_out_718;
assign col_out_719 = (sel_data_in)? u0_col_out_719 : u1_col_out_719;
assign col_out_720 = (sel_data_in)? u0_col_out_720 : u1_col_out_720;
assign col_out_721 = (sel_data_in)? u0_col_out_721 : u1_col_out_721;
assign col_out_722 = (sel_data_in)? u0_col_out_722 : u1_col_out_722;
assign col_out_723 = (sel_data_in)? u0_col_out_723 : u1_col_out_723;
assign col_out_724 = (sel_data_in)? u0_col_out_724 : u1_col_out_724;
assign col_out_725 = (sel_data_in)? u0_col_out_725 : u1_col_out_725;
assign col_out_726 = (sel_data_in)? u0_col_out_726 : u1_col_out_726;
assign col_out_727 = (sel_data_in)? u0_col_out_727 : u1_col_out_727;
assign col_out_728 = (sel_data_in)? u0_col_out_728 : u1_col_out_728;
assign col_out_729 = (sel_data_in)? u0_col_out_729 : u1_col_out_729;
assign col_out_730 = (sel_data_in)? u0_col_out_730 : u1_col_out_730;
assign col_out_731 = (sel_data_in)? u0_col_out_731 : u1_col_out_731;
assign col_out_732 = (sel_data_in)? u0_col_out_732 : u1_col_out_732;
assign col_out_733 = (sel_data_in)? u0_col_out_733 : u1_col_out_733;
assign col_out_734 = (sel_data_in)? u0_col_out_734 : u1_col_out_734;
assign col_out_735 = (sel_data_in)? u0_col_out_735 : u1_col_out_735;
assign col_out_736 = (sel_data_in)? u0_col_out_736 : u1_col_out_736;
assign col_out_737 = (sel_data_in)? u0_col_out_737 : u1_col_out_737;
assign col_out_738 = (sel_data_in)? u0_col_out_738 : u1_col_out_738;
assign col_out_739 = (sel_data_in)? u0_col_out_739 : u1_col_out_739;
assign col_out_740 = (sel_data_in)? u0_col_out_740 : u1_col_out_740;
assign col_out_741 = (sel_data_in)? u0_col_out_741 : u1_col_out_741;
assign col_out_742 = (sel_data_in)? u0_col_out_742 : u1_col_out_742;
assign col_out_743 = (sel_data_in)? u0_col_out_743 : u1_col_out_743;
assign col_out_744 = (sel_data_in)? u0_col_out_744 : u1_col_out_744;
assign col_out_745 = (sel_data_in)? u0_col_out_745 : u1_col_out_745;
assign col_out_746 = (sel_data_in)? u0_col_out_746 : u1_col_out_746;
assign col_out_747 = (sel_data_in)? u0_col_out_747 : u1_col_out_747;
assign col_out_748 = (sel_data_in)? u0_col_out_748 : u1_col_out_748;
assign col_out_749 = (sel_data_in)? u0_col_out_749 : u1_col_out_749;
assign col_out_750 = (sel_data_in)? u0_col_out_750 : u1_col_out_750;
assign col_out_751 = (sel_data_in)? u0_col_out_751 : u1_col_out_751;
assign col_out_752 = (sel_data_in)? u0_col_out_752 : u1_col_out_752;
assign col_out_753 = (sel_data_in)? u0_col_out_753 : u1_col_out_753;
assign col_out_754 = (sel_data_in)? u0_col_out_754 : u1_col_out_754;
assign col_out_755 = (sel_data_in)? u0_col_out_755 : u1_col_out_755;
assign col_out_756 = (sel_data_in)? u0_col_out_756 : u1_col_out_756;
assign col_out_757 = (sel_data_in)? u0_col_out_757 : u1_col_out_757;
assign col_out_758 = (sel_data_in)? u0_col_out_758 : u1_col_out_758;
assign col_out_759 = (sel_data_in)? u0_col_out_759 : u1_col_out_759;
assign col_out_760 = (sel_data_in)? u0_col_out_760 : u1_col_out_760;
assign col_out_761 = (sel_data_in)? u0_col_out_761 : u1_col_out_761;
assign col_out_762 = (sel_data_in)? u0_col_out_762 : u1_col_out_762;
assign col_out_763 = (sel_data_in)? u0_col_out_763 : u1_col_out_763;
assign col_out_764 = (sel_data_in)? u0_col_out_764 : u1_col_out_764;
assign col_out_765 = (sel_data_in)? u0_col_out_765 : u1_col_out_765;
assign col_out_766 = (sel_data_in)? u0_col_out_766 : u1_col_out_766;
assign col_out_767 = (sel_data_in)? u0_col_out_767 : u1_col_out_767;
assign col_out_768 = (sel_data_in)? u0_col_out_768 : u1_col_out_768;
assign col_out_769 = (sel_data_in)? u0_col_out_769 : u1_col_out_769;
assign col_out_770 = (sel_data_in)? u0_col_out_770 : u1_col_out_770;
assign col_out_771 = (sel_data_in)? u0_col_out_771 : u1_col_out_771;
assign col_out_772 = (sel_data_in)? u0_col_out_772 : u1_col_out_772;
assign col_out_773 = (sel_data_in)? u0_col_out_773 : u1_col_out_773;
assign col_out_774 = (sel_data_in)? u0_col_out_774 : u1_col_out_774;
assign col_out_775 = (sel_data_in)? u0_col_out_775 : u1_col_out_775;
assign col_out_776 = (sel_data_in)? u0_col_out_776 : u1_col_out_776;
assign col_out_777 = (sel_data_in)? u0_col_out_777 : u1_col_out_777;
assign col_out_778 = (sel_data_in)? u0_col_out_778 : u1_col_out_778;
assign col_out_779 = (sel_data_in)? u0_col_out_779 : u1_col_out_779;
assign col_out_780 = (sel_data_in)? u0_col_out_780 : u1_col_out_780;
assign col_out_781 = (sel_data_in)? u0_col_out_781 : u1_col_out_781;
assign col_out_782 = (sel_data_in)? u0_col_out_782 : u1_col_out_782;
assign col_out_783 = (sel_data_in)? u0_col_out_783 : u1_col_out_783;
assign col_out_784 = (sel_data_in)? u0_col_out_784 : u1_col_out_784;
assign col_out_785 = (sel_data_in)? u0_col_out_785 : u1_col_out_785;
assign col_out_786 = (sel_data_in)? u0_col_out_786 : u1_col_out_786;
assign col_out_787 = (sel_data_in)? u0_col_out_787 : u1_col_out_787;
assign col_out_788 = (sel_data_in)? u0_col_out_788 : u1_col_out_788;
assign col_out_789 = (sel_data_in)? u0_col_out_789 : u1_col_out_789;
assign col_out_790 = (sel_data_in)? u0_col_out_790 : u1_col_out_790;
assign col_out_791 = (sel_data_in)? u0_col_out_791 : u1_col_out_791;
assign col_out_792 = (sel_data_in)? u0_col_out_792 : u1_col_out_792;
assign col_out_793 = (sel_data_in)? u0_col_out_793 : u1_col_out_793;
assign col_out_794 = (sel_data_in)? u0_col_out_794 : u1_col_out_794;
assign col_out_795 = (sel_data_in)? u0_col_out_795 : u1_col_out_795;
assign col_out_796 = (sel_data_in)? u0_col_out_796 : u1_col_out_796;
assign col_out_797 = (sel_data_in)? u0_col_out_797 : u1_col_out_797;
assign col_out_798 = (sel_data_in)? u0_col_out_798 : u1_col_out_798;
assign col_out_799 = (sel_data_in)? u0_col_out_799 : u1_col_out_799;
assign col_out_800 = (sel_data_in)? u0_col_out_800 : u1_col_out_800;
assign col_out_801 = (sel_data_in)? u0_col_out_801 : u1_col_out_801;
assign col_out_802 = (sel_data_in)? u0_col_out_802 : u1_col_out_802;
assign col_out_803 = (sel_data_in)? u0_col_out_803 : u1_col_out_803;
assign col_out_804 = (sel_data_in)? u0_col_out_804 : u1_col_out_804;
assign col_out_805 = (sel_data_in)? u0_col_out_805 : u1_col_out_805;
assign col_out_806 = (sel_data_in)? u0_col_out_806 : u1_col_out_806;
assign col_out_807 = (sel_data_in)? u0_col_out_807 : u1_col_out_807;
assign col_out_808 = (sel_data_in)? u0_col_out_808 : u1_col_out_808;
assign col_out_809 = (sel_data_in)? u0_col_out_809 : u1_col_out_809;
assign col_out_810 = (sel_data_in)? u0_col_out_810 : u1_col_out_810;
assign col_out_811 = (sel_data_in)? u0_col_out_811 : u1_col_out_811;
assign col_out_812 = (sel_data_in)? u0_col_out_812 : u1_col_out_812;
assign col_out_813 = (sel_data_in)? u0_col_out_813 : u1_col_out_813;
assign col_out_814 = (sel_data_in)? u0_col_out_814 : u1_col_out_814;
assign col_out_815 = (sel_data_in)? u0_col_out_815 : u1_col_out_815;
assign col_out_816 = (sel_data_in)? u0_col_out_816 : u1_col_out_816;
assign col_out_817 = (sel_data_in)? u0_col_out_817 : u1_col_out_817;
assign col_out_818 = (sel_data_in)? u0_col_out_818 : u1_col_out_818;
assign col_out_819 = (sel_data_in)? u0_col_out_819 : u1_col_out_819;
assign col_out_820 = (sel_data_in)? u0_col_out_820 : u1_col_out_820;
assign col_out_821 = (sel_data_in)? u0_col_out_821 : u1_col_out_821;
assign col_out_822 = (sel_data_in)? u0_col_out_822 : u1_col_out_822;
assign col_out_823 = (sel_data_in)? u0_col_out_823 : u1_col_out_823;
assign col_out_824 = (sel_data_in)? u0_col_out_824 : u1_col_out_824;
assign col_out_825 = (sel_data_in)? u0_col_out_825 : u1_col_out_825;
assign col_out_826 = (sel_data_in)? u0_col_out_826 : u1_col_out_826;
assign col_out_827 = (sel_data_in)? u0_col_out_827 : u1_col_out_827;
assign col_out_828 = (sel_data_in)? u0_col_out_828 : u1_col_out_828;
assign col_out_829 = (sel_data_in)? u0_col_out_829 : u1_col_out_829;
assign col_out_830 = (sel_data_in)? u0_col_out_830 : u1_col_out_830;
assign col_out_831 = (sel_data_in)? u0_col_out_831 : u1_col_out_831;
assign col_out_832 = (sel_data_in)? u0_col_out_832 : u1_col_out_832;
assign col_out_833 = (sel_data_in)? u0_col_out_833 : u1_col_out_833;
assign col_out_834 = (sel_data_in)? u0_col_out_834 : u1_col_out_834;
assign col_out_835 = (sel_data_in)? u0_col_out_835 : u1_col_out_835;
assign col_out_836 = (sel_data_in)? u0_col_out_836 : u1_col_out_836;
assign col_out_837 = (sel_data_in)? u0_col_out_837 : u1_col_out_837;
assign col_out_838 = (sel_data_in)? u0_col_out_838 : u1_col_out_838;
assign col_out_839 = (sel_data_in)? u0_col_out_839 : u1_col_out_839;
assign col_out_840 = (sel_data_in)? u0_col_out_840 : u1_col_out_840;
assign col_out_841 = (sel_data_in)? u0_col_out_841 : u1_col_out_841;
assign col_out_842 = (sel_data_in)? u0_col_out_842 : u1_col_out_842;
assign col_out_843 = (sel_data_in)? u0_col_out_843 : u1_col_out_843;
assign col_out_844 = (sel_data_in)? u0_col_out_844 : u1_col_out_844;
assign col_out_845 = (sel_data_in)? u0_col_out_845 : u1_col_out_845;
assign col_out_846 = (sel_data_in)? u0_col_out_846 : u1_col_out_846;
assign col_out_847 = (sel_data_in)? u0_col_out_847 : u1_col_out_847;
assign col_out_848 = (sel_data_in)? u0_col_out_848 : u1_col_out_848;
assign col_out_849 = (sel_data_in)? u0_col_out_849 : u1_col_out_849;
assign col_out_850 = (sel_data_in)? u0_col_out_850 : u1_col_out_850;
assign col_out_851 = (sel_data_in)? u0_col_out_851 : u1_col_out_851;
assign col_out_852 = (sel_data_in)? u0_col_out_852 : u1_col_out_852;
assign col_out_853 = (sel_data_in)? u0_col_out_853 : u1_col_out_853;
assign col_out_854 = (sel_data_in)? u0_col_out_854 : u1_col_out_854;
assign col_out_855 = (sel_data_in)? u0_col_out_855 : u1_col_out_855;
assign col_out_856 = (sel_data_in)? u0_col_out_856 : u1_col_out_856;
assign col_out_857 = (sel_data_in)? u0_col_out_857 : u1_col_out_857;
assign col_out_858 = (sel_data_in)? u0_col_out_858 : u1_col_out_858;
assign col_out_859 = (sel_data_in)? u0_col_out_859 : u1_col_out_859;
assign col_out_860 = (sel_data_in)? u0_col_out_860 : u1_col_out_860;
assign col_out_861 = (sel_data_in)? u0_col_out_861 : u1_col_out_861;
assign col_out_862 = (sel_data_in)? u0_col_out_862 : u1_col_out_862;
assign col_out_863 = (sel_data_in)? u0_col_out_863 : u1_col_out_863;
assign col_out_864 = (sel_data_in)? u0_col_out_864 : u1_col_out_864;
assign col_out_865 = (sel_data_in)? u0_col_out_865 : u1_col_out_865;
assign col_out_866 = (sel_data_in)? u0_col_out_866 : u1_col_out_866;
assign col_out_867 = (sel_data_in)? u0_col_out_867 : u1_col_out_867;
assign col_out_868 = (sel_data_in)? u0_col_out_868 : u1_col_out_868;
assign col_out_869 = (sel_data_in)? u0_col_out_869 : u1_col_out_869;
assign col_out_870 = (sel_data_in)? u0_col_out_870 : u1_col_out_870;
assign col_out_871 = (sel_data_in)? u0_col_out_871 : u1_col_out_871;
assign col_out_872 = (sel_data_in)? u0_col_out_872 : u1_col_out_872;
assign col_out_873 = (sel_data_in)? u0_col_out_873 : u1_col_out_873;
assign col_out_874 = (sel_data_in)? u0_col_out_874 : u1_col_out_874;
assign col_out_875 = (sel_data_in)? u0_col_out_875 : u1_col_out_875;
assign col_out_876 = (sel_data_in)? u0_col_out_876 : u1_col_out_876;
assign col_out_877 = (sel_data_in)? u0_col_out_877 : u1_col_out_877;
assign col_out_878 = (sel_data_in)? u0_col_out_878 : u1_col_out_878;
assign col_out_879 = (sel_data_in)? u0_col_out_879 : u1_col_out_879;
assign col_out_880 = (sel_data_in)? u0_col_out_880 : u1_col_out_880;
assign col_out_881 = (sel_data_in)? u0_col_out_881 : u1_col_out_881;
assign col_out_882 = (sel_data_in)? u0_col_out_882 : u1_col_out_882;
assign col_out_883 = (sel_data_in)? u0_col_out_883 : u1_col_out_883;
assign col_out_884 = (sel_data_in)? u0_col_out_884 : u1_col_out_884;
assign col_out_885 = (sel_data_in)? u0_col_out_885 : u1_col_out_885;
assign col_out_886 = (sel_data_in)? u0_col_out_886 : u1_col_out_886;
assign col_out_887 = (sel_data_in)? u0_col_out_887 : u1_col_out_887;
assign col_out_888 = (sel_data_in)? u0_col_out_888 : u1_col_out_888;
assign col_out_889 = (sel_data_in)? u0_col_out_889 : u1_col_out_889;
assign col_out_890 = (sel_data_in)? u0_col_out_890 : u1_col_out_890;
assign col_out_891 = (sel_data_in)? u0_col_out_891 : u1_col_out_891;
assign col_out_892 = (sel_data_in)? u0_col_out_892 : u1_col_out_892;
assign col_out_893 = (sel_data_in)? u0_col_out_893 : u1_col_out_893;
assign col_out_894 = (sel_data_in)? u0_col_out_894 : u1_col_out_894;
assign col_out_895 = (sel_data_in)? u0_col_out_895 : u1_col_out_895;
assign col_out_896 = (sel_data_in)? u0_col_out_896 : u1_col_out_896;
assign col_out_897 = (sel_data_in)? u0_col_out_897 : u1_col_out_897;
assign col_out_898 = (sel_data_in)? u0_col_out_898 : u1_col_out_898;
assign col_out_899 = (sel_data_in)? u0_col_out_899 : u1_col_out_899;
assign col_out_900 = (sel_data_in)? u0_col_out_900 : u1_col_out_900;
assign col_out_901 = (sel_data_in)? u0_col_out_901 : u1_col_out_901;
assign col_out_902 = (sel_data_in)? u0_col_out_902 : u1_col_out_902;
assign col_out_903 = (sel_data_in)? u0_col_out_903 : u1_col_out_903;
assign col_out_904 = (sel_data_in)? u0_col_out_904 : u1_col_out_904;
assign col_out_905 = (sel_data_in)? u0_col_out_905 : u1_col_out_905;
assign col_out_906 = (sel_data_in)? u0_col_out_906 : u1_col_out_906;
assign col_out_907 = (sel_data_in)? u0_col_out_907 : u1_col_out_907;
assign col_out_908 = (sel_data_in)? u0_col_out_908 : u1_col_out_908;
assign col_out_909 = (sel_data_in)? u0_col_out_909 : u1_col_out_909;
assign col_out_910 = (sel_data_in)? u0_col_out_910 : u1_col_out_910;
assign col_out_911 = (sel_data_in)? u0_col_out_911 : u1_col_out_911;
assign col_out_912 = (sel_data_in)? u0_col_out_912 : u1_col_out_912;
assign col_out_913 = (sel_data_in)? u0_col_out_913 : u1_col_out_913;
assign col_out_914 = (sel_data_in)? u0_col_out_914 : u1_col_out_914;
assign col_out_915 = (sel_data_in)? u0_col_out_915 : u1_col_out_915;
assign col_out_916 = (sel_data_in)? u0_col_out_916 : u1_col_out_916;
assign col_out_917 = (sel_data_in)? u0_col_out_917 : u1_col_out_917;
assign col_out_918 = (sel_data_in)? u0_col_out_918 : u1_col_out_918;
assign col_out_919 = (sel_data_in)? u0_col_out_919 : u1_col_out_919;
assign col_out_920 = (sel_data_in)? u0_col_out_920 : u1_col_out_920;
assign col_out_921 = (sel_data_in)? u0_col_out_921 : u1_col_out_921;
assign col_out_922 = (sel_data_in)? u0_col_out_922 : u1_col_out_922;
assign col_out_923 = (sel_data_in)? u0_col_out_923 : u1_col_out_923;
assign col_out_924 = (sel_data_in)? u0_col_out_924 : u1_col_out_924;
assign col_out_925 = (sel_data_in)? u0_col_out_925 : u1_col_out_925;
assign col_out_926 = (sel_data_in)? u0_col_out_926 : u1_col_out_926;
assign col_out_927 = (sel_data_in)? u0_col_out_927 : u1_col_out_927;
assign col_out_928 = (sel_data_in)? u0_col_out_928 : u1_col_out_928;
assign col_out_929 = (sel_data_in)? u0_col_out_929 : u1_col_out_929;
assign col_out_930 = (sel_data_in)? u0_col_out_930 : u1_col_out_930;
assign col_out_931 = (sel_data_in)? u0_col_out_931 : u1_col_out_931;
assign col_out_932 = (sel_data_in)? u0_col_out_932 : u1_col_out_932;
assign col_out_933 = (sel_data_in)? u0_col_out_933 : u1_col_out_933;
assign col_out_934 = (sel_data_in)? u0_col_out_934 : u1_col_out_934;
assign col_out_935 = (sel_data_in)? u0_col_out_935 : u1_col_out_935;
assign col_out_936 = (sel_data_in)? u0_col_out_936 : u1_col_out_936;
assign col_out_937 = (sel_data_in)? u0_col_out_937 : u1_col_out_937;
assign col_out_938 = (sel_data_in)? u0_col_out_938 : u1_col_out_938;
assign col_out_939 = (sel_data_in)? u0_col_out_939 : u1_col_out_939;
assign col_out_940 = (sel_data_in)? u0_col_out_940 : u1_col_out_940;
assign col_out_941 = (sel_data_in)? u0_col_out_941 : u1_col_out_941;
assign col_out_942 = (sel_data_in)? u0_col_out_942 : u1_col_out_942;
assign col_out_943 = (sel_data_in)? u0_col_out_943 : u1_col_out_943;
assign col_out_944 = (sel_data_in)? u0_col_out_944 : u1_col_out_944;
assign col_out_945 = (sel_data_in)? u0_col_out_945 : u1_col_out_945;
assign col_out_946 = (sel_data_in)? u0_col_out_946 : u1_col_out_946;
assign col_out_947 = (sel_data_in)? u0_col_out_947 : u1_col_out_947;
assign col_out_948 = (sel_data_in)? u0_col_out_948 : u1_col_out_948;
assign col_out_949 = (sel_data_in)? u0_col_out_949 : u1_col_out_949;
assign col_out_950 = (sel_data_in)? u0_col_out_950 : u1_col_out_950;
assign col_out_951 = (sel_data_in)? u0_col_out_951 : u1_col_out_951;
assign col_out_952 = (sel_data_in)? u0_col_out_952 : u1_col_out_952;
assign col_out_953 = (sel_data_in)? u0_col_out_953 : u1_col_out_953;
assign col_out_954 = (sel_data_in)? u0_col_out_954 : u1_col_out_954;
assign col_out_955 = (sel_data_in)? u0_col_out_955 : u1_col_out_955;
assign col_out_956 = (sel_data_in)? u0_col_out_956 : u1_col_out_956;
assign col_out_957 = (sel_data_in)? u0_col_out_957 : u1_col_out_957;
assign col_out_958 = (sel_data_in)? u0_col_out_958 : u1_col_out_958;
assign col_out_959 = (sel_data_in)? u0_col_out_959 : u1_col_out_959;
assign col_out_960 = (sel_data_in)? u0_col_out_960 : u1_col_out_960;
assign col_out_961 = (sel_data_in)? u0_col_out_961 : u1_col_out_961;
assign col_out_962 = (sel_data_in)? u0_col_out_962 : u1_col_out_962;
assign col_out_963 = (sel_data_in)? u0_col_out_963 : u1_col_out_963;
assign col_out_964 = (sel_data_in)? u0_col_out_964 : u1_col_out_964;
assign col_out_965 = (sel_data_in)? u0_col_out_965 : u1_col_out_965;
assign col_out_966 = (sel_data_in)? u0_col_out_966 : u1_col_out_966;
assign col_out_967 = (sel_data_in)? u0_col_out_967 : u1_col_out_967;
assign col_out_968 = (sel_data_in)? u0_col_out_968 : u1_col_out_968;
assign col_out_969 = (sel_data_in)? u0_col_out_969 : u1_col_out_969;
assign col_out_970 = (sel_data_in)? u0_col_out_970 : u1_col_out_970;
assign col_out_971 = (sel_data_in)? u0_col_out_971 : u1_col_out_971;
assign col_out_972 = (sel_data_in)? u0_col_out_972 : u1_col_out_972;
assign col_out_973 = (sel_data_in)? u0_col_out_973 : u1_col_out_973;
assign col_out_974 = (sel_data_in)? u0_col_out_974 : u1_col_out_974;
assign col_out_975 = (sel_data_in)? u0_col_out_975 : u1_col_out_975;
assign col_out_976 = (sel_data_in)? u0_col_out_976 : u1_col_out_976;
assign col_out_977 = (sel_data_in)? u0_col_out_977 : u1_col_out_977;
assign col_out_978 = (sel_data_in)? u0_col_out_978 : u1_col_out_978;
assign col_out_979 = (sel_data_in)? u0_col_out_979 : u1_col_out_979;
assign col_out_980 = (sel_data_in)? u0_col_out_980 : u1_col_out_980;
assign col_out_981 = (sel_data_in)? u0_col_out_981 : u1_col_out_981;
assign col_out_982 = (sel_data_in)? u0_col_out_982 : u1_col_out_982;
assign col_out_983 = (sel_data_in)? u0_col_out_983 : u1_col_out_983;
assign col_out_984 = (sel_data_in)? u0_col_out_984 : u1_col_out_984;
assign col_out_985 = (sel_data_in)? u0_col_out_985 : u1_col_out_985;
assign col_out_986 = (sel_data_in)? u0_col_out_986 : u1_col_out_986;
assign col_out_987 = (sel_data_in)? u0_col_out_987 : u1_col_out_987;
assign col_out_988 = (sel_data_in)? u0_col_out_988 : u1_col_out_988;
assign col_out_989 = (sel_data_in)? u0_col_out_989 : u1_col_out_989;
assign col_out_990 = (sel_data_in)? u0_col_out_990 : u1_col_out_990;
assign col_out_991 = (sel_data_in)? u0_col_out_991 : u1_col_out_991;
assign col_out_992 = (sel_data_in)? u0_col_out_992 : u1_col_out_992;
assign col_out_993 = (sel_data_in)? u0_col_out_993 : u1_col_out_993;
assign col_out_994 = (sel_data_in)? u0_col_out_994 : u1_col_out_994;
assign col_out_995 = (sel_data_in)? u0_col_out_995 : u1_col_out_995;
assign col_out_996 = (sel_data_in)? u0_col_out_996 : u1_col_out_996;
assign col_out_997 = (sel_data_in)? u0_col_out_997 : u1_col_out_997;
assign col_out_998 = (sel_data_in)? u0_col_out_998 : u1_col_out_998;
assign col_out_999 = (sel_data_in)? u0_col_out_999 : u1_col_out_999;
assign col_out_1000 = (sel_data_in)? u0_col_out_1000 : u1_col_out_1000;
assign col_out_1001 = (sel_data_in)? u0_col_out_1001 : u1_col_out_1001;
assign col_out_1002 = (sel_data_in)? u0_col_out_1002 : u1_col_out_1002;
assign col_out_1003 = (sel_data_in)? u0_col_out_1003 : u1_col_out_1003;
assign col_out_1004 = (sel_data_in)? u0_col_out_1004 : u1_col_out_1004;
assign col_out_1005 = (sel_data_in)? u0_col_out_1005 : u1_col_out_1005;
assign col_out_1006 = (sel_data_in)? u0_col_out_1006 : u1_col_out_1006;
assign col_out_1007 = (sel_data_in)? u0_col_out_1007 : u1_col_out_1007;
assign col_out_1008 = (sel_data_in)? u0_col_out_1008 : u1_col_out_1008;
assign col_out_1009 = (sel_data_in)? u0_col_out_1009 : u1_col_out_1009;
assign col_out_1010 = (sel_data_in)? u0_col_out_1010 : u1_col_out_1010;
assign col_out_1011 = (sel_data_in)? u0_col_out_1011 : u1_col_out_1011;
assign col_out_1012 = (sel_data_in)? u0_col_out_1012 : u1_col_out_1012;
assign col_out_1013 = (sel_data_in)? u0_col_out_1013 : u1_col_out_1013;
assign col_out_1014 = (sel_data_in)? u0_col_out_1014 : u1_col_out_1014;
assign col_out_1015 = (sel_data_in)? u0_col_out_1015 : u1_col_out_1015;
assign col_out_1016 = (sel_data_in)? u0_col_out_1016 : u1_col_out_1016;
assign col_out_1017 = (sel_data_in)? u0_col_out_1017 : u1_col_out_1017;
assign col_out_1018 = (sel_data_in)? u0_col_out_1018 : u1_col_out_1018;
assign col_out_1019 = (sel_data_in)? u0_col_out_1019 : u1_col_out_1019;
assign col_out_1020 = (sel_data_in)? u0_col_out_1020 : u1_col_out_1020;
assign col_out_1021 = (sel_data_in)? u0_col_out_1021 : u1_col_out_1021;
assign col_out_1022 = (sel_data_in)? u0_col_out_1022 : u1_col_out_1022;
assign col_out_1023 = (sel_data_in)? u0_col_out_1023 : u1_col_out_1023;










endmodule
module xpb_5_825
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h9f8d426013718949489b07217d9f0e18a2bc0cdc8d90db967f8fc75ed7229440ef9f3872de4ab455077bc4970f48735b8393895d9c7bc74ab27ae43e399ba8b44da310d31e92c0721f45aab5addcac1e57bb0e6ef83af0de6b27000e4e8a29e5929ff0a854fdd7aa65572324dfa07c19fb7314d1baf51a8f5a87f07966eca351;
    5'b00010 : xpb = 1024'h8e6d3f6a64f4ddc9c630966beae3d4dfd402168845aa16b58142d567fb427b79dbf5f36cf26eea1b6f9949e73b32d5eca30cead51644be49b456891e3864dcb726f6ecf78d94839f2bf152c8c2dd940bbb71234563efb4ac20c16e21e2e9b138f6384f26f932b6c743ee5f6ac770d20aa80c4ac1259ed7ee6ea065ee44f6e037;
    5'b00011 : xpb = 1024'h7d4d3c74b678324a43c625b658289ba705482033fdc351d482f5e3711f6262b2c84cae6706931fe1d7b6cf37671d387dc2864c4c900db548b6322dfe372e10ba004ac91bfc9646cc389cfadbd7de7bf91f27381bcfa47879d65bdc357749388c59d0ada59d6795e422859bb0af4127fb54a580b09048954d82b8db6323011d1d;
    5'b00100 : xpb = 1024'h6c2d397f07fb86cac15bb500c56d626e368e29dfb5dc8cf384a8f17a438249ebb4a369611ab755a83fd4548793079b0ee1ffadc409d6ac47b80dd2de35f744bcd99ea5406b9809f94548a2eeecdf63e682dd4cf23b593c478bf64a490ba8bfdfbd690c24419c7501011cd7f697117dec013eb69ffaf252ac96d150d8010b5a03;
    5'b00101 : xpb = 1024'h5b0d3689597edb4b3ef1444b32b2293567d4338b6df5c812865bff8367a23124a0fa245b2edb8b6ea7f1d9d7bef1fda001790f3b839fa346b9e977be34c078bfb2f28164da99cd2651f44b0201e04bd3e69361c8a70e00154190b85ca008473321016aa2e5d1541ddfb4143c7ee1d3dcadd7ec8f659c100baae9c64cdf1596e9;
    5'b00110 : xpb = 1024'h49ed3393ab022fcbbc86d3959ff6effc991a3d37260f0331880f0d8c8bc2185d8d50df5542ffc135100f5f27eadc603120f270b2fd689a45bbc51c9e3389acc28c465d89499b90535e9ff31516e133c14a49769f12c2c3e2f72b26703467ce868499c9218a06333abe4b508266b229cd5a71227ed045cd6abf023bc1bd1fd3cf;
    5'b00111 : xpb = 1024'h38cd309dfc85844c3a1c62e00d3bb6c3ca6046e2de283e5089c21b95afe1ff9679a79a4f5723f6fb782ce47816c6c2c2406bd22a77319144bda0c17e3252e0c5659a39adb89d53806b4b9b282be21baeadff8b757e7787b0acc59483c8c755d9e83227a02e3b12579ce28cc84e827fbe070a586e3aef8ac9d31ab1369b2a10b5;
    5'b01000 : xpb = 1024'h27ad2da84e08d8ccb7b1f22a7a807d8afba6508e9641796f8b75299ed401e6cf65fe55496b482cc1e04a69c842b125535fe533a1f0fa8843bf7c665e311c14c83eee15d2279f16ad77f7433b40e3039c11b5a04bea2c4b7e626002975d26dd2d4bca861ed26ff1747b79c90e3652d5aeb3a38e5da5994828e73326ab79344d9b;
    5'b01001 : xpb = 1024'h168d2ab29f8c2d4d35478174e7c544522cec5a3a4e5ab48e8d2837a7f821ce08525510437f6c62884867ef186e9b87e47f5e95196ac37f42c1580b3e2fe548cb1841f1f696a0d9da84a2eb4e55e3eb89756bb52255e10f4c17fa70aaf1866480af62e49d76a4d0915a1105541e232b9f603cc44d10430587fb4b9c20573e8a81;
    5'b01010 : xpb = 1024'h56d27bcf10f81cdb2dd10bf550a0b195e3263e60673efad8edb45b11c41b5413eabcb3d9390984eb08574689a85ea759ed7f690e48c7641c333b01e2eae7ccdf195ce1b05a29d07914e93616ae4d376d921c9f8c195d319cd94debe85e5ebd412fb431c1ad9afae38a8419a05f381900cd5fa3c7aecc2e70f6411953548c767;
    5'b01011 : xpb = 1024'ha4fa6a1d04810b16fb7817e0d2a9193200ee70c29404cb440e6b0d0ff36449822e4b03b071db4ca3b80138ffa9ce5dd1226b7fee81083d8c75ae945c684a25823f38deee24355d79b0943e1718c17f9530dcd867b9d0c3f838bbdeccd47015b9a59b33c46fd787589dff64bee593fdaa08490f0e35e1dd7669ec020e9c356ab8;
    5'b01100 : xpb = 1024'h93da672756045f97790da72b3feddff932347a6e4c1e0663101e1b19178430bb1aa1beaa85ff826a201ebe4fd5b8c06241e4e165fad1348b778a393c67135985188cbb12933720a6bd3fe62a2dc267829492ed3e258587c5ee564ce068cf9d0d09339243140c66757c96a104cd64539ab4e244fda08b9ad57e0477837a3fa79e;
    5'b01101 : xpb = 1024'h82ba6431a787b417f6a33675ad32a6c0637a841a0437418211d129223ba417f406f879a49a23b830883c43a001a322f3615e42dd749a2b8a7965de1c65dc8d87f1e097370238e3d3c9eb8e3d42c34f6ff8490214913a4b93a3f0baf3fd2f24606ccbf0c1b84145925b2ddd4ab534a98b617b7aed0b355834921cecf85849e484;
    5'b01110 : xpb = 1024'h719a613bf90b08987438c5c01a776d8794c08dc5bc507ca11384372b5fc3ff2cf34f349eae47edf6f059c8f02d8d858480d7a454ee6322897b4182fc64a5c18acb34735b713aa700d697365057c4375d5bff16eafcef0f61598b2907918eabb3d0644f405c7624af39c519909d04ff7c0e14b0dc75df1593a635626d3654216a;
    5'b01111 : xpb = 1024'h607a5e464a8e5d18f1ce550a87bc344ec60697717469b7c01537453483e3e665dfa5ef98c26c23bd58774e405977e815a05105cc682c19887d1d27dc636ef58da4884f7fe03c6a2de342de636cc51f4abfb52bc168a3d32f0f25971b25ee330733fcadbf00ab03cc185c55d684d5556cbaade6cbe088d2f2ba4dd7e2145e5e50;
    5'b10000 : xpb = 1024'h4f5a5b509c11b1996f63e454f500fb15f74ca11d2c82f2df16ea533da803cd9ecbfcaa92d6905983c094d39085624aa6bfca6743e1f510877ef8ccbc623829907ddc2ba44f3e2d5aefee867681c60738236b4097d45896fcc4c0052eba4dba5a97950c3da4dfe2e8f6f3921c6ca5ab5d67471cbb4b329051ce664d56f2689b36;
    5'b10001 : xpb = 1024'h3e3a585aed950619ecf9739f6245c1dd2892aac8e49c2dfe189d6146cc23b4d7b853658ceab48f4a28b258e0b14cad37df43c8bb5bbe078680d4719c61015d93573007c8be3ff087fc9a2e8996c6ef258721556e400d5aca7a5a73424ead41adfb2d6abc4914c205d58ace625476014e13e052aab5dc4db0e27ec2cbd072d81c;
    5'b10010 : xpb = 1024'h2d1a55653f185a9a6a8f02e9cf8a88a459d8b4749cb5691d1a506f4ff0439c10a4aa2086fed8c51090cfde30dd370fc8febd2a32d586fe8582b0167c5fca91963083e3ed2d41b3b50945d69cabc7d712ead76a44abc21e982ff4e155e30cc9015ec5c93aed49a122b4220aa83c46573ec079889a20860b0ff6973840ae7d1502;
    5'b10011 : xpb = 1024'h1bfa526f909baf1ae82492343ccf4f6b8b1ebe2054cea43c1c037d59146383499100db8112fcfad6f8ed63810921725a1e368baa4f4ff584848bbb5c5e93c59909d7c0119c4376e215f17eafc0c8bf004e8d7f1b1776e265e58f4f69776c5054c25e27b9917e803f92b946ee2416ad2f6d12be898b2fc86f0aafadb58c8751e8;
    5'b10100 : xpb = 1024'hada4f79e21f039b65ba217eaa141632bc64c7cc0ce7df5b1db68b6238836a827d57967b2721309d610ae8d1350bd4eb3dafed21c918ec838667603c5d5cf99be32b9c360b453a0f229d26c2d5c9a6edb24393f1832ba6339b29bd7d0bcbd7a825f6863835b35f5c715083340be7032019abf478f5d985ce1ec8232a6a918ece;
    5'b10101 : xpb = 1024'haa6791d9f5908ce4ae5528a027b3244b5f20d4a89a78baf19d4652c10fa5fec36cf6ceee056be4f26886ad6844544846c143767f6594b3ce38e2447a96f8a25030cead0929d7fa8141e2d17883a6530c09fea2607b6697120650bd8b5a56018db89676e08ab13706d6a7a658eb877f3a151f094ab0cea05d795013a3d17e321f;
    5'b10110 : xpb = 1024'h99478ee44713e1652beab7ea94f7eb129066de545291f6109ef960ca33c5e5fc594d89e819901ab8d0a432b8703eaad7e0bcd7f6df5daacd3abde95a95c1d6530a22892d98d9bdae4e8e798b98a73af96db4b736e71b5adfbbeb2b9eeeb588e11c2ed55f2ee61623b53ee29ed357d52ac1b83f3a1b785dbc8d688918af886f05;
    5'b10111 : xpb = 1024'h88278bee989735e5a9804735023cb1d9c1ace8000aab312fa0ac6ed357e5cd3545a444e22db4507f38c1b8089c290d690036396e5926a1cc3c998e3a948b0a55e376655207db80db5b3a219eada822e6d16acc0d52d01ead718599b2831510347fc733ddd31af54093d61ee4bb282b1b6e51752986221b1ba180fe8d8d92abeb;
    5'b11000 : xpb = 1024'h770788f8ea1a8a662715d67f6f8178a0f2f2f1abc2c46c4ea25f7cdc7c05b46e31faffdc41d88645a0df3d58c8136ffa1faf9ae5d2ef98cb3e75331a93543e58bcca417676dd440867e5c9b1c2a90ad43520e0e3be84e27b272007c617749787e35f925c774fd45d726d5b2aa2f8810c1aeaab18f0cbd87ab59974026b9ce8d1;
    5'b11001 : xpb = 1024'h65e786033b9ddee6a4ab65c9dcc63f682438fb577adda76da4128ae5a0259ba71e51bad655fcbc0c08fcc2a8f3fdd28b3f28fc5d4cb88fca4050d7fa921d725b961e1d9ae5df0735749171c4d7a9f2c198d6f5ba2a39a648dcba75d9abd41edb46f7f0db1b84b37a510497708ac8d6fcc783e1085b7595d9c9b1e97749a725b7;
    5'b11010 : xpb = 1024'h54c7830d8d2133672240f5144a0b062f557f050332f6e28ca5c598eec44582e00aa875d06a20f1d2711a47f91fe8351c5ea25dd4c68186c9422c7cda90e6a65e6f71f9bf54e0ca62813d19d7ecaadaaefc8d0a9095ee6a169254e3ed4033a62eaa904f59bfb992972f9bd3b672992ced741d16f7c61f5338ddca5eec27b1629d;
    5'b11011 : xpb = 1024'h43a78017dea487e79fd6845eb74fccf686c50eaeeb101daba778a6f7e8656a18f6ff30ca7e452798d937cd494bd297ad7e1bbf4c404a7dc8440821ba8fafda6148c5d5e3c3e28d8f8de8c1eb01abc29c60431f6701a32de447ef5200d4932d820e28add863ee71b40e330ffc5a6982de20b64ce730c91097f1e2d46105bb9f83;
    5'b11100 : xpb = 1024'h32877d223027dc681d6c13a9249493bdb80b185aa32958caa92bb5010c855151e355ebc492695d5f4155529977bcfa3e9d9520c3ba1374c745e3c69a8e790e642219b20832e450bc9a9469fe16acaa89c3f9343d6d57f1b1fd89c01468f2b4d571c10c57082350d0ecca4c424239d8cecd4f82d69b72cdf705fb49d5e3c5dc69;
    5'b11101 : xpb = 1024'h21677a2c81ab30e89b01a2f391d95a84e95122065b4293e9aadec30a30a5388acfaca6bea68d9325a972d7e9a3a75ccfbd0e823b33dc6bc647bf6b7a8d424266fb6d8e2ca1e613e9a74012112bad927727af4913d90cb57fb3242e27fd523c28d5596ad5ac582fedcb6188882a0a2ebf79e8b8c6061c8b561a13bf4ac1d0194f;
    5'b11110 : xpb = 1024'h10477736d32e85691897323dff1e214c1a972bb2135bcf08ac91d11354c51fc3bc0361b8bab1c8ec11905d39cf91bf60dc87e3b2ada562c5499b105a8c0b7669d4c16a5110e7d716b3ebba2440ae7a648b655dea44c1794d68be9c3b91b1c37c38f1c954508d0f0aa9f8c4ce11da84b02681eeb570c648b52e2c34bf9fda5635;
    5'b11111 : xpb = 1024'hafd4b996e6a00eb26132395f7cbd2f64bd53388ea0ecaa9f2c2198722be7b404aba29a2b98fc7d41190c21d0deda32bc601b6d104a212a0ffc15f498c5a71f1e22647b242f7a9788d33164d9ee8b2682e3206c593cfc6a2bd3e59c49e03bed61cb91b9fca58ae6b50f4fe7f2f17b00ca21f503872bbb634488b4253906c6f986;
    endcase
end

endmodule

module xpb_5_145
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h10ec13be8c5966e3c2213e0bb9ccf58346a581ae4dbf43a9590a482b027701f2341e874e6aca6b8f4be6da91cd3518a0df560ef20db2bf61702c28e974eb2d638746c22eb9f3995fbcbf222e92a987ed41e5ec88524abe87a3cdcf9f46ba0e609c3fdc9aa939948117fbd571fbcaf04dd90ba7cc4250f7f5cd40bbae885cff7;
    5'b00010 : xpb = 1024'h21d8277d18b2cdc784427c177399eb068d4b035c9b7e8752b214905604ee03e4683d0e9cd594d71e97cdb5239a6a3141beac1de41b657ec2e05851d2e9d65ac70e8d845d73e732bf797e445d25530fda83cbd910a4957d0f479b9f3e8d741cc1387fb935527329022ff7aae3f795e09bb2174f9884a1efeb9a81775d10b9fee;
    5'b00011 : xpb = 1024'h32c43b3ba50c34ab4663ba232d66e089d3f0850ae93dcafc0b1ed881076505d69c5b95eb405f42ade3b48fb5679f49e29e022cd629183e2450847abc5ec1882a95d4468c2ddacc1f363d668bb7fc97c7c5b1c598f6e03b96eb696eddd42e2b21d4bf95cffbacbd8347f38055f360d0e98b22f764c6f2e7e167c2330b9916fe5;
    5'b00100 : xpb = 1024'h43b04efa31659b8f0884f82ee733d60d1a9606b936fd0ea5642920ac09dc07c8d07a1d39ab29ae3d2f9b6a4734d462837d583bc836cafd85c0b0a3a5d3acb58e1d1b08bae7ce657ef2fc88ba4aa61fb50797b221492afa1e8f373e7d1ae8398270ff726aa4e652045fef55c7ef2bc137642e9f310943dfd73502eeba2173fdc;
    5'b00101 : xpb = 1024'h549c62b8bdbf0272caa6363aa100cb90613b886784bc524ebd3368d70c5309bb0498a48815f419cc7b8244d902097b245cae4aba447dbce730dccc8f4897e2f1a461cae9a1c1fedeafbbaae8dd4fa7a2497d9ea99b75b8a633050e1c61a247e30d3f4f054e1fe68577eb2b39eaf6b1853d3a46fd4b94d7cd0243aa68a9d0fd3;
    5'b00110 : xpb = 1024'h658876774a1869568cc774465acdc113a7e10a15d27b95f8163db1020eca0bad38b72bd680be855bc7691f6acf3e93c53c0459ac52307c48a108f578bd8310552ba88d185bb5983e6c7acd176ff92f8f8b638b31edc0772dd6d2ddbba85c5643a97f2b9ff7597b068fe700abe6c1a1d31645eec98de5cfc2cf846617322dfca;
    5'b00111 : xpb = 1024'h76748a35d671d03a4ee8b252149ab696ee868bc4203ad9a16f47f92d11410d9f6cd5b324eb88f0eb134ff9fc9c73ac661b5a689e5fe33baa11351e62326e3db8b2ef4f4715a9319e2939ef4602a2b77ccd4977ba400b35b57aa0ad5aef1664a445bf083aa0930f87a7e2d61de28c9220ef519695d036c7b89cc521c5ba8afc1;
    5'b01000 : xpb = 1024'h87609df462cb371e1109f05dce67ac1a352c0d726dfa1d4ac852415813b80f91a0f43a7356535c7a5f36d48e69a8c506fab077906d95fb0b8161474ba7596b1c3a361175cf9ccafde5f91174954c3f6a0f2f64429255f43d1e6e7cfa35d07304e1fee4d549cca408bfdeab8fde57826ec85d3e621287bfae6a05dd7442e7fb8;
    5'b01001 : xpb = 1024'h984cb1b2ef249e01d32b2e698834a19d7bd18f20bbb960f4215c8983162f1183d512c1c1c11dc809ab1daf2036dddda7da0686827b48ba6cf18d70351c44987fc17cd3a48990645da2b833a327f5c757511550cae4a0b2c4c23c4c997c8a81657e3ec16ff3063889d7da8101da2272bca168e62e54d8b7a437469922cb44faf;
    5'b01010 : xpb = 1024'ha938c5717b7e04e5954c6c7542019720c27710cf0978a49d7a66d1ae18a61376093149102be83398f70489b20412f648b95c957488fb79ce61b9991e912fc5e348c395d34383fdbd5f7755d1ba9f4f4492fb3d5336eb714c660a1c38c3448fc61a7e9e0a9c3fcd0aefd65673d5ed630a7a748dfa9729af9a048754d153a1fa6;
    5'b01011 : xpb = 1024'hba24d93007d76bc9576daa80fbce8ca4091c927d5737e846d37119d91b1d15683d4fd05e96b29f2842eb6443d1480ee998b2a46696ae392fd1e5c208061af346d00a5801fd77971d1c3678004d48d731d4e129db89362fd409d7ebd809fe9e26b6be7aa54579618c07d22be5d1b85358538035c6d97aa78fd1c8107fdbfef9d;
    5'b01100 : xpb = 1024'hcb10ecee9430d2ad198ee88cb59b82274fc2142ba4f72bf02c7b62041d94175a716e57ad017d0ab78ed23ed59e7d278a7808b358a460f8914211eaf17b0620aa57511a30b76b307cd8f59a2edff25f1f16c71663db80ee5bada5bb7750b8ac8752fe573feeb2f60d1fce0157cd8343a62c8bdd931bcb9f859f08cc2e645bf94;
    5'b01101 : xpb = 1024'hdbfd00ad208a3990dbb026986f6877aa966795d9f2b66f998585aa2f200b194ca58cdefb6c477646dab919676bb2402b575ec24ab213b7f2b23e13daeff14e0dde97dc5f715ec9dc95b4bc5d729be70c58ad02ec2dcbace351738b169772bae7ef3e33da97ec8a8e37c9d6c9c94e33f40597855f5e1c977b6c4987dcecb8f8b;
    5'b01110 : xpb = 1024'hece9146bace3a0749dd164a429356d2ddd0d17884075b342de8ff25a22821b3ed9ab6649d711e1d6269ff3f938e758cc36b4d13cbfc67754226a3cc464dc7b7165de9e8e2b52633c5273de8c05456ef99a92ef7480166b6af5415ab5de2cc9488b7e107541261f0f4fc5ac3bc5192441dea32d2ba06d8f71398a438b7515f82;
    5'b01111 : xpb = 1024'hfdd5282a393d07585ff2a2afe30262b123b299368e34f6ec379a3a8524f91d310dc9ed9841dc4d657286ce8b061c716d160ae02ecd7936b5929665add9c7a8d4ed2560bce545fc9c0f3300ba97eef6e6dc78dbfcd26129f2990f2a5524e6d7a927bded0fea5fb39067c181adc0e4148fb7aed4f7e2be876706caff39fd72f79;
    5'b10000 : xpb = 1024'h10ec13be8c5966e3c2213e0bb9ccf58346a581ae4dbf43a9590a482b027701f2341e874e6aca6b8f4be6da91cd3518a0df560ef20db2bf61702c28e974eb2d638746c22eb9f3995fbcbf222e92a987ed41e5ec88524abe87a3cdcf9f46ba0e609c3fdc9aa939948117fbd571fbcaf04dd90ba7cc4250f7f5cd40bbae885cff70;
    5'b10001 : xpb = 1024'h11fad4fa751efd51fe4351ec7569c4db7b0fd9c9329b37e3ee9aecadb29e721157606fc35177124840a5483aea086a2aed4b6fe12e8deb57872eeb780c39e039bfbb2e51a592d2f5b88b14517bd4206c16044b50d76f6a701e0aac993b25af46a603da6453cd2dc9297b92c91b879f52b69c6249067607752a14c76970e2cf67;
    5'b10010 : xpb = 1024'h130996365de493c03a6565cd31069433af7a31e417772c1e842b913062c5e2307aa258383823b9013563b5e406dbbbb4fb40d0d04f69174d9e31ae06a388930ff82f9a7491320c8bb457067464feb8eaea22aa195c941658984789932f91502cafc7d82dfe60c7113afb50203b444e57942d1cc5ca9b16f486e8d32459689f5e;
    5'b10011 : xpb = 1024'h1418577246aa2a2e768779adeca3638be3e489fefc53205919bc35b312ed524f9de440ad1ed05fba2a22238d23af0d3f093631bf70444343b53470953ad745e630a406977cd14621b022f8974e295169be4108e1e1b8c2411284668d23fcf112b98bd5f7a8f460594c7b0d775b00fd5c71bdd7428ec02673e3bcdedf41ee6f55;
    5'b10100 : xpb = 1024'h152718ae2f6fc09cb2a98d8ea84032e4184ee219e12f1493af4cda35c314c26ec1262922057d06731ee0913640825ec9172b92ae911f6f39cc373323d225f8bc691872ba68707fb7abeeeaba3753e9e8925f67aa66dd6e298cc14387186891f8c34fd3c15387f9a15dfacace7abdac614f4e91bf52e535f34090ea9a2a743f4c;
    5'b10101 : xpb = 1024'h1635d9ea1835570aeecba16f63dd023c4cb93a34c60b08ce44dd7eb8733c328de4681196ec29ad2c139efedf5d55b0532520f39db1fa9b2fe339f5b26974ab92a18cdedd540fb94da7badcdd207e8267667dc672ec021a1206fe20810cd432decd13d18afe1b92e96f7a88259a7a5b662cdf4c3c170a45729d64f65512fa0f43;
    5'b10110 : xpb = 1024'h17449b2600faed792aedb5501f79d1948123924faae6fd08da6e233b2363a2ad07a9fa0bd2d653e5085d6c887a2901dd3316548cd2d5c725fa3cb84100c35e68da014b003faef2e3a386cf0009a91ae63a9c253b7126c5fa813afd7b013fd3c4d6d7cf54a8af2c3180fa457cba370a6b0a7006b8db2f54f1fa39020ffb7fdf3a;
    5'b10111 : xpb = 1024'h18535c61e9c083e7670fc930db16a0ecb58dea6a8fc2f1436ffec7bdd38b12cc2aebe280b982fa9dfd1bda3196fc5367410bb57bf3b0f31c113f7acf9812113f1275b7232b4e2c799f52c122f2d3b3650eba8403f64b71e2fb77da74f5ab74aae09bcd1e5342c579927a02d3d9f3b96fe800c1359f546471570d0dcae405af31;
    5'b11000 : xpb = 1024'h19621d9dd2861a55a331dd1196b37044e9f84285749ee57e058f6c4083b282eb4e2dcaf5a02fa156f1da47dab3cfa4f14f01166b148c1f1228423d5e2f60c4154aea234616ed660f9b1eb345dbfe4be3e2d8e2cc7b701dcb75b4b76eea171590ea5fcae7fdd65ec1a3f9c02af9b06874c5917bb2637973f0b3e11985cc8b7f28;
    5'b11001 : xpb = 1024'h1a70ded9bb4bb0c3df53f0f252503f9d1e629aa0597ad9b89b2010c333d9f30a716fb36a86dc480fe698b583d0a2f67b5cf6775a35674b083f44ffecc6af76eb835e8f69028c9fa596eaa568c528e462b6f741950094c9b3eff19468de82b676f423c8b1a869f809b5797d82196d1779a322362f279e837010b52540b5114f1f;
    5'b11010 : xpb = 1024'h1b7fa015a41147321b7604d30ded0ef552ccf2bb3e56cdf330b0b545e401632994b19bdf6d88eec8db57232ced7648056aebd849564276fe5647c27b5dfe29c1bbd2fb8bee2bd93b92b6978bae537ce18b15a05d85b9759c6a2e7162d2ee575cfde7c67b52fd9151c6f93ad93929c67e80b2f0abebc392ef6d8930fb9d971f16;
    5'b11011 : xpb = 1024'h1c8e61518cd6dda0579818b3c989de4d87374ad62332c22dc64159c89428d348b7f3845454359581d01590d60a49998f78e13938771da2f46d4a8509f54cdc97f44767aed9cb12d18e8289ae977e15605f33ff260ade2184e46b4e5cc759f84307abc444fd912a99d878f83058e675835e43ab28afe8a26eca5d3cb6861cef0d;
    5'b11100 : xpb = 1024'h1d9d228d759c740e93ba2c948526ada5bba1a2f1080eb6685bd1fe4b44504367db356cc93ae23c3ac4d3fe7f271ceb1986d69a2797f8ceea844d47988c9b8f6e2cbbd3d1c56a4c678a4e7bd180a8addf33525dee9002cd6d5ea82b56bbc59929116fc20ea824c3e1e9f8b58778a324883bd465a5740db1ee273148716ea2bf04;
    5'b11101 : xpb = 1024'h1eabe3c95e620a7ccfdc407540c37cfdf00bfb0beceaaaa2f162a2cdf477b386fe77553e218ee2f3b9926c2843f03ca394cbfb16b8d3fae09b500a2723ea424465303ff4b10985fd861a6df469d3465e0770bcb715277955d8e50850b0313a0f1b33bfd852b85d29fb7872de985fd38d196520223832c16d8405542c57288efb;
    5'b11110 : xpb = 1024'h1fbaa5054727a0eb0bfe5455fc604c5624765326d1c69edd86f34750a49f23a621b93db3083b89acae50d9d160c38e2da2c15c05d9af26d6b252ccb5bb38f51a9da4ac179ca8bf9381e6601752fddedcdb8f1b7f9a4c253e5321e54aa49cdaf524f7bda1fd4bf6720cf83035b81c8291f6f5da9efc57d0ece0d95fe73fae5ef2;
    5'b11111 : xpb = 1024'h20c966412fed375948206836b7fd1bae58e0ab41b6a293181c83ebd354c693c544fb2627eee83065a30f477a7d96dfb7b0b6bcf4fa8a52ccc9558f445287a7f0d619183a8847f9297db2523a3c28775bafad7a481f70d126cd5ec24499087bdb2ebbbb6ba7df8fba1e77ed8cd7d93196d486951bc07ce06c3dad6ba228342ee9;
    endcase
end

endmodule

module xpb_5_45
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h531b4da555074852e49aae7ac4081938c236f783b60ee12bcd6ab660d2d6b10381ec6a88e97ab0b6a9821be7ffa401c3ddfa3f0308ff9a7c5aaf416407cad6bd286bcc9a9f9e83ad78c3cbdc7381696bf58553491b62df315aaf39095e0cdd6631aa7702efb0ac3623884cdae47d13a44e2e5372c49b5122934964a977b6ea7d;
    5'b00010 : xpb = 1024'ha6369b4aaa0e90a5c9355cf588103271846def076c1dc2579ad56cc1a5ad620703d8d511d2f5616d530437cfff480387bbf47e0611ff34f8b55e82c80f95ad7a50d799353f3d075af18797b8e702d2d7eb0aa69236c5be62b55e7212bc19bacc6354ee05df61586c471099b5c8fa27489c5ca6e58936a2452692c952ef6dd4fa;
    5'b00011 : xpb = 1024'h48a4a39a3d27a42fe2ca93993bbe0458d52ee35a4cb5030bea6369ccc5816602827cc221f24993955d2814711b8df48135d49522f84bff295f6e84cddc8e0f8604f431212f4a8dc357b160f2c1a87812ec8b0042c5a270835a8119215ffbf5a065f7d2df1e490c14e3d8ffb1b5a714c39bb11b75fd869637736cb2f7de42590c;
    5'b00100 : xpb = 1024'h9bbff13f922eec82c7654213ffc61d919765dade02c3e437b7ce202d9858170604692caadbc4444c06aa30591b31f64513ced426014b99a5ba1dc631e458e6432d5ffdbbcee91170d0752ccf3529e17ee210538be1054fb4b530522abe08d30697a249e20df9b84b07614c8c9a242867e9df6ee8c221e75a06b617a155f94389;
    5'b00101 : xpb = 1024'h3e2df98f2548000ce0fa78b7b373ef78e826cf30e35b24ec075c1d38b82c1b01830d19bafb18767410ce0cfa3777e73e8daeeb42e79863d6642dc837b151484ee17c95a7bef697d9369ef6090fcf86b9e390ad3c6fe201d55a52f93961eb0dda9a452ebb4ce16bf3a429b28886d115e2e933e3793671db4c5390014644cdc79b;
    5'b00110 : xpb = 1024'h914947347a4f485fc5952732777c08b1aa5dc6b4996a0617d4c6d3998b02cc0504f98443e493272aba5028e2371be9026ba92a45f097fe52bedd099bb91c1f0c09e862425e951b86af62c1e58350f025d91600858b44e106b5023242bff7eb40cbefa5be3c921829c7b1ff636b4e2987376236ebfb0d2c6ee6d965efbc84b218;
    5'b00111 : xpb = 1024'h33b74f840d685be9df2a5dd62b29da98fb1ebb077a0146cc2454d0a4aad6d000839d715403e75952c47405835361d9fbe5894162d6e4c88368ed0ba186148117be04fa2e4ea2a1ef158c8b1f5df69560da965a361a2193275a24d95163da2614ce928a977b79cbd2647a655f57fb170236b6ab7c6f5d206133b34f94ab59362a;
    5'b01000 : xpb = 1024'h86d29d29626fa43cc3c50c50ef31f3d1bd55b28b301027f7f1bf87057dad81040589dbdced620a096df6216b5305dbbfc3838065dfe462ffc39c4d058ddf57d4e670c6c8ee41259c8e5056fbd177feccd01bad7f35847258b4d4125ac1e7037b003d019a6b2a78088802b23a3c782aa684e4feef33f87183c6fcb43e231020a7;
    5'b01001 : xpb = 1024'h2940a578f588b7c6dd5a42f4a2dfc5b90e16a6de10a768ac414d84109d8184ff842dc8ed0cb63c317819fe0c6f4bccb93d639782c6312d306dac4f0b5ad7b9e09a8d5eb4de4eac04f47a2035ac1da407d19c072fc461247959f6b96965c93e4f02dfe673aa122bb124cb1836292518218439737fa848657613d69de311e4a4b9;
    5'b01010 : xpb = 1024'h7c5bf31e4a900019c1f4f16f66e7def1d04d9e61c6b649d80eb83a7170583603061a3375f630ece8219c19f46eefce7d1b5dd685cf30c7acc85b906f62a2909dc2f92b4f7ded2fb26d3dec121f9f0d73c7215a78dfc403aab4a5f272c3d61bb5348a5d7699c2d7e7485365110da22bc5d267c6f26ce3b698a720028c899b8f36;
    5'b01011 : xpb = 1024'h1ec9fb6ddda913a3db8a28131a95b0d9210e92b4a74d8a8c5e46377c902c39fe84be208615851f102bbff6958b35bf76953deda2b57d91dd726b92752f9af2a97715c33b6dfab61ad367b54bfa44b2aec8a1b4296ea0b5cb59c8998167b85689372d424fd8aa8b8fe51bcb0cfa4f1940d1bc3b82e133aa8af3f9ec3178701348;
    5'b01100 : xpb = 1024'h71e5491332b05bf6c024d68dde9dca11e3458a385d5c6bb82bb0eddd6302eb0206aa8b0efeffcfc6d542127d8ad9c13a73382ca5be7d2c59cd1ad3d93765c9669f818fd60d9939c84c2b81286dc61c1abe2707728a0394fcb477d28ac5c533ef68d7b952c85b37c608a417e7decc2ce51fea8ef5a5cefbad874350daf026fdc5;
    5'b01101 : xpb = 1024'h14535162c5c96f80d9ba0d31924b9bf934067e8b3df3ac6c7b3eeae882d6eefd854e781f1e5401eedf65ef1ea71fb233ed1843c2a4c9f68a772ad5df045e2b72539e27c1fda6c030b2554a62486bc155bfa7612318e0471d599a799969a76ec36b7a9e2c0742eb6ea56c7de3cb791a601f3f03861a1eef9fd41d3a7fdefb81d7;
    5'b01110 : xpb = 1024'h676e9f081ad0b7d3be54bbac5653b531f63d760ef4028d9848a9a14955ada001073ae2a807ceb2a588e80b06a6c3b3f7cb1282c5adc99106d1da17430c29022f7c09f45c9d4543de2b19163ebbed2ac1b52cb46c3443264eb449b2a2c7b44c299d25152ef6f397a4c8f4cabeaff62e046d6d56f8deba40c267669f2956b26c54;
    5'b01111 : xpb = 1024'h9dca757ade9cb5dd7e9f2500a01871946fe6a61d499ce4c98379e547581a3fc85decfb82722e4cd930be7a7c309a4f144f299e294165b377bea1948d921643b30268c488d52ca469142df789692cffcb6ad0e1cc31fd86f596c59b16b9686fd9fc7fa0835db4b4d65bd30ba9ca31b7f6cc1cb89530a34b4b44088ce4586f066;
    5'b10000 : xpb = 1024'h5cf7f4fd02f113b0bc84a0cace09a052093561e58aa8af7865a254b54858550007cb3a41109d95843c8e038fc2ada6b522ecd8e59d15f5b3d6995aace0ec3af8589258e32cf14df40a06ab550a143968ac326165de82b7a0b41b92bac9a36463d172710b258bf78389457d9581202f23baf01efc17a585d74789ed77bd3ddae3;
    5'b10001 : xpb = 1024'hb01342a257f85c03a11f4f459211b98acb6c596940b790a4330d0b161b2f060389b7a4c9fa18463ae6101f77c251a87900e717e8a615903031489c10e8b711b580fe257dcc8fd1a182ca77317d95a2d4a1b7b4aef9e596d20ecacbc427b041ca031ce80e153ca3b9accdca70659d42c8091e726edc40d6f9dad3522134f4c560;
    5'b10010 : xpb = 1024'h52814af1eb116f8dbab485e945bf8b721c2d4dbc214ed158829b08213b0309ff085b91da196c7862f033fc18de9799727ac72f058c625a60db589e16b5af73c1351abd69bc9d5809e8f4406b583b480fa3380e5f88c248f2b3ed72d2cb927c9e05bfcce7542457624996306c524a30430872e6ff5090caec27ad3bc623c94972;
    5'b10011 : xpb = 1024'ha59c98974018b7e09f4f346409c7a4aade64453fd75db2845005be820dd9bb028a47fc6302e7291999b61800de3b9b3658c16e089561f4dd3607df7abd7a4a7e5d868a045c3bdbb761b80c47cbbcb17b98bd61a8a42528240e9cabdc299f5a04376a43ea43d503986d1e7d4736c743e756a13a72152c1c0ebaf6a06f9b8033ef;
    5'b10100 : xpb = 1024'h480aa0e6d331cb6ab8e46b07bd7576922f253992b7f4f3389f93bb8d2dadbefe08ebe973223b5b41a3d9f4a1fa818c2fd2a185257baebf0de017e1808a72ac8a11a321f04c49621fc7e1d581a66256b69a3dbb593301da44b3bf52eacd8194d83a0d28c382bcb74109e6e3432374316255f5af02897c100107d08a148a54b801;
    5'b10101 : xpb = 1024'h9b25ee8c283913bd9d7f1982817d8fcaf15c31166e03d4646cfe71ee008470018ad853fc0bb60bf84d5c1089fa258df3b09bc42884ae598a3ac722e4923d83473a0eee8aebe7e5cd40a5a15e19e3c0228fc30ea24e64b9760e6e8bf42b8e723e6bb79fc6726d63772d6f301e07f14506a42402754e1761239b19eebe020ba27e;
    5'b10110 : xpb = 1024'h3d93f6dbbb522747b7145026352b61b2421d25694e9b1518bc8c6ef9205873fd097c410c2b0a3e20577fed2b166b7eed2a7bdb456afb23bae4d724ea5f35e552ee2b8676dbf56c35a6cf6a97f489655d91436852dd416b96b3913302cf70ad126e5a849fb155171fca379619f49e3281a3787705c2675515e7f3d862f0e02690;
    5'b10111 : xpb = 1024'h90af448110596f9a9baefea0f9337aeb04541ced04a9f64489f72559f32f25008b68ab951484eed701020913160f80b108761a4873fabe373f86664e6700bc10169753117b93efe31f933674680acec986c8bb9bf8a44ac80e406c0c2d7d8a78a004fba2a105c355edbfe2f4d91b4625f1a6ca788702a6387b3d3d0c6897110d;
    5'b11000 : xpb = 1024'h331d4cd0a3728324b5443544ace14cd25515113fe54136f8d9852265130328fc0a0c98a533d920ff0b25e5b4325571aa825631655a478867e996685433f91e1bcab3eafd6ba1764b85bcffae42b074048849154c8780fce8b363131ad15fc54ca2a7e07bdfed76fe8a8848f0c5c833a0f0fb3f08fb529a2ac81726b1576b951f;
    5'b11001 : xpb = 1024'h86389a75f879cb7799dee3bf70e9660b174c08c39b501824a6efd8c5e5d9d9ff8bf9032e1d53d1b5b4a8019c31f9736e60507068634722e44445a9b83bc3f4d8f31fb7980b3ff9f8fe80cb8ab631dd707dce6895a2e3dc1a0e124c242f6ca2b2d452577ecf9e2334ae1095cbaa4547453f29927bbfedeb4d5b608b5acf227f9c;
    5'b11010 : xpb = 1024'h28a6a2c58b92df01b3741a63249737f2680cfd167be758d8f67dd5d105adddfb0a9cf03e3ca803ddbecbde3d4e3f6467da3087854993ed14ee55abbe08bc56e4a73c4f83fb4d806164aa94c490d782ab7f4ec24631c08e3ab334f332d34edd86d6f53c580e85d6dd4ad8fbc796f234c03e7e070c343ddf3fa83a74ffbdf703ae;
    5'b11011 : xpb = 1024'h7bc1f06ae09a2754980ec8dde89f512b2a43f49a31f63a04c3e88c31d8848efe8c895ac72622b494684dfa254de3662bb82ac688529387914904ed2210872da1cfa81c1e9aec040edd6e60a10458ec1774d4158f4d236d6c0de42c3c315bbaed089fb35afe3683136e6148a27b6f48648cac5a7ef8d930623b83d9a935adee2b;
    5'b11100 : xpb = 1024'h1e2ff8ba73b33adeb1a3ff819c4d23127b04e8ed128d7ab91376893cf85892fa0b2d47d74576e6bc7271d6c66a295725320adda538e051c1f314ef27dd7f8fad83c4b40a8af98a77439829dadefe915276546f3fdc001f8cb306d34ad53df5c10b4298343d1e36bc0b29ae9e681c35df8c00cf0f6d292454885dc34e2482723d;
    5'b11101 : xpb = 1024'h714b465fc8ba8331963eadfc60553c4b3d3be070c89c5be4e0e13f9dcb2f43fd8d19b2602ef197731bf3f2ae69cd58e910051ca841dfec3e4dc4308be54a666aac3080a52a980e24bc5bf5b7527ffabe6bd9c288f762febe0db60c54334ad3273ced0f372ccee2f22eb1fb794c994983da2f228231c475771ba727f79c395cba;
    5'b11110 : xpb = 1024'h13b94eaf5bd396bbafd3e4a014030e328dfcd4c3a9339c99306f3ca8eb0347f90bbd9f704e45c99b2617cf4f861349e289e533c5282cb66ef7d43291b242c876604d18911aa5948d2285bef12d259ff96d5a1c39863fb0deb2d8b362d72d0dfb3f8ff4106bb6969acb7a6175394636fed9839712a61469696881119c8b0de0cc;
    5'b11111 : xpb = 1024'h66d49c54b0dadf0e946e931ad80b276b5033cc475f427dc4fdd9f309bdd9f8fc8daa09f937c07a51cf99eb3785b74ba667df72c8312c50eb528373f5ba0d9f3388b8e52bba44183a9b498acda0a7096562df6f82a1a290100d87ec6c3539eb61713a6b135b6742d0ef02ae501dc34aa327b1ea856aafba8bfbca764602c4cb49;
    endcase
end

endmodule

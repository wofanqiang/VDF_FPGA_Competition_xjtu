module alu
(
    input  [511:0] col_in_0,
    input  [511:0] col_in_1,
    input  [511:0] col_in_2,
    input  [511:0] col_in_3,
    input  [511:0] col_in_4,
    input  [511:0] col_in_5,
    input  [511:0] col_in_6,
    input  [511:0] col_in_7,
    input  [511:0] col_in_8,
    input  [511:0] col_in_9,
    input  [511:0] col_in_10,
    input  [511:0] col_in_11,
    input  [511:0] col_in_12,
    input  [511:0] col_in_13,
    input  [511:0] col_in_14,
    input  [511:0] col_in_15,
    input  [511:0] col_in_16,
    input  [511:0] col_in_17,
    input  [511:0] col_in_18,
    input  [511:0] col_in_19,
    input  [511:0] col_in_20,
    input  [511:0] col_in_21,
    input  [511:0] col_in_22,
    input  [511:0] col_in_23,
    input  [511:0] col_in_24,
    input  [511:0] col_in_25,
    input  [511:0] col_in_26,
    input  [511:0] col_in_27,
    input  [511:0] col_in_28,
    input  [511:0] col_in_29,
    input  [511:0] col_in_30,
    input  [511:0] col_in_31,
    input  [511:0] col_in_32,
    input  [511:0] col_in_33,
    input  [511:0] col_in_34,
    input  [511:0] col_in_35,
    input  [511:0] col_in_36,
    input  [511:0] col_in_37,
    input  [511:0] col_in_38,
    input  [511:0] col_in_39,
    input  [511:0] col_in_40,
    input  [511:0] col_in_41,
    input  [511:0] col_in_42,
    input  [511:0] col_in_43,
    input  [511:0] col_in_44,
    input  [511:0] col_in_45,
    input  [511:0] col_in_46,
    input  [511:0] col_in_47,
    input  [511:0] col_in_48,
    input  [511:0] col_in_49,
    input  [511:0] col_in_50,
    input  [511:0] col_in_51,
    input  [511:0] col_in_52,
    input  [511:0] col_in_53,
    input  [511:0] col_in_54,
    input  [511:0] col_in_55,
    input  [511:0] col_in_56,
    input  [511:0] col_in_57,
    input  [511:0] col_in_58,
    input  [511:0] col_in_59,
    input  [511:0] col_in_60,
    input  [511:0] col_in_61,
    input  [511:0] col_in_62,
    input  [511:0] col_in_63,
    input  [511:0] col_in_64,
    input  [511:0] col_in_65,
    input  [511:0] col_in_66,
    input  [511:0] col_in_67,
    input  [511:0] col_in_68,
    input  [511:0] col_in_69,
    input  [511:0] col_in_70,
    input  [511:0] col_in_71,
    input  [511:0] col_in_72,
    input  [511:0] col_in_73,
    input  [511:0] col_in_74,
    input  [511:0] col_in_75,
    input  [511:0] col_in_76,
    input  [511:0] col_in_77,
    input  [511:0] col_in_78,
    input  [511:0] col_in_79,
    input  [511:0] col_in_80,
    input  [511:0] col_in_81,
    input  [511:0] col_in_82,
    input  [511:0] col_in_83,
    input  [511:0] col_in_84,
    input  [511:0] col_in_85,
    input  [511:0] col_in_86,
    input  [511:0] col_in_87,
    input  [511:0] col_in_88,
    input  [511:0] col_in_89,
    input  [511:0] col_in_90,
    input  [511:0] col_in_91,
    input  [511:0] col_in_92,
    input  [511:0] col_in_93,
    input  [511:0] col_in_94,
    input  [511:0] col_in_95,
    input  [511:0] col_in_96,
    input  [511:0] col_in_97,
    input  [511:0] col_in_98,
    input  [511:0] col_in_99,
    input  [511:0] col_in_100,
    input  [511:0] col_in_101,
    input  [511:0] col_in_102,
    input  [511:0] col_in_103,
    input  [511:0] col_in_104,
    input  [511:0] col_in_105,
    input  [511:0] col_in_106,
    input  [511:0] col_in_107,
    input  [511:0] col_in_108,
    input  [511:0] col_in_109,
    input  [511:0] col_in_110,
    input  [511:0] col_in_111,
    input  [511:0] col_in_112,
    input  [511:0] col_in_113,
    input  [511:0] col_in_114,
    input  [511:0] col_in_115,
    input  [511:0] col_in_116,
    input  [511:0] col_in_117,
    input  [511:0] col_in_118,
    input  [511:0] col_in_119,
    input  [511:0] col_in_120,
    input  [511:0] col_in_121,
    input  [511:0] col_in_122,
    input  [511:0] col_in_123,
    input  [511:0] col_in_124,
    input  [511:0] col_in_125,
    input  [511:0] col_in_126,
    input  [511:0] col_in_127,
    input  [511:0] col_in_128,
    input  [511:0] col_in_129,
    input  [511:0] col_in_130,
    input  [511:0] col_in_131,
    input  [511:0] col_in_132,
    input  [511:0] col_in_133,
    input  [511:0] col_in_134,
    input  [511:0] col_in_135,
    input  [511:0] col_in_136,
    input  [511:0] col_in_137,
    input  [511:0] col_in_138,
    input  [511:0] col_in_139,
    input  [511:0] col_in_140,
    input  [511:0] col_in_141,
    input  [511:0] col_in_142,
    input  [511:0] col_in_143,
    input  [511:0] col_in_144,
    input  [511:0] col_in_145,
    input  [511:0] col_in_146,
    input  [511:0] col_in_147,
    input  [511:0] col_in_148,
    input  [511:0] col_in_149,
    input  [511:0] col_in_150,
    input  [511:0] col_in_151,
    input  [511:0] col_in_152,
    input  [511:0] col_in_153,
    input  [511:0] col_in_154,
    input  [511:0] col_in_155,
    input  [511:0] col_in_156,
    input  [511:0] col_in_157,
    input  [511:0] col_in_158,
    input  [511:0] col_in_159,
    input  [511:0] col_in_160,
    input  [511:0] col_in_161,
    input  [511:0] col_in_162,
    input  [511:0] col_in_163,
    input  [511:0] col_in_164,
    input  [511:0] col_in_165,
    input  [511:0] col_in_166,
    input  [511:0] col_in_167,
    input  [511:0] col_in_168,
    input  [511:0] col_in_169,
    input  [511:0] col_in_170,
    input  [511:0] col_in_171,
    input  [511:0] col_in_172,
    input  [511:0] col_in_173,
    input  [511:0] col_in_174,
    input  [511:0] col_in_175,
    input  [511:0] col_in_176,
    input  [511:0] col_in_177,
    input  [511:0] col_in_178,
    input  [511:0] col_in_179,
    input  [511:0] col_in_180,
    input  [511:0] col_in_181,
    input  [511:0] col_in_182,
    input  [511:0] col_in_183,
    input  [511:0] col_in_184,
    input  [511:0] col_in_185,
    input  [511:0] col_in_186,
    input  [511:0] col_in_187,
    input  [511:0] col_in_188,
    input  [511:0] col_in_189,
    input  [511:0] col_in_190,
    input  [511:0] col_in_191,
    input  [511:0] col_in_192,
    input  [511:0] col_in_193,
    input  [511:0] col_in_194,
    input  [511:0] col_in_195,
    input  [511:0] col_in_196,
    input  [511:0] col_in_197,
    input  [511:0] col_in_198,
    input  [511:0] col_in_199,
    input  [511:0] col_in_200,
    input  [511:0] col_in_201,
    input  [511:0] col_in_202,
    input  [511:0] col_in_203,
    input  [511:0] col_in_204,
    input  [511:0] col_in_205,
    input  [511:0] col_in_206,
    input  [511:0] col_in_207,
    input  [511:0] col_in_208,
    input  [511:0] col_in_209,
    input  [511:0] col_in_210,
    input  [511:0] col_in_211,
    input  [511:0] col_in_212,
    input  [511:0] col_in_213,
    input  [511:0] col_in_214,
    input  [511:0] col_in_215,
    input  [511:0] col_in_216,
    input  [511:0] col_in_217,
    input  [511:0] col_in_218,
    input  [511:0] col_in_219,
    input  [511:0] col_in_220,
    input  [511:0] col_in_221,
    input  [511:0] col_in_222,
    input  [511:0] col_in_223,
    input  [511:0] col_in_224,
    input  [511:0] col_in_225,
    input  [511:0] col_in_226,
    input  [511:0] col_in_227,
    input  [511:0] col_in_228,
    input  [511:0] col_in_229,
    input  [511:0] col_in_230,
    input  [511:0] col_in_231,
    input  [511:0] col_in_232,
    input  [511:0] col_in_233,
    input  [511:0] col_in_234,
    input  [511:0] col_in_235,
    input  [511:0] col_in_236,
    input  [511:0] col_in_237,
    input  [511:0] col_in_238,
    input  [511:0] col_in_239,
    input  [511:0] col_in_240,
    input  [511:0] col_in_241,
    input  [511:0] col_in_242,
    input  [511:0] col_in_243,
    input  [511:0] col_in_244,
    input  [511:0] col_in_245,
    input  [511:0] col_in_246,
    input  [511:0] col_in_247,
    input  [511:0] col_in_248,
    input  [511:0] col_in_249,
    input  [511:0] col_in_250,
    input  [511:0] col_in_251,
    input  [511:0] col_in_252,
    input  [511:0] col_in_253,
    input  [511:0] col_in_254,
    input  [511:0] col_in_255,
    input  [511:0] col_in_256,
    input  [511:0] col_in_257,
    input  [511:0] col_in_258,
    input  [511:0] col_in_259,
    input  [511:0] col_in_260,
    input  [511:0] col_in_261,
    input  [511:0] col_in_262,
    input  [511:0] col_in_263,
    input  [511:0] col_in_264,
    input  [511:0] col_in_265,
    input  [511:0] col_in_266,
    input  [511:0] col_in_267,
    input  [511:0] col_in_268,
    input  [511:0] col_in_269,
    input  [511:0] col_in_270,
    input  [511:0] col_in_271,
    input  [511:0] col_in_272,
    input  [511:0] col_in_273,
    input  [511:0] col_in_274,
    input  [511:0] col_in_275,
    input  [511:0] col_in_276,
    input  [511:0] col_in_277,
    input  [511:0] col_in_278,
    input  [511:0] col_in_279,
    input  [511:0] col_in_280,
    input  [511:0] col_in_281,
    input  [511:0] col_in_282,
    input  [511:0] col_in_283,
    input  [511:0] col_in_284,
    input  [511:0] col_in_285,
    input  [511:0] col_in_286,
    input  [511:0] col_in_287,
    input  [511:0] col_in_288,
    input  [511:0] col_in_289,
    input  [511:0] col_in_290,
    input  [511:0] col_in_291,
    input  [511:0] col_in_292,
    input  [511:0] col_in_293,
    input  [511:0] col_in_294,
    input  [511:0] col_in_295,
    input  [511:0] col_in_296,
    input  [511:0] col_in_297,
    input  [511:0] col_in_298,
    input  [511:0] col_in_299,
    input  [511:0] col_in_300,
    input  [511:0] col_in_301,
    input  [511:0] col_in_302,
    input  [511:0] col_in_303,
    input  [511:0] col_in_304,
    input  [511:0] col_in_305,
    input  [511:0] col_in_306,
    input  [511:0] col_in_307,
    input  [511:0] col_in_308,
    input  [511:0] col_in_309,
    input  [511:0] col_in_310,
    input  [511:0] col_in_311,
    input  [511:0] col_in_312,
    input  [511:0] col_in_313,
    input  [511:0] col_in_314,
    input  [511:0] col_in_315,
    input  [511:0] col_in_316,
    input  [511:0] col_in_317,
    input  [511:0] col_in_318,
    input  [511:0] col_in_319,
    input  [511:0] col_in_320,
    input  [511:0] col_in_321,
    input  [511:0] col_in_322,
    input  [511:0] col_in_323,
    input  [511:0] col_in_324,
    input  [511:0] col_in_325,
    input  [511:0] col_in_326,
    input  [511:0] col_in_327,
    input  [511:0] col_in_328,
    input  [511:0] col_in_329,
    input  [511:0] col_in_330,
    input  [511:0] col_in_331,
    input  [511:0] col_in_332,
    input  [511:0] col_in_333,
    input  [511:0] col_in_334,
    input  [511:0] col_in_335,
    input  [511:0] col_in_336,
    input  [511:0] col_in_337,
    input  [511:0] col_in_338,
    input  [511:0] col_in_339,
    input  [511:0] col_in_340,
    input  [511:0] col_in_341,
    input  [511:0] col_in_342,
    input  [511:0] col_in_343,
    input  [511:0] col_in_344,
    input  [511:0] col_in_345,
    input  [511:0] col_in_346,
    input  [511:0] col_in_347,
    input  [511:0] col_in_348,
    input  [511:0] col_in_349,
    input  [511:0] col_in_350,
    input  [511:0] col_in_351,
    input  [511:0] col_in_352,
    input  [511:0] col_in_353,
    input  [511:0] col_in_354,
    input  [511:0] col_in_355,
    input  [511:0] col_in_356,
    input  [511:0] col_in_357,
    input  [511:0] col_in_358,
    input  [511:0] col_in_359,
    input  [511:0] col_in_360,
    input  [511:0] col_in_361,
    input  [511:0] col_in_362,
    input  [511:0] col_in_363,
    input  [511:0] col_in_364,
    input  [511:0] col_in_365,
    input  [511:0] col_in_366,
    input  [511:0] col_in_367,
    input  [511:0] col_in_368,
    input  [511:0] col_in_369,
    input  [511:0] col_in_370,
    input  [511:0] col_in_371,
    input  [511:0] col_in_372,
    input  [511:0] col_in_373,
    input  [511:0] col_in_374,
    input  [511:0] col_in_375,
    input  [511:0] col_in_376,
    input  [511:0] col_in_377,
    input  [511:0] col_in_378,
    input  [511:0] col_in_379,
    input  [511:0] col_in_380,
    input  [511:0] col_in_381,
    input  [511:0] col_in_382,
    input  [511:0] col_in_383,
    input  [511:0] col_in_384,
    input  [511:0] col_in_385,
    input  [511:0] col_in_386,
    input  [511:0] col_in_387,
    input  [511:0] col_in_388,
    input  [511:0] col_in_389,
    input  [511:0] col_in_390,
    input  [511:0] col_in_391,
    input  [511:0] col_in_392,
    input  [511:0] col_in_393,
    input  [511:0] col_in_394,
    input  [511:0] col_in_395,
    input  [511:0] col_in_396,
    input  [511:0] col_in_397,
    input  [511:0] col_in_398,
    input  [511:0] col_in_399,
    input  [511:0] col_in_400,
    input  [511:0] col_in_401,
    input  [511:0] col_in_402,
    input  [511:0] col_in_403,
    input  [511:0] col_in_404,
    input  [511:0] col_in_405,
    input  [511:0] col_in_406,
    input  [511:0] col_in_407,
    input  [511:0] col_in_408,
    input  [511:0] col_in_409,
    input  [511:0] col_in_410,
    input  [511:0] col_in_411,
    input  [511:0] col_in_412,
    input  [511:0] col_in_413,
    input  [511:0] col_in_414,
    input  [511:0] col_in_415,
    input  [511:0] col_in_416,
    input  [511:0] col_in_417,
    input  [511:0] col_in_418,
    input  [511:0] col_in_419,
    input  [511:0] col_in_420,
    input  [511:0] col_in_421,
    input  [511:0] col_in_422,
    input  [511:0] col_in_423,
    input  [511:0] col_in_424,
    input  [511:0] col_in_425,
    input  [511:0] col_in_426,
    input  [511:0] col_in_427,
    input  [511:0] col_in_428,
    input  [511:0] col_in_429,
    input  [511:0] col_in_430,
    input  [511:0] col_in_431,
    input  [511:0] col_in_432,
    input  [511:0] col_in_433,
    input  [511:0] col_in_434,
    input  [511:0] col_in_435,
    input  [511:0] col_in_436,
    input  [511:0] col_in_437,
    input  [511:0] col_in_438,
    input  [511:0] col_in_439,
    input  [511:0] col_in_440,
    input  [511:0] col_in_441,
    input  [511:0] col_in_442,
    input  [511:0] col_in_443,
    input  [511:0] col_in_444,
    input  [511:0] col_in_445,
    input  [511:0] col_in_446,
    input  [511:0] col_in_447,
    input  [511:0] col_in_448,
    input  [511:0] col_in_449,
    input  [511:0] col_in_450,
    input  [511:0] col_in_451,
    input  [511:0] col_in_452,
    input  [511:0] col_in_453,
    input  [511:0] col_in_454,
    input  [511:0] col_in_455,
    input  [511:0] col_in_456,
    input  [511:0] col_in_457,
    input  [511:0] col_in_458,
    input  [511:0] col_in_459,
    input  [511:0] col_in_460,
    input  [511:0] col_in_461,
    input  [511:0] col_in_462,
    input  [511:0] col_in_463,
    input  [511:0] col_in_464,
    input  [511:0] col_in_465,
    input  [511:0] col_in_466,
    input  [511:0] col_in_467,
    input  [511:0] col_in_468,
    input  [511:0] col_in_469,
    input  [511:0] col_in_470,
    input  [511:0] col_in_471,
    input  [511:0] col_in_472,
    input  [511:0] col_in_473,
    input  [511:0] col_in_474,
    input  [511:0] col_in_475,
    input  [511:0] col_in_476,
    input  [511:0] col_in_477,
    input  [511:0] col_in_478,
    input  [511:0] col_in_479,
    input  [511:0] col_in_480,
    input  [511:0] col_in_481,
    input  [511:0] col_in_482,
    input  [511:0] col_in_483,
    input  [511:0] col_in_484,
    input  [511:0] col_in_485,
    input  [511:0] col_in_486,
    input  [511:0] col_in_487,
    input  [511:0] col_in_488,
    input  [511:0] col_in_489,
    input  [511:0] col_in_490,
    input  [511:0] col_in_491,
    input  [511:0] col_in_492,
    input  [511:0] col_in_493,
    input  [511:0] col_in_494,
    input  [511:0] col_in_495,
    input  [511:0] col_in_496,
    input  [511:0] col_in_497,
    input  [511:0] col_in_498,
    input  [511:0] col_in_499,
    input  [511:0] col_in_500,
    input  [511:0] col_in_501,
    input  [511:0] col_in_502,
    input  [511:0] col_in_503,
    input  [511:0] col_in_504,
    input  [511:0] col_in_505,
    input  [511:0] col_in_506,
    input  [511:0] col_in_507,
    input  [511:0] col_in_508,
    input  [511:0] col_in_509,
    input  [511:0] col_in_510,
    input  [511:0] col_in_511,
    input  [511:0] col_in_512,
    input  [511:0] col_in_513,
    input  [511:0] col_in_514,
    input  [511:0] col_in_515,
    input  [511:0] col_in_516,
    input  [511:0] col_in_517,
    input  [511:0] col_in_518,
    input  [511:0] col_in_519,
    input  [511:0] col_in_520,
    input  [511:0] col_in_521,
    input  [511:0] col_in_522,
    input  [511:0] col_in_523,
    input  [511:0] col_in_524,
    input  [511:0] col_in_525,
    input  [511:0] col_in_526,
    input  [511:0] col_in_527,
    input  [511:0] col_in_528,
    input  [511:0] col_in_529,
    input  [511:0] col_in_530,
    input  [511:0] col_in_531,
    input  [511:0] col_in_532,
    input  [511:0] col_in_533,
    input  [511:0] col_in_534,
    input  [511:0] col_in_535,
    input  [511:0] col_in_536,
    input  [511:0] col_in_537,
    input  [511:0] col_in_538,
    input  [511:0] col_in_539,
    input  [511:0] col_in_540,
    input  [511:0] col_in_541,
    input  [511:0] col_in_542,
    input  [511:0] col_in_543,
    input  [511:0] col_in_544,
    input  [511:0] col_in_545,
    input  [511:0] col_in_546,
    input  [511:0] col_in_547,
    input  [511:0] col_in_548,
    input  [511:0] col_in_549,
    input  [511:0] col_in_550,
    input  [511:0] col_in_551,
    input  [511:0] col_in_552,
    input  [511:0] col_in_553,
    input  [511:0] col_in_554,
    input  [511:0] col_in_555,
    input  [511:0] col_in_556,
    input  [511:0] col_in_557,
    input  [511:0] col_in_558,
    input  [511:0] col_in_559,
    input  [511:0] col_in_560,
    input  [511:0] col_in_561,
    input  [511:0] col_in_562,
    input  [511:0] col_in_563,
    input  [511:0] col_in_564,
    input  [511:0] col_in_565,
    input  [511:0] col_in_566,
    input  [511:0] col_in_567,
    input  [511:0] col_in_568,
    input  [511:0] col_in_569,
    input  [511:0] col_in_570,
    input  [511:0] col_in_571,
    input  [511:0] col_in_572,
    input  [511:0] col_in_573,
    input  [511:0] col_in_574,
    input  [511:0] col_in_575,
    input  [511:0] col_in_576,
    input  [511:0] col_in_577,
    input  [511:0] col_in_578,
    input  [511:0] col_in_579,
    input  [511:0] col_in_580,
    input  [511:0] col_in_581,
    input  [511:0] col_in_582,
    input  [511:0] col_in_583,
    input  [511:0] col_in_584,
    input  [511:0] col_in_585,
    input  [511:0] col_in_586,
    input  [511:0] col_in_587,
    input  [511:0] col_in_588,
    input  [511:0] col_in_589,
    input  [511:0] col_in_590,
    input  [511:0] col_in_591,
    input  [511:0] col_in_592,
    input  [511:0] col_in_593,
    input  [511:0] col_in_594,
    input  [511:0] col_in_595,
    input  [511:0] col_in_596,
    input  [511:0] col_in_597,
    input  [511:0] col_in_598,
    input  [511:0] col_in_599,
    input  [511:0] col_in_600,
    input  [511:0] col_in_601,
    input  [511:0] col_in_602,
    input  [511:0] col_in_603,
    input  [511:0] col_in_604,
    input  [511:0] col_in_605,
    input  [511:0] col_in_606,
    input  [511:0] col_in_607,
    input  [511:0] col_in_608,
    input  [511:0] col_in_609,
    input  [511:0] col_in_610,
    input  [511:0] col_in_611,
    input  [511:0] col_in_612,
    input  [511:0] col_in_613,
    input  [511:0] col_in_614,
    input  [511:0] col_in_615,
    input  [511:0] col_in_616,
    input  [511:0] col_in_617,
    input  [511:0] col_in_618,
    input  [511:0] col_in_619,
    input  [511:0] col_in_620,
    input  [511:0] col_in_621,
    input  [511:0] col_in_622,
    input  [511:0] col_in_623,
    input  [511:0] col_in_624,
    input  [511:0] col_in_625,
    input  [511:0] col_in_626,
    input  [511:0] col_in_627,
    input  [511:0] col_in_628,
    input  [511:0] col_in_629,
    input  [511:0] col_in_630,
    input  [511:0] col_in_631,
    input  [511:0] col_in_632,
    input  [511:0] col_in_633,
    input  [511:0] col_in_634,
    input  [511:0] col_in_635,
    input  [511:0] col_in_636,
    input  [511:0] col_in_637,
    input  [511:0] col_in_638,
    input  [511:0] col_in_639,
    input  [511:0] col_in_640,
    input  [511:0] col_in_641,
    input  [511:0] col_in_642,
    input  [511:0] col_in_643,
    input  [511:0] col_in_644,
    input  [511:0] col_in_645,
    input  [511:0] col_in_646,
    input  [511:0] col_in_647,
    input  [511:0] col_in_648,
    input  [511:0] col_in_649,
    input  [511:0] col_in_650,
    input  [511:0] col_in_651,
    input  [511:0] col_in_652,
    input  [511:0] col_in_653,
    input  [511:0] col_in_654,
    input  [511:0] col_in_655,
    input  [511:0] col_in_656,
    input  [511:0] col_in_657,
    input  [511:0] col_in_658,
    input  [511:0] col_in_659,
    input  [511:0] col_in_660,
    input  [511:0] col_in_661,
    input  [511:0] col_in_662,
    input  [511:0] col_in_663,
    input  [511:0] col_in_664,
    input  [511:0] col_in_665,
    input  [511:0] col_in_666,
    input  [511:0] col_in_667,
    input  [511:0] col_in_668,
    input  [511:0] col_in_669,
    input  [511:0] col_in_670,
    input  [511:0] col_in_671,
    input  [511:0] col_in_672,
    input  [511:0] col_in_673,
    input  [511:0] col_in_674,
    input  [511:0] col_in_675,
    input  [511:0] col_in_676,
    input  [511:0] col_in_677,
    input  [511:0] col_in_678,
    input  [511:0] col_in_679,
    input  [511:0] col_in_680,
    input  [511:0] col_in_681,
    input  [511:0] col_in_682,
    input  [511:0] col_in_683,
    input  [511:0] col_in_684,
    input  [511:0] col_in_685,
    input  [511:0] col_in_686,
    input  [511:0] col_in_687,
    input  [511:0] col_in_688,
    input  [511:0] col_in_689,
    input  [511:0] col_in_690,
    input  [511:0] col_in_691,
    input  [511:0] col_in_692,
    input  [511:0] col_in_693,
    input  [511:0] col_in_694,
    input  [511:0] col_in_695,
    input  [511:0] col_in_696,
    input  [511:0] col_in_697,
    input  [511:0] col_in_698,
    input  [511:0] col_in_699,
    input  [511:0] col_in_700,
    input  [511:0] col_in_701,
    input  [511:0] col_in_702,
    input  [511:0] col_in_703,
    input  [511:0] col_in_704,
    input  [511:0] col_in_705,
    input  [511:0] col_in_706,
    input  [511:0] col_in_707,
    input  [511:0] col_in_708,
    input  [511:0] col_in_709,
    input  [511:0] col_in_710,
    input  [511:0] col_in_711,
    input  [511:0] col_in_712,
    input  [511:0] col_in_713,
    input  [511:0] col_in_714,
    input  [511:0] col_in_715,
    input  [511:0] col_in_716,
    input  [511:0] col_in_717,
    input  [511:0] col_in_718,
    input  [511:0] col_in_719,
    input  [511:0] col_in_720,
    input  [511:0] col_in_721,
    input  [511:0] col_in_722,
    input  [511:0] col_in_723,
    input  [511:0] col_in_724,
    input  [511:0] col_in_725,
    input  [511:0] col_in_726,
    input  [511:0] col_in_727,
    input  [511:0] col_in_728,
    input  [511:0] col_in_729,
    input  [511:0] col_in_730,
    input  [511:0] col_in_731,
    input  [511:0] col_in_732,
    input  [511:0] col_in_733,
    input  [511:0] col_in_734,
    input  [511:0] col_in_735,
    input  [511:0] col_in_736,
    input  [511:0] col_in_737,
    input  [511:0] col_in_738,
    input  [511:0] col_in_739,
    input  [511:0] col_in_740,
    input  [511:0] col_in_741,
    input  [511:0] col_in_742,
    input  [511:0] col_in_743,
    input  [511:0] col_in_744,
    input  [511:0] col_in_745,
    input  [511:0] col_in_746,
    input  [511:0] col_in_747,
    input  [511:0] col_in_748,
    input  [511:0] col_in_749,
    input  [511:0] col_in_750,
    input  [511:0] col_in_751,
    input  [511:0] col_in_752,
    input  [511:0] col_in_753,
    input  [511:0] col_in_754,
    input  [511:0] col_in_755,
    input  [511:0] col_in_756,
    input  [511:0] col_in_757,
    input  [511:0] col_in_758,
    input  [511:0] col_in_759,
    input  [511:0] col_in_760,
    input  [511:0] col_in_761,
    input  [511:0] col_in_762,
    input  [511:0] col_in_763,
    input  [511:0] col_in_764,
    input  [511:0] col_in_765,
    input  [511:0] col_in_766,
    input  [511:0] col_in_767,
    input  [511:0] col_in_768,
    input  [511:0] col_in_769,
    input  [511:0] col_in_770,
    input  [511:0] col_in_771,
    input  [511:0] col_in_772,
    input  [511:0] col_in_773,
    input  [511:0] col_in_774,
    input  [511:0] col_in_775,
    input  [511:0] col_in_776,
    input  [511:0] col_in_777,
    input  [511:0] col_in_778,
    input  [511:0] col_in_779,
    input  [511:0] col_in_780,
    input  [511:0] col_in_781,
    input  [511:0] col_in_782,
    input  [511:0] col_in_783,
    input  [511:0] col_in_784,
    input  [511:0] col_in_785,
    input  [511:0] col_in_786,
    input  [511:0] col_in_787,
    input  [511:0] col_in_788,
    input  [511:0] col_in_789,
    input  [511:0] col_in_790,
    input  [511:0] col_in_791,
    input  [511:0] col_in_792,
    input  [511:0] col_in_793,
    input  [511:0] col_in_794,
    input  [511:0] col_in_795,
    input  [511:0] col_in_796,
    input  [511:0] col_in_797,
    input  [511:0] col_in_798,
    input  [511:0] col_in_799,
    input  [511:0] col_in_800,
    input  [511:0] col_in_801,
    input  [511:0] col_in_802,
    input  [511:0] col_in_803,
    input  [511:0] col_in_804,
    input  [511:0] col_in_805,
    input  [511:0] col_in_806,
    input  [511:0] col_in_807,
    input  [511:0] col_in_808,
    input  [511:0] col_in_809,
    input  [511:0] col_in_810,
    input  [511:0] col_in_811,
    input  [511:0] col_in_812,
    input  [511:0] col_in_813,
    input  [511:0] col_in_814,
    input  [511:0] col_in_815,
    input  [511:0] col_in_816,
    input  [511:0] col_in_817,
    input  [511:0] col_in_818,
    input  [511:0] col_in_819,
    input  [511:0] col_in_820,
    input  [511:0] col_in_821,
    input  [511:0] col_in_822,
    input  [511:0] col_in_823,
    input  [511:0] col_in_824,
    input  [511:0] col_in_825,
    input  [511:0] col_in_826,
    input  [511:0] col_in_827,
    input  [511:0] col_in_828,
    input  [511:0] col_in_829,
    input  [511:0] col_in_830,
    input  [511:0] col_in_831,
    input  [511:0] col_in_832,
    input  [511:0] col_in_833,
    input  [511:0] col_in_834,
    input  [511:0] col_in_835,
    input  [511:0] col_in_836,
    input  [511:0] col_in_837,
    input  [511:0] col_in_838,
    input  [511:0] col_in_839,
    input  [511:0] col_in_840,
    input  [511:0] col_in_841,
    input  [511:0] col_in_842,
    input  [511:0] col_in_843,
    input  [511:0] col_in_844,
    input  [511:0] col_in_845,
    input  [511:0] col_in_846,
    input  [511:0] col_in_847,
    input  [511:0] col_in_848,
    input  [511:0] col_in_849,
    input  [511:0] col_in_850,
    input  [511:0] col_in_851,
    input  [511:0] col_in_852,
    input  [511:0] col_in_853,
    input  [511:0] col_in_854,
    input  [511:0] col_in_855,
    input  [511:0] col_in_856,
    input  [511:0] col_in_857,
    input  [511:0] col_in_858,
    input  [511:0] col_in_859,
    input  [511:0] col_in_860,
    input  [511:0] col_in_861,
    input  [511:0] col_in_862,
    input  [511:0] col_in_863,
    input  [511:0] col_in_864,
    input  [511:0] col_in_865,
    input  [511:0] col_in_866,
    input  [511:0] col_in_867,
    input  [511:0] col_in_868,
    input  [511:0] col_in_869,
    input  [511:0] col_in_870,
    input  [511:0] col_in_871,
    input  [511:0] col_in_872,
    input  [511:0] col_in_873,
    input  [511:0] col_in_874,
    input  [511:0] col_in_875,
    input  [511:0] col_in_876,
    input  [511:0] col_in_877,
    input  [511:0] col_in_878,
    input  [511:0] col_in_879,
    input  [511:0] col_in_880,
    input  [511:0] col_in_881,
    input  [511:0] col_in_882,
    input  [511:0] col_in_883,
    input  [511:0] col_in_884,
    input  [511:0] col_in_885,
    input  [511:0] col_in_886,
    input  [511:0] col_in_887,
    input  [511:0] col_in_888,
    input  [511:0] col_in_889,
    input  [511:0] col_in_890,
    input  [511:0] col_in_891,
    input  [511:0] col_in_892,
    input  [511:0] col_in_893,
    input  [511:0] col_in_894,
    input  [511:0] col_in_895,
    input  [511:0] col_in_896,
    input  [511:0] col_in_897,
    input  [511:0] col_in_898,
    input  [511:0] col_in_899,
    input  [511:0] col_in_900,
    input  [511:0] col_in_901,
    input  [511:0] col_in_902,
    input  [511:0] col_in_903,
    input  [511:0] col_in_904,
    input  [511:0] col_in_905,
    input  [511:0] col_in_906,
    input  [511:0] col_in_907,
    input  [511:0] col_in_908,
    input  [511:0] col_in_909,
    input  [511:0] col_in_910,
    input  [511:0] col_in_911,
    input  [511:0] col_in_912,
    input  [511:0] col_in_913,
    input  [511:0] col_in_914,
    input  [511:0] col_in_915,
    input  [511:0] col_in_916,
    input  [511:0] col_in_917,
    input  [511:0] col_in_918,
    input  [511:0] col_in_919,
    input  [511:0] col_in_920,
    input  [511:0] col_in_921,
    input  [511:0] col_in_922,
    input  [511:0] col_in_923,
    input  [511:0] col_in_924,
    input  [511:0] col_in_925,
    input  [511:0] col_in_926,
    input  [511:0] col_in_927,
    input  [511:0] col_in_928,
    input  [511:0] col_in_929,
    input  [511:0] col_in_930,
    input  [511:0] col_in_931,
    input  [511:0] col_in_932,
    input  [511:0] col_in_933,
    input  [511:0] col_in_934,
    input  [511:0] col_in_935,
    input  [511:0] col_in_936,
    input  [511:0] col_in_937,
    input  [511:0] col_in_938,
    input  [511:0] col_in_939,
    input  [511:0] col_in_940,
    input  [511:0] col_in_941,
    input  [511:0] col_in_942,
    input  [511:0] col_in_943,
    input  [511:0] col_in_944,
    input  [511:0] col_in_945,
    input  [511:0] col_in_946,
    input  [511:0] col_in_947,
    input  [511:0] col_in_948,
    input  [511:0] col_in_949,
    input  [511:0] col_in_950,
    input  [511:0] col_in_951,
    input  [511:0] col_in_952,
    input  [511:0] col_in_953,
    input  [511:0] col_in_954,
    input  [511:0] col_in_955,
    input  [511:0] col_in_956,
    input  [511:0] col_in_957,
    input  [511:0] col_in_958,
    input  [511:0] col_in_959,
    input  [511:0] col_in_960,
    input  [511:0] col_in_961,
    input  [511:0] col_in_962,
    input  [511:0] col_in_963,
    input  [511:0] col_in_964,
    input  [511:0] col_in_965,
    input  [511:0] col_in_966,
    input  [511:0] col_in_967,
    input  [511:0] col_in_968,
    input  [511:0] col_in_969,
    input  [511:0] col_in_970,
    input  [511:0] col_in_971,
    input  [511:0] col_in_972,
    input  [511:0] col_in_973,
    input  [511:0] col_in_974,
    input  [511:0] col_in_975,
    input  [511:0] col_in_976,
    input  [511:0] col_in_977,
    input  [511:0] col_in_978,
    input  [511:0] col_in_979,
    input  [511:0] col_in_980,
    input  [511:0] col_in_981,
    input  [511:0] col_in_982,
    input  [511:0] col_in_983,
    input  [511:0] col_in_984,
    input  [511:0] col_in_985,
    input  [511:0] col_in_986,
    input  [511:0] col_in_987,
    input  [511:0] col_in_988,
    input  [511:0] col_in_989,
    input  [511:0] col_in_990,
    input  [511:0] col_in_991,
    input  [511:0] col_in_992,
    input  [511:0] col_in_993,
    input  [511:0] col_in_994,
    input  [511:0] col_in_995,
    input  [511:0] col_in_996,
    input  [511:0] col_in_997,
    input  [511:0] col_in_998,
    input  [511:0] col_in_999,
    input  [511:0] col_in_1000,
    input  [511:0] col_in_1001,
    input  [511:0] col_in_1002,
    input  [511:0] col_in_1003,
    input  [511:0] col_in_1004,
    input  [511:0] col_in_1005,
    input  [511:0] col_in_1006,
    input  [511:0] col_in_1007,
    input  [511:0] col_in_1008,
    input  [511:0] col_in_1009,
    input  [511:0] col_in_1010,
    input  [511:0] col_in_1011,
    input  [511:0] col_in_1012,
    input  [511:0] col_in_1013,
    input  [511:0] col_in_1014,
    input  [511:0] col_in_1015,
    input  [511:0] col_in_1016,
    input  [511:0] col_in_1017,
    input  [511:0] col_in_1018,
    input  [511:0] col_in_1019,
    input  [511:0] col_in_1020,
    input  [511:0] col_in_1021,
    input  [511:0] col_in_1022,
    input  [511:0] col_in_1023,

    output  [1032:0]  compressor_array_512_out0,
    output  [1032:0]  compressor_array_512_out1,

    output  [1024:0]  data_out_0,
    output  [1024:0]  data_out_1
);










compressor_array_512_2_1024_row  u0_compressor_array_512_2_1024_row (
    .col_in_0                ( col_in_0      ),
    .col_in_1                ( col_in_1      ),
    .col_in_2                ( col_in_2      ),
    .col_in_3                ( col_in_3      ),
    .col_in_4                ( col_in_4      ),
    .col_in_5                ( col_in_5      ),
    .col_in_6                ( col_in_6      ),
    .col_in_7                ( col_in_7      ),
    .col_in_8                ( col_in_8      ),
    .col_in_9                ( col_in_9      ),
    .col_in_10               ( col_in_10     ),
    .col_in_11               ( col_in_11     ),
    .col_in_12               ( col_in_12     ),
    .col_in_13               ( col_in_13     ),
    .col_in_14               ( col_in_14     ),
    .col_in_15               ( col_in_15     ),
    .col_in_16               ( col_in_16     ),
    .col_in_17               ( col_in_17     ),
    .col_in_18               ( col_in_18     ),
    .col_in_19               ( col_in_19     ),
    .col_in_20               ( col_in_20     ),
    .col_in_21               ( col_in_21     ),
    .col_in_22               ( col_in_22     ),
    .col_in_23               ( col_in_23     ),
    .col_in_24               ( col_in_24     ),
    .col_in_25               ( col_in_25     ),
    .col_in_26               ( col_in_26     ),
    .col_in_27               ( col_in_27     ),
    .col_in_28               ( col_in_28     ),
    .col_in_29               ( col_in_29     ),
    .col_in_30               ( col_in_30     ),
    .col_in_31               ( col_in_31     ),
    .col_in_32               ( col_in_32     ),
    .col_in_33               ( col_in_33     ),
    .col_in_34               ( col_in_34     ),
    .col_in_35               ( col_in_35     ),
    .col_in_36               ( col_in_36     ),
    .col_in_37               ( col_in_37     ),
    .col_in_38               ( col_in_38     ),
    .col_in_39               ( col_in_39     ),
    .col_in_40               ( col_in_40     ),
    .col_in_41               ( col_in_41     ),
    .col_in_42               ( col_in_42     ),
    .col_in_43               ( col_in_43     ),
    .col_in_44               ( col_in_44     ),
    .col_in_45               ( col_in_45     ),
    .col_in_46               ( col_in_46     ),
    .col_in_47               ( col_in_47     ),
    .col_in_48               ( col_in_48     ),
    .col_in_49               ( col_in_49     ),
    .col_in_50               ( col_in_50     ),
    .col_in_51               ( col_in_51     ),
    .col_in_52               ( col_in_52     ),
    .col_in_53               ( col_in_53     ),
    .col_in_54               ( col_in_54     ),
    .col_in_55               ( col_in_55     ),
    .col_in_56               ( col_in_56     ),
    .col_in_57               ( col_in_57     ),
    .col_in_58               ( col_in_58     ),
    .col_in_59               ( col_in_59     ),
    .col_in_60               ( col_in_60     ),
    .col_in_61               ( col_in_61     ),
    .col_in_62               ( col_in_62     ),
    .col_in_63               ( col_in_63     ),
    .col_in_64               ( col_in_64     ),
    .col_in_65               ( col_in_65     ),
    .col_in_66               ( col_in_66     ),
    .col_in_67               ( col_in_67     ),
    .col_in_68               ( col_in_68     ),
    .col_in_69               ( col_in_69     ),
    .col_in_70               ( col_in_70     ),
    .col_in_71               ( col_in_71     ),
    .col_in_72               ( col_in_72     ),
    .col_in_73               ( col_in_73     ),
    .col_in_74               ( col_in_74     ),
    .col_in_75               ( col_in_75     ),
    .col_in_76               ( col_in_76     ),
    .col_in_77               ( col_in_77     ),
    .col_in_78               ( col_in_78     ),
    .col_in_79               ( col_in_79     ),
    .col_in_80               ( col_in_80     ),
    .col_in_81               ( col_in_81     ),
    .col_in_82               ( col_in_82     ),
    .col_in_83               ( col_in_83     ),
    .col_in_84               ( col_in_84     ),
    .col_in_85               ( col_in_85     ),
    .col_in_86               ( col_in_86     ),
    .col_in_87               ( col_in_87     ),
    .col_in_88               ( col_in_88     ),
    .col_in_89               ( col_in_89     ),
    .col_in_90               ( col_in_90     ),
    .col_in_91               ( col_in_91     ),
    .col_in_92               ( col_in_92     ),
    .col_in_93               ( col_in_93     ),
    .col_in_94               ( col_in_94     ),
    .col_in_95               ( col_in_95     ),
    .col_in_96               ( col_in_96     ),
    .col_in_97               ( col_in_97     ),
    .col_in_98               ( col_in_98     ),
    .col_in_99               ( col_in_99     ),
    .col_in_100              ( col_in_100    ),
    .col_in_101              ( col_in_101    ),
    .col_in_102              ( col_in_102    ),
    .col_in_103              ( col_in_103    ),
    .col_in_104              ( col_in_104    ),
    .col_in_105              ( col_in_105    ),
    .col_in_106              ( col_in_106    ),
    .col_in_107              ( col_in_107    ),
    .col_in_108              ( col_in_108    ),
    .col_in_109              ( col_in_109    ),
    .col_in_110              ( col_in_110    ),
    .col_in_111              ( col_in_111    ),
    .col_in_112              ( col_in_112    ),
    .col_in_113              ( col_in_113    ),
    .col_in_114              ( col_in_114    ),
    .col_in_115              ( col_in_115    ),
    .col_in_116              ( col_in_116    ),
    .col_in_117              ( col_in_117    ),
    .col_in_118              ( col_in_118    ),
    .col_in_119              ( col_in_119    ),
    .col_in_120              ( col_in_120    ),
    .col_in_121              ( col_in_121    ),
    .col_in_122              ( col_in_122    ),
    .col_in_123              ( col_in_123    ),
    .col_in_124              ( col_in_124    ),
    .col_in_125              ( col_in_125    ),
    .col_in_126              ( col_in_126    ),
    .col_in_127              ( col_in_127    ),
    .col_in_128              ( col_in_128    ),
    .col_in_129              ( col_in_129    ),
    .col_in_130              ( col_in_130    ),
    .col_in_131              ( col_in_131    ),
    .col_in_132              ( col_in_132    ),
    .col_in_133              ( col_in_133    ),
    .col_in_134              ( col_in_134    ),
    .col_in_135              ( col_in_135    ),
    .col_in_136              ( col_in_136    ),
    .col_in_137              ( col_in_137    ),
    .col_in_138              ( col_in_138    ),
    .col_in_139              ( col_in_139    ),
    .col_in_140              ( col_in_140    ),
    .col_in_141              ( col_in_141    ),
    .col_in_142              ( col_in_142    ),
    .col_in_143              ( col_in_143    ),
    .col_in_144              ( col_in_144    ),
    .col_in_145              ( col_in_145    ),
    .col_in_146              ( col_in_146    ),
    .col_in_147              ( col_in_147    ),
    .col_in_148              ( col_in_148    ),
    .col_in_149              ( col_in_149    ),
    .col_in_150              ( col_in_150    ),
    .col_in_151              ( col_in_151    ),
    .col_in_152              ( col_in_152    ),
    .col_in_153              ( col_in_153    ),
    .col_in_154              ( col_in_154    ),
    .col_in_155              ( col_in_155    ),
    .col_in_156              ( col_in_156    ),
    .col_in_157              ( col_in_157    ),
    .col_in_158              ( col_in_158    ),
    .col_in_159              ( col_in_159    ),
    .col_in_160              ( col_in_160    ),
    .col_in_161              ( col_in_161    ),
    .col_in_162              ( col_in_162    ),
    .col_in_163              ( col_in_163    ),
    .col_in_164              ( col_in_164    ),
    .col_in_165              ( col_in_165    ),
    .col_in_166              ( col_in_166    ),
    .col_in_167              ( col_in_167    ),
    .col_in_168              ( col_in_168    ),
    .col_in_169              ( col_in_169    ),
    .col_in_170              ( col_in_170    ),
    .col_in_171              ( col_in_171    ),
    .col_in_172              ( col_in_172    ),
    .col_in_173              ( col_in_173    ),
    .col_in_174              ( col_in_174    ),
    .col_in_175              ( col_in_175    ),
    .col_in_176              ( col_in_176    ),
    .col_in_177              ( col_in_177    ),
    .col_in_178              ( col_in_178    ),
    .col_in_179              ( col_in_179    ),
    .col_in_180              ( col_in_180    ),
    .col_in_181              ( col_in_181    ),
    .col_in_182              ( col_in_182    ),
    .col_in_183              ( col_in_183    ),
    .col_in_184              ( col_in_184    ),
    .col_in_185              ( col_in_185    ),
    .col_in_186              ( col_in_186    ),
    .col_in_187              ( col_in_187    ),
    .col_in_188              ( col_in_188    ),
    .col_in_189              ( col_in_189    ),
    .col_in_190              ( col_in_190    ),
    .col_in_191              ( col_in_191    ),
    .col_in_192              ( col_in_192    ),
    .col_in_193              ( col_in_193    ),
    .col_in_194              ( col_in_194    ),
    .col_in_195              ( col_in_195    ),
    .col_in_196              ( col_in_196    ),
    .col_in_197              ( col_in_197    ),
    .col_in_198              ( col_in_198    ),
    .col_in_199              ( col_in_199    ),
    .col_in_200              ( col_in_200    ),
    .col_in_201              ( col_in_201    ),
    .col_in_202              ( col_in_202    ),
    .col_in_203              ( col_in_203    ),
    .col_in_204              ( col_in_204    ),
    .col_in_205              ( col_in_205    ),
    .col_in_206              ( col_in_206    ),
    .col_in_207              ( col_in_207    ),
    .col_in_208              ( col_in_208    ),
    .col_in_209              ( col_in_209    ),
    .col_in_210              ( col_in_210    ),
    .col_in_211              ( col_in_211    ),
    .col_in_212              ( col_in_212    ),
    .col_in_213              ( col_in_213    ),
    .col_in_214              ( col_in_214    ),
    .col_in_215              ( col_in_215    ),
    .col_in_216              ( col_in_216    ),
    .col_in_217              ( col_in_217    ),
    .col_in_218              ( col_in_218    ),
    .col_in_219              ( col_in_219    ),
    .col_in_220              ( col_in_220    ),
    .col_in_221              ( col_in_221    ),
    .col_in_222              ( col_in_222    ),
    .col_in_223              ( col_in_223    ),
    .col_in_224              ( col_in_224    ),
    .col_in_225              ( col_in_225    ),
    .col_in_226              ( col_in_226    ),
    .col_in_227              ( col_in_227    ),
    .col_in_228              ( col_in_228    ),
    .col_in_229              ( col_in_229    ),
    .col_in_230              ( col_in_230    ),
    .col_in_231              ( col_in_231    ),
    .col_in_232              ( col_in_232    ),
    .col_in_233              ( col_in_233    ),
    .col_in_234              ( col_in_234    ),
    .col_in_235              ( col_in_235    ),
    .col_in_236              ( col_in_236    ),
    .col_in_237              ( col_in_237    ),
    .col_in_238              ( col_in_238    ),
    .col_in_239              ( col_in_239    ),
    .col_in_240              ( col_in_240    ),
    .col_in_241              ( col_in_241    ),
    .col_in_242              ( col_in_242    ),
    .col_in_243              ( col_in_243    ),
    .col_in_244              ( col_in_244    ),
    .col_in_245              ( col_in_245    ),
    .col_in_246              ( col_in_246    ),
    .col_in_247              ( col_in_247    ),
    .col_in_248              ( col_in_248    ),
    .col_in_249              ( col_in_249    ),
    .col_in_250              ( col_in_250    ),
    .col_in_251              ( col_in_251    ),
    .col_in_252              ( col_in_252    ),
    .col_in_253              ( col_in_253    ),
    .col_in_254              ( col_in_254    ),
    .col_in_255              ( col_in_255    ),
    .col_in_256              ( col_in_256    ),
    .col_in_257              ( col_in_257    ),
    .col_in_258              ( col_in_258    ),
    .col_in_259              ( col_in_259    ),
    .col_in_260              ( col_in_260    ),
    .col_in_261              ( col_in_261    ),
    .col_in_262              ( col_in_262    ),
    .col_in_263              ( col_in_263    ),
    .col_in_264              ( col_in_264    ),
    .col_in_265              ( col_in_265    ),
    .col_in_266              ( col_in_266    ),
    .col_in_267              ( col_in_267    ),
    .col_in_268              ( col_in_268    ),
    .col_in_269              ( col_in_269    ),
    .col_in_270              ( col_in_270    ),
    .col_in_271              ( col_in_271    ),
    .col_in_272              ( col_in_272    ),
    .col_in_273              ( col_in_273    ),
    .col_in_274              ( col_in_274    ),
    .col_in_275              ( col_in_275    ),
    .col_in_276              ( col_in_276    ),
    .col_in_277              ( col_in_277    ),
    .col_in_278              ( col_in_278    ),
    .col_in_279              ( col_in_279    ),
    .col_in_280              ( col_in_280    ),
    .col_in_281              ( col_in_281    ),
    .col_in_282              ( col_in_282    ),
    .col_in_283              ( col_in_283    ),
    .col_in_284              ( col_in_284    ),
    .col_in_285              ( col_in_285    ),
    .col_in_286              ( col_in_286    ),
    .col_in_287              ( col_in_287    ),
    .col_in_288              ( col_in_288    ),
    .col_in_289              ( col_in_289    ),
    .col_in_290              ( col_in_290    ),
    .col_in_291              ( col_in_291    ),
    .col_in_292              ( col_in_292    ),
    .col_in_293              ( col_in_293    ),
    .col_in_294              ( col_in_294    ),
    .col_in_295              ( col_in_295    ),
    .col_in_296              ( col_in_296    ),
    .col_in_297              ( col_in_297    ),
    .col_in_298              ( col_in_298    ),
    .col_in_299              ( col_in_299    ),
    .col_in_300              ( col_in_300    ),
    .col_in_301              ( col_in_301    ),
    .col_in_302              ( col_in_302    ),
    .col_in_303              ( col_in_303    ),
    .col_in_304              ( col_in_304    ),
    .col_in_305              ( col_in_305    ),
    .col_in_306              ( col_in_306    ),
    .col_in_307              ( col_in_307    ),
    .col_in_308              ( col_in_308    ),
    .col_in_309              ( col_in_309    ),
    .col_in_310              ( col_in_310    ),
    .col_in_311              ( col_in_311    ),
    .col_in_312              ( col_in_312    ),
    .col_in_313              ( col_in_313    ),
    .col_in_314              ( col_in_314    ),
    .col_in_315              ( col_in_315    ),
    .col_in_316              ( col_in_316    ),
    .col_in_317              ( col_in_317    ),
    .col_in_318              ( col_in_318    ),
    .col_in_319              ( col_in_319    ),
    .col_in_320              ( col_in_320    ),
    .col_in_321              ( col_in_321    ),
    .col_in_322              ( col_in_322    ),
    .col_in_323              ( col_in_323    ),
    .col_in_324              ( col_in_324    ),
    .col_in_325              ( col_in_325    ),
    .col_in_326              ( col_in_326    ),
    .col_in_327              ( col_in_327    ),
    .col_in_328              ( col_in_328    ),
    .col_in_329              ( col_in_329    ),
    .col_in_330              ( col_in_330    ),
    .col_in_331              ( col_in_331    ),
    .col_in_332              ( col_in_332    ),
    .col_in_333              ( col_in_333    ),
    .col_in_334              ( col_in_334    ),
    .col_in_335              ( col_in_335    ),
    .col_in_336              ( col_in_336    ),
    .col_in_337              ( col_in_337    ),
    .col_in_338              ( col_in_338    ),
    .col_in_339              ( col_in_339    ),
    .col_in_340              ( col_in_340    ),
    .col_in_341              ( col_in_341    ),
    .col_in_342              ( col_in_342    ),
    .col_in_343              ( col_in_343    ),
    .col_in_344              ( col_in_344    ),
    .col_in_345              ( col_in_345    ),
    .col_in_346              ( col_in_346    ),
    .col_in_347              ( col_in_347    ),
    .col_in_348              ( col_in_348    ),
    .col_in_349              ( col_in_349    ),
    .col_in_350              ( col_in_350    ),
    .col_in_351              ( col_in_351    ),
    .col_in_352              ( col_in_352    ),
    .col_in_353              ( col_in_353    ),
    .col_in_354              ( col_in_354    ),
    .col_in_355              ( col_in_355    ),
    .col_in_356              ( col_in_356    ),
    .col_in_357              ( col_in_357    ),
    .col_in_358              ( col_in_358    ),
    .col_in_359              ( col_in_359    ),
    .col_in_360              ( col_in_360    ),
    .col_in_361              ( col_in_361    ),
    .col_in_362              ( col_in_362    ),
    .col_in_363              ( col_in_363    ),
    .col_in_364              ( col_in_364    ),
    .col_in_365              ( col_in_365    ),
    .col_in_366              ( col_in_366    ),
    .col_in_367              ( col_in_367    ),
    .col_in_368              ( col_in_368    ),
    .col_in_369              ( col_in_369    ),
    .col_in_370              ( col_in_370    ),
    .col_in_371              ( col_in_371    ),
    .col_in_372              ( col_in_372    ),
    .col_in_373              ( col_in_373    ),
    .col_in_374              ( col_in_374    ),
    .col_in_375              ( col_in_375    ),
    .col_in_376              ( col_in_376    ),
    .col_in_377              ( col_in_377    ),
    .col_in_378              ( col_in_378    ),
    .col_in_379              ( col_in_379    ),
    .col_in_380              ( col_in_380    ),
    .col_in_381              ( col_in_381    ),
    .col_in_382              ( col_in_382    ),
    .col_in_383              ( col_in_383    ),
    .col_in_384              ( col_in_384    ),
    .col_in_385              ( col_in_385    ),
    .col_in_386              ( col_in_386    ),
    .col_in_387              ( col_in_387    ),
    .col_in_388              ( col_in_388    ),
    .col_in_389              ( col_in_389    ),
    .col_in_390              ( col_in_390    ),
    .col_in_391              ( col_in_391    ),
    .col_in_392              ( col_in_392    ),
    .col_in_393              ( col_in_393    ),
    .col_in_394              ( col_in_394    ),
    .col_in_395              ( col_in_395    ),
    .col_in_396              ( col_in_396    ),
    .col_in_397              ( col_in_397    ),
    .col_in_398              ( col_in_398    ),
    .col_in_399              ( col_in_399    ),
    .col_in_400              ( col_in_400    ),
    .col_in_401              ( col_in_401    ),
    .col_in_402              ( col_in_402    ),
    .col_in_403              ( col_in_403    ),
    .col_in_404              ( col_in_404    ),
    .col_in_405              ( col_in_405    ),
    .col_in_406              ( col_in_406    ),
    .col_in_407              ( col_in_407    ),
    .col_in_408              ( col_in_408    ),
    .col_in_409              ( col_in_409    ),
    .col_in_410              ( col_in_410    ),
    .col_in_411              ( col_in_411    ),
    .col_in_412              ( col_in_412    ),
    .col_in_413              ( col_in_413    ),
    .col_in_414              ( col_in_414    ),
    .col_in_415              ( col_in_415    ),
    .col_in_416              ( col_in_416    ),
    .col_in_417              ( col_in_417    ),
    .col_in_418              ( col_in_418    ),
    .col_in_419              ( col_in_419    ),
    .col_in_420              ( col_in_420    ),
    .col_in_421              ( col_in_421    ),
    .col_in_422              ( col_in_422    ),
    .col_in_423              ( col_in_423    ),
    .col_in_424              ( col_in_424    ),
    .col_in_425              ( col_in_425    ),
    .col_in_426              ( col_in_426    ),
    .col_in_427              ( col_in_427    ),
    .col_in_428              ( col_in_428    ),
    .col_in_429              ( col_in_429    ),
    .col_in_430              ( col_in_430    ),
    .col_in_431              ( col_in_431    ),
    .col_in_432              ( col_in_432    ),
    .col_in_433              ( col_in_433    ),
    .col_in_434              ( col_in_434    ),
    .col_in_435              ( col_in_435    ),
    .col_in_436              ( col_in_436    ),
    .col_in_437              ( col_in_437    ),
    .col_in_438              ( col_in_438    ),
    .col_in_439              ( col_in_439    ),
    .col_in_440              ( col_in_440    ),
    .col_in_441              ( col_in_441    ),
    .col_in_442              ( col_in_442    ),
    .col_in_443              ( col_in_443    ),
    .col_in_444              ( col_in_444    ),
    .col_in_445              ( col_in_445    ),
    .col_in_446              ( col_in_446    ),
    .col_in_447              ( col_in_447    ),
    .col_in_448              ( col_in_448    ),
    .col_in_449              ( col_in_449    ),
    .col_in_450              ( col_in_450    ),
    .col_in_451              ( col_in_451    ),
    .col_in_452              ( col_in_452    ),
    .col_in_453              ( col_in_453    ),
    .col_in_454              ( col_in_454    ),
    .col_in_455              ( col_in_455    ),
    .col_in_456              ( col_in_456    ),
    .col_in_457              ( col_in_457    ),
    .col_in_458              ( col_in_458    ),
    .col_in_459              ( col_in_459    ),
    .col_in_460              ( col_in_460    ),
    .col_in_461              ( col_in_461    ),
    .col_in_462              ( col_in_462    ),
    .col_in_463              ( col_in_463    ),
    .col_in_464              ( col_in_464    ),
    .col_in_465              ( col_in_465    ),
    .col_in_466              ( col_in_466    ),
    .col_in_467              ( col_in_467    ),
    .col_in_468              ( col_in_468    ),
    .col_in_469              ( col_in_469    ),
    .col_in_470              ( col_in_470    ),
    .col_in_471              ( col_in_471    ),
    .col_in_472              ( col_in_472    ),
    .col_in_473              ( col_in_473    ),
    .col_in_474              ( col_in_474    ),
    .col_in_475              ( col_in_475    ),
    .col_in_476              ( col_in_476    ),
    .col_in_477              ( col_in_477    ),
    .col_in_478              ( col_in_478    ),
    .col_in_479              ( col_in_479    ),
    .col_in_480              ( col_in_480    ),
    .col_in_481              ( col_in_481    ),
    .col_in_482              ( col_in_482    ),
    .col_in_483              ( col_in_483    ),
    .col_in_484              ( col_in_484    ),
    .col_in_485              ( col_in_485    ),
    .col_in_486              ( col_in_486    ),
    .col_in_487              ( col_in_487    ),
    .col_in_488              ( col_in_488    ),
    .col_in_489              ( col_in_489    ),
    .col_in_490              ( col_in_490    ),
    .col_in_491              ( col_in_491    ),
    .col_in_492              ( col_in_492    ),
    .col_in_493              ( col_in_493    ),
    .col_in_494              ( col_in_494    ),
    .col_in_495              ( col_in_495    ),
    .col_in_496              ( col_in_496    ),
    .col_in_497              ( col_in_497    ),
    .col_in_498              ( col_in_498    ),
    .col_in_499              ( col_in_499    ),
    .col_in_500              ( col_in_500    ),
    .col_in_501              ( col_in_501    ),
    .col_in_502              ( col_in_502    ),
    .col_in_503              ( col_in_503    ),
    .col_in_504              ( col_in_504    ),
    .col_in_505              ( col_in_505    ),
    .col_in_506              ( col_in_506    ),
    .col_in_507              ( col_in_507    ),
    .col_in_508              ( col_in_508    ),
    .col_in_509              ( col_in_509    ),
    .col_in_510              ( col_in_510    ),
    .col_in_511              ( col_in_511    ),
    .col_in_512              ( col_in_512    ),
    .col_in_513              ( col_in_513    ),
    .col_in_514              ( col_in_514    ),
    .col_in_515              ( col_in_515    ),
    .col_in_516              ( col_in_516    ),
    .col_in_517              ( col_in_517    ),
    .col_in_518              ( col_in_518    ),
    .col_in_519              ( col_in_519    ),
    .col_in_520              ( col_in_520    ),
    .col_in_521              ( col_in_521    ),
    .col_in_522              ( col_in_522    ),
    .col_in_523              ( col_in_523    ),
    .col_in_524              ( col_in_524    ),
    .col_in_525              ( col_in_525    ),
    .col_in_526              ( col_in_526    ),
    .col_in_527              ( col_in_527    ),
    .col_in_528              ( col_in_528    ),
    .col_in_529              ( col_in_529    ),
    .col_in_530              ( col_in_530    ),
    .col_in_531              ( col_in_531    ),
    .col_in_532              ( col_in_532    ),
    .col_in_533              ( col_in_533    ),
    .col_in_534              ( col_in_534    ),
    .col_in_535              ( col_in_535    ),
    .col_in_536              ( col_in_536    ),
    .col_in_537              ( col_in_537    ),
    .col_in_538              ( col_in_538    ),
    .col_in_539              ( col_in_539    ),
    .col_in_540              ( col_in_540    ),
    .col_in_541              ( col_in_541    ),
    .col_in_542              ( col_in_542    ),
    .col_in_543              ( col_in_543    ),
    .col_in_544              ( col_in_544    ),
    .col_in_545              ( col_in_545    ),
    .col_in_546              ( col_in_546    ),
    .col_in_547              ( col_in_547    ),
    .col_in_548              ( col_in_548    ),
    .col_in_549              ( col_in_549    ),
    .col_in_550              ( col_in_550    ),
    .col_in_551              ( col_in_551    ),
    .col_in_552              ( col_in_552    ),
    .col_in_553              ( col_in_553    ),
    .col_in_554              ( col_in_554    ),
    .col_in_555              ( col_in_555    ),
    .col_in_556              ( col_in_556    ),
    .col_in_557              ( col_in_557    ),
    .col_in_558              ( col_in_558    ),
    .col_in_559              ( col_in_559    ),
    .col_in_560              ( col_in_560    ),
    .col_in_561              ( col_in_561    ),
    .col_in_562              ( col_in_562    ),
    .col_in_563              ( col_in_563    ),
    .col_in_564              ( col_in_564    ),
    .col_in_565              ( col_in_565    ),
    .col_in_566              ( col_in_566    ),
    .col_in_567              ( col_in_567    ),
    .col_in_568              ( col_in_568    ),
    .col_in_569              ( col_in_569    ),
    .col_in_570              ( col_in_570    ),
    .col_in_571              ( col_in_571    ),
    .col_in_572              ( col_in_572    ),
    .col_in_573              ( col_in_573    ),
    .col_in_574              ( col_in_574    ),
    .col_in_575              ( col_in_575    ),
    .col_in_576              ( col_in_576    ),
    .col_in_577              ( col_in_577    ),
    .col_in_578              ( col_in_578    ),
    .col_in_579              ( col_in_579    ),
    .col_in_580              ( col_in_580    ),
    .col_in_581              ( col_in_581    ),
    .col_in_582              ( col_in_582    ),
    .col_in_583              ( col_in_583    ),
    .col_in_584              ( col_in_584    ),
    .col_in_585              ( col_in_585    ),
    .col_in_586              ( col_in_586    ),
    .col_in_587              ( col_in_587    ),
    .col_in_588              ( col_in_588    ),
    .col_in_589              ( col_in_589    ),
    .col_in_590              ( col_in_590    ),
    .col_in_591              ( col_in_591    ),
    .col_in_592              ( col_in_592    ),
    .col_in_593              ( col_in_593    ),
    .col_in_594              ( col_in_594    ),
    .col_in_595              ( col_in_595    ),
    .col_in_596              ( col_in_596    ),
    .col_in_597              ( col_in_597    ),
    .col_in_598              ( col_in_598    ),
    .col_in_599              ( col_in_599    ),
    .col_in_600              ( col_in_600    ),
    .col_in_601              ( col_in_601    ),
    .col_in_602              ( col_in_602    ),
    .col_in_603              ( col_in_603    ),
    .col_in_604              ( col_in_604    ),
    .col_in_605              ( col_in_605    ),
    .col_in_606              ( col_in_606    ),
    .col_in_607              ( col_in_607    ),
    .col_in_608              ( col_in_608    ),
    .col_in_609              ( col_in_609    ),
    .col_in_610              ( col_in_610    ),
    .col_in_611              ( col_in_611    ),
    .col_in_612              ( col_in_612    ),
    .col_in_613              ( col_in_613    ),
    .col_in_614              ( col_in_614    ),
    .col_in_615              ( col_in_615    ),
    .col_in_616              ( col_in_616    ),
    .col_in_617              ( col_in_617    ),
    .col_in_618              ( col_in_618    ),
    .col_in_619              ( col_in_619    ),
    .col_in_620              ( col_in_620    ),
    .col_in_621              ( col_in_621    ),
    .col_in_622              ( col_in_622    ),
    .col_in_623              ( col_in_623    ),
    .col_in_624              ( col_in_624    ),
    .col_in_625              ( col_in_625    ),
    .col_in_626              ( col_in_626    ),
    .col_in_627              ( col_in_627    ),
    .col_in_628              ( col_in_628    ),
    .col_in_629              ( col_in_629    ),
    .col_in_630              ( col_in_630    ),
    .col_in_631              ( col_in_631    ),
    .col_in_632              ( col_in_632    ),
    .col_in_633              ( col_in_633    ),
    .col_in_634              ( col_in_634    ),
    .col_in_635              ( col_in_635    ),
    .col_in_636              ( col_in_636    ),
    .col_in_637              ( col_in_637    ),
    .col_in_638              ( col_in_638    ),
    .col_in_639              ( col_in_639    ),
    .col_in_640              ( col_in_640    ),
    .col_in_641              ( col_in_641    ),
    .col_in_642              ( col_in_642    ),
    .col_in_643              ( col_in_643    ),
    .col_in_644              ( col_in_644    ),
    .col_in_645              ( col_in_645    ),
    .col_in_646              ( col_in_646    ),
    .col_in_647              ( col_in_647    ),
    .col_in_648              ( col_in_648    ),
    .col_in_649              ( col_in_649    ),
    .col_in_650              ( col_in_650    ),
    .col_in_651              ( col_in_651    ),
    .col_in_652              ( col_in_652    ),
    .col_in_653              ( col_in_653    ),
    .col_in_654              ( col_in_654    ),
    .col_in_655              ( col_in_655    ),
    .col_in_656              ( col_in_656    ),
    .col_in_657              ( col_in_657    ),
    .col_in_658              ( col_in_658    ),
    .col_in_659              ( col_in_659    ),
    .col_in_660              ( col_in_660    ),
    .col_in_661              ( col_in_661    ),
    .col_in_662              ( col_in_662    ),
    .col_in_663              ( col_in_663    ),
    .col_in_664              ( col_in_664    ),
    .col_in_665              ( col_in_665    ),
    .col_in_666              ( col_in_666    ),
    .col_in_667              ( col_in_667    ),
    .col_in_668              ( col_in_668    ),
    .col_in_669              ( col_in_669    ),
    .col_in_670              ( col_in_670    ),
    .col_in_671              ( col_in_671    ),
    .col_in_672              ( col_in_672    ),
    .col_in_673              ( col_in_673    ),
    .col_in_674              ( col_in_674    ),
    .col_in_675              ( col_in_675    ),
    .col_in_676              ( col_in_676    ),
    .col_in_677              ( col_in_677    ),
    .col_in_678              ( col_in_678    ),
    .col_in_679              ( col_in_679    ),
    .col_in_680              ( col_in_680    ),
    .col_in_681              ( col_in_681    ),
    .col_in_682              ( col_in_682    ),
    .col_in_683              ( col_in_683    ),
    .col_in_684              ( col_in_684    ),
    .col_in_685              ( col_in_685    ),
    .col_in_686              ( col_in_686    ),
    .col_in_687              ( col_in_687    ),
    .col_in_688              ( col_in_688    ),
    .col_in_689              ( col_in_689    ),
    .col_in_690              ( col_in_690    ),
    .col_in_691              ( col_in_691    ),
    .col_in_692              ( col_in_692    ),
    .col_in_693              ( col_in_693    ),
    .col_in_694              ( col_in_694    ),
    .col_in_695              ( col_in_695    ),
    .col_in_696              ( col_in_696    ),
    .col_in_697              ( col_in_697    ),
    .col_in_698              ( col_in_698    ),
    .col_in_699              ( col_in_699    ),
    .col_in_700              ( col_in_700    ),
    .col_in_701              ( col_in_701    ),
    .col_in_702              ( col_in_702    ),
    .col_in_703              ( col_in_703    ),
    .col_in_704              ( col_in_704    ),
    .col_in_705              ( col_in_705    ),
    .col_in_706              ( col_in_706    ),
    .col_in_707              ( col_in_707    ),
    .col_in_708              ( col_in_708    ),
    .col_in_709              ( col_in_709    ),
    .col_in_710              ( col_in_710    ),
    .col_in_711              ( col_in_711    ),
    .col_in_712              ( col_in_712    ),
    .col_in_713              ( col_in_713    ),
    .col_in_714              ( col_in_714    ),
    .col_in_715              ( col_in_715    ),
    .col_in_716              ( col_in_716    ),
    .col_in_717              ( col_in_717    ),
    .col_in_718              ( col_in_718    ),
    .col_in_719              ( col_in_719    ),
    .col_in_720              ( col_in_720    ),
    .col_in_721              ( col_in_721    ),
    .col_in_722              ( col_in_722    ),
    .col_in_723              ( col_in_723    ),
    .col_in_724              ( col_in_724    ),
    .col_in_725              ( col_in_725    ),
    .col_in_726              ( col_in_726    ),
    .col_in_727              ( col_in_727    ),
    .col_in_728              ( col_in_728    ),
    .col_in_729              ( col_in_729    ),
    .col_in_730              ( col_in_730    ),
    .col_in_731              ( col_in_731    ),
    .col_in_732              ( col_in_732    ),
    .col_in_733              ( col_in_733    ),
    .col_in_734              ( col_in_734    ),
    .col_in_735              ( col_in_735    ),
    .col_in_736              ( col_in_736    ),
    .col_in_737              ( col_in_737    ),
    .col_in_738              ( col_in_738    ),
    .col_in_739              ( col_in_739    ),
    .col_in_740              ( col_in_740    ),
    .col_in_741              ( col_in_741    ),
    .col_in_742              ( col_in_742    ),
    .col_in_743              ( col_in_743    ),
    .col_in_744              ( col_in_744    ),
    .col_in_745              ( col_in_745    ),
    .col_in_746              ( col_in_746    ),
    .col_in_747              ( col_in_747    ),
    .col_in_748              ( col_in_748    ),
    .col_in_749              ( col_in_749    ),
    .col_in_750              ( col_in_750    ),
    .col_in_751              ( col_in_751    ),
    .col_in_752              ( col_in_752    ),
    .col_in_753              ( col_in_753    ),
    .col_in_754              ( col_in_754    ),
    .col_in_755              ( col_in_755    ),
    .col_in_756              ( col_in_756    ),
    .col_in_757              ( col_in_757    ),
    .col_in_758              ( col_in_758    ),
    .col_in_759              ( col_in_759    ),
    .col_in_760              ( col_in_760    ),
    .col_in_761              ( col_in_761    ),
    .col_in_762              ( col_in_762    ),
    .col_in_763              ( col_in_763    ),
    .col_in_764              ( col_in_764    ),
    .col_in_765              ( col_in_765    ),
    .col_in_766              ( col_in_766    ),
    .col_in_767              ( col_in_767    ),
    .col_in_768              ( col_in_768    ),
    .col_in_769              ( col_in_769    ),
    .col_in_770              ( col_in_770    ),
    .col_in_771              ( col_in_771    ),
    .col_in_772              ( col_in_772    ),
    .col_in_773              ( col_in_773    ),
    .col_in_774              ( col_in_774    ),
    .col_in_775              ( col_in_775    ),
    .col_in_776              ( col_in_776    ),
    .col_in_777              ( col_in_777    ),
    .col_in_778              ( col_in_778    ),
    .col_in_779              ( col_in_779    ),
    .col_in_780              ( col_in_780    ),
    .col_in_781              ( col_in_781    ),
    .col_in_782              ( col_in_782    ),
    .col_in_783              ( col_in_783    ),
    .col_in_784              ( col_in_784    ),
    .col_in_785              ( col_in_785    ),
    .col_in_786              ( col_in_786    ),
    .col_in_787              ( col_in_787    ),
    .col_in_788              ( col_in_788    ),
    .col_in_789              ( col_in_789    ),
    .col_in_790              ( col_in_790    ),
    .col_in_791              ( col_in_791    ),
    .col_in_792              ( col_in_792    ),
    .col_in_793              ( col_in_793    ),
    .col_in_794              ( col_in_794    ),
    .col_in_795              ( col_in_795    ),
    .col_in_796              ( col_in_796    ),
    .col_in_797              ( col_in_797    ),
    .col_in_798              ( col_in_798    ),
    .col_in_799              ( col_in_799    ),
    .col_in_800              ( col_in_800    ),
    .col_in_801              ( col_in_801    ),
    .col_in_802              ( col_in_802    ),
    .col_in_803              ( col_in_803    ),
    .col_in_804              ( col_in_804    ),
    .col_in_805              ( col_in_805    ),
    .col_in_806              ( col_in_806    ),
    .col_in_807              ( col_in_807    ),
    .col_in_808              ( col_in_808    ),
    .col_in_809              ( col_in_809    ),
    .col_in_810              ( col_in_810    ),
    .col_in_811              ( col_in_811    ),
    .col_in_812              ( col_in_812    ),
    .col_in_813              ( col_in_813    ),
    .col_in_814              ( col_in_814    ),
    .col_in_815              ( col_in_815    ),
    .col_in_816              ( col_in_816    ),
    .col_in_817              ( col_in_817    ),
    .col_in_818              ( col_in_818    ),
    .col_in_819              ( col_in_819    ),
    .col_in_820              ( col_in_820    ),
    .col_in_821              ( col_in_821    ),
    .col_in_822              ( col_in_822    ),
    .col_in_823              ( col_in_823    ),
    .col_in_824              ( col_in_824    ),
    .col_in_825              ( col_in_825    ),
    .col_in_826              ( col_in_826    ),
    .col_in_827              ( col_in_827    ),
    .col_in_828              ( col_in_828    ),
    .col_in_829              ( col_in_829    ),
    .col_in_830              ( col_in_830    ),
    .col_in_831              ( col_in_831    ),
    .col_in_832              ( col_in_832    ),
    .col_in_833              ( col_in_833    ),
    .col_in_834              ( col_in_834    ),
    .col_in_835              ( col_in_835    ),
    .col_in_836              ( col_in_836    ),
    .col_in_837              ( col_in_837    ),
    .col_in_838              ( col_in_838    ),
    .col_in_839              ( col_in_839    ),
    .col_in_840              ( col_in_840    ),
    .col_in_841              ( col_in_841    ),
    .col_in_842              ( col_in_842    ),
    .col_in_843              ( col_in_843    ),
    .col_in_844              ( col_in_844    ),
    .col_in_845              ( col_in_845    ),
    .col_in_846              ( col_in_846    ),
    .col_in_847              ( col_in_847    ),
    .col_in_848              ( col_in_848    ),
    .col_in_849              ( col_in_849    ),
    .col_in_850              ( col_in_850    ),
    .col_in_851              ( col_in_851    ),
    .col_in_852              ( col_in_852    ),
    .col_in_853              ( col_in_853    ),
    .col_in_854              ( col_in_854    ),
    .col_in_855              ( col_in_855    ),
    .col_in_856              ( col_in_856    ),
    .col_in_857              ( col_in_857    ),
    .col_in_858              ( col_in_858    ),
    .col_in_859              ( col_in_859    ),
    .col_in_860              ( col_in_860    ),
    .col_in_861              ( col_in_861    ),
    .col_in_862              ( col_in_862    ),
    .col_in_863              ( col_in_863    ),
    .col_in_864              ( col_in_864    ),
    .col_in_865              ( col_in_865    ),
    .col_in_866              ( col_in_866    ),
    .col_in_867              ( col_in_867    ),
    .col_in_868              ( col_in_868    ),
    .col_in_869              ( col_in_869    ),
    .col_in_870              ( col_in_870    ),
    .col_in_871              ( col_in_871    ),
    .col_in_872              ( col_in_872    ),
    .col_in_873              ( col_in_873    ),
    .col_in_874              ( col_in_874    ),
    .col_in_875              ( col_in_875    ),
    .col_in_876              ( col_in_876    ),
    .col_in_877              ( col_in_877    ),
    .col_in_878              ( col_in_878    ),
    .col_in_879              ( col_in_879    ),
    .col_in_880              ( col_in_880    ),
    .col_in_881              ( col_in_881    ),
    .col_in_882              ( col_in_882    ),
    .col_in_883              ( col_in_883    ),
    .col_in_884              ( col_in_884    ),
    .col_in_885              ( col_in_885    ),
    .col_in_886              ( col_in_886    ),
    .col_in_887              ( col_in_887    ),
    .col_in_888              ( col_in_888    ),
    .col_in_889              ( col_in_889    ),
    .col_in_890              ( col_in_890    ),
    .col_in_891              ( col_in_891    ),
    .col_in_892              ( col_in_892    ),
    .col_in_893              ( col_in_893    ),
    .col_in_894              ( col_in_894    ),
    .col_in_895              ( col_in_895    ),
    .col_in_896              ( col_in_896    ),
    .col_in_897              ( col_in_897    ),
    .col_in_898              ( col_in_898    ),
    .col_in_899              ( col_in_899    ),
    .col_in_900              ( col_in_900    ),
    .col_in_901              ( col_in_901    ),
    .col_in_902              ( col_in_902    ),
    .col_in_903              ( col_in_903    ),
    .col_in_904              ( col_in_904    ),
    .col_in_905              ( col_in_905    ),
    .col_in_906              ( col_in_906    ),
    .col_in_907              ( col_in_907    ),
    .col_in_908              ( col_in_908    ),
    .col_in_909              ( col_in_909    ),
    .col_in_910              ( col_in_910    ),
    .col_in_911              ( col_in_911    ),
    .col_in_912              ( col_in_912    ),
    .col_in_913              ( col_in_913    ),
    .col_in_914              ( col_in_914    ),
    .col_in_915              ( col_in_915    ),
    .col_in_916              ( col_in_916    ),
    .col_in_917              ( col_in_917    ),
    .col_in_918              ( col_in_918    ),
    .col_in_919              ( col_in_919    ),
    .col_in_920              ( col_in_920    ),
    .col_in_921              ( col_in_921    ),
    .col_in_922              ( col_in_922    ),
    .col_in_923              ( col_in_923    ),
    .col_in_924              ( col_in_924    ),
    .col_in_925              ( col_in_925    ),
    .col_in_926              ( col_in_926    ),
    .col_in_927              ( col_in_927    ),
    .col_in_928              ( col_in_928    ),
    .col_in_929              ( col_in_929    ),
    .col_in_930              ( col_in_930    ),
    .col_in_931              ( col_in_931    ),
    .col_in_932              ( col_in_932    ),
    .col_in_933              ( col_in_933    ),
    .col_in_934              ( col_in_934    ),
    .col_in_935              ( col_in_935    ),
    .col_in_936              ( col_in_936    ),
    .col_in_937              ( col_in_937    ),
    .col_in_938              ( col_in_938    ),
    .col_in_939              ( col_in_939    ),
    .col_in_940              ( col_in_940    ),
    .col_in_941              ( col_in_941    ),
    .col_in_942              ( col_in_942    ),
    .col_in_943              ( col_in_943    ),
    .col_in_944              ( col_in_944    ),
    .col_in_945              ( col_in_945    ),
    .col_in_946              ( col_in_946    ),
    .col_in_947              ( col_in_947    ),
    .col_in_948              ( col_in_948    ),
    .col_in_949              ( col_in_949    ),
    .col_in_950              ( col_in_950    ),
    .col_in_951              ( col_in_951    ),
    .col_in_952              ( col_in_952    ),
    .col_in_953              ( col_in_953    ),
    .col_in_954              ( col_in_954    ),
    .col_in_955              ( col_in_955    ),
    .col_in_956              ( col_in_956    ),
    .col_in_957              ( col_in_957    ),
    .col_in_958              ( col_in_958    ),
    .col_in_959              ( col_in_959    ),
    .col_in_960              ( col_in_960    ),
    .col_in_961              ( col_in_961    ),
    .col_in_962              ( col_in_962    ),
    .col_in_963              ( col_in_963    ),
    .col_in_964              ( col_in_964    ),
    .col_in_965              ( col_in_965    ),
    .col_in_966              ( col_in_966    ),
    .col_in_967              ( col_in_967    ),
    .col_in_968              ( col_in_968    ),
    .col_in_969              ( col_in_969    ),
    .col_in_970              ( col_in_970    ),
    .col_in_971              ( col_in_971    ),
    .col_in_972              ( col_in_972    ),
    .col_in_973              ( col_in_973    ),
    .col_in_974              ( col_in_974    ),
    .col_in_975              ( col_in_975    ),
    .col_in_976              ( col_in_976    ),
    .col_in_977              ( col_in_977    ),
    .col_in_978              ( col_in_978    ),
    .col_in_979              ( col_in_979    ),
    .col_in_980              ( col_in_980    ),
    .col_in_981              ( col_in_981    ),
    .col_in_982              ( col_in_982    ),
    .col_in_983              ( col_in_983    ),
    .col_in_984              ( col_in_984    ),
    .col_in_985              ( col_in_985    ),
    .col_in_986              ( col_in_986    ),
    .col_in_987              ( col_in_987    ),
    .col_in_988              ( col_in_988    ),
    .col_in_989              ( col_in_989    ),
    .col_in_990              ( col_in_990    ),
    .col_in_991              ( col_in_991    ),
    .col_in_992              ( col_in_992    ),
    .col_in_993              ( col_in_993    ),
    .col_in_994              ( col_in_994    ),
    .col_in_995              ( col_in_995    ),
    .col_in_996              ( col_in_996    ),
    .col_in_997              ( col_in_997    ),
    .col_in_998              ( col_in_998    ),
    .col_in_999              ( col_in_999    ),
    .col_in_1000             ( col_in_1000   ),
    .col_in_1001             ( col_in_1001   ),
    .col_in_1002             ( col_in_1002   ),
    .col_in_1003             ( col_in_1003   ),
    .col_in_1004             ( col_in_1004   ),
    .col_in_1005             ( col_in_1005   ),
    .col_in_1006             ( col_in_1006   ),
    .col_in_1007             ( col_in_1007   ),
    .col_in_1008             ( col_in_1008   ),
    .col_in_1009             ( col_in_1009   ),
    .col_in_1010             ( col_in_1010   ),
    .col_in_1011             ( col_in_1011   ),
    .col_in_1012             ( col_in_1012   ),
    .col_in_1013             ( col_in_1013   ),
    .col_in_1014             ( col_in_1014   ),
    .col_in_1015             ( col_in_1015   ),
    .col_in_1016             ( col_in_1016   ),
    .col_in_1017             ( col_in_1017   ),
    .col_in_1018             ( col_in_1018   ),
    .col_in_1019             ( col_in_1019   ),
    .col_in_1020             ( col_in_1020   ),
    .col_in_1021             ( col_in_1021   ),
    .col_in_1022             ( col_in_1022   ),
    .col_in_1023             ( col_in_1023   ),

    .row_out_0               ( compressor_array_512_out0     ),
    .row_out_1               ( compressor_array_512_out1     )
);








// xpb_18 Inputs
wire   [8:0]  u1_data_in0;
wire   [8:0]  u1_data_in1;

// xpb_18 Outputs
wire  [1023:0]  u1_data_out_0;
wire  [1023:0]  u1_data_out_1;
wire  [1023:0]  u1_data_out_2;
wire  [1023:0]  u1_data_out_3;

assign u1_data_in0 = compressor_array_512_out0[1032:1024];
assign u1_data_in1 = compressor_array_512_out1[1032:1024];

xpb_18  u1_xpb_18 (
    .data_in0                ( u1_data_in0     ),
    .data_in1                ( u1_data_in1     ),

    .data_out_0              ( u1_data_out_0   ),
    .data_out_1              ( u1_data_out_1   ),
    .data_out_2              ( u1_data_out_2   ),
    .data_out_3              ( u1_data_out_3   )
);



// compressor_array_6_2_1024_row Inputs
wire   [1023:0]  u2_row_in_0;
wire   [1023:0]  u2_row_in_1;
wire   [1023:0]  u2_row_in_2;
wire   [1023:0]  u2_row_in_3;
wire   [1023:0]  u2_row_in_4;
wire   [1023:0]  u2_row_in_5;

// compressor_array_6_2_1024_row Outputs
wire  [1026:0]  u2_row_out_0;
wire  [1026:0]  u2_row_out_1;


assign u2_row_in_0 = u1_data_out_0;
assign u2_row_in_1 = u1_data_out_1;
assign u2_row_in_2 = u1_data_out_2;
assign u2_row_in_3 = u1_data_out_3;
assign u2_row_in_4 = compressor_array_512_out0[1023:0];
assign u2_row_in_5 = compressor_array_512_out1[1023:0];

compressor_array_6_2_1024_row  u2_compressor_array_6_2_1024_row (
    .row_in_0                ( u2_row_in_0    ),
    .row_in_1                ( u2_row_in_1    ),
    .row_in_2                ( u2_row_in_2    ),
    .row_in_3                ( u2_row_in_3    ),
    .row_in_4                ( u2_row_in_4    ),
    .row_in_5                ( u2_row_in_5    ),

    .row_out_0               ( u2_row_out_0   ),
    .row_out_1               ( u2_row_out_1   )
);






// xpb_6_0 Inputs
wire   [3:1]  u3_data_in0;
wire   [3:1]  u3_data_in1;

// xpb_6_0 Outputs
wire  [1024:1]  u3_data_out;

assign u3_data_in0 = u2_row_out_0[1026:1024];
assign u3_data_in1 = u2_row_out_1[1026:1024];


xpb_6_0  u3_xpb_6_0 (
    .data_in0                ( u3_data_in0   ),
    .data_in1                ( u3_data_in1   ),

    .data_out                ( u3_data_out   )
);








// compressor_array_3_2_1024 Inputs
wire   [1023:0]  u4_row_in_0;
wire   [1023:0]  u4_row_in_1;
wire   [1023:0]  u4_row_in_2;

// compressor_array_3_2_1024 Outputs
wire  [1024:0]  u4_row_out_0;
wire  [1024:0]  u4_row_out_1;


assign u4_row_in_0 = u2_row_out_0[1023:0];
assign u4_row_in_1 = u2_row_out_1[1023:0];
assign u4_row_in_2 = u3_data_out;


compressor_array_3_2_1024_row  u4_compressor_array_3_2_1024_row (
    .row_in_0                ( u4_row_in_0    ),
    .row_in_1                ( u4_row_in_1    ),
    .row_in_2                ( u4_row_in_2    ),

    .row_out_0               ( u4_row_out_0   ),
    .row_out_1               ( u4_row_out_1   )
);


assign data_out_0 = u4_row_out_0;
assign data_out_1 = u4_row_out_1;



endmodule
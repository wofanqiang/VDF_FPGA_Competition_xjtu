module xpb_5_530
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h17f946a51904a256b82e5937d3db4734d76f64fa056b93d3ed4ba1db2dcfa8059a3cbd52c9d5bc4f98a2a74b34395d656916b3d228f404d052cb477252f62bd95b1c8ae2b6a483f9f2f7d78578e450ab82c1ddf869519466e60654d583d0a19aa6347de395c666e8df3d85685be324a0225abe2286acff57456f904efcd914cc;
    5'b00010 : xpb = 1024'h2ff28d4a320944ad705cb26fa7b68e69aedec9f40ad727a7da9743b65b9f500b34797aa593ab789f31454e966872bacad22d67a451e809a0a5968ee4a5ec57b2b63915c56d4907f3e5efaf0af1c8a1570583bbf0d2a328cdcc0ca9ab07a143354c68fbc72b8ccdd1be7b0ad0b7c6494044b57c450d59feae8adf209df9b22998;
    5'b00011 : xpb = 1024'h47ebd3ef4b0de704288b0ba77b91d59e864e2eee1042bb7bc7e2e591896ef810ceb637f85d8134eec9e7f5e19cac18303b441b767adc0e70f861d656f8e2838c1155a0a823ed8bedd8e786906aacf202884599e93bf4bd34b212fe808b71e4cff29d79aac15334ba9db8903913a96de067103a679406fe05d04eb0ecf68b3e64;
    5'b00100 : xpb = 1024'h5fe51a946412895ae0b964df4f6d1cd35dbd93e815ae4f4fb52e876cb73ea01668f2f54b2756f13e628a9d2cd0e57595a45acf48a3d013414b2d1dc94bd8af656c722b8ada920fe7cbdf5e15e39142ae0b0777e1a546519b981953560f42866a98d1f78e57199ba37cf615a16f8c9280896af88a1ab3fd5d15be413bf3645330;
    5'b00101 : xpb = 1024'h77de61397d172bb198e7be1723486408352cf8e21b19e323a27a2947e50e481c032fb29df12cad8dfb2d4478051ed2fb0d71831accc418119df8653b9ecedb3ec78eb66d913693e1bed7359b5c7593598dc955da0e97e6027e1fa82b931328053f067571ece0028c5c339b09cb6fb720abc5b6aca160fcb45b2dd18af03d67fc;
    5'b00110 : xpb = 1024'h8fd7a7de961bce085116174ef723ab3d0c9c5ddc208576f78fc5cb2312ddf0219d6c6ff0bb0269dd93cfebc339583060768836ecf5b81ce1f0c3acadf1c5071822ab415047db17dbb1cf0d20d559e405108b33d277e97a696425fd0116e3c99fe53af35582a669753b7120722752dbc0ce2074cf280dfc0ba09d61d9ed167cc8;
    5'b00111 : xpb = 1024'ha7d0ee83af20705f09447086cafef271e40bc2d625f10acb7d116cfe40ad982737a92d4384d8262d2c72930e6d918dc5df9eeabf1eac21b2438ef42044bb32f17dc7cc32fe7f9bd5a4c6e4a64e3e34b0934d11cae13b0ed04a2c51d69ab46b3a8b6f7139186cd05e1aaea5da83360060f07b32f1aebafb62e60cf228e9ef9194;
    5'b01000 : xpb = 1024'hf1cefd30636ddecf66d51e78e7ff2554a05249f55e4fe27ec805583bb7a9324ce9d6d1d848763ee25b6fb12be6cda60e49b76ab24ed5636e5bafc345cdeea19649522670593228a8524b9892e46c12b2209f62abe0676267aa614b1645a6a43029c5cf2fd6a3eb9732c4463e748fed7c3fc1231e51c9d89e50d07735de63ff5;
    5'b01001 : xpb = 1024'h271636781f3b8043ae9bab1f625b398a217489995b5091fbd9cbf75ee94a3b2a68da2a704e5d203dbe59a25df2a637c64db22a7d4de15b07388643a6afd515f2bfb1ad49bc37a684781c910ea72b11d6a4cbd42327580a8d60ac6986e82b0bdda8d0dad69330a5a25269c9cc432c2377e656d0546bc99ce12a7c97c25abf54c1;
    5'b01010 : xpb = 1024'h3f0f7d1d3840229a66ca0457363680bef8e3ee9360bc25cfc717993a1719e3300316e7c31832dc8d56fc49a926df952bb6c8de4f76d55fd78b518b1902cb41cc1ace382c72dc2a7e6b146894200f6282278db21b90a99ef446b2be5c6bfbad784f0558ba28f70c8b31a74f349f0f481808b18e76f2769c386fec28115798698d;
    5'b01011 : xpb = 1024'h5708c3c25144c4f11ef85d8f0a11c7f3d053538d6627b9a3b4633b1544e98b359d53a515e20898dcef9ef0f45b18f2911fdf92219fc964a7de1cd28b55c16da575eac30f2980ae785e0c401998f3b32daa4f9013f9fb335b2cb91331efcc4f12f539d69dbebd737410e4d49cfaf26cb82b0c4c9979239b8fb55bb86054717e59;
    5'b01100 : xpb = 1024'h6f020a676a496747d726b6c6dded0f28a7c2b8876b934d77a1aedcf072b9333b37906268abde552c8841983f8f524ff688f645f3c8bd697830e819fda8b7997ed1074df1e02532725104179f11d803d92d116e0c634cc7c212bf6807739cf0ad9b6e54815483da5cf0225a0556d591584d670abbffd09ae6facb48af514a9325;
    5'b01101 : xpb = 1024'h86fb510c834e099e8f550ffeb1c8565d7f321d8170fee14b8efa7ecba088db40d1cd1fbb75b4117c20e43f8ac38bad5bf20cf9c5f1b16e4883b3616ffbadc5582c23d8d496c9b66c43fbef248abc5484afd34c04cc9e5c28f8c5bcdcf76d924841a2d264ea4a4145cf5fdf6db2b8b5f86fc1c8de867d9a3e403ad8fe4e23a7f1;
    5'b01110 : xpb = 1024'h9ef497b19c52abf54783693685a39d9256a1827b766a751f7c4620a6ce5883466c09dd0e3f89cdcbb986e6d5f7c50ac15b23ad981aa57318d67ea8e24ea3f131874063b74d6e3a6636f3c6aa03a0a530329529fd35eff08fdecc11b27b3e33e2e7d750488010a82eae9d64d60e9bda98921c87010d2a999585aa694d4afcbcbd;
    5'b01111 : xpb = 1024'h6409900f369198334ac4a9749249d75bc9ae444a65e687bebb5092c49257e4402fe1ce83f390b8cb2cb4eda48a0575c6020398420e6a79d78aab0f666c7a8596e0db9eb5481c11b17519b8ce3a931aac1520e5d12bb57e60f45d48d44e432eb5f043c02650e168a071b035f72aed90f659d6641438c3bbc84aa7e97bef36b1e;
    5'b10000 : xpb = 1024'h1e39dfa60c6dbbd9ecdaa3cf1cffe4aa940a493eabc9fc4fd900ab0776f526499d3ada3b090ec7dc4b6df6257cd9b4c1c936ed5649daac6dcb75f868b9bdd432c92a44ce0b2645150a4973125c8d82564413ec557c0cec4cf54c2962c8b4d4860538b9e5fad47d72e65888c7ce91fdaf87f82463ca393b13ca1a0ee6bbcc7fea;
    5'b10001 : xpb = 1024'h3633264b25725e30a508fd06f0db2bdf6b79ae38b1359023c64c4ce2a4c4ce4f3777978dd2e4842be4109d70b1131227324da12872ceb13e1e413fdb0cb4000c2446cfb0c1cac90efd414a97d571d301c6d5ca4de55e80b3db527e384c857620ab6d37c9909ae45bc5960e302a75224faa52e28650e63a6b0f899f35b8a594b6;
    5'b10010 : xpb = 1024'h4e2c6cf03e7700875d37563ec4b6731442e91332b6a123f7b397eebdd2947654d1b454e09cba407b7cb344bbe54c6f8c9b6454fa9bc2b60e710c874d5faa2be57f635a93786f4d08f039221d4e5623ad4997a8464eb0151ac158d30dd05617bb51a1b5ad26614b44a4d39398865846efccada0a8d79339c254f92f84b57ea982;
    5'b10011 : xpb = 1024'h6625b395577ba2de1565af769891ba491a58782cbc0cb7cba0e3909900641e5a6bf11233668ffccb1555ec071985ccf2047b08ccc4b6badec3d7cebfb2a057beda7fe5762f13d102e330f9a2c73a7458cc59863eb801a981a75f27e35426b955f7d63390bc27b22d84111900e23b6b8fef085ecb5e4039199a68bfd3b257be4e;
    5'b10100 : xpb = 1024'h7e1efa3a70804534cd9408ae6c6d017df1c7dd26c1784b9f8e2f32742e33c660062dcf863065b91aadf893524dbf2a576d91bc9eedaabfaf16a3163205968398359c7058e5b854fcd628d128401ec5044f1b643721533de88d657cb8d7f75af09e0ab17451ee1916634e9e693e1e903011631cede4ed3870dfd85022af30d31a;
    5'b10101 : xpb = 1024'h961840df8984e78b85c261e6404848b2c9374220c6e3df737b7ad44f5c036e65a06a8cd8fa3b756a469b3a9d81f887bcd6a87071169ec47f696e5da4588caf7190b8fb3b9c5cd8f6c920a8adb90315afd1dd422f8aa4d24f736bd18e5bc7fc8b443f2f57e7b47fff428c23d19a01b4d033bddb106b9a37c82547e071ac09e7e6;
    5'b10110 : xpb = 1024'hae118784a28989e23df0bb1e14238fe7a0a6a71acc4f734768c6762a89d3166b3aa74a2bc41131b9df3de1e8b631e5223fbf24433f92c94fbc39a516ab82db4aebd5861e53015cf0bc18803331e7665b549f2027f3f666b659722663df989e25ea73ad3b7d7ae6e821c9a939f5e4d97056189932f247371f6ab770c0a8e2fcb2;
    5'b10111 : xpb = 1024'h155d88d3f99ff7702b199c7ed7a48fcb06a008e3fc4366a3d8355eb004a01168d19b8a05c3c06f7ad88249ed070d31bd44bbb02f45d3fdd45e65ad2ac3a69272d2a2dc525a14e3a59c76551611eff2d5e35c0487d0c1ce0c89ebe93ea93e9d2e61a098f5627855437a4747c359f7d7e72999787328a8d94669b7860b1cd9ab13;
    5'b11000 : xpb = 1024'h2d56cf7912a499c6e347f5b6ab7fd6ffde0f6dde01aefa77c581008b326fb96e6bd847588d962bca7124f1383b468f22add264016ec802a4b130f49d169cbe4c2dbf673510b9679f8f6e2c9b8ad44381661de2803a1362736ff23e142d0f3ec907d516d8f83ebc2c5984cd2bb5dafc874bf43695af55d89daf27165a19b2bfdf;
    5'b11001 : xpb = 1024'h4550161e2ba93c1d9b764eee7f5b1e34b57ed2d8071a8e4bb2cca266603f6174061504ab576be81a09c798836f7fec8816e917d397bc077503fc3c0f6992ea2588dbf217c75deb998266042103b8942ce8dfc078a364f6da55f892e9b0dfe063ae0994bc8e05231538c2529411be21276e4ef4b83602d7f4f496a6a9168bd4ab;
    5'b11010 : xpb = 1024'h5d495cc344adde7453a4a826533665698cee37d20c86221fa01844418e0f0979a051c1fe2141a469a26a3fcea3b949ed7fffcba5c0b00c4556c78381bc8915fee3f87cfa7e026f93755ddba67c9ce4d86ba19e710cb68b413bfee7bf34b081fe543e12a023cb89fe17ffd7fc6da145c790a9b2dabcafd74c3a0636f81364e977;
    5'b11011 : xpb = 1024'h7542a3685db280cb0bd3015e2711ac9e645d9ccc11f1b5f38d63e61cbbdeb17f3a8e7f50eb1760b93b0ce719d7f2a752e9167f77e9a41115a992caf40f7f41d83f1507dd34a6f38d6855b32bf5813583ee637c6976081fa822053c94b8812398fa729083b991f0e6f73d5d64c9846a67b30470fd435cd6a37f75c747103dfe43;
    5'b11100 : xpb = 1024'h8d3bea0d76b72321c4015a95faecf3d33bcd01c6175d49c77aaf87f7e9ae5984d4cb3ca3b4ed1d08d3af8e650c2c04b8522d334a129815e5fc5e126662756db19a3192bfeb4b77875b4d8ab16e65862f71255a61df59b40f080b916a3c51c533a0a70e674f5857cfd67ae2cd25678f07d55f2f1fca09d5fac4e557960d17130f;
    5'b11101 : xpb = 1024'ha53530b28fbbc5787c2fb3cdcec83b08133c66c01cc8dd9b67fb29d3177e018a6f07f9f67ec2d9586c5235b04065621dbb43e71c3b8c1ab64f2959d8b56b998af54e1da2a1effb814e456236e749d6daf3e7385a48ab4875ee11e63fc02266ce46db8c4ae51ebeb8b5b86835814ab3a7f7b9ed4250b6d5520a54e7e509f027db;
    5'b11110 : xpb = 1024'hc813201e6d233066958952e92493aeb7935c8894cbcd0f7d76a1258924afc8805fc39d07e72171965969db49140aeb8c040730841cd4f3af15561eccd8f50b2dc1b73d6a90382362ea33719c752635582a41cba2576afcc1e8ba91a89c865d6be087804ca1c2d140e3606bee55db21ecb3acc82871877790954fd2f7de6d63c;
    5'b11111 : xpb = 1024'h247a78a6ffd6d55d2186ee666624822050a52d83522864cbc4b5b433c01aa48da038f7234847d368fe3944ffc57a0c1e295726da6ac1540b4420a95f20857c8c3737feb95fa80630219b0e9f4036b4010565fab28ec844330491fdf00d990771643cf5e85fe293fced738c274140d6beed958aa50dc576d04ec48d7e7abfeb08;
    endcase
end

endmodule

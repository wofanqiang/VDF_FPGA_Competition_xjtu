module xpb_5_325
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h2bd6ed8bd69639939736aebfc3a7b447c72945431a0a7bd2d85d01a2ab64288e7a20c1422d86437d8a6328f83de4be7a4fe0efb4032060be5e9ffe871e27940091371943fb9ad38cddd7a17eb11540f007d51e42b885c609cbee73b9e2aa62635ff74901a2ab11218b524419a2eeb20234f65d39eb2035c0449daa291c825834;
    5'b00010 : xpb = 1024'h57addb17ad2c73272e6d5d7f874f688f8e528a863414f7a5b0ba034556c8511cf44182845b0c86fb14c651f07bc97cf49fc1df680640c17cbd3ffd0e3c4f2801226e3287f735a719bbaf42fd622a81e00faa3c85710b8c1397dce773c554c4c6bfee92034556224316a4883345dd640469ecba73d6406b80893b54523904b068;
    5'b00011 : xpb = 1024'h8384c8a383c2acbac5a40c3f4af71cd7557bcfc94e1f7378891704e8022c79ab6e6243c68892ca789f297ae8b9ae3b6eefa2cf1c0961223b1bdffb955a76bc01b3a54bcbf2d07aa69986e47c133fc2d0177f5ac82991521d63cb5b2da7ff272a1fe5db04e8013364a1f6cc4ce8cc16069ee317adc160a140cdd8fe7b5587089c;
    5'b00100 : xpb = 1024'haf5bb62f5a58e64e5cdabaff0e9ed11f1ca5150c6829ef4b6174068aad90a239e8830508b6190df6298ca3e0f792f9e93f83bed00c8182f97a7ffa1c789e500244dc650fee6b4e33775e85fac45503c01f54790ae21718272fb9cee78aa9898d7fdd24068aac44862d4910668bbac808d3d974e7ac80d7011276a8a4720960d0;
    5'b00101 : xpb = 1024'h2a855e656f00eb19290bf1e7c1ec3e157258571eacbccaa6bbf44ed7a5f21dc05f5b48d21978d2e514918d925219a7992b4a869decef136c2880b9455bf36f5161c449a53a75247b429c24d6dc8e807f33249db50e16b120461bb0a6b329495eb0ccdade7c8e5d1a31db6da136d953e1b9f5f33f4755af9110a4d7c905a95299;
    5'b00110 : xpb = 1024'h565c4bf1459724acc042a0a78593f25d39819c61c6c746799451507a5156464ed97c0a1446ff16629ef4b68a8ffe66137b2b7651f00f742a8720b7cc7a1b0351f2fb62e9360ff8082073c6558da3c16f3af9bbf7c69c772a120a246095d3abc210c423e01f396e3bbd2db1bad9c805e3eeec50793275e551554281f2222baacd;
    5'b00111 : xpb = 1024'h8233397d1c2d5e4057794f67493ba6a500aae1a4e0d1c24c6cae521cfcba6edd539ccb56748559e02957df82cde3248dcb0c6605f32fd4e8e5c0b6539842975284327c2d31aacb94fe4b67d43eb9025f42ceda3a7f223d33ddf8981a787e0e2570bb6ce1c1e47f5d487ff5d47cb6b7e623e2adb31d961b1199e02c1b3eae0301;
    5'b01000 : xpb = 1024'hae0a2708f2c397d3eeaffe270ce35aecc7d426e7fadc3e1f450b53bfa81e976bcdbd8c98a20b9d5db3bb087b0bc7e3081aed55b9f65035a74460b4dab66a2b53156995712d459f21dc230952efce434f4aa3f87d37a8033da9e70bd45b287088d0b2b5e3648f907ed3d239ee1fa569e858d90aed08b650d1de7dd6445b305b35;
    5'b01001 : xpb = 1024'h2933cf3f076b9c9ebae1350fc030c7e31d8768fa3f6f197a9f8b9c0ca08012f24495d062056b624c9ebff22c664e90b806b41d87d6bdc619f261740399bf4aa232517a06794f7569a760a82f0807c00e5e741d2763a79c36c048ed9383a8305a01a26cbb5671a912d8649728cac3f5c13ef58944a38b2961dcac0568eed04cfe;
    5'b01010 : xpb = 1024'h550abccade01d6325217e3cf83d87c2ae4b0ae3d5979954d77e89daf4be43b80beb691a432f1a5ca29231b24a4334f3256950d3bd9de26d85101728ab7e6dea2c388934a74ea48f6853849adb91d00fe66493b6a1c2d62408c37614d665292bd6199b5bcf91cba3463b6db426db2a7c373ebe67e8eab5f222149af920b52a532;
    5'b01011 : xpb = 1024'h80e1aa56b4980fc5e94e928f47803072abd9f3807384112050459f51f748640f38d752e66077e947b386441ce2180daca675fcefdcfe8796afa17111d60e72a354bfac8e70851c83630feb2c6a3241ee6e1e59acd4b3284a5825d50748fcf520c190febe9bc7cb55ef091f5c10a159c5a8e243b879cb94e265e759bb27d4fd66;
    5'b01100 : xpb = 1024'hacb897e28b2e49598085414f0b27e4ba730338c38d8e8cf328a2a0f4a2ac8c9db2f814288dfe2cc53de96d151ffccc26f656eca3e01ee8550e416f98f43606a3e5f6c5d26c1ff01040e78cab1b4782de75f377ef8d38ee54241448c12ba75784218847c03e72dc777a5b6375b3900bc7ddd8a0f264ebcaa2aa8503e44457559a;
    5'b01101 : xpb = 1024'h27e240189fd64e244cb67837be7551b0c8b67ad5d221684e8322e9419b0e082429d057f1f15df1b428ee56c67a8379d6e21db471c08c78c7bc422ec1d78b25f302deaa67b829c6580c252b873380ff9d89c39c99b938874d3a762a80542717555277fe983054f50b7eedc0b05eae97a0c3f51f49ffc0a332a8b33308d7f74763;
    5'b01110 : xpb = 1024'h53b92da4766c87b7e3ed26f7821d05f88fdfc018ec2be4215b7feae4467230b2a3f119341ee43531b3517fbeb868385131fea425c3acd9861ae22d48f5b2b9f39415c3abb3c499e4e9fccd05e496408d9198badc71be4d5706649e3a36d179b8b26f4799d300062d0a4004ca019d49a2f8eb7c83eae0d8f2ed50dd31f4799f97;
    5'b01111 : xpb = 1024'h7f901b304d02c14b7b23d5b745c4ba405709055c06365ff433dcec86f1d659411e11da764c6a78af3db4a8b6f64cf6cb81df93d9c6cd3a4479822bd013da4df4254cdcefaf5f6d71c7d46e8495ab817d996dd91f2a441360d25311f4197bdc1c1266909b75ab174e959248e3a48bfba52de1d9bdd6010eb331ee875b10fbf7cb;
    5'b10000 : xpb = 1024'hab6708bc2398fadf125a8477096c6e881e324a9f2040dbc70c39ee299d3a81cf98329bb879f0bc2cc817d1af3431b545d1c0838dc9ed9b02d8222a573201e1f4b683f633aafa40fea5ac100346c0c26da142f761e2c9d96a9e4185adfc263e7f725dd99d1856287020e48cfd477aada762d836f7c1214473768c31842d7e4fff;
    5'b10001 : xpb = 1024'h2690b0f23840ffa9de8bbb5fbcb9db7e73e58cb164d3b72266ba3676959bfd560f0adf81dd50811bb31cbb608eb862f5bd874b5baa5b2b758622e98015570143d36bdac8f704174670e9aedf5efa3f2cb5131c0c0ec97263b4a3676d24a5fe50a34d90750a3841042576ea37f299398048f4b54f5bf61d0374ba60a8c11e41c8;
    5'b10010 : xpb = 1024'h52679e7e0ed7393d75c26a1f80618fc63b0ed1f47ede32f53f173819410025e4892ba0c40ad6c4993d7fe458cc9d21700d683b0fad7b8c33e4c2e807337e954464a2f40cf29eead34ec1505e100f801cbce83a4ec74f386d8091db27075060b40344d976ace35225b0c92e519587eb827deb1289471652c3b9580ad1dda099fc;
    5'b10011 : xpb = 1024'h7e3e8c09e56d72d10cf918df4409440e0238173798e8aec8177439bbec644e73034c6206385d0816c7e30d510a81dfea5d492ac3b09becf24362e68e51a62944f5da0d50ee39be602c98f1dcc124c10cc4bd58917fd4fe774c804ee0e9fac317633c22784f8e63473c1b726b38769d84b2e16fc332368883fdf5b4fafa22f230;
    5'b10100 : xpb = 1024'haa157995bc03ac64a42fc79f07b0f855c9615c7ab2f32a9aefd13b5e97c877017d6d234865e34b945246364948669e64ad2a1a77b3bc4db0a202e5156fcdbd4587112694e9d491ed0a70935b723a01fccc9276d4385ac481186ec29acca5257ac3336b79f2397468c76db684db654f86e7d7ccfd1d56be4442935f2416a54a64;
    5'b10101 : xpb = 1024'h253f21cbd0abb12f7060fe87bafe654c1f149e8cf78605f64a5183ab9029f287f4456711c94310833d4b1ffaa2ed4c1498f0e2459429de235003a43e5322dc94a3f90b2a35de6834d5ae32378a737ebbe0629b7e645a5d7a2ed0a459f524e54bf4232251e41b8cfccc0013bf8683db5fcdf44b54b82b96d440c18e48aa453c2d;
    5'b10110 : xpb = 1024'h51160f57a741eac30797ad477ea61993e63de3d0119081c922ae854e3b8e1b166e662853f6c95400c7ae48f2e0d20a8ee8d1d1f9974a3ee1aea3a2c5714a70953530246e31793bc1b385d3b63b88bfabe837b9c11ce02383fabf1813d7cf47af541a6b5386c69e1e575257d929728d6202eaa88ea34bcc94855f3871c6c79461;
    5'b10111 : xpb = 1024'h7cecfce37dd824569ece5c07424dcddbad6729132b9afd9bfb0b86f0e6f243a4e886e996244f977e521171eb1eb6c90938b2c1ad9a6a9fa00d43a14c8f720495c6673db22d140f4e915d7534ec9e009bf00cd803d565e98dc6ad8bcdba79aa12b411b4552971af3fe2a49bf2cc613f6437e105c88e6c0254c9fce29ae349ec95;
    5'b11000 : xpb = 1024'ha8c3ea6f546e5dea36050ac705f5822374906e5645a5796ed368889392566c3362a7aad851d5dafbdc749ae35c9b87838893b1619d8b005e6be39fd3ad999896579e56f628aee2db6f3516b39db3418bf7e1f6468debaf97929bff879d240c761408fd56cc1cc0616df6e00c6f4ff1666cd76302798c38150e9a8cc3ffcc44c9;
    5'b11001 : xpb = 1024'h23ed92a5691662b5023641afb942ef19ca43b0688a3854ca2de8d0e08ab7e7b9d97feea1b5359feac7798494b7223533745a792f7df890d119e45efc90eeb7e574863b8b74b8b9233a72b58fb5ecbe4b0bb21af0b9eb4890a8fde146c5a3cc4744f8b42ebdfed8f572893d471a6e7d3f52f3e15a146110a50cc8bbe8936c3692;
    5'b11010 : xpb = 1024'h4fc480313fac9c48996cf06f7ceaa361916cf5aba442d09d0645d283361c104853a0afe3e2bbe36851dcad8cf506f3adc43b68e38118f18f78845d83af164be605bd54cf70538cb0184a570e6701ff3b1387393372710e9a74ec5500a84e2eaaa4effd3060a9ea16fddb8160bd5d2f4187ea3e93ff81466551666611afee8ec6;
    5'b11011 : xpb = 1024'h7b9b6dbd1642d5dc30a39f2f409257a958963aeebe4d4c6fdea2d425e18038d6cdc17126104226e5dc3fd68532ebb228141c58978439524dd7245c0acd3ddfe696f46e136bee603cf621f88d1817402b1b5c57762af6d4a440dac8ba8af8910e04e746320354fb38892dc57a604be143bce09bcdeaa17c259604103acc70e6fa;
    5'b11100 : xpb = 1024'ha7725b48ecd90f6fc7da4def043a0bf11fbf8031d857c842b6ffd5c88ce4616547e232683dc86a6366a2ff7d70d070a263fd484b8759b30c35c45a91eb6573e7282b8757678933c9d3f99a0bc92c811b233175b8e37c9aae0cc93c746da2f37164de8f33a6000c5a14800994033a9345f1d6f907d5c1b1e5daa1ba63e8f33f2e;
    5'b11101 : xpb = 1024'h229c037f0181143a940b84d7b78778e77572c2441ceaa39e11801e158545dcebbeba7631a1282f5251a7e92ecb571e524fc4101967c7437ee3c519baceba933645136becb3930a119f3738e7e165fdda37019a630f7c33a7232b1e339622b34295ce460b97e224ee191266ceae591f1ed7f3775f70968a75d8cfe9887c9330f7;
    5'b11110 : xpb = 1024'h4e72f10ad8174dce2b4233977b2f2d2f3c9c078736f51f70e9dd1fb830aa057a38db3773ceae72cfdc0b1227093bdccc9fa4ffcd6ae7a43d42651841ece22736d64a8530af2ddd9e7d0eda66927b3eca3ed6b8a5c801f9b0ef1991ed78cd15a5f5c58f0d3a8d360fa464aae85147d1210ce9d4995bb6c0361d6d93b19915892b;
    5'b11111 : xpb = 1024'h7a49de96aead8761c278e2573ed6e17703c54cca50ff9b43c23a215adc0e2e08b2fbf8b5fc34b64d666e3b1f47209b46ef85ef816e0804fba10516c90b09bb3767819e74aac8b12b5ae67be543907fba46abd6e88087bfbabb0805a75b77780955bcd80edd3847312fb6ef01f436832341e031d346d6f5f6620b3ddab597e15f;
    endcase
end

endmodule

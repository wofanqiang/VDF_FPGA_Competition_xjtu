module xpb_5_210
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h2efe2687a3db34bdbaffc194d84e6edb1ce088f1b87459e50649d9de8651ac70bbf1a1bc5c14bc5e1c8579c387ac5e2f18d22f38d28592caff6b33c7a1e4cbfa8e3aabe66629798f6f623978ae1084526ddff4e76e6c2fa03c3089fa35533b39092bf28721b4240d4612259e187e409b20e1e3bfcc76375623bd0531c63ed06c;
    5'b00010 : xpb = 1024'h5dfc4d0f47b6697b75ff8329b09cddb639c111e370e8b3ca0c93b3bd0ca358e177e34378b82978bc390af3870f58bc5e31a45e71a50b2595fed6678f43c997f51c7557cccc52f31edec472f15c2108a4dbbfe9cedcd85f40786113f46aa676721257e50e4368481a8c244b3c30fc813641c3c77f98ec6eac477a0a638c7da0d8;
    5'b00011 : xpb = 1024'h8cfa7396eb919e3930ff44be88eb4c9156a19ad5295d0daf12dd8d9b92f5055233d4e535143e351a55906d4a97051a8d4a768daa7790b860fe419b56e5ae63efaab003b3327c6cae4e26ac6a0a318cf7499fdeb64b448ee0b4919dee9ff9b1ab1b83d795651c6c27d23670da497ac1d162a5ab3f6562a6026b370f9552bc7144;
    5'b00100 : xpb = 1024'hb4b54c8cd7e9e2e20f98e7c50df741b020c20960c59c71c9b4aae24664404baec7e0978a62c72e9d2b7a7c73b5367f1ff2e94fd27637ae04d0d8fc04cc0bb38c49b7aeae914e8f8aaeee3401f664d18c37ada052d2a91703b3595ee1b224a51f5a837f2d60797a79188af996a28dc4334adb01ce18d8028488499c29018db45;
    5'b00101 : xpb = 1024'h3a497b507159d2ebdbf95011292de2f61eeca987c4ce2101a1948802ec95b12ba86fab3502412f47ef3d218ac2ffc6211800c435f9e90dab4c78c387eea5873352d626d14f3e62881a511cb8cd76d16b315aceec9b96c11077661fe85075858afed42a79f7bbbbb4d79ad53782a71cde558f93dcae03b77e6c419ef45657abb1;
    5'b00110 : xpb = 1024'h6947a1d8153507a996f911a6017c51d13bcd32797d427ae6a7de61e172e75d9c64614cf15e55eba60bc29b4e4aac245030d2f36ecc6ea0764be3f74f908a532de110d2b7b567dc1789b356317b8755bd9f3ac3d40a02f0b0b396a9e285c8c0c408001d01196fdfc21dacfad59b255d797671779c7a79eed48ffea4261c967c1d;
    5'b00111 : xpb = 1024'h9845c85fb9103c6751f8d33ad9cac0ac58adbb6b35b6d4cbae283bbff9390a0d2052eeadba6aa80428481511d258827f49a522a79ef433414b4f2b17326f1f286f4b7e9e1b9155a6f9158faa2997da100d1ab8bb786f2050efc733dcbb1bfbfd112c0f883b2403cf63bf2073b3a39e1497535b5c46f0262ab3bba957e2d54c89;
    5'b01000 : xpb = 1024'h1696a9919afd3c5c41f31cf8a1bee8360418412c18b38e3936955c48cc880975d8fc12f14c58e5d3a56f4f8e76a6cfe3fe5d29fa4ec6f5c09a1b1f80998176718936f5d5d229d1f155ddc6803ecc9a3186f5b40a5a5522e0766b2bdc364494a3eb506fe5ac0f2f4f23115f32d451b886695b6039c31b0050910933852031b68a;
    5'b01001 : xpb = 1024'h4594d0193ed87119fcf2de8d7a0d571120f8ca1dd127e81e3cdf362752d9b5e694edb4ada86da231c1f4c951fe532e13172f5933214c888b998653483b66426c1771a1bc38534b80c53ffff8ecdd1e83f4d5a8f1c8c15280b29bb5d66b97cfdcf47c626ccdc3535c692384d0eccff9218a3d43f98f9137a6b4c638b6e67086f6;
    5'b01010 : xpb = 1024'h7492f6a0e2b3a5d7b7f2a022525bc5ec3dd9530f899c420343291005d92b625750df566a04825e8fde7a431585ff8c423001886bf3d21b5698f1870fdd4b0e66a5ac4da29e7cc51034a239719aeda2d662b59dd9372d8220eecc3fd0a0eb0b15fda854f3ef777769af35aa6f054e39bcab1f27b95c076efcd8833de8acaf5762;
    5'b01011 : xpb = 1024'ha3911d28868eda9572f261b72aaa34c75ab9dc0142109be84972e9e45f7d0ec80cd0f82660971aedfaffbcd90dabea7148d3b7a4c657ae21985cbad77f2fda6133e6f98904a63e9fa40472ea48fe2728d09592c0a599b1c12afcc9cad63e464f06d4477b112b9b76f547d00d1dcc7a57cc010b79287da652fc40431a72ee27ce;
    5'b01100 : xpb = 1024'h21e1fe5a687bda8a62ecab74f29e5c51062461c2250d5555d1e00a6d32cc0e30c57a1c69f28558bd7826f755b1fa37d5fd8bbef7762a70a0e728af40e64231aa4dd270c0bb3ebaea00cca9c05e32e74a4a708e0f877fb450b1a0c1ca5166def5e0f8a7d88216c6f6b49a0ecc3e7a94c99e091056a4a88078d98dcd47b04a91cf;
    5'b01101 : xpb = 1024'h50e024e20c570f481dec6d09caeccb2c2304eab3dd81af3ad829e44bb91dbaa1816bbe264e9a151b94ac711939a69605165dee3048b0036be693e3088826fda4dc0d1ca721683479702ee3390c436b9cb85082f6f5ebe3f0edd14bc486ba1a2eea249a5fa3caeb03faac346a56f8d564beeaf416711eb7cefd4ad2797689623b;
    5'b01110 : xpb = 1024'h7fde4b69b0324405d8ec2e9ea33b3a073fe573a595f6091fde73be2a3f6f67123d5d5fe2aaaed179b131eadcc152f4342f301d691b359636e5ff16d02a0bc99f6a47c88d8791ae08df911cb1ba53efef263077de645813912a01d5bebc0d5567f3508ce6c57f0f1140be5a086f7715ffdfccd7d63d94ef252107d7ab3cc832a7;
    5'b01111 : xpb = 1024'haedc71f1540d78c393ebf0337b89a8e25cc5fc974e6a6304e4bd9808c5c11382f94f019f06c38dd7cdb764a048ff526348024ca1edbb2901e56a4a97cbf09599f8827473edbb27984ef3562a6864744194106cc5d2c4433166325fb8f16090a0fc7c7f6de733331e86d07fa687f5569b00aebb960a0b267b44c4dcdd03070313;
    5'b10000 : xpb = 1024'h2d2d532335fa78b883e639f1437dd06c0830825831671c726d2ab891991012ebb1f825e298b1cba74ade9f1ced4d9fc7fcba53f49d8deb8134363f013302ece3126debaba453a3e2abbb8d007d9934630deb6814b4aa45c0ecd657b86c892947d6a0dfcb581e5e9e4622be65a8a3710cd2b6c073863600a12212670a40636d14;
    5'b10001 : xpb = 1024'h5c2b79aad9d5ad763ee5fb861bcc3f4725110b49e9db7657737492701f61bf5c6de9c79ef4c68805676418e074f9fdf7158c832d70137e4c33a172c8d4e7b8dda0a897920a7d1d721b1dc6792ba9b8b57bcb5cfc231675612906e1b2a1dc6480dfccd25279d282ab8c34e403c121b1a7f398a43352ac37f745cf6c3c06a23d80;
    5'b10010 : xpb = 1024'h8b29a0327db0e233f9e5bd1af41aae2241f1943ba24fd03c79be6c4ea5b36bcd29db695b50db446383e992a3fca65c262e5eb26642991117330ca69076cc84d82ee3437870a697018a7ffff1d9ba3d07e9ab51e39182a50165376bacd72f9fb9e8f8c4d99b86a6b8d24709a1d99ff243147a87f31f226f4d698c716dcce10dec;
    5'b10011 : xpb = 1024'h97a81645f9de228e9e006d8bc0ed5abed5c19fc854c89aa022b8cd779026b35e2848d9ee2c982330110cd20a0f4a98ae316b9b8f26bd39681d89af9dddedc2148cebab0273f134be74836c7eeeefd2963864d327368a790ebdb63ac52583860c31d25370c71d23891994860fa4e0cb4e6828cd09b4d497346d9fb9b0a3d77ed;
    5'b10100 : xpb = 1024'h3878a7ec037916e6a4dfc86d945d44870a3ca2ee3dc0e38f087566b5ff5417a69e762f5b3ede3e911d9646e428a107b9fbe8e8f1c4f166618143cec17fc3a81bd70966968d688cdb56aa70409cff817bd1664219e1d4d731280beda687ab7399cc4917be2e25f645d7ab6dff12cc4d500764709067c380c96a9700ccd07c4859;
    5'b10101 : xpb = 1024'h6776ce73a7544ba45fdf8a026cabb362271d2bdff6353d740ebf409485a5c4175a67d1179af2faef3a1bc0a7b04d65e914bb182a9776f92c80af028921a874166544127cf392066ac60ca9b94b1005ce3f463701504106d1643c77a0bcfeaed2d5750a454fda1a531dbd939d2b4a8deb284654503439b81f8e5405fe96bb18c5;
    5'b10110 : xpb = 1024'h9674f4fb4b2f80621adf4b9744fa223d43fdb4d1aea9975915091a730bf77088165972d3f707b74d56a13a6b37f9c4182d8d476369fc8bf7801a3650c38d4010f37ebe6359bb7ffa356ee331f9208a20ad262be8bead3671a06d019af251ea0bdea0fccc718e3e6063cfb93b43c8ce864928381000afef75b2110b305cf9e931;
    5'b10111 : xpb = 1024'h14c5d62d2d1c80570ad995550cee49c6ef683a9291a650c69d763afbdf466ff0cf02971788f5f51cd3c874e7dc48117ce2454eb619cf4e76cee62aba2a9f975a0d6a359b1053fc4492371a080e554a4227012737a09339012710f99a6d7a82b2b8c55d29e27969e02321f7fa6476e8f81b303ced7cdac99b8f5e955d9a565332;
    5'b11000 : xpb = 1024'h43c3fcb4d0f7b514c5d956e9e53cb8a20c48c3844a1aaaaba3c014da65981c618af438d3e50ab17af04deeab63f46fabfb177deeec54e141ce515e81cc8463549ba4e181767d75d401995380bc65ce9494e11c1f0eff68a163418394a2cdbdebc1f14fb1042d8ded69341d987cf529933c1220ad495100f1b31b9a8f6095239e;
    5'b11001 : xpb = 1024'h72c2233c74d2e9d280d9187ebd8b277d29294c76028f0490aa09eeb8ebe9c8d246e5da90411f6dd90cd3686eeba0cddb13e9ad27beda740ccdbc92496e692f4f29df8d67dca6ef6370fb8cf96a7652e702c111067d6b98419f720d8ed820f924cb1d423825e1b1faaf46433695736a2e5cf4046d15c73847d6d89fc126d3f40a;
    5'b11010 : xpb = 1024'ha1c049c418ae1e903bd8da1395d996584609d567bb035e75b053c897723b754302d77c4c9d342a372958e232734d2c0a2cbbdc60916006d7cd27c611104dfb49b81a394e42d068f2e05dc6721886d73970a105edebd7c7e1dba297890d74345dd44934bf4795d607f55868d4adf1aac97dd5e82ce23d6f9dfa95a4f2ed12c476;
    5'b11011 : xpb = 1024'h20112af5fa9b1e852bd323d15dcdbde1f1745b289e0017e338c0e920458a74abbb80a0902f226806a6801caf179b796ee173e3b34132c9571bf3ba7a77605292d205b085f968e53d3d25fd482dbb975aea7c013ccdbdca7162468f88889ccd04ae6d951cb8810187b4aaa793ce9fc53b4fdded0a5e6849c3d7e32f202a6f2e77;
    5'b11100 : xpb = 1024'h4f0f517d9e765342e6d2e566361c2cbd0e54e41a567471c83f0ac2fecbdc211c7772424c8b372464c30596729f47d79dfa4612ec13b85c221b5eee4219451e8d60405c6c5f925eccac8836c0dbcc1bad585bf6243c29fa119e771982bdf0083db79987a3da352594fabccd31e71e05d670bfd0ca2ade8119fba03451f0adfee3;
    5'b11101 : xpb = 1024'h7e0d780542518800a1d2a6fb0e6a9b982b356d0c0ee8cbad45549cdd522dcd8d3363e408e74be0c2df8b103626f435cd13184224e63deeed1aca2209bb29ea87ee7b0852c5bbd85c1bea703989dc9fffc63beb0baa9629b1daa7a37cf3434376c0c57a2afbe949a240cef2cfff9c467191a1b489f754b8701f5d3983b6eccf4f;
    5'b11110 : xpb = 1024'had0b9e8ce62cbcbe5cd2688fe6b90a734815f5fdc75d25924b9e76bbd87f79fdef5585c543609d20fc1089f9aea093fc2bea715db8c381b81a3555d15d0eb6827cb5b4392be551eb8b4ca9b237ed2452341bdff31902595216d82d7728967eafc9f16cb21d9d6daf86e1186e181a870cb2839849c3caefc6431a3eb57d2b9fbb;
    5'b11111 : xpb = 1024'h2b5c7fbec819bcb34cccb24daead31fcf3807bbeaa59deffd40b9744abce7966a7feaa08d54edaf07937c47652eee160e0a278b06896443769014a3ac4210dcb96a12b70e27dce35e814e0884d21e473adf6db41fae85be19d7c2576a3bf1756a415cd0f8e88992f4633572d38c8a17e848b9d273ff5c9ec2067c8e2ba8809bc;
    endcase
end

endmodule

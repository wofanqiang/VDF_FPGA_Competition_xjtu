module xpb_5_115
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h9af3a9ec43d7f289d38af60f1a49d8be5a2664d4c9cfcd76e1ea4fdb57c292d13157eb8f47ca0a1e046f4cc6ab7cb342d415eff874e9092159a757e195a92fb6d231fe872e922eb3b4c857d9c76236e729aad4134c5bfde03cca593bfdb9109ee25d8be946fc1e9e5cb3cc99e01bb7dae1ad169819765a8b2664fc9a491603f0;
    5'b00010 : xpb = 1024'h853a0e82c5c1b04adc10744724396a2b42d6c678be27fa7645f7e660fc82789a5f6759a5c56d95ad69805a46739b55bb4411b80ac71f41f702af7064f07feabc3014c85fad93602256f6ad10f5e8a99d5f50ae8e0c31ceafc408207d41477eab95b385a8dd2f44af32a7b254c867498c74804e4de2a157e6065a7e300949a175;
    5'b00011 : xpb = 1024'h6f80731947ab6e0be495f27f2e28fb982b87281cb2802775aa057ce6a1425e638d76c7bc4311213cce9167c63bb9f833b40d801d19557accabb788e84b56a5c18df792382c949190f9250248246f1c5394f68908cc079f7f4b45e7be84d5ecb849097f6873626ac0089b980fb0b2db3e07538603abcc5540e64fffc5c97d3efa;
    5'b00100 : xpb = 1024'h59c6d7afc9952bcced1b70b738188d05143789c0a6d854750e13136c4602442cbb8635d2c0b4accc33a2754603d89aac2409482f6b8bb3a254bfa16ba62d60c6ebda5c10ab95c2ff9b53577f52f58f09ca9c63838bdd704ed283aeffc8645ac4fc5f7928099590d0de8f7dca98fe6cef9a26bdb974f7529bc645815b89b0dc7f;
    5'b00101 : xpb = 1024'h440d3c464b7ee98df5a0eeef42081e71fce7eb649b3081747220a9f1eac229f5e995a3e93e58385b98b382c5cbf73d2494051041bdc1ec77fdc7b9ef01041bcc49bd25e92a96f46e3d81acb6817c01c000423dfe4bb3411e59c176410bf2c8d1afb572e79fc8b6e1b48363858149fea12cf9f56f3e224ff6a63b02f149e47a04;
    5'b00110 : xpb = 1024'h2e53a0dccd68a74efe266d274bf7afdee5984d088f88ae73d62e40778f820fbf17a511ffbbfbc3eafdc490459415df9d0400d8540ff8254da6cfd2725bdad6d1a79fefc1a99825dcdfb001edb002747635e818790b8911ede0ff3d824f8136de630b6ca735fbdcf28a77494069959052bfcd2d25074d4d51863084870a181789;
    5'b00111 : xpb = 1024'h189a05734f52651006abeb5f55e7414bce48aeac83e0db733a3bd6fd3441f58845b48016399f4f7a62d59dc55c34821573fca066622e5e234fd7eaf5b6b191d70582b99a2899574b81de5724de88e72c6b8df2f3cb5ee2bd683d04c3930fa4eb16616666cc2f0303606b2efb51e1220452a064dad0784aac6626061cca4bb50e;
    5'b01000 : xpb = 1024'h2e06a09d13c22d10f3169975fd6d2b8b6f91050783908729e496d82d901db5173c3ee2cb742db09c7e6ab452453248de3f86878b46496f8f8e0037911884cdc63658372a79a88ba240cac5c0d0f59e2a133cd6e8b34b38cef7acc04d69e12f7c9b7602662622914365f14b63a2cb3b5e5739c9099a34807461b87b28a7f5293;
    5'b01001 : xpb = 1024'h9dd413f61514155ae2bc5fa67a20ab77111f75254208d5e98033bd5e30c46e22a51bd9bbff0ce527cc55f80bcfcfd7d0b80e5871294da01a52875b5aa7317c93359781f9d62cb76dd8d50435d47190c9cadea181d790b16d2c452540d4572396ac14ec0fa95e47b29312e1501a486b90c720b328b319a2926c80844cd3955683;
    5'b01010 : xpb = 1024'h881a788c96fdd31beb41ddde84103ce3f9cfd6c9366102e8e44153e3d58453ebd32b47d27cb070b73167058b97ee7a49280a20837b83d8effb8f73de02083798937a4bd2552de8dc7b03596d02f8038000847bfc9766823cb382ec8217e591a35f6ae5cf3f916dc36906c70b0293fd4259f3eade7c449fed4c7605e293c8f408;
    5'b01011 : xpb = 1024'h7260dd2318e790dcf3c75c168dffce50e280386d2ab92fe8484eea697a4439b5013ab5e8fa53fc469678130b600d1cc19805e895cdba11c5a4978c615cdef29df15d15aad42f1a4b1d31aea4317e7636362a5677573c530c3ac0b3c35b73ffb012c0df8ed5c493d43efaacc5eadf8ef3ecc72294456f9d482c6b877853fc918d;
    5'b01100 : xpb = 1024'h5ca741b99ad14e9dfc4cda4e97ef5fbdcb309a111f115ce7ac5c80ef1f041f7e2f4a23ff77f787d5fb89208b282bbf3a0801b0a81ff04a9b4d9fa4e4b7b5ada34f3fdf8353304bb9bf6003db6004e8ec6bd030f2171223dbc1fe7b049f026dbcc616d94e6bf7b9e514ee9280d32b20a57f9a5a4a0e9a9aa30c61090e14302f12;
    5'b01101 : xpb = 1024'h46eda6501cbb0c5f04d25886a1def12ab3e0fbb5136989e7106a1774c3c405475d599215f59b1365609a2e0af04a61b277fd78ba72268370f6a7bd68128c68a8ad22a95bd2317d28618e59128e8b5ba2a1760b6cd6e7f4ab493c4245e290dbc9796cd30e022adff5eae2783bbb76b257126d91ffd7c597fdec568aa3d463cc97;
    5'b01110 : xpb = 1024'h31340ae69ea4ca200d57d6beabce82979c915d5907c1b6e67477adfa6883eb108b69002c733e9ef4c5ab3b8ab869042ae7f940ccc45cbc469fafd5eb6d6323ae0b0573345132ae9703bcae49bd11ce58d71be5e796bdc57ad07a0987261f49d62cc2cccd985e0606c0d65df6a3c24408a540c9b5a0f09558cc4c0c3994976a1c;
    5'b01111 : xpb = 1024'h1b7a6f7d208e87e115dd54f6b5be14048541befcfc19e3e5d88544800d43d0d9b9786e42f0e22a842abc490a8087a6a357f508df1692f51c48b7ee6ec839deb368e83d0cd033e005a5eb0380eb98410f0cc1c0625693964a57b7d0c869adb7e2e018c68d2e912c1796ca43b18c0dd5ba3814016b6a1b92b3ac418dcf54cb07a1;
    5'b10000 : xpb = 1024'h5c0d413a27845a21e62d32ebfada5716df220a0f07210e53c92db05b203b6a2e787dc596e85b6138fcd568a48a6491bc7f0d0f168c92df1f1c006f2231099b8c6cb06e54f351174481958b81a1eb3c542679add16696719def59809ad3c25ef936ec04cc4c452286cbe296c7459676bcae739213346900e8c370f6514fea526;
    5'b10001 : xpb = 1024'ha0b47dffe650382bf1edc93dd9f77e2fc8188575ba41de5c1e7d2ae109c6497418dfc7e8b64fc031943ca350f422fc5e9c06c0e9ddb237134b675ed3b8b9c96f98fd056c7dc74027fce1b091e180eaac6c126ef062c564fa1bbff145aaf5368e75cc4c360bc070c6c971f60654751f46ac944fb94cbcea99b29c0bff5e14a916;
    5'b10010 : xpb = 1024'h8afae2966839f5ecfa734775e3e70f9cb0c8e719ae9a0b5b828ac166ae862f3d46ef35ff33f34bc0f94db0d0bc419ed70c0288fc2fe86fe8f46f775713908474f6dfcf44fcc871969f1005c910075d62a1b8496b229b35c9a2fdb886ee83a49b292245f5a1f396d79f65dbc13cc0b0f83f67876f15e7e7f492918d951e48469b;
    5'b10011 : xpb = 1024'h7541472cea23b3ae02f8c5adedd6a109997948bda2f2385ae69857ec5346150674fea415b196d7505e5ebe508460414f7bfe510e821ea8be9d778fda6e673f7a54c2991d7bc9a305413e5b003e8dd018d75e23e5e27106992a3b7fc8321212a7dc783fb53826bce87559c17c250c42a9d23abf24df12e54f72870f2ade7be420;
    5'b10100 : xpb = 1024'h5f87abc36c0d716f0b7e43e5f7c632768229aa61974a655a4aa5ee71f805facfa30e122c2f3a62dfc36fcbd04c7ee3c7ebfa1920d454e194467fa85dc93dfa7fb2a562f5facad473e36cb0376d1442cf0d03fe60a246d768b179470975a080b48fce3974ce59e2f94b4da7370d57d45b650df6daa83de2aa527c90c09eaf81a5;
    5'b10101 : xpb = 1024'h49ce1059edf72f301403c21e01b5c3e36ada0c058ba29259aeb384f79cc5e098d11d8042acddee6f2880d950149d86405bf5e133268b1a69ef87c0e12414b58510882cce79cc05e2859b056e9b9ab58542a9d8db621ca83838b70e4ab92eeec143243334648d090a21418cf1f5a3660cf7e12e907168e005327212565ee31f2a;
    5'b10110 : xpb = 1024'h341474f06fe0ecf11c8940560ba55550538a6da97ffabf5912c11b7d4185c661ff2cee592a8179fe8d91e6cfdcbc28b8cbf1a94578c1533f988fd9647eeb708a6e6af6a6f8cd375127c95aa5ca21283b784fb35621f27907bff4d58bfcbd5ccdf67a2cf3fac02f1af73572acddeef7be8ab466463a93dd60126793ec1f16bcaf;
    5'b10111 : xpb = 1024'h1e5ad986f1caaab2250ebe8e1594e6bd3c3acf4d7452ec5876ceb202e645ac2b2d3c5c6fa825058df2a2f44fa4dacb313bed7157caf78c154197f1e7d9c22b8fcc4dc07f77ce68bfc9f7afdcf8a79af1adf58dd0e1c849d747329ccd404bcadaa9d026b390f3552bcd295867c63a89701d879dfc03bedabaf25d1581df4a5a34;
    5'b11000 : xpb = 1024'h8a13e1d73b468732d943cc61f84782a24eb30f168ab1957dadc48888b0591f45b4bca8625c8911d57b401cf6cf96da9abe9396a1d2dc4eaeaa00a6b3498e6952a308a57f6cf9a2e6c260514272e0da7e39b684ba19e1aa6ce70640e83da38e75d26207327267b3ca31d3e22ae861b21b05ad5b1cce9d815d25297179f7df7b9;
    5'b11001 : xpb = 1024'ha394e809b78c5afd011f32d539ce50e87f1195c6327ae6cebcc69863e2c824c58ca3b6156d929b3b5c234e96187620ec7fff29629216ce0c4447624cca42164bfc6288df2561c8e220ee5cedee90448f0d463c5eedfa18870b3abd4a819349863f83ac5c6e2299daffd10abc8ea1d2fc9207ec49e66032a0f8b793b1e893fba9;
    5'b11010 : xpb = 1024'h8ddb4ca0397618be09a4b10d43bde25567c1f76a26d313ce20d42ee987880a8ebab3242beb3626cac1345c15e094c364effaf174e44d06e1ed4f7ad02518d1515a4552b7a462fa50c31cb2251d16b74542ec16d9adcfe9569278848bc521b792f2d9a61c0455bfebd5c4f07776ed64ae24db23ffaf8b2ffbd8ad1547a8c7992e;
    5'b11011 : xpb = 1024'h7821b136bb5fd67f122a2f454dad73c25072590e1b2b40cd84e1c56f2c47f057e8c2924268d9b25a26456995a8b365dd5ff6b98736833fb7965793537fef8c56b8281c9023642bbf654b075c4b9d29fb7891f1546da5ba2619b64bcd08b0259fa62f9fdb9a88e5fcabb8d6325f38f65fb7ae5bb578b62d56b8a296dd68fb36b3;
    5'b11100 : xpb = 1024'h626815cd3d4994401aafad7d579d052f3922bab20f836dcce8ef5bf4d107d62116d20058e67d3de98b56771570d20855cff2819988b9788d3f5fabd6dac6475c160ae668a2655d2e07795c937a239cb1ae37cbcf2d7b8af5a0f4130e4c3e93ac5985999b30bc0c0d81acbbed478488114a81936b41e12ab198981873292ed438;
    5'b11101 : xpb = 1024'h4cae7a63bf33520123352bb5618c969c21d31c5603db9acc4cfcf27a75c7bbea44e16e6f6420c978f067849538f0aace3fee49abdaefb162e867c45a359d026173edb04121668e9ca9a7b1caa8aa0f67e3dda649ed515bc52831da4f8fcd01b90cdb935ac6ef321e57a0a1a82fd019c2dd54cb210b0c280c788d9a08e96271bd;
    5'b11110 : xpb = 1024'h36f4defa411d0fc22bbaa9ed6b7c28090a837df9f833c7cbb10a89001a87a1b372f0dc85e1c4550855789215010f4d46afea11be2d25ea38916fdcdd9073bd66d1d07a19a067c00b4bd60701d730821e198380c4ad272c94af6fa190d35b6fc5c0318d1a5d22582f2d948763181bab74702802d6d437256758831b9ea9960f42;
    5'b11111 : xpb = 1024'h213b4390c306cd8334402825756bb975f333df9dec8bf4cb15181f85bf47877ca1004a9c5f67e097ba899f94c92defbf1fe5d9d07f5c230e3a77f560eb4a786c2fb343f21f68f179ee045c3905b6f4d44f295b3f6cfcfd6436ad68d216e9ddd2738786d9f3557e4003886d1e00673d2602fb3a8c9d6222c238789d3469c9acc7;
    endcase
end

endmodule

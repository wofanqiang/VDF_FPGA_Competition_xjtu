module xpb_5_270
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h9df7a0f7e484979cf2a53face20c45c1de896529d7b3da2cdab0f66006a933b9cd68e436dd1a80e4f686611ef1b5d3314a8f4f901523fddafaf3eec3db9c295af25f0447fc0c49f8d91f7191527c938075c1e36d684d7cfa5936cc5d73f8424dbf6cab424155a8000122cec3e684303d7ee935ce968a5c92c37f0968ddca1065;
    5'b00010 : xpb = 1024'h8b41fc9a071afa711a450782b3be44324b9cc722d9f013e23785336a5a4fba6b97894af4f00e833b4dae82f7000d95983104773a07952b6a45489e297c65de04706ed3e1488796ac9fa4e0800c1d62cff77ecd424414cce3fce106c02dc5e2094fd1c45ad1e257727b85b6a8d5383a51aef88cbadcc95bf5408e97cd32b1ba5f;
    5'b00011 : xpb = 1024'h788c583c29b15d4541e4cf58857042a2b8b0291bdc2c4d9794597074adf6411d61a9b1b303028591a4d6a4cf0e6557ff17799ee3fa0658f98f9d4d8f1d2f92adee7ea37a9502e360662a4f6ec5be321f793bb7171fdc1ccda08b4122e79381c4e036dd73626f06e4f5e89e8dc3ec4465df07e3a723085b57bd9e263187996459;
    5'b00100 : xpb = 1024'h65d6b3de4c47c0196984972e5722411325c38b14de68874cf12dad7f019cc7cf2bca187115f687e7fbfec6a71cbd1a65fdeec68dec778688d9f1fcf4bdf947576c8e7313e17e30142cafbe5d7f5f016efaf8a0ebfba36cb744357b85a1612180709bf68bf2fbb657704b8672b2a04e7a0f173a9369475aba3aadb495dc810e53;
    5'b00101 : xpb = 1024'h53210f806ede22ed91245f0428d43f8392d6ed0de0a4c1024e01ea8955434e80f5ea7f2f28ea8a3e5326e87f2b14dccce463ee37dee8b4182446ac5a5ec2fc00ea9e42ad2df97cc7f3352d4c38ffd0be7cb58ac0d76abca0e7dfb5e85b2ec13c01010fa4838865c9eaae6e57a154588e3f26917faf865a1cb7bd42fa3168b84d;
    5'b00110 : xpb = 1024'h406b6b22917485c1b8c426d9fa863df3ffea4f06e2e0fab7aad62793a8e9d532c00ae5ed3bde8c94aa4f0a57396c9f33cad915e1d159e1a76e9b5bbfff8cb0aa68ae12467a74c97bb9ba9c3af2a0a00dfe727495b3320c8a8b89f04b14fc60f7916628bd1415153c6511563c900862a26f35e86bf5c5597f34ccd15e86506247;
    5'b00111 : xpb = 1024'h2db5c6c4b40ae895e063eeafcc383c646cfdb0ffe51d346d07aa649dfc905be48a2b4cab4ed28eeb01772c2f47c4619ab14e3d8bc3cb0f36b8f00b25a0566553e6bde1dfc6f0162f80400b29ac416f5d802f5e6a8ef95c742f342aadceca00b321cb41d5a4a1c4aedf743e217ebc6cb69f453f583c0458e1b1dc5fc2db380c41;
    5'b01000 : xpb = 1024'h1b002266d6a14b6a0803b6859dea3ad4da1112f8e7596e22647ea1a85036e296544bb36961c69141589f4e07561c240197c36535b63c3cc60344ba8b412019fd64cdb179136b62e346c57a1865e23ead01ec483f6ac0ac5dd2de65108897a06eb2305aee352e742159d726066d7076cacf549644824358442eebee27301fb63b;
    5'b01001 : xpb = 1024'h84a7e08f937ae3e2fa37e5b6f9c3945472474f1e995a7d7c152deb2a3dd69481e6c1a2774ba9397afc76fdf6473e6687e388cdfa8ad6a554d9969f0e1e9cea6e2dd81125fe6af970d4ae9071f830dfc83a932144687fc4776889f734265402a42957406c5bb2393d43a0deb5c2480deff63ed30c88257a6abfb7c8b85076035;
    5'b01010 : xpb = 1024'ha6421f00ddbc45db2248be0851a87f0725adda1bc14982049c03d512aa869d01ebd4fe5e51d5147ca64dd0fe5629b999c8c7dc6fbdd16830488d58b4bd85f801d53c855a5bf2f98fe66a5a9871ffa17cf96b1581aed57941cfbf6bd0b65d827802021f490710cb93d55cdcaf42a8b11c7e4d22ff5f0cb4396f7a85f462d1709a;
    5'b01011 : xpb = 1024'h938c7aa30052a8af49e885de235a7d7792c13c14c385bbb9f8d8121cfe2d23b3b5f5651c64c916d2fd75f2d664817c00af3d0419b04295bf92e2081a5e4facab534c54f3a86e4643acefc9872ba070cc7b27ff568a9cc92b7369a633702b223392673861979d7b064fbfc494315cbb30ae5c79eba54bb39bec8a1458b7b91a94;
    5'b01100 : xpb = 1024'h80d6d64522e90b8371884db3f50c7be7ffd49e0dc5c1f56f55ac4f2751d3aa658015cbda77bd1929549e14ae72d93e6795b22bc3a2b3c34edd36b77fff196154d15c248cf4e992f773753875e541401bfce4e92b666419151713e09629f8c1ef22cc517a282a2a78ca22ac792010c544de6bd0d7eb8ab2fe6999a2bd0ca0c48e;
    5'b01101 : xpb = 1024'h6e2131e7457f6e5799281589c6be7a586ce80006c7fe2f24b2808c31a57a31174a3632988ab11b7fabc63686813100ce7c27536d9524f0de278b66e59fe315fe4f6bf4264164dfab39faa7649ee20f6b7ea1d300422b68febabe1af8e3c661aab3316a92b8b6d9eb4485945e0ec4cf590e7b27c431c9b260e6a9312161886e88;
    5'b01110 : xpb = 1024'h5b6b8d896815d12bc0c7dd5f987078c8d9fb61ffca3a68da0f54c93bf920b7c9145699569da51dd602ee585e8f88c335629c7b1787961e6d71e0164b40accaa7cd7bc3bf8de02c5f008016535882debb005ebcd51df2b8e85e68555b9d940166439683ab4943895dbee87c42fd78d96d3e8a7eb07808b1c363b8bf85b6701882;
    5'b01111 : xpb = 1024'h48b5e92b8aac33ffe867a5356a227739470ec3f8cc76a28f6c2906464cc73e7ade770014b099202c5a167a369de0859c4911a2c17a074bfcbc34c5b0e1767f514b8b9358da5b7912c70585421223ae0a821ba6a9f9ba08d202128fbe5761a121d3fb9cc3d9d038d0394b6427ec2ce3816e99d59cbe47b125e0c84dea0b57c27c;
    5'b10000 : xpb = 1024'h360044cdad4296d410076d0b3bd475a9b42225f1ceb2dc44c8fd4350a06dc52ca89766d2c38d2282b13e9c0eac3848032f86ca6b6c78798c06897516824033fac99b62f226d6c5c68d8af430cbc47d5a03d8907ed58158bba5bcca21112f40dd6460b5dc6a5ce842b3ae4c0cdae0ed959ea92c890486b0885dd7dc4e603f6c76;
    5'b10001 : xpb = 1024'h234aa06fcfd8f9a837a734e10d86741a213587ead0ef15fa25d1805af4144bde72b7cd90d68124d90866bde6ba900a6a15fbf2155ee9a71b50de247c2309e8a447ab328b7352127a5410631f85654ca985957a53b148a8a549670483cafce098f4c5cef4fae997b52e1133f1c994f7a9ceb883754ac5afeadae76ab2b5271670;
    5'b10010 : xpb = 1024'h1094fc11f26f5c7c5f46fcb6df38728a8e48e9e3d32b4faf82a5bd6547bad2903cd8344ee975272f5f8edfbec8e7ccd0fc7119bf515ad4aa9b32d3e1c3d39d4dc5bb0224bfcd5f2e1a95d20e3f061bf9075264288d0ff88eed113ee684ca8054852ae80d8b764727a8741bd6b84901bdfec7da619104af4d57f6f9170a0ec06a;
    5'b10011 : xpb = 1024'hae8c9d09d6f3f41951ec3c63c144b84c6cd24f0daadf29dc5d56b3c54e64064a0a411885c68fa814561540ddba9da0024700694f667ed2859626c2a59f6fc6a8b81a066cbbd9a926f3b5439f9182af797d144795f55d758946480b43f8c2c2a24497934fcccbef27a996ea9a9ecd31fb7db11030278f0be01b76027fe7d8d0cf;
    5'b10100 : xpb = 1024'h9bd6f8abf98a56ed798c043992f6b6bcd9e5b106ad1b6391ba2af0cfa20a8cfbd4617f43d983aa6aad3d62b5c8f562692d7590f958f00014e07b720b40397b523629d6060854f5daba3ab28e4b237ec8fed1316ad124c572e9f245a6b290625dd4fcac685d589e9a23f9d27f8d813c0fadc0671c6dce0b42988590e43cc07ac9;
    5'b10101 : xpb = 1024'h8921544e1c20b9c1a12bcc0f64a8b52d46f912ffaf579d4716ff2dd9f5b113ad9e81e601ec77acc10465848dd74d24d013eab8a34b612da42ad02170e1032ffbb439a59f54d0428e80c0217d04c44e18808e1b3facec155c8d9c80096c5e02196561c580ede54e0c9e5cba647c354623ddcfbe08b40d0aa515951f4891a824c3;
    5'b10110 : xpb = 1024'h766baff03eb71c95c8cb93e5365ab39db40c74f8b193d6fc73d36ae449579a5f68a24cbfff6baf175b8da665e5a4e736fa5fe04d3dd25b337524d0d681cce4a532497538a14b8f424745906bbe651d68024b051488b365463146ba6c262ba1d4f5c6de997e71fd7f18bfa2496ae950380ddf14f4fa4c0a0792a4adace68fcebd;
    5'b10111 : xpb = 1024'h63b60b92614d7f69f06b5bbb080cb20e211fd6f1b3d010b1d0a7a7ee9cfe211132c2b37e125fb16db2b5c83df3fca99de0d507f7304388c2bf79803c2296994eb05944d1edc6dbf60dcaff5a7805ecb78407eee9647ab52fd4f0f4cedff94190862bf7b20efeacf193228a2e599d5a4c3dee6be1408b096a0fb43c113b7778b7;
    5'b11000 : xpb = 1024'h5100673483e3e23e180b2390d9beb07e8e3338eab60c4a672d7be4f8f0a4a7c2fce31a3c2553b3c409ddea1602546c04c74a2fa122b4b65209ce2fa1c3604df82e69146b3a4228a9d4506e4931a6bc0705c4d8be40420519789b2f3199c6e14c169110ca9f8b5c640d857213485164606dfdc2cd86ca08cc8cc3ca75905f22b1;
    5'b11001 : xpb = 1024'h3e4ac2d6a67a45123faaeb66ab70aeeefb469ae3b848841c8a502203444b2e74c70380fa3847b61a61060bee10ac2e6badbf574b1525e3e15422df07642a02a1ac78e40486bd755d9ad5dd37eb478b568781c2931c0955031c45699453948107a6f629e330180bd687e859f837056e749e0d19b9cd09082f09d358d9e546ccab;
    5'b11010 : xpb = 1024'h2b951e78c910a7e6674ab33c7d22ad5f6859fcdcba84bdd1e7245f0d97f1b5269123e7b84b3bb870b82e2dc61f03f0d294347ef5079711709e778e6d04f3b74b2a88b39dd338c211615b4c26a4e85aa6093eac67f7d0a4ecbfefa3f70d6220c3375b42fbc0a4bb49024b41dd25b97888ce1c70a61348079186e2e73e3a2e76a5;
    5'b11011 : xpb = 1024'h18df7a1aeba70aba8eea7b124ed4abcfd56d5ed5bcc0f78743f89c17eb983bd85b444e765e2fbac70f564f9e2d5bb3397aa9a69efa083effe8cc3dd2a5bd6bf4a89883371fb40ec527e0bb155e8929f58afb963cd397f4d66399de59c72fc07ec7c05c1451316abb7cae29c2146d829cfe2bc792598706f403f275a28f16209f;
    5'b11100 : xpb = 1024'h629d5bd0e3d6d8eb68a42e82086aa404280c0cebefd313ca0ccd9223f3ec28a2564b5347123bd1d667e71763bb375a0611ece48ec796c8f3320ed384687209e26a852d06c2f5b78ee662a041829f9450cb88011af5f44c0074418bc80fd603a5825752ce1be1a2df71111a703218cb12e3b1e7e9fc6065681020406e3fdca99;
    5'b11101 : xpb = 1024'ha42176b4f2c2052ba92f82950292f002210a25f896b10b697b7dcf8245e7f643f2cd996b4e3e3e025d04d2952d6948d1abae1dd9019d6a6a2e14dbfc222349f919075718683ba571c7859b956aa68cc5827a637f17acc1ba607ae519f4f5a2881792206f2313c22df833e06ae9a5bceead24544d365062e944810d6fc1c7dafe;
    5'b11110 : xpb = 1024'h916bd257155867ffd0cf4a6ad444ee728e1d87f198ed451ed8520c8c998e7cf5bcee002961324058b42cf46d3bc10b3892234582f40e97f978698b61c2ecfea2971726b1b4b6f2258e0b0a8424475c1504374d53f37411a404251f7caec34243a7f73987b3a071a07296c84fd859c702dd33ab397c8f624bc1909bd416af84f8;
    5'b11111 : xpb = 1024'h7eb62df937eecad3f86f1240a5f6ece2fb30e9ea9b297ed435264996ed3503a7870e66e7742642af0b5516454a18cd9f78986d2ce67fc588c2be3ac763b6b34c1526f64b01323ed954907972dde82b6485f43728cf3b618da7cf59df6890e1ff385c52a0442d2112ecf9b034c70dd1170d430225c2ce61ae3ea02a386b972ef2;
    endcase
end

endmodule

module xpb_5_190
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h9c7a8d393141bf4a2cc994be7c833eb09b12d6ebfc1345acb25dbaa332404e5c944d72edc1e8033685907703d492838a42b0f2f5109d5baf6e9c0eb29c85e8fc0a92a27cc4d9a88f516d51bd1d492941629881dcb8fdfa171041427a709b4f9efbee3d68ff4d44ec7d01d16f8b25e22058719d1b1f98e85199cb751849be5ed9;
    5'b00010 : xpb = 1024'h8847d51ca09549cb8e8db1a5e8ac360fc4afaaa722aeeae1e6debbf0b17defb125526862b9a987de6bc2aec0c5c6f64a2147be03fe87e7132c98de06fe395d46a0d6104ada2253d99040a0d7a1b68e51d12c0a20e575c71d6af5f2fa270bfcabc8d4e8a84dd1914b7343bc001e7b9e1762095b53eee67372ed276f2c0a9a5747;
    5'b00011 : xpb = 1024'h74151d000fe8d44cf051ce8d54d52d6eee4c7e62494a90171b5fbd3e30bb9105b6575dd7b16b0c8651f4e67db6fb6909ffde8912ec727276ea95ad5b5fecd19137197e18ef6aff23cf13eff22623f3623fbf926511ed9423c5aaa379dd7ca9b895bb93e79c55ddaa6985a690b1d15a0e6ba1198cbe33fe944083693fcb764fb5;
    5'b00100 : xpb = 1024'h5fe264e37f3c5ece5215eb74c0fe24ce17e9521d6fe6354c4fe0be8baff9325a475c534ca92c912e38271e3aa82fdbc9de755421da5cfddaa8927cafc1a045dbcd5cebe704b3aa6e0de73f0caa915872ae531aa93e65612a205f53f993ed56c562a23f26eada2a095fc79121452716057538d7c58d8189b593df63538c524823;
    5'b00101 : xpb = 1024'h4bafacc6ee8fe94fb3da085c2d271c2d418625d89681da818461bfd92f36d3aed86148c1a0ee15d61e5955f799644e89bd0c1f30c847893e668f4c042353ba2663a059b519fc55b84cba8e272efebd831ce6a2ed6add2e307b1404794a5e03d22f88ea66395e766856097bb1d87cd1fc7ed095fe5ccf14d6e73b5d674d2e4091;
    5'b00110 : xpb = 1024'h377cf4aa5de373d1159e25439950138c6b22f993bd1d7fb6b8e2c126ae74750369663e3698af9a7e048b8db48a98c1499ba2ea3fb63214a2248c1b5885072e70f9e3c7832f4501028b8ddd41b36c22938b7a2b319754fb36d5c8b4f900ceb0defc6f95a587e2c2c74c4b66426bd28df3886854372c1c9ff83a97577b0e0a38ff;
    5'b00111 : xpb = 1024'h234a3c8dcd36fe527762422b05790aeb94bfcd4ee3b924ebed63c2742db21657fa6b33ab90711f25eabdc5717bcd34097a39b54ea41ca005e288eaace6baa2bb90273551448dac4cca612c5c37d987a3fa0db375c3ccc83d307d6578b73f5debc95640e4d6670f26428d50d2ff2849ea9200126ffb6a2b198df3518ecee6316d;
    5'b01000 : xpb = 1024'hf1784713c8a88d3d9265f1271a2024abe5ca10a0a54ca2121e4c3c1acefb7ac8b7029208832a3cdd0effd2e6d01a6c958d0805d92072b69a085ba01486e1706266aa31f59d6579709347b76bc46ecb468a13bb9f04495438b3215f86db00af8963cec2424eb5b8538cf3b63927e05e19b97d0a8cab7b63ae14f4ba28fc229db;
    5'b01001 : xpb = 1024'hab9211aa6dcc481e05eff3d0ee2540fb596f77f606680fcdd4427e64df3006091fbd9c0e4a1aa7045680743241942a539b817352a2a487190f21c8b3e4f4000230fd459c1eb000265aa1cd33d99015f5cb39bd96a9428f5a9b735872de4b5a97922b298d2438a071b5d10cd31da3e801f4096dc3ea509e8c7b1ac0bad98088b4;
    5'b01010 : xpb = 1024'h975f598ddd1fd29f67b410b85a4e385a830c4bb12d03b50308c37fb25e6da75db0c2918341dc2bac3cb2abef32c89d137a183e61908f127ccd1e980846a7744cc740b36a33f8ab7099751c4e5dfd7b0639cd45dad5ba5c60f62808f294bc07a45f11d4cc72bcecd0ac12f763b0f9a3f8fda12bfcb99e29adce76bace9a5c8122;
    5'b01011 : xpb = 1024'h832ca1714c735d20c9782d9fc6772fb9aca91f6c539f5a383d4480ffddab48b241c786f8399db05422e4e3ac23fd0fd358af09707e799de08b1b675ca85ae8975d842138494156bad8486b68e26ae016a860ce1f0232296750dcb9724b2cb4b12bf8800bc141392fa254e1f4444f5ff00738ea3588ebb4cf21d2b4e25b387990;
    5'b01100 : xpb = 1024'h6ef9e954bbc6e7a22b3c4a8732a02718d645f3277a3aff6d71c5824d5ce8ea06d2cc7c6d315f34fc09171b69153182933745d47f6c642944491836b10a0e5ce1f3c78f065e8a0205171bba8366d8452716f456632ea9f66dab9169f2019d61bdf8df2b4b0fc5858e9896cc84d7a51be710d0a86e58393ff0752eaef61c1471fe;
    5'b01101 : xpb = 1024'h5ac731382b1a72238d00676e9ec91e77ffe2c6e2a0d6a4a2a646839adc268b5b63d171e22920b9a3ef4953260665f55315dc9f8e5a4eb4a8071506056bc1d12c8a0afcd473d2ad4f55ef099deb45aa378587dea75b21c37406461a71b80e0ecac5c5d68a5e49d1ed8ed8b7156afad7de1a6866a72786cb11c88aa909dcf06a6c;
    5'b01110 : xpb = 1024'h4694791b9a6dfca4eec484560af215d7297f9a9dc77249d7dac784e85b642caff4d6675720e23e4bd57b8ae2f79a6812f4736a9d4839400bc511d559cd754577204e6aa2891b589994c258b86fb30f47f41b66eb8799907a60facaf16e7ebbd792ac81c9acce1e4c851aa1a5fe5093d5240024dff6d456331be6a31d9dcc62da;
    5'b01111 : xpb = 1024'h3261c0ff09c187265088a13d771b0d36531c6e58ee0def0d0f488635daa1ce0485db5ccc18a3c2f3bbadc29fe8cedad2d30a35ac3623cb6f830ea4ae2f28b9c1b691d8709e6403e3d395a7d2f420745862aeef2fb4115d80bbaf7b7124ef68e45f932d08fb526aab7b5c8c3691a64fcc2d97e318c621e1546f429d315ea85b48;
    5'b10000 : xpb = 1024'h1e2f08e2791511a7b24cbe24e34404957cb9421414a9944243c9878359df6f5916e052411065479ba1dffa5cda034d92b1a100bb240e56d3410b740290dc2e0c4cd5463eb3acaf2e1268f6ed788dd968d1427773e0892a8716642bf0db6015f12c79d84849d6b70a719e76c724fc0bc3372fa151956f6c75c29e97451f8453b6;
    5'b10001 : xpb = 1024'h9fc50c5e8689c291410db0c4f6cfbf4a65615cf3b453977784a88d0d91d10ada7e547b60826cc4388123219cb37c0529037cbca11f8e236ff084356f28fa256e318b40cc8f55a78513c4607fcfb3e793fd5ffb80d00f78d7118dc7091d0c2fdf9608387985b036967e06157b851c7ba40c75f8a64bcf79715fa9158e0604c24;
    5'b10010 : xpb = 1024'ha676ddff19aa5b7340da6fcacbf03aa54168ecbb37587f242aa843740b5d5f0a3c32baa3ca0ecf7a0da2a91d9fca43dcd2e8bebf22963de66da452098f158b52edab56898dcf0307a2a997c51a4467baa26e8194c5fef1a4815a1eeb026c129cf54ec0f097a84855e4e232c74377a9da9938fca58455dfe8afc606712a1eaafd;
    5'b10011 : xpb = 1024'h924425e288fde5f4a29e8cb2381932046b05c0765df424595f2944c18a9b005ecd37b018c1d05421f3d4e0da90feb69cb17f89ce1080c94a2ba1215df0c8ff9d83eec457a317ae51e17ce6df9eb1cccb110209d8f276beaadc0ecf6ab8dcbfa9c2356c2fe62c94b4db241d57d6cd65d1a2d0bade53a36b0a03220084eafaa36b;
    5'b10100 : xpb = 1024'h7e116dc5f85170760462a999a442296394a29431848fc98e93aa460f09d8a1b35e3ca58db991d8c9da0718978233295c901654dcfe6b54ade99df0b2527c73e81a323225b860599c205035fa231f31db7f95921d1eee8bb136c37fea6f4d6cb68f1c176f34b0e113d16607e86a2321c8ac68791722f0f62b567dfa98abd69bd9;
    5'b10101 : xpb = 1024'h69deb5a967a4faf76626c681106b20c2be3f67ecab2b6ec3c82b475c89164307ef419b02b1535d71c039505473679c1c6ead1febec55e011a79ac006b42fe832b0759ff3cda904e65f238514a78c96ebee291a614b6658b79178306a25be19c35c02c2ae83352d72c7a7f278fd78ddbfb600374ff23e814ca9d9f4ac6cb29447;
    5'b10110 : xpb = 1024'h55abfd8cd6f88578c7eae3687c941821e7dc3ba7d1c713f8fcac48aa0853e45c80469077a914e219a66b8811649c0edc4d43eafada406b7565978f5b15e35c7d46b90dc1e2f1b0309df6d42f2bf9fbfc5cbca2a577de25bdec2ce0e9dc2ec6d028e96dedd1b979d1bde9dd0990ce99b6bf97f588c18c0c6dfd35eec02d8e8cb5;
    5'b10111 : xpb = 1024'h41794570464c0ffa29af004fe8bd0f8111790f62f862b92e312d49f7879185b1114b85eca0d666c18c9dbfce55d0819c2bdab609c82af6d923945eaf7796d0c7dcfc7b8ff83a5b7adcca2349b067610ccb502ae9a455f2c446e19169929f73dcf5d0192d203dc630b42bc79a242455adc92fb3c190d9978f5091e8d3ee6a8523;
    5'b11000 : xpb = 1024'h2d468d53b59f9a7b8b731d3754e606e03b15e31e1efe5e6365ae4b4506cf2705a2507b619897eb6972cff78b4704f45c0a718118b615823ce1912e03d94a4512733fe95e0d8306c51b9d726434d4c61d39e3b32dd0cdbfcaa19641e9491020e9c2b6c46c6ec2128faa6db22ab77a11a4d2c771fa602722b0a3ede2e7af467d91;
    5'b11001 : xpb = 1024'h1913d53724f324fced373a1ec10efe3f64b2b6d9459a03989a2f4c92860cc85a335570d69059701159022f483839671be9084c27a4000da09f8dfd583afdb95d0983572c22cbb20f5a70c17eb9422b2da8773b71fd458cd0fc4af268ff80cdf68f9d6fabbd465eeea0af9cbb4acfcd9bdc5f30332f74add1f749dcfb702275ff;
    5'b11010 : xpb = 1024'h4e11d1a9446af7e4efb57062d37f59e8e4f8a946c35a8cdceb04de0054a69aec45a664b881af4b93f346705296dd9dbc79f173691ea99045d8accac9cb12da79fc6c4fa38145d59994410993daf903e170ac3b629bd59d756ffa2e8b5f17b035c841aeb0bcaab4d96f1874bde258992e5f6ee6bfec238f34aa5d70f30fe6e6d;
    5'b11011 : xpb = 1024'ha15baa53c5886ec87bc4ebc4a9bb344f296261806848ee7a810e0883378ab80b58a7d9394a02f7efc4c4de08fe005d660a500a2ba287f4b3cc26db5f393716a3aa596776fcee05e8eab162565af8b97f79a34592e2bb53ee6740e563268ccaa2587258540b17f03a13f358bb694b6bb33e688b871e5b2144e4714c277abccd46;
    5'b11100 : xpb = 1024'h8d28f23734dbf949dd8908ac15e42bae52ff353b8ee493afb58f09d0b6c8595fe9acceae41c47c97aaf715c5ef34d025e8e6d53a907280178a23aab39aea8aee409cd5451236b1332984b170df661e8fe836cdd70f3320f4c1f595e2dcfd77af25590393599c3c990a35434bfca127aa480049bfeda8ac6637cd463b3b98c5b4;
    5'b11101 : xpb = 1024'h78f63a1aa42f83cb3f4d2593820d230d7c9c08f6b58038e4ea100b1e3605fab47ab1c4233986013f91294d82e06942e5c77da0497e5d0b7b48207a07fc9dff38d6e04313277f5c7d6858008b63d383a056ca561b3baaedfb1caa4662936e24bbf23faed2a82088f800772ddc8ff6e3a1519807f8bcf637878b29404efc74be22;
    5'b11110 : xpb = 1024'h64c381fe13830e4ca111427aee361a6ca638dcb1dc1bde1a1e910c6bb5439c090bb6b998314785e7775b853fd19db5a5a6146b586c4796df061d495c5e5173836d23b0e13cc807c7a72b4fa5e840e8b0c55dde5f6822bb01775ef6e249ded1c8bf265a11f6a4d556f6b9186d234c9f985b2fc6318c43c2a8de853a62bd50b690;
    5'b11111 : xpb = 1024'h5090c9e182d698ce02d55f625a5f11cbcfd5b06d02b7834f53120db934813d5d9cbbaf0d29090a8f5d8dbcfcc2d2286584ab36675a322242c41a18b0c004e7ce03671eaf5210b311e5fe9ec06cae4dc133f166a3949a8807d213a762004f7ed58c0d0551452921b5ecfb02fdb6a25b8f64c7846a5b914dca31e134767e2caefe;
    endcase
end

endmodule

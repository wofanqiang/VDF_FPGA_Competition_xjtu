module xpb_5_680
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h20a53948e0f026bcc7b1818d7744e73ada17e1e65ea27b6d0f9dab2a63839582484c4792d33f5bba727698259867a9dc973058632d39f5caf15dc511ea43745ef0d91de5776de3beb6f8467bca21126b5957cc79e79825f2ed1016136a88da0fca3cddb58d927fe1f5fdde114c4f00832ffe01893e2432a936db9955a8d400ce;
    5'b00010 : xpb = 1024'h414a7291c1e04d798f63031aee89ce75b42fc3ccbd44f6da1f3b5654c7072b0490988f25a67eb774e4ed304b30cf53b92e60b0c65a73eb95e2bb8a23d486e8bde1b23bcaeedbc77d6df08cf7944224d6b2af98f3cf304be5da202c26d511b41f9479bb6b1b24ffc3ebfbbc22989e01065ffc03127c4865526db732ab51a8019c;
    5'b00011 : xpb = 1024'h61efabdaa2d07436571484a865ceb5b08e47a5b31be772472ed9017f2a8ac086d8e4d6b879be132f5763c870c936fd95c591092987ade160d4194f35beca5d1cd28b59b06649ab3c24e8d3735e6337420c07656db6c871d8c730423a3f9a8e2f5eb69920a8b77fa5e1f99a33e4ed01898ffa049bba6c97fba492cc00fa7c026a;
    5'b00100 : xpb = 1024'h8294e52383c09af31ec60635dd139ceb685f87997a89edb43e76aca98e0e560921311e4b4cfd6ee9c9da6096619ea7725cc1618cb4e7d72bc5771447a90dd17bc3647795ddb78efadbe119ef288449ad655f31e79e6097cbb440584daa23683f28f376d63649ff87d7f77845313c020cbff80624f890caa4db6e6556a3500338;
    5'b00101 : xpb = 1024'ha33a1e6c64b0c1afe67787c3545884264277697fd92c69214e1457d3f191eb8b697d65de203ccaa43c50f8bbfa06514ef3f1b9efe221ccf6b6d4d959935145dab43d957b552572b992d9606af2a55c18beb6fe6185f8bdbea1506e6114ac424ef330548bc3dc7f69cdf556567d8b028feff607ae36b4fd4e1249feac4c240406;
    5'b00110 : xpb = 1024'h1332125f83b2b3a3e3239179bb43240fab19483562574416dfd549a8a212d405ae812ff82955a7d00f69519aaf0fea612707ea6ceca8f275f7935f0d42c2458830c77eb21d0259333737a44423eaaa532409d142e10ab6a0d8d3f279c50a79cc8e65a017a0a606be3d334d88d209dce9d11a2a55248dd2c702b61cfd6c159e69;
    5'b00111 : xpb = 1024'h33d74ba864a2da60aad5130732880b4a85312a1bc0f9bf83ef72f4d305966987f6cd778afc95038a81dfe9c04777943dbe3842d019e2e840e8f1241f2d05b9e721a09c9794703cf1ee2feabfee0bbcbe7d619dbcc8a2dc93c5e4088d2f9353dc58a27dcd2e3886a033312b9a1e58dd6d01182bde62b205703991b65314e99f37;
    5'b01000 : xpb = 1024'h547c84f14593011d72869494a9ccf2855f490c021f9c3af0ff109ffd6919ff0a3f19bf1dcfd45f44f45681e5dfdf3e1a55689b33471cde0bda4ee93117492e461279ba7d0bde20b0a528313bb82ccf29d6b96a36b03b0286b2f41ea09a1c2dec22df5b82bbcb0682292f09ab6aa7ddf031162d67a0d63819706d4fa8bdbda005;
    5'b01001 : xpb = 1024'h7521be3a268327da3a3816222111d9c03960ede87e3eb65e0eae4b27cc9d948c876606b0a313baff66cd1a0b7846e7f6ec98f3967456d3d6cbacae43018ca2a50352d862834c046f5c2077b7824de195301136b097d32879a00434b404a507fbed1c3938495d86641f2ce7bcb6f6de7361142ef0defa6ac2a748e8fe6691a0d3;
    5'b01010 : xpb = 1024'h95c6f78307734e9701e997af9856c0fb1378cfcedce131cb1e4bf65230212a0ecfb24e43765316b9d943b23110ae91d383c94bf9a190c9a1bd0a7354ebd01703f42bf647fab9e82e1318be334c6ef4008969032a7f6b4e6c8d144ac76f2de20bb75916edd6f00646152ac5ce0345def69112307a1d1e9d6bde2482540f65a1a1;
    5'b01011 : xpb = 1024'h5beeb762675408afe95a165ff4160e47c1aae84660c0cc0b00ce826e0a2128914b6185d7f6bf3e5ac5c0b0fc5b82ae5b6df7c76ac17ef20fdc8f9089b4116b170b5df7ec296cea7b777020c7db4423aeebbd60bda7d474ec497cee01f8c1989528e6279b3b98d9a8468bd0057c4b950723653210af772e4ce90a0a52f573c04;
    5'b01100 : xpb = 1024'h266424bf07656747c64722f37686481f5632906ac4ae882dbfaa93514425a80b5d025ff052ab4fa01ed2a3355e1fd4c24e0fd4d9d951e4ebef26be1a85848b10618efd643a04b2666e6f488847d554a64813a285c2156d41b1a7e4f38a14f3991ccb402f414c0d7c7a669b11a413b9d3a23454aa491ba58e056c39fad82b3cd2;
    5'b01101 : xpb = 1024'h47095e07e8558e048df8a480edcb2f5a304a72512351039acf483e7ba7a93d8da54ea78325eaab5a91493b5af6877e9ee5402d3d068bdab6e084832c6fc7ff6f52681b49b172962525678f0411f66711a16b6effa9ad93349eb7fb06f49dcda8e7081de4cede8d5e70647922f062ba56d2325633873fd8373c47d35080ff3da0;
    5'b01110 : xpb = 1024'h67ae9750c945b4c155aa260e651016950a62543781f37f07dee5e9a60b2cd30fed9aef15f92a071503bfd3808eef287b7c7085a033c5d081d1e2483e5a0b73ce4341392f28e079e3dc5fd57fdc17797cfac33b799145b9278bc8111a5f26a7b8b144fb9a5c710d40666257343cb1bada023057bcc5640ae073236ca629d33e6e;
    5'b01111 : xpb = 1024'h8853d099aa35db7e1d5ba79bdc54fdcfe47a361de095fa74ee8394d06eb0689235e736a8cc6962cf76366ba62756d25813a0de0360ffc64cc3400d50444ee82d341a5714a04e5da293581bfba6388be8541b07f378dddf1a78d8272dc9af81c87b81d94fea038d225c6035458900bb5d322e594603883d89a9ff05fbd2a73f3c;
    5'b10000 : xpb = 1024'ha8f909e28b26023ae50d29295399e50abe9218043f3875e1fe213ffad233fe147e337e3b9fa8be89e8ad03cbbfbe7c34aad136668e39bc17b49dd2622e925c8c24f374fa17bc41614a50627770599e53ad72d46d6076050d65e83d4134385bd845beb70577960d04525e1356d54fbbe0622c5acf41ac7032e0da9f517b7b400a;
    5'b10001 : xpb = 1024'h18f0fdd5aa27f42ee1b932dfba8484f42733f6b9c86350d78fe231cf82b4e68ec3374855a8c19bb5bbc55caa74c81546dde766e398c0e196f55c5815de035c39a17d5e30df9927daeeaea650a19eec8e12c5a74ebb87fdef9d6bc159e4969355e0f40291545f9458c19c0a8929ce963a43507d762f8545abd146bda29b6cda6d;
    5'b10010 : xpb = 1024'h3996371e8b181aeba96ab46d31c96c2f014bd8a02705cc449f7fdcf9e6387c110b838fe87c00f7702e3bf4d00d2fbf237517bf46c5fad761e6ba1d27c846d09892567c1657070b99a5a6eccc6bbffef96c1d73c8a32023e28a7bd76d4f1f6d65ab30e046e1f2143ab799e89a761d96bd734e7eff6da97855082256f84440db3b;
    5'b10011 : xpb = 1024'h5a3b70676c0841a8711c35faa90e5369db63ba8685a847b1af1d882449bc119353cfd77b4f40532aa0b28cf5a59769000c4817a9f334cd2cd817e239b28a44f7832f99fbce74ef585c9f334835e11164c57540428ab849d5778bed80b9a84775756dbdfc6f84941cad97c6abc26c9740a34c8088abcdaafe3efdf04ded14dc09;
    5'b10100 : xpb = 1024'h7ae0a9b04cf8686538cdb78820533aa4b57b9c6ce44ac31ebebb334ead3fa7159c1c1f0e227faee51329251b3dff12dca378700d206ec2f7c975a74b9ccdb9567408b7e145e2d317139779c4000223d01ecd0cbc72506fc8649c0394243121853faa9bb1fd1713fea395a4bd0ebb97c3d34a8211e9f1dda775d989a395e8dcd7;
    5'b10101 : xpb = 1024'h9b85e2f92de88f22007f3915979821df8f937e5342ed3e8bce58de7910c33c97e46866a0f5bf0a9f859fbd40d666bcb93aa8c8704da8b8c2bad36c5d87112db564e1d5c6bd50b6d5ca8fc03fca23363b7824d93659e895bb51ac19a78eb9fb9509e779678aa993e0999382ce5b0a98470348839b28161050acb522f93ebcdda5;
    5'b10110 : xpb = 1024'hb7dd6ec4cea8115fd2b42cbfe82c1c8f8355d08cc1819816019d04dc1442512296c30bafed7e7cb58b8161f8b7055cb6dbef8ed582fde41fb91f21136822d62e16bbefd852d9d4f6eee0418fb688475dd77ac17b4fa8e9d892f9dc03f183312a51cc4f367731b3508d17a00af8972a0e46ca64215eee5c99d21414a5eae7808;
    5'b10111 : xpb = 1024'h2c2310352ddaa7d2c4dcc45975c7a903d24d3eef2aba94ee6fb77b7824c7ba9471b8784dd2174385cb2eae4523d7ffa804ef51508569d40cecefb72320c5a1c1d244dce2fc9b810e25e64a94c58996e136cf78919c92b490763fb3d3a9a10d226f59a2a8f5059b16fecf5811fbd87324146aa7cb54131872d3fcdaa0078278d6;
    5'b11000 : xpb = 1024'h4cc8497e0ecace8f8c8e45e6ed0c903eac6520d5895d105b7f5526a2884b5016ba04bfe0a5569f403da5466abc3fa9849c1fa9b3b2a3c9d7de4d7c350b091620c31dfac8740964ccdcde91108faaa94c9027450b842ada83634fc9e71429e7323996805e82981af8f4cd3623482773a74468a95492374b1c0ad873f5b05679a4;
    5'b11001 : xpb = 1024'h6d6d82c6efbaf54c543fc77464517779867d02bbe7ff8bc88ef2d1ccebcee599025107737895fafab01bde9054a7536133500216dfddbfa2cfab4146f54c8a7fb3f718adeb77488b93d6d78c59cbbbb7e97f11856bc30076505fdffa7eb2c14203d35e14102a9adaeacb14349476742a7466aaddd05b7dc541b40d4b592a7a72;
    5'b11010 : xpb = 1024'h8e12bc0fd0ab1c091bf14901db965eb46094e4a246a207359e907cf74f527b1b4a9d4f064bd556b5229276b5ed0efd3dca805a7a0d17b56dc1090658df8ffedea4d0369362e52c4a4acf1e0823ecce2342d6ddff535b26693d6ff60de93b9b51ce103bc99dbd1abce0c8f245e0c574ada464ac670e7fb06e788fa6a101fe7b40;
    5'b11011 : xpb = 1024'haeb7f558b19b42c5e3a2ca8f52db45ef3aacc688a54482a2ae2e2821b2d6109d92e996991f14b26f95090edb8576a71a61b0b2dd3a51ab38b266cb6ac9d3733d95a95478da53100901c76483ee0de08e9c2eaa793af34c5c2a800c2153c47561984d197f2b4f9a9ed6c6d0572d147530d462adf04ca3e317af6b3ff6aad27c0e;
    5'b11100 : xpb = 1024'h1eafe94bd09d34b9e04ed445b9c5e5d8a34ea53e2e6f5d983fef19f66356f917d7ed60b3282d8f9b682167ba3a80402c94c6e35a44d8d0b7f325511e794472eb12333dafa22ff682a625a85d1f532ec901817d5a9605453e6203903a0422acdf3382650b081921f34604c78981934f8ab586d0973a7cb8909fd75e47cac41671;
    5'b11101 : xpb = 1024'h3f552294b18d5b76a80055d3310acd137d6687248d11d9054f8cc520c6da8e9a2039a845fb6ceb55da97ffdfd2e7ea092bf73bbd7212c682e48316306387e74a030c5b95199dda415d1deed8e97441345ad949d47d9d6b314f13a64d6eab86eefdbf42c095aba1d53c02a59acde2500de584d22078a0eb39d6b2f79d7398173f;
    5'b11110 : xpb = 1024'h5ffa5bdd927d82336fb1d760a84fb44e577e690aebb454725f2a704b2a5e241c6885efd8ceac47104d0e98056b4f93e5c32794209f4cbc4dd5e0db424dcb5ba8f3e5797a910bbe0014163554b395539fb431164e653591243c23bc60d93460fec7fc2076233e21b7320083ac1a3150911582d3a9b6c51de30d8e90f31c6c180d;
    5'b11111 : xpb = 1024'h809f9526736da8f0376358ee1f949b8931964af14a56cfdf6ec81b758de1b99eb0d2376ba1eba2cabf85302b03b73dc25a57ec83cc86b218c73ea054380ed007e4be97600879a1becb0e7bd07db6660b0d88e2c84ccdb7172933d27443bd3b0e9238fe2bb0d0a19927fe61bd668051144580d532f4e9508c446a2a48c54018db;
    endcase
end

endmodule

module xpb_5_675
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h7a7c49753c5b457ff1d14e7046f83841d4d1e140c5b7522d8f04acc43e2df3a19484387fa19471dfe1248041e913e8da098b7e315144bee260f869b957c2cbdcf77d3d27446f1d3d7281a403a7681f75028e29fcafd9002b1439250cfb519694fea71b6a55f6bee05c53dda9d4c192407fb5b947e124f1a67a23815dcb624670;
    5'b00010 : xpb = 1024'h444b4d94b6c85637189d25097d962932382dbf50b5f703e3a02ca032c9593a3b25bff3867902653122eac13ceec9c0e9aefcd47c7fd6ad791151941474b323087aab459fd94d3d35d2694564b5f47ab911175a60d32bd34572e5b81f3c788a97ce46a4aafb24853331e7d474b1b2fe57b09193ad71fe861cadd787b70de22675;
    5'b00011 : xpb = 1024'he1a51b4313566ee3f68fba2b4341a229b899d60a636b599b15493a1548480d4b6fbae8d5070588264b10237f47f98f9546e2ac7ae689c0fc1aabe6f91a37a33fdd94e186e2b5d2e3250e6c5c480d5fd1fa08ac4f67ea65fd1924b317d9f7e9a9de62deba0524b86077bcb3f8ea46a6ee16d6e1302d81a92e18b8e105062067a;
    5'b00100 : xpb = 1024'h88969b296d90ac6e313a4a12fb2c5264705b7ea16bee07c74059406592b274764b7fe70cf204ca6245d58279dd9381d35df9a8f8ffad5af222a32828e9664610f5568b3fb29a7a6ba4d28ac96be8f572222eb4c1a657a68ae5cb703e78f1152f9c8d4955f6490a6663cfa8e96365fcaf6123275ae3fd0c395baf0f6e1bc44cea;
    5'b00101 : xpb = 1024'h52659f48e7fdbd25580620ac31ca4354d3b75cb15c2db97d518133d41dddbb0fdcbba213c972bdb3879bc374e34959e3036aff442e3f4988d2fc528406569d3c788493b847789a6404ba2c2a7a7550b630b7e525c9aa79a544780350ba1809326c2cd2969b76d0b939639fb4405768c691ff01c074d6a0af8f6315c75e442cef;
    5'b00110 : xpb = 1024'h1c34a368626acddc7ed1f7456868344537133ac14c6d6b3362a92742a90901a96df75d1aa0e0b104c962046fe8ff31f2a8dc558f5cd1381f83557cdf2346f467fbb29c30dc56ba5c64a1cd8b8901abfa3f411589ecfd4cbfa3249662fb3efd353bcc5bd740a4970c0ef7967f1d48d4ddc2dadc2605b03525c3171c20a0c40cf4;
    5'b00111 : xpb = 1024'h96b0ecdd9ec6135c70a345b5af606c870be51c021224bd60f1add406e736f54b027b959a427522e4aa8684b1d2131accb267d3c0ae15f701e44de6987b09c044f32fd95820c5d799d723718f3069cb6f41cf3f869cd64ceab75dbb6ff69093ca3a737741969b55ec6b4b7428f20a671e4290956de6d526cc3d3a9d7e6c265364;
    5'b01000 : xpb = 1024'h607ff0fd19332413976f1c4ee5fe5d776f40fa1202646f1702d5c77572623be493b750a119e31635ec4cc5acd7c8f2dc57d92a0bdca7e59894a710f397fa1770765de1d0b5a3f792370b12f03ef626b350586feac0292005160a4e8237b787cd0a1300823bc91c3f40df6af3cefbd335736c6fd377aebb4270eea3d7aea63369;
    5'b01001 : xpb = 1024'h2a4ef51c93a034cabe3af2e81c9c4e67d29cd821f2a420cd13fdbae3fd8d827e24f30ba7f15109872e1306a7dd7ecaebfd4a80570b39d42f45003b4eb4ea6e9bf98bea494a82178a96f2b4514d8281f75ee1a04ee37bf31f74b6e19478de7bcfd9b289c2e0f6e292167361beabed3f4ca4484a3908884fb8a4a2aa30f126136e;
    5'b01010 : xpb = 1024'ha4cb3e91cffb7a4ab00c4158639486a9a76eb962b85b72faa30267a83bbb761fb977442792e57b670f3786e9c692b3c606d5fe885c7e9311a5f8a5080cad3a78f10927708ef134c809745854f4eaa16c616fca4b9354f34a88f006a174301264d859a52d36eda17272c73f6880aed18d23fe0380e9ad415f1ec62b8ebc8859de;
    5'b01011 : xpb = 1024'h6e9a42b14a688b01d6d817f19a32779a0aca9772a89b24b0b42a5b16c6e6bcb94ab2ff2e6a536eb850fdc7e4cc488bd5ac4754d38b1081a85651cf63299d91a474372fe923cf54c0695bf9b60376fcb06ff8faafb6a7c664e79c99b3b5570667a7f92e6ddc1b67c5485b36335da03da454d9dde67a86d5d5527a31e7ff0839e3;
    5'b01100 : xpb = 1024'h386946d0c4d59bb8fda3ee8ad0d0688a6e26758298dad666c5524e8552120352dbeeba3541c1620992c408dfd1fe63e551b8ab1eb9a2703f06aaf9be468de8cff7653861b8ad74b8c9439b17120357f47e822b13d9fa997f46492cc5f67dfa6a7798b7ae81492e181def2cfe3a91a9bb85b5b84c0b606a4b862e3841418819e8;
    5'b01101 : xpb = 1024'h2384af03f42ac70246fc524076e597ad1825392891a881cd67a41f3dd3d49ec6d2a753c192f555ad48a49dad7b43bf4f72a0169e8345ed5b7042419637e3ffb7a9340da4d8b94b1292b3c78208fb3388d0b5b77fd4d6c99a4f5bfd837a4ee6d473840ef2676f46af38323c9178315d2b69192b19c39fec1b9e23e9a8407f9ed;
    5'b01110 : xpb = 1024'h7cb494657b9df1f0164113944e6691bca65434d34ed1da4a657eeeb81b6b3d8e01aeadbbbac3c73ab5aeca1cc0c824cf00b57f9b39791db817fc8dd2bb410bd872107e0191fab1ee9bace07bc7f7d2ad8f998574ad266cc4b92ee4e532f6850245df5c597c6db34b4fd70172ec44a81336474bf97d5ef0683405bff84f6a405d;
    5'b01111 : xpb = 1024'h46839884f60b02a73d0cea2d850482ad09b012e33f118c0076a6e226a696842792ea68c29231ba8bf7750b17c67dfcdea626d5e6680b0c4ec855b82dd8316303f53e867a26d8d1e6fb9481dcd6842df19e22b5d8d0793fdf17db77f7741d7905157ee59a219b799e256af83dc936142a6723265f0e3884de67b9c65191ea2062;
    5'b10000 : xpb = 1024'h10529ca47078135e63d8c0c6bba2739d6d0bf0f32f513db687ced59531c1cac1242623c9699faddd393b4c12cc33d4ee4b982c31969cfae578aee288f521ba2f786c8ef2bbb6f1df5b7c233de5108935acabe63cf3cc12f976880b09b5446d07e51e6edac6c93ff0fafeef08a627804197ff00c49f1219549b6dccaad46a0067;
    5'b10001 : xpb = 1024'h8acee619acd358de55aa0f37029aabdf41ddd233f5088fe416d382596fefbe62b8aa5c490b341fbd1a5fcc54b547bdc85523aa62e7e1b9c7d9a74c424ce4860c6fe9cc1a00260f1ccdfdc7418c78a8aaaf3a1039a3a513248ac13016b096039ce3c58a451cbffed15752ccb27ae9128217b4ba0c80370afb15914e089fcc46d7;
    5'b10010 : xpb = 1024'h549dea39274069957c75e5d039389ccfa539b043e548419a27fb75c7fb1b04fc49e6174fe2a2130e5c260d4fbafd95d7fa9500ae1673a85e8a00769d69d4dd37f317d49295042f152de568a29b0503eebdc3409dc6f7e63ee96dc328f1bcf79fb3651385c1edc5242ce6c37d57da7e994890947211109f7149455461e24c26dc;
    5'b10011 : xpb = 1024'h1e6cee58a1ad7a4ca341bc696fd68dc008958e53d587f3503923693686464b95db21d256ba10065f9dec4e4ac0b36de7a00656f9450596f53a59a0f886c534637645dd0b29e24f0d8dcd0a03a9915f32cc4c7101ea4ab959481a563b32e3eba283049cc6671b8b77027aba4834cbeab0796c6ed7a1ea33e77cf95abb24cc06e1;
    5'b10100 : xpb = 1024'h98e937cdde08bfcc95130ad9b6cec601dd676f949b3f457dc82815fac4743f376fa60ad65ba4783f7f10ce8ca9c756c1a991d52a964a55d79b520ab1de8800406dc31a326e516c4b004eae0750f97ea7ceda9afe9a23b9845c537b482e35823781abb830bd124a575ece97f2098d7cf0f922281f830f258df71cdc18f02e4d51;
    5'b10101 : xpb = 1024'h62b83bed5875d083bbdee172ed6cb6f240c34da48b7ef733d95009694f9f85d100e1c5dd33126b90c0d70f87af7d2ed14f032b75c4dc446e4bab350cfb78576bf0f122ab032f8c4360364f685f85d9ebdd63cb62bd768c9ebb000e5a6f5c763a514b4171624010aa34628ebce67ee90829fe028513e8ba042ad0e27232ae2d56;
    5'b10110 : xpb = 1024'h2c87400cd2e2e13ae2aab80c240aa7e2a41f2bb47bbea8e9ea77fcd7dacacc6a921d80e40a805ee2029d5082b53306e0f47481c0f36e3304fc045f681868ae97741f2b23980dac3bc01df0c96e12352febecfbc6e0c95fb919aca16cb0836a3d20eacab2076dd6fd09f68587c370551f5ad9dceaa4c24e7a5e84e8cb752e0d5b;
    5'b10111 : xpb = 1024'ha70389820f3e26bad47c067c6b02e02478f10cf54175fb17797ca99c18f8c00c26a1b963ac14d0c1e3c1d0c49e46efbafdfffff244b2f1e75cfcc921702b7a746b9c684adc7cc979329f94cd157a54a4ee7b25c390a25fe42de5c679abd500d21f91e61c5d6495dd664a63319831e75fda8f963285e74020d8a86a29409053cb;
    5'b11000 : xpb = 1024'h70d28da189ab3771fb47dd15a1a0d114dc4ceb0531b5accd8aa49d0aa42406a5b7dd746a8382c413258811bfa3fcc7caa371563d7344e07e0d55f37c8d1bd19feeca70c3715ae9719287362e2406afe8fd045627b3f532fe8c92598becfbf4d4ef316f5d02925c303bde59fc752353770b6b709816c0d4970c5c7082831033d0;
    5'b11001 : xpb = 1024'h3aa191c1041848292213b3aed83ec2053fa8c91521f55e839bcc90792f4f4d3f49192f715af0b764674e52baa9b29fda48e2ac88a1d6cf14bdaf1dd7aa0c28cb71f8793c06390969f26ed78f32930b2d0b8d868bd7480618eb3eec9e2e22e8d7bed0f89da7c02283117250c75214bf8e3c474afda79a690d401076dbc59013d5;
    5'b11010 : xpb = 1024'h47095e07e8558e048df8a480edcb2f5a304a72512351039acf483e7ba7a93d8da54ea78325eaab5a91493b5af6877e9ee5402d3d068bdab6e084832c6fc7ff6f52681b49b172962525678f0411f66711a16b6effa9ad93349eb7fb06f49dcda8e7081de4cede8d5e70647922f062ba56d2325633873fd8373c47d35080ff3da;
    5'b11011 : xpb = 1024'h7eecdf55bae09e603ab0d8b855d4eb3777d68865d7ec62673bf930abf8a8877a6ed922f7d3f31c958a3913f7987c60c3f7df810521ad7c8dcf00b1ec1ebf4bd3eca3bedbdf86469fc4d81cf3e88785e61ca4e0ecaa73d95e5e24a4bd6a9b736f8d179d48a2e4a7b6435a253c03c7bde5ecd8deab1998ef29ede7fe92d3723a4a;
    5'b11100 : xpb = 1024'h48bbe375354daf17617caf518c72dc27db326675c82c141d4d21241a83d3ce140014ddfeab610fe6cbff54f29e3238d39d50d750503f6b247f59dc473bafa2ff6fd1c7547464669824bfbe54f713e12a2b2e1150cdc6ac78bcd137cfabc267725cb7268948126e0918ee1c06e0b929fd1db4b910aa7283a0219c04ec15f21a4f;
    5'b11101 : xpb = 1024'h128ae794afbabfce884885eac310cd183e8e4485b86bc5d35e4917890eff14ad9150990582cf03380dc595eda3e810e342c22d9b7ed159bb2fb306a2589ffa2af2ffcfcd0942869084a75fb605a03c6e39b741b4f1197f931b7dcae1ece95b752c56afc9ed40345bee8212d1bdaa96144e9093763b4c181655500b455871fa54;
    5'b11110 : xpb = 1024'h8d073109ec16054e7a19d45b0a09055a136025c67e231800ed4dc44d4d2d084f25d4d18524637517eeea162f8cfbf9bd4c4dabccd016189d90ab705bb062c607ea7d0cf44db1a3cdf72903b9ad085be33c456bb1a0f27fbe2fb6efeee83af20a2afdcb344336f33c4ad5f07b926c2854ce464cbe1c7109bccf738ca323d440c4;
    5'b11111 : xpb = 1024'h56d6352966831605a0e5aaf440a6f64a76bc03d66e62c9b6fe75b7bbd8584ee8b7108c8bfbd1686930b0572a92b1d1ccf1bf0217fea8073441049ab6cd531d336dab156ce28fc3c65710a51abb94b7274ace9c15c44552d88e6383012961e60cfa9d5474e864b98f2069e7466f5d946bff222723ad4a9e33032792fc665420c9;
    endcase
end

endmodule

module xpb_5_415
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h4da6f10d9313d2e3bcf2395c1f3ce89e132b3ea75ab846109977a53a051b008c0253b0f3a1735ad8f1d949473a082b4839bfdff17204b622a93179cfb9f3e768bb2ba5909b95b2e98147e275df3254a49b7a3d16722c0fc623492501bceeb96e6ea1992577e75bf53893626ac9a6d64a82e4c0de098a259ed362250c3c960471;
    5'b00010 : xpb = 1024'h9b4de21b2627a5c779e472b83e79d13c26567d4eb5708c2132ef4a740a36011804a761e742e6b5b1e3b2928e74105690737fbfe2e4096c455262f39f73e7ced176574b21372b65d3028fc4ebbe64a94936f47a2ce4581f8c46924a0379dd72dcdd43324aefceb7ea7126c4d5934dac9505c981bc13144b3da6c44a18792c08e2;
    5'b00011 : xpb = 1024'h38478dd2f74d43e26bd1343d4d5c7288c80bb8c53ab131ba4e8a36585c4e549c03b295621a3391fc362d9c8ecaba710e492577ee335b521c4af52e10f3094188bd33bc0323301b77713da4bf04bb39bcde69bdaac9fe0241b44edd0a7ca189b91cdd3946b6ed1b5222fa406165245cb639d463b7cc5313ac33b6f4202cdfa6e8;
    5'b00100 : xpb = 1024'h85ee7ee08a6116c628c36d996c995b26db36f76c956977cae801db926169552806064655bba6ecd52806e5d604c29c5682e557dfa560083ef426a7e0acfd28f1785f6193bec5ce60f2858734e3ed8e6179e3fac13c2a1207d798020c399043278b7ed26c2ed477475b8da2cc2ecb3300bcb92495d5dd394b0719192c6975ab59;
    5'b00101 : xpb = 1024'h22e82a985b86b4e11ab02f1e7b7bfc737cec32e31aaa1d64039cc776b381a8ac051179d092f3c91f7a81efd65b6cb6d4588b0feaf4b1ee15ecb8e2522c1e9ba8bf3bd275aaca8405613367082a441ed521593e3f21cff4bd455495133c545a03cb18d967f5f2daaf0d611e5800a1e321f0c406918f1c01b9940bc3341d29495f;
    5'b00110 : xpb = 1024'h708f1ba5ee9a87c4d7a2687a9ab8e5119017718a756263749d146cb0b89ca93807652ac4346723f86c5b391d9574e21c924aefdc66b6a43895ea5c21e61283117a677806466036eee27b497e09767379bcd37b5593fc0483689dba14f943137239ba728d6dda36a445f480c2ca48b96c73a8c76f98a62758676de84059bf4dd0;
    5'b00111 : xpb = 1024'hd88c75dbfc025dfc98f29ffa99b865e31ccad00faa3090db8af58950ab4fcbc06705e3f0bb40042bed6431dec1efc9a67f0a7e7b6088a0f8e7c96936533f5c8c143e8e83264ec93512929514fcd03ed6448bed379a1e738d65a4d1bfc072a4e7954798934f89a0bf7c7fc4e9c1f698da7b3a96b51e4efc6f46092480d72ebd6;
    5'b01000 : xpb = 1024'h5b2fb86b52d3f8c38681635bc8d86efc44f7eba8555b4f1e5226fdcf0fcffd4808c40f32ad275b1bb0af8c65262727e2a1b087d9280d403237ae10631f27dd317c6f8e78cdfa9f7cd2710bc72eff5891ffc2fbe9ebcdf6fef9a3721db8f5e3bce7f612aeacdff601305b5eb965c63fd82a986a495b6f1565c7c2b7544a08f047;
    5'b01001 : xpb = 1024'ha8d6a978e5e7cba743739cb7e815579a58232a4fb013952eeb9ea30914eafdd40b17c0264e9ab5f4a288d5ac602f532adb7067ca9a11f654e0df8a32d91bc49a379b34096990526653b8ee3d0e31ad369b3d39005dfa06c51cec971f75e49d2b5697abd424c751f668eec1242f6d1622ad7d2b2764f93b049b24dc60869ef4b8;
    5'b01010 : xpb = 1024'h45d05530b70d69c235605e3cf6f7f8e6f9d865c635543ac807398eed670351580a22f3a125e7923ef503dfacb6d96da8b1161fd5e963dc2bd971c4a4583d37517e77a4eb5595080ac266ce1054883daa42b27c7e439fe97a8aa92a2678a8b4079631b2cfebe5b55e1ac23cb00143c643e1880d231e380373281786683a5292be;
    5'b01011 : xpb = 1024'h9377463e4a213ca5f25297991634e1850d03a46d900c80d8a0b134276c1e51e40c76a494c75aed17e6dd28f3f0e198f0ead5ffc75b68924e82a33e7412311eba39a34a7bf12abaf443aeb08633ba924ede2cb994b5cbf940adf24f2835976d7604d34bf563cd115353559f1acaea9c8e646cce0127c22911fb79ab7476e8972f;
    5'b01100 : xpb = 1024'h3070f1f61b46dac0e43f591e251782d1aeb8dfe4154d2671bc4c200bbe36a5680b81d80f9ea7c962395832f4478bb36ec07bb7d2aaba78257b3578e591529171807fbb5ddd2f7098b25c90597a1122c285a1fd129b71dbf61baee22f385b8452446d52f12aeb74bb05291aa69cc14caf9877affce100f180886c557c2a9c3535;
    5'b01101 : xpb = 1024'h7e17e303ae5aada4a131927a44546b6fc1e41e8b70056c8255c3c545c351a5f40dd58903401b243b2b317c3b8193deb6fa3b97c41cbf2e482466f2b54b4678da3bab60ee78c5238233a472cf59437767211c3a290d9debbc3ef80730f54a3dc0b30eec16a2d2d0b03dbc7d11666822fa1b5c70daea8b171f5bce7a88673239a6;
    5'b01110 : xpb = 1024'h1b118ebb7f804bbf931e53ff53370cbc63995a01f546121b715eb12a1569f9780ce0bc7e176800857dac863bd83df934cfe14fcf6c11141f1cf92d26ca67eb918287d1d064c9d926a25252a29f9a07dac8917da6f343ce71acb49a37f80e549cf2a8f31269f13417ef8ff89d383ed31b4f6752d6a3c9df8de8c124901ae5d7ac;
    5'b01111 : xpb = 1024'h68b87fc912941ea350108d5b7273f55a76c498a94ffe582c0ad656641a84fa040f346d71b8db5b5e6f85cf831246247d09a12fc0de15ca41c62aa6f6845bd2fa3db37761005f8c10239a35187ecc5c7f640bbabd656fde37cffdbf39b4fd0e0b614a8c37e1d8900d28235b0801e5a965d24c13b4ad54052cbc23499c577bdc1d;
    5'b10000 : xpb = 1024'h5b22b80e3b9bcbe41fd4ee0815696a71879d41fd53efdc5267142486c9d4d880e3fa0ec902837a8c200d98368f03efadf46e7cc2d67b018bebce168037d45b1848fe842ec6441b4924814ebc522ecf30b80fe3b4b15c0ed3dba5240b7c124e7a0e49333a8f6f374d9f6d693d3bc59870656f5b06692cd9b4915f3a40b2f7a23;
    5'b10001 : xpb = 1024'h53591c8e76cd8fa1feef883ca0937f452ba512c72ff743d5bfe8e78271b84e14109351e0319b9281b3da22caa2f86a431906c7bd9f6c663b67ee5b37bd712d1a3fbb8dd387f9f49e138ff761a4554197a6fb3b51bd41d0b36103774274afde560f862c5920de4f6a128a38fe9d632fd1893bb68e701cf33a1c7818b047c57e94;
    5'b10010 : xpb = 1024'ha1000d9c09e16285bbe1c198bfd067e33ed0516e8aaf89e659608cbc76d34ea012e702d3d30eed5aa5b36c11dd00958b52c6a7af11711c5e111fd50777651482fae73364238fa78794d7d9d78387963c427578682f6de079844c9c44319e97c47e27c57e98c5ab5f4b1d9b69670a061c0c20776c79a718d8efda3dbc845b8305;
    5'b10011 : xpb = 1024'h3df9b953db0700a0adce831dceb3092fe0858ce50ff02f7f74fb78a0c8eba22411f2364eaa5bc9a4f82e761233aab009286c5fba60c3023509b20f78f686873a41c3a4460f945d2c0385b9aac9de26afe9eabbe61513c32ef2092f4b3462aea0bdc1cc7a5fe40ec6fcf116f538e0b63d402b596832e5e1477ccce7c4380f210b;
    5'b10100 : xpb = 1024'h8ba0aa616e1ad3846ac0bc79edeff1cdf3b0cb8c6aa875900e731ddace06a2b01445e7424bcf247dea07bf596db2db51622c3fabd2c7b857b2e38948b07a6ea2fcef49d6ab2a101584cd9c20a9107b548564f8fc873fd2f51552544cf151680f2c63659fd7cb6abc3584796002878c87c3101a463c7006e6502f0cd074a5257c;
    5'b10101 : xpb = 1024'h289a56193f40719f5cad7dfefcd2931a95660702efe91b292a0e09bf201ef63413511abd231c00c83c82c959c45cf5cf37d1f7b722199e2eab75c3ba2f9be15a43cbbab8972ec5b9f37b7bf3ef670bc82cda3c7a6ce5b5aa830ee753f4157eeb6bfd6c9b9ee9ce23e757f4ebd45e3ca8f71afc41f5aecf54dd21b6d82858c382;
    5'b10110 : xpb = 1024'h76414726d2544483199fb75b1c0f7bb8a89145aa4aa16139c385aef92539f6c015a4cbb0c48f5ba12e5c12a0fe6521177191d7a8941e545154a73d89e98fc8c2fef7604932c478a374c35e69ce99606cc8547990df11c570a6580c55b1043859da9f05c116d12a191feb57569e0512f379ffbd1fff38f4f3b083dbe464eec7f3;
    5'b10111 : xpb = 1024'h133af2dea379e29e0b8c78e02af21d054a468120cfe206d2df209add77524a4414afff2b9bdc37eb80d71ca1550f3b9547378fb3e3703a284d3977fb68b13b7a45d3d12b1ec92e47e3713e3d14eff0e06fc9bd0ec4b7a82614149f5cb3c84f361a390cbcddef8d80d1bed2e26fdbc314ae0a9f1bb877bd623d7685ec18a265f9;
    5'b11000 : xpb = 1024'h60e1e3ec368db581c87eb23c4a2f05a35d71bfc82a9a4ce3789840177c6d4ad01703b01f3d4f92c472b065e88f1766dd80f76fa55574f04af66af1cb22a522e300ff76bbba5ee13164b920b2f42245850b43fa2536e3b7ec375dc45e70b708a488daa5e255d6e9760a52354d3982995f30ef5ff9c201e30110d8aaf855386a6a;
    5'b11001 : xpb = 1024'hae88d4f9c9a188658570eb98696bee41709cfe6f855292f4120fe55181884b5c19576112dec2ed9d6489af2fc91f9225bab74f96c779a66d9f9c6b9adc990a4bbc2b1c4c55f4941ae6010328d3549a29a6be373ba90fc7b25aa6e9602da5c212f77c3f07cdbe456b42e597b803296fa9b3d420d7cb8c089fe43ad00491ce6edb;
    5'b11010 : xpb = 1024'h4b8280b19ac72680775dad1d784e8f8e125239e60a93388d2daad135d3a09ee01862948db60fc9e7b704b9301fc9aca3905d07a216cb8c44982ea60c5bba7d0303078d2e41f949bf54aee2fc19ab2a9d4e337ab98eb5aa67c8637c673069d8ef3716460394dca8d2f4b91343d5001fcae7df02d384cad10e712d7a0c45820ce1;
    5'b11011 : xpb = 1024'h992971bf2ddaf964344fe679978b782c257d788d654b7e9dc722766fd8bb9f6c1ab64581578324c0a8de027759d1d7ebca1ce79388d0426741601fdc15ae646bbe3332bedd8efca8d5f6c571f8dd7f41e9adb7d000e1ba2debaca168ed58925da5b7df290cc404c82d4c75ae9ea6f6156ac3c3b18e54f6ad448f9f1882181152;
    5'b11100 : xpb = 1024'h36231d76ff00977f263ca7fea66e1978c732b403ea8c2436e2bd62542ad3f2f019c178fc2ed0010afb590c77b07bf2699fc29f9ed822283e39f25a4d94cfd723050fa3a0c993b24d44a4a5453f340fb59122fb4de6879ce35969346ff01ca939e551e624d3e2682fdf1ff13a707da6369ecea5ad4793bf1bd182492035cbaf58;
    5'b11101 : xpb = 1024'h83ca0e8492146a62e32ee15ac5ab0216da5df2ab45446a477c35078e2feef37c1c1529efd0435be3ed3255beea841db1d9827f904a26de60e323d41d4ec3be8bc03b493165296536c5ec87bb1e66645a2c9d386458b3aca97cb25971ad0b62a853f37f4a4bc9c42517b353a53a247c8121b3668b511de4baa4e46e2c7261b3c9;
    5'b11110 : xpb = 1024'h20c3ba3c633a087dd51ba2dfd48da3637c132e21ca850fe097cff372820747001b205d6aa790382e3fad5fbf412e382faf28379b9978c437dbb60e8ecde531430717ba13512e1adb349a678e64bcf4cdd4127be23e598f5eea6eec78afcf7984938d864612e8278cc986cf310bfb2ca255be48870a5cad2931d71834261551cf;
    5'b11111 : xpb = 1024'h6e6aab49f64ddb61920ddc3bf3ca8c018f3e6cc9253d55f1314798ac8722478c1d740e5e490393073186a9067b366377e8e8178d0b7d7a5a84e7885e87d918abc2435fa3ecc3cdc4b5e24a0443ef49726f8cb8f8b0859f250db8117a6cbe32f3022f1f6b8acf8382021a319bd5a202ecd8a3096513e6d2c805393d4062ab5640;
    endcase
end

endmodule

module xpb_5_595
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h4a8c537924508ce3a4987205568d5a11c163cb3dbc84c3a9e16291c478d919bed62b6a7865209f4a43a04e4e21be90f1437ecf85f60905346966f593fd0db50c2a16afeee04fa17c3086277b6d475ee2d5231e8ddcea9a26dca3b6759f0d41bc1b1244901a08829e030448ee4767e089c7cd35594e027697ad47f5baa1efc905;
    5'b00010 : xpb = 1024'h9518a6f248a119c74930e40aad1ab42382c7967b79098753c2c52388f1b2337dac56d4f0ca413e9487409c9c437d21e286fd9f0bec120a68d2cdeb27fa1b6a18542d5fddc09f42f8610c4ef6da8ebdc5aa463d1bb9d5344db9476ceb3e1a8378362489203411053c060891dc8ecfc1138f9a6ab29c04ed2f5a8feb7543df920a;
    5'b00011 : xpb = 1024'h2ef7b515ab0371e222c3de38f34dc6e3d2b55e886016aa86264afbf7b788a0347f39c1f0653b5f502b82aba381dda209666246abbf683f518b95a15dbc56aa7309f4db1df15de72f7ef873cfaefa58778b6462110a39a163e05e916622fd22a2222f3b869d508f4c824cf3ebde677b74088dc12999bc0696c168662b5cecf4a4;
    5'b00100 : xpb = 1024'h7984088ecf53fec5c75c503e49db20f5941929c61c9b6e3007ad8dbc3061b9f355652c68ca5bfe9a6f22f9f1a39c32faa9e11631b5714485f4fc96f1b9645f7f340b8b0cd1ad88abaf7e9b4b1c41b75a6087809ee7243b8abd0247dbc20a645e3d418016b75911ea85513cda25cf5bfdd05af682e7be7d2e6eb05be5fedcbda9;
    5'b00101 : xpb = 1024'h136316b231b656e0a0ef4a6c900e33b5e406f1d303a891626b33662af63826aa2848196865561f56136508f8e1fcb3218945bdd188c7796eadc44d277b9f9fd9e9d3064d026c2ce2cd6ac023f0ad520c41a5a5943788a8a0e4196c56a6ed0388294c327d20989bfb01959ee97567165e494e4cf9e5759695d588d69c17ea2043;
    5'b00110 : xpb = 1024'h5def6a2b5606e3c44587bc71e69b8dc7a56abd10c02d550c4c95f7ef6f114068fe7383e0ca76bea05705574703bb4412ccc48d577ed07ea3172b42bb78ad54e613e9b63be2bbce5efdf0e79f5df4b0ef16c8c422147342c7c0bd22cc45fa4544445e770d3aa11e990499e7d7bccef6e8111b825333780d2d82d0cc56b9d9e948;
    5'b00111 : xpb = 1024'ha87bbda47a5770a7ea202e773d28e7d966ce884e7cb218b62df889b3e7ea5a27d49eee592f975dea9aa5a5952579d50410435cdd74d983d78092384f75bb09f23e00662ac30b6fdb2e770f1acb3c0fd1ebebe2aff15ddcee9d60d941e50787005f70bb9d54a9a137079e30c60436d771d8e8b7ac817a83c53018c2115bc9b24d;
    5'b01000 : xpb = 1024'h425acbc7dcb9c8c2c3b328a5835bfa99b6bc505b63bf3be8917e6222adc0c6dea781db58ca917ea63ee7b49c63da552aefa8047d482fb8c03959ee8537f64a4cf3c7e16af3ca14124c6333f39fa7aa83cd0a07a541c24a04c477fdbcc9ea262a4b7b6e03bde92b4783e292d553ce91d251dc0e237f319d2c96f13cc774d714e7;
    5'b01001 : xpb = 1024'h8ce71f41010a55a6684b9aaad9e954ab78201b992043ff9272e0f3e72699e09d7dad45d12fb21df0828802ea8598e61c3326d4033e38bdf4a2c0e4193503ff591dde9159d419b58e7ce95b6f0cef0966a22d26331eace42ba11bb43268f767e6668db293d7f1ade586e6dbc39b36725c19a9437ccd3413c44439328216c6ddec;
    5'b01010 : xpb = 1024'h26c62d64636cadc141de94d9201c676bc80de3a6075122c4d666cc55ec704d54509032d0caac3eac26ca11f1c3f96643128b7ba3118ef2dd5b889a4ef73f3fb3d3a60c9a04d859c59ad58047e15aa418834b4b286f115141c832d8ad4dda0710529864fa413137f6032b3dd2eace2cbc929c99f3caeb2d2bab11ad382fd44086;
    5'b01011 : xpb = 1024'h715280dd87bd3aa4e67706de76a9c17d8971aee3c3d5e66eb7c95e1a6549671326bb9d492fccddf66a6a603fe5b7f734560a4b290797f811c4ef8fe2f44cf4bffdbcbc88e527fb41cb5ba7c34ea202fb586e69b64bfbeb68a4d68f22ece748cc6daaa98a5b39ba94062f86c132360d465a69cf4d18eda3c35859a2f2d1c4098b;
    5'b01100 : xpb = 1024'hb318f00ea1f92bfc00a010cbcdcd43dd95f76f0aae309a11b4f36892b1fd3c9f99e8a48cac6feb20eac6f472418775b356ef2c8daee2cfa7db74618b688351ab38437c915e69f78e947cc9c230d9dad398c8eab9c60587ecbedb39dd1c9e7f659b55bf0c47944a48273e8d081cdc7a6d35d25c416a4bd2abf321da8ead16c25;
    5'b01101 : xpb = 1024'h55bde27a0e701fa364a27312136a2e4f9ac3422e6767cd4afcb1c84da3f8ed88cfc9f4c12fe79dfc524cbd9545d7084c78edc24ed0f7322ee71e3bacb395ea26dd9ae7b7f63640f519cdf4179054fc900eafad39794af2a5a8916a1370d729b274c7a080de81c742857831bec935a8309b2a5b1d64a733c26c7a13638cc1352a;
    5'b01110 : xpb = 1024'ha04a35f332c0ac87093ae51769f788615c270d6c23ec90f4de145a121cd20747a5f55f3995083d4695ed0be36795993dbc6c91d4c700376350853140b0a39f3307b197a6d685e2714a541b92fd9c5b72e3d2cbc756358ccc853520890fe46b6e8fd9e510f88a49e0887c7aad109d88ba62f79076b2a9aa5a19c2091e2eb0fe2f;
    5'b01111 : xpb = 1024'h3a294416952304a1e2cddf45b02a9b21ac14d5790af9b427419a3280e2a873fe78d84c3930025e023a2f1aeaa5f619649bd139749a566c4c094ce77672dedf8dbd7912e7074486a86840406bd207f624c4f0f0bca699f9e2ac4c4503f4c70a987be4977761c9d3f104c0dcbc6035431adbeae6edb060c3c1809a83d447be60c9;
    5'b10000 : xpb = 1024'h84b5978fb97391858766514b06b7f5336d78a0b6c77e77d122fcc4455b818dbd4f03b6b19522fd4c7dcf6938c7b4aa55df5008fa905f718072b3dd0a6fec9499e78fc2d5e794282498c667e73f4f55079a140f4a8384940988effb7993d44c5496f6dc077bd2568f07c525aaa79d23a4a3b81c46fe633a592de2798ee9ae29ce;
    5'b10001 : xpb = 1024'h1e94a5b31bd5e9a060f94b794ceb07f3bd6668c3ae8b9b0386829cb42157fa7421e6a3b1301d1e082211784006152a7cbeb4b09a63b5a6692b7b93403227d4f49d573e161852cc5bb6b28cc013baefb97b32343fd3e9011fb0071ff478b6eb7e83018e6de511e09f840987b9f734de051cab72bdfc1a53c094baf44502bb8c68;
    5'b10010 : xpb = 1024'h6920f92c402676840591bd7ea37862057eca34016b105ead67e52e789a311432f8120e29953dbd5265b1c68e27d3bb6e0233802059beab9d94e288d42f358a00c76dee04f8a26dd7e738b43b81024e9c505552cdb0d39b468caad66a17c42d3a9e13d2fdff1a633d870dd0a83e9cbe8ee478a8174a1cca584202e9ffa4ab556d;
    5'b10011 : xpb = 1024'h300074fa288ce9edf24b7ace9ab74c5ceb7fc0e521d81dfcb6b06e7600780e9caf4fb293037de0e09f3d59566343b94e19827c02d14e0864daa3f09f170ca5b7d3569452961120f0524d914556de94e317377c30138085cb3c1fae4fca6cc648a1e85646859ed4e035232b78e3478ef5d6bfe8e47d3e3bfa8db64b5bdb8b807;
    5'b10100 : xpb = 1024'h4d8c5ac8c6d95b8283bd29b24038ced7901bc74c0ea24589accd98abd8e09aa8a12065a195587d584d9423e387f2cc862516f746231de5bab711349dee7e7f67a74c193409b0b38b35ab008fc2b5483106969650de22a2839065b15a9bb40e20a530c9f482626fec06567ba5d59c5979253933e795d65a5756235a705fa8810c;
    5'b10101 : xpb = 1024'h9818ae41eb29e86628559bb796c628e9517f9289cb2709338e302a7051b9b467774bd019fa791ca291347231a9b15d776895c6cc1926eaef20782a31eb8c3473d162c922ea0055076631280b2ffca713dbb9b4debb0d3caa6d0967d03ac14fdcc0430e849c6af28a095ac4941d043a02ed066940e3d8d0ef036b502b01984a11;
    5'b10110 : xpb = 1024'h31f7bc654d8c408101e895e5dcf93ba9a16d5a96b2342c65f1b602df1790211e4a2ebd1995733d5e35768138e811dd9e47fa6e6bec7d1fd7d93fe067adc774ce872a44631abef93e841d4ce4046841c5bcd7d9d40b71a9c094208c4b1fa3ef06ac4dc0eb05aa7c9a859f26a36c9bf46365f9bfb7e18fea566a43cae11aa5acab;
    5'b10111 : xpb = 1024'h7c840fde71dccd64a68107eb338695bb62d125d46eb8f00fd31894a390693add205a2791fa93dca87916cf8709d06e8f8b793df1e286250c42a6d5fbaad529dab140f451fb0e9abab4a3745f71afa0a891faf861e85c43e770c442c0beb130c2c760057b1fb2ff3888a36f91b403d4ed2dc6f5112f9260ee178bc09bbc9575b0;
    5'b11000 : xpb = 1024'h16631e01d43f257f8014021979b9a87bb2beede155c61342369e6d12563fa793f33d1491958dfd641d58de8e4830eeb66adde591b5dc59f4fb6e8c316d106a3567086f922bcd3ef1d28f9938461b3b5a73191d5738c0b0fd97db673ba393cfecb36ab7e188f2894904e7d1a1039b8f4da6ba4b882d497a557e643b51d5a2d84a;
    5'b11001 : xpb = 1024'h60ef717af88fb26324ac741ed047028d7422b91f124ad6ec1800fed6cf18c152c9687f09faae9cae60f92cdc69ef7fa7ae5cb517abe55f2964d581c56a1e1f41911f1f810c1ce06e0315c0b3b3629a3d483c3be515ab4b24747f1db142a111a8ce7cfc71a2fb0be707ec1a8f4b036fd76e8780e17b4bf0ed2bac310c7792a14f;
    5'b11010 : xpb = 1024'hab7bc4f41ce03f46c944e62426d45c9f3586845ccecf9a95f963909b47f1db119f93e9825fcf3bf8a4997b2a8bae1098f1db849da1ee645dce3c7759672bd44dbb35cf6fec6c81ea339be82f20a9f9201d5f5a72f295e54b5122d426e1ae5364e98f4101bd038e850af0637d926b50613654b63ac94e6784d8f426c719826a54;
    5'b11011 : xpb = 1024'h455ad3177f429761a2d7e0526d076f5f85744c69b5dcbdc85ce9690a0dc847c87276d681fac95cb448db8a31ca0e90bfd1402c3d7544994687042d8f296714a870fd4ab01d2b262151880d07f51593d1fe7d7f6842fa52617839f8a1c690f28ed599f368264318958734c58ce2030ac1af480cb1c70580ec3fcca17d328fccee;
    5'b11100 : xpb = 1024'h8fe72690a393244547705257c394c97146d817a7726181723e4bface86a1618748a240fa5fe9fbfe8c7bd87febcd21b114befbc36b4d9e7af06b23232674c9b49b13fa9efd7ac79d820e3483625cf2b4d3a09df61fe4ec8854ddaf17659e344af0ac37f8404b9b338a390e7b296aeb4b7715420b1507f783ed149737d47f95f3;
    5'b11101 : xpb = 1024'h29c634b405f57c6021034c8609c7dc3196c5dfb4596ea4a4a1d1d33d4c77ce3e1b852df9fae41cba30bde7872a2da1d7f423a3633ea3d363a932d958e8b00a0f50db75df2e396bd49ffa595c36c88d66b4bec2eb7049599e7bf4d3924a80d374dcb6ea5ea98b2544067d708a7902a5abf008988212bf10eb53ed11eded8cf88d;
    5'b11110 : xpb = 1024'h7452882d2a460943c59bbe8b605536435829aaf215f3684e83346501c550e7fcf1b098726004bc04745e35d54bec32c937a272e934acd8981299ceece5bdbf1b7af225ce0e890d50d08080d7a40fec4989e1e1794d33f3c558988a07e98e1530f7c92eeec393a7e20981b978c06a8635b7d5cddb60c18783013507a88f7cc192;
    5'b11111 : xpb = 1024'he3196508ca8615e9f2eb8b9a6884903a81772fefd008b80e6ba3d708b2754b3c4938571fafedcc018a044dc8a4cb2f017071a8908030d80cb618522a7f8ff7630b9a10e3f47b187ee6ca5b0787b86fb6b00066e9d9860db7fafae82ce70b45ae3d3e1552cd331f285c61b881002409630c924525e78a0ea680d825ea88a242c;
    endcase
end

endmodule

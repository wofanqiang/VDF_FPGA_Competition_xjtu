module xpb_5_450
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h906a5455549e65f8d23c3003187bc6b8682a28fc41d857df8cb9629fc63e9b93e255822fe6fa5941fbef12171063ab6c0aae597bff098d8db173ec7c672f8b08393f354a5d41091a5376864d06d2262f27943c6c0f346a42c8f311a5f5b57c9990abbba482f1f6197f8b0f2ee162b49ffcc759588e935c3f64c81551f0a6d8db;
    5'b00010 : xpb = 1024'h70276354e74e9728d972e82f209d461f5ede4ec7ae390f479b960be9d97a8a1fc16286e703ce33f5587fe4e73d69460db1428b11db604acfb248999a938ca15efe2f35e60af114ef945309f774c8882d5b237f3f91e2a774dc599151314056a0f24fe51f551af3a57856377ecaf54316aab4d3ceccdb5b4e8320af9f586b4b4b;
    5'b00011 : xpb = 1024'h4fe4725479fec858e0a9a05b28bec586559274931a99c6afaa72b533ecb678aba06f8b9e20a20ea8b510b7b76a6ee0af57d6bca7b7b70811b31d46b8bfe9b7b5c31f3681b8a120c4d52f8da1e2beea2b8eb2c2131490e4a6efc010fc6ccb30a853f40e9a2743f13171215fceb487d18d58a24e450b235a5da17949ecc02fbdbb;
    5'b00100 : xpb = 1024'h2fa181540caef988e7e0588730e044ed4c469a5e86fa7e17b94f5e7dfff267377f7c90553d75e95c11a18a8797747b50fe6aee3d940dc553b3f1f3d6ec46ce0c880f371d66512c9a160c114c50b54c29c24204e6973f21d9032690a7a8560aafb5983814f96ceebd69ec881e9e1a6004068fc8bb496b596cbfd1e43a27f4302b;
    5'b00101 : xpb = 1024'hf5e90539f5f2ab8ef1710b33901c45442fac029f35b357fc82c07c8132e55c35e89950c5a49c40f6e325d57c47a15f2a4ff1fd370648295b4c6a0f518a3e4634cff37b91401386f56e894f6beabae27f5d147ba19ed5f0b168d1052e3e0e4b7173c618fcb95ec4962b7b06e87acee7ab47d433187b3587bde2a7e878fb8a29b;
    5'b00110 : xpb = 1024'h9fc8e4a8f3fd90b1c15340b6517d8b0cab24e92635338d5f54e56a67d96cf15740df173c41441d516a216f6ed4ddc15eafad794f6f6e1023663a8d717fd36f6b863e6d0371424189aa5f1b43c57dd4571d6584262921c94ddf8021f8d9966150a7e81d344e87e262e242bf9d690fa31ab1449c8a1646b4bb42f293d9805f7b76;
    5'b00111 : xpb = 1024'h7f85f3a886adc1e1c889f8e2599f0a73a1d90ef1a19444c763c213b1eca8dfe31fec1bf35e17f804c6b2423f01e35c005641aae54bc4cd65670f3a8fac3085c24b2e6d9f1ef24d5eeb3b9eee3374365550f4c6f9abd0067ff2e6a1a415213b58098c46af20b0dfeedb0de7ed52a231915f321700548eb3ca614b2e26e823ede6;
    5'b01000 : xpb = 1024'h5f4302a8195df311cfc0b10e61c089da988d34bd0df4fc2f729ebcfbffe4ce6efef920aa7aebd2b82343150f2ee8f6a1fcd5dc7b281b8aa767e3e7add88d9c19101e6e3acca259342c182298a16a9853848409cd2e7e43b2064d214f50ac155f6b307029f2d9dd7ad3d9103d3c34c0080d1f917692d6b2d97fa3c8744fe86056;
    5'b01001 : xpb = 1024'h3f0011a7ac0e2441d6f7693a69e209418f415a887a55b397817b66461320bcfade06256197bfad6b7fd3e7df5bee9143a36a0e11047247e968b894cc04eab26fd50e6ed67a5265096cf4a6430f60fa51b8134ca0b12c80e419b3a0fa8c36ef66ccd499a4c502db06cca4388d25c74e7ebb0d0becd11eb1e89dfc62c1b7acd2c6;
    5'b01010 : xpb = 1024'h1ebd20a73ebe5571de2e2166720388a885f58053e6b66aff90580f90265cab86bd132a18b493881edc64baaf88f42be549fe3fa6e0c9052b698d41ea3147c8c699fe6f72280270deadd129ed7d575c4feba28f7433dabe162d1a20a5c7c1c96e2e78c31f972bd892c56f60dd0f59dcf568fa86630f66b0f7bc54fd0f1f714536;
    5'b01011 : xpb = 1024'haf2774fc935cbb6ab06a51698a7f4f60ee1fa950288ec2df1d11722fec9b471a9f68ac489b8de160d853ccc69957d75154ac9922dfd292b91b012e66987753ced33da4bc854379f90147b03a8429827f1336cbe0430f2858f60d324bbd774607bf247ec41a1dceac44fa700bf0bc919565c1dfbb9dfa0d37211d126110181e11;
    5'b01100 : xpb = 1024'h8ee483fc260cec9ab7a1099592a0cec7e4d3cf1b94ef7a472bee1b79ffd735a67e75b0ffb861bc1434e49f96c65d71f2fb40cab8bc294ffb1bd5db84c4d46a25982da55832f385ce422433e4f21fe47d46c60eb3c5bd658b0973b1f6f902200f20c8a83eec46cc383dc5985bda4f200c13af5a31dc420c463f75acae77dc9081;
    5'b01101 : xpb = 1024'h6ea192fbb8bd1dcabed7c1c19ac24e2edb87f4e7015031af3acac4c4131324325d82b5b6d53596c791757266f3630c94a1d4fc4e98800d3d1caa88a2f131807c5d1da5f3e0a391a38300b78f6016467b7a555187486ba2bd1cda31a2348cfa16826cd1b9be6fc9c43690c0abc3e1ae82c19cd4a81a8a0b555dce46fbdfa102f1;
    5'b01110 : xpb = 1024'h4e5ea1fb4b6d4efac60e79eda2e3cd95d23c1ab26db0e91749a76e0e264f12be3c8fba6df209717aee0645372068a73648692de474d6ca7f1d7f35c11d8e96d3220da68f8e539d78c3dd3b39ce0ca879ade4945acb19dfef3040b14d7017d41de410fb349098c7502f5be8fbad743cf96f8a4f1e58d20a647c26e14947657561;
    5'b01111 : xpb = 1024'h2e1bb0fade1d802acd453219ab054cfcc8f0407dda11a07f58841758398b014a1b9cbf250edd4c2e4a9718074d6e41d7eefd5f7a512d87c11e53e2df49ebad29e6fda72b3c03a94e04b9bee43c030a77e173d72e4dc81d2143a730f8aba2ae2545b524af62c1c4dc2827114b9706cb701d77c994971a09739a7f7b96af29e7d1;
    5'b10000 : xpb = 1024'hdd8bffa70cdb15ad47bea45b326cc63bfa46649467257e76760c0a24cc6efd5faa9c3dc2bb126e1a727ead77a73dc79959191102d8445031f288ffd7648c380abeda7c6e9b3b5234596428ea9f96c7615031a01d0765a53570db0a3e72d882ca7594e2a34eac26820f2399b809959e6cb65440ad5620882b8d815e416ee5a41;
    5'b10001 : xpb = 1024'h9e43144fc56c1753a6b81a48cba2931c27ce8f45884aafc6f41a234213058b69dcff460c12ab8023a316fcee8ad787e5a03fea8c2c8dd290d09c7c79dd784e88e52cdd1146f4be3d990cc8dbb0cb92a53c97566ddfaac4962000c249dce304c6380509ceb7dcb881a07d48ca61fc0e86c82c9d6363f564c21da02b360795331c;
    5'b10010 : xpb = 1024'h7e00234f581c4883adeed274d3c412831e82b510f4ab672f02f6cc8c264179f5bc0c4ac32f7f5ad6ffa7cfbeb7dd228746d41c2208e48fd2d171299809d564dfaa1cddacf4a4ca12d9e94c861ec1f4a370269941625901c8336741f5186ddecd99a933498a05b60d9948711a4b8e9cfd761a17d9a23d63d13bf8c5836f59a58c;
    5'b10011 : xpb = 1024'h5dbd324eeacc79b3b5258aa0dbe591ea1536dadc610c1e9711d375d6397d68819b194f7a4c53358a5c38a28ee4e2bd28ed684db7e53b4d14d245d6b636327b366f0cde48a254d5e81ac5d0308cb856a1a3b5dc14e5073efa46cdc1a053f8b8d4fb4d5cc45c2eb3999213996a35212b742407924fe08562e05a515fd0d71e17fc;
    5'b10100 : xpb = 1024'h3d7a414e7d7caae3bc5c42cce40711510beb00a7cd6cd5ff20b01f204cb9570d7a2654316927103db8c9755f11e857ca93fc7f4dc1920a56d31a83d4628f918d33fcdee45004e1bd5ba253dafaaeb89fd7451ee867b57c2c5a34414b8f8392dc5cf1863f2e57b1258adec1ba1eb3b9ead1f50cc61ecd61ef78a9fa1e3ee28a6c;
    5'b10101 : xpb = 1024'h1d37504e102cdc13c392faf8ec2890b8029f267339cd8d672f8cc86a5ff54599593358e885faeaf1155a482f3eedf26c3a90b0e39de8c798d3ef30f28eeca7e3f8ecdf7ffdb4ed929c7ed78568a51a9e0ad461bbea63b95e6d9ac0f6cb0e6ce3be95afba0080aeb183a9ea0a084648617fe2873c5d1560fe9702946ba6a6fcdc;
    5'b10110 : xpb = 1024'hada1a4a364cb420c95cf2afc04a457706ac94f6f7ba5e546bc462b0a2633e12d3b88db186cf5443311495a464f519dd8453f0a5f9cf2552685631d6ef61c32ec322c14ca5af5f6aceff55dd26f7740cd32689e27f99823a1368dd29cc0c3e97d4f416b5e8372a4cb0334f938e9a8fd017ca9e094eba8bd3dfbcaa9bd974dd5b7;
    5'b10111 : xpb = 1024'h8d5eb3a2f77b733c9d05e3280cc5d6d7617d753ae8069caecb22d454396fcfb91a95dfcf89c91ee66dda2d167c573879ebd33bf5794912688637ca8d22794942f71c156608a6028230d1e17cdd6da2cb65f7e0fb7c4660d349f45247fc4ec384b0e594d9559ba256fc002188d33b8b782a975b0b29f0bc4d1a23440aff124827;
    5'b11000 : xpb = 1024'h6d1bc2a28a2ba46ca43c9b5414e7563e58319b0654675416d9ff7d9e4cabbe44f9a2e486a69cf999ca6affe6a95cd31b92676d8b559fcfaa870c77ab4ed65f99bc0c1601b6560e5771ae65274b6404c9998723cefef49e055d5ad1f337d99d8c1289be5427c49fe2f4cb49d8bcce19eed884d5816838bb5c387bde5866d6ba97;
    5'b11001 : xpb = 1024'h4cd8d1a21cdbd59cab7353801d08d5a54ee5c0d1c0c80b7ee8dc26e85fe7acd0d8afe93dc370d44d26fbd2b6d6626dbd38fb9f2131f68cec87e124c97b3375f080fc169d64061a2cb28ae8d1b95a66c7cd1666a281a2db3770c1519e73647793742de7cef9ed9d6eed967228a660a86586724ff7a680ba6b56d478a5ce9b2d07;
    5'b11010 : xpb = 1024'h2c95e0a1af8c06ccb2aa0bac252a550c4599e69d2d28c2e6f7b8d03273239b5cb7bcedf4e044af00838ca5870368085edf8fd0b70e4d4a2e88b5d1e7a7908c4745ec173911b62601f3676c7c2750c8c600a5a976045118698427d149aeef519ad5d21149cc169afae6619a788ff336dc345fca6de4c8b97a752d12f3365f9f77;
    5'b11011 : xpb = 1024'hc52efa1423c37fcb9e0c3d82d4bd4733c4e0c6899897a4f0695797c865f89e896c9f2abfd1889b3e01d7857306da3008624024ceaa40770898a7f05d3eda29e0adc17d4bf6631d73443f02695472ac43434ec4986ff559b978e50f4ea7a2ba237763ac49e3f9886df2cc2c87985c552e24d44e42310b8899385ad409e2411e7;
    5'b11100 : xpb = 1024'h9cbd43f696da9df58c1cf3db45c79b2ba4783564db61d22e934edc1c4c9e257c791f74dbe412e2f5dc0c8a6e40d14e6c90d25bc8e9ad94fe3afe6b823b1d2da6441b4d1f1ca73af187ba76739c1950f35bc928b59633bfde6081629ae02fa83bc821f66921318ea05eb7d1f75ae879f2df149e3cb1a414c8f84dc2928ecaeac2;
    5'b11101 : xpb = 1024'h7c7a52f6298acf259353ac074de91a929b2c5b3047c28996a22b85665fda1408582c799300e6bda9389d5d3e6dd6e90e37668d5ec60452403bd318a0677a43fd090b4dbaca5746c6c896fa1e0a0fb2f18f586b8918e1fd1073e7e2461bba824329c61fe3f35a8c2c5782fa47447b08698d0218b2efec13d816a65cdff68f5d32;
    5'b11110 : xpb = 1024'h5c3761f5bc3b00559a8a6433560a99f991e080fbb42340feb1082eb07316029437397e4a1dba985c952e300e9adc83afddfabef4a25b0f823ca7c5be93d75a53cdfb4e567807529c09737dc8780614efc2e7ae5c9b903a42874e61f157455c4a8b6a495ec58389b8504e22972e0d96e03aef93292e3412e734fef72d5e53cfa2;
    5'b11111 : xpb = 1024'h3bf470f54eeb3185a1c11c5f5e2c19608894a6c72083f866bfe4d7fa8651f120164683013a8e730ff1bf02dec7e21e51848ef08a7eb1ccc43d7c72dcc03470aa92eb4ef225b75e714a500172e5fc76edf676f1301e3e77749ab4e19c92d03651ed0e72d997ac874449194ae717a02556e8dd0d9f6c7c11f65357917ac6184212;
    endcase
end

endmodule

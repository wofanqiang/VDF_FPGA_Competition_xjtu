module xpb_5_575
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h6dfa7b5b827bd0d96593575a0b38a8d16981d41c13d8175007e7ea861056ee29384f9e49ddfcd73e038bbdfd6e438f2f76398e8dadd2267acaf2b2977056c2c7b4ed63c6976d4ed5f8075893ef5eb55b5727115cfa03b046722650c5a247adb41371501a770a467d58b2cf37d02932a4b9138a4b3b95138ff924c64402ad38c4;
    5'b00010 : xpb = 1024'h2b47b16143096cea002136dd06170a51618da50752388e2891f31bb66dab2f4a6d56bf1af1d32fed67b93cb3f9290d948858f53538f17ca9e54625d0a5db10ddf58b92de7f49a066dd74ae8545e1a685ba4929216781337c2ec00f908a64b8d5f7db0e0b3d4b946d2aa5b790a8823f20234d35b426dec9efabda11837c780b1d;
    5'b00011 : xpb = 1024'h99422cbcc5853dc365b48e37114fb322cb0f79236610a57899db063c7e021d73a5a65d64cfd0072b6b44fab1676c9cc3fe9283c2e6c3a324b038d8681631d3a5aa78f6a516b6ef3cd57c071935405be111703a7e6184e3c2a0e660562cac668a0b4c5e25b455daea835886c878ab71c4dc60bfff6273dd7fa4fed7c77f2543e1;
    5'b00100 : xpb = 1024'h568f62c28612d9d400426dba0c2e14a2c31b4a0ea4711c5123e6376cdb565e94daad7e35e3a65fdacf727967f2521b2910b1ea6a71e2f953ca8c4ba14bb621bbeb1725bcfe9340cdbae95d0a8bc34d0b74925242cf0266f85d801f2114c971abefb61c167a9728da554b6f2151047e40469a6b684dbd93df57b42306f8f0163a;
    5'b00101 : xpb = 1024'h13dc98c846a075e49ad04d3d070c7622bb271af9e2d19329adf1689d38aa9fb60fb49f06f77cb88a339ff81e7d37998e22d15111fd024f82e4dfbeda813a6fd22bb554d4e66f925ea056b2fbe2463e35d7b46a073c7fea2e1a19ddebfce67ccdd41fda0740d876ca273e577a295d8abbb0d416d139074a3f0a696e4672bae893;
    5'b00110 : xpb = 1024'h81d71423c91c46be0063a49712451ef424a8ef15f6a9aa79b5d9532349018ddf48043d50d5798fc8372bb61beb7b28bd990adf9faad475fdafd27171f1913299e0a2b89b7ddce134985e0b8fd1a4f3912edb7b6436839a748c402eb19f2e2a81e7912a21b7e2bd477ff126b1f986bd6069e7a11c749c5dcf038e348a75682157;
    5'b00111 : xpb = 1024'h3f244a2989a9e2ce9af1841a0d2380741cb4c001350a21523fe48453a655cf007d0b5e21e94fe8779b5934d27660a722ab2a464735f3cc2cca25e4ab271580b02140e7b365b932c57dcb61812827e4bb91fd9328a4011daa48d9ed7c874b35a3cbfae8127e240b3751e40f0ad1dfc9dbd4214c855fe6142eb6437fc9ef32f3b0;
    5'b01000 : xpb = 1024'had1ec5850c25b3a80084db74185c29458636941d48e238a247cc6ed9b6acbd29b55afc6bc74cbfb59ee4f2cfe4a436522163d4d4e3c5f2a795189742976c4377d62e4b79fd26819b75d2ba1517869a16e924a4859e04cdf0bb003e422992e357df6c382cf52e51b4aa96de42a208fc808d34d6d09b7b27beaf68460df1e02c74;
    5'b01001 : xpb = 1024'h6a6bfb8accb34fb89b12baf7133a8ac57e4265088742af7ad1d7a00a1400fe4aea621d3cdb231865031271866f89b4b733833b7c6ee548d6af6c0a7bccf0918e16cc7a91e502d32c5b4010066e098b414c46bc4a0b8251267799fd0d11afee79c3d5f61dbb6f9fa47c89c69b7a6208fbf76e823986c4de1e621d914d6baafecd;
    5'b01010 : xpb = 1024'h27b931908d40ebc935a09a7a0e18ec45764e35f3c5a326535be2d13a71553f6c1f693e0deef97114673ff03cfa6f331c45a2a223fa049f05c9bf7db50274dfa4576aa9a9ccdf24bd40ad65f7c48c7c6baf68d40e78ffd45c3433bbd7f9ccf99ba83fb40e81b0ed944e7caef452bb157761a82da2720e947e14d2dc8ce575d126;
    5'b01011 : xpb = 1024'h95b3acec0fbcbca29b33f1d419519516dfd00a0fd97b3da363cabbc081ac2d9557b8dc57ccf648526acbae3a68b2c24bbbdc30b1a7d6c58094b2304c72cba26c0c580d70644c739338b4be8bb3eb31c7068fe56b730384a2a65a0c9d9c14a74fbbb10428f8bb3411a72f7e2c22e4481c1abbb7edada3a80e0df7a2d0e82309ea;
    5'b01100 : xpb = 1024'h5300e2f1d04a58b335c1d157142ff696d7dbdafb17dbb47bedd5ecf0df006eb68cbffd28e0cca101cef92cf0f39840b0cdfb975932f61bafaf05a385a84ff0824cf63c884c28c5241e22147d0a6e22f169b1fd2fe08107d862f3cb688431b271a01ac219befc820179226684fb3d549784f5635698ed5e6dc0acee1061eddc43;
    5'b01101 : xpb = 1024'h104e18f790d7f4c3d04fb0da0f0e5816cfe7abe6563c2b5477e11e213c54afd7c1c71df9f4a2f9b13326aba77e7dbf15e01afe00be1571dec95916beddd43e988d946ba0340516b5038f6a6e60f1141bccd414f44dfe8b0e1f8d8a336c4ebd938484800a853dcff14b154eddd3966112ef2f0ebf843714cd7362394fdbb8ae9c;
    5'b01110 : xpb = 1024'h7e4894531353c59d35e308341a4700e8396980026a1442a47fc908a74cab9e00fa16bc43d29fd0ef36b269a4ecc14e4556548c8e6be79859944bc9564e2b01604281cf66cb72658afb96c302504fc97723fb265148023b5491b3daf90e966b4797f5d024fc48166ea3c81e15a3bf93b7a842990abfcc285d6c86ff93de65e760;
    5'b01111 : xpb = 1024'h3b95ca58d3e161add070e7b715256268317550eda874b97d09d439d7a9ffdf222f1ddd14e676299e9adfe85b77a6ccaa6873f335f706ee88ae9f3c8f83af4f76831ffe7eb34eb71be10418f3a6d2baa1871d3e15b57fbe8a4e4d99c3f6b376697c5f8e15c289645e75bb066e7c18a033127c4473ab15debd1f3c4ad35830b9b9;
    5'b10000 : xpb = 1024'ha99045b4565d328736043f11205e0b399af72509bc4cd0cd11bc245dba56cd4b676d7b5ec47300dc9e6ba658e5ea5bd9dead81c3a4d915037991ef26f406123e380d62454abc05f1d90b718796316ffcde444f72af836ed0c073ea8998fb241d8fd0de303993aadbce6dd5a64c41d2d7cb8fcebee6aaf24d186111175addf27d;
    5'b10001 : xpb = 1024'h66dd7bba16eace97d0921e941b3c6cb99302f5f4faad47a59bc7558e17ab0e6c9c749c2fd849598c0299250f70cfda3ef0cce86b2ff86b3293e56260298a605478ab915d32985782be78c778ecb46127416667371d00f2067d0da95481182f3f743a9c20ffd4f8cba060bdff249adf5335c97a27d1f4a8accb165c56d4a8c4d6;
    5'b10010 : xpb = 1024'h242ab1bfd7786aa86b1ffe17161ace398b0ec6e0390dbe7e25d286be74ff4f8dd17bbd00ec1fb23b66c6a3c5fbb558a402ec4f12bb17c161ae38d5995f0eae6ab949c0751a74a913a3e61d6a43375251a4887efb8a7e753c39a7681f69353a6158a45a11c61646bb7253a657fcf3ebcea0032590bd3e5f0c7dcba7964e73972f;
    5'b10011 : xpb = 1024'h92252d1b59f43b81d0b355712153770af4909afc4ce5d5ce2dba714485563db709cb5b4aca1c89796a5261c369f8e7d37925dda068e9e7dc792b8830cf6571326e37243bb1e1f7e99bed75fe329607acfbaf905884822582abcdb8e50b7ce8156c15aa2c3d208d38cb06758fcd1d1e735916afdbf8d3729c76f06dda5120cff3;
    5'b10100 : xpb = 1024'h4f7263211a81d7926b4134f41c31d88aec9c6be78b464ca6b7c5a274e2aa7ed83ed27c1bddf2e228ce7fe079f4de66388b454447f4093e0b937efb6a04e9bf48aed5535399be497a815acbef8918f8d75ed1a81cf1ffa8b8686777aff399f337507f681d0361db289cf95de8a5762aeec3505b44e41d28fc29a5b919caeba24c;
    5'b10101 : xpb = 1024'hcbf9926db0f73a305cf147717103a0ae4a83cd2c9a6c37f41d0d3a53ffebff973d99cecf1c93ad832ad5f307fc3e49d9d64aaef7f28943aadd26ea33a6e0d5eef73826b819a9b0b66c821e0df9bea01c1f3bfe15f7d2bee2501367adbb6fe5934e9260dc9a329186eec46417dcf376a2d8a06adcf66df5bdc5b045944b674a5;
    5'b10110 : xpb = 1024'h7aba14825d8b447c6b626bd12248e2dc4e2a10eedd7edacf49b8be2b5055ae22ac293b36cfc6121636391d2dee0773cd139e397d2cfabab578c5213aaac4d026a460e6321907e9e15ecf7a74cefa9f5d191ad13e5980dc34972787407dfeac0d485a762840ad6f95c79f15794df86a0ee69d90f90afbf2ebd57fca9d4763ad69;
    5'b10111 : xpb = 1024'h38074a881e18e08d05f04b541d27445c4635e1da1bdf51a7d3c3ef5bada9ef43e1305c07e39c6ac59a669be478ecf23225bda024b81a10e493189473e0491e3ce4ff154a00e43b72443cd066257d90877c3ce902c6fe5f6a53c1460b661bb72f2cc4341906eebd859991fdd22651768a50d73c61f645a94b883515dcc12e7fc2;
    5'b11000 : xpb = 1024'ha601c5e3a094b1666b83a2ae285fed2dafb7b5f62fb768f7dbabd9e1be00dd6d197ffa51c19942039df259e1e73081619bf72eb265ec375f5e0b470b509fe10499ec791098518a483c4428fa14dc45e2d363fa5fc1020fb0c5e796d1086364e3403584337df90402f244cd09f67aa92f09eac6ad31dabcdb8159dc20c3dbb886;
    5'b11001 : xpb = 1024'h634efbe961224d7706118231233e4eada7c386e16e17dfd065b70b121b551e8e4e871b22d56f9ab3021fd8987215ffc6ae169559f10b8d8e785eba4486242f1ada8aa828802ddbd921b17eeb6b5f370d368612242e7f92e68281559bf0807005249f4224443a51f2c437b562ced3b5aa742472161d24733b340f27603da68adf;
    5'b11010 : xpb = 1024'h209c31ef21afe987a09f61b41e1cb02d9fcf57ccac7856a8efc23c4278a95faf838e3bf3e945f362664d574efcfb7e2bc035fc017c2ae3bd92b22d7dbba87d311b28d740680a2d6a071ed4dcc1e2283799a829e89bfd161c3f1b1466d89d7b27090900150a7b9fe2962a9dbba72cc225de5e1d7f086e299ae6c4729fb7715d38;
    5'b11011 : xpb = 1024'h8e96ad4aa42bba610632b90e295558ff09512be8c0506df8f7aa26c889004dd8bbddda3dc742caa069d9154c6b3f0d5b366f8a8f29fd0a385da4e0152bff3ff8d0163b06ff777c3fff262d70b140dd92f0cf3b459600c662b141652c7ae528db1c7a502f8185e65feedd6cf37755f4ca9771a7ca44033d2adfe938e3ba1e95fc;
    5'b11100 : xpb = 1024'h4be3e35064b95671a0c098912433ba7f015cfcd3feb0e4d181b557f8e6548ef9f0e4fb0edb19234fce069402f6248bc0488ef136b51c606777f8534e61838e0f10b46a1ee753cdd0e493836207c3cebd53f1530a037e49986ddb23f7630233fd00e40e2047c7344fc0d0554c4faf014601ab53332f4cf38a929e842333e96855;
    5'b11101 : xpb = 1024'h93119562546f2823b4e78141f121bfef968cdbf3d115baa0bc0892943a8d01b25ec1bdfeeef7bff323412b9810a0a255aae57de403bb696924bc6879707dc2551529936cf301f61ca00d9535e46bfe7b7136ace70fbccce2a74e2c24b1f3f1ee54dcc110e08823f92c33da528080dc16be4fe9c1a96a9ea4553cf62adb43aae;
    5'b11110 : xpb = 1024'h772b94b1a7c2c35ba0e1cf6e2a4ac4d062eaa1db50e972fa13a873af53ffbe445e3bba29ccec533d35bfd0b6ef4d9954d0e7e66bee0ddd115d3e791f075e9eed063ffcfd669d6e37c20831e74da575430e3a7c2b6aff7d149c9b3387ed66ecd2f8bf1c2b8512c8bceb760cdcf831406624f888e7562bbd7a3e7895a6b0617372;
    5'b11111 : xpb = 1024'h3478cab768505f6c3b6faef1252926505af672c68f49e9d29db3a4dfb153ff659342dafae0c2abec99ed4f6d7a3317b9e3074d13792d33407791ec583ce2ed0346de2c154e79bfc8a77587d8a428666d715c93efd87d004a5934f252d583f7f4dd28da1c4b5416acbd68f535d08a4ce18f323450417573d9f12de0e62a2c45cb;
    endcase
end

endmodule

module xpb_5_535
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h3c73bf4c18db77b3d9b5479e39ffc9552814927d5793f89fb201560eedea4c933a75b476121d8fb896dbec4af9b36983926ddaac93b558db96ebf0d1737ba8659254899c164c8a2a1492e624b91b04ac8827d8aaf819d899ea9852c59169a90c0a7173cbf5a8fae5ccb1118f9d23fb5f0ff048c79472762794341dcd7798ffd4;
    5'b00010 : xpb = 1024'h78e77e9831b6ef67b36a8f3c73ff92aa502924faaf27f13f6402ac1ddbd4992674eb68ec243b1f712db7d895f366d30724dbb559276ab1b72dd7e1a2e6f750cb24a913382c9914542925cc4972360959104fb155f033b133d530a58b22d3521814e2e797eb51f5cb9962231f3a47f6be1fe0918f28e4ec4f28683b9aef31ffa8;
    5'b00011 : xpb = 1024'h4adf88e88a43252c21a5f039da514ae06c7b44731444967982748d716bc38b1ac189fe96c32309b2535859a09bc2bc0532f681f986d3a47142493161fa0847f42ae68259354a1392b1eafcb927549d4a47290685bc75cbd0a3c6655fa125891f04cc93a3031f823df534dcfdf9bcbf3e0f6fb746d0c0546762cde63dde89911;
    5'b00100 : xpb = 1024'h4121b7daa17faa069bcfa6a1d7a4de032edc46c488d842074a289ee604a68544e68e545f7e4fc053bc1171e5036f9543e59d42cc2c229322ab1083e7931c2ce4d502f1c1a9a12b633fb195f04b904e812c9a691353e13556f4d4b91b8b7c019dfabe3d0625daf309ac045f5f7cbfc752f0e7443c017e7b6e0a60fc31558198e5;
    5'b00101 : xpb = 1024'h7d957726ba5b21ba7584ee4011a4a75856f0d941e06c3aa6fc29f4f4f290d1d8210408d5906d500c52ed5e2ffd22fec7780b1d78bfd7ebfe41fc74b90697d54a67577b5dbfedb58d54447c1504ab532db4c241be4bfb0df0df6d0be11ce5aaaa052fb0d21b83edef78b570ef19e3c2b200d78d0395f0f1959e9519fecd1a98b9;
    5'b00110 : xpb = 1024'h95bf11d114864a58434be073b4a295c0d8f688e628892cf304e91ae2d78716358313fd2d86461364a6b0b3413785780a65ed03f30da748e2849262c3f4108fe855cd04b26a94272563d5f9724ea93a948e520d0b78eb97a1478ccabf424b123e09992746063f047bea69b9fbf3797e7c1edf6e8da180a8cec59bcc7bbd13222;
    5'b00111 : xpb = 1024'h45cfb0692a23dc595dea05a57549f2b135a3fb0bba1c8b6ee24fe7bd1b62bdf692a6f448ea81f0eee146f77f0d2bc10438ccaaebc48fcd69bf3516fdb2bcb16417b159e73cf5cc9c6ad045bbde059855d10cf97bafa89213ff111f71858e5a2feb0b0640560ceb2d8b57ad2f5c5b9346d1de3fb06e8a80b4808dda95336a31f6;
    5'b01000 : xpb = 1024'h82436fb542ff540d379f4d43af49bc065db88d8911b0840e94513dcc094d0a89cd1ca8befc9f80a77822e3ca06df2a87cb3a859858452645562107cf263859c9aa05e383534256c67f632be097209d025934d226a7c26aade9a9723716f8033bf57c7a0c4bb5e6135808bebef97f8ea5e1ce887802fcf6dc14c1f862ab0331ca;
    5'b01001 : xpb = 1024'he09e9ab99ec96f8464f1d0ad8ef3e0a14571cd593ccdc36c875da854434aa150449dfbc449691d16fa090ce1d348340f98e385ec947aed53c6db9425ee18d7dc80b3870b9fde3ab815c0f62b75fdd7ded57b139135616371eb53301ee3709b5d0e65bae9095e86b9df9e96f9ed363dba2e4f25d47240fd362869b2b99b9cb33;
    5'b01010 : xpb = 1024'h4a7da8f7b2c80eac200464a912ef075f3c6baf52eb60d4d67a773094321ef6a83ebf943256b4218a067c7d1916e7ecc48bfc130b5cfd07b0d359aa13d25d35e35a5fc20cd04a6dd595eef587707ae22a757f89e40b6feed1094d85c77fa0b2c1db57cf7a863ee3516aaafaff3bf75f3ab2d53b24db9685faf6bab8f91152cb07;
    5'b01011 : xpb = 1024'h86f16843cba3865ff9b9ac474ceed0b4648041d042f4cd762c7886a32009433b793548a868d1b1429d586964109b56481e69edb7f0b2608c6a459ae545d8de48ecb44ba8e696f7ffaa81dbac2995e6d6fda7628f0389c76af3e5d88d110a5bcde5c943467be7de37375c0c8ed91b5a99c2c583ec7008fc228aeed6c688ebcadb;
    5'b01100 : xpb = 1024'h12b7e23a2290c94b08697c0e769452b81b1ed11cc511259e609d235c5af0e2c6b0627fa5b0c8c26c94d6166826f0af014cbda07e61b4e91c50924c587e8211fd0ab9a0964d5284e4ac7abf2e49d5275291ca41a16f1d72f428f19957e8496247c13324e8c0c7e08f7d4d373f7e6f2fcf83dbedd1b4301519d8b3798f77a26444;
    5'b01101 : xpb = 1024'h4f2ba1863b6c40fee21ec3acb0941c0d4333639a1ca51e3e129e796b48db2f59ead8341bc2e652252bb202b320a41884df2b7b2af56a41f7e77e3d29f1fdba629d0e2a32639f0f0ec10da55302f02bff19f21a4c67374b8e1389ec1d79b30b53cba498b4b670db7549fe48cf1b932b2e93cc369948a28b416ce7975cef3b6418;
    5'b01110 : xpb = 1024'h8b9f60d25447b8b2bbd40b4aea93e5626b47f617743916ddc49fcf7a36c57bed254de891d503e1ddc28deefe1a578208719955d7891f9ad37e6a2dfb657962c82f62b3ce79eb9938d5a08b77bc0b30aba219f2f75f512427fe223ee30b1cb45fd6160c80ac19d65b16af5a5eb8b7268da3bc7f60dd150169011bb52a66d463ec;
    5'b01111 : xpb = 1024'h1765dac8ab34fb9dca83db121439676621e68563f6556f05f8c46c3371ad1b785c7b1f8f1cfaf307ba0b9c0230acdac19fed089dfa22236364b6df6e9e22967c4d6808bbe0a7261dd7996ef9dc4a7127363cd209cae4cfb1332dffade25bbad9b17fee22f0f9d8b35ca0850f5e0afbc364d2e946213c1a604ee057f3558afd55;
    5'b10000 : xpb = 1024'h53d99a14c4107351a43922b04e3930bb49fb17e14de967a5aac5c2425f97680b96f0d4052f1882c050e7884d2a604445325ae34a8dd77c3efba2d040119e3ee1dfbc9257f6f3b047ec2c551e956575d3be64aab4c2fea84b1dc6527373c563e5bbf161eee6a2d3992951969efb2ef72274c3320db5ae9087e31475c0cd23fd29;
    5'b10001 : xpb = 1024'h904d5960dcebeb057dee6a4e8838fa10720faa5ea57d60455cc718514d81b49ed166887b41361278e7c374982413adc8c4c8bdf7218cd51a928ec1118519e74772111bf40d403a7200bf3b434e807a80468c835fbb1880e5085ea539052f0cf1c662d5badc4bce7ef602a82e9852f28184b37ad54a2106af7748938e44bcfcfd;
    5'b10010 : xpb = 1024'h1c13d35733d92df08c9e3a15b1de7c1428ae39ab2799b86d90ebb50a8869542a0893bf78892d23a2df41219c3a690681f31c70bd928f5daa78db7284bdc31afb901670e173fbc75702b81ec56ebfbafbdaaf627226ac2c6e3d6a6603dc6e136ba1ccb75d212bd0d73bf3d2df3da6c7b745c9e4ba8e481fa6c50d365733739666;
    5'b10011 : xpb = 1024'h588792a34cb4a5a4665381b3ebde456950c2cc287f2db10d42ed0b197653a0bd430973ee9b4ab35b761d0de7341c7005858a4b6a2644b6860fc76356313ec361226afa7d8a485181174b04ea27dabfa862d73b1d1ec605082802b8c96dd7bc77ac3e2b2916d4cbbd08a4e46edacac31655ba2d8222ba95ce59415424ab0c963a;
    5'b10100 : xpb = 1024'h94fb51ef65901d584008c95225de0ebe78d75ea5d6c1a9acf4ee6128643ded507d7f2864ad6843140cf8fa322dcfd98917f82616b9fa0f61a6b35427a4ba6bc6b4bf8419a094dbab2bddeb0ee0f5c454eaff13c816dfdda2129b0b8eff416583b6af9ef50c7dc6a2d555f5fe77eebe7565aa7649b72d0bf5ed7571f222a5960e;
    5'b10101 : xpb = 1024'h20c1cbe5bc7d60434eb899194f8390c22f75edf258de01d52912fde19f258cdbb4ac5f61f55f543e0476a73644253242464bd8dd2afc97f18d00059add639f7ad2c4d907075068902dd6ce91013504d07f21f2da8273892b47a6cc59d6806bfd92198097515dc8fb1b4720af1d4293ab26c0e02efb5424ed3b3a14bb115c2f77;
    5'b10110 : xpb = 1024'h5d358b31d558d7f7286de0b789835a17578a806fb071fa74db1453f08d0fd96eef2213d8077ce3f69b5293813dd89bc5d8b9b389beb1f0cd23ebf66c50df47e0651962a31d9cf2ba4269b4b5ba50097d0749cb857a8d61c5323f1f1f67ea15099c8af4634706c3e0e7f8323eba668f0a36b128f68fc69b14cf6e328888f52f4b;
    5'b10111 : xpb = 1024'h99a94a7dee344fab02232855c383236c7f9f12ed0805f3148d15a9ff7afa26022997c84e199a73af322e7fcc378c05496b278e36526749a8bad7e73dc45af045f76dec3f33e97ce456fc9ada736b0e298f71a43072a73a5f1cd771e4f953be15a6fc682f3cafbec6b4a943ce578a8a6946a171be2439113c63a25056008e2f1f;
    5'b11000 : xpb = 1024'h256fc4744521929610d2f81ced28a570363da2398a224b3cc13a46b8b5e1c58d60c4ff4b619184d929ac2cd04de15e02997b40fcc369d238a12498b0fd0423fa1573412c9aa509c958f57e5c93aa4ea523948342de3ae5e851e332afd092c48f826649d1818fc11efa9a6e7efcde5f9f07b7dba368602a33b166f31eef44c888;
    5'b11001 : xpb = 1024'h61e383c05dfd0a49ea883fbb27286ec55e5234b6e1b643dc733b9cc7a3cc12209b3ab3c173af1491c088191b4794c7862be91ba9571f2b1438108982707fcc5fa7c7cac8b0f193f36d8864814cc55351abbc5bedd654be823c7b857561fc6d9b8cd7bd9d7738bc04c74b800e9a025afe17a8246afcd2a05b459b10ec66ddc85c;
    5'b11010 : xpb = 1024'h9e57430c76d881fdc43d87596128381a8666c734394a3c7c253cf2d691b65eb3d5b0683785cca44a5764056641483109be56f655ead483efcefc7a53e3fb74c53a1c5464c73e1e1d821b4aa605e057fe33e43498ce6e971c2713d83af36616a7974931696ce1b6ea93fc919e3726565d27986d3291451682d9cf2eb9de76c830;
    5'b11011 : xpb = 1024'h2a1dbd02cdc5c4e8d2ed57208acdba1e3d055680bb6694a459618f8fcc9dfe3f0cdd9f34cdc3b5744ee1b26a579d89c2ecaaa91c5bd70c7fb5492bc71ca4a8795821a9522df9ab0284142e28261f9879c80713ab3a0242a55c1f9905caa51d2172b3130bb1c1b942d9edbc4edc7a2b92e8aed717d56c2f7a2793d182cd2d6199;
    5'b11100 : xpb = 1024'h66917c4ee6a13c9caca29ebec4cd83736519e8fe12fa8d440b62e59eba884ad2475353aadfe1452ce5bd9eb55150f3467f1883c8ef8c655b4c351c98902050deea7632ee4446352c98a7144cdf3a9d26502eec56321c1b3f46b7ebcb5c0ec62d7d2486d7a76ab428a69ecdde799e26f1f89f1fdf69dea5a1bbc7ef5044c6616d;
    5'b11101 : xpb = 1024'ha3053b9aff7cb4508657e65cfecd4cc88d2e7b7b6a8e85e3bd643bada872976581c90820f1fed4e57c998b004b045cca11865e758341be36e3210d6a039bf9447ccabc8a5a92bf56ad39fa719855a1d2d856c5012a35f3d931503e90ed786f398795faa39d13af0e734fdf6e16c22251088f68a6fe511bc94ffc0d1dbc5f6141;
    5'b11110 : xpb = 1024'h2ecbb5915669f73b9507b6242872cecc43cd0ac7ecaade0bf188d866e35a36f0b8f63f1e39f5e60f741738046159b5833fda113bf44446c6c96dbedd3c452cf89ad01177c14e4c3baf32ddf3b894e24e6c79a41395c99f62665bff5bc4b775b362ffdc45e1f3b166b9410a1ebc15f786c9a5d28c427834c09dc0afe6ab15faaa;
    5'b11111 : xpb = 1024'h6b3f74dd6f456eef6ebcfdc2627298216be19d45443ed6aba38a2e75d1448383f36bf3944c1375c80af3244f5b0d1f06d247ebe887f99fa26059afaeafc0d55e2d249b13d79ad665c3c5c41871afe6faf4a17cbe8de377fc50f4522156211ebf6d715011d79cac4c85f21bae5939f2e5d9961b53d6eaaae831f4cdb422aefa7e;
    endcase
end

endmodule

module compressor_array_236_72_1280
(
    input  [235:0] col_in_0,
    input  [235:0] col_in_1,
    input  [235:0] col_in_2,
    input  [235:0] col_in_3,
    input  [235:0] col_in_4,
    input  [235:0] col_in_5,
    input  [235:0] col_in_6,
    input  [235:0] col_in_7,
    input  [235:0] col_in_8,
    input  [235:0] col_in_9,
    input  [235:0] col_in_10,
    input  [235:0] col_in_11,
    input  [235:0] col_in_12,
    input  [235:0] col_in_13,
    input  [235:0] col_in_14,
    input  [235:0] col_in_15,
    input  [235:0] col_in_16,
    input  [235:0] col_in_17,
    input  [235:0] col_in_18,
    input  [235:0] col_in_19,
    input  [235:0] col_in_20,
    input  [235:0] col_in_21,
    input  [235:0] col_in_22,
    input  [235:0] col_in_23,
    input  [235:0] col_in_24,
    input  [235:0] col_in_25,
    input  [235:0] col_in_26,
    input  [235:0] col_in_27,
    input  [235:0] col_in_28,
    input  [235:0] col_in_29,
    input  [235:0] col_in_30,
    input  [235:0] col_in_31,
    input  [235:0] col_in_32,
    input  [235:0] col_in_33,
    input  [235:0] col_in_34,
    input  [235:0] col_in_35,
    input  [235:0] col_in_36,
    input  [235:0] col_in_37,
    input  [235:0] col_in_38,
    input  [235:0] col_in_39,
    input  [235:0] col_in_40,
    input  [235:0] col_in_41,
    input  [235:0] col_in_42,
    input  [235:0] col_in_43,
    input  [235:0] col_in_44,
    input  [235:0] col_in_45,
    input  [235:0] col_in_46,
    input  [235:0] col_in_47,
    input  [235:0] col_in_48,
    input  [235:0] col_in_49,
    input  [235:0] col_in_50,
    input  [235:0] col_in_51,
    input  [235:0] col_in_52,
    input  [235:0] col_in_53,
    input  [235:0] col_in_54,
    input  [235:0] col_in_55,
    input  [235:0] col_in_56,
    input  [235:0] col_in_57,
    input  [235:0] col_in_58,
    input  [235:0] col_in_59,
    input  [235:0] col_in_60,
    input  [235:0] col_in_61,
    input  [235:0] col_in_62,
    input  [235:0] col_in_63,
    input  [235:0] col_in_64,
    input  [235:0] col_in_65,
    input  [235:0] col_in_66,
    input  [235:0] col_in_67,
    input  [235:0] col_in_68,
    input  [235:0] col_in_69,
    input  [235:0] col_in_70,
    input  [235:0] col_in_71,
    input  [235:0] col_in_72,
    input  [235:0] col_in_73,
    input  [235:0] col_in_74,
    input  [235:0] col_in_75,
    input  [235:0] col_in_76,
    input  [235:0] col_in_77,
    input  [235:0] col_in_78,
    input  [235:0] col_in_79,
    input  [235:0] col_in_80,
    input  [235:0] col_in_81,
    input  [235:0] col_in_82,
    input  [235:0] col_in_83,
    input  [235:0] col_in_84,
    input  [235:0] col_in_85,
    input  [235:0] col_in_86,
    input  [235:0] col_in_87,
    input  [235:0] col_in_88,
    input  [235:0] col_in_89,
    input  [235:0] col_in_90,
    input  [235:0] col_in_91,
    input  [235:0] col_in_92,
    input  [235:0] col_in_93,
    input  [235:0] col_in_94,
    input  [235:0] col_in_95,
    input  [235:0] col_in_96,
    input  [235:0] col_in_97,
    input  [235:0] col_in_98,
    input  [235:0] col_in_99,
    input  [235:0] col_in_100,
    input  [235:0] col_in_101,
    input  [235:0] col_in_102,
    input  [235:0] col_in_103,
    input  [235:0] col_in_104,
    input  [235:0] col_in_105,
    input  [235:0] col_in_106,
    input  [235:0] col_in_107,
    input  [235:0] col_in_108,
    input  [235:0] col_in_109,
    input  [235:0] col_in_110,
    input  [235:0] col_in_111,
    input  [235:0] col_in_112,
    input  [235:0] col_in_113,
    input  [235:0] col_in_114,
    input  [235:0] col_in_115,
    input  [235:0] col_in_116,
    input  [235:0] col_in_117,
    input  [235:0] col_in_118,
    input  [235:0] col_in_119,
    input  [235:0] col_in_120,
    input  [235:0] col_in_121,
    input  [235:0] col_in_122,
    input  [235:0] col_in_123,
    input  [235:0] col_in_124,
    input  [235:0] col_in_125,
    input  [235:0] col_in_126,
    input  [235:0] col_in_127,
    input  [235:0] col_in_128,
    input  [235:0] col_in_129,
    input  [235:0] col_in_130,
    input  [235:0] col_in_131,
    input  [235:0] col_in_132,
    input  [235:0] col_in_133,
    input  [235:0] col_in_134,
    input  [235:0] col_in_135,
    input  [235:0] col_in_136,
    input  [235:0] col_in_137,
    input  [235:0] col_in_138,
    input  [235:0] col_in_139,
    input  [235:0] col_in_140,
    input  [235:0] col_in_141,
    input  [235:0] col_in_142,
    input  [235:0] col_in_143,
    input  [235:0] col_in_144,
    input  [235:0] col_in_145,
    input  [235:0] col_in_146,
    input  [235:0] col_in_147,
    input  [235:0] col_in_148,
    input  [235:0] col_in_149,
    input  [235:0] col_in_150,
    input  [235:0] col_in_151,
    input  [235:0] col_in_152,
    input  [235:0] col_in_153,
    input  [235:0] col_in_154,
    input  [235:0] col_in_155,
    input  [235:0] col_in_156,
    input  [235:0] col_in_157,
    input  [235:0] col_in_158,
    input  [235:0] col_in_159,
    input  [235:0] col_in_160,
    input  [235:0] col_in_161,
    input  [235:0] col_in_162,
    input  [235:0] col_in_163,
    input  [235:0] col_in_164,
    input  [235:0] col_in_165,
    input  [235:0] col_in_166,
    input  [235:0] col_in_167,
    input  [235:0] col_in_168,
    input  [235:0] col_in_169,
    input  [235:0] col_in_170,
    input  [235:0] col_in_171,
    input  [235:0] col_in_172,
    input  [235:0] col_in_173,
    input  [235:0] col_in_174,
    input  [235:0] col_in_175,
    input  [235:0] col_in_176,
    input  [235:0] col_in_177,
    input  [235:0] col_in_178,
    input  [235:0] col_in_179,
    input  [235:0] col_in_180,
    input  [235:0] col_in_181,
    input  [235:0] col_in_182,
    input  [235:0] col_in_183,
    input  [235:0] col_in_184,
    input  [235:0] col_in_185,
    input  [235:0] col_in_186,
    input  [235:0] col_in_187,
    input  [235:0] col_in_188,
    input  [235:0] col_in_189,
    input  [235:0] col_in_190,
    input  [235:0] col_in_191,
    input  [235:0] col_in_192,
    input  [235:0] col_in_193,
    input  [235:0] col_in_194,
    input  [235:0] col_in_195,
    input  [235:0] col_in_196,
    input  [235:0] col_in_197,
    input  [235:0] col_in_198,
    input  [235:0] col_in_199,
    input  [235:0] col_in_200,
    input  [235:0] col_in_201,
    input  [235:0] col_in_202,
    input  [235:0] col_in_203,
    input  [235:0] col_in_204,
    input  [235:0] col_in_205,
    input  [235:0] col_in_206,
    input  [235:0] col_in_207,
    input  [235:0] col_in_208,
    input  [235:0] col_in_209,
    input  [235:0] col_in_210,
    input  [235:0] col_in_211,
    input  [235:0] col_in_212,
    input  [235:0] col_in_213,
    input  [235:0] col_in_214,
    input  [235:0] col_in_215,
    input  [235:0] col_in_216,
    input  [235:0] col_in_217,
    input  [235:0] col_in_218,
    input  [235:0] col_in_219,
    input  [235:0] col_in_220,
    input  [235:0] col_in_221,
    input  [235:0] col_in_222,
    input  [235:0] col_in_223,
    input  [235:0] col_in_224,
    input  [235:0] col_in_225,
    input  [235:0] col_in_226,
    input  [235:0] col_in_227,
    input  [235:0] col_in_228,
    input  [235:0] col_in_229,
    input  [235:0] col_in_230,
    input  [235:0] col_in_231,
    input  [235:0] col_in_232,
    input  [235:0] col_in_233,
    input  [235:0] col_in_234,
    input  [235:0] col_in_235,
    input  [235:0] col_in_236,
    input  [235:0] col_in_237,
    input  [235:0] col_in_238,
    input  [235:0] col_in_239,
    input  [235:0] col_in_240,
    input  [235:0] col_in_241,
    input  [235:0] col_in_242,
    input  [235:0] col_in_243,
    input  [235:0] col_in_244,
    input  [235:0] col_in_245,
    input  [235:0] col_in_246,
    input  [235:0] col_in_247,
    input  [235:0] col_in_248,
    input  [235:0] col_in_249,
    input  [235:0] col_in_250,
    input  [235:0] col_in_251,
    input  [235:0] col_in_252,
    input  [235:0] col_in_253,
    input  [235:0] col_in_254,
    input  [235:0] col_in_255,
    input  [235:0] col_in_256,
    input  [235:0] col_in_257,
    input  [235:0] col_in_258,
    input  [235:0] col_in_259,
    input  [235:0] col_in_260,
    input  [235:0] col_in_261,
    input  [235:0] col_in_262,
    input  [235:0] col_in_263,
    input  [235:0] col_in_264,
    input  [235:0] col_in_265,
    input  [235:0] col_in_266,
    input  [235:0] col_in_267,
    input  [235:0] col_in_268,
    input  [235:0] col_in_269,
    input  [235:0] col_in_270,
    input  [235:0] col_in_271,
    input  [235:0] col_in_272,
    input  [235:0] col_in_273,
    input  [235:0] col_in_274,
    input  [235:0] col_in_275,
    input  [235:0] col_in_276,
    input  [235:0] col_in_277,
    input  [235:0] col_in_278,
    input  [235:0] col_in_279,
    input  [235:0] col_in_280,
    input  [235:0] col_in_281,
    input  [235:0] col_in_282,
    input  [235:0] col_in_283,
    input  [235:0] col_in_284,
    input  [235:0] col_in_285,
    input  [235:0] col_in_286,
    input  [235:0] col_in_287,
    input  [235:0] col_in_288,
    input  [235:0] col_in_289,
    input  [235:0] col_in_290,
    input  [235:0] col_in_291,
    input  [235:0] col_in_292,
    input  [235:0] col_in_293,
    input  [235:0] col_in_294,
    input  [235:0] col_in_295,
    input  [235:0] col_in_296,
    input  [235:0] col_in_297,
    input  [235:0] col_in_298,
    input  [235:0] col_in_299,
    input  [235:0] col_in_300,
    input  [235:0] col_in_301,
    input  [235:0] col_in_302,
    input  [235:0] col_in_303,
    input  [235:0] col_in_304,
    input  [235:0] col_in_305,
    input  [235:0] col_in_306,
    input  [235:0] col_in_307,
    input  [235:0] col_in_308,
    input  [235:0] col_in_309,
    input  [235:0] col_in_310,
    input  [235:0] col_in_311,
    input  [235:0] col_in_312,
    input  [235:0] col_in_313,
    input  [235:0] col_in_314,
    input  [235:0] col_in_315,
    input  [235:0] col_in_316,
    input  [235:0] col_in_317,
    input  [235:0] col_in_318,
    input  [235:0] col_in_319,
    input  [235:0] col_in_320,
    input  [235:0] col_in_321,
    input  [235:0] col_in_322,
    input  [235:0] col_in_323,
    input  [235:0] col_in_324,
    input  [235:0] col_in_325,
    input  [235:0] col_in_326,
    input  [235:0] col_in_327,
    input  [235:0] col_in_328,
    input  [235:0] col_in_329,
    input  [235:0] col_in_330,
    input  [235:0] col_in_331,
    input  [235:0] col_in_332,
    input  [235:0] col_in_333,
    input  [235:0] col_in_334,
    input  [235:0] col_in_335,
    input  [235:0] col_in_336,
    input  [235:0] col_in_337,
    input  [235:0] col_in_338,
    input  [235:0] col_in_339,
    input  [235:0] col_in_340,
    input  [235:0] col_in_341,
    input  [235:0] col_in_342,
    input  [235:0] col_in_343,
    input  [235:0] col_in_344,
    input  [235:0] col_in_345,
    input  [235:0] col_in_346,
    input  [235:0] col_in_347,
    input  [235:0] col_in_348,
    input  [235:0] col_in_349,
    input  [235:0] col_in_350,
    input  [235:0] col_in_351,
    input  [235:0] col_in_352,
    input  [235:0] col_in_353,
    input  [235:0] col_in_354,
    input  [235:0] col_in_355,
    input  [235:0] col_in_356,
    input  [235:0] col_in_357,
    input  [235:0] col_in_358,
    input  [235:0] col_in_359,
    input  [235:0] col_in_360,
    input  [235:0] col_in_361,
    input  [235:0] col_in_362,
    input  [235:0] col_in_363,
    input  [235:0] col_in_364,
    input  [235:0] col_in_365,
    input  [235:0] col_in_366,
    input  [235:0] col_in_367,
    input  [235:0] col_in_368,
    input  [235:0] col_in_369,
    input  [235:0] col_in_370,
    input  [235:0] col_in_371,
    input  [235:0] col_in_372,
    input  [235:0] col_in_373,
    input  [235:0] col_in_374,
    input  [235:0] col_in_375,
    input  [235:0] col_in_376,
    input  [235:0] col_in_377,
    input  [235:0] col_in_378,
    input  [235:0] col_in_379,
    input  [235:0] col_in_380,
    input  [235:0] col_in_381,
    input  [235:0] col_in_382,
    input  [235:0] col_in_383,
    input  [235:0] col_in_384,
    input  [235:0] col_in_385,
    input  [235:0] col_in_386,
    input  [235:0] col_in_387,
    input  [235:0] col_in_388,
    input  [235:0] col_in_389,
    input  [235:0] col_in_390,
    input  [235:0] col_in_391,
    input  [235:0] col_in_392,
    input  [235:0] col_in_393,
    input  [235:0] col_in_394,
    input  [235:0] col_in_395,
    input  [235:0] col_in_396,
    input  [235:0] col_in_397,
    input  [235:0] col_in_398,
    input  [235:0] col_in_399,
    input  [235:0] col_in_400,
    input  [235:0] col_in_401,
    input  [235:0] col_in_402,
    input  [235:0] col_in_403,
    input  [235:0] col_in_404,
    input  [235:0] col_in_405,
    input  [235:0] col_in_406,
    input  [235:0] col_in_407,
    input  [235:0] col_in_408,
    input  [235:0] col_in_409,
    input  [235:0] col_in_410,
    input  [235:0] col_in_411,
    input  [235:0] col_in_412,
    input  [235:0] col_in_413,
    input  [235:0] col_in_414,
    input  [235:0] col_in_415,
    input  [235:0] col_in_416,
    input  [235:0] col_in_417,
    input  [235:0] col_in_418,
    input  [235:0] col_in_419,
    input  [235:0] col_in_420,
    input  [235:0] col_in_421,
    input  [235:0] col_in_422,
    input  [235:0] col_in_423,
    input  [235:0] col_in_424,
    input  [235:0] col_in_425,
    input  [235:0] col_in_426,
    input  [235:0] col_in_427,
    input  [235:0] col_in_428,
    input  [235:0] col_in_429,
    input  [235:0] col_in_430,
    input  [235:0] col_in_431,
    input  [235:0] col_in_432,
    input  [235:0] col_in_433,
    input  [235:0] col_in_434,
    input  [235:0] col_in_435,
    input  [235:0] col_in_436,
    input  [235:0] col_in_437,
    input  [235:0] col_in_438,
    input  [235:0] col_in_439,
    input  [235:0] col_in_440,
    input  [235:0] col_in_441,
    input  [235:0] col_in_442,
    input  [235:0] col_in_443,
    input  [235:0] col_in_444,
    input  [235:0] col_in_445,
    input  [235:0] col_in_446,
    input  [235:0] col_in_447,
    input  [235:0] col_in_448,
    input  [235:0] col_in_449,
    input  [235:0] col_in_450,
    input  [235:0] col_in_451,
    input  [235:0] col_in_452,
    input  [235:0] col_in_453,
    input  [235:0] col_in_454,
    input  [235:0] col_in_455,
    input  [235:0] col_in_456,
    input  [235:0] col_in_457,
    input  [235:0] col_in_458,
    input  [235:0] col_in_459,
    input  [235:0] col_in_460,
    input  [235:0] col_in_461,
    input  [235:0] col_in_462,
    input  [235:0] col_in_463,
    input  [235:0] col_in_464,
    input  [235:0] col_in_465,
    input  [235:0] col_in_466,
    input  [235:0] col_in_467,
    input  [235:0] col_in_468,
    input  [235:0] col_in_469,
    input  [235:0] col_in_470,
    input  [235:0] col_in_471,
    input  [235:0] col_in_472,
    input  [235:0] col_in_473,
    input  [235:0] col_in_474,
    input  [235:0] col_in_475,
    input  [235:0] col_in_476,
    input  [235:0] col_in_477,
    input  [235:0] col_in_478,
    input  [235:0] col_in_479,
    input  [235:0] col_in_480,
    input  [235:0] col_in_481,
    input  [235:0] col_in_482,
    input  [235:0] col_in_483,
    input  [235:0] col_in_484,
    input  [235:0] col_in_485,
    input  [235:0] col_in_486,
    input  [235:0] col_in_487,
    input  [235:0] col_in_488,
    input  [235:0] col_in_489,
    input  [235:0] col_in_490,
    input  [235:0] col_in_491,
    input  [235:0] col_in_492,
    input  [235:0] col_in_493,
    input  [235:0] col_in_494,
    input  [235:0] col_in_495,
    input  [235:0] col_in_496,
    input  [235:0] col_in_497,
    input  [235:0] col_in_498,
    input  [235:0] col_in_499,
    input  [235:0] col_in_500,
    input  [235:0] col_in_501,
    input  [235:0] col_in_502,
    input  [235:0] col_in_503,
    input  [235:0] col_in_504,
    input  [235:0] col_in_505,
    input  [235:0] col_in_506,
    input  [235:0] col_in_507,
    input  [235:0] col_in_508,
    input  [235:0] col_in_509,
    input  [235:0] col_in_510,
    input  [235:0] col_in_511,
    input  [235:0] col_in_512,
    input  [235:0] col_in_513,
    input  [235:0] col_in_514,
    input  [235:0] col_in_515,
    input  [235:0] col_in_516,
    input  [235:0] col_in_517,
    input  [235:0] col_in_518,
    input  [235:0] col_in_519,
    input  [235:0] col_in_520,
    input  [235:0] col_in_521,
    input  [235:0] col_in_522,
    input  [235:0] col_in_523,
    input  [235:0] col_in_524,
    input  [235:0] col_in_525,
    input  [235:0] col_in_526,
    input  [235:0] col_in_527,
    input  [235:0] col_in_528,
    input  [235:0] col_in_529,
    input  [235:0] col_in_530,
    input  [235:0] col_in_531,
    input  [235:0] col_in_532,
    input  [235:0] col_in_533,
    input  [235:0] col_in_534,
    input  [235:0] col_in_535,
    input  [235:0] col_in_536,
    input  [235:0] col_in_537,
    input  [235:0] col_in_538,
    input  [235:0] col_in_539,
    input  [235:0] col_in_540,
    input  [235:0] col_in_541,
    input  [235:0] col_in_542,
    input  [235:0] col_in_543,
    input  [235:0] col_in_544,
    input  [235:0] col_in_545,
    input  [235:0] col_in_546,
    input  [235:0] col_in_547,
    input  [235:0] col_in_548,
    input  [235:0] col_in_549,
    input  [235:0] col_in_550,
    input  [235:0] col_in_551,
    input  [235:0] col_in_552,
    input  [235:0] col_in_553,
    input  [235:0] col_in_554,
    input  [235:0] col_in_555,
    input  [235:0] col_in_556,
    input  [235:0] col_in_557,
    input  [235:0] col_in_558,
    input  [235:0] col_in_559,
    input  [235:0] col_in_560,
    input  [235:0] col_in_561,
    input  [235:0] col_in_562,
    input  [235:0] col_in_563,
    input  [235:0] col_in_564,
    input  [235:0] col_in_565,
    input  [235:0] col_in_566,
    input  [235:0] col_in_567,
    input  [235:0] col_in_568,
    input  [235:0] col_in_569,
    input  [235:0] col_in_570,
    input  [235:0] col_in_571,
    input  [235:0] col_in_572,
    input  [235:0] col_in_573,
    input  [235:0] col_in_574,
    input  [235:0] col_in_575,
    input  [235:0] col_in_576,
    input  [235:0] col_in_577,
    input  [235:0] col_in_578,
    input  [235:0] col_in_579,
    input  [235:0] col_in_580,
    input  [235:0] col_in_581,
    input  [235:0] col_in_582,
    input  [235:0] col_in_583,
    input  [235:0] col_in_584,
    input  [235:0] col_in_585,
    input  [235:0] col_in_586,
    input  [235:0] col_in_587,
    input  [235:0] col_in_588,
    input  [235:0] col_in_589,
    input  [235:0] col_in_590,
    input  [235:0] col_in_591,
    input  [235:0] col_in_592,
    input  [235:0] col_in_593,
    input  [235:0] col_in_594,
    input  [235:0] col_in_595,
    input  [235:0] col_in_596,
    input  [235:0] col_in_597,
    input  [235:0] col_in_598,
    input  [235:0] col_in_599,
    input  [235:0] col_in_600,
    input  [235:0] col_in_601,
    input  [235:0] col_in_602,
    input  [235:0] col_in_603,
    input  [235:0] col_in_604,
    input  [235:0] col_in_605,
    input  [235:0] col_in_606,
    input  [235:0] col_in_607,
    input  [235:0] col_in_608,
    input  [235:0] col_in_609,
    input  [235:0] col_in_610,
    input  [235:0] col_in_611,
    input  [235:0] col_in_612,
    input  [235:0] col_in_613,
    input  [235:0] col_in_614,
    input  [235:0] col_in_615,
    input  [235:0] col_in_616,
    input  [235:0] col_in_617,
    input  [235:0] col_in_618,
    input  [235:0] col_in_619,
    input  [235:0] col_in_620,
    input  [235:0] col_in_621,
    input  [235:0] col_in_622,
    input  [235:0] col_in_623,
    input  [235:0] col_in_624,
    input  [235:0] col_in_625,
    input  [235:0] col_in_626,
    input  [235:0] col_in_627,
    input  [235:0] col_in_628,
    input  [235:0] col_in_629,
    input  [235:0] col_in_630,
    input  [235:0] col_in_631,
    input  [235:0] col_in_632,
    input  [235:0] col_in_633,
    input  [235:0] col_in_634,
    input  [235:0] col_in_635,
    input  [235:0] col_in_636,
    input  [235:0] col_in_637,
    input  [235:0] col_in_638,
    input  [235:0] col_in_639,
    input  [235:0] col_in_640,
    input  [235:0] col_in_641,
    input  [235:0] col_in_642,
    input  [235:0] col_in_643,
    input  [235:0] col_in_644,
    input  [235:0] col_in_645,
    input  [235:0] col_in_646,
    input  [235:0] col_in_647,
    input  [235:0] col_in_648,
    input  [235:0] col_in_649,
    input  [235:0] col_in_650,
    input  [235:0] col_in_651,
    input  [235:0] col_in_652,
    input  [235:0] col_in_653,
    input  [235:0] col_in_654,
    input  [235:0] col_in_655,
    input  [235:0] col_in_656,
    input  [235:0] col_in_657,
    input  [235:0] col_in_658,
    input  [235:0] col_in_659,
    input  [235:0] col_in_660,
    input  [235:0] col_in_661,
    input  [235:0] col_in_662,
    input  [235:0] col_in_663,
    input  [235:0] col_in_664,
    input  [235:0] col_in_665,
    input  [235:0] col_in_666,
    input  [235:0] col_in_667,
    input  [235:0] col_in_668,
    input  [235:0] col_in_669,
    input  [235:0] col_in_670,
    input  [235:0] col_in_671,
    input  [235:0] col_in_672,
    input  [235:0] col_in_673,
    input  [235:0] col_in_674,
    input  [235:0] col_in_675,
    input  [235:0] col_in_676,
    input  [235:0] col_in_677,
    input  [235:0] col_in_678,
    input  [235:0] col_in_679,
    input  [235:0] col_in_680,
    input  [235:0] col_in_681,
    input  [235:0] col_in_682,
    input  [235:0] col_in_683,
    input  [235:0] col_in_684,
    input  [235:0] col_in_685,
    input  [235:0] col_in_686,
    input  [235:0] col_in_687,
    input  [235:0] col_in_688,
    input  [235:0] col_in_689,
    input  [235:0] col_in_690,
    input  [235:0] col_in_691,
    input  [235:0] col_in_692,
    input  [235:0] col_in_693,
    input  [235:0] col_in_694,
    input  [235:0] col_in_695,
    input  [235:0] col_in_696,
    input  [235:0] col_in_697,
    input  [235:0] col_in_698,
    input  [235:0] col_in_699,
    input  [235:0] col_in_700,
    input  [235:0] col_in_701,
    input  [235:0] col_in_702,
    input  [235:0] col_in_703,
    input  [235:0] col_in_704,
    input  [235:0] col_in_705,
    input  [235:0] col_in_706,
    input  [235:0] col_in_707,
    input  [235:0] col_in_708,
    input  [235:0] col_in_709,
    input  [235:0] col_in_710,
    input  [235:0] col_in_711,
    input  [235:0] col_in_712,
    input  [235:0] col_in_713,
    input  [235:0] col_in_714,
    input  [235:0] col_in_715,
    input  [235:0] col_in_716,
    input  [235:0] col_in_717,
    input  [235:0] col_in_718,
    input  [235:0] col_in_719,
    input  [235:0] col_in_720,
    input  [235:0] col_in_721,
    input  [235:0] col_in_722,
    input  [235:0] col_in_723,
    input  [235:0] col_in_724,
    input  [235:0] col_in_725,
    input  [235:0] col_in_726,
    input  [235:0] col_in_727,
    input  [235:0] col_in_728,
    input  [235:0] col_in_729,
    input  [235:0] col_in_730,
    input  [235:0] col_in_731,
    input  [235:0] col_in_732,
    input  [235:0] col_in_733,
    input  [235:0] col_in_734,
    input  [235:0] col_in_735,
    input  [235:0] col_in_736,
    input  [235:0] col_in_737,
    input  [235:0] col_in_738,
    input  [235:0] col_in_739,
    input  [235:0] col_in_740,
    input  [235:0] col_in_741,
    input  [235:0] col_in_742,
    input  [235:0] col_in_743,
    input  [235:0] col_in_744,
    input  [235:0] col_in_745,
    input  [235:0] col_in_746,
    input  [235:0] col_in_747,
    input  [235:0] col_in_748,
    input  [235:0] col_in_749,
    input  [235:0] col_in_750,
    input  [235:0] col_in_751,
    input  [235:0] col_in_752,
    input  [235:0] col_in_753,
    input  [235:0] col_in_754,
    input  [235:0] col_in_755,
    input  [235:0] col_in_756,
    input  [235:0] col_in_757,
    input  [235:0] col_in_758,
    input  [235:0] col_in_759,
    input  [235:0] col_in_760,
    input  [235:0] col_in_761,
    input  [235:0] col_in_762,
    input  [235:0] col_in_763,
    input  [235:0] col_in_764,
    input  [235:0] col_in_765,
    input  [235:0] col_in_766,
    input  [235:0] col_in_767,
    input  [235:0] col_in_768,
    input  [235:0] col_in_769,
    input  [235:0] col_in_770,
    input  [235:0] col_in_771,
    input  [235:0] col_in_772,
    input  [235:0] col_in_773,
    input  [235:0] col_in_774,
    input  [235:0] col_in_775,
    input  [235:0] col_in_776,
    input  [235:0] col_in_777,
    input  [235:0] col_in_778,
    input  [235:0] col_in_779,
    input  [235:0] col_in_780,
    input  [235:0] col_in_781,
    input  [235:0] col_in_782,
    input  [235:0] col_in_783,
    input  [235:0] col_in_784,
    input  [235:0] col_in_785,
    input  [235:0] col_in_786,
    input  [235:0] col_in_787,
    input  [235:0] col_in_788,
    input  [235:0] col_in_789,
    input  [235:0] col_in_790,
    input  [235:0] col_in_791,
    input  [235:0] col_in_792,
    input  [235:0] col_in_793,
    input  [235:0] col_in_794,
    input  [235:0] col_in_795,
    input  [235:0] col_in_796,
    input  [235:0] col_in_797,
    input  [235:0] col_in_798,
    input  [235:0] col_in_799,
    input  [235:0] col_in_800,
    input  [235:0] col_in_801,
    input  [235:0] col_in_802,
    input  [235:0] col_in_803,
    input  [235:0] col_in_804,
    input  [235:0] col_in_805,
    input  [235:0] col_in_806,
    input  [235:0] col_in_807,
    input  [235:0] col_in_808,
    input  [235:0] col_in_809,
    input  [235:0] col_in_810,
    input  [235:0] col_in_811,
    input  [235:0] col_in_812,
    input  [235:0] col_in_813,
    input  [235:0] col_in_814,
    input  [235:0] col_in_815,
    input  [235:0] col_in_816,
    input  [235:0] col_in_817,
    input  [235:0] col_in_818,
    input  [235:0] col_in_819,
    input  [235:0] col_in_820,
    input  [235:0] col_in_821,
    input  [235:0] col_in_822,
    input  [235:0] col_in_823,
    input  [235:0] col_in_824,
    input  [235:0] col_in_825,
    input  [235:0] col_in_826,
    input  [235:0] col_in_827,
    input  [235:0] col_in_828,
    input  [235:0] col_in_829,
    input  [235:0] col_in_830,
    input  [235:0] col_in_831,
    input  [235:0] col_in_832,
    input  [235:0] col_in_833,
    input  [235:0] col_in_834,
    input  [235:0] col_in_835,
    input  [235:0] col_in_836,
    input  [235:0] col_in_837,
    input  [235:0] col_in_838,
    input  [235:0] col_in_839,
    input  [235:0] col_in_840,
    input  [235:0] col_in_841,
    input  [235:0] col_in_842,
    input  [235:0] col_in_843,
    input  [235:0] col_in_844,
    input  [235:0] col_in_845,
    input  [235:0] col_in_846,
    input  [235:0] col_in_847,
    input  [235:0] col_in_848,
    input  [235:0] col_in_849,
    input  [235:0] col_in_850,
    input  [235:0] col_in_851,
    input  [235:0] col_in_852,
    input  [235:0] col_in_853,
    input  [235:0] col_in_854,
    input  [235:0] col_in_855,
    input  [235:0] col_in_856,
    input  [235:0] col_in_857,
    input  [235:0] col_in_858,
    input  [235:0] col_in_859,
    input  [235:0] col_in_860,
    input  [235:0] col_in_861,
    input  [235:0] col_in_862,
    input  [235:0] col_in_863,
    input  [235:0] col_in_864,
    input  [235:0] col_in_865,
    input  [235:0] col_in_866,
    input  [235:0] col_in_867,
    input  [235:0] col_in_868,
    input  [235:0] col_in_869,
    input  [235:0] col_in_870,
    input  [235:0] col_in_871,
    input  [235:0] col_in_872,
    input  [235:0] col_in_873,
    input  [235:0] col_in_874,
    input  [235:0] col_in_875,
    input  [235:0] col_in_876,
    input  [235:0] col_in_877,
    input  [235:0] col_in_878,
    input  [235:0] col_in_879,
    input  [235:0] col_in_880,
    input  [235:0] col_in_881,
    input  [235:0] col_in_882,
    input  [235:0] col_in_883,
    input  [235:0] col_in_884,
    input  [235:0] col_in_885,
    input  [235:0] col_in_886,
    input  [235:0] col_in_887,
    input  [235:0] col_in_888,
    input  [235:0] col_in_889,
    input  [235:0] col_in_890,
    input  [235:0] col_in_891,
    input  [235:0] col_in_892,
    input  [235:0] col_in_893,
    input  [235:0] col_in_894,
    input  [235:0] col_in_895,
    input  [235:0] col_in_896,
    input  [235:0] col_in_897,
    input  [235:0] col_in_898,
    input  [235:0] col_in_899,
    input  [235:0] col_in_900,
    input  [235:0] col_in_901,
    input  [235:0] col_in_902,
    input  [235:0] col_in_903,
    input  [235:0] col_in_904,
    input  [235:0] col_in_905,
    input  [235:0] col_in_906,
    input  [235:0] col_in_907,
    input  [235:0] col_in_908,
    input  [235:0] col_in_909,
    input  [235:0] col_in_910,
    input  [235:0] col_in_911,
    input  [235:0] col_in_912,
    input  [235:0] col_in_913,
    input  [235:0] col_in_914,
    input  [235:0] col_in_915,
    input  [235:0] col_in_916,
    input  [235:0] col_in_917,
    input  [235:0] col_in_918,
    input  [235:0] col_in_919,
    input  [235:0] col_in_920,
    input  [235:0] col_in_921,
    input  [235:0] col_in_922,
    input  [235:0] col_in_923,
    input  [235:0] col_in_924,
    input  [235:0] col_in_925,
    input  [235:0] col_in_926,
    input  [235:0] col_in_927,
    input  [235:0] col_in_928,
    input  [235:0] col_in_929,
    input  [235:0] col_in_930,
    input  [235:0] col_in_931,
    input  [235:0] col_in_932,
    input  [235:0] col_in_933,
    input  [235:0] col_in_934,
    input  [235:0] col_in_935,
    input  [235:0] col_in_936,
    input  [235:0] col_in_937,
    input  [235:0] col_in_938,
    input  [235:0] col_in_939,
    input  [235:0] col_in_940,
    input  [235:0] col_in_941,
    input  [235:0] col_in_942,
    input  [235:0] col_in_943,
    input  [235:0] col_in_944,
    input  [235:0] col_in_945,
    input  [235:0] col_in_946,
    input  [235:0] col_in_947,
    input  [235:0] col_in_948,
    input  [235:0] col_in_949,
    input  [235:0] col_in_950,
    input  [235:0] col_in_951,
    input  [235:0] col_in_952,
    input  [235:0] col_in_953,
    input  [235:0] col_in_954,
    input  [235:0] col_in_955,
    input  [235:0] col_in_956,
    input  [235:0] col_in_957,
    input  [235:0] col_in_958,
    input  [235:0] col_in_959,
    input  [235:0] col_in_960,
    input  [235:0] col_in_961,
    input  [235:0] col_in_962,
    input  [235:0] col_in_963,
    input  [235:0] col_in_964,
    input  [235:0] col_in_965,
    input  [235:0] col_in_966,
    input  [235:0] col_in_967,
    input  [235:0] col_in_968,
    input  [235:0] col_in_969,
    input  [235:0] col_in_970,
    input  [235:0] col_in_971,
    input  [235:0] col_in_972,
    input  [235:0] col_in_973,
    input  [235:0] col_in_974,
    input  [235:0] col_in_975,
    input  [235:0] col_in_976,
    input  [235:0] col_in_977,
    input  [235:0] col_in_978,
    input  [235:0] col_in_979,
    input  [235:0] col_in_980,
    input  [235:0] col_in_981,
    input  [235:0] col_in_982,
    input  [235:0] col_in_983,
    input  [235:0] col_in_984,
    input  [235:0] col_in_985,
    input  [235:0] col_in_986,
    input  [235:0] col_in_987,
    input  [235:0] col_in_988,
    input  [235:0] col_in_989,
    input  [235:0] col_in_990,
    input  [235:0] col_in_991,
    input  [235:0] col_in_992,
    input  [235:0] col_in_993,
    input  [235:0] col_in_994,
    input  [235:0] col_in_995,
    input  [235:0] col_in_996,
    input  [235:0] col_in_997,
    input  [235:0] col_in_998,
    input  [235:0] col_in_999,
    input  [235:0] col_in_1000,
    input  [235:0] col_in_1001,
    input  [235:0] col_in_1002,
    input  [235:0] col_in_1003,
    input  [235:0] col_in_1004,
    input  [235:0] col_in_1005,
    input  [235:0] col_in_1006,
    input  [235:0] col_in_1007,
    input  [235:0] col_in_1008,
    input  [235:0] col_in_1009,
    input  [235:0] col_in_1010,
    input  [235:0] col_in_1011,
    input  [235:0] col_in_1012,
    input  [235:0] col_in_1013,
    input  [235:0] col_in_1014,
    input  [235:0] col_in_1015,
    input  [235:0] col_in_1016,
    input  [235:0] col_in_1017,
    input  [235:0] col_in_1018,
    input  [235:0] col_in_1019,
    input  [235:0] col_in_1020,
    input  [235:0] col_in_1021,
    input  [235:0] col_in_1022,
    input  [235:0] col_in_1023,
    input  [235:0] col_in_1024,
    input  [235:0] col_in_1025,
    input  [235:0] col_in_1026,
    input  [235:0] col_in_1027,
    input  [235:0] col_in_1028,
    input  [235:0] col_in_1029,
    input  [235:0] col_in_1030,
    input  [235:0] col_in_1031,
    input  [235:0] col_in_1032,
    input  [235:0] col_in_1033,
    input  [235:0] col_in_1034,
    input  [235:0] col_in_1035,
    input  [235:0] col_in_1036,
    input  [235:0] col_in_1037,
    input  [235:0] col_in_1038,
    input  [235:0] col_in_1039,
    input  [235:0] col_in_1040,
    input  [235:0] col_in_1041,
    input  [235:0] col_in_1042,
    input  [235:0] col_in_1043,
    input  [235:0] col_in_1044,
    input  [235:0] col_in_1045,
    input  [235:0] col_in_1046,
    input  [235:0] col_in_1047,
    input  [235:0] col_in_1048,
    input  [235:0] col_in_1049,
    input  [235:0] col_in_1050,
    input  [235:0] col_in_1051,
    input  [235:0] col_in_1052,
    input  [235:0] col_in_1053,
    input  [235:0] col_in_1054,
    input  [235:0] col_in_1055,
    input  [235:0] col_in_1056,
    input  [235:0] col_in_1057,
    input  [235:0] col_in_1058,
    input  [235:0] col_in_1059,
    input  [235:0] col_in_1060,
    input  [235:0] col_in_1061,
    input  [235:0] col_in_1062,
    input  [235:0] col_in_1063,
    input  [235:0] col_in_1064,
    input  [235:0] col_in_1065,
    input  [235:0] col_in_1066,
    input  [235:0] col_in_1067,
    input  [235:0] col_in_1068,
    input  [235:0] col_in_1069,
    input  [235:0] col_in_1070,
    input  [235:0] col_in_1071,
    input  [235:0] col_in_1072,
    input  [235:0] col_in_1073,
    input  [235:0] col_in_1074,
    input  [235:0] col_in_1075,
    input  [235:0] col_in_1076,
    input  [235:0] col_in_1077,
    input  [235:0] col_in_1078,
    input  [235:0] col_in_1079,
    input  [235:0] col_in_1080,
    input  [235:0] col_in_1081,
    input  [235:0] col_in_1082,
    input  [235:0] col_in_1083,
    input  [235:0] col_in_1084,
    input  [235:0] col_in_1085,
    input  [235:0] col_in_1086,
    input  [235:0] col_in_1087,
    input  [235:0] col_in_1088,
    input  [235:0] col_in_1089,
    input  [235:0] col_in_1090,
    input  [235:0] col_in_1091,
    input  [235:0] col_in_1092,
    input  [235:0] col_in_1093,
    input  [235:0] col_in_1094,
    input  [235:0] col_in_1095,
    input  [235:0] col_in_1096,
    input  [235:0] col_in_1097,
    input  [235:0] col_in_1098,
    input  [235:0] col_in_1099,
    input  [235:0] col_in_1100,
    input  [235:0] col_in_1101,
    input  [235:0] col_in_1102,
    input  [235:0] col_in_1103,
    input  [235:0] col_in_1104,
    input  [235:0] col_in_1105,
    input  [235:0] col_in_1106,
    input  [235:0] col_in_1107,
    input  [235:0] col_in_1108,
    input  [235:0] col_in_1109,
    input  [235:0] col_in_1110,
    input  [235:0] col_in_1111,
    input  [235:0] col_in_1112,
    input  [235:0] col_in_1113,
    input  [235:0] col_in_1114,
    input  [235:0] col_in_1115,
    input  [235:0] col_in_1116,
    input  [235:0] col_in_1117,
    input  [235:0] col_in_1118,
    input  [235:0] col_in_1119,
    input  [235:0] col_in_1120,
    input  [235:0] col_in_1121,
    input  [235:0] col_in_1122,
    input  [235:0] col_in_1123,
    input  [235:0] col_in_1124,
    input  [235:0] col_in_1125,
    input  [235:0] col_in_1126,
    input  [235:0] col_in_1127,
    input  [235:0] col_in_1128,
    input  [235:0] col_in_1129,
    input  [235:0] col_in_1130,
    input  [235:0] col_in_1131,
    input  [235:0] col_in_1132,
    input  [235:0] col_in_1133,
    input  [235:0] col_in_1134,
    input  [235:0] col_in_1135,
    input  [235:0] col_in_1136,
    input  [235:0] col_in_1137,
    input  [235:0] col_in_1138,
    input  [235:0] col_in_1139,
    input  [235:0] col_in_1140,
    input  [235:0] col_in_1141,
    input  [235:0] col_in_1142,
    input  [235:0] col_in_1143,
    input  [235:0] col_in_1144,
    input  [235:0] col_in_1145,
    input  [235:0] col_in_1146,
    input  [235:0] col_in_1147,
    input  [235:0] col_in_1148,
    input  [235:0] col_in_1149,
    input  [235:0] col_in_1150,
    input  [235:0] col_in_1151,
    input  [235:0] col_in_1152,
    input  [235:0] col_in_1153,
    input  [235:0] col_in_1154,
    input  [235:0] col_in_1155,
    input  [235:0] col_in_1156,
    input  [235:0] col_in_1157,
    input  [235:0] col_in_1158,
    input  [235:0] col_in_1159,
    input  [235:0] col_in_1160,
    input  [235:0] col_in_1161,
    input  [235:0] col_in_1162,
    input  [235:0] col_in_1163,
    input  [235:0] col_in_1164,
    input  [235:0] col_in_1165,
    input  [235:0] col_in_1166,
    input  [235:0] col_in_1167,
    input  [235:0] col_in_1168,
    input  [235:0] col_in_1169,
    input  [235:0] col_in_1170,
    input  [235:0] col_in_1171,
    input  [235:0] col_in_1172,
    input  [235:0] col_in_1173,
    input  [235:0] col_in_1174,
    input  [235:0] col_in_1175,
    input  [235:0] col_in_1176,
    input  [235:0] col_in_1177,
    input  [235:0] col_in_1178,
    input  [235:0] col_in_1179,
    input  [235:0] col_in_1180,
    input  [235:0] col_in_1181,
    input  [235:0] col_in_1182,
    input  [235:0] col_in_1183,
    input  [235:0] col_in_1184,
    input  [235:0] col_in_1185,
    input  [235:0] col_in_1186,
    input  [235:0] col_in_1187,
    input  [235:0] col_in_1188,
    input  [235:0] col_in_1189,
    input  [235:0] col_in_1190,
    input  [235:0] col_in_1191,
    input  [235:0] col_in_1192,
    input  [235:0] col_in_1193,
    input  [235:0] col_in_1194,
    input  [235:0] col_in_1195,
    input  [235:0] col_in_1196,
    input  [235:0] col_in_1197,
    input  [235:0] col_in_1198,
    input  [235:0] col_in_1199,
    input  [235:0] col_in_1200,
    input  [235:0] col_in_1201,
    input  [235:0] col_in_1202,
    input  [235:0] col_in_1203,
    input  [235:0] col_in_1204,
    input  [235:0] col_in_1205,
    input  [235:0] col_in_1206,
    input  [235:0] col_in_1207,
    input  [235:0] col_in_1208,
    input  [235:0] col_in_1209,
    input  [235:0] col_in_1210,
    input  [235:0] col_in_1211,
    input  [235:0] col_in_1212,
    input  [235:0] col_in_1213,
    input  [235:0] col_in_1214,
    input  [235:0] col_in_1215,
    input  [235:0] col_in_1216,
    input  [235:0] col_in_1217,
    input  [235:0] col_in_1218,
    input  [235:0] col_in_1219,
    input  [235:0] col_in_1220,
    input  [235:0] col_in_1221,
    input  [235:0] col_in_1222,
    input  [235:0] col_in_1223,
    input  [235:0] col_in_1224,
    input  [235:0] col_in_1225,
    input  [235:0] col_in_1226,
    input  [235:0] col_in_1227,
    input  [235:0] col_in_1228,
    input  [235:0] col_in_1229,
    input  [235:0] col_in_1230,
    input  [235:0] col_in_1231,
    input  [235:0] col_in_1232,
    input  [235:0] col_in_1233,
    input  [235:0] col_in_1234,
    input  [235:0] col_in_1235,
    input  [235:0] col_in_1236,
    input  [235:0] col_in_1237,
    input  [235:0] col_in_1238,
    input  [235:0] col_in_1239,
    input  [235:0] col_in_1240,
    input  [235:0] col_in_1241,
    input  [235:0] col_in_1242,
    input  [235:0] col_in_1243,
    input  [235:0] col_in_1244,
    input  [235:0] col_in_1245,
    input  [235:0] col_in_1246,
    input  [235:0] col_in_1247,
    input  [235:0] col_in_1248,
    input  [235:0] col_in_1249,
    input  [235:0] col_in_1250,
    input  [235:0] col_in_1251,
    input  [235:0] col_in_1252,
    input  [235:0] col_in_1253,
    input  [235:0] col_in_1254,
    input  [235:0] col_in_1255,
    input  [235:0] col_in_1256,
    input  [235:0] col_in_1257,
    input  [235:0] col_in_1258,
    input  [235:0] col_in_1259,
    input  [235:0] col_in_1260,
    input  [235:0] col_in_1261,
    input  [235:0] col_in_1262,
    input  [235:0] col_in_1263,
    input  [235:0] col_in_1264,
    input  [235:0] col_in_1265,
    input  [235:0] col_in_1266,
    input  [235:0] col_in_1267,
    input  [235:0] col_in_1268,
    input  [235:0] col_in_1269,
    input  [235:0] col_in_1270,
    input  [235:0] col_in_1271,
    input  [235:0] col_in_1272,
    input  [235:0] col_in_1273,
    input  [235:0] col_in_1274,
    input  [235:0] col_in_1275,
    input  [235:0] col_in_1276,
    input  [235:0] col_in_1277,
    input  [235:0] col_in_1278,
    input  [235:0] col_in_1279,

    output [71:0] col_out_0,
    output [71:0] col_out_1,
    output [71:0] col_out_2,
    output [71:0] col_out_3,
    output [71:0] col_out_4,
    output [71:0] col_out_5,
    output [71:0] col_out_6,
    output [71:0] col_out_7,
    output [71:0] col_out_8,
    output [71:0] col_out_9,
    output [71:0] col_out_10,
    output [71:0] col_out_11,
    output [71:0] col_out_12,
    output [71:0] col_out_13,
    output [71:0] col_out_14,
    output [71:0] col_out_15,
    output [71:0] col_out_16,
    output [71:0] col_out_17,
    output [71:0] col_out_18,
    output [71:0] col_out_19,
    output [71:0] col_out_20,
    output [71:0] col_out_21,
    output [71:0] col_out_22,
    output [71:0] col_out_23,
    output [71:0] col_out_24,
    output [71:0] col_out_25,
    output [71:0] col_out_26,
    output [71:0] col_out_27,
    output [71:0] col_out_28,
    output [71:0] col_out_29,
    output [71:0] col_out_30,
    output [71:0] col_out_31,
    output [71:0] col_out_32,
    output [71:0] col_out_33,
    output [71:0] col_out_34,
    output [71:0] col_out_35,
    output [71:0] col_out_36,
    output [71:0] col_out_37,
    output [71:0] col_out_38,
    output [71:0] col_out_39,
    output [71:0] col_out_40,
    output [71:0] col_out_41,
    output [71:0] col_out_42,
    output [71:0] col_out_43,
    output [71:0] col_out_44,
    output [71:0] col_out_45,
    output [71:0] col_out_46,
    output [71:0] col_out_47,
    output [71:0] col_out_48,
    output [71:0] col_out_49,
    output [71:0] col_out_50,
    output [71:0] col_out_51,
    output [71:0] col_out_52,
    output [71:0] col_out_53,
    output [71:0] col_out_54,
    output [71:0] col_out_55,
    output [71:0] col_out_56,
    output [71:0] col_out_57,
    output [71:0] col_out_58,
    output [71:0] col_out_59,
    output [71:0] col_out_60,
    output [71:0] col_out_61,
    output [71:0] col_out_62,
    output [71:0] col_out_63,
    output [71:0] col_out_64,
    output [71:0] col_out_65,
    output [71:0] col_out_66,
    output [71:0] col_out_67,
    output [71:0] col_out_68,
    output [71:0] col_out_69,
    output [71:0] col_out_70,
    output [71:0] col_out_71,
    output [71:0] col_out_72,
    output [71:0] col_out_73,
    output [71:0] col_out_74,
    output [71:0] col_out_75,
    output [71:0] col_out_76,
    output [71:0] col_out_77,
    output [71:0] col_out_78,
    output [71:0] col_out_79,
    output [71:0] col_out_80,
    output [71:0] col_out_81,
    output [71:0] col_out_82,
    output [71:0] col_out_83,
    output [71:0] col_out_84,
    output [71:0] col_out_85,
    output [71:0] col_out_86,
    output [71:0] col_out_87,
    output [71:0] col_out_88,
    output [71:0] col_out_89,
    output [71:0] col_out_90,
    output [71:0] col_out_91,
    output [71:0] col_out_92,
    output [71:0] col_out_93,
    output [71:0] col_out_94,
    output [71:0] col_out_95,
    output [71:0] col_out_96,
    output [71:0] col_out_97,
    output [71:0] col_out_98,
    output [71:0] col_out_99,
    output [71:0] col_out_100,
    output [71:0] col_out_101,
    output [71:0] col_out_102,
    output [71:0] col_out_103,
    output [71:0] col_out_104,
    output [71:0] col_out_105,
    output [71:0] col_out_106,
    output [71:0] col_out_107,
    output [71:0] col_out_108,
    output [71:0] col_out_109,
    output [71:0] col_out_110,
    output [71:0] col_out_111,
    output [71:0] col_out_112,
    output [71:0] col_out_113,
    output [71:0] col_out_114,
    output [71:0] col_out_115,
    output [71:0] col_out_116,
    output [71:0] col_out_117,
    output [71:0] col_out_118,
    output [71:0] col_out_119,
    output [71:0] col_out_120,
    output [71:0] col_out_121,
    output [71:0] col_out_122,
    output [71:0] col_out_123,
    output [71:0] col_out_124,
    output [71:0] col_out_125,
    output [71:0] col_out_126,
    output [71:0] col_out_127,
    output [71:0] col_out_128,
    output [71:0] col_out_129,
    output [71:0] col_out_130,
    output [71:0] col_out_131,
    output [71:0] col_out_132,
    output [71:0] col_out_133,
    output [71:0] col_out_134,
    output [71:0] col_out_135,
    output [71:0] col_out_136,
    output [71:0] col_out_137,
    output [71:0] col_out_138,
    output [71:0] col_out_139,
    output [71:0] col_out_140,
    output [71:0] col_out_141,
    output [71:0] col_out_142,
    output [71:0] col_out_143,
    output [71:0] col_out_144,
    output [71:0] col_out_145,
    output [71:0] col_out_146,
    output [71:0] col_out_147,
    output [71:0] col_out_148,
    output [71:0] col_out_149,
    output [71:0] col_out_150,
    output [71:0] col_out_151,
    output [71:0] col_out_152,
    output [71:0] col_out_153,
    output [71:0] col_out_154,
    output [71:0] col_out_155,
    output [71:0] col_out_156,
    output [71:0] col_out_157,
    output [71:0] col_out_158,
    output [71:0] col_out_159,
    output [71:0] col_out_160,
    output [71:0] col_out_161,
    output [71:0] col_out_162,
    output [71:0] col_out_163,
    output [71:0] col_out_164,
    output [71:0] col_out_165,
    output [71:0] col_out_166,
    output [71:0] col_out_167,
    output [71:0] col_out_168,
    output [71:0] col_out_169,
    output [71:0] col_out_170,
    output [71:0] col_out_171,
    output [71:0] col_out_172,
    output [71:0] col_out_173,
    output [71:0] col_out_174,
    output [71:0] col_out_175,
    output [71:0] col_out_176,
    output [71:0] col_out_177,
    output [71:0] col_out_178,
    output [71:0] col_out_179,
    output [71:0] col_out_180,
    output [71:0] col_out_181,
    output [71:0] col_out_182,
    output [71:0] col_out_183,
    output [71:0] col_out_184,
    output [71:0] col_out_185,
    output [71:0] col_out_186,
    output [71:0] col_out_187,
    output [71:0] col_out_188,
    output [71:0] col_out_189,
    output [71:0] col_out_190,
    output [71:0] col_out_191,
    output [71:0] col_out_192,
    output [71:0] col_out_193,
    output [71:0] col_out_194,
    output [71:0] col_out_195,
    output [71:0] col_out_196,
    output [71:0] col_out_197,
    output [71:0] col_out_198,
    output [71:0] col_out_199,
    output [71:0] col_out_200,
    output [71:0] col_out_201,
    output [71:0] col_out_202,
    output [71:0] col_out_203,
    output [71:0] col_out_204,
    output [71:0] col_out_205,
    output [71:0] col_out_206,
    output [71:0] col_out_207,
    output [71:0] col_out_208,
    output [71:0] col_out_209,
    output [71:0] col_out_210,
    output [71:0] col_out_211,
    output [71:0] col_out_212,
    output [71:0] col_out_213,
    output [71:0] col_out_214,
    output [71:0] col_out_215,
    output [71:0] col_out_216,
    output [71:0] col_out_217,
    output [71:0] col_out_218,
    output [71:0] col_out_219,
    output [71:0] col_out_220,
    output [71:0] col_out_221,
    output [71:0] col_out_222,
    output [71:0] col_out_223,
    output [71:0] col_out_224,
    output [71:0] col_out_225,
    output [71:0] col_out_226,
    output [71:0] col_out_227,
    output [71:0] col_out_228,
    output [71:0] col_out_229,
    output [71:0] col_out_230,
    output [71:0] col_out_231,
    output [71:0] col_out_232,
    output [71:0] col_out_233,
    output [71:0] col_out_234,
    output [71:0] col_out_235,
    output [71:0] col_out_236,
    output [71:0] col_out_237,
    output [71:0] col_out_238,
    output [71:0] col_out_239,
    output [71:0] col_out_240,
    output [71:0] col_out_241,
    output [71:0] col_out_242,
    output [71:0] col_out_243,
    output [71:0] col_out_244,
    output [71:0] col_out_245,
    output [71:0] col_out_246,
    output [71:0] col_out_247,
    output [71:0] col_out_248,
    output [71:0] col_out_249,
    output [71:0] col_out_250,
    output [71:0] col_out_251,
    output [71:0] col_out_252,
    output [71:0] col_out_253,
    output [71:0] col_out_254,
    output [71:0] col_out_255,
    output [71:0] col_out_256,
    output [71:0] col_out_257,
    output [71:0] col_out_258,
    output [71:0] col_out_259,
    output [71:0] col_out_260,
    output [71:0] col_out_261,
    output [71:0] col_out_262,
    output [71:0] col_out_263,
    output [71:0] col_out_264,
    output [71:0] col_out_265,
    output [71:0] col_out_266,
    output [71:0] col_out_267,
    output [71:0] col_out_268,
    output [71:0] col_out_269,
    output [71:0] col_out_270,
    output [71:0] col_out_271,
    output [71:0] col_out_272,
    output [71:0] col_out_273,
    output [71:0] col_out_274,
    output [71:0] col_out_275,
    output [71:0] col_out_276,
    output [71:0] col_out_277,
    output [71:0] col_out_278,
    output [71:0] col_out_279,
    output [71:0] col_out_280,
    output [71:0] col_out_281,
    output [71:0] col_out_282,
    output [71:0] col_out_283,
    output [71:0] col_out_284,
    output [71:0] col_out_285,
    output [71:0] col_out_286,
    output [71:0] col_out_287,
    output [71:0] col_out_288,
    output [71:0] col_out_289,
    output [71:0] col_out_290,
    output [71:0] col_out_291,
    output [71:0] col_out_292,
    output [71:0] col_out_293,
    output [71:0] col_out_294,
    output [71:0] col_out_295,
    output [71:0] col_out_296,
    output [71:0] col_out_297,
    output [71:0] col_out_298,
    output [71:0] col_out_299,
    output [71:0] col_out_300,
    output [71:0] col_out_301,
    output [71:0] col_out_302,
    output [71:0] col_out_303,
    output [71:0] col_out_304,
    output [71:0] col_out_305,
    output [71:0] col_out_306,
    output [71:0] col_out_307,
    output [71:0] col_out_308,
    output [71:0] col_out_309,
    output [71:0] col_out_310,
    output [71:0] col_out_311,
    output [71:0] col_out_312,
    output [71:0] col_out_313,
    output [71:0] col_out_314,
    output [71:0] col_out_315,
    output [71:0] col_out_316,
    output [71:0] col_out_317,
    output [71:0] col_out_318,
    output [71:0] col_out_319,
    output [71:0] col_out_320,
    output [71:0] col_out_321,
    output [71:0] col_out_322,
    output [71:0] col_out_323,
    output [71:0] col_out_324,
    output [71:0] col_out_325,
    output [71:0] col_out_326,
    output [71:0] col_out_327,
    output [71:0] col_out_328,
    output [71:0] col_out_329,
    output [71:0] col_out_330,
    output [71:0] col_out_331,
    output [71:0] col_out_332,
    output [71:0] col_out_333,
    output [71:0] col_out_334,
    output [71:0] col_out_335,
    output [71:0] col_out_336,
    output [71:0] col_out_337,
    output [71:0] col_out_338,
    output [71:0] col_out_339,
    output [71:0] col_out_340,
    output [71:0] col_out_341,
    output [71:0] col_out_342,
    output [71:0] col_out_343,
    output [71:0] col_out_344,
    output [71:0] col_out_345,
    output [71:0] col_out_346,
    output [71:0] col_out_347,
    output [71:0] col_out_348,
    output [71:0] col_out_349,
    output [71:0] col_out_350,
    output [71:0] col_out_351,
    output [71:0] col_out_352,
    output [71:0] col_out_353,
    output [71:0] col_out_354,
    output [71:0] col_out_355,
    output [71:0] col_out_356,
    output [71:0] col_out_357,
    output [71:0] col_out_358,
    output [71:0] col_out_359,
    output [71:0] col_out_360,
    output [71:0] col_out_361,
    output [71:0] col_out_362,
    output [71:0] col_out_363,
    output [71:0] col_out_364,
    output [71:0] col_out_365,
    output [71:0] col_out_366,
    output [71:0] col_out_367,
    output [71:0] col_out_368,
    output [71:0] col_out_369,
    output [71:0] col_out_370,
    output [71:0] col_out_371,
    output [71:0] col_out_372,
    output [71:0] col_out_373,
    output [71:0] col_out_374,
    output [71:0] col_out_375,
    output [71:0] col_out_376,
    output [71:0] col_out_377,
    output [71:0] col_out_378,
    output [71:0] col_out_379,
    output [71:0] col_out_380,
    output [71:0] col_out_381,
    output [71:0] col_out_382,
    output [71:0] col_out_383,
    output [71:0] col_out_384,
    output [71:0] col_out_385,
    output [71:0] col_out_386,
    output [71:0] col_out_387,
    output [71:0] col_out_388,
    output [71:0] col_out_389,
    output [71:0] col_out_390,
    output [71:0] col_out_391,
    output [71:0] col_out_392,
    output [71:0] col_out_393,
    output [71:0] col_out_394,
    output [71:0] col_out_395,
    output [71:0] col_out_396,
    output [71:0] col_out_397,
    output [71:0] col_out_398,
    output [71:0] col_out_399,
    output [71:0] col_out_400,
    output [71:0] col_out_401,
    output [71:0] col_out_402,
    output [71:0] col_out_403,
    output [71:0] col_out_404,
    output [71:0] col_out_405,
    output [71:0] col_out_406,
    output [71:0] col_out_407,
    output [71:0] col_out_408,
    output [71:0] col_out_409,
    output [71:0] col_out_410,
    output [71:0] col_out_411,
    output [71:0] col_out_412,
    output [71:0] col_out_413,
    output [71:0] col_out_414,
    output [71:0] col_out_415,
    output [71:0] col_out_416,
    output [71:0] col_out_417,
    output [71:0] col_out_418,
    output [71:0] col_out_419,
    output [71:0] col_out_420,
    output [71:0] col_out_421,
    output [71:0] col_out_422,
    output [71:0] col_out_423,
    output [71:0] col_out_424,
    output [71:0] col_out_425,
    output [71:0] col_out_426,
    output [71:0] col_out_427,
    output [71:0] col_out_428,
    output [71:0] col_out_429,
    output [71:0] col_out_430,
    output [71:0] col_out_431,
    output [71:0] col_out_432,
    output [71:0] col_out_433,
    output [71:0] col_out_434,
    output [71:0] col_out_435,
    output [71:0] col_out_436,
    output [71:0] col_out_437,
    output [71:0] col_out_438,
    output [71:0] col_out_439,
    output [71:0] col_out_440,
    output [71:0] col_out_441,
    output [71:0] col_out_442,
    output [71:0] col_out_443,
    output [71:0] col_out_444,
    output [71:0] col_out_445,
    output [71:0] col_out_446,
    output [71:0] col_out_447,
    output [71:0] col_out_448,
    output [71:0] col_out_449,
    output [71:0] col_out_450,
    output [71:0] col_out_451,
    output [71:0] col_out_452,
    output [71:0] col_out_453,
    output [71:0] col_out_454,
    output [71:0] col_out_455,
    output [71:0] col_out_456,
    output [71:0] col_out_457,
    output [71:0] col_out_458,
    output [71:0] col_out_459,
    output [71:0] col_out_460,
    output [71:0] col_out_461,
    output [71:0] col_out_462,
    output [71:0] col_out_463,
    output [71:0] col_out_464,
    output [71:0] col_out_465,
    output [71:0] col_out_466,
    output [71:0] col_out_467,
    output [71:0] col_out_468,
    output [71:0] col_out_469,
    output [71:0] col_out_470,
    output [71:0] col_out_471,
    output [71:0] col_out_472,
    output [71:0] col_out_473,
    output [71:0] col_out_474,
    output [71:0] col_out_475,
    output [71:0] col_out_476,
    output [71:0] col_out_477,
    output [71:0] col_out_478,
    output [71:0] col_out_479,
    output [71:0] col_out_480,
    output [71:0] col_out_481,
    output [71:0] col_out_482,
    output [71:0] col_out_483,
    output [71:0] col_out_484,
    output [71:0] col_out_485,
    output [71:0] col_out_486,
    output [71:0] col_out_487,
    output [71:0] col_out_488,
    output [71:0] col_out_489,
    output [71:0] col_out_490,
    output [71:0] col_out_491,
    output [71:0] col_out_492,
    output [71:0] col_out_493,
    output [71:0] col_out_494,
    output [71:0] col_out_495,
    output [71:0] col_out_496,
    output [71:0] col_out_497,
    output [71:0] col_out_498,
    output [71:0] col_out_499,
    output [71:0] col_out_500,
    output [71:0] col_out_501,
    output [71:0] col_out_502,
    output [71:0] col_out_503,
    output [71:0] col_out_504,
    output [71:0] col_out_505,
    output [71:0] col_out_506,
    output [71:0] col_out_507,
    output [71:0] col_out_508,
    output [71:0] col_out_509,
    output [71:0] col_out_510,
    output [71:0] col_out_511,
    output [71:0] col_out_512,
    output [71:0] col_out_513,
    output [71:0] col_out_514,
    output [71:0] col_out_515,
    output [71:0] col_out_516,
    output [71:0] col_out_517,
    output [71:0] col_out_518,
    output [71:0] col_out_519,
    output [71:0] col_out_520,
    output [71:0] col_out_521,
    output [71:0] col_out_522,
    output [71:0] col_out_523,
    output [71:0] col_out_524,
    output [71:0] col_out_525,
    output [71:0] col_out_526,
    output [71:0] col_out_527,
    output [71:0] col_out_528,
    output [71:0] col_out_529,
    output [71:0] col_out_530,
    output [71:0] col_out_531,
    output [71:0] col_out_532,
    output [71:0] col_out_533,
    output [71:0] col_out_534,
    output [71:0] col_out_535,
    output [71:0] col_out_536,
    output [71:0] col_out_537,
    output [71:0] col_out_538,
    output [71:0] col_out_539,
    output [71:0] col_out_540,
    output [71:0] col_out_541,
    output [71:0] col_out_542,
    output [71:0] col_out_543,
    output [71:0] col_out_544,
    output [71:0] col_out_545,
    output [71:0] col_out_546,
    output [71:0] col_out_547,
    output [71:0] col_out_548,
    output [71:0] col_out_549,
    output [71:0] col_out_550,
    output [71:0] col_out_551,
    output [71:0] col_out_552,
    output [71:0] col_out_553,
    output [71:0] col_out_554,
    output [71:0] col_out_555,
    output [71:0] col_out_556,
    output [71:0] col_out_557,
    output [71:0] col_out_558,
    output [71:0] col_out_559,
    output [71:0] col_out_560,
    output [71:0] col_out_561,
    output [71:0] col_out_562,
    output [71:0] col_out_563,
    output [71:0] col_out_564,
    output [71:0] col_out_565,
    output [71:0] col_out_566,
    output [71:0] col_out_567,
    output [71:0] col_out_568,
    output [71:0] col_out_569,
    output [71:0] col_out_570,
    output [71:0] col_out_571,
    output [71:0] col_out_572,
    output [71:0] col_out_573,
    output [71:0] col_out_574,
    output [71:0] col_out_575,
    output [71:0] col_out_576,
    output [71:0] col_out_577,
    output [71:0] col_out_578,
    output [71:0] col_out_579,
    output [71:0] col_out_580,
    output [71:0] col_out_581,
    output [71:0] col_out_582,
    output [71:0] col_out_583,
    output [71:0] col_out_584,
    output [71:0] col_out_585,
    output [71:0] col_out_586,
    output [71:0] col_out_587,
    output [71:0] col_out_588,
    output [71:0] col_out_589,
    output [71:0] col_out_590,
    output [71:0] col_out_591,
    output [71:0] col_out_592,
    output [71:0] col_out_593,
    output [71:0] col_out_594,
    output [71:0] col_out_595,
    output [71:0] col_out_596,
    output [71:0] col_out_597,
    output [71:0] col_out_598,
    output [71:0] col_out_599,
    output [71:0] col_out_600,
    output [71:0] col_out_601,
    output [71:0] col_out_602,
    output [71:0] col_out_603,
    output [71:0] col_out_604,
    output [71:0] col_out_605,
    output [71:0] col_out_606,
    output [71:0] col_out_607,
    output [71:0] col_out_608,
    output [71:0] col_out_609,
    output [71:0] col_out_610,
    output [71:0] col_out_611,
    output [71:0] col_out_612,
    output [71:0] col_out_613,
    output [71:0] col_out_614,
    output [71:0] col_out_615,
    output [71:0] col_out_616,
    output [71:0] col_out_617,
    output [71:0] col_out_618,
    output [71:0] col_out_619,
    output [71:0] col_out_620,
    output [71:0] col_out_621,
    output [71:0] col_out_622,
    output [71:0] col_out_623,
    output [71:0] col_out_624,
    output [71:0] col_out_625,
    output [71:0] col_out_626,
    output [71:0] col_out_627,
    output [71:0] col_out_628,
    output [71:0] col_out_629,
    output [71:0] col_out_630,
    output [71:0] col_out_631,
    output [71:0] col_out_632,
    output [71:0] col_out_633,
    output [71:0] col_out_634,
    output [71:0] col_out_635,
    output [71:0] col_out_636,
    output [71:0] col_out_637,
    output [71:0] col_out_638,
    output [71:0] col_out_639,
    output [71:0] col_out_640,
    output [71:0] col_out_641,
    output [71:0] col_out_642,
    output [71:0] col_out_643,
    output [71:0] col_out_644,
    output [71:0] col_out_645,
    output [71:0] col_out_646,
    output [71:0] col_out_647,
    output [71:0] col_out_648,
    output [71:0] col_out_649,
    output [71:0] col_out_650,
    output [71:0] col_out_651,
    output [71:0] col_out_652,
    output [71:0] col_out_653,
    output [71:0] col_out_654,
    output [71:0] col_out_655,
    output [71:0] col_out_656,
    output [71:0] col_out_657,
    output [71:0] col_out_658,
    output [71:0] col_out_659,
    output [71:0] col_out_660,
    output [71:0] col_out_661,
    output [71:0] col_out_662,
    output [71:0] col_out_663,
    output [71:0] col_out_664,
    output [71:0] col_out_665,
    output [71:0] col_out_666,
    output [71:0] col_out_667,
    output [71:0] col_out_668,
    output [71:0] col_out_669,
    output [71:0] col_out_670,
    output [71:0] col_out_671,
    output [71:0] col_out_672,
    output [71:0] col_out_673,
    output [71:0] col_out_674,
    output [71:0] col_out_675,
    output [71:0] col_out_676,
    output [71:0] col_out_677,
    output [71:0] col_out_678,
    output [71:0] col_out_679,
    output [71:0] col_out_680,
    output [71:0] col_out_681,
    output [71:0] col_out_682,
    output [71:0] col_out_683,
    output [71:0] col_out_684,
    output [71:0] col_out_685,
    output [71:0] col_out_686,
    output [71:0] col_out_687,
    output [71:0] col_out_688,
    output [71:0] col_out_689,
    output [71:0] col_out_690,
    output [71:0] col_out_691,
    output [71:0] col_out_692,
    output [71:0] col_out_693,
    output [71:0] col_out_694,
    output [71:0] col_out_695,
    output [71:0] col_out_696,
    output [71:0] col_out_697,
    output [71:0] col_out_698,
    output [71:0] col_out_699,
    output [71:0] col_out_700,
    output [71:0] col_out_701,
    output [71:0] col_out_702,
    output [71:0] col_out_703,
    output [71:0] col_out_704,
    output [71:0] col_out_705,
    output [71:0] col_out_706,
    output [71:0] col_out_707,
    output [71:0] col_out_708,
    output [71:0] col_out_709,
    output [71:0] col_out_710,
    output [71:0] col_out_711,
    output [71:0] col_out_712,
    output [71:0] col_out_713,
    output [71:0] col_out_714,
    output [71:0] col_out_715,
    output [71:0] col_out_716,
    output [71:0] col_out_717,
    output [71:0] col_out_718,
    output [71:0] col_out_719,
    output [71:0] col_out_720,
    output [71:0] col_out_721,
    output [71:0] col_out_722,
    output [71:0] col_out_723,
    output [71:0] col_out_724,
    output [71:0] col_out_725,
    output [71:0] col_out_726,
    output [71:0] col_out_727,
    output [71:0] col_out_728,
    output [71:0] col_out_729,
    output [71:0] col_out_730,
    output [71:0] col_out_731,
    output [71:0] col_out_732,
    output [71:0] col_out_733,
    output [71:0] col_out_734,
    output [71:0] col_out_735,
    output [71:0] col_out_736,
    output [71:0] col_out_737,
    output [71:0] col_out_738,
    output [71:0] col_out_739,
    output [71:0] col_out_740,
    output [71:0] col_out_741,
    output [71:0] col_out_742,
    output [71:0] col_out_743,
    output [71:0] col_out_744,
    output [71:0] col_out_745,
    output [71:0] col_out_746,
    output [71:0] col_out_747,
    output [71:0] col_out_748,
    output [71:0] col_out_749,
    output [71:0] col_out_750,
    output [71:0] col_out_751,
    output [71:0] col_out_752,
    output [71:0] col_out_753,
    output [71:0] col_out_754,
    output [71:0] col_out_755,
    output [71:0] col_out_756,
    output [71:0] col_out_757,
    output [71:0] col_out_758,
    output [71:0] col_out_759,
    output [71:0] col_out_760,
    output [71:0] col_out_761,
    output [71:0] col_out_762,
    output [71:0] col_out_763,
    output [71:0] col_out_764,
    output [71:0] col_out_765,
    output [71:0] col_out_766,
    output [71:0] col_out_767,
    output [71:0] col_out_768,
    output [71:0] col_out_769,
    output [71:0] col_out_770,
    output [71:0] col_out_771,
    output [71:0] col_out_772,
    output [71:0] col_out_773,
    output [71:0] col_out_774,
    output [71:0] col_out_775,
    output [71:0] col_out_776,
    output [71:0] col_out_777,
    output [71:0] col_out_778,
    output [71:0] col_out_779,
    output [71:0] col_out_780,
    output [71:0] col_out_781,
    output [71:0] col_out_782,
    output [71:0] col_out_783,
    output [71:0] col_out_784,
    output [71:0] col_out_785,
    output [71:0] col_out_786,
    output [71:0] col_out_787,
    output [71:0] col_out_788,
    output [71:0] col_out_789,
    output [71:0] col_out_790,
    output [71:0] col_out_791,
    output [71:0] col_out_792,
    output [71:0] col_out_793,
    output [71:0] col_out_794,
    output [71:0] col_out_795,
    output [71:0] col_out_796,
    output [71:0] col_out_797,
    output [71:0] col_out_798,
    output [71:0] col_out_799,
    output [71:0] col_out_800,
    output [71:0] col_out_801,
    output [71:0] col_out_802,
    output [71:0] col_out_803,
    output [71:0] col_out_804,
    output [71:0] col_out_805,
    output [71:0] col_out_806,
    output [71:0] col_out_807,
    output [71:0] col_out_808,
    output [71:0] col_out_809,
    output [71:0] col_out_810,
    output [71:0] col_out_811,
    output [71:0] col_out_812,
    output [71:0] col_out_813,
    output [71:0] col_out_814,
    output [71:0] col_out_815,
    output [71:0] col_out_816,
    output [71:0] col_out_817,
    output [71:0] col_out_818,
    output [71:0] col_out_819,
    output [71:0] col_out_820,
    output [71:0] col_out_821,
    output [71:0] col_out_822,
    output [71:0] col_out_823,
    output [71:0] col_out_824,
    output [71:0] col_out_825,
    output [71:0] col_out_826,
    output [71:0] col_out_827,
    output [71:0] col_out_828,
    output [71:0] col_out_829,
    output [71:0] col_out_830,
    output [71:0] col_out_831,
    output [71:0] col_out_832,
    output [71:0] col_out_833,
    output [71:0] col_out_834,
    output [71:0] col_out_835,
    output [71:0] col_out_836,
    output [71:0] col_out_837,
    output [71:0] col_out_838,
    output [71:0] col_out_839,
    output [71:0] col_out_840,
    output [71:0] col_out_841,
    output [71:0] col_out_842,
    output [71:0] col_out_843,
    output [71:0] col_out_844,
    output [71:0] col_out_845,
    output [71:0] col_out_846,
    output [71:0] col_out_847,
    output [71:0] col_out_848,
    output [71:0] col_out_849,
    output [71:0] col_out_850,
    output [71:0] col_out_851,
    output [71:0] col_out_852,
    output [71:0] col_out_853,
    output [71:0] col_out_854,
    output [71:0] col_out_855,
    output [71:0] col_out_856,
    output [71:0] col_out_857,
    output [71:0] col_out_858,
    output [71:0] col_out_859,
    output [71:0] col_out_860,
    output [71:0] col_out_861,
    output [71:0] col_out_862,
    output [71:0] col_out_863,
    output [71:0] col_out_864,
    output [71:0] col_out_865,
    output [71:0] col_out_866,
    output [71:0] col_out_867,
    output [71:0] col_out_868,
    output [71:0] col_out_869,
    output [71:0] col_out_870,
    output [71:0] col_out_871,
    output [71:0] col_out_872,
    output [71:0] col_out_873,
    output [71:0] col_out_874,
    output [71:0] col_out_875,
    output [71:0] col_out_876,
    output [71:0] col_out_877,
    output [71:0] col_out_878,
    output [71:0] col_out_879,
    output [71:0] col_out_880,
    output [71:0] col_out_881,
    output [71:0] col_out_882,
    output [71:0] col_out_883,
    output [71:0] col_out_884,
    output [71:0] col_out_885,
    output [71:0] col_out_886,
    output [71:0] col_out_887,
    output [71:0] col_out_888,
    output [71:0] col_out_889,
    output [71:0] col_out_890,
    output [71:0] col_out_891,
    output [71:0] col_out_892,
    output [71:0] col_out_893,
    output [71:0] col_out_894,
    output [71:0] col_out_895,
    output [71:0] col_out_896,
    output [71:0] col_out_897,
    output [71:0] col_out_898,
    output [71:0] col_out_899,
    output [71:0] col_out_900,
    output [71:0] col_out_901,
    output [71:0] col_out_902,
    output [71:0] col_out_903,
    output [71:0] col_out_904,
    output [71:0] col_out_905,
    output [71:0] col_out_906,
    output [71:0] col_out_907,
    output [71:0] col_out_908,
    output [71:0] col_out_909,
    output [71:0] col_out_910,
    output [71:0] col_out_911,
    output [71:0] col_out_912,
    output [71:0] col_out_913,
    output [71:0] col_out_914,
    output [71:0] col_out_915,
    output [71:0] col_out_916,
    output [71:0] col_out_917,
    output [71:0] col_out_918,
    output [71:0] col_out_919,
    output [71:0] col_out_920,
    output [71:0] col_out_921,
    output [71:0] col_out_922,
    output [71:0] col_out_923,
    output [71:0] col_out_924,
    output [71:0] col_out_925,
    output [71:0] col_out_926,
    output [71:0] col_out_927,
    output [71:0] col_out_928,
    output [71:0] col_out_929,
    output [71:0] col_out_930,
    output [71:0] col_out_931,
    output [71:0] col_out_932,
    output [71:0] col_out_933,
    output [71:0] col_out_934,
    output [71:0] col_out_935,
    output [71:0] col_out_936,
    output [71:0] col_out_937,
    output [71:0] col_out_938,
    output [71:0] col_out_939,
    output [71:0] col_out_940,
    output [71:0] col_out_941,
    output [71:0] col_out_942,
    output [71:0] col_out_943,
    output [71:0] col_out_944,
    output [71:0] col_out_945,
    output [71:0] col_out_946,
    output [71:0] col_out_947,
    output [71:0] col_out_948,
    output [71:0] col_out_949,
    output [71:0] col_out_950,
    output [71:0] col_out_951,
    output [71:0] col_out_952,
    output [71:0] col_out_953,
    output [71:0] col_out_954,
    output [71:0] col_out_955,
    output [71:0] col_out_956,
    output [71:0] col_out_957,
    output [71:0] col_out_958,
    output [71:0] col_out_959,
    output [71:0] col_out_960,
    output [71:0] col_out_961,
    output [71:0] col_out_962,
    output [71:0] col_out_963,
    output [71:0] col_out_964,
    output [71:0] col_out_965,
    output [71:0] col_out_966,
    output [71:0] col_out_967,
    output [71:0] col_out_968,
    output [71:0] col_out_969,
    output [71:0] col_out_970,
    output [71:0] col_out_971,
    output [71:0] col_out_972,
    output [71:0] col_out_973,
    output [71:0] col_out_974,
    output [71:0] col_out_975,
    output [71:0] col_out_976,
    output [71:0] col_out_977,
    output [71:0] col_out_978,
    output [71:0] col_out_979,
    output [71:0] col_out_980,
    output [71:0] col_out_981,
    output [71:0] col_out_982,
    output [71:0] col_out_983,
    output [71:0] col_out_984,
    output [71:0] col_out_985,
    output [71:0] col_out_986,
    output [71:0] col_out_987,
    output [71:0] col_out_988,
    output [71:0] col_out_989,
    output [71:0] col_out_990,
    output [71:0] col_out_991,
    output [71:0] col_out_992,
    output [71:0] col_out_993,
    output [71:0] col_out_994,
    output [71:0] col_out_995,
    output [71:0] col_out_996,
    output [71:0] col_out_997,
    output [71:0] col_out_998,
    output [71:0] col_out_999,
    output [71:0] col_out_1000,
    output [71:0] col_out_1001,
    output [71:0] col_out_1002,
    output [71:0] col_out_1003,
    output [71:0] col_out_1004,
    output [71:0] col_out_1005,
    output [71:0] col_out_1006,
    output [71:0] col_out_1007,
    output [71:0] col_out_1008,
    output [71:0] col_out_1009,
    output [71:0] col_out_1010,
    output [71:0] col_out_1011,
    output [71:0] col_out_1012,
    output [71:0] col_out_1013,
    output [71:0] col_out_1014,
    output [71:0] col_out_1015,
    output [71:0] col_out_1016,
    output [71:0] col_out_1017,
    output [71:0] col_out_1018,
    output [71:0] col_out_1019,
    output [71:0] col_out_1020,
    output [71:0] col_out_1021,
    output [71:0] col_out_1022,
    output [71:0] col_out_1023,
    output [71:0] col_out_1024,
    output [71:0] col_out_1025,
    output [71:0] col_out_1026,
    output [71:0] col_out_1027,
    output [71:0] col_out_1028,
    output [71:0] col_out_1029,
    output [71:0] col_out_1030,
    output [71:0] col_out_1031,
    output [71:0] col_out_1032,
    output [71:0] col_out_1033,
    output [71:0] col_out_1034,
    output [71:0] col_out_1035,
    output [71:0] col_out_1036,
    output [71:0] col_out_1037,
    output [71:0] col_out_1038,
    output [71:0] col_out_1039,
    output [71:0] col_out_1040,
    output [71:0] col_out_1041,
    output [71:0] col_out_1042,
    output [71:0] col_out_1043,
    output [71:0] col_out_1044,
    output [71:0] col_out_1045,
    output [71:0] col_out_1046,
    output [71:0] col_out_1047,
    output [71:0] col_out_1048,
    output [71:0] col_out_1049,
    output [71:0] col_out_1050,
    output [71:0] col_out_1051,
    output [71:0] col_out_1052,
    output [71:0] col_out_1053,
    output [71:0] col_out_1054,
    output [71:0] col_out_1055,
    output [71:0] col_out_1056,
    output [71:0] col_out_1057,
    output [71:0] col_out_1058,
    output [71:0] col_out_1059,
    output [71:0] col_out_1060,
    output [71:0] col_out_1061,
    output [71:0] col_out_1062,
    output [71:0] col_out_1063,
    output [71:0] col_out_1064,
    output [71:0] col_out_1065,
    output [71:0] col_out_1066,
    output [71:0] col_out_1067,
    output [71:0] col_out_1068,
    output [71:0] col_out_1069,
    output [71:0] col_out_1070,
    output [71:0] col_out_1071,
    output [71:0] col_out_1072,
    output [71:0] col_out_1073,
    output [71:0] col_out_1074,
    output [71:0] col_out_1075,
    output [71:0] col_out_1076,
    output [71:0] col_out_1077,
    output [71:0] col_out_1078,
    output [71:0] col_out_1079,
    output [71:0] col_out_1080,
    output [71:0] col_out_1081,
    output [71:0] col_out_1082,
    output [71:0] col_out_1083,
    output [71:0] col_out_1084,
    output [71:0] col_out_1085,
    output [71:0] col_out_1086,
    output [71:0] col_out_1087,
    output [71:0] col_out_1088,
    output [71:0] col_out_1089,
    output [71:0] col_out_1090,
    output [71:0] col_out_1091,
    output [71:0] col_out_1092,
    output [71:0] col_out_1093,
    output [71:0] col_out_1094,
    output [71:0] col_out_1095,
    output [71:0] col_out_1096,
    output [71:0] col_out_1097,
    output [71:0] col_out_1098,
    output [71:0] col_out_1099,
    output [71:0] col_out_1100,
    output [71:0] col_out_1101,
    output [71:0] col_out_1102,
    output [71:0] col_out_1103,
    output [71:0] col_out_1104,
    output [71:0] col_out_1105,
    output [71:0] col_out_1106,
    output [71:0] col_out_1107,
    output [71:0] col_out_1108,
    output [71:0] col_out_1109,
    output [71:0] col_out_1110,
    output [71:0] col_out_1111,
    output [71:0] col_out_1112,
    output [71:0] col_out_1113,
    output [71:0] col_out_1114,
    output [71:0] col_out_1115,
    output [71:0] col_out_1116,
    output [71:0] col_out_1117,
    output [71:0] col_out_1118,
    output [71:0] col_out_1119,
    output [71:0] col_out_1120,
    output [71:0] col_out_1121,
    output [71:0] col_out_1122,
    output [71:0] col_out_1123,
    output [71:0] col_out_1124,
    output [71:0] col_out_1125,
    output [71:0] col_out_1126,
    output [71:0] col_out_1127,
    output [71:0] col_out_1128,
    output [71:0] col_out_1129,
    output [71:0] col_out_1130,
    output [71:0] col_out_1131,
    output [71:0] col_out_1132,
    output [71:0] col_out_1133,
    output [71:0] col_out_1134,
    output [71:0] col_out_1135,
    output [71:0] col_out_1136,
    output [71:0] col_out_1137,
    output [71:0] col_out_1138,
    output [71:0] col_out_1139,
    output [71:0] col_out_1140,
    output [71:0] col_out_1141,
    output [71:0] col_out_1142,
    output [71:0] col_out_1143,
    output [71:0] col_out_1144,
    output [71:0] col_out_1145,
    output [71:0] col_out_1146,
    output [71:0] col_out_1147,
    output [71:0] col_out_1148,
    output [71:0] col_out_1149,
    output [71:0] col_out_1150,
    output [71:0] col_out_1151,
    output [71:0] col_out_1152,
    output [71:0] col_out_1153,
    output [71:0] col_out_1154,
    output [71:0] col_out_1155,
    output [71:0] col_out_1156,
    output [71:0] col_out_1157,
    output [71:0] col_out_1158,
    output [71:0] col_out_1159,
    output [71:0] col_out_1160,
    output [71:0] col_out_1161,
    output [71:0] col_out_1162,
    output [71:0] col_out_1163,
    output [71:0] col_out_1164,
    output [71:0] col_out_1165,
    output [71:0] col_out_1166,
    output [71:0] col_out_1167,
    output [71:0] col_out_1168,
    output [71:0] col_out_1169,
    output [71:0] col_out_1170,
    output [71:0] col_out_1171,
    output [71:0] col_out_1172,
    output [71:0] col_out_1173,
    output [71:0] col_out_1174,
    output [71:0] col_out_1175,
    output [71:0] col_out_1176,
    output [71:0] col_out_1177,
    output [71:0] col_out_1178,
    output [71:0] col_out_1179,
    output [71:0] col_out_1180,
    output [71:0] col_out_1181,
    output [71:0] col_out_1182,
    output [71:0] col_out_1183,
    output [71:0] col_out_1184,
    output [71:0] col_out_1185,
    output [71:0] col_out_1186,
    output [71:0] col_out_1187,
    output [71:0] col_out_1188,
    output [71:0] col_out_1189,
    output [71:0] col_out_1190,
    output [71:0] col_out_1191,
    output [71:0] col_out_1192,
    output [71:0] col_out_1193,
    output [71:0] col_out_1194,
    output [71:0] col_out_1195,
    output [71:0] col_out_1196,
    output [71:0] col_out_1197,
    output [71:0] col_out_1198,
    output [71:0] col_out_1199,
    output [71:0] col_out_1200,
    output [71:0] col_out_1201,
    output [71:0] col_out_1202,
    output [71:0] col_out_1203,
    output [71:0] col_out_1204,
    output [71:0] col_out_1205,
    output [71:0] col_out_1206,
    output [71:0] col_out_1207,
    output [71:0] col_out_1208,
    output [71:0] col_out_1209,
    output [71:0] col_out_1210,
    output [71:0] col_out_1211,
    output [71:0] col_out_1212,
    output [71:0] col_out_1213,
    output [71:0] col_out_1214,
    output [71:0] col_out_1215,
    output [71:0] col_out_1216,
    output [71:0] col_out_1217,
    output [71:0] col_out_1218,
    output [71:0] col_out_1219,
    output [71:0] col_out_1220,
    output [71:0] col_out_1221,
    output [71:0] col_out_1222,
    output [71:0] col_out_1223,
    output [71:0] col_out_1224,
    output [71:0] col_out_1225,
    output [71:0] col_out_1226,
    output [71:0] col_out_1227,
    output [71:0] col_out_1228,
    output [71:0] col_out_1229,
    output [71:0] col_out_1230,
    output [71:0] col_out_1231,
    output [71:0] col_out_1232,
    output [71:0] col_out_1233,
    output [71:0] col_out_1234,
    output [71:0] col_out_1235,
    output [71:0] col_out_1236,
    output [71:0] col_out_1237,
    output [71:0] col_out_1238,
    output [71:0] col_out_1239,
    output [71:0] col_out_1240,
    output [71:0] col_out_1241,
    output [71:0] col_out_1242,
    output [71:0] col_out_1243,
    output [71:0] col_out_1244,
    output [71:0] col_out_1245,
    output [71:0] col_out_1246,
    output [71:0] col_out_1247,
    output [71:0] col_out_1248,
    output [71:0] col_out_1249,
    output [71:0] col_out_1250,
    output [71:0] col_out_1251,
    output [71:0] col_out_1252,
    output [71:0] col_out_1253,
    output [71:0] col_out_1254,
    output [71:0] col_out_1255,
    output [71:0] col_out_1256,
    output [71:0] col_out_1257,
    output [71:0] col_out_1258,
    output [71:0] col_out_1259,
    output [71:0] col_out_1260,
    output [71:0] col_out_1261,
    output [71:0] col_out_1262,
    output [71:0] col_out_1263,
    output [71:0] col_out_1264,
    output [71:0] col_out_1265,
    output [71:0] col_out_1266,
    output [71:0] col_out_1267,
    output [71:0] col_out_1268,
    output [71:0] col_out_1269,
    output [71:0] col_out_1270,
    output [71:0] col_out_1271,
    output [71:0] col_out_1272,
    output [71:0] col_out_1273,
    output [71:0] col_out_1274,
    output [71:0] col_out_1275,
    output [71:0] col_out_1276,
    output [71:0] col_out_1277,
    output [71:0] col_out_1278,
    output [71:0] col_out_1279,
    output [71:0] col_out_1280,
    output [71:0] col_out_1281,
    output [71:0] col_out_1282
);



//--compressor_array input and output----------------------

wire [242:0] u_ca_in_0;
wire [242:0] u_ca_in_1;
wire [242:0] u_ca_in_2;
wire [242:0] u_ca_in_3;
wire [242:0] u_ca_in_4;
wire [242:0] u_ca_in_5;
wire [242:0] u_ca_in_6;
wire [242:0] u_ca_in_7;
wire [242:0] u_ca_in_8;
wire [242:0] u_ca_in_9;
wire [242:0] u_ca_in_10;
wire [242:0] u_ca_in_11;
wire [242:0] u_ca_in_12;
wire [242:0] u_ca_in_13;
wire [242:0] u_ca_in_14;
wire [242:0] u_ca_in_15;
wire [242:0] u_ca_in_16;
wire [242:0] u_ca_in_17;
wire [242:0] u_ca_in_18;
wire [242:0] u_ca_in_19;
wire [242:0] u_ca_in_20;
wire [242:0] u_ca_in_21;
wire [242:0] u_ca_in_22;
wire [242:0] u_ca_in_23;
wire [242:0] u_ca_in_24;
wire [242:0] u_ca_in_25;
wire [242:0] u_ca_in_26;
wire [242:0] u_ca_in_27;
wire [242:0] u_ca_in_28;
wire [242:0] u_ca_in_29;
wire [242:0] u_ca_in_30;
wire [242:0] u_ca_in_31;
wire [242:0] u_ca_in_32;
wire [242:0] u_ca_in_33;
wire [242:0] u_ca_in_34;
wire [242:0] u_ca_in_35;
wire [242:0] u_ca_in_36;
wire [242:0] u_ca_in_37;
wire [242:0] u_ca_in_38;
wire [242:0] u_ca_in_39;
wire [242:0] u_ca_in_40;
wire [242:0] u_ca_in_41;
wire [242:0] u_ca_in_42;
wire [242:0] u_ca_in_43;
wire [242:0] u_ca_in_44;
wire [242:0] u_ca_in_45;
wire [242:0] u_ca_in_46;
wire [242:0] u_ca_in_47;
wire [242:0] u_ca_in_48;
wire [242:0] u_ca_in_49;
wire [242:0] u_ca_in_50;
wire [242:0] u_ca_in_51;
wire [242:0] u_ca_in_52;
wire [242:0] u_ca_in_53;
wire [242:0] u_ca_in_54;
wire [242:0] u_ca_in_55;
wire [242:0] u_ca_in_56;
wire [242:0] u_ca_in_57;
wire [242:0] u_ca_in_58;
wire [242:0] u_ca_in_59;
wire [242:0] u_ca_in_60;
wire [242:0] u_ca_in_61;
wire [242:0] u_ca_in_62;
wire [242:0] u_ca_in_63;
wire [242:0] u_ca_in_64;
wire [242:0] u_ca_in_65;
wire [242:0] u_ca_in_66;
wire [242:0] u_ca_in_67;
wire [242:0] u_ca_in_68;
wire [242:0] u_ca_in_69;
wire [242:0] u_ca_in_70;
wire [242:0] u_ca_in_71;
wire [242:0] u_ca_in_72;
wire [242:0] u_ca_in_73;
wire [242:0] u_ca_in_74;
wire [242:0] u_ca_in_75;
wire [242:0] u_ca_in_76;
wire [242:0] u_ca_in_77;
wire [242:0] u_ca_in_78;
wire [242:0] u_ca_in_79;
wire [242:0] u_ca_in_80;
wire [242:0] u_ca_in_81;
wire [242:0] u_ca_in_82;
wire [242:0] u_ca_in_83;
wire [242:0] u_ca_in_84;
wire [242:0] u_ca_in_85;
wire [242:0] u_ca_in_86;
wire [242:0] u_ca_in_87;
wire [242:0] u_ca_in_88;
wire [242:0] u_ca_in_89;
wire [242:0] u_ca_in_90;
wire [242:0] u_ca_in_91;
wire [242:0] u_ca_in_92;
wire [242:0] u_ca_in_93;
wire [242:0] u_ca_in_94;
wire [242:0] u_ca_in_95;
wire [242:0] u_ca_in_96;
wire [242:0] u_ca_in_97;
wire [242:0] u_ca_in_98;
wire [242:0] u_ca_in_99;
wire [242:0] u_ca_in_100;
wire [242:0] u_ca_in_101;
wire [242:0] u_ca_in_102;
wire [242:0] u_ca_in_103;
wire [242:0] u_ca_in_104;
wire [242:0] u_ca_in_105;
wire [242:0] u_ca_in_106;
wire [242:0] u_ca_in_107;
wire [242:0] u_ca_in_108;
wire [242:0] u_ca_in_109;
wire [242:0] u_ca_in_110;
wire [242:0] u_ca_in_111;
wire [242:0] u_ca_in_112;
wire [242:0] u_ca_in_113;
wire [242:0] u_ca_in_114;
wire [242:0] u_ca_in_115;
wire [242:0] u_ca_in_116;
wire [242:0] u_ca_in_117;
wire [242:0] u_ca_in_118;
wire [242:0] u_ca_in_119;
wire [242:0] u_ca_in_120;
wire [242:0] u_ca_in_121;
wire [242:0] u_ca_in_122;
wire [242:0] u_ca_in_123;
wire [242:0] u_ca_in_124;
wire [242:0] u_ca_in_125;
wire [242:0] u_ca_in_126;
wire [242:0] u_ca_in_127;
wire [242:0] u_ca_in_128;
wire [242:0] u_ca_in_129;
wire [242:0] u_ca_in_130;
wire [242:0] u_ca_in_131;
wire [242:0] u_ca_in_132;
wire [242:0] u_ca_in_133;
wire [242:0] u_ca_in_134;
wire [242:0] u_ca_in_135;
wire [242:0] u_ca_in_136;
wire [242:0] u_ca_in_137;
wire [242:0] u_ca_in_138;
wire [242:0] u_ca_in_139;
wire [242:0] u_ca_in_140;
wire [242:0] u_ca_in_141;
wire [242:0] u_ca_in_142;
wire [242:0] u_ca_in_143;
wire [242:0] u_ca_in_144;
wire [242:0] u_ca_in_145;
wire [242:0] u_ca_in_146;
wire [242:0] u_ca_in_147;
wire [242:0] u_ca_in_148;
wire [242:0] u_ca_in_149;
wire [242:0] u_ca_in_150;
wire [242:0] u_ca_in_151;
wire [242:0] u_ca_in_152;
wire [242:0] u_ca_in_153;
wire [242:0] u_ca_in_154;
wire [242:0] u_ca_in_155;
wire [242:0] u_ca_in_156;
wire [242:0] u_ca_in_157;
wire [242:0] u_ca_in_158;
wire [242:0] u_ca_in_159;
wire [242:0] u_ca_in_160;
wire [242:0] u_ca_in_161;
wire [242:0] u_ca_in_162;
wire [242:0] u_ca_in_163;
wire [242:0] u_ca_in_164;
wire [242:0] u_ca_in_165;
wire [242:0] u_ca_in_166;
wire [242:0] u_ca_in_167;
wire [242:0] u_ca_in_168;
wire [242:0] u_ca_in_169;
wire [242:0] u_ca_in_170;
wire [242:0] u_ca_in_171;
wire [242:0] u_ca_in_172;
wire [242:0] u_ca_in_173;
wire [242:0] u_ca_in_174;
wire [242:0] u_ca_in_175;
wire [242:0] u_ca_in_176;
wire [242:0] u_ca_in_177;
wire [242:0] u_ca_in_178;
wire [242:0] u_ca_in_179;
wire [242:0] u_ca_in_180;
wire [242:0] u_ca_in_181;
wire [242:0] u_ca_in_182;
wire [242:0] u_ca_in_183;
wire [242:0] u_ca_in_184;
wire [242:0] u_ca_in_185;
wire [242:0] u_ca_in_186;
wire [242:0] u_ca_in_187;
wire [242:0] u_ca_in_188;
wire [242:0] u_ca_in_189;
wire [242:0] u_ca_in_190;
wire [242:0] u_ca_in_191;
wire [242:0] u_ca_in_192;
wire [242:0] u_ca_in_193;
wire [242:0] u_ca_in_194;
wire [242:0] u_ca_in_195;
wire [242:0] u_ca_in_196;
wire [242:0] u_ca_in_197;
wire [242:0] u_ca_in_198;
wire [242:0] u_ca_in_199;
wire [242:0] u_ca_in_200;
wire [242:0] u_ca_in_201;
wire [242:0] u_ca_in_202;
wire [242:0] u_ca_in_203;
wire [242:0] u_ca_in_204;
wire [242:0] u_ca_in_205;
wire [242:0] u_ca_in_206;
wire [242:0] u_ca_in_207;
wire [242:0] u_ca_in_208;
wire [242:0] u_ca_in_209;
wire [242:0] u_ca_in_210;
wire [242:0] u_ca_in_211;
wire [242:0] u_ca_in_212;
wire [242:0] u_ca_in_213;
wire [242:0] u_ca_in_214;
wire [242:0] u_ca_in_215;
wire [242:0] u_ca_in_216;
wire [242:0] u_ca_in_217;
wire [242:0] u_ca_in_218;
wire [242:0] u_ca_in_219;
wire [242:0] u_ca_in_220;
wire [242:0] u_ca_in_221;
wire [242:0] u_ca_in_222;
wire [242:0] u_ca_in_223;
wire [242:0] u_ca_in_224;
wire [242:0] u_ca_in_225;
wire [242:0] u_ca_in_226;
wire [242:0] u_ca_in_227;
wire [242:0] u_ca_in_228;
wire [242:0] u_ca_in_229;
wire [242:0] u_ca_in_230;
wire [242:0] u_ca_in_231;
wire [242:0] u_ca_in_232;
wire [242:0] u_ca_in_233;
wire [242:0] u_ca_in_234;
wire [242:0] u_ca_in_235;
wire [242:0] u_ca_in_236;
wire [242:0] u_ca_in_237;
wire [242:0] u_ca_in_238;
wire [242:0] u_ca_in_239;
wire [242:0] u_ca_in_240;
wire [242:0] u_ca_in_241;
wire [242:0] u_ca_in_242;
wire [242:0] u_ca_in_243;
wire [242:0] u_ca_in_244;
wire [242:0] u_ca_in_245;
wire [242:0] u_ca_in_246;
wire [242:0] u_ca_in_247;
wire [242:0] u_ca_in_248;
wire [242:0] u_ca_in_249;
wire [242:0] u_ca_in_250;
wire [242:0] u_ca_in_251;
wire [242:0] u_ca_in_252;
wire [242:0] u_ca_in_253;
wire [242:0] u_ca_in_254;
wire [242:0] u_ca_in_255;
wire [242:0] u_ca_in_256;
wire [242:0] u_ca_in_257;
wire [242:0] u_ca_in_258;
wire [242:0] u_ca_in_259;
wire [242:0] u_ca_in_260;
wire [242:0] u_ca_in_261;
wire [242:0] u_ca_in_262;
wire [242:0] u_ca_in_263;
wire [242:0] u_ca_in_264;
wire [242:0] u_ca_in_265;
wire [242:0] u_ca_in_266;
wire [242:0] u_ca_in_267;
wire [242:0] u_ca_in_268;
wire [242:0] u_ca_in_269;
wire [242:0] u_ca_in_270;
wire [242:0] u_ca_in_271;
wire [242:0] u_ca_in_272;
wire [242:0] u_ca_in_273;
wire [242:0] u_ca_in_274;
wire [242:0] u_ca_in_275;
wire [242:0] u_ca_in_276;
wire [242:0] u_ca_in_277;
wire [242:0] u_ca_in_278;
wire [242:0] u_ca_in_279;
wire [242:0] u_ca_in_280;
wire [242:0] u_ca_in_281;
wire [242:0] u_ca_in_282;
wire [242:0] u_ca_in_283;
wire [242:0] u_ca_in_284;
wire [242:0] u_ca_in_285;
wire [242:0] u_ca_in_286;
wire [242:0] u_ca_in_287;
wire [242:0] u_ca_in_288;
wire [242:0] u_ca_in_289;
wire [242:0] u_ca_in_290;
wire [242:0] u_ca_in_291;
wire [242:0] u_ca_in_292;
wire [242:0] u_ca_in_293;
wire [242:0] u_ca_in_294;
wire [242:0] u_ca_in_295;
wire [242:0] u_ca_in_296;
wire [242:0] u_ca_in_297;
wire [242:0] u_ca_in_298;
wire [242:0] u_ca_in_299;
wire [242:0] u_ca_in_300;
wire [242:0] u_ca_in_301;
wire [242:0] u_ca_in_302;
wire [242:0] u_ca_in_303;
wire [242:0] u_ca_in_304;
wire [242:0] u_ca_in_305;
wire [242:0] u_ca_in_306;
wire [242:0] u_ca_in_307;
wire [242:0] u_ca_in_308;
wire [242:0] u_ca_in_309;
wire [242:0] u_ca_in_310;
wire [242:0] u_ca_in_311;
wire [242:0] u_ca_in_312;
wire [242:0] u_ca_in_313;
wire [242:0] u_ca_in_314;
wire [242:0] u_ca_in_315;
wire [242:0] u_ca_in_316;
wire [242:0] u_ca_in_317;
wire [242:0] u_ca_in_318;
wire [242:0] u_ca_in_319;
wire [242:0] u_ca_in_320;
wire [242:0] u_ca_in_321;
wire [242:0] u_ca_in_322;
wire [242:0] u_ca_in_323;
wire [242:0] u_ca_in_324;
wire [242:0] u_ca_in_325;
wire [242:0] u_ca_in_326;
wire [242:0] u_ca_in_327;
wire [242:0] u_ca_in_328;
wire [242:0] u_ca_in_329;
wire [242:0] u_ca_in_330;
wire [242:0] u_ca_in_331;
wire [242:0] u_ca_in_332;
wire [242:0] u_ca_in_333;
wire [242:0] u_ca_in_334;
wire [242:0] u_ca_in_335;
wire [242:0] u_ca_in_336;
wire [242:0] u_ca_in_337;
wire [242:0] u_ca_in_338;
wire [242:0] u_ca_in_339;
wire [242:0] u_ca_in_340;
wire [242:0] u_ca_in_341;
wire [242:0] u_ca_in_342;
wire [242:0] u_ca_in_343;
wire [242:0] u_ca_in_344;
wire [242:0] u_ca_in_345;
wire [242:0] u_ca_in_346;
wire [242:0] u_ca_in_347;
wire [242:0] u_ca_in_348;
wire [242:0] u_ca_in_349;
wire [242:0] u_ca_in_350;
wire [242:0] u_ca_in_351;
wire [242:0] u_ca_in_352;
wire [242:0] u_ca_in_353;
wire [242:0] u_ca_in_354;
wire [242:0] u_ca_in_355;
wire [242:0] u_ca_in_356;
wire [242:0] u_ca_in_357;
wire [242:0] u_ca_in_358;
wire [242:0] u_ca_in_359;
wire [242:0] u_ca_in_360;
wire [242:0] u_ca_in_361;
wire [242:0] u_ca_in_362;
wire [242:0] u_ca_in_363;
wire [242:0] u_ca_in_364;
wire [242:0] u_ca_in_365;
wire [242:0] u_ca_in_366;
wire [242:0] u_ca_in_367;
wire [242:0] u_ca_in_368;
wire [242:0] u_ca_in_369;
wire [242:0] u_ca_in_370;
wire [242:0] u_ca_in_371;
wire [242:0] u_ca_in_372;
wire [242:0] u_ca_in_373;
wire [242:0] u_ca_in_374;
wire [242:0] u_ca_in_375;
wire [242:0] u_ca_in_376;
wire [242:0] u_ca_in_377;
wire [242:0] u_ca_in_378;
wire [242:0] u_ca_in_379;
wire [242:0] u_ca_in_380;
wire [242:0] u_ca_in_381;
wire [242:0] u_ca_in_382;
wire [242:0] u_ca_in_383;
wire [242:0] u_ca_in_384;
wire [242:0] u_ca_in_385;
wire [242:0] u_ca_in_386;
wire [242:0] u_ca_in_387;
wire [242:0] u_ca_in_388;
wire [242:0] u_ca_in_389;
wire [242:0] u_ca_in_390;
wire [242:0] u_ca_in_391;
wire [242:0] u_ca_in_392;
wire [242:0] u_ca_in_393;
wire [242:0] u_ca_in_394;
wire [242:0] u_ca_in_395;
wire [242:0] u_ca_in_396;
wire [242:0] u_ca_in_397;
wire [242:0] u_ca_in_398;
wire [242:0] u_ca_in_399;
wire [242:0] u_ca_in_400;
wire [242:0] u_ca_in_401;
wire [242:0] u_ca_in_402;
wire [242:0] u_ca_in_403;
wire [242:0] u_ca_in_404;
wire [242:0] u_ca_in_405;
wire [242:0] u_ca_in_406;
wire [242:0] u_ca_in_407;
wire [242:0] u_ca_in_408;
wire [242:0] u_ca_in_409;
wire [242:0] u_ca_in_410;
wire [242:0] u_ca_in_411;
wire [242:0] u_ca_in_412;
wire [242:0] u_ca_in_413;
wire [242:0] u_ca_in_414;
wire [242:0] u_ca_in_415;
wire [242:0] u_ca_in_416;
wire [242:0] u_ca_in_417;
wire [242:0] u_ca_in_418;
wire [242:0] u_ca_in_419;
wire [242:0] u_ca_in_420;
wire [242:0] u_ca_in_421;
wire [242:0] u_ca_in_422;
wire [242:0] u_ca_in_423;
wire [242:0] u_ca_in_424;
wire [242:0] u_ca_in_425;
wire [242:0] u_ca_in_426;
wire [242:0] u_ca_in_427;
wire [242:0] u_ca_in_428;
wire [242:0] u_ca_in_429;
wire [242:0] u_ca_in_430;
wire [242:0] u_ca_in_431;
wire [242:0] u_ca_in_432;
wire [242:0] u_ca_in_433;
wire [242:0] u_ca_in_434;
wire [242:0] u_ca_in_435;
wire [242:0] u_ca_in_436;
wire [242:0] u_ca_in_437;
wire [242:0] u_ca_in_438;
wire [242:0] u_ca_in_439;
wire [242:0] u_ca_in_440;
wire [242:0] u_ca_in_441;
wire [242:0] u_ca_in_442;
wire [242:0] u_ca_in_443;
wire [242:0] u_ca_in_444;
wire [242:0] u_ca_in_445;
wire [242:0] u_ca_in_446;
wire [242:0] u_ca_in_447;
wire [242:0] u_ca_in_448;
wire [242:0] u_ca_in_449;
wire [242:0] u_ca_in_450;
wire [242:0] u_ca_in_451;
wire [242:0] u_ca_in_452;
wire [242:0] u_ca_in_453;
wire [242:0] u_ca_in_454;
wire [242:0] u_ca_in_455;
wire [242:0] u_ca_in_456;
wire [242:0] u_ca_in_457;
wire [242:0] u_ca_in_458;
wire [242:0] u_ca_in_459;
wire [242:0] u_ca_in_460;
wire [242:0] u_ca_in_461;
wire [242:0] u_ca_in_462;
wire [242:0] u_ca_in_463;
wire [242:0] u_ca_in_464;
wire [242:0] u_ca_in_465;
wire [242:0] u_ca_in_466;
wire [242:0] u_ca_in_467;
wire [242:0] u_ca_in_468;
wire [242:0] u_ca_in_469;
wire [242:0] u_ca_in_470;
wire [242:0] u_ca_in_471;
wire [242:0] u_ca_in_472;
wire [242:0] u_ca_in_473;
wire [242:0] u_ca_in_474;
wire [242:0] u_ca_in_475;
wire [242:0] u_ca_in_476;
wire [242:0] u_ca_in_477;
wire [242:0] u_ca_in_478;
wire [242:0] u_ca_in_479;
wire [242:0] u_ca_in_480;
wire [242:0] u_ca_in_481;
wire [242:0] u_ca_in_482;
wire [242:0] u_ca_in_483;
wire [242:0] u_ca_in_484;
wire [242:0] u_ca_in_485;
wire [242:0] u_ca_in_486;
wire [242:0] u_ca_in_487;
wire [242:0] u_ca_in_488;
wire [242:0] u_ca_in_489;
wire [242:0] u_ca_in_490;
wire [242:0] u_ca_in_491;
wire [242:0] u_ca_in_492;
wire [242:0] u_ca_in_493;
wire [242:0] u_ca_in_494;
wire [242:0] u_ca_in_495;
wire [242:0] u_ca_in_496;
wire [242:0] u_ca_in_497;
wire [242:0] u_ca_in_498;
wire [242:0] u_ca_in_499;
wire [242:0] u_ca_in_500;
wire [242:0] u_ca_in_501;
wire [242:0] u_ca_in_502;
wire [242:0] u_ca_in_503;
wire [242:0] u_ca_in_504;
wire [242:0] u_ca_in_505;
wire [242:0] u_ca_in_506;
wire [242:0] u_ca_in_507;
wire [242:0] u_ca_in_508;
wire [242:0] u_ca_in_509;
wire [242:0] u_ca_in_510;
wire [242:0] u_ca_in_511;
wire [242:0] u_ca_in_512;
wire [242:0] u_ca_in_513;
wire [242:0] u_ca_in_514;
wire [242:0] u_ca_in_515;
wire [242:0] u_ca_in_516;
wire [242:0] u_ca_in_517;
wire [242:0] u_ca_in_518;
wire [242:0] u_ca_in_519;
wire [242:0] u_ca_in_520;
wire [242:0] u_ca_in_521;
wire [242:0] u_ca_in_522;
wire [242:0] u_ca_in_523;
wire [242:0] u_ca_in_524;
wire [242:0] u_ca_in_525;
wire [242:0] u_ca_in_526;
wire [242:0] u_ca_in_527;
wire [242:0] u_ca_in_528;
wire [242:0] u_ca_in_529;
wire [242:0] u_ca_in_530;
wire [242:0] u_ca_in_531;
wire [242:0] u_ca_in_532;
wire [242:0] u_ca_in_533;
wire [242:0] u_ca_in_534;
wire [242:0] u_ca_in_535;
wire [242:0] u_ca_in_536;
wire [242:0] u_ca_in_537;
wire [242:0] u_ca_in_538;
wire [242:0] u_ca_in_539;
wire [242:0] u_ca_in_540;
wire [242:0] u_ca_in_541;
wire [242:0] u_ca_in_542;
wire [242:0] u_ca_in_543;
wire [242:0] u_ca_in_544;
wire [242:0] u_ca_in_545;
wire [242:0] u_ca_in_546;
wire [242:0] u_ca_in_547;
wire [242:0] u_ca_in_548;
wire [242:0] u_ca_in_549;
wire [242:0] u_ca_in_550;
wire [242:0] u_ca_in_551;
wire [242:0] u_ca_in_552;
wire [242:0] u_ca_in_553;
wire [242:0] u_ca_in_554;
wire [242:0] u_ca_in_555;
wire [242:0] u_ca_in_556;
wire [242:0] u_ca_in_557;
wire [242:0] u_ca_in_558;
wire [242:0] u_ca_in_559;
wire [242:0] u_ca_in_560;
wire [242:0] u_ca_in_561;
wire [242:0] u_ca_in_562;
wire [242:0] u_ca_in_563;
wire [242:0] u_ca_in_564;
wire [242:0] u_ca_in_565;
wire [242:0] u_ca_in_566;
wire [242:0] u_ca_in_567;
wire [242:0] u_ca_in_568;
wire [242:0] u_ca_in_569;
wire [242:0] u_ca_in_570;
wire [242:0] u_ca_in_571;
wire [242:0] u_ca_in_572;
wire [242:0] u_ca_in_573;
wire [242:0] u_ca_in_574;
wire [242:0] u_ca_in_575;
wire [242:0] u_ca_in_576;
wire [242:0] u_ca_in_577;
wire [242:0] u_ca_in_578;
wire [242:0] u_ca_in_579;
wire [242:0] u_ca_in_580;
wire [242:0] u_ca_in_581;
wire [242:0] u_ca_in_582;
wire [242:0] u_ca_in_583;
wire [242:0] u_ca_in_584;
wire [242:0] u_ca_in_585;
wire [242:0] u_ca_in_586;
wire [242:0] u_ca_in_587;
wire [242:0] u_ca_in_588;
wire [242:0] u_ca_in_589;
wire [242:0] u_ca_in_590;
wire [242:0] u_ca_in_591;
wire [242:0] u_ca_in_592;
wire [242:0] u_ca_in_593;
wire [242:0] u_ca_in_594;
wire [242:0] u_ca_in_595;
wire [242:0] u_ca_in_596;
wire [242:0] u_ca_in_597;
wire [242:0] u_ca_in_598;
wire [242:0] u_ca_in_599;
wire [242:0] u_ca_in_600;
wire [242:0] u_ca_in_601;
wire [242:0] u_ca_in_602;
wire [242:0] u_ca_in_603;
wire [242:0] u_ca_in_604;
wire [242:0] u_ca_in_605;
wire [242:0] u_ca_in_606;
wire [242:0] u_ca_in_607;
wire [242:0] u_ca_in_608;
wire [242:0] u_ca_in_609;
wire [242:0] u_ca_in_610;
wire [242:0] u_ca_in_611;
wire [242:0] u_ca_in_612;
wire [242:0] u_ca_in_613;
wire [242:0] u_ca_in_614;
wire [242:0] u_ca_in_615;
wire [242:0] u_ca_in_616;
wire [242:0] u_ca_in_617;
wire [242:0] u_ca_in_618;
wire [242:0] u_ca_in_619;
wire [242:0] u_ca_in_620;
wire [242:0] u_ca_in_621;
wire [242:0] u_ca_in_622;
wire [242:0] u_ca_in_623;
wire [242:0] u_ca_in_624;
wire [242:0] u_ca_in_625;
wire [242:0] u_ca_in_626;
wire [242:0] u_ca_in_627;
wire [242:0] u_ca_in_628;
wire [242:0] u_ca_in_629;
wire [242:0] u_ca_in_630;
wire [242:0] u_ca_in_631;
wire [242:0] u_ca_in_632;
wire [242:0] u_ca_in_633;
wire [242:0] u_ca_in_634;
wire [242:0] u_ca_in_635;
wire [242:0] u_ca_in_636;
wire [242:0] u_ca_in_637;
wire [242:0] u_ca_in_638;
wire [242:0] u_ca_in_639;
wire [242:0] u_ca_in_640;
wire [242:0] u_ca_in_641;
wire [242:0] u_ca_in_642;
wire [242:0] u_ca_in_643;
wire [242:0] u_ca_in_644;
wire [242:0] u_ca_in_645;
wire [242:0] u_ca_in_646;
wire [242:0] u_ca_in_647;
wire [242:0] u_ca_in_648;
wire [242:0] u_ca_in_649;
wire [242:0] u_ca_in_650;
wire [242:0] u_ca_in_651;
wire [242:0] u_ca_in_652;
wire [242:0] u_ca_in_653;
wire [242:0] u_ca_in_654;
wire [242:0] u_ca_in_655;
wire [242:0] u_ca_in_656;
wire [242:0] u_ca_in_657;
wire [242:0] u_ca_in_658;
wire [242:0] u_ca_in_659;
wire [242:0] u_ca_in_660;
wire [242:0] u_ca_in_661;
wire [242:0] u_ca_in_662;
wire [242:0] u_ca_in_663;
wire [242:0] u_ca_in_664;
wire [242:0] u_ca_in_665;
wire [242:0] u_ca_in_666;
wire [242:0] u_ca_in_667;
wire [242:0] u_ca_in_668;
wire [242:0] u_ca_in_669;
wire [242:0] u_ca_in_670;
wire [242:0] u_ca_in_671;
wire [242:0] u_ca_in_672;
wire [242:0] u_ca_in_673;
wire [242:0] u_ca_in_674;
wire [242:0] u_ca_in_675;
wire [242:0] u_ca_in_676;
wire [242:0] u_ca_in_677;
wire [242:0] u_ca_in_678;
wire [242:0] u_ca_in_679;
wire [242:0] u_ca_in_680;
wire [242:0] u_ca_in_681;
wire [242:0] u_ca_in_682;
wire [242:0] u_ca_in_683;
wire [242:0] u_ca_in_684;
wire [242:0] u_ca_in_685;
wire [242:0] u_ca_in_686;
wire [242:0] u_ca_in_687;
wire [242:0] u_ca_in_688;
wire [242:0] u_ca_in_689;
wire [242:0] u_ca_in_690;
wire [242:0] u_ca_in_691;
wire [242:0] u_ca_in_692;
wire [242:0] u_ca_in_693;
wire [242:0] u_ca_in_694;
wire [242:0] u_ca_in_695;
wire [242:0] u_ca_in_696;
wire [242:0] u_ca_in_697;
wire [242:0] u_ca_in_698;
wire [242:0] u_ca_in_699;
wire [242:0] u_ca_in_700;
wire [242:0] u_ca_in_701;
wire [242:0] u_ca_in_702;
wire [242:0] u_ca_in_703;
wire [242:0] u_ca_in_704;
wire [242:0] u_ca_in_705;
wire [242:0] u_ca_in_706;
wire [242:0] u_ca_in_707;
wire [242:0] u_ca_in_708;
wire [242:0] u_ca_in_709;
wire [242:0] u_ca_in_710;
wire [242:0] u_ca_in_711;
wire [242:0] u_ca_in_712;
wire [242:0] u_ca_in_713;
wire [242:0] u_ca_in_714;
wire [242:0] u_ca_in_715;
wire [242:0] u_ca_in_716;
wire [242:0] u_ca_in_717;
wire [242:0] u_ca_in_718;
wire [242:0] u_ca_in_719;
wire [242:0] u_ca_in_720;
wire [242:0] u_ca_in_721;
wire [242:0] u_ca_in_722;
wire [242:0] u_ca_in_723;
wire [242:0] u_ca_in_724;
wire [242:0] u_ca_in_725;
wire [242:0] u_ca_in_726;
wire [242:0] u_ca_in_727;
wire [242:0] u_ca_in_728;
wire [242:0] u_ca_in_729;
wire [242:0] u_ca_in_730;
wire [242:0] u_ca_in_731;
wire [242:0] u_ca_in_732;
wire [242:0] u_ca_in_733;
wire [242:0] u_ca_in_734;
wire [242:0] u_ca_in_735;
wire [242:0] u_ca_in_736;
wire [242:0] u_ca_in_737;
wire [242:0] u_ca_in_738;
wire [242:0] u_ca_in_739;
wire [242:0] u_ca_in_740;
wire [242:0] u_ca_in_741;
wire [242:0] u_ca_in_742;
wire [242:0] u_ca_in_743;
wire [242:0] u_ca_in_744;
wire [242:0] u_ca_in_745;
wire [242:0] u_ca_in_746;
wire [242:0] u_ca_in_747;
wire [242:0] u_ca_in_748;
wire [242:0] u_ca_in_749;
wire [242:0] u_ca_in_750;
wire [242:0] u_ca_in_751;
wire [242:0] u_ca_in_752;
wire [242:0] u_ca_in_753;
wire [242:0] u_ca_in_754;
wire [242:0] u_ca_in_755;
wire [242:0] u_ca_in_756;
wire [242:0] u_ca_in_757;
wire [242:0] u_ca_in_758;
wire [242:0] u_ca_in_759;
wire [242:0] u_ca_in_760;
wire [242:0] u_ca_in_761;
wire [242:0] u_ca_in_762;
wire [242:0] u_ca_in_763;
wire [242:0] u_ca_in_764;
wire [242:0] u_ca_in_765;
wire [242:0] u_ca_in_766;
wire [242:0] u_ca_in_767;
wire [242:0] u_ca_in_768;
wire [242:0] u_ca_in_769;
wire [242:0] u_ca_in_770;
wire [242:0] u_ca_in_771;
wire [242:0] u_ca_in_772;
wire [242:0] u_ca_in_773;
wire [242:0] u_ca_in_774;
wire [242:0] u_ca_in_775;
wire [242:0] u_ca_in_776;
wire [242:0] u_ca_in_777;
wire [242:0] u_ca_in_778;
wire [242:0] u_ca_in_779;
wire [242:0] u_ca_in_780;
wire [242:0] u_ca_in_781;
wire [242:0] u_ca_in_782;
wire [242:0] u_ca_in_783;
wire [242:0] u_ca_in_784;
wire [242:0] u_ca_in_785;
wire [242:0] u_ca_in_786;
wire [242:0] u_ca_in_787;
wire [242:0] u_ca_in_788;
wire [242:0] u_ca_in_789;
wire [242:0] u_ca_in_790;
wire [242:0] u_ca_in_791;
wire [242:0] u_ca_in_792;
wire [242:0] u_ca_in_793;
wire [242:0] u_ca_in_794;
wire [242:0] u_ca_in_795;
wire [242:0] u_ca_in_796;
wire [242:0] u_ca_in_797;
wire [242:0] u_ca_in_798;
wire [242:0] u_ca_in_799;
wire [242:0] u_ca_in_800;
wire [242:0] u_ca_in_801;
wire [242:0] u_ca_in_802;
wire [242:0] u_ca_in_803;
wire [242:0] u_ca_in_804;
wire [242:0] u_ca_in_805;
wire [242:0] u_ca_in_806;
wire [242:0] u_ca_in_807;
wire [242:0] u_ca_in_808;
wire [242:0] u_ca_in_809;
wire [242:0] u_ca_in_810;
wire [242:0] u_ca_in_811;
wire [242:0] u_ca_in_812;
wire [242:0] u_ca_in_813;
wire [242:0] u_ca_in_814;
wire [242:0] u_ca_in_815;
wire [242:0] u_ca_in_816;
wire [242:0] u_ca_in_817;
wire [242:0] u_ca_in_818;
wire [242:0] u_ca_in_819;
wire [242:0] u_ca_in_820;
wire [242:0] u_ca_in_821;
wire [242:0] u_ca_in_822;
wire [242:0] u_ca_in_823;
wire [242:0] u_ca_in_824;
wire [242:0] u_ca_in_825;
wire [242:0] u_ca_in_826;
wire [242:0] u_ca_in_827;
wire [242:0] u_ca_in_828;
wire [242:0] u_ca_in_829;
wire [242:0] u_ca_in_830;
wire [242:0] u_ca_in_831;
wire [242:0] u_ca_in_832;
wire [242:0] u_ca_in_833;
wire [242:0] u_ca_in_834;
wire [242:0] u_ca_in_835;
wire [242:0] u_ca_in_836;
wire [242:0] u_ca_in_837;
wire [242:0] u_ca_in_838;
wire [242:0] u_ca_in_839;
wire [242:0] u_ca_in_840;
wire [242:0] u_ca_in_841;
wire [242:0] u_ca_in_842;
wire [242:0] u_ca_in_843;
wire [242:0] u_ca_in_844;
wire [242:0] u_ca_in_845;
wire [242:0] u_ca_in_846;
wire [242:0] u_ca_in_847;
wire [242:0] u_ca_in_848;
wire [242:0] u_ca_in_849;
wire [242:0] u_ca_in_850;
wire [242:0] u_ca_in_851;
wire [242:0] u_ca_in_852;
wire [242:0] u_ca_in_853;
wire [242:0] u_ca_in_854;
wire [242:0] u_ca_in_855;
wire [242:0] u_ca_in_856;
wire [242:0] u_ca_in_857;
wire [242:0] u_ca_in_858;
wire [242:0] u_ca_in_859;
wire [242:0] u_ca_in_860;
wire [242:0] u_ca_in_861;
wire [242:0] u_ca_in_862;
wire [242:0] u_ca_in_863;
wire [242:0] u_ca_in_864;
wire [242:0] u_ca_in_865;
wire [242:0] u_ca_in_866;
wire [242:0] u_ca_in_867;
wire [242:0] u_ca_in_868;
wire [242:0] u_ca_in_869;
wire [242:0] u_ca_in_870;
wire [242:0] u_ca_in_871;
wire [242:0] u_ca_in_872;
wire [242:0] u_ca_in_873;
wire [242:0] u_ca_in_874;
wire [242:0] u_ca_in_875;
wire [242:0] u_ca_in_876;
wire [242:0] u_ca_in_877;
wire [242:0] u_ca_in_878;
wire [242:0] u_ca_in_879;
wire [242:0] u_ca_in_880;
wire [242:0] u_ca_in_881;
wire [242:0] u_ca_in_882;
wire [242:0] u_ca_in_883;
wire [242:0] u_ca_in_884;
wire [242:0] u_ca_in_885;
wire [242:0] u_ca_in_886;
wire [242:0] u_ca_in_887;
wire [242:0] u_ca_in_888;
wire [242:0] u_ca_in_889;
wire [242:0] u_ca_in_890;
wire [242:0] u_ca_in_891;
wire [242:0] u_ca_in_892;
wire [242:0] u_ca_in_893;
wire [242:0] u_ca_in_894;
wire [242:0] u_ca_in_895;
wire [242:0] u_ca_in_896;
wire [242:0] u_ca_in_897;
wire [242:0] u_ca_in_898;
wire [242:0] u_ca_in_899;
wire [242:0] u_ca_in_900;
wire [242:0] u_ca_in_901;
wire [242:0] u_ca_in_902;
wire [242:0] u_ca_in_903;
wire [242:0] u_ca_in_904;
wire [242:0] u_ca_in_905;
wire [242:0] u_ca_in_906;
wire [242:0] u_ca_in_907;
wire [242:0] u_ca_in_908;
wire [242:0] u_ca_in_909;
wire [242:0] u_ca_in_910;
wire [242:0] u_ca_in_911;
wire [242:0] u_ca_in_912;
wire [242:0] u_ca_in_913;
wire [242:0] u_ca_in_914;
wire [242:0] u_ca_in_915;
wire [242:0] u_ca_in_916;
wire [242:0] u_ca_in_917;
wire [242:0] u_ca_in_918;
wire [242:0] u_ca_in_919;
wire [242:0] u_ca_in_920;
wire [242:0] u_ca_in_921;
wire [242:0] u_ca_in_922;
wire [242:0] u_ca_in_923;
wire [242:0] u_ca_in_924;
wire [242:0] u_ca_in_925;
wire [242:0] u_ca_in_926;
wire [242:0] u_ca_in_927;
wire [242:0] u_ca_in_928;
wire [242:0] u_ca_in_929;
wire [242:0] u_ca_in_930;
wire [242:0] u_ca_in_931;
wire [242:0] u_ca_in_932;
wire [242:0] u_ca_in_933;
wire [242:0] u_ca_in_934;
wire [242:0] u_ca_in_935;
wire [242:0] u_ca_in_936;
wire [242:0] u_ca_in_937;
wire [242:0] u_ca_in_938;
wire [242:0] u_ca_in_939;
wire [242:0] u_ca_in_940;
wire [242:0] u_ca_in_941;
wire [242:0] u_ca_in_942;
wire [242:0] u_ca_in_943;
wire [242:0] u_ca_in_944;
wire [242:0] u_ca_in_945;
wire [242:0] u_ca_in_946;
wire [242:0] u_ca_in_947;
wire [242:0] u_ca_in_948;
wire [242:0] u_ca_in_949;
wire [242:0] u_ca_in_950;
wire [242:0] u_ca_in_951;
wire [242:0] u_ca_in_952;
wire [242:0] u_ca_in_953;
wire [242:0] u_ca_in_954;
wire [242:0] u_ca_in_955;
wire [242:0] u_ca_in_956;
wire [242:0] u_ca_in_957;
wire [242:0] u_ca_in_958;
wire [242:0] u_ca_in_959;
wire [242:0] u_ca_in_960;
wire [242:0] u_ca_in_961;
wire [242:0] u_ca_in_962;
wire [242:0] u_ca_in_963;
wire [242:0] u_ca_in_964;
wire [242:0] u_ca_in_965;
wire [242:0] u_ca_in_966;
wire [242:0] u_ca_in_967;
wire [242:0] u_ca_in_968;
wire [242:0] u_ca_in_969;
wire [242:0] u_ca_in_970;
wire [242:0] u_ca_in_971;
wire [242:0] u_ca_in_972;
wire [242:0] u_ca_in_973;
wire [242:0] u_ca_in_974;
wire [242:0] u_ca_in_975;
wire [242:0] u_ca_in_976;
wire [242:0] u_ca_in_977;
wire [242:0] u_ca_in_978;
wire [242:0] u_ca_in_979;
wire [242:0] u_ca_in_980;
wire [242:0] u_ca_in_981;
wire [242:0] u_ca_in_982;
wire [242:0] u_ca_in_983;
wire [242:0] u_ca_in_984;
wire [242:0] u_ca_in_985;
wire [242:0] u_ca_in_986;
wire [242:0] u_ca_in_987;
wire [242:0] u_ca_in_988;
wire [242:0] u_ca_in_989;
wire [242:0] u_ca_in_990;
wire [242:0] u_ca_in_991;
wire [242:0] u_ca_in_992;
wire [242:0] u_ca_in_993;
wire [242:0] u_ca_in_994;
wire [242:0] u_ca_in_995;
wire [242:0] u_ca_in_996;
wire [242:0] u_ca_in_997;
wire [242:0] u_ca_in_998;
wire [242:0] u_ca_in_999;
wire [242:0] u_ca_in_1000;
wire [242:0] u_ca_in_1001;
wire [242:0] u_ca_in_1002;
wire [242:0] u_ca_in_1003;
wire [242:0] u_ca_in_1004;
wire [242:0] u_ca_in_1005;
wire [242:0] u_ca_in_1006;
wire [242:0] u_ca_in_1007;
wire [242:0] u_ca_in_1008;
wire [242:0] u_ca_in_1009;
wire [242:0] u_ca_in_1010;
wire [242:0] u_ca_in_1011;
wire [242:0] u_ca_in_1012;
wire [242:0] u_ca_in_1013;
wire [242:0] u_ca_in_1014;
wire [242:0] u_ca_in_1015;
wire [242:0] u_ca_in_1016;
wire [242:0] u_ca_in_1017;
wire [242:0] u_ca_in_1018;
wire [242:0] u_ca_in_1019;
wire [242:0] u_ca_in_1020;
wire [242:0] u_ca_in_1021;
wire [242:0] u_ca_in_1022;
wire [242:0] u_ca_in_1023;
wire [242:0] u_ca_in_1024;
wire [242:0] u_ca_in_1025;
wire [242:0] u_ca_in_1026;
wire [242:0] u_ca_in_1027;
wire [242:0] u_ca_in_1028;
wire [242:0] u_ca_in_1029;
wire [242:0] u_ca_in_1030;
wire [242:0] u_ca_in_1031;
wire [242:0] u_ca_in_1032;
wire [242:0] u_ca_in_1033;
wire [242:0] u_ca_in_1034;
wire [242:0] u_ca_in_1035;
wire [242:0] u_ca_in_1036;
wire [242:0] u_ca_in_1037;
wire [242:0] u_ca_in_1038;
wire [242:0] u_ca_in_1039;
wire [242:0] u_ca_in_1040;
wire [242:0] u_ca_in_1041;
wire [242:0] u_ca_in_1042;
wire [242:0] u_ca_in_1043;
wire [242:0] u_ca_in_1044;
wire [242:0] u_ca_in_1045;
wire [242:0] u_ca_in_1046;
wire [242:0] u_ca_in_1047;
wire [242:0] u_ca_in_1048;
wire [242:0] u_ca_in_1049;
wire [242:0] u_ca_in_1050;
wire [242:0] u_ca_in_1051;
wire [242:0] u_ca_in_1052;
wire [242:0] u_ca_in_1053;
wire [242:0] u_ca_in_1054;
wire [242:0] u_ca_in_1055;
wire [242:0] u_ca_in_1056;
wire [242:0] u_ca_in_1057;
wire [242:0] u_ca_in_1058;
wire [242:0] u_ca_in_1059;
wire [242:0] u_ca_in_1060;
wire [242:0] u_ca_in_1061;
wire [242:0] u_ca_in_1062;
wire [242:0] u_ca_in_1063;
wire [242:0] u_ca_in_1064;
wire [242:0] u_ca_in_1065;
wire [242:0] u_ca_in_1066;
wire [242:0] u_ca_in_1067;
wire [242:0] u_ca_in_1068;
wire [242:0] u_ca_in_1069;
wire [242:0] u_ca_in_1070;
wire [242:0] u_ca_in_1071;
wire [242:0] u_ca_in_1072;
wire [242:0] u_ca_in_1073;
wire [242:0] u_ca_in_1074;
wire [242:0] u_ca_in_1075;
wire [242:0] u_ca_in_1076;
wire [242:0] u_ca_in_1077;
wire [242:0] u_ca_in_1078;
wire [242:0] u_ca_in_1079;
wire [242:0] u_ca_in_1080;
wire [242:0] u_ca_in_1081;
wire [242:0] u_ca_in_1082;
wire [242:0] u_ca_in_1083;
wire [242:0] u_ca_in_1084;
wire [242:0] u_ca_in_1085;
wire [242:0] u_ca_in_1086;
wire [242:0] u_ca_in_1087;
wire [242:0] u_ca_in_1088;
wire [242:0] u_ca_in_1089;
wire [242:0] u_ca_in_1090;
wire [242:0] u_ca_in_1091;
wire [242:0] u_ca_in_1092;
wire [242:0] u_ca_in_1093;
wire [242:0] u_ca_in_1094;
wire [242:0] u_ca_in_1095;
wire [242:0] u_ca_in_1096;
wire [242:0] u_ca_in_1097;
wire [242:0] u_ca_in_1098;
wire [242:0] u_ca_in_1099;
wire [242:0] u_ca_in_1100;
wire [242:0] u_ca_in_1101;
wire [242:0] u_ca_in_1102;
wire [242:0] u_ca_in_1103;
wire [242:0] u_ca_in_1104;
wire [242:0] u_ca_in_1105;
wire [242:0] u_ca_in_1106;
wire [242:0] u_ca_in_1107;
wire [242:0] u_ca_in_1108;
wire [242:0] u_ca_in_1109;
wire [242:0] u_ca_in_1110;
wire [242:0] u_ca_in_1111;
wire [242:0] u_ca_in_1112;
wire [242:0] u_ca_in_1113;
wire [242:0] u_ca_in_1114;
wire [242:0] u_ca_in_1115;
wire [242:0] u_ca_in_1116;
wire [242:0] u_ca_in_1117;
wire [242:0] u_ca_in_1118;
wire [242:0] u_ca_in_1119;
wire [242:0] u_ca_in_1120;
wire [242:0] u_ca_in_1121;
wire [242:0] u_ca_in_1122;
wire [242:0] u_ca_in_1123;
wire [242:0] u_ca_in_1124;
wire [242:0] u_ca_in_1125;
wire [242:0] u_ca_in_1126;
wire [242:0] u_ca_in_1127;
wire [242:0] u_ca_in_1128;
wire [242:0] u_ca_in_1129;
wire [242:0] u_ca_in_1130;
wire [242:0] u_ca_in_1131;
wire [242:0] u_ca_in_1132;
wire [242:0] u_ca_in_1133;
wire [242:0] u_ca_in_1134;
wire [242:0] u_ca_in_1135;
wire [242:0] u_ca_in_1136;
wire [242:0] u_ca_in_1137;
wire [242:0] u_ca_in_1138;
wire [242:0] u_ca_in_1139;
wire [242:0] u_ca_in_1140;
wire [242:0] u_ca_in_1141;
wire [242:0] u_ca_in_1142;
wire [242:0] u_ca_in_1143;
wire [242:0] u_ca_in_1144;
wire [242:0] u_ca_in_1145;
wire [242:0] u_ca_in_1146;
wire [242:0] u_ca_in_1147;
wire [242:0] u_ca_in_1148;
wire [242:0] u_ca_in_1149;
wire [242:0] u_ca_in_1150;
wire [242:0] u_ca_in_1151;
wire [242:0] u_ca_in_1152;
wire [242:0] u_ca_in_1153;
wire [242:0] u_ca_in_1154;
wire [242:0] u_ca_in_1155;
wire [242:0] u_ca_in_1156;
wire [242:0] u_ca_in_1157;
wire [242:0] u_ca_in_1158;
wire [242:0] u_ca_in_1159;
wire [242:0] u_ca_in_1160;
wire [242:0] u_ca_in_1161;
wire [242:0] u_ca_in_1162;
wire [242:0] u_ca_in_1163;
wire [242:0] u_ca_in_1164;
wire [242:0] u_ca_in_1165;
wire [242:0] u_ca_in_1166;
wire [242:0] u_ca_in_1167;
wire [242:0] u_ca_in_1168;
wire [242:0] u_ca_in_1169;
wire [242:0] u_ca_in_1170;
wire [242:0] u_ca_in_1171;
wire [242:0] u_ca_in_1172;
wire [242:0] u_ca_in_1173;
wire [242:0] u_ca_in_1174;
wire [242:0] u_ca_in_1175;
wire [242:0] u_ca_in_1176;
wire [242:0] u_ca_in_1177;
wire [242:0] u_ca_in_1178;
wire [242:0] u_ca_in_1179;
wire [242:0] u_ca_in_1180;
wire [242:0] u_ca_in_1181;
wire [242:0] u_ca_in_1182;
wire [242:0] u_ca_in_1183;
wire [242:0] u_ca_in_1184;
wire [242:0] u_ca_in_1185;
wire [242:0] u_ca_in_1186;
wire [242:0] u_ca_in_1187;
wire [242:0] u_ca_in_1188;
wire [242:0] u_ca_in_1189;
wire [242:0] u_ca_in_1190;
wire [242:0] u_ca_in_1191;
wire [242:0] u_ca_in_1192;
wire [242:0] u_ca_in_1193;
wire [242:0] u_ca_in_1194;
wire [242:0] u_ca_in_1195;
wire [242:0] u_ca_in_1196;
wire [242:0] u_ca_in_1197;
wire [242:0] u_ca_in_1198;
wire [242:0] u_ca_in_1199;
wire [242:0] u_ca_in_1200;
wire [242:0] u_ca_in_1201;
wire [242:0] u_ca_in_1202;
wire [242:0] u_ca_in_1203;
wire [242:0] u_ca_in_1204;
wire [242:0] u_ca_in_1205;
wire [242:0] u_ca_in_1206;
wire [242:0] u_ca_in_1207;
wire [242:0] u_ca_in_1208;
wire [242:0] u_ca_in_1209;
wire [242:0] u_ca_in_1210;
wire [242:0] u_ca_in_1211;
wire [242:0] u_ca_in_1212;
wire [242:0] u_ca_in_1213;
wire [242:0] u_ca_in_1214;
wire [242:0] u_ca_in_1215;
wire [242:0] u_ca_in_1216;
wire [242:0] u_ca_in_1217;
wire [242:0] u_ca_in_1218;
wire [242:0] u_ca_in_1219;
wire [242:0] u_ca_in_1220;
wire [242:0] u_ca_in_1221;
wire [242:0] u_ca_in_1222;
wire [242:0] u_ca_in_1223;
wire [242:0] u_ca_in_1224;
wire [242:0] u_ca_in_1225;
wire [242:0] u_ca_in_1226;
wire [242:0] u_ca_in_1227;
wire [242:0] u_ca_in_1228;
wire [242:0] u_ca_in_1229;
wire [242:0] u_ca_in_1230;
wire [242:0] u_ca_in_1231;
wire [242:0] u_ca_in_1232;
wire [242:0] u_ca_in_1233;
wire [242:0] u_ca_in_1234;
wire [242:0] u_ca_in_1235;
wire [242:0] u_ca_in_1236;
wire [242:0] u_ca_in_1237;
wire [242:0] u_ca_in_1238;
wire [242:0] u_ca_in_1239;
wire [242:0] u_ca_in_1240;
wire [242:0] u_ca_in_1241;
wire [242:0] u_ca_in_1242;
wire [242:0] u_ca_in_1243;
wire [242:0] u_ca_in_1244;
wire [242:0] u_ca_in_1245;
wire [242:0] u_ca_in_1246;
wire [242:0] u_ca_in_1247;
wire [242:0] u_ca_in_1248;
wire [242:0] u_ca_in_1249;
wire [242:0] u_ca_in_1250;
wire [242:0] u_ca_in_1251;
wire [242:0] u_ca_in_1252;
wire [242:0] u_ca_in_1253;
wire [242:0] u_ca_in_1254;
wire [242:0] u_ca_in_1255;
wire [242:0] u_ca_in_1256;
wire [242:0] u_ca_in_1257;
wire [242:0] u_ca_in_1258;
wire [242:0] u_ca_in_1259;
wire [242:0] u_ca_in_1260;
wire [242:0] u_ca_in_1261;
wire [242:0] u_ca_in_1262;
wire [242:0] u_ca_in_1263;
wire [242:0] u_ca_in_1264;
wire [242:0] u_ca_in_1265;
wire [242:0] u_ca_in_1266;
wire [242:0] u_ca_in_1267;
wire [242:0] u_ca_in_1268;
wire [242:0] u_ca_in_1269;
wire [242:0] u_ca_in_1270;
wire [242:0] u_ca_in_1271;
wire [242:0] u_ca_in_1272;
wire [242:0] u_ca_in_1273;
wire [242:0] u_ca_in_1274;
wire [242:0] u_ca_in_1275;
wire [242:0] u_ca_in_1276;
wire [242:0] u_ca_in_1277;
wire [242:0] u_ca_in_1278;
wire [242:0] u_ca_in_1279;


wire [71:0] u_ca_out_0;
wire [71:0] u_ca_out_1;
wire [71:0] u_ca_out_2;
wire [71:0] u_ca_out_3;
wire [71:0] u_ca_out_4;
wire [71:0] u_ca_out_5;
wire [71:0] u_ca_out_6;
wire [71:0] u_ca_out_7;
wire [71:0] u_ca_out_8;
wire [71:0] u_ca_out_9;
wire [71:0] u_ca_out_10;
wire [71:0] u_ca_out_11;
wire [71:0] u_ca_out_12;
wire [71:0] u_ca_out_13;
wire [71:0] u_ca_out_14;
wire [71:0] u_ca_out_15;
wire [71:0] u_ca_out_16;
wire [71:0] u_ca_out_17;
wire [71:0] u_ca_out_18;
wire [71:0] u_ca_out_19;
wire [71:0] u_ca_out_20;
wire [71:0] u_ca_out_21;
wire [71:0] u_ca_out_22;
wire [71:0] u_ca_out_23;
wire [71:0] u_ca_out_24;
wire [71:0] u_ca_out_25;
wire [71:0] u_ca_out_26;
wire [71:0] u_ca_out_27;
wire [71:0] u_ca_out_28;
wire [71:0] u_ca_out_29;
wire [71:0] u_ca_out_30;
wire [71:0] u_ca_out_31;
wire [71:0] u_ca_out_32;
wire [71:0] u_ca_out_33;
wire [71:0] u_ca_out_34;
wire [71:0] u_ca_out_35;
wire [71:0] u_ca_out_36;
wire [71:0] u_ca_out_37;
wire [71:0] u_ca_out_38;
wire [71:0] u_ca_out_39;
wire [71:0] u_ca_out_40;
wire [71:0] u_ca_out_41;
wire [71:0] u_ca_out_42;
wire [71:0] u_ca_out_43;
wire [71:0] u_ca_out_44;
wire [71:0] u_ca_out_45;
wire [71:0] u_ca_out_46;
wire [71:0] u_ca_out_47;
wire [71:0] u_ca_out_48;
wire [71:0] u_ca_out_49;
wire [71:0] u_ca_out_50;
wire [71:0] u_ca_out_51;
wire [71:0] u_ca_out_52;
wire [71:0] u_ca_out_53;
wire [71:0] u_ca_out_54;
wire [71:0] u_ca_out_55;
wire [71:0] u_ca_out_56;
wire [71:0] u_ca_out_57;
wire [71:0] u_ca_out_58;
wire [71:0] u_ca_out_59;
wire [71:0] u_ca_out_60;
wire [71:0] u_ca_out_61;
wire [71:0] u_ca_out_62;
wire [71:0] u_ca_out_63;
wire [71:0] u_ca_out_64;
wire [71:0] u_ca_out_65;
wire [71:0] u_ca_out_66;
wire [71:0] u_ca_out_67;
wire [71:0] u_ca_out_68;
wire [71:0] u_ca_out_69;
wire [71:0] u_ca_out_70;
wire [71:0] u_ca_out_71;
wire [71:0] u_ca_out_72;
wire [71:0] u_ca_out_73;
wire [71:0] u_ca_out_74;
wire [71:0] u_ca_out_75;
wire [71:0] u_ca_out_76;
wire [71:0] u_ca_out_77;
wire [71:0] u_ca_out_78;
wire [71:0] u_ca_out_79;
wire [71:0] u_ca_out_80;
wire [71:0] u_ca_out_81;
wire [71:0] u_ca_out_82;
wire [71:0] u_ca_out_83;
wire [71:0] u_ca_out_84;
wire [71:0] u_ca_out_85;
wire [71:0] u_ca_out_86;
wire [71:0] u_ca_out_87;
wire [71:0] u_ca_out_88;
wire [71:0] u_ca_out_89;
wire [71:0] u_ca_out_90;
wire [71:0] u_ca_out_91;
wire [71:0] u_ca_out_92;
wire [71:0] u_ca_out_93;
wire [71:0] u_ca_out_94;
wire [71:0] u_ca_out_95;
wire [71:0] u_ca_out_96;
wire [71:0] u_ca_out_97;
wire [71:0] u_ca_out_98;
wire [71:0] u_ca_out_99;
wire [71:0] u_ca_out_100;
wire [71:0] u_ca_out_101;
wire [71:0] u_ca_out_102;
wire [71:0] u_ca_out_103;
wire [71:0] u_ca_out_104;
wire [71:0] u_ca_out_105;
wire [71:0] u_ca_out_106;
wire [71:0] u_ca_out_107;
wire [71:0] u_ca_out_108;
wire [71:0] u_ca_out_109;
wire [71:0] u_ca_out_110;
wire [71:0] u_ca_out_111;
wire [71:0] u_ca_out_112;
wire [71:0] u_ca_out_113;
wire [71:0] u_ca_out_114;
wire [71:0] u_ca_out_115;
wire [71:0] u_ca_out_116;
wire [71:0] u_ca_out_117;
wire [71:0] u_ca_out_118;
wire [71:0] u_ca_out_119;
wire [71:0] u_ca_out_120;
wire [71:0] u_ca_out_121;
wire [71:0] u_ca_out_122;
wire [71:0] u_ca_out_123;
wire [71:0] u_ca_out_124;
wire [71:0] u_ca_out_125;
wire [71:0] u_ca_out_126;
wire [71:0] u_ca_out_127;
wire [71:0] u_ca_out_128;
wire [71:0] u_ca_out_129;
wire [71:0] u_ca_out_130;
wire [71:0] u_ca_out_131;
wire [71:0] u_ca_out_132;
wire [71:0] u_ca_out_133;
wire [71:0] u_ca_out_134;
wire [71:0] u_ca_out_135;
wire [71:0] u_ca_out_136;
wire [71:0] u_ca_out_137;
wire [71:0] u_ca_out_138;
wire [71:0] u_ca_out_139;
wire [71:0] u_ca_out_140;
wire [71:0] u_ca_out_141;
wire [71:0] u_ca_out_142;
wire [71:0] u_ca_out_143;
wire [71:0] u_ca_out_144;
wire [71:0] u_ca_out_145;
wire [71:0] u_ca_out_146;
wire [71:0] u_ca_out_147;
wire [71:0] u_ca_out_148;
wire [71:0] u_ca_out_149;
wire [71:0] u_ca_out_150;
wire [71:0] u_ca_out_151;
wire [71:0] u_ca_out_152;
wire [71:0] u_ca_out_153;
wire [71:0] u_ca_out_154;
wire [71:0] u_ca_out_155;
wire [71:0] u_ca_out_156;
wire [71:0] u_ca_out_157;
wire [71:0] u_ca_out_158;
wire [71:0] u_ca_out_159;
wire [71:0] u_ca_out_160;
wire [71:0] u_ca_out_161;
wire [71:0] u_ca_out_162;
wire [71:0] u_ca_out_163;
wire [71:0] u_ca_out_164;
wire [71:0] u_ca_out_165;
wire [71:0] u_ca_out_166;
wire [71:0] u_ca_out_167;
wire [71:0] u_ca_out_168;
wire [71:0] u_ca_out_169;
wire [71:0] u_ca_out_170;
wire [71:0] u_ca_out_171;
wire [71:0] u_ca_out_172;
wire [71:0] u_ca_out_173;
wire [71:0] u_ca_out_174;
wire [71:0] u_ca_out_175;
wire [71:0] u_ca_out_176;
wire [71:0] u_ca_out_177;
wire [71:0] u_ca_out_178;
wire [71:0] u_ca_out_179;
wire [71:0] u_ca_out_180;
wire [71:0] u_ca_out_181;
wire [71:0] u_ca_out_182;
wire [71:0] u_ca_out_183;
wire [71:0] u_ca_out_184;
wire [71:0] u_ca_out_185;
wire [71:0] u_ca_out_186;
wire [71:0] u_ca_out_187;
wire [71:0] u_ca_out_188;
wire [71:0] u_ca_out_189;
wire [71:0] u_ca_out_190;
wire [71:0] u_ca_out_191;
wire [71:0] u_ca_out_192;
wire [71:0] u_ca_out_193;
wire [71:0] u_ca_out_194;
wire [71:0] u_ca_out_195;
wire [71:0] u_ca_out_196;
wire [71:0] u_ca_out_197;
wire [71:0] u_ca_out_198;
wire [71:0] u_ca_out_199;
wire [71:0] u_ca_out_200;
wire [71:0] u_ca_out_201;
wire [71:0] u_ca_out_202;
wire [71:0] u_ca_out_203;
wire [71:0] u_ca_out_204;
wire [71:0] u_ca_out_205;
wire [71:0] u_ca_out_206;
wire [71:0] u_ca_out_207;
wire [71:0] u_ca_out_208;
wire [71:0] u_ca_out_209;
wire [71:0] u_ca_out_210;
wire [71:0] u_ca_out_211;
wire [71:0] u_ca_out_212;
wire [71:0] u_ca_out_213;
wire [71:0] u_ca_out_214;
wire [71:0] u_ca_out_215;
wire [71:0] u_ca_out_216;
wire [71:0] u_ca_out_217;
wire [71:0] u_ca_out_218;
wire [71:0] u_ca_out_219;
wire [71:0] u_ca_out_220;
wire [71:0] u_ca_out_221;
wire [71:0] u_ca_out_222;
wire [71:0] u_ca_out_223;
wire [71:0] u_ca_out_224;
wire [71:0] u_ca_out_225;
wire [71:0] u_ca_out_226;
wire [71:0] u_ca_out_227;
wire [71:0] u_ca_out_228;
wire [71:0] u_ca_out_229;
wire [71:0] u_ca_out_230;
wire [71:0] u_ca_out_231;
wire [71:0] u_ca_out_232;
wire [71:0] u_ca_out_233;
wire [71:0] u_ca_out_234;
wire [71:0] u_ca_out_235;
wire [71:0] u_ca_out_236;
wire [71:0] u_ca_out_237;
wire [71:0] u_ca_out_238;
wire [71:0] u_ca_out_239;
wire [71:0] u_ca_out_240;
wire [71:0] u_ca_out_241;
wire [71:0] u_ca_out_242;
wire [71:0] u_ca_out_243;
wire [71:0] u_ca_out_244;
wire [71:0] u_ca_out_245;
wire [71:0] u_ca_out_246;
wire [71:0] u_ca_out_247;
wire [71:0] u_ca_out_248;
wire [71:0] u_ca_out_249;
wire [71:0] u_ca_out_250;
wire [71:0] u_ca_out_251;
wire [71:0] u_ca_out_252;
wire [71:0] u_ca_out_253;
wire [71:0] u_ca_out_254;
wire [71:0] u_ca_out_255;
wire [71:0] u_ca_out_256;
wire [71:0] u_ca_out_257;
wire [71:0] u_ca_out_258;
wire [71:0] u_ca_out_259;
wire [71:0] u_ca_out_260;
wire [71:0] u_ca_out_261;
wire [71:0] u_ca_out_262;
wire [71:0] u_ca_out_263;
wire [71:0] u_ca_out_264;
wire [71:0] u_ca_out_265;
wire [71:0] u_ca_out_266;
wire [71:0] u_ca_out_267;
wire [71:0] u_ca_out_268;
wire [71:0] u_ca_out_269;
wire [71:0] u_ca_out_270;
wire [71:0] u_ca_out_271;
wire [71:0] u_ca_out_272;
wire [71:0] u_ca_out_273;
wire [71:0] u_ca_out_274;
wire [71:0] u_ca_out_275;
wire [71:0] u_ca_out_276;
wire [71:0] u_ca_out_277;
wire [71:0] u_ca_out_278;
wire [71:0] u_ca_out_279;
wire [71:0] u_ca_out_280;
wire [71:0] u_ca_out_281;
wire [71:0] u_ca_out_282;
wire [71:0] u_ca_out_283;
wire [71:0] u_ca_out_284;
wire [71:0] u_ca_out_285;
wire [71:0] u_ca_out_286;
wire [71:0] u_ca_out_287;
wire [71:0] u_ca_out_288;
wire [71:0] u_ca_out_289;
wire [71:0] u_ca_out_290;
wire [71:0] u_ca_out_291;
wire [71:0] u_ca_out_292;
wire [71:0] u_ca_out_293;
wire [71:0] u_ca_out_294;
wire [71:0] u_ca_out_295;
wire [71:0] u_ca_out_296;
wire [71:0] u_ca_out_297;
wire [71:0] u_ca_out_298;
wire [71:0] u_ca_out_299;
wire [71:0] u_ca_out_300;
wire [71:0] u_ca_out_301;
wire [71:0] u_ca_out_302;
wire [71:0] u_ca_out_303;
wire [71:0] u_ca_out_304;
wire [71:0] u_ca_out_305;
wire [71:0] u_ca_out_306;
wire [71:0] u_ca_out_307;
wire [71:0] u_ca_out_308;
wire [71:0] u_ca_out_309;
wire [71:0] u_ca_out_310;
wire [71:0] u_ca_out_311;
wire [71:0] u_ca_out_312;
wire [71:0] u_ca_out_313;
wire [71:0] u_ca_out_314;
wire [71:0] u_ca_out_315;
wire [71:0] u_ca_out_316;
wire [71:0] u_ca_out_317;
wire [71:0] u_ca_out_318;
wire [71:0] u_ca_out_319;
wire [71:0] u_ca_out_320;
wire [71:0] u_ca_out_321;
wire [71:0] u_ca_out_322;
wire [71:0] u_ca_out_323;
wire [71:0] u_ca_out_324;
wire [71:0] u_ca_out_325;
wire [71:0] u_ca_out_326;
wire [71:0] u_ca_out_327;
wire [71:0] u_ca_out_328;
wire [71:0] u_ca_out_329;
wire [71:0] u_ca_out_330;
wire [71:0] u_ca_out_331;
wire [71:0] u_ca_out_332;
wire [71:0] u_ca_out_333;
wire [71:0] u_ca_out_334;
wire [71:0] u_ca_out_335;
wire [71:0] u_ca_out_336;
wire [71:0] u_ca_out_337;
wire [71:0] u_ca_out_338;
wire [71:0] u_ca_out_339;
wire [71:0] u_ca_out_340;
wire [71:0] u_ca_out_341;
wire [71:0] u_ca_out_342;
wire [71:0] u_ca_out_343;
wire [71:0] u_ca_out_344;
wire [71:0] u_ca_out_345;
wire [71:0] u_ca_out_346;
wire [71:0] u_ca_out_347;
wire [71:0] u_ca_out_348;
wire [71:0] u_ca_out_349;
wire [71:0] u_ca_out_350;
wire [71:0] u_ca_out_351;
wire [71:0] u_ca_out_352;
wire [71:0] u_ca_out_353;
wire [71:0] u_ca_out_354;
wire [71:0] u_ca_out_355;
wire [71:0] u_ca_out_356;
wire [71:0] u_ca_out_357;
wire [71:0] u_ca_out_358;
wire [71:0] u_ca_out_359;
wire [71:0] u_ca_out_360;
wire [71:0] u_ca_out_361;
wire [71:0] u_ca_out_362;
wire [71:0] u_ca_out_363;
wire [71:0] u_ca_out_364;
wire [71:0] u_ca_out_365;
wire [71:0] u_ca_out_366;
wire [71:0] u_ca_out_367;
wire [71:0] u_ca_out_368;
wire [71:0] u_ca_out_369;
wire [71:0] u_ca_out_370;
wire [71:0] u_ca_out_371;
wire [71:0] u_ca_out_372;
wire [71:0] u_ca_out_373;
wire [71:0] u_ca_out_374;
wire [71:0] u_ca_out_375;
wire [71:0] u_ca_out_376;
wire [71:0] u_ca_out_377;
wire [71:0] u_ca_out_378;
wire [71:0] u_ca_out_379;
wire [71:0] u_ca_out_380;
wire [71:0] u_ca_out_381;
wire [71:0] u_ca_out_382;
wire [71:0] u_ca_out_383;
wire [71:0] u_ca_out_384;
wire [71:0] u_ca_out_385;
wire [71:0] u_ca_out_386;
wire [71:0] u_ca_out_387;
wire [71:0] u_ca_out_388;
wire [71:0] u_ca_out_389;
wire [71:0] u_ca_out_390;
wire [71:0] u_ca_out_391;
wire [71:0] u_ca_out_392;
wire [71:0] u_ca_out_393;
wire [71:0] u_ca_out_394;
wire [71:0] u_ca_out_395;
wire [71:0] u_ca_out_396;
wire [71:0] u_ca_out_397;
wire [71:0] u_ca_out_398;
wire [71:0] u_ca_out_399;
wire [71:0] u_ca_out_400;
wire [71:0] u_ca_out_401;
wire [71:0] u_ca_out_402;
wire [71:0] u_ca_out_403;
wire [71:0] u_ca_out_404;
wire [71:0] u_ca_out_405;
wire [71:0] u_ca_out_406;
wire [71:0] u_ca_out_407;
wire [71:0] u_ca_out_408;
wire [71:0] u_ca_out_409;
wire [71:0] u_ca_out_410;
wire [71:0] u_ca_out_411;
wire [71:0] u_ca_out_412;
wire [71:0] u_ca_out_413;
wire [71:0] u_ca_out_414;
wire [71:0] u_ca_out_415;
wire [71:0] u_ca_out_416;
wire [71:0] u_ca_out_417;
wire [71:0] u_ca_out_418;
wire [71:0] u_ca_out_419;
wire [71:0] u_ca_out_420;
wire [71:0] u_ca_out_421;
wire [71:0] u_ca_out_422;
wire [71:0] u_ca_out_423;
wire [71:0] u_ca_out_424;
wire [71:0] u_ca_out_425;
wire [71:0] u_ca_out_426;
wire [71:0] u_ca_out_427;
wire [71:0] u_ca_out_428;
wire [71:0] u_ca_out_429;
wire [71:0] u_ca_out_430;
wire [71:0] u_ca_out_431;
wire [71:0] u_ca_out_432;
wire [71:0] u_ca_out_433;
wire [71:0] u_ca_out_434;
wire [71:0] u_ca_out_435;
wire [71:0] u_ca_out_436;
wire [71:0] u_ca_out_437;
wire [71:0] u_ca_out_438;
wire [71:0] u_ca_out_439;
wire [71:0] u_ca_out_440;
wire [71:0] u_ca_out_441;
wire [71:0] u_ca_out_442;
wire [71:0] u_ca_out_443;
wire [71:0] u_ca_out_444;
wire [71:0] u_ca_out_445;
wire [71:0] u_ca_out_446;
wire [71:0] u_ca_out_447;
wire [71:0] u_ca_out_448;
wire [71:0] u_ca_out_449;
wire [71:0] u_ca_out_450;
wire [71:0] u_ca_out_451;
wire [71:0] u_ca_out_452;
wire [71:0] u_ca_out_453;
wire [71:0] u_ca_out_454;
wire [71:0] u_ca_out_455;
wire [71:0] u_ca_out_456;
wire [71:0] u_ca_out_457;
wire [71:0] u_ca_out_458;
wire [71:0] u_ca_out_459;
wire [71:0] u_ca_out_460;
wire [71:0] u_ca_out_461;
wire [71:0] u_ca_out_462;
wire [71:0] u_ca_out_463;
wire [71:0] u_ca_out_464;
wire [71:0] u_ca_out_465;
wire [71:0] u_ca_out_466;
wire [71:0] u_ca_out_467;
wire [71:0] u_ca_out_468;
wire [71:0] u_ca_out_469;
wire [71:0] u_ca_out_470;
wire [71:0] u_ca_out_471;
wire [71:0] u_ca_out_472;
wire [71:0] u_ca_out_473;
wire [71:0] u_ca_out_474;
wire [71:0] u_ca_out_475;
wire [71:0] u_ca_out_476;
wire [71:0] u_ca_out_477;
wire [71:0] u_ca_out_478;
wire [71:0] u_ca_out_479;
wire [71:0] u_ca_out_480;
wire [71:0] u_ca_out_481;
wire [71:0] u_ca_out_482;
wire [71:0] u_ca_out_483;
wire [71:0] u_ca_out_484;
wire [71:0] u_ca_out_485;
wire [71:0] u_ca_out_486;
wire [71:0] u_ca_out_487;
wire [71:0] u_ca_out_488;
wire [71:0] u_ca_out_489;
wire [71:0] u_ca_out_490;
wire [71:0] u_ca_out_491;
wire [71:0] u_ca_out_492;
wire [71:0] u_ca_out_493;
wire [71:0] u_ca_out_494;
wire [71:0] u_ca_out_495;
wire [71:0] u_ca_out_496;
wire [71:0] u_ca_out_497;
wire [71:0] u_ca_out_498;
wire [71:0] u_ca_out_499;
wire [71:0] u_ca_out_500;
wire [71:0] u_ca_out_501;
wire [71:0] u_ca_out_502;
wire [71:0] u_ca_out_503;
wire [71:0] u_ca_out_504;
wire [71:0] u_ca_out_505;
wire [71:0] u_ca_out_506;
wire [71:0] u_ca_out_507;
wire [71:0] u_ca_out_508;
wire [71:0] u_ca_out_509;
wire [71:0] u_ca_out_510;
wire [71:0] u_ca_out_511;
wire [71:0] u_ca_out_512;
wire [71:0] u_ca_out_513;
wire [71:0] u_ca_out_514;
wire [71:0] u_ca_out_515;
wire [71:0] u_ca_out_516;
wire [71:0] u_ca_out_517;
wire [71:0] u_ca_out_518;
wire [71:0] u_ca_out_519;
wire [71:0] u_ca_out_520;
wire [71:0] u_ca_out_521;
wire [71:0] u_ca_out_522;
wire [71:0] u_ca_out_523;
wire [71:0] u_ca_out_524;
wire [71:0] u_ca_out_525;
wire [71:0] u_ca_out_526;
wire [71:0] u_ca_out_527;
wire [71:0] u_ca_out_528;
wire [71:0] u_ca_out_529;
wire [71:0] u_ca_out_530;
wire [71:0] u_ca_out_531;
wire [71:0] u_ca_out_532;
wire [71:0] u_ca_out_533;
wire [71:0] u_ca_out_534;
wire [71:0] u_ca_out_535;
wire [71:0] u_ca_out_536;
wire [71:0] u_ca_out_537;
wire [71:0] u_ca_out_538;
wire [71:0] u_ca_out_539;
wire [71:0] u_ca_out_540;
wire [71:0] u_ca_out_541;
wire [71:0] u_ca_out_542;
wire [71:0] u_ca_out_543;
wire [71:0] u_ca_out_544;
wire [71:0] u_ca_out_545;
wire [71:0] u_ca_out_546;
wire [71:0] u_ca_out_547;
wire [71:0] u_ca_out_548;
wire [71:0] u_ca_out_549;
wire [71:0] u_ca_out_550;
wire [71:0] u_ca_out_551;
wire [71:0] u_ca_out_552;
wire [71:0] u_ca_out_553;
wire [71:0] u_ca_out_554;
wire [71:0] u_ca_out_555;
wire [71:0] u_ca_out_556;
wire [71:0] u_ca_out_557;
wire [71:0] u_ca_out_558;
wire [71:0] u_ca_out_559;
wire [71:0] u_ca_out_560;
wire [71:0] u_ca_out_561;
wire [71:0] u_ca_out_562;
wire [71:0] u_ca_out_563;
wire [71:0] u_ca_out_564;
wire [71:0] u_ca_out_565;
wire [71:0] u_ca_out_566;
wire [71:0] u_ca_out_567;
wire [71:0] u_ca_out_568;
wire [71:0] u_ca_out_569;
wire [71:0] u_ca_out_570;
wire [71:0] u_ca_out_571;
wire [71:0] u_ca_out_572;
wire [71:0] u_ca_out_573;
wire [71:0] u_ca_out_574;
wire [71:0] u_ca_out_575;
wire [71:0] u_ca_out_576;
wire [71:0] u_ca_out_577;
wire [71:0] u_ca_out_578;
wire [71:0] u_ca_out_579;
wire [71:0] u_ca_out_580;
wire [71:0] u_ca_out_581;
wire [71:0] u_ca_out_582;
wire [71:0] u_ca_out_583;
wire [71:0] u_ca_out_584;
wire [71:0] u_ca_out_585;
wire [71:0] u_ca_out_586;
wire [71:0] u_ca_out_587;
wire [71:0] u_ca_out_588;
wire [71:0] u_ca_out_589;
wire [71:0] u_ca_out_590;
wire [71:0] u_ca_out_591;
wire [71:0] u_ca_out_592;
wire [71:0] u_ca_out_593;
wire [71:0] u_ca_out_594;
wire [71:0] u_ca_out_595;
wire [71:0] u_ca_out_596;
wire [71:0] u_ca_out_597;
wire [71:0] u_ca_out_598;
wire [71:0] u_ca_out_599;
wire [71:0] u_ca_out_600;
wire [71:0] u_ca_out_601;
wire [71:0] u_ca_out_602;
wire [71:0] u_ca_out_603;
wire [71:0] u_ca_out_604;
wire [71:0] u_ca_out_605;
wire [71:0] u_ca_out_606;
wire [71:0] u_ca_out_607;
wire [71:0] u_ca_out_608;
wire [71:0] u_ca_out_609;
wire [71:0] u_ca_out_610;
wire [71:0] u_ca_out_611;
wire [71:0] u_ca_out_612;
wire [71:0] u_ca_out_613;
wire [71:0] u_ca_out_614;
wire [71:0] u_ca_out_615;
wire [71:0] u_ca_out_616;
wire [71:0] u_ca_out_617;
wire [71:0] u_ca_out_618;
wire [71:0] u_ca_out_619;
wire [71:0] u_ca_out_620;
wire [71:0] u_ca_out_621;
wire [71:0] u_ca_out_622;
wire [71:0] u_ca_out_623;
wire [71:0] u_ca_out_624;
wire [71:0] u_ca_out_625;
wire [71:0] u_ca_out_626;
wire [71:0] u_ca_out_627;
wire [71:0] u_ca_out_628;
wire [71:0] u_ca_out_629;
wire [71:0] u_ca_out_630;
wire [71:0] u_ca_out_631;
wire [71:0] u_ca_out_632;
wire [71:0] u_ca_out_633;
wire [71:0] u_ca_out_634;
wire [71:0] u_ca_out_635;
wire [71:0] u_ca_out_636;
wire [71:0] u_ca_out_637;
wire [71:0] u_ca_out_638;
wire [71:0] u_ca_out_639;
wire [71:0] u_ca_out_640;
wire [71:0] u_ca_out_641;
wire [71:0] u_ca_out_642;
wire [71:0] u_ca_out_643;
wire [71:0] u_ca_out_644;
wire [71:0] u_ca_out_645;
wire [71:0] u_ca_out_646;
wire [71:0] u_ca_out_647;
wire [71:0] u_ca_out_648;
wire [71:0] u_ca_out_649;
wire [71:0] u_ca_out_650;
wire [71:0] u_ca_out_651;
wire [71:0] u_ca_out_652;
wire [71:0] u_ca_out_653;
wire [71:0] u_ca_out_654;
wire [71:0] u_ca_out_655;
wire [71:0] u_ca_out_656;
wire [71:0] u_ca_out_657;
wire [71:0] u_ca_out_658;
wire [71:0] u_ca_out_659;
wire [71:0] u_ca_out_660;
wire [71:0] u_ca_out_661;
wire [71:0] u_ca_out_662;
wire [71:0] u_ca_out_663;
wire [71:0] u_ca_out_664;
wire [71:0] u_ca_out_665;
wire [71:0] u_ca_out_666;
wire [71:0] u_ca_out_667;
wire [71:0] u_ca_out_668;
wire [71:0] u_ca_out_669;
wire [71:0] u_ca_out_670;
wire [71:0] u_ca_out_671;
wire [71:0] u_ca_out_672;
wire [71:0] u_ca_out_673;
wire [71:0] u_ca_out_674;
wire [71:0] u_ca_out_675;
wire [71:0] u_ca_out_676;
wire [71:0] u_ca_out_677;
wire [71:0] u_ca_out_678;
wire [71:0] u_ca_out_679;
wire [71:0] u_ca_out_680;
wire [71:0] u_ca_out_681;
wire [71:0] u_ca_out_682;
wire [71:0] u_ca_out_683;
wire [71:0] u_ca_out_684;
wire [71:0] u_ca_out_685;
wire [71:0] u_ca_out_686;
wire [71:0] u_ca_out_687;
wire [71:0] u_ca_out_688;
wire [71:0] u_ca_out_689;
wire [71:0] u_ca_out_690;
wire [71:0] u_ca_out_691;
wire [71:0] u_ca_out_692;
wire [71:0] u_ca_out_693;
wire [71:0] u_ca_out_694;
wire [71:0] u_ca_out_695;
wire [71:0] u_ca_out_696;
wire [71:0] u_ca_out_697;
wire [71:0] u_ca_out_698;
wire [71:0] u_ca_out_699;
wire [71:0] u_ca_out_700;
wire [71:0] u_ca_out_701;
wire [71:0] u_ca_out_702;
wire [71:0] u_ca_out_703;
wire [71:0] u_ca_out_704;
wire [71:0] u_ca_out_705;
wire [71:0] u_ca_out_706;
wire [71:0] u_ca_out_707;
wire [71:0] u_ca_out_708;
wire [71:0] u_ca_out_709;
wire [71:0] u_ca_out_710;
wire [71:0] u_ca_out_711;
wire [71:0] u_ca_out_712;
wire [71:0] u_ca_out_713;
wire [71:0] u_ca_out_714;
wire [71:0] u_ca_out_715;
wire [71:0] u_ca_out_716;
wire [71:0] u_ca_out_717;
wire [71:0] u_ca_out_718;
wire [71:0] u_ca_out_719;
wire [71:0] u_ca_out_720;
wire [71:0] u_ca_out_721;
wire [71:0] u_ca_out_722;
wire [71:0] u_ca_out_723;
wire [71:0] u_ca_out_724;
wire [71:0] u_ca_out_725;
wire [71:0] u_ca_out_726;
wire [71:0] u_ca_out_727;
wire [71:0] u_ca_out_728;
wire [71:0] u_ca_out_729;
wire [71:0] u_ca_out_730;
wire [71:0] u_ca_out_731;
wire [71:0] u_ca_out_732;
wire [71:0] u_ca_out_733;
wire [71:0] u_ca_out_734;
wire [71:0] u_ca_out_735;
wire [71:0] u_ca_out_736;
wire [71:0] u_ca_out_737;
wire [71:0] u_ca_out_738;
wire [71:0] u_ca_out_739;
wire [71:0] u_ca_out_740;
wire [71:0] u_ca_out_741;
wire [71:0] u_ca_out_742;
wire [71:0] u_ca_out_743;
wire [71:0] u_ca_out_744;
wire [71:0] u_ca_out_745;
wire [71:0] u_ca_out_746;
wire [71:0] u_ca_out_747;
wire [71:0] u_ca_out_748;
wire [71:0] u_ca_out_749;
wire [71:0] u_ca_out_750;
wire [71:0] u_ca_out_751;
wire [71:0] u_ca_out_752;
wire [71:0] u_ca_out_753;
wire [71:0] u_ca_out_754;
wire [71:0] u_ca_out_755;
wire [71:0] u_ca_out_756;
wire [71:0] u_ca_out_757;
wire [71:0] u_ca_out_758;
wire [71:0] u_ca_out_759;
wire [71:0] u_ca_out_760;
wire [71:0] u_ca_out_761;
wire [71:0] u_ca_out_762;
wire [71:0] u_ca_out_763;
wire [71:0] u_ca_out_764;
wire [71:0] u_ca_out_765;
wire [71:0] u_ca_out_766;
wire [71:0] u_ca_out_767;
wire [71:0] u_ca_out_768;
wire [71:0] u_ca_out_769;
wire [71:0] u_ca_out_770;
wire [71:0] u_ca_out_771;
wire [71:0] u_ca_out_772;
wire [71:0] u_ca_out_773;
wire [71:0] u_ca_out_774;
wire [71:0] u_ca_out_775;
wire [71:0] u_ca_out_776;
wire [71:0] u_ca_out_777;
wire [71:0] u_ca_out_778;
wire [71:0] u_ca_out_779;
wire [71:0] u_ca_out_780;
wire [71:0] u_ca_out_781;
wire [71:0] u_ca_out_782;
wire [71:0] u_ca_out_783;
wire [71:0] u_ca_out_784;
wire [71:0] u_ca_out_785;
wire [71:0] u_ca_out_786;
wire [71:0] u_ca_out_787;
wire [71:0] u_ca_out_788;
wire [71:0] u_ca_out_789;
wire [71:0] u_ca_out_790;
wire [71:0] u_ca_out_791;
wire [71:0] u_ca_out_792;
wire [71:0] u_ca_out_793;
wire [71:0] u_ca_out_794;
wire [71:0] u_ca_out_795;
wire [71:0] u_ca_out_796;
wire [71:0] u_ca_out_797;
wire [71:0] u_ca_out_798;
wire [71:0] u_ca_out_799;
wire [71:0] u_ca_out_800;
wire [71:0] u_ca_out_801;
wire [71:0] u_ca_out_802;
wire [71:0] u_ca_out_803;
wire [71:0] u_ca_out_804;
wire [71:0] u_ca_out_805;
wire [71:0] u_ca_out_806;
wire [71:0] u_ca_out_807;
wire [71:0] u_ca_out_808;
wire [71:0] u_ca_out_809;
wire [71:0] u_ca_out_810;
wire [71:0] u_ca_out_811;
wire [71:0] u_ca_out_812;
wire [71:0] u_ca_out_813;
wire [71:0] u_ca_out_814;
wire [71:0] u_ca_out_815;
wire [71:0] u_ca_out_816;
wire [71:0] u_ca_out_817;
wire [71:0] u_ca_out_818;
wire [71:0] u_ca_out_819;
wire [71:0] u_ca_out_820;
wire [71:0] u_ca_out_821;
wire [71:0] u_ca_out_822;
wire [71:0] u_ca_out_823;
wire [71:0] u_ca_out_824;
wire [71:0] u_ca_out_825;
wire [71:0] u_ca_out_826;
wire [71:0] u_ca_out_827;
wire [71:0] u_ca_out_828;
wire [71:0] u_ca_out_829;
wire [71:0] u_ca_out_830;
wire [71:0] u_ca_out_831;
wire [71:0] u_ca_out_832;
wire [71:0] u_ca_out_833;
wire [71:0] u_ca_out_834;
wire [71:0] u_ca_out_835;
wire [71:0] u_ca_out_836;
wire [71:0] u_ca_out_837;
wire [71:0] u_ca_out_838;
wire [71:0] u_ca_out_839;
wire [71:0] u_ca_out_840;
wire [71:0] u_ca_out_841;
wire [71:0] u_ca_out_842;
wire [71:0] u_ca_out_843;
wire [71:0] u_ca_out_844;
wire [71:0] u_ca_out_845;
wire [71:0] u_ca_out_846;
wire [71:0] u_ca_out_847;
wire [71:0] u_ca_out_848;
wire [71:0] u_ca_out_849;
wire [71:0] u_ca_out_850;
wire [71:0] u_ca_out_851;
wire [71:0] u_ca_out_852;
wire [71:0] u_ca_out_853;
wire [71:0] u_ca_out_854;
wire [71:0] u_ca_out_855;
wire [71:0] u_ca_out_856;
wire [71:0] u_ca_out_857;
wire [71:0] u_ca_out_858;
wire [71:0] u_ca_out_859;
wire [71:0] u_ca_out_860;
wire [71:0] u_ca_out_861;
wire [71:0] u_ca_out_862;
wire [71:0] u_ca_out_863;
wire [71:0] u_ca_out_864;
wire [71:0] u_ca_out_865;
wire [71:0] u_ca_out_866;
wire [71:0] u_ca_out_867;
wire [71:0] u_ca_out_868;
wire [71:0] u_ca_out_869;
wire [71:0] u_ca_out_870;
wire [71:0] u_ca_out_871;
wire [71:0] u_ca_out_872;
wire [71:0] u_ca_out_873;
wire [71:0] u_ca_out_874;
wire [71:0] u_ca_out_875;
wire [71:0] u_ca_out_876;
wire [71:0] u_ca_out_877;
wire [71:0] u_ca_out_878;
wire [71:0] u_ca_out_879;
wire [71:0] u_ca_out_880;
wire [71:0] u_ca_out_881;
wire [71:0] u_ca_out_882;
wire [71:0] u_ca_out_883;
wire [71:0] u_ca_out_884;
wire [71:0] u_ca_out_885;
wire [71:0] u_ca_out_886;
wire [71:0] u_ca_out_887;
wire [71:0] u_ca_out_888;
wire [71:0] u_ca_out_889;
wire [71:0] u_ca_out_890;
wire [71:0] u_ca_out_891;
wire [71:0] u_ca_out_892;
wire [71:0] u_ca_out_893;
wire [71:0] u_ca_out_894;
wire [71:0] u_ca_out_895;
wire [71:0] u_ca_out_896;
wire [71:0] u_ca_out_897;
wire [71:0] u_ca_out_898;
wire [71:0] u_ca_out_899;
wire [71:0] u_ca_out_900;
wire [71:0] u_ca_out_901;
wire [71:0] u_ca_out_902;
wire [71:0] u_ca_out_903;
wire [71:0] u_ca_out_904;
wire [71:0] u_ca_out_905;
wire [71:0] u_ca_out_906;
wire [71:0] u_ca_out_907;
wire [71:0] u_ca_out_908;
wire [71:0] u_ca_out_909;
wire [71:0] u_ca_out_910;
wire [71:0] u_ca_out_911;
wire [71:0] u_ca_out_912;
wire [71:0] u_ca_out_913;
wire [71:0] u_ca_out_914;
wire [71:0] u_ca_out_915;
wire [71:0] u_ca_out_916;
wire [71:0] u_ca_out_917;
wire [71:0] u_ca_out_918;
wire [71:0] u_ca_out_919;
wire [71:0] u_ca_out_920;
wire [71:0] u_ca_out_921;
wire [71:0] u_ca_out_922;
wire [71:0] u_ca_out_923;
wire [71:0] u_ca_out_924;
wire [71:0] u_ca_out_925;
wire [71:0] u_ca_out_926;
wire [71:0] u_ca_out_927;
wire [71:0] u_ca_out_928;
wire [71:0] u_ca_out_929;
wire [71:0] u_ca_out_930;
wire [71:0] u_ca_out_931;
wire [71:0] u_ca_out_932;
wire [71:0] u_ca_out_933;
wire [71:0] u_ca_out_934;
wire [71:0] u_ca_out_935;
wire [71:0] u_ca_out_936;
wire [71:0] u_ca_out_937;
wire [71:0] u_ca_out_938;
wire [71:0] u_ca_out_939;
wire [71:0] u_ca_out_940;
wire [71:0] u_ca_out_941;
wire [71:0] u_ca_out_942;
wire [71:0] u_ca_out_943;
wire [71:0] u_ca_out_944;
wire [71:0] u_ca_out_945;
wire [71:0] u_ca_out_946;
wire [71:0] u_ca_out_947;
wire [71:0] u_ca_out_948;
wire [71:0] u_ca_out_949;
wire [71:0] u_ca_out_950;
wire [71:0] u_ca_out_951;
wire [71:0] u_ca_out_952;
wire [71:0] u_ca_out_953;
wire [71:0] u_ca_out_954;
wire [71:0] u_ca_out_955;
wire [71:0] u_ca_out_956;
wire [71:0] u_ca_out_957;
wire [71:0] u_ca_out_958;
wire [71:0] u_ca_out_959;
wire [71:0] u_ca_out_960;
wire [71:0] u_ca_out_961;
wire [71:0] u_ca_out_962;
wire [71:0] u_ca_out_963;
wire [71:0] u_ca_out_964;
wire [71:0] u_ca_out_965;
wire [71:0] u_ca_out_966;
wire [71:0] u_ca_out_967;
wire [71:0] u_ca_out_968;
wire [71:0] u_ca_out_969;
wire [71:0] u_ca_out_970;
wire [71:0] u_ca_out_971;
wire [71:0] u_ca_out_972;
wire [71:0] u_ca_out_973;
wire [71:0] u_ca_out_974;
wire [71:0] u_ca_out_975;
wire [71:0] u_ca_out_976;
wire [71:0] u_ca_out_977;
wire [71:0] u_ca_out_978;
wire [71:0] u_ca_out_979;
wire [71:0] u_ca_out_980;
wire [71:0] u_ca_out_981;
wire [71:0] u_ca_out_982;
wire [71:0] u_ca_out_983;
wire [71:0] u_ca_out_984;
wire [71:0] u_ca_out_985;
wire [71:0] u_ca_out_986;
wire [71:0] u_ca_out_987;
wire [71:0] u_ca_out_988;
wire [71:0] u_ca_out_989;
wire [71:0] u_ca_out_990;
wire [71:0] u_ca_out_991;
wire [71:0] u_ca_out_992;
wire [71:0] u_ca_out_993;
wire [71:0] u_ca_out_994;
wire [71:0] u_ca_out_995;
wire [71:0] u_ca_out_996;
wire [71:0] u_ca_out_997;
wire [71:0] u_ca_out_998;
wire [71:0] u_ca_out_999;
wire [71:0] u_ca_out_1000;
wire [71:0] u_ca_out_1001;
wire [71:0] u_ca_out_1002;
wire [71:0] u_ca_out_1003;
wire [71:0] u_ca_out_1004;
wire [71:0] u_ca_out_1005;
wire [71:0] u_ca_out_1006;
wire [71:0] u_ca_out_1007;
wire [71:0] u_ca_out_1008;
wire [71:0] u_ca_out_1009;
wire [71:0] u_ca_out_1010;
wire [71:0] u_ca_out_1011;
wire [71:0] u_ca_out_1012;
wire [71:0] u_ca_out_1013;
wire [71:0] u_ca_out_1014;
wire [71:0] u_ca_out_1015;
wire [71:0] u_ca_out_1016;
wire [71:0] u_ca_out_1017;
wire [71:0] u_ca_out_1018;
wire [71:0] u_ca_out_1019;
wire [71:0] u_ca_out_1020;
wire [71:0] u_ca_out_1021;
wire [71:0] u_ca_out_1022;
wire [71:0] u_ca_out_1023;
wire [71:0] u_ca_out_1024;
wire [71:0] u_ca_out_1025;
wire [71:0] u_ca_out_1026;
wire [71:0] u_ca_out_1027;
wire [71:0] u_ca_out_1028;
wire [71:0] u_ca_out_1029;
wire [71:0] u_ca_out_1030;
wire [71:0] u_ca_out_1031;
wire [71:0] u_ca_out_1032;
wire [71:0] u_ca_out_1033;
wire [71:0] u_ca_out_1034;
wire [71:0] u_ca_out_1035;
wire [71:0] u_ca_out_1036;
wire [71:0] u_ca_out_1037;
wire [71:0] u_ca_out_1038;
wire [71:0] u_ca_out_1039;
wire [71:0] u_ca_out_1040;
wire [71:0] u_ca_out_1041;
wire [71:0] u_ca_out_1042;
wire [71:0] u_ca_out_1043;
wire [71:0] u_ca_out_1044;
wire [71:0] u_ca_out_1045;
wire [71:0] u_ca_out_1046;
wire [71:0] u_ca_out_1047;
wire [71:0] u_ca_out_1048;
wire [71:0] u_ca_out_1049;
wire [71:0] u_ca_out_1050;
wire [71:0] u_ca_out_1051;
wire [71:0] u_ca_out_1052;
wire [71:0] u_ca_out_1053;
wire [71:0] u_ca_out_1054;
wire [71:0] u_ca_out_1055;
wire [71:0] u_ca_out_1056;
wire [71:0] u_ca_out_1057;
wire [71:0] u_ca_out_1058;
wire [71:0] u_ca_out_1059;
wire [71:0] u_ca_out_1060;
wire [71:0] u_ca_out_1061;
wire [71:0] u_ca_out_1062;
wire [71:0] u_ca_out_1063;
wire [71:0] u_ca_out_1064;
wire [71:0] u_ca_out_1065;
wire [71:0] u_ca_out_1066;
wire [71:0] u_ca_out_1067;
wire [71:0] u_ca_out_1068;
wire [71:0] u_ca_out_1069;
wire [71:0] u_ca_out_1070;
wire [71:0] u_ca_out_1071;
wire [71:0] u_ca_out_1072;
wire [71:0] u_ca_out_1073;
wire [71:0] u_ca_out_1074;
wire [71:0] u_ca_out_1075;
wire [71:0] u_ca_out_1076;
wire [71:0] u_ca_out_1077;
wire [71:0] u_ca_out_1078;
wire [71:0] u_ca_out_1079;
wire [71:0] u_ca_out_1080;
wire [71:0] u_ca_out_1081;
wire [71:0] u_ca_out_1082;
wire [71:0] u_ca_out_1083;
wire [71:0] u_ca_out_1084;
wire [71:0] u_ca_out_1085;
wire [71:0] u_ca_out_1086;
wire [71:0] u_ca_out_1087;
wire [71:0] u_ca_out_1088;
wire [71:0] u_ca_out_1089;
wire [71:0] u_ca_out_1090;
wire [71:0] u_ca_out_1091;
wire [71:0] u_ca_out_1092;
wire [71:0] u_ca_out_1093;
wire [71:0] u_ca_out_1094;
wire [71:0] u_ca_out_1095;
wire [71:0] u_ca_out_1096;
wire [71:0] u_ca_out_1097;
wire [71:0] u_ca_out_1098;
wire [71:0] u_ca_out_1099;
wire [71:0] u_ca_out_1100;
wire [71:0] u_ca_out_1101;
wire [71:0] u_ca_out_1102;
wire [71:0] u_ca_out_1103;
wire [71:0] u_ca_out_1104;
wire [71:0] u_ca_out_1105;
wire [71:0] u_ca_out_1106;
wire [71:0] u_ca_out_1107;
wire [71:0] u_ca_out_1108;
wire [71:0] u_ca_out_1109;
wire [71:0] u_ca_out_1110;
wire [71:0] u_ca_out_1111;
wire [71:0] u_ca_out_1112;
wire [71:0] u_ca_out_1113;
wire [71:0] u_ca_out_1114;
wire [71:0] u_ca_out_1115;
wire [71:0] u_ca_out_1116;
wire [71:0] u_ca_out_1117;
wire [71:0] u_ca_out_1118;
wire [71:0] u_ca_out_1119;
wire [71:0] u_ca_out_1120;
wire [71:0] u_ca_out_1121;
wire [71:0] u_ca_out_1122;
wire [71:0] u_ca_out_1123;
wire [71:0] u_ca_out_1124;
wire [71:0] u_ca_out_1125;
wire [71:0] u_ca_out_1126;
wire [71:0] u_ca_out_1127;
wire [71:0] u_ca_out_1128;
wire [71:0] u_ca_out_1129;
wire [71:0] u_ca_out_1130;
wire [71:0] u_ca_out_1131;
wire [71:0] u_ca_out_1132;
wire [71:0] u_ca_out_1133;
wire [71:0] u_ca_out_1134;
wire [71:0] u_ca_out_1135;
wire [71:0] u_ca_out_1136;
wire [71:0] u_ca_out_1137;
wire [71:0] u_ca_out_1138;
wire [71:0] u_ca_out_1139;
wire [71:0] u_ca_out_1140;
wire [71:0] u_ca_out_1141;
wire [71:0] u_ca_out_1142;
wire [71:0] u_ca_out_1143;
wire [71:0] u_ca_out_1144;
wire [71:0] u_ca_out_1145;
wire [71:0] u_ca_out_1146;
wire [71:0] u_ca_out_1147;
wire [71:0] u_ca_out_1148;
wire [71:0] u_ca_out_1149;
wire [71:0] u_ca_out_1150;
wire [71:0] u_ca_out_1151;
wire [71:0] u_ca_out_1152;
wire [71:0] u_ca_out_1153;
wire [71:0] u_ca_out_1154;
wire [71:0] u_ca_out_1155;
wire [71:0] u_ca_out_1156;
wire [71:0] u_ca_out_1157;
wire [71:0] u_ca_out_1158;
wire [71:0] u_ca_out_1159;
wire [71:0] u_ca_out_1160;
wire [71:0] u_ca_out_1161;
wire [71:0] u_ca_out_1162;
wire [71:0] u_ca_out_1163;
wire [71:0] u_ca_out_1164;
wire [71:0] u_ca_out_1165;
wire [71:0] u_ca_out_1166;
wire [71:0] u_ca_out_1167;
wire [71:0] u_ca_out_1168;
wire [71:0] u_ca_out_1169;
wire [71:0] u_ca_out_1170;
wire [71:0] u_ca_out_1171;
wire [71:0] u_ca_out_1172;
wire [71:0] u_ca_out_1173;
wire [71:0] u_ca_out_1174;
wire [71:0] u_ca_out_1175;
wire [71:0] u_ca_out_1176;
wire [71:0] u_ca_out_1177;
wire [71:0] u_ca_out_1178;
wire [71:0] u_ca_out_1179;
wire [71:0] u_ca_out_1180;
wire [71:0] u_ca_out_1181;
wire [71:0] u_ca_out_1182;
wire [71:0] u_ca_out_1183;
wire [71:0] u_ca_out_1184;
wire [71:0] u_ca_out_1185;
wire [71:0] u_ca_out_1186;
wire [71:0] u_ca_out_1187;
wire [71:0] u_ca_out_1188;
wire [71:0] u_ca_out_1189;
wire [71:0] u_ca_out_1190;
wire [71:0] u_ca_out_1191;
wire [71:0] u_ca_out_1192;
wire [71:0] u_ca_out_1193;
wire [71:0] u_ca_out_1194;
wire [71:0] u_ca_out_1195;
wire [71:0] u_ca_out_1196;
wire [71:0] u_ca_out_1197;
wire [71:0] u_ca_out_1198;
wire [71:0] u_ca_out_1199;
wire [71:0] u_ca_out_1200;
wire [71:0] u_ca_out_1201;
wire [71:0] u_ca_out_1202;
wire [71:0] u_ca_out_1203;
wire [71:0] u_ca_out_1204;
wire [71:0] u_ca_out_1205;
wire [71:0] u_ca_out_1206;
wire [71:0] u_ca_out_1207;
wire [71:0] u_ca_out_1208;
wire [71:0] u_ca_out_1209;
wire [71:0] u_ca_out_1210;
wire [71:0] u_ca_out_1211;
wire [71:0] u_ca_out_1212;
wire [71:0] u_ca_out_1213;
wire [71:0] u_ca_out_1214;
wire [71:0] u_ca_out_1215;
wire [71:0] u_ca_out_1216;
wire [71:0] u_ca_out_1217;
wire [71:0] u_ca_out_1218;
wire [71:0] u_ca_out_1219;
wire [71:0] u_ca_out_1220;
wire [71:0] u_ca_out_1221;
wire [71:0] u_ca_out_1222;
wire [71:0] u_ca_out_1223;
wire [71:0] u_ca_out_1224;
wire [71:0] u_ca_out_1225;
wire [71:0] u_ca_out_1226;
wire [71:0] u_ca_out_1227;
wire [71:0] u_ca_out_1228;
wire [71:0] u_ca_out_1229;
wire [71:0] u_ca_out_1230;
wire [71:0] u_ca_out_1231;
wire [71:0] u_ca_out_1232;
wire [71:0] u_ca_out_1233;
wire [71:0] u_ca_out_1234;
wire [71:0] u_ca_out_1235;
wire [71:0] u_ca_out_1236;
wire [71:0] u_ca_out_1237;
wire [71:0] u_ca_out_1238;
wire [71:0] u_ca_out_1239;
wire [71:0] u_ca_out_1240;
wire [71:0] u_ca_out_1241;
wire [71:0] u_ca_out_1242;
wire [71:0] u_ca_out_1243;
wire [71:0] u_ca_out_1244;
wire [71:0] u_ca_out_1245;
wire [71:0] u_ca_out_1246;
wire [71:0] u_ca_out_1247;
wire [71:0] u_ca_out_1248;
wire [71:0] u_ca_out_1249;
wire [71:0] u_ca_out_1250;
wire [71:0] u_ca_out_1251;
wire [71:0] u_ca_out_1252;
wire [71:0] u_ca_out_1253;
wire [71:0] u_ca_out_1254;
wire [71:0] u_ca_out_1255;
wire [71:0] u_ca_out_1256;
wire [71:0] u_ca_out_1257;
wire [71:0] u_ca_out_1258;
wire [71:0] u_ca_out_1259;
wire [71:0] u_ca_out_1260;
wire [71:0] u_ca_out_1261;
wire [71:0] u_ca_out_1262;
wire [71:0] u_ca_out_1263;
wire [71:0] u_ca_out_1264;
wire [71:0] u_ca_out_1265;
wire [71:0] u_ca_out_1266;
wire [71:0] u_ca_out_1267;
wire [71:0] u_ca_out_1268;
wire [71:0] u_ca_out_1269;
wire [71:0] u_ca_out_1270;
wire [71:0] u_ca_out_1271;
wire [71:0] u_ca_out_1272;
wire [71:0] u_ca_out_1273;
wire [71:0] u_ca_out_1274;
wire [71:0] u_ca_out_1275;
wire [71:0] u_ca_out_1276;
wire [71:0] u_ca_out_1277;
wire [71:0] u_ca_out_1278;
wire [71:0] u_ca_out_1279;

assign u_ca_in_0 = {{7{1'b0}}, col_in_0};
assign u_ca_in_1 = {{7{1'b0}}, col_in_1};
assign u_ca_in_2 = {{7{1'b0}}, col_in_2};
assign u_ca_in_3 = {{7{1'b0}}, col_in_3};
assign u_ca_in_4 = {{7{1'b0}}, col_in_4};
assign u_ca_in_5 = {{7{1'b0}}, col_in_5};
assign u_ca_in_6 = {{7{1'b0}}, col_in_6};
assign u_ca_in_7 = {{7{1'b0}}, col_in_7};
assign u_ca_in_8 = {{7{1'b0}}, col_in_8};
assign u_ca_in_9 = {{7{1'b0}}, col_in_9};
assign u_ca_in_10 = {{7{1'b0}}, col_in_10};
assign u_ca_in_11 = {{7{1'b0}}, col_in_11};
assign u_ca_in_12 = {{7{1'b0}}, col_in_12};
assign u_ca_in_13 = {{7{1'b0}}, col_in_13};
assign u_ca_in_14 = {{7{1'b0}}, col_in_14};
assign u_ca_in_15 = {{7{1'b0}}, col_in_15};
assign u_ca_in_16 = {{7{1'b0}}, col_in_16};
assign u_ca_in_17 = {{7{1'b0}}, col_in_17};
assign u_ca_in_18 = {{7{1'b0}}, col_in_18};
assign u_ca_in_19 = {{7{1'b0}}, col_in_19};
assign u_ca_in_20 = {{7{1'b0}}, col_in_20};
assign u_ca_in_21 = {{7{1'b0}}, col_in_21};
assign u_ca_in_22 = {{7{1'b0}}, col_in_22};
assign u_ca_in_23 = {{7{1'b0}}, col_in_23};
assign u_ca_in_24 = {{7{1'b0}}, col_in_24};
assign u_ca_in_25 = {{7{1'b0}}, col_in_25};
assign u_ca_in_26 = {{7{1'b0}}, col_in_26};
assign u_ca_in_27 = {{7{1'b0}}, col_in_27};
assign u_ca_in_28 = {{7{1'b0}}, col_in_28};
assign u_ca_in_29 = {{7{1'b0}}, col_in_29};
assign u_ca_in_30 = {{7{1'b0}}, col_in_30};
assign u_ca_in_31 = {{7{1'b0}}, col_in_31};
assign u_ca_in_32 = {{7{1'b0}}, col_in_32};
assign u_ca_in_33 = {{7{1'b0}}, col_in_33};
assign u_ca_in_34 = {{7{1'b0}}, col_in_34};
assign u_ca_in_35 = {{7{1'b0}}, col_in_35};
assign u_ca_in_36 = {{7{1'b0}}, col_in_36};
assign u_ca_in_37 = {{7{1'b0}}, col_in_37};
assign u_ca_in_38 = {{7{1'b0}}, col_in_38};
assign u_ca_in_39 = {{7{1'b0}}, col_in_39};
assign u_ca_in_40 = {{7{1'b0}}, col_in_40};
assign u_ca_in_41 = {{7{1'b0}}, col_in_41};
assign u_ca_in_42 = {{7{1'b0}}, col_in_42};
assign u_ca_in_43 = {{7{1'b0}}, col_in_43};
assign u_ca_in_44 = {{7{1'b0}}, col_in_44};
assign u_ca_in_45 = {{7{1'b0}}, col_in_45};
assign u_ca_in_46 = {{7{1'b0}}, col_in_46};
assign u_ca_in_47 = {{7{1'b0}}, col_in_47};
assign u_ca_in_48 = {{7{1'b0}}, col_in_48};
assign u_ca_in_49 = {{7{1'b0}}, col_in_49};
assign u_ca_in_50 = {{7{1'b0}}, col_in_50};
assign u_ca_in_51 = {{7{1'b0}}, col_in_51};
assign u_ca_in_52 = {{7{1'b0}}, col_in_52};
assign u_ca_in_53 = {{7{1'b0}}, col_in_53};
assign u_ca_in_54 = {{7{1'b0}}, col_in_54};
assign u_ca_in_55 = {{7{1'b0}}, col_in_55};
assign u_ca_in_56 = {{7{1'b0}}, col_in_56};
assign u_ca_in_57 = {{7{1'b0}}, col_in_57};
assign u_ca_in_58 = {{7{1'b0}}, col_in_58};
assign u_ca_in_59 = {{7{1'b0}}, col_in_59};
assign u_ca_in_60 = {{7{1'b0}}, col_in_60};
assign u_ca_in_61 = {{7{1'b0}}, col_in_61};
assign u_ca_in_62 = {{7{1'b0}}, col_in_62};
assign u_ca_in_63 = {{7{1'b0}}, col_in_63};
assign u_ca_in_64 = {{7{1'b0}}, col_in_64};
assign u_ca_in_65 = {{7{1'b0}}, col_in_65};
assign u_ca_in_66 = {{7{1'b0}}, col_in_66};
assign u_ca_in_67 = {{7{1'b0}}, col_in_67};
assign u_ca_in_68 = {{7{1'b0}}, col_in_68};
assign u_ca_in_69 = {{7{1'b0}}, col_in_69};
assign u_ca_in_70 = {{7{1'b0}}, col_in_70};
assign u_ca_in_71 = {{7{1'b0}}, col_in_71};
assign u_ca_in_72 = {{7{1'b0}}, col_in_72};
assign u_ca_in_73 = {{7{1'b0}}, col_in_73};
assign u_ca_in_74 = {{7{1'b0}}, col_in_74};
assign u_ca_in_75 = {{7{1'b0}}, col_in_75};
assign u_ca_in_76 = {{7{1'b0}}, col_in_76};
assign u_ca_in_77 = {{7{1'b0}}, col_in_77};
assign u_ca_in_78 = {{7{1'b0}}, col_in_78};
assign u_ca_in_79 = {{7{1'b0}}, col_in_79};
assign u_ca_in_80 = {{7{1'b0}}, col_in_80};
assign u_ca_in_81 = {{7{1'b0}}, col_in_81};
assign u_ca_in_82 = {{7{1'b0}}, col_in_82};
assign u_ca_in_83 = {{7{1'b0}}, col_in_83};
assign u_ca_in_84 = {{7{1'b0}}, col_in_84};
assign u_ca_in_85 = {{7{1'b0}}, col_in_85};
assign u_ca_in_86 = {{7{1'b0}}, col_in_86};
assign u_ca_in_87 = {{7{1'b0}}, col_in_87};
assign u_ca_in_88 = {{7{1'b0}}, col_in_88};
assign u_ca_in_89 = {{7{1'b0}}, col_in_89};
assign u_ca_in_90 = {{7{1'b0}}, col_in_90};
assign u_ca_in_91 = {{7{1'b0}}, col_in_91};
assign u_ca_in_92 = {{7{1'b0}}, col_in_92};
assign u_ca_in_93 = {{7{1'b0}}, col_in_93};
assign u_ca_in_94 = {{7{1'b0}}, col_in_94};
assign u_ca_in_95 = {{7{1'b0}}, col_in_95};
assign u_ca_in_96 = {{7{1'b0}}, col_in_96};
assign u_ca_in_97 = {{7{1'b0}}, col_in_97};
assign u_ca_in_98 = {{7{1'b0}}, col_in_98};
assign u_ca_in_99 = {{7{1'b0}}, col_in_99};
assign u_ca_in_100 = {{7{1'b0}}, col_in_100};
assign u_ca_in_101 = {{7{1'b0}}, col_in_101};
assign u_ca_in_102 = {{7{1'b0}}, col_in_102};
assign u_ca_in_103 = {{7{1'b0}}, col_in_103};
assign u_ca_in_104 = {{7{1'b0}}, col_in_104};
assign u_ca_in_105 = {{7{1'b0}}, col_in_105};
assign u_ca_in_106 = {{7{1'b0}}, col_in_106};
assign u_ca_in_107 = {{7{1'b0}}, col_in_107};
assign u_ca_in_108 = {{7{1'b0}}, col_in_108};
assign u_ca_in_109 = {{7{1'b0}}, col_in_109};
assign u_ca_in_110 = {{7{1'b0}}, col_in_110};
assign u_ca_in_111 = {{7{1'b0}}, col_in_111};
assign u_ca_in_112 = {{7{1'b0}}, col_in_112};
assign u_ca_in_113 = {{7{1'b0}}, col_in_113};
assign u_ca_in_114 = {{7{1'b0}}, col_in_114};
assign u_ca_in_115 = {{7{1'b0}}, col_in_115};
assign u_ca_in_116 = {{7{1'b0}}, col_in_116};
assign u_ca_in_117 = {{7{1'b0}}, col_in_117};
assign u_ca_in_118 = {{7{1'b0}}, col_in_118};
assign u_ca_in_119 = {{7{1'b0}}, col_in_119};
assign u_ca_in_120 = {{7{1'b0}}, col_in_120};
assign u_ca_in_121 = {{7{1'b0}}, col_in_121};
assign u_ca_in_122 = {{7{1'b0}}, col_in_122};
assign u_ca_in_123 = {{7{1'b0}}, col_in_123};
assign u_ca_in_124 = {{7{1'b0}}, col_in_124};
assign u_ca_in_125 = {{7{1'b0}}, col_in_125};
assign u_ca_in_126 = {{7{1'b0}}, col_in_126};
assign u_ca_in_127 = {{7{1'b0}}, col_in_127};
assign u_ca_in_128 = {{7{1'b0}}, col_in_128};
assign u_ca_in_129 = {{7{1'b0}}, col_in_129};
assign u_ca_in_130 = {{7{1'b0}}, col_in_130};
assign u_ca_in_131 = {{7{1'b0}}, col_in_131};
assign u_ca_in_132 = {{7{1'b0}}, col_in_132};
assign u_ca_in_133 = {{7{1'b0}}, col_in_133};
assign u_ca_in_134 = {{7{1'b0}}, col_in_134};
assign u_ca_in_135 = {{7{1'b0}}, col_in_135};
assign u_ca_in_136 = {{7{1'b0}}, col_in_136};
assign u_ca_in_137 = {{7{1'b0}}, col_in_137};
assign u_ca_in_138 = {{7{1'b0}}, col_in_138};
assign u_ca_in_139 = {{7{1'b0}}, col_in_139};
assign u_ca_in_140 = {{7{1'b0}}, col_in_140};
assign u_ca_in_141 = {{7{1'b0}}, col_in_141};
assign u_ca_in_142 = {{7{1'b0}}, col_in_142};
assign u_ca_in_143 = {{7{1'b0}}, col_in_143};
assign u_ca_in_144 = {{7{1'b0}}, col_in_144};
assign u_ca_in_145 = {{7{1'b0}}, col_in_145};
assign u_ca_in_146 = {{7{1'b0}}, col_in_146};
assign u_ca_in_147 = {{7{1'b0}}, col_in_147};
assign u_ca_in_148 = {{7{1'b0}}, col_in_148};
assign u_ca_in_149 = {{7{1'b0}}, col_in_149};
assign u_ca_in_150 = {{7{1'b0}}, col_in_150};
assign u_ca_in_151 = {{7{1'b0}}, col_in_151};
assign u_ca_in_152 = {{7{1'b0}}, col_in_152};
assign u_ca_in_153 = {{7{1'b0}}, col_in_153};
assign u_ca_in_154 = {{7{1'b0}}, col_in_154};
assign u_ca_in_155 = {{7{1'b0}}, col_in_155};
assign u_ca_in_156 = {{7{1'b0}}, col_in_156};
assign u_ca_in_157 = {{7{1'b0}}, col_in_157};
assign u_ca_in_158 = {{7{1'b0}}, col_in_158};
assign u_ca_in_159 = {{7{1'b0}}, col_in_159};
assign u_ca_in_160 = {{7{1'b0}}, col_in_160};
assign u_ca_in_161 = {{7{1'b0}}, col_in_161};
assign u_ca_in_162 = {{7{1'b0}}, col_in_162};
assign u_ca_in_163 = {{7{1'b0}}, col_in_163};
assign u_ca_in_164 = {{7{1'b0}}, col_in_164};
assign u_ca_in_165 = {{7{1'b0}}, col_in_165};
assign u_ca_in_166 = {{7{1'b0}}, col_in_166};
assign u_ca_in_167 = {{7{1'b0}}, col_in_167};
assign u_ca_in_168 = {{7{1'b0}}, col_in_168};
assign u_ca_in_169 = {{7{1'b0}}, col_in_169};
assign u_ca_in_170 = {{7{1'b0}}, col_in_170};
assign u_ca_in_171 = {{7{1'b0}}, col_in_171};
assign u_ca_in_172 = {{7{1'b0}}, col_in_172};
assign u_ca_in_173 = {{7{1'b0}}, col_in_173};
assign u_ca_in_174 = {{7{1'b0}}, col_in_174};
assign u_ca_in_175 = {{7{1'b0}}, col_in_175};
assign u_ca_in_176 = {{7{1'b0}}, col_in_176};
assign u_ca_in_177 = {{7{1'b0}}, col_in_177};
assign u_ca_in_178 = {{7{1'b0}}, col_in_178};
assign u_ca_in_179 = {{7{1'b0}}, col_in_179};
assign u_ca_in_180 = {{7{1'b0}}, col_in_180};
assign u_ca_in_181 = {{7{1'b0}}, col_in_181};
assign u_ca_in_182 = {{7{1'b0}}, col_in_182};
assign u_ca_in_183 = {{7{1'b0}}, col_in_183};
assign u_ca_in_184 = {{7{1'b0}}, col_in_184};
assign u_ca_in_185 = {{7{1'b0}}, col_in_185};
assign u_ca_in_186 = {{7{1'b0}}, col_in_186};
assign u_ca_in_187 = {{7{1'b0}}, col_in_187};
assign u_ca_in_188 = {{7{1'b0}}, col_in_188};
assign u_ca_in_189 = {{7{1'b0}}, col_in_189};
assign u_ca_in_190 = {{7{1'b0}}, col_in_190};
assign u_ca_in_191 = {{7{1'b0}}, col_in_191};
assign u_ca_in_192 = {{7{1'b0}}, col_in_192};
assign u_ca_in_193 = {{7{1'b0}}, col_in_193};
assign u_ca_in_194 = {{7{1'b0}}, col_in_194};
assign u_ca_in_195 = {{7{1'b0}}, col_in_195};
assign u_ca_in_196 = {{7{1'b0}}, col_in_196};
assign u_ca_in_197 = {{7{1'b0}}, col_in_197};
assign u_ca_in_198 = {{7{1'b0}}, col_in_198};
assign u_ca_in_199 = {{7{1'b0}}, col_in_199};
assign u_ca_in_200 = {{7{1'b0}}, col_in_200};
assign u_ca_in_201 = {{7{1'b0}}, col_in_201};
assign u_ca_in_202 = {{7{1'b0}}, col_in_202};
assign u_ca_in_203 = {{7{1'b0}}, col_in_203};
assign u_ca_in_204 = {{7{1'b0}}, col_in_204};
assign u_ca_in_205 = {{7{1'b0}}, col_in_205};
assign u_ca_in_206 = {{7{1'b0}}, col_in_206};
assign u_ca_in_207 = {{7{1'b0}}, col_in_207};
assign u_ca_in_208 = {{7{1'b0}}, col_in_208};
assign u_ca_in_209 = {{7{1'b0}}, col_in_209};
assign u_ca_in_210 = {{7{1'b0}}, col_in_210};
assign u_ca_in_211 = {{7{1'b0}}, col_in_211};
assign u_ca_in_212 = {{7{1'b0}}, col_in_212};
assign u_ca_in_213 = {{7{1'b0}}, col_in_213};
assign u_ca_in_214 = {{7{1'b0}}, col_in_214};
assign u_ca_in_215 = {{7{1'b0}}, col_in_215};
assign u_ca_in_216 = {{7{1'b0}}, col_in_216};
assign u_ca_in_217 = {{7{1'b0}}, col_in_217};
assign u_ca_in_218 = {{7{1'b0}}, col_in_218};
assign u_ca_in_219 = {{7{1'b0}}, col_in_219};
assign u_ca_in_220 = {{7{1'b0}}, col_in_220};
assign u_ca_in_221 = {{7{1'b0}}, col_in_221};
assign u_ca_in_222 = {{7{1'b0}}, col_in_222};
assign u_ca_in_223 = {{7{1'b0}}, col_in_223};
assign u_ca_in_224 = {{7{1'b0}}, col_in_224};
assign u_ca_in_225 = {{7{1'b0}}, col_in_225};
assign u_ca_in_226 = {{7{1'b0}}, col_in_226};
assign u_ca_in_227 = {{7{1'b0}}, col_in_227};
assign u_ca_in_228 = {{7{1'b0}}, col_in_228};
assign u_ca_in_229 = {{7{1'b0}}, col_in_229};
assign u_ca_in_230 = {{7{1'b0}}, col_in_230};
assign u_ca_in_231 = {{7{1'b0}}, col_in_231};
assign u_ca_in_232 = {{7{1'b0}}, col_in_232};
assign u_ca_in_233 = {{7{1'b0}}, col_in_233};
assign u_ca_in_234 = {{7{1'b0}}, col_in_234};
assign u_ca_in_235 = {{7{1'b0}}, col_in_235};
assign u_ca_in_236 = {{7{1'b0}}, col_in_236};
assign u_ca_in_237 = {{7{1'b0}}, col_in_237};
assign u_ca_in_238 = {{7{1'b0}}, col_in_238};
assign u_ca_in_239 = {{7{1'b0}}, col_in_239};
assign u_ca_in_240 = {{7{1'b0}}, col_in_240};
assign u_ca_in_241 = {{7{1'b0}}, col_in_241};
assign u_ca_in_242 = {{7{1'b0}}, col_in_242};
assign u_ca_in_243 = {{7{1'b0}}, col_in_243};
assign u_ca_in_244 = {{7{1'b0}}, col_in_244};
assign u_ca_in_245 = {{7{1'b0}}, col_in_245};
assign u_ca_in_246 = {{7{1'b0}}, col_in_246};
assign u_ca_in_247 = {{7{1'b0}}, col_in_247};
assign u_ca_in_248 = {{7{1'b0}}, col_in_248};
assign u_ca_in_249 = {{7{1'b0}}, col_in_249};
assign u_ca_in_250 = {{7{1'b0}}, col_in_250};
assign u_ca_in_251 = {{7{1'b0}}, col_in_251};
assign u_ca_in_252 = {{7{1'b0}}, col_in_252};
assign u_ca_in_253 = {{7{1'b0}}, col_in_253};
assign u_ca_in_254 = {{7{1'b0}}, col_in_254};
assign u_ca_in_255 = {{7{1'b0}}, col_in_255};
assign u_ca_in_256 = {{7{1'b0}}, col_in_256};
assign u_ca_in_257 = {{7{1'b0}}, col_in_257};
assign u_ca_in_258 = {{7{1'b0}}, col_in_258};
assign u_ca_in_259 = {{7{1'b0}}, col_in_259};
assign u_ca_in_260 = {{7{1'b0}}, col_in_260};
assign u_ca_in_261 = {{7{1'b0}}, col_in_261};
assign u_ca_in_262 = {{7{1'b0}}, col_in_262};
assign u_ca_in_263 = {{7{1'b0}}, col_in_263};
assign u_ca_in_264 = {{7{1'b0}}, col_in_264};
assign u_ca_in_265 = {{7{1'b0}}, col_in_265};
assign u_ca_in_266 = {{7{1'b0}}, col_in_266};
assign u_ca_in_267 = {{7{1'b0}}, col_in_267};
assign u_ca_in_268 = {{7{1'b0}}, col_in_268};
assign u_ca_in_269 = {{7{1'b0}}, col_in_269};
assign u_ca_in_270 = {{7{1'b0}}, col_in_270};
assign u_ca_in_271 = {{7{1'b0}}, col_in_271};
assign u_ca_in_272 = {{7{1'b0}}, col_in_272};
assign u_ca_in_273 = {{7{1'b0}}, col_in_273};
assign u_ca_in_274 = {{7{1'b0}}, col_in_274};
assign u_ca_in_275 = {{7{1'b0}}, col_in_275};
assign u_ca_in_276 = {{7{1'b0}}, col_in_276};
assign u_ca_in_277 = {{7{1'b0}}, col_in_277};
assign u_ca_in_278 = {{7{1'b0}}, col_in_278};
assign u_ca_in_279 = {{7{1'b0}}, col_in_279};
assign u_ca_in_280 = {{7{1'b0}}, col_in_280};
assign u_ca_in_281 = {{7{1'b0}}, col_in_281};
assign u_ca_in_282 = {{7{1'b0}}, col_in_282};
assign u_ca_in_283 = {{7{1'b0}}, col_in_283};
assign u_ca_in_284 = {{7{1'b0}}, col_in_284};
assign u_ca_in_285 = {{7{1'b0}}, col_in_285};
assign u_ca_in_286 = {{7{1'b0}}, col_in_286};
assign u_ca_in_287 = {{7{1'b0}}, col_in_287};
assign u_ca_in_288 = {{7{1'b0}}, col_in_288};
assign u_ca_in_289 = {{7{1'b0}}, col_in_289};
assign u_ca_in_290 = {{7{1'b0}}, col_in_290};
assign u_ca_in_291 = {{7{1'b0}}, col_in_291};
assign u_ca_in_292 = {{7{1'b0}}, col_in_292};
assign u_ca_in_293 = {{7{1'b0}}, col_in_293};
assign u_ca_in_294 = {{7{1'b0}}, col_in_294};
assign u_ca_in_295 = {{7{1'b0}}, col_in_295};
assign u_ca_in_296 = {{7{1'b0}}, col_in_296};
assign u_ca_in_297 = {{7{1'b0}}, col_in_297};
assign u_ca_in_298 = {{7{1'b0}}, col_in_298};
assign u_ca_in_299 = {{7{1'b0}}, col_in_299};
assign u_ca_in_300 = {{7{1'b0}}, col_in_300};
assign u_ca_in_301 = {{7{1'b0}}, col_in_301};
assign u_ca_in_302 = {{7{1'b0}}, col_in_302};
assign u_ca_in_303 = {{7{1'b0}}, col_in_303};
assign u_ca_in_304 = {{7{1'b0}}, col_in_304};
assign u_ca_in_305 = {{7{1'b0}}, col_in_305};
assign u_ca_in_306 = {{7{1'b0}}, col_in_306};
assign u_ca_in_307 = {{7{1'b0}}, col_in_307};
assign u_ca_in_308 = {{7{1'b0}}, col_in_308};
assign u_ca_in_309 = {{7{1'b0}}, col_in_309};
assign u_ca_in_310 = {{7{1'b0}}, col_in_310};
assign u_ca_in_311 = {{7{1'b0}}, col_in_311};
assign u_ca_in_312 = {{7{1'b0}}, col_in_312};
assign u_ca_in_313 = {{7{1'b0}}, col_in_313};
assign u_ca_in_314 = {{7{1'b0}}, col_in_314};
assign u_ca_in_315 = {{7{1'b0}}, col_in_315};
assign u_ca_in_316 = {{7{1'b0}}, col_in_316};
assign u_ca_in_317 = {{7{1'b0}}, col_in_317};
assign u_ca_in_318 = {{7{1'b0}}, col_in_318};
assign u_ca_in_319 = {{7{1'b0}}, col_in_319};
assign u_ca_in_320 = {{7{1'b0}}, col_in_320};
assign u_ca_in_321 = {{7{1'b0}}, col_in_321};
assign u_ca_in_322 = {{7{1'b0}}, col_in_322};
assign u_ca_in_323 = {{7{1'b0}}, col_in_323};
assign u_ca_in_324 = {{7{1'b0}}, col_in_324};
assign u_ca_in_325 = {{7{1'b0}}, col_in_325};
assign u_ca_in_326 = {{7{1'b0}}, col_in_326};
assign u_ca_in_327 = {{7{1'b0}}, col_in_327};
assign u_ca_in_328 = {{7{1'b0}}, col_in_328};
assign u_ca_in_329 = {{7{1'b0}}, col_in_329};
assign u_ca_in_330 = {{7{1'b0}}, col_in_330};
assign u_ca_in_331 = {{7{1'b0}}, col_in_331};
assign u_ca_in_332 = {{7{1'b0}}, col_in_332};
assign u_ca_in_333 = {{7{1'b0}}, col_in_333};
assign u_ca_in_334 = {{7{1'b0}}, col_in_334};
assign u_ca_in_335 = {{7{1'b0}}, col_in_335};
assign u_ca_in_336 = {{7{1'b0}}, col_in_336};
assign u_ca_in_337 = {{7{1'b0}}, col_in_337};
assign u_ca_in_338 = {{7{1'b0}}, col_in_338};
assign u_ca_in_339 = {{7{1'b0}}, col_in_339};
assign u_ca_in_340 = {{7{1'b0}}, col_in_340};
assign u_ca_in_341 = {{7{1'b0}}, col_in_341};
assign u_ca_in_342 = {{7{1'b0}}, col_in_342};
assign u_ca_in_343 = {{7{1'b0}}, col_in_343};
assign u_ca_in_344 = {{7{1'b0}}, col_in_344};
assign u_ca_in_345 = {{7{1'b0}}, col_in_345};
assign u_ca_in_346 = {{7{1'b0}}, col_in_346};
assign u_ca_in_347 = {{7{1'b0}}, col_in_347};
assign u_ca_in_348 = {{7{1'b0}}, col_in_348};
assign u_ca_in_349 = {{7{1'b0}}, col_in_349};
assign u_ca_in_350 = {{7{1'b0}}, col_in_350};
assign u_ca_in_351 = {{7{1'b0}}, col_in_351};
assign u_ca_in_352 = {{7{1'b0}}, col_in_352};
assign u_ca_in_353 = {{7{1'b0}}, col_in_353};
assign u_ca_in_354 = {{7{1'b0}}, col_in_354};
assign u_ca_in_355 = {{7{1'b0}}, col_in_355};
assign u_ca_in_356 = {{7{1'b0}}, col_in_356};
assign u_ca_in_357 = {{7{1'b0}}, col_in_357};
assign u_ca_in_358 = {{7{1'b0}}, col_in_358};
assign u_ca_in_359 = {{7{1'b0}}, col_in_359};
assign u_ca_in_360 = {{7{1'b0}}, col_in_360};
assign u_ca_in_361 = {{7{1'b0}}, col_in_361};
assign u_ca_in_362 = {{7{1'b0}}, col_in_362};
assign u_ca_in_363 = {{7{1'b0}}, col_in_363};
assign u_ca_in_364 = {{7{1'b0}}, col_in_364};
assign u_ca_in_365 = {{7{1'b0}}, col_in_365};
assign u_ca_in_366 = {{7{1'b0}}, col_in_366};
assign u_ca_in_367 = {{7{1'b0}}, col_in_367};
assign u_ca_in_368 = {{7{1'b0}}, col_in_368};
assign u_ca_in_369 = {{7{1'b0}}, col_in_369};
assign u_ca_in_370 = {{7{1'b0}}, col_in_370};
assign u_ca_in_371 = {{7{1'b0}}, col_in_371};
assign u_ca_in_372 = {{7{1'b0}}, col_in_372};
assign u_ca_in_373 = {{7{1'b0}}, col_in_373};
assign u_ca_in_374 = {{7{1'b0}}, col_in_374};
assign u_ca_in_375 = {{7{1'b0}}, col_in_375};
assign u_ca_in_376 = {{7{1'b0}}, col_in_376};
assign u_ca_in_377 = {{7{1'b0}}, col_in_377};
assign u_ca_in_378 = {{7{1'b0}}, col_in_378};
assign u_ca_in_379 = {{7{1'b0}}, col_in_379};
assign u_ca_in_380 = {{7{1'b0}}, col_in_380};
assign u_ca_in_381 = {{7{1'b0}}, col_in_381};
assign u_ca_in_382 = {{7{1'b0}}, col_in_382};
assign u_ca_in_383 = {{7{1'b0}}, col_in_383};
assign u_ca_in_384 = {{7{1'b0}}, col_in_384};
assign u_ca_in_385 = {{7{1'b0}}, col_in_385};
assign u_ca_in_386 = {{7{1'b0}}, col_in_386};
assign u_ca_in_387 = {{7{1'b0}}, col_in_387};
assign u_ca_in_388 = {{7{1'b0}}, col_in_388};
assign u_ca_in_389 = {{7{1'b0}}, col_in_389};
assign u_ca_in_390 = {{7{1'b0}}, col_in_390};
assign u_ca_in_391 = {{7{1'b0}}, col_in_391};
assign u_ca_in_392 = {{7{1'b0}}, col_in_392};
assign u_ca_in_393 = {{7{1'b0}}, col_in_393};
assign u_ca_in_394 = {{7{1'b0}}, col_in_394};
assign u_ca_in_395 = {{7{1'b0}}, col_in_395};
assign u_ca_in_396 = {{7{1'b0}}, col_in_396};
assign u_ca_in_397 = {{7{1'b0}}, col_in_397};
assign u_ca_in_398 = {{7{1'b0}}, col_in_398};
assign u_ca_in_399 = {{7{1'b0}}, col_in_399};
assign u_ca_in_400 = {{7{1'b0}}, col_in_400};
assign u_ca_in_401 = {{7{1'b0}}, col_in_401};
assign u_ca_in_402 = {{7{1'b0}}, col_in_402};
assign u_ca_in_403 = {{7{1'b0}}, col_in_403};
assign u_ca_in_404 = {{7{1'b0}}, col_in_404};
assign u_ca_in_405 = {{7{1'b0}}, col_in_405};
assign u_ca_in_406 = {{7{1'b0}}, col_in_406};
assign u_ca_in_407 = {{7{1'b0}}, col_in_407};
assign u_ca_in_408 = {{7{1'b0}}, col_in_408};
assign u_ca_in_409 = {{7{1'b0}}, col_in_409};
assign u_ca_in_410 = {{7{1'b0}}, col_in_410};
assign u_ca_in_411 = {{7{1'b0}}, col_in_411};
assign u_ca_in_412 = {{7{1'b0}}, col_in_412};
assign u_ca_in_413 = {{7{1'b0}}, col_in_413};
assign u_ca_in_414 = {{7{1'b0}}, col_in_414};
assign u_ca_in_415 = {{7{1'b0}}, col_in_415};
assign u_ca_in_416 = {{7{1'b0}}, col_in_416};
assign u_ca_in_417 = {{7{1'b0}}, col_in_417};
assign u_ca_in_418 = {{7{1'b0}}, col_in_418};
assign u_ca_in_419 = {{7{1'b0}}, col_in_419};
assign u_ca_in_420 = {{7{1'b0}}, col_in_420};
assign u_ca_in_421 = {{7{1'b0}}, col_in_421};
assign u_ca_in_422 = {{7{1'b0}}, col_in_422};
assign u_ca_in_423 = {{7{1'b0}}, col_in_423};
assign u_ca_in_424 = {{7{1'b0}}, col_in_424};
assign u_ca_in_425 = {{7{1'b0}}, col_in_425};
assign u_ca_in_426 = {{7{1'b0}}, col_in_426};
assign u_ca_in_427 = {{7{1'b0}}, col_in_427};
assign u_ca_in_428 = {{7{1'b0}}, col_in_428};
assign u_ca_in_429 = {{7{1'b0}}, col_in_429};
assign u_ca_in_430 = {{7{1'b0}}, col_in_430};
assign u_ca_in_431 = {{7{1'b0}}, col_in_431};
assign u_ca_in_432 = {{7{1'b0}}, col_in_432};
assign u_ca_in_433 = {{7{1'b0}}, col_in_433};
assign u_ca_in_434 = {{7{1'b0}}, col_in_434};
assign u_ca_in_435 = {{7{1'b0}}, col_in_435};
assign u_ca_in_436 = {{7{1'b0}}, col_in_436};
assign u_ca_in_437 = {{7{1'b0}}, col_in_437};
assign u_ca_in_438 = {{7{1'b0}}, col_in_438};
assign u_ca_in_439 = {{7{1'b0}}, col_in_439};
assign u_ca_in_440 = {{7{1'b0}}, col_in_440};
assign u_ca_in_441 = {{7{1'b0}}, col_in_441};
assign u_ca_in_442 = {{7{1'b0}}, col_in_442};
assign u_ca_in_443 = {{7{1'b0}}, col_in_443};
assign u_ca_in_444 = {{7{1'b0}}, col_in_444};
assign u_ca_in_445 = {{7{1'b0}}, col_in_445};
assign u_ca_in_446 = {{7{1'b0}}, col_in_446};
assign u_ca_in_447 = {{7{1'b0}}, col_in_447};
assign u_ca_in_448 = {{7{1'b0}}, col_in_448};
assign u_ca_in_449 = {{7{1'b0}}, col_in_449};
assign u_ca_in_450 = {{7{1'b0}}, col_in_450};
assign u_ca_in_451 = {{7{1'b0}}, col_in_451};
assign u_ca_in_452 = {{7{1'b0}}, col_in_452};
assign u_ca_in_453 = {{7{1'b0}}, col_in_453};
assign u_ca_in_454 = {{7{1'b0}}, col_in_454};
assign u_ca_in_455 = {{7{1'b0}}, col_in_455};
assign u_ca_in_456 = {{7{1'b0}}, col_in_456};
assign u_ca_in_457 = {{7{1'b0}}, col_in_457};
assign u_ca_in_458 = {{7{1'b0}}, col_in_458};
assign u_ca_in_459 = {{7{1'b0}}, col_in_459};
assign u_ca_in_460 = {{7{1'b0}}, col_in_460};
assign u_ca_in_461 = {{7{1'b0}}, col_in_461};
assign u_ca_in_462 = {{7{1'b0}}, col_in_462};
assign u_ca_in_463 = {{7{1'b0}}, col_in_463};
assign u_ca_in_464 = {{7{1'b0}}, col_in_464};
assign u_ca_in_465 = {{7{1'b0}}, col_in_465};
assign u_ca_in_466 = {{7{1'b0}}, col_in_466};
assign u_ca_in_467 = {{7{1'b0}}, col_in_467};
assign u_ca_in_468 = {{7{1'b0}}, col_in_468};
assign u_ca_in_469 = {{7{1'b0}}, col_in_469};
assign u_ca_in_470 = {{7{1'b0}}, col_in_470};
assign u_ca_in_471 = {{7{1'b0}}, col_in_471};
assign u_ca_in_472 = {{7{1'b0}}, col_in_472};
assign u_ca_in_473 = {{7{1'b0}}, col_in_473};
assign u_ca_in_474 = {{7{1'b0}}, col_in_474};
assign u_ca_in_475 = {{7{1'b0}}, col_in_475};
assign u_ca_in_476 = {{7{1'b0}}, col_in_476};
assign u_ca_in_477 = {{7{1'b0}}, col_in_477};
assign u_ca_in_478 = {{7{1'b0}}, col_in_478};
assign u_ca_in_479 = {{7{1'b0}}, col_in_479};
assign u_ca_in_480 = {{7{1'b0}}, col_in_480};
assign u_ca_in_481 = {{7{1'b0}}, col_in_481};
assign u_ca_in_482 = {{7{1'b0}}, col_in_482};
assign u_ca_in_483 = {{7{1'b0}}, col_in_483};
assign u_ca_in_484 = {{7{1'b0}}, col_in_484};
assign u_ca_in_485 = {{7{1'b0}}, col_in_485};
assign u_ca_in_486 = {{7{1'b0}}, col_in_486};
assign u_ca_in_487 = {{7{1'b0}}, col_in_487};
assign u_ca_in_488 = {{7{1'b0}}, col_in_488};
assign u_ca_in_489 = {{7{1'b0}}, col_in_489};
assign u_ca_in_490 = {{7{1'b0}}, col_in_490};
assign u_ca_in_491 = {{7{1'b0}}, col_in_491};
assign u_ca_in_492 = {{7{1'b0}}, col_in_492};
assign u_ca_in_493 = {{7{1'b0}}, col_in_493};
assign u_ca_in_494 = {{7{1'b0}}, col_in_494};
assign u_ca_in_495 = {{7{1'b0}}, col_in_495};
assign u_ca_in_496 = {{7{1'b0}}, col_in_496};
assign u_ca_in_497 = {{7{1'b0}}, col_in_497};
assign u_ca_in_498 = {{7{1'b0}}, col_in_498};
assign u_ca_in_499 = {{7{1'b0}}, col_in_499};
assign u_ca_in_500 = {{7{1'b0}}, col_in_500};
assign u_ca_in_501 = {{7{1'b0}}, col_in_501};
assign u_ca_in_502 = {{7{1'b0}}, col_in_502};
assign u_ca_in_503 = {{7{1'b0}}, col_in_503};
assign u_ca_in_504 = {{7{1'b0}}, col_in_504};
assign u_ca_in_505 = {{7{1'b0}}, col_in_505};
assign u_ca_in_506 = {{7{1'b0}}, col_in_506};
assign u_ca_in_507 = {{7{1'b0}}, col_in_507};
assign u_ca_in_508 = {{7{1'b0}}, col_in_508};
assign u_ca_in_509 = {{7{1'b0}}, col_in_509};
assign u_ca_in_510 = {{7{1'b0}}, col_in_510};
assign u_ca_in_511 = {{7{1'b0}}, col_in_511};
assign u_ca_in_512 = {{7{1'b0}}, col_in_512};
assign u_ca_in_513 = {{7{1'b0}}, col_in_513};
assign u_ca_in_514 = {{7{1'b0}}, col_in_514};
assign u_ca_in_515 = {{7{1'b0}}, col_in_515};
assign u_ca_in_516 = {{7{1'b0}}, col_in_516};
assign u_ca_in_517 = {{7{1'b0}}, col_in_517};
assign u_ca_in_518 = {{7{1'b0}}, col_in_518};
assign u_ca_in_519 = {{7{1'b0}}, col_in_519};
assign u_ca_in_520 = {{7{1'b0}}, col_in_520};
assign u_ca_in_521 = {{7{1'b0}}, col_in_521};
assign u_ca_in_522 = {{7{1'b0}}, col_in_522};
assign u_ca_in_523 = {{7{1'b0}}, col_in_523};
assign u_ca_in_524 = {{7{1'b0}}, col_in_524};
assign u_ca_in_525 = {{7{1'b0}}, col_in_525};
assign u_ca_in_526 = {{7{1'b0}}, col_in_526};
assign u_ca_in_527 = {{7{1'b0}}, col_in_527};
assign u_ca_in_528 = {{7{1'b0}}, col_in_528};
assign u_ca_in_529 = {{7{1'b0}}, col_in_529};
assign u_ca_in_530 = {{7{1'b0}}, col_in_530};
assign u_ca_in_531 = {{7{1'b0}}, col_in_531};
assign u_ca_in_532 = {{7{1'b0}}, col_in_532};
assign u_ca_in_533 = {{7{1'b0}}, col_in_533};
assign u_ca_in_534 = {{7{1'b0}}, col_in_534};
assign u_ca_in_535 = {{7{1'b0}}, col_in_535};
assign u_ca_in_536 = {{7{1'b0}}, col_in_536};
assign u_ca_in_537 = {{7{1'b0}}, col_in_537};
assign u_ca_in_538 = {{7{1'b0}}, col_in_538};
assign u_ca_in_539 = {{7{1'b0}}, col_in_539};
assign u_ca_in_540 = {{7{1'b0}}, col_in_540};
assign u_ca_in_541 = {{7{1'b0}}, col_in_541};
assign u_ca_in_542 = {{7{1'b0}}, col_in_542};
assign u_ca_in_543 = {{7{1'b0}}, col_in_543};
assign u_ca_in_544 = {{7{1'b0}}, col_in_544};
assign u_ca_in_545 = {{7{1'b0}}, col_in_545};
assign u_ca_in_546 = {{7{1'b0}}, col_in_546};
assign u_ca_in_547 = {{7{1'b0}}, col_in_547};
assign u_ca_in_548 = {{7{1'b0}}, col_in_548};
assign u_ca_in_549 = {{7{1'b0}}, col_in_549};
assign u_ca_in_550 = {{7{1'b0}}, col_in_550};
assign u_ca_in_551 = {{7{1'b0}}, col_in_551};
assign u_ca_in_552 = {{7{1'b0}}, col_in_552};
assign u_ca_in_553 = {{7{1'b0}}, col_in_553};
assign u_ca_in_554 = {{7{1'b0}}, col_in_554};
assign u_ca_in_555 = {{7{1'b0}}, col_in_555};
assign u_ca_in_556 = {{7{1'b0}}, col_in_556};
assign u_ca_in_557 = {{7{1'b0}}, col_in_557};
assign u_ca_in_558 = {{7{1'b0}}, col_in_558};
assign u_ca_in_559 = {{7{1'b0}}, col_in_559};
assign u_ca_in_560 = {{7{1'b0}}, col_in_560};
assign u_ca_in_561 = {{7{1'b0}}, col_in_561};
assign u_ca_in_562 = {{7{1'b0}}, col_in_562};
assign u_ca_in_563 = {{7{1'b0}}, col_in_563};
assign u_ca_in_564 = {{7{1'b0}}, col_in_564};
assign u_ca_in_565 = {{7{1'b0}}, col_in_565};
assign u_ca_in_566 = {{7{1'b0}}, col_in_566};
assign u_ca_in_567 = {{7{1'b0}}, col_in_567};
assign u_ca_in_568 = {{7{1'b0}}, col_in_568};
assign u_ca_in_569 = {{7{1'b0}}, col_in_569};
assign u_ca_in_570 = {{7{1'b0}}, col_in_570};
assign u_ca_in_571 = {{7{1'b0}}, col_in_571};
assign u_ca_in_572 = {{7{1'b0}}, col_in_572};
assign u_ca_in_573 = {{7{1'b0}}, col_in_573};
assign u_ca_in_574 = {{7{1'b0}}, col_in_574};
assign u_ca_in_575 = {{7{1'b0}}, col_in_575};
assign u_ca_in_576 = {{7{1'b0}}, col_in_576};
assign u_ca_in_577 = {{7{1'b0}}, col_in_577};
assign u_ca_in_578 = {{7{1'b0}}, col_in_578};
assign u_ca_in_579 = {{7{1'b0}}, col_in_579};
assign u_ca_in_580 = {{7{1'b0}}, col_in_580};
assign u_ca_in_581 = {{7{1'b0}}, col_in_581};
assign u_ca_in_582 = {{7{1'b0}}, col_in_582};
assign u_ca_in_583 = {{7{1'b0}}, col_in_583};
assign u_ca_in_584 = {{7{1'b0}}, col_in_584};
assign u_ca_in_585 = {{7{1'b0}}, col_in_585};
assign u_ca_in_586 = {{7{1'b0}}, col_in_586};
assign u_ca_in_587 = {{7{1'b0}}, col_in_587};
assign u_ca_in_588 = {{7{1'b0}}, col_in_588};
assign u_ca_in_589 = {{7{1'b0}}, col_in_589};
assign u_ca_in_590 = {{7{1'b0}}, col_in_590};
assign u_ca_in_591 = {{7{1'b0}}, col_in_591};
assign u_ca_in_592 = {{7{1'b0}}, col_in_592};
assign u_ca_in_593 = {{7{1'b0}}, col_in_593};
assign u_ca_in_594 = {{7{1'b0}}, col_in_594};
assign u_ca_in_595 = {{7{1'b0}}, col_in_595};
assign u_ca_in_596 = {{7{1'b0}}, col_in_596};
assign u_ca_in_597 = {{7{1'b0}}, col_in_597};
assign u_ca_in_598 = {{7{1'b0}}, col_in_598};
assign u_ca_in_599 = {{7{1'b0}}, col_in_599};
assign u_ca_in_600 = {{7{1'b0}}, col_in_600};
assign u_ca_in_601 = {{7{1'b0}}, col_in_601};
assign u_ca_in_602 = {{7{1'b0}}, col_in_602};
assign u_ca_in_603 = {{7{1'b0}}, col_in_603};
assign u_ca_in_604 = {{7{1'b0}}, col_in_604};
assign u_ca_in_605 = {{7{1'b0}}, col_in_605};
assign u_ca_in_606 = {{7{1'b0}}, col_in_606};
assign u_ca_in_607 = {{7{1'b0}}, col_in_607};
assign u_ca_in_608 = {{7{1'b0}}, col_in_608};
assign u_ca_in_609 = {{7{1'b0}}, col_in_609};
assign u_ca_in_610 = {{7{1'b0}}, col_in_610};
assign u_ca_in_611 = {{7{1'b0}}, col_in_611};
assign u_ca_in_612 = {{7{1'b0}}, col_in_612};
assign u_ca_in_613 = {{7{1'b0}}, col_in_613};
assign u_ca_in_614 = {{7{1'b0}}, col_in_614};
assign u_ca_in_615 = {{7{1'b0}}, col_in_615};
assign u_ca_in_616 = {{7{1'b0}}, col_in_616};
assign u_ca_in_617 = {{7{1'b0}}, col_in_617};
assign u_ca_in_618 = {{7{1'b0}}, col_in_618};
assign u_ca_in_619 = {{7{1'b0}}, col_in_619};
assign u_ca_in_620 = {{7{1'b0}}, col_in_620};
assign u_ca_in_621 = {{7{1'b0}}, col_in_621};
assign u_ca_in_622 = {{7{1'b0}}, col_in_622};
assign u_ca_in_623 = {{7{1'b0}}, col_in_623};
assign u_ca_in_624 = {{7{1'b0}}, col_in_624};
assign u_ca_in_625 = {{7{1'b0}}, col_in_625};
assign u_ca_in_626 = {{7{1'b0}}, col_in_626};
assign u_ca_in_627 = {{7{1'b0}}, col_in_627};
assign u_ca_in_628 = {{7{1'b0}}, col_in_628};
assign u_ca_in_629 = {{7{1'b0}}, col_in_629};
assign u_ca_in_630 = {{7{1'b0}}, col_in_630};
assign u_ca_in_631 = {{7{1'b0}}, col_in_631};
assign u_ca_in_632 = {{7{1'b0}}, col_in_632};
assign u_ca_in_633 = {{7{1'b0}}, col_in_633};
assign u_ca_in_634 = {{7{1'b0}}, col_in_634};
assign u_ca_in_635 = {{7{1'b0}}, col_in_635};
assign u_ca_in_636 = {{7{1'b0}}, col_in_636};
assign u_ca_in_637 = {{7{1'b0}}, col_in_637};
assign u_ca_in_638 = {{7{1'b0}}, col_in_638};
assign u_ca_in_639 = {{7{1'b0}}, col_in_639};
assign u_ca_in_640 = {{7{1'b0}}, col_in_640};
assign u_ca_in_641 = {{7{1'b0}}, col_in_641};
assign u_ca_in_642 = {{7{1'b0}}, col_in_642};
assign u_ca_in_643 = {{7{1'b0}}, col_in_643};
assign u_ca_in_644 = {{7{1'b0}}, col_in_644};
assign u_ca_in_645 = {{7{1'b0}}, col_in_645};
assign u_ca_in_646 = {{7{1'b0}}, col_in_646};
assign u_ca_in_647 = {{7{1'b0}}, col_in_647};
assign u_ca_in_648 = {{7{1'b0}}, col_in_648};
assign u_ca_in_649 = {{7{1'b0}}, col_in_649};
assign u_ca_in_650 = {{7{1'b0}}, col_in_650};
assign u_ca_in_651 = {{7{1'b0}}, col_in_651};
assign u_ca_in_652 = {{7{1'b0}}, col_in_652};
assign u_ca_in_653 = {{7{1'b0}}, col_in_653};
assign u_ca_in_654 = {{7{1'b0}}, col_in_654};
assign u_ca_in_655 = {{7{1'b0}}, col_in_655};
assign u_ca_in_656 = {{7{1'b0}}, col_in_656};
assign u_ca_in_657 = {{7{1'b0}}, col_in_657};
assign u_ca_in_658 = {{7{1'b0}}, col_in_658};
assign u_ca_in_659 = {{7{1'b0}}, col_in_659};
assign u_ca_in_660 = {{7{1'b0}}, col_in_660};
assign u_ca_in_661 = {{7{1'b0}}, col_in_661};
assign u_ca_in_662 = {{7{1'b0}}, col_in_662};
assign u_ca_in_663 = {{7{1'b0}}, col_in_663};
assign u_ca_in_664 = {{7{1'b0}}, col_in_664};
assign u_ca_in_665 = {{7{1'b0}}, col_in_665};
assign u_ca_in_666 = {{7{1'b0}}, col_in_666};
assign u_ca_in_667 = {{7{1'b0}}, col_in_667};
assign u_ca_in_668 = {{7{1'b0}}, col_in_668};
assign u_ca_in_669 = {{7{1'b0}}, col_in_669};
assign u_ca_in_670 = {{7{1'b0}}, col_in_670};
assign u_ca_in_671 = {{7{1'b0}}, col_in_671};
assign u_ca_in_672 = {{7{1'b0}}, col_in_672};
assign u_ca_in_673 = {{7{1'b0}}, col_in_673};
assign u_ca_in_674 = {{7{1'b0}}, col_in_674};
assign u_ca_in_675 = {{7{1'b0}}, col_in_675};
assign u_ca_in_676 = {{7{1'b0}}, col_in_676};
assign u_ca_in_677 = {{7{1'b0}}, col_in_677};
assign u_ca_in_678 = {{7{1'b0}}, col_in_678};
assign u_ca_in_679 = {{7{1'b0}}, col_in_679};
assign u_ca_in_680 = {{7{1'b0}}, col_in_680};
assign u_ca_in_681 = {{7{1'b0}}, col_in_681};
assign u_ca_in_682 = {{7{1'b0}}, col_in_682};
assign u_ca_in_683 = {{7{1'b0}}, col_in_683};
assign u_ca_in_684 = {{7{1'b0}}, col_in_684};
assign u_ca_in_685 = {{7{1'b0}}, col_in_685};
assign u_ca_in_686 = {{7{1'b0}}, col_in_686};
assign u_ca_in_687 = {{7{1'b0}}, col_in_687};
assign u_ca_in_688 = {{7{1'b0}}, col_in_688};
assign u_ca_in_689 = {{7{1'b0}}, col_in_689};
assign u_ca_in_690 = {{7{1'b0}}, col_in_690};
assign u_ca_in_691 = {{7{1'b0}}, col_in_691};
assign u_ca_in_692 = {{7{1'b0}}, col_in_692};
assign u_ca_in_693 = {{7{1'b0}}, col_in_693};
assign u_ca_in_694 = {{7{1'b0}}, col_in_694};
assign u_ca_in_695 = {{7{1'b0}}, col_in_695};
assign u_ca_in_696 = {{7{1'b0}}, col_in_696};
assign u_ca_in_697 = {{7{1'b0}}, col_in_697};
assign u_ca_in_698 = {{7{1'b0}}, col_in_698};
assign u_ca_in_699 = {{7{1'b0}}, col_in_699};
assign u_ca_in_700 = {{7{1'b0}}, col_in_700};
assign u_ca_in_701 = {{7{1'b0}}, col_in_701};
assign u_ca_in_702 = {{7{1'b0}}, col_in_702};
assign u_ca_in_703 = {{7{1'b0}}, col_in_703};
assign u_ca_in_704 = {{7{1'b0}}, col_in_704};
assign u_ca_in_705 = {{7{1'b0}}, col_in_705};
assign u_ca_in_706 = {{7{1'b0}}, col_in_706};
assign u_ca_in_707 = {{7{1'b0}}, col_in_707};
assign u_ca_in_708 = {{7{1'b0}}, col_in_708};
assign u_ca_in_709 = {{7{1'b0}}, col_in_709};
assign u_ca_in_710 = {{7{1'b0}}, col_in_710};
assign u_ca_in_711 = {{7{1'b0}}, col_in_711};
assign u_ca_in_712 = {{7{1'b0}}, col_in_712};
assign u_ca_in_713 = {{7{1'b0}}, col_in_713};
assign u_ca_in_714 = {{7{1'b0}}, col_in_714};
assign u_ca_in_715 = {{7{1'b0}}, col_in_715};
assign u_ca_in_716 = {{7{1'b0}}, col_in_716};
assign u_ca_in_717 = {{7{1'b0}}, col_in_717};
assign u_ca_in_718 = {{7{1'b0}}, col_in_718};
assign u_ca_in_719 = {{7{1'b0}}, col_in_719};
assign u_ca_in_720 = {{7{1'b0}}, col_in_720};
assign u_ca_in_721 = {{7{1'b0}}, col_in_721};
assign u_ca_in_722 = {{7{1'b0}}, col_in_722};
assign u_ca_in_723 = {{7{1'b0}}, col_in_723};
assign u_ca_in_724 = {{7{1'b0}}, col_in_724};
assign u_ca_in_725 = {{7{1'b0}}, col_in_725};
assign u_ca_in_726 = {{7{1'b0}}, col_in_726};
assign u_ca_in_727 = {{7{1'b0}}, col_in_727};
assign u_ca_in_728 = {{7{1'b0}}, col_in_728};
assign u_ca_in_729 = {{7{1'b0}}, col_in_729};
assign u_ca_in_730 = {{7{1'b0}}, col_in_730};
assign u_ca_in_731 = {{7{1'b0}}, col_in_731};
assign u_ca_in_732 = {{7{1'b0}}, col_in_732};
assign u_ca_in_733 = {{7{1'b0}}, col_in_733};
assign u_ca_in_734 = {{7{1'b0}}, col_in_734};
assign u_ca_in_735 = {{7{1'b0}}, col_in_735};
assign u_ca_in_736 = {{7{1'b0}}, col_in_736};
assign u_ca_in_737 = {{7{1'b0}}, col_in_737};
assign u_ca_in_738 = {{7{1'b0}}, col_in_738};
assign u_ca_in_739 = {{7{1'b0}}, col_in_739};
assign u_ca_in_740 = {{7{1'b0}}, col_in_740};
assign u_ca_in_741 = {{7{1'b0}}, col_in_741};
assign u_ca_in_742 = {{7{1'b0}}, col_in_742};
assign u_ca_in_743 = {{7{1'b0}}, col_in_743};
assign u_ca_in_744 = {{7{1'b0}}, col_in_744};
assign u_ca_in_745 = {{7{1'b0}}, col_in_745};
assign u_ca_in_746 = {{7{1'b0}}, col_in_746};
assign u_ca_in_747 = {{7{1'b0}}, col_in_747};
assign u_ca_in_748 = {{7{1'b0}}, col_in_748};
assign u_ca_in_749 = {{7{1'b0}}, col_in_749};
assign u_ca_in_750 = {{7{1'b0}}, col_in_750};
assign u_ca_in_751 = {{7{1'b0}}, col_in_751};
assign u_ca_in_752 = {{7{1'b0}}, col_in_752};
assign u_ca_in_753 = {{7{1'b0}}, col_in_753};
assign u_ca_in_754 = {{7{1'b0}}, col_in_754};
assign u_ca_in_755 = {{7{1'b0}}, col_in_755};
assign u_ca_in_756 = {{7{1'b0}}, col_in_756};
assign u_ca_in_757 = {{7{1'b0}}, col_in_757};
assign u_ca_in_758 = {{7{1'b0}}, col_in_758};
assign u_ca_in_759 = {{7{1'b0}}, col_in_759};
assign u_ca_in_760 = {{7{1'b0}}, col_in_760};
assign u_ca_in_761 = {{7{1'b0}}, col_in_761};
assign u_ca_in_762 = {{7{1'b0}}, col_in_762};
assign u_ca_in_763 = {{7{1'b0}}, col_in_763};
assign u_ca_in_764 = {{7{1'b0}}, col_in_764};
assign u_ca_in_765 = {{7{1'b0}}, col_in_765};
assign u_ca_in_766 = {{7{1'b0}}, col_in_766};
assign u_ca_in_767 = {{7{1'b0}}, col_in_767};
assign u_ca_in_768 = {{7{1'b0}}, col_in_768};
assign u_ca_in_769 = {{7{1'b0}}, col_in_769};
assign u_ca_in_770 = {{7{1'b0}}, col_in_770};
assign u_ca_in_771 = {{7{1'b0}}, col_in_771};
assign u_ca_in_772 = {{7{1'b0}}, col_in_772};
assign u_ca_in_773 = {{7{1'b0}}, col_in_773};
assign u_ca_in_774 = {{7{1'b0}}, col_in_774};
assign u_ca_in_775 = {{7{1'b0}}, col_in_775};
assign u_ca_in_776 = {{7{1'b0}}, col_in_776};
assign u_ca_in_777 = {{7{1'b0}}, col_in_777};
assign u_ca_in_778 = {{7{1'b0}}, col_in_778};
assign u_ca_in_779 = {{7{1'b0}}, col_in_779};
assign u_ca_in_780 = {{7{1'b0}}, col_in_780};
assign u_ca_in_781 = {{7{1'b0}}, col_in_781};
assign u_ca_in_782 = {{7{1'b0}}, col_in_782};
assign u_ca_in_783 = {{7{1'b0}}, col_in_783};
assign u_ca_in_784 = {{7{1'b0}}, col_in_784};
assign u_ca_in_785 = {{7{1'b0}}, col_in_785};
assign u_ca_in_786 = {{7{1'b0}}, col_in_786};
assign u_ca_in_787 = {{7{1'b0}}, col_in_787};
assign u_ca_in_788 = {{7{1'b0}}, col_in_788};
assign u_ca_in_789 = {{7{1'b0}}, col_in_789};
assign u_ca_in_790 = {{7{1'b0}}, col_in_790};
assign u_ca_in_791 = {{7{1'b0}}, col_in_791};
assign u_ca_in_792 = {{7{1'b0}}, col_in_792};
assign u_ca_in_793 = {{7{1'b0}}, col_in_793};
assign u_ca_in_794 = {{7{1'b0}}, col_in_794};
assign u_ca_in_795 = {{7{1'b0}}, col_in_795};
assign u_ca_in_796 = {{7{1'b0}}, col_in_796};
assign u_ca_in_797 = {{7{1'b0}}, col_in_797};
assign u_ca_in_798 = {{7{1'b0}}, col_in_798};
assign u_ca_in_799 = {{7{1'b0}}, col_in_799};
assign u_ca_in_800 = {{7{1'b0}}, col_in_800};
assign u_ca_in_801 = {{7{1'b0}}, col_in_801};
assign u_ca_in_802 = {{7{1'b0}}, col_in_802};
assign u_ca_in_803 = {{7{1'b0}}, col_in_803};
assign u_ca_in_804 = {{7{1'b0}}, col_in_804};
assign u_ca_in_805 = {{7{1'b0}}, col_in_805};
assign u_ca_in_806 = {{7{1'b0}}, col_in_806};
assign u_ca_in_807 = {{7{1'b0}}, col_in_807};
assign u_ca_in_808 = {{7{1'b0}}, col_in_808};
assign u_ca_in_809 = {{7{1'b0}}, col_in_809};
assign u_ca_in_810 = {{7{1'b0}}, col_in_810};
assign u_ca_in_811 = {{7{1'b0}}, col_in_811};
assign u_ca_in_812 = {{7{1'b0}}, col_in_812};
assign u_ca_in_813 = {{7{1'b0}}, col_in_813};
assign u_ca_in_814 = {{7{1'b0}}, col_in_814};
assign u_ca_in_815 = {{7{1'b0}}, col_in_815};
assign u_ca_in_816 = {{7{1'b0}}, col_in_816};
assign u_ca_in_817 = {{7{1'b0}}, col_in_817};
assign u_ca_in_818 = {{7{1'b0}}, col_in_818};
assign u_ca_in_819 = {{7{1'b0}}, col_in_819};
assign u_ca_in_820 = {{7{1'b0}}, col_in_820};
assign u_ca_in_821 = {{7{1'b0}}, col_in_821};
assign u_ca_in_822 = {{7{1'b0}}, col_in_822};
assign u_ca_in_823 = {{7{1'b0}}, col_in_823};
assign u_ca_in_824 = {{7{1'b0}}, col_in_824};
assign u_ca_in_825 = {{7{1'b0}}, col_in_825};
assign u_ca_in_826 = {{7{1'b0}}, col_in_826};
assign u_ca_in_827 = {{7{1'b0}}, col_in_827};
assign u_ca_in_828 = {{7{1'b0}}, col_in_828};
assign u_ca_in_829 = {{7{1'b0}}, col_in_829};
assign u_ca_in_830 = {{7{1'b0}}, col_in_830};
assign u_ca_in_831 = {{7{1'b0}}, col_in_831};
assign u_ca_in_832 = {{7{1'b0}}, col_in_832};
assign u_ca_in_833 = {{7{1'b0}}, col_in_833};
assign u_ca_in_834 = {{7{1'b0}}, col_in_834};
assign u_ca_in_835 = {{7{1'b0}}, col_in_835};
assign u_ca_in_836 = {{7{1'b0}}, col_in_836};
assign u_ca_in_837 = {{7{1'b0}}, col_in_837};
assign u_ca_in_838 = {{7{1'b0}}, col_in_838};
assign u_ca_in_839 = {{7{1'b0}}, col_in_839};
assign u_ca_in_840 = {{7{1'b0}}, col_in_840};
assign u_ca_in_841 = {{7{1'b0}}, col_in_841};
assign u_ca_in_842 = {{7{1'b0}}, col_in_842};
assign u_ca_in_843 = {{7{1'b0}}, col_in_843};
assign u_ca_in_844 = {{7{1'b0}}, col_in_844};
assign u_ca_in_845 = {{7{1'b0}}, col_in_845};
assign u_ca_in_846 = {{7{1'b0}}, col_in_846};
assign u_ca_in_847 = {{7{1'b0}}, col_in_847};
assign u_ca_in_848 = {{7{1'b0}}, col_in_848};
assign u_ca_in_849 = {{7{1'b0}}, col_in_849};
assign u_ca_in_850 = {{7{1'b0}}, col_in_850};
assign u_ca_in_851 = {{7{1'b0}}, col_in_851};
assign u_ca_in_852 = {{7{1'b0}}, col_in_852};
assign u_ca_in_853 = {{7{1'b0}}, col_in_853};
assign u_ca_in_854 = {{7{1'b0}}, col_in_854};
assign u_ca_in_855 = {{7{1'b0}}, col_in_855};
assign u_ca_in_856 = {{7{1'b0}}, col_in_856};
assign u_ca_in_857 = {{7{1'b0}}, col_in_857};
assign u_ca_in_858 = {{7{1'b0}}, col_in_858};
assign u_ca_in_859 = {{7{1'b0}}, col_in_859};
assign u_ca_in_860 = {{7{1'b0}}, col_in_860};
assign u_ca_in_861 = {{7{1'b0}}, col_in_861};
assign u_ca_in_862 = {{7{1'b0}}, col_in_862};
assign u_ca_in_863 = {{7{1'b0}}, col_in_863};
assign u_ca_in_864 = {{7{1'b0}}, col_in_864};
assign u_ca_in_865 = {{7{1'b0}}, col_in_865};
assign u_ca_in_866 = {{7{1'b0}}, col_in_866};
assign u_ca_in_867 = {{7{1'b0}}, col_in_867};
assign u_ca_in_868 = {{7{1'b0}}, col_in_868};
assign u_ca_in_869 = {{7{1'b0}}, col_in_869};
assign u_ca_in_870 = {{7{1'b0}}, col_in_870};
assign u_ca_in_871 = {{7{1'b0}}, col_in_871};
assign u_ca_in_872 = {{7{1'b0}}, col_in_872};
assign u_ca_in_873 = {{7{1'b0}}, col_in_873};
assign u_ca_in_874 = {{7{1'b0}}, col_in_874};
assign u_ca_in_875 = {{7{1'b0}}, col_in_875};
assign u_ca_in_876 = {{7{1'b0}}, col_in_876};
assign u_ca_in_877 = {{7{1'b0}}, col_in_877};
assign u_ca_in_878 = {{7{1'b0}}, col_in_878};
assign u_ca_in_879 = {{7{1'b0}}, col_in_879};
assign u_ca_in_880 = {{7{1'b0}}, col_in_880};
assign u_ca_in_881 = {{7{1'b0}}, col_in_881};
assign u_ca_in_882 = {{7{1'b0}}, col_in_882};
assign u_ca_in_883 = {{7{1'b0}}, col_in_883};
assign u_ca_in_884 = {{7{1'b0}}, col_in_884};
assign u_ca_in_885 = {{7{1'b0}}, col_in_885};
assign u_ca_in_886 = {{7{1'b0}}, col_in_886};
assign u_ca_in_887 = {{7{1'b0}}, col_in_887};
assign u_ca_in_888 = {{7{1'b0}}, col_in_888};
assign u_ca_in_889 = {{7{1'b0}}, col_in_889};
assign u_ca_in_890 = {{7{1'b0}}, col_in_890};
assign u_ca_in_891 = {{7{1'b0}}, col_in_891};
assign u_ca_in_892 = {{7{1'b0}}, col_in_892};
assign u_ca_in_893 = {{7{1'b0}}, col_in_893};
assign u_ca_in_894 = {{7{1'b0}}, col_in_894};
assign u_ca_in_895 = {{7{1'b0}}, col_in_895};
assign u_ca_in_896 = {{7{1'b0}}, col_in_896};
assign u_ca_in_897 = {{7{1'b0}}, col_in_897};
assign u_ca_in_898 = {{7{1'b0}}, col_in_898};
assign u_ca_in_899 = {{7{1'b0}}, col_in_899};
assign u_ca_in_900 = {{7{1'b0}}, col_in_900};
assign u_ca_in_901 = {{7{1'b0}}, col_in_901};
assign u_ca_in_902 = {{7{1'b0}}, col_in_902};
assign u_ca_in_903 = {{7{1'b0}}, col_in_903};
assign u_ca_in_904 = {{7{1'b0}}, col_in_904};
assign u_ca_in_905 = {{7{1'b0}}, col_in_905};
assign u_ca_in_906 = {{7{1'b0}}, col_in_906};
assign u_ca_in_907 = {{7{1'b0}}, col_in_907};
assign u_ca_in_908 = {{7{1'b0}}, col_in_908};
assign u_ca_in_909 = {{7{1'b0}}, col_in_909};
assign u_ca_in_910 = {{7{1'b0}}, col_in_910};
assign u_ca_in_911 = {{7{1'b0}}, col_in_911};
assign u_ca_in_912 = {{7{1'b0}}, col_in_912};
assign u_ca_in_913 = {{7{1'b0}}, col_in_913};
assign u_ca_in_914 = {{7{1'b0}}, col_in_914};
assign u_ca_in_915 = {{7{1'b0}}, col_in_915};
assign u_ca_in_916 = {{7{1'b0}}, col_in_916};
assign u_ca_in_917 = {{7{1'b0}}, col_in_917};
assign u_ca_in_918 = {{7{1'b0}}, col_in_918};
assign u_ca_in_919 = {{7{1'b0}}, col_in_919};
assign u_ca_in_920 = {{7{1'b0}}, col_in_920};
assign u_ca_in_921 = {{7{1'b0}}, col_in_921};
assign u_ca_in_922 = {{7{1'b0}}, col_in_922};
assign u_ca_in_923 = {{7{1'b0}}, col_in_923};
assign u_ca_in_924 = {{7{1'b0}}, col_in_924};
assign u_ca_in_925 = {{7{1'b0}}, col_in_925};
assign u_ca_in_926 = {{7{1'b0}}, col_in_926};
assign u_ca_in_927 = {{7{1'b0}}, col_in_927};
assign u_ca_in_928 = {{7{1'b0}}, col_in_928};
assign u_ca_in_929 = {{7{1'b0}}, col_in_929};
assign u_ca_in_930 = {{7{1'b0}}, col_in_930};
assign u_ca_in_931 = {{7{1'b0}}, col_in_931};
assign u_ca_in_932 = {{7{1'b0}}, col_in_932};
assign u_ca_in_933 = {{7{1'b0}}, col_in_933};
assign u_ca_in_934 = {{7{1'b0}}, col_in_934};
assign u_ca_in_935 = {{7{1'b0}}, col_in_935};
assign u_ca_in_936 = {{7{1'b0}}, col_in_936};
assign u_ca_in_937 = {{7{1'b0}}, col_in_937};
assign u_ca_in_938 = {{7{1'b0}}, col_in_938};
assign u_ca_in_939 = {{7{1'b0}}, col_in_939};
assign u_ca_in_940 = {{7{1'b0}}, col_in_940};
assign u_ca_in_941 = {{7{1'b0}}, col_in_941};
assign u_ca_in_942 = {{7{1'b0}}, col_in_942};
assign u_ca_in_943 = {{7{1'b0}}, col_in_943};
assign u_ca_in_944 = {{7{1'b0}}, col_in_944};
assign u_ca_in_945 = {{7{1'b0}}, col_in_945};
assign u_ca_in_946 = {{7{1'b0}}, col_in_946};
assign u_ca_in_947 = {{7{1'b0}}, col_in_947};
assign u_ca_in_948 = {{7{1'b0}}, col_in_948};
assign u_ca_in_949 = {{7{1'b0}}, col_in_949};
assign u_ca_in_950 = {{7{1'b0}}, col_in_950};
assign u_ca_in_951 = {{7{1'b0}}, col_in_951};
assign u_ca_in_952 = {{7{1'b0}}, col_in_952};
assign u_ca_in_953 = {{7{1'b0}}, col_in_953};
assign u_ca_in_954 = {{7{1'b0}}, col_in_954};
assign u_ca_in_955 = {{7{1'b0}}, col_in_955};
assign u_ca_in_956 = {{7{1'b0}}, col_in_956};
assign u_ca_in_957 = {{7{1'b0}}, col_in_957};
assign u_ca_in_958 = {{7{1'b0}}, col_in_958};
assign u_ca_in_959 = {{7{1'b0}}, col_in_959};
assign u_ca_in_960 = {{7{1'b0}}, col_in_960};
assign u_ca_in_961 = {{7{1'b0}}, col_in_961};
assign u_ca_in_962 = {{7{1'b0}}, col_in_962};
assign u_ca_in_963 = {{7{1'b0}}, col_in_963};
assign u_ca_in_964 = {{7{1'b0}}, col_in_964};
assign u_ca_in_965 = {{7{1'b0}}, col_in_965};
assign u_ca_in_966 = {{7{1'b0}}, col_in_966};
assign u_ca_in_967 = {{7{1'b0}}, col_in_967};
assign u_ca_in_968 = {{7{1'b0}}, col_in_968};
assign u_ca_in_969 = {{7{1'b0}}, col_in_969};
assign u_ca_in_970 = {{7{1'b0}}, col_in_970};
assign u_ca_in_971 = {{7{1'b0}}, col_in_971};
assign u_ca_in_972 = {{7{1'b0}}, col_in_972};
assign u_ca_in_973 = {{7{1'b0}}, col_in_973};
assign u_ca_in_974 = {{7{1'b0}}, col_in_974};
assign u_ca_in_975 = {{7{1'b0}}, col_in_975};
assign u_ca_in_976 = {{7{1'b0}}, col_in_976};
assign u_ca_in_977 = {{7{1'b0}}, col_in_977};
assign u_ca_in_978 = {{7{1'b0}}, col_in_978};
assign u_ca_in_979 = {{7{1'b0}}, col_in_979};
assign u_ca_in_980 = {{7{1'b0}}, col_in_980};
assign u_ca_in_981 = {{7{1'b0}}, col_in_981};
assign u_ca_in_982 = {{7{1'b0}}, col_in_982};
assign u_ca_in_983 = {{7{1'b0}}, col_in_983};
assign u_ca_in_984 = {{7{1'b0}}, col_in_984};
assign u_ca_in_985 = {{7{1'b0}}, col_in_985};
assign u_ca_in_986 = {{7{1'b0}}, col_in_986};
assign u_ca_in_987 = {{7{1'b0}}, col_in_987};
assign u_ca_in_988 = {{7{1'b0}}, col_in_988};
assign u_ca_in_989 = {{7{1'b0}}, col_in_989};
assign u_ca_in_990 = {{7{1'b0}}, col_in_990};
assign u_ca_in_991 = {{7{1'b0}}, col_in_991};
assign u_ca_in_992 = {{7{1'b0}}, col_in_992};
assign u_ca_in_993 = {{7{1'b0}}, col_in_993};
assign u_ca_in_994 = {{7{1'b0}}, col_in_994};
assign u_ca_in_995 = {{7{1'b0}}, col_in_995};
assign u_ca_in_996 = {{7{1'b0}}, col_in_996};
assign u_ca_in_997 = {{7{1'b0}}, col_in_997};
assign u_ca_in_998 = {{7{1'b0}}, col_in_998};
assign u_ca_in_999 = {{7{1'b0}}, col_in_999};
assign u_ca_in_1000 = {{7{1'b0}}, col_in_1000};
assign u_ca_in_1001 = {{7{1'b0}}, col_in_1001};
assign u_ca_in_1002 = {{7{1'b0}}, col_in_1002};
assign u_ca_in_1003 = {{7{1'b0}}, col_in_1003};
assign u_ca_in_1004 = {{7{1'b0}}, col_in_1004};
assign u_ca_in_1005 = {{7{1'b0}}, col_in_1005};
assign u_ca_in_1006 = {{7{1'b0}}, col_in_1006};
assign u_ca_in_1007 = {{7{1'b0}}, col_in_1007};
assign u_ca_in_1008 = {{7{1'b0}}, col_in_1008};
assign u_ca_in_1009 = {{7{1'b0}}, col_in_1009};
assign u_ca_in_1010 = {{7{1'b0}}, col_in_1010};
assign u_ca_in_1011 = {{7{1'b0}}, col_in_1011};
assign u_ca_in_1012 = {{7{1'b0}}, col_in_1012};
assign u_ca_in_1013 = {{7{1'b0}}, col_in_1013};
assign u_ca_in_1014 = {{7{1'b0}}, col_in_1014};
assign u_ca_in_1015 = {{7{1'b0}}, col_in_1015};
assign u_ca_in_1016 = {{7{1'b0}}, col_in_1016};
assign u_ca_in_1017 = {{7{1'b0}}, col_in_1017};
assign u_ca_in_1018 = {{7{1'b0}}, col_in_1018};
assign u_ca_in_1019 = {{7{1'b0}}, col_in_1019};
assign u_ca_in_1020 = {{7{1'b0}}, col_in_1020};
assign u_ca_in_1021 = {{7{1'b0}}, col_in_1021};
assign u_ca_in_1022 = {{7{1'b0}}, col_in_1022};
assign u_ca_in_1023 = {{7{1'b0}}, col_in_1023};
assign u_ca_in_1024 = {{7{1'b0}}, col_in_1024};
assign u_ca_in_1025 = {{7{1'b0}}, col_in_1025};
assign u_ca_in_1026 = {{7{1'b0}}, col_in_1026};
assign u_ca_in_1027 = {{7{1'b0}}, col_in_1027};
assign u_ca_in_1028 = {{7{1'b0}}, col_in_1028};
assign u_ca_in_1029 = {{7{1'b0}}, col_in_1029};
assign u_ca_in_1030 = {{7{1'b0}}, col_in_1030};
assign u_ca_in_1031 = {{7{1'b0}}, col_in_1031};
assign u_ca_in_1032 = {{7{1'b0}}, col_in_1032};
assign u_ca_in_1033 = {{7{1'b0}}, col_in_1033};
assign u_ca_in_1034 = {{7{1'b0}}, col_in_1034};
assign u_ca_in_1035 = {{7{1'b0}}, col_in_1035};
assign u_ca_in_1036 = {{7{1'b0}}, col_in_1036};
assign u_ca_in_1037 = {{7{1'b0}}, col_in_1037};
assign u_ca_in_1038 = {{7{1'b0}}, col_in_1038};
assign u_ca_in_1039 = {{7{1'b0}}, col_in_1039};
assign u_ca_in_1040 = {{7{1'b0}}, col_in_1040};
assign u_ca_in_1041 = {{7{1'b0}}, col_in_1041};
assign u_ca_in_1042 = {{7{1'b0}}, col_in_1042};
assign u_ca_in_1043 = {{7{1'b0}}, col_in_1043};
assign u_ca_in_1044 = {{7{1'b0}}, col_in_1044};
assign u_ca_in_1045 = {{7{1'b0}}, col_in_1045};
assign u_ca_in_1046 = {{7{1'b0}}, col_in_1046};
assign u_ca_in_1047 = {{7{1'b0}}, col_in_1047};
assign u_ca_in_1048 = {{7{1'b0}}, col_in_1048};
assign u_ca_in_1049 = {{7{1'b0}}, col_in_1049};
assign u_ca_in_1050 = {{7{1'b0}}, col_in_1050};
assign u_ca_in_1051 = {{7{1'b0}}, col_in_1051};
assign u_ca_in_1052 = {{7{1'b0}}, col_in_1052};
assign u_ca_in_1053 = {{7{1'b0}}, col_in_1053};
assign u_ca_in_1054 = {{7{1'b0}}, col_in_1054};
assign u_ca_in_1055 = {{7{1'b0}}, col_in_1055};
assign u_ca_in_1056 = {{7{1'b0}}, col_in_1056};
assign u_ca_in_1057 = {{7{1'b0}}, col_in_1057};
assign u_ca_in_1058 = {{7{1'b0}}, col_in_1058};
assign u_ca_in_1059 = {{7{1'b0}}, col_in_1059};
assign u_ca_in_1060 = {{7{1'b0}}, col_in_1060};
assign u_ca_in_1061 = {{7{1'b0}}, col_in_1061};
assign u_ca_in_1062 = {{7{1'b0}}, col_in_1062};
assign u_ca_in_1063 = {{7{1'b0}}, col_in_1063};
assign u_ca_in_1064 = {{7{1'b0}}, col_in_1064};
assign u_ca_in_1065 = {{7{1'b0}}, col_in_1065};
assign u_ca_in_1066 = {{7{1'b0}}, col_in_1066};
assign u_ca_in_1067 = {{7{1'b0}}, col_in_1067};
assign u_ca_in_1068 = {{7{1'b0}}, col_in_1068};
assign u_ca_in_1069 = {{7{1'b0}}, col_in_1069};
assign u_ca_in_1070 = {{7{1'b0}}, col_in_1070};
assign u_ca_in_1071 = {{7{1'b0}}, col_in_1071};
assign u_ca_in_1072 = {{7{1'b0}}, col_in_1072};
assign u_ca_in_1073 = {{7{1'b0}}, col_in_1073};
assign u_ca_in_1074 = {{7{1'b0}}, col_in_1074};
assign u_ca_in_1075 = {{7{1'b0}}, col_in_1075};
assign u_ca_in_1076 = {{7{1'b0}}, col_in_1076};
assign u_ca_in_1077 = {{7{1'b0}}, col_in_1077};
assign u_ca_in_1078 = {{7{1'b0}}, col_in_1078};
assign u_ca_in_1079 = {{7{1'b0}}, col_in_1079};
assign u_ca_in_1080 = {{7{1'b0}}, col_in_1080};
assign u_ca_in_1081 = {{7{1'b0}}, col_in_1081};
assign u_ca_in_1082 = {{7{1'b0}}, col_in_1082};
assign u_ca_in_1083 = {{7{1'b0}}, col_in_1083};
assign u_ca_in_1084 = {{7{1'b0}}, col_in_1084};
assign u_ca_in_1085 = {{7{1'b0}}, col_in_1085};
assign u_ca_in_1086 = {{7{1'b0}}, col_in_1086};
assign u_ca_in_1087 = {{7{1'b0}}, col_in_1087};
assign u_ca_in_1088 = {{7{1'b0}}, col_in_1088};
assign u_ca_in_1089 = {{7{1'b0}}, col_in_1089};
assign u_ca_in_1090 = {{7{1'b0}}, col_in_1090};
assign u_ca_in_1091 = {{7{1'b0}}, col_in_1091};
assign u_ca_in_1092 = {{7{1'b0}}, col_in_1092};
assign u_ca_in_1093 = {{7{1'b0}}, col_in_1093};
assign u_ca_in_1094 = {{7{1'b0}}, col_in_1094};
assign u_ca_in_1095 = {{7{1'b0}}, col_in_1095};
assign u_ca_in_1096 = {{7{1'b0}}, col_in_1096};
assign u_ca_in_1097 = {{7{1'b0}}, col_in_1097};
assign u_ca_in_1098 = {{7{1'b0}}, col_in_1098};
assign u_ca_in_1099 = {{7{1'b0}}, col_in_1099};
assign u_ca_in_1100 = {{7{1'b0}}, col_in_1100};
assign u_ca_in_1101 = {{7{1'b0}}, col_in_1101};
assign u_ca_in_1102 = {{7{1'b0}}, col_in_1102};
assign u_ca_in_1103 = {{7{1'b0}}, col_in_1103};
assign u_ca_in_1104 = {{7{1'b0}}, col_in_1104};
assign u_ca_in_1105 = {{7{1'b0}}, col_in_1105};
assign u_ca_in_1106 = {{7{1'b0}}, col_in_1106};
assign u_ca_in_1107 = {{7{1'b0}}, col_in_1107};
assign u_ca_in_1108 = {{7{1'b0}}, col_in_1108};
assign u_ca_in_1109 = {{7{1'b0}}, col_in_1109};
assign u_ca_in_1110 = {{7{1'b0}}, col_in_1110};
assign u_ca_in_1111 = {{7{1'b0}}, col_in_1111};
assign u_ca_in_1112 = {{7{1'b0}}, col_in_1112};
assign u_ca_in_1113 = {{7{1'b0}}, col_in_1113};
assign u_ca_in_1114 = {{7{1'b0}}, col_in_1114};
assign u_ca_in_1115 = {{7{1'b0}}, col_in_1115};
assign u_ca_in_1116 = {{7{1'b0}}, col_in_1116};
assign u_ca_in_1117 = {{7{1'b0}}, col_in_1117};
assign u_ca_in_1118 = {{7{1'b0}}, col_in_1118};
assign u_ca_in_1119 = {{7{1'b0}}, col_in_1119};
assign u_ca_in_1120 = {{7{1'b0}}, col_in_1120};
assign u_ca_in_1121 = {{7{1'b0}}, col_in_1121};
assign u_ca_in_1122 = {{7{1'b0}}, col_in_1122};
assign u_ca_in_1123 = {{7{1'b0}}, col_in_1123};
assign u_ca_in_1124 = {{7{1'b0}}, col_in_1124};
assign u_ca_in_1125 = {{7{1'b0}}, col_in_1125};
assign u_ca_in_1126 = {{7{1'b0}}, col_in_1126};
assign u_ca_in_1127 = {{7{1'b0}}, col_in_1127};
assign u_ca_in_1128 = {{7{1'b0}}, col_in_1128};
assign u_ca_in_1129 = {{7{1'b0}}, col_in_1129};
assign u_ca_in_1130 = {{7{1'b0}}, col_in_1130};
assign u_ca_in_1131 = {{7{1'b0}}, col_in_1131};
assign u_ca_in_1132 = {{7{1'b0}}, col_in_1132};
assign u_ca_in_1133 = {{7{1'b0}}, col_in_1133};
assign u_ca_in_1134 = {{7{1'b0}}, col_in_1134};
assign u_ca_in_1135 = {{7{1'b0}}, col_in_1135};
assign u_ca_in_1136 = {{7{1'b0}}, col_in_1136};
assign u_ca_in_1137 = {{7{1'b0}}, col_in_1137};
assign u_ca_in_1138 = {{7{1'b0}}, col_in_1138};
assign u_ca_in_1139 = {{7{1'b0}}, col_in_1139};
assign u_ca_in_1140 = {{7{1'b0}}, col_in_1140};
assign u_ca_in_1141 = {{7{1'b0}}, col_in_1141};
assign u_ca_in_1142 = {{7{1'b0}}, col_in_1142};
assign u_ca_in_1143 = {{7{1'b0}}, col_in_1143};
assign u_ca_in_1144 = {{7{1'b0}}, col_in_1144};
assign u_ca_in_1145 = {{7{1'b0}}, col_in_1145};
assign u_ca_in_1146 = {{7{1'b0}}, col_in_1146};
assign u_ca_in_1147 = {{7{1'b0}}, col_in_1147};
assign u_ca_in_1148 = {{7{1'b0}}, col_in_1148};
assign u_ca_in_1149 = {{7{1'b0}}, col_in_1149};
assign u_ca_in_1150 = {{7{1'b0}}, col_in_1150};
assign u_ca_in_1151 = {{7{1'b0}}, col_in_1151};
assign u_ca_in_1152 = {{7{1'b0}}, col_in_1152};
assign u_ca_in_1153 = {{7{1'b0}}, col_in_1153};
assign u_ca_in_1154 = {{7{1'b0}}, col_in_1154};
assign u_ca_in_1155 = {{7{1'b0}}, col_in_1155};
assign u_ca_in_1156 = {{7{1'b0}}, col_in_1156};
assign u_ca_in_1157 = {{7{1'b0}}, col_in_1157};
assign u_ca_in_1158 = {{7{1'b0}}, col_in_1158};
assign u_ca_in_1159 = {{7{1'b0}}, col_in_1159};
assign u_ca_in_1160 = {{7{1'b0}}, col_in_1160};
assign u_ca_in_1161 = {{7{1'b0}}, col_in_1161};
assign u_ca_in_1162 = {{7{1'b0}}, col_in_1162};
assign u_ca_in_1163 = {{7{1'b0}}, col_in_1163};
assign u_ca_in_1164 = {{7{1'b0}}, col_in_1164};
assign u_ca_in_1165 = {{7{1'b0}}, col_in_1165};
assign u_ca_in_1166 = {{7{1'b0}}, col_in_1166};
assign u_ca_in_1167 = {{7{1'b0}}, col_in_1167};
assign u_ca_in_1168 = {{7{1'b0}}, col_in_1168};
assign u_ca_in_1169 = {{7{1'b0}}, col_in_1169};
assign u_ca_in_1170 = {{7{1'b0}}, col_in_1170};
assign u_ca_in_1171 = {{7{1'b0}}, col_in_1171};
assign u_ca_in_1172 = {{7{1'b0}}, col_in_1172};
assign u_ca_in_1173 = {{7{1'b0}}, col_in_1173};
assign u_ca_in_1174 = {{7{1'b0}}, col_in_1174};
assign u_ca_in_1175 = {{7{1'b0}}, col_in_1175};
assign u_ca_in_1176 = {{7{1'b0}}, col_in_1176};
assign u_ca_in_1177 = {{7{1'b0}}, col_in_1177};
assign u_ca_in_1178 = {{7{1'b0}}, col_in_1178};
assign u_ca_in_1179 = {{7{1'b0}}, col_in_1179};
assign u_ca_in_1180 = {{7{1'b0}}, col_in_1180};
assign u_ca_in_1181 = {{7{1'b0}}, col_in_1181};
assign u_ca_in_1182 = {{7{1'b0}}, col_in_1182};
assign u_ca_in_1183 = {{7{1'b0}}, col_in_1183};
assign u_ca_in_1184 = {{7{1'b0}}, col_in_1184};
assign u_ca_in_1185 = {{7{1'b0}}, col_in_1185};
assign u_ca_in_1186 = {{7{1'b0}}, col_in_1186};
assign u_ca_in_1187 = {{7{1'b0}}, col_in_1187};
assign u_ca_in_1188 = {{7{1'b0}}, col_in_1188};
assign u_ca_in_1189 = {{7{1'b0}}, col_in_1189};
assign u_ca_in_1190 = {{7{1'b0}}, col_in_1190};
assign u_ca_in_1191 = {{7{1'b0}}, col_in_1191};
assign u_ca_in_1192 = {{7{1'b0}}, col_in_1192};
assign u_ca_in_1193 = {{7{1'b0}}, col_in_1193};
assign u_ca_in_1194 = {{7{1'b0}}, col_in_1194};
assign u_ca_in_1195 = {{7{1'b0}}, col_in_1195};
assign u_ca_in_1196 = {{7{1'b0}}, col_in_1196};
assign u_ca_in_1197 = {{7{1'b0}}, col_in_1197};
assign u_ca_in_1198 = {{7{1'b0}}, col_in_1198};
assign u_ca_in_1199 = {{7{1'b0}}, col_in_1199};
assign u_ca_in_1200 = {{7{1'b0}}, col_in_1200};
assign u_ca_in_1201 = {{7{1'b0}}, col_in_1201};
assign u_ca_in_1202 = {{7{1'b0}}, col_in_1202};
assign u_ca_in_1203 = {{7{1'b0}}, col_in_1203};
assign u_ca_in_1204 = {{7{1'b0}}, col_in_1204};
assign u_ca_in_1205 = {{7{1'b0}}, col_in_1205};
assign u_ca_in_1206 = {{7{1'b0}}, col_in_1206};
assign u_ca_in_1207 = {{7{1'b0}}, col_in_1207};
assign u_ca_in_1208 = {{7{1'b0}}, col_in_1208};
assign u_ca_in_1209 = {{7{1'b0}}, col_in_1209};
assign u_ca_in_1210 = {{7{1'b0}}, col_in_1210};
assign u_ca_in_1211 = {{7{1'b0}}, col_in_1211};
assign u_ca_in_1212 = {{7{1'b0}}, col_in_1212};
assign u_ca_in_1213 = {{7{1'b0}}, col_in_1213};
assign u_ca_in_1214 = {{7{1'b0}}, col_in_1214};
assign u_ca_in_1215 = {{7{1'b0}}, col_in_1215};
assign u_ca_in_1216 = {{7{1'b0}}, col_in_1216};
assign u_ca_in_1217 = {{7{1'b0}}, col_in_1217};
assign u_ca_in_1218 = {{7{1'b0}}, col_in_1218};
assign u_ca_in_1219 = {{7{1'b0}}, col_in_1219};
assign u_ca_in_1220 = {{7{1'b0}}, col_in_1220};
assign u_ca_in_1221 = {{7{1'b0}}, col_in_1221};
assign u_ca_in_1222 = {{7{1'b0}}, col_in_1222};
assign u_ca_in_1223 = {{7{1'b0}}, col_in_1223};
assign u_ca_in_1224 = {{7{1'b0}}, col_in_1224};
assign u_ca_in_1225 = {{7{1'b0}}, col_in_1225};
assign u_ca_in_1226 = {{7{1'b0}}, col_in_1226};
assign u_ca_in_1227 = {{7{1'b0}}, col_in_1227};
assign u_ca_in_1228 = {{7{1'b0}}, col_in_1228};
assign u_ca_in_1229 = {{7{1'b0}}, col_in_1229};
assign u_ca_in_1230 = {{7{1'b0}}, col_in_1230};
assign u_ca_in_1231 = {{7{1'b0}}, col_in_1231};
assign u_ca_in_1232 = {{7{1'b0}}, col_in_1232};
assign u_ca_in_1233 = {{7{1'b0}}, col_in_1233};
assign u_ca_in_1234 = {{7{1'b0}}, col_in_1234};
assign u_ca_in_1235 = {{7{1'b0}}, col_in_1235};
assign u_ca_in_1236 = {{7{1'b0}}, col_in_1236};
assign u_ca_in_1237 = {{7{1'b0}}, col_in_1237};
assign u_ca_in_1238 = {{7{1'b0}}, col_in_1238};
assign u_ca_in_1239 = {{7{1'b0}}, col_in_1239};
assign u_ca_in_1240 = {{7{1'b0}}, col_in_1240};
assign u_ca_in_1241 = {{7{1'b0}}, col_in_1241};
assign u_ca_in_1242 = {{7{1'b0}}, col_in_1242};
assign u_ca_in_1243 = {{7{1'b0}}, col_in_1243};
assign u_ca_in_1244 = {{7{1'b0}}, col_in_1244};
assign u_ca_in_1245 = {{7{1'b0}}, col_in_1245};
assign u_ca_in_1246 = {{7{1'b0}}, col_in_1246};
assign u_ca_in_1247 = {{7{1'b0}}, col_in_1247};
assign u_ca_in_1248 = {{7{1'b0}}, col_in_1248};
assign u_ca_in_1249 = {{7{1'b0}}, col_in_1249};
assign u_ca_in_1250 = {{7{1'b0}}, col_in_1250};
assign u_ca_in_1251 = {{7{1'b0}}, col_in_1251};
assign u_ca_in_1252 = {{7{1'b0}}, col_in_1252};
assign u_ca_in_1253 = {{7{1'b0}}, col_in_1253};
assign u_ca_in_1254 = {{7{1'b0}}, col_in_1254};
assign u_ca_in_1255 = {{7{1'b0}}, col_in_1255};
assign u_ca_in_1256 = {{7{1'b0}}, col_in_1256};
assign u_ca_in_1257 = {{7{1'b0}}, col_in_1257};
assign u_ca_in_1258 = {{7{1'b0}}, col_in_1258};
assign u_ca_in_1259 = {{7{1'b0}}, col_in_1259};
assign u_ca_in_1260 = {{7{1'b0}}, col_in_1260};
assign u_ca_in_1261 = {{7{1'b0}}, col_in_1261};
assign u_ca_in_1262 = {{7{1'b0}}, col_in_1262};
assign u_ca_in_1263 = {{7{1'b0}}, col_in_1263};
assign u_ca_in_1264 = {{7{1'b0}}, col_in_1264};
assign u_ca_in_1265 = {{7{1'b0}}, col_in_1265};
assign u_ca_in_1266 = {{7{1'b0}}, col_in_1266};
assign u_ca_in_1267 = {{7{1'b0}}, col_in_1267};
assign u_ca_in_1268 = {{7{1'b0}}, col_in_1268};
assign u_ca_in_1269 = {{7{1'b0}}, col_in_1269};
assign u_ca_in_1270 = {{7{1'b0}}, col_in_1270};
assign u_ca_in_1271 = {{7{1'b0}}, col_in_1271};
assign u_ca_in_1272 = {{7{1'b0}}, col_in_1272};
assign u_ca_in_1273 = {{7{1'b0}}, col_in_1273};
assign u_ca_in_1274 = {{7{1'b0}}, col_in_1274};
assign u_ca_in_1275 = {{7{1'b0}}, col_in_1275};
assign u_ca_in_1276 = {{7{1'b0}}, col_in_1276};
assign u_ca_in_1277 = {{7{1'b0}}, col_in_1277};
assign u_ca_in_1278 = {{7{1'b0}}, col_in_1278};
assign u_ca_in_1279 = {{7{1'b0}}, col_in_1279};

//---------------------------------------------------------


compressor_243_72 u_ca_243_72_0(.d_in(u_ca_in_0), .d_out(u_ca_out_0));
compressor_243_72 u_ca_243_72_1(.d_in(u_ca_in_1), .d_out(u_ca_out_1));
compressor_243_72 u_ca_243_72_2(.d_in(u_ca_in_2), .d_out(u_ca_out_2));
compressor_243_72 u_ca_243_72_3(.d_in(u_ca_in_3), .d_out(u_ca_out_3));
compressor_243_72 u_ca_243_72_4(.d_in(u_ca_in_4), .d_out(u_ca_out_4));
compressor_243_72 u_ca_243_72_5(.d_in(u_ca_in_5), .d_out(u_ca_out_5));
compressor_243_72 u_ca_243_72_6(.d_in(u_ca_in_6), .d_out(u_ca_out_6));
compressor_243_72 u_ca_243_72_7(.d_in(u_ca_in_7), .d_out(u_ca_out_7));
compressor_243_72 u_ca_243_72_8(.d_in(u_ca_in_8), .d_out(u_ca_out_8));
compressor_243_72 u_ca_243_72_9(.d_in(u_ca_in_9), .d_out(u_ca_out_9));
compressor_243_72 u_ca_243_72_10(.d_in(u_ca_in_10), .d_out(u_ca_out_10));
compressor_243_72 u_ca_243_72_11(.d_in(u_ca_in_11), .d_out(u_ca_out_11));
compressor_243_72 u_ca_243_72_12(.d_in(u_ca_in_12), .d_out(u_ca_out_12));
compressor_243_72 u_ca_243_72_13(.d_in(u_ca_in_13), .d_out(u_ca_out_13));
compressor_243_72 u_ca_243_72_14(.d_in(u_ca_in_14), .d_out(u_ca_out_14));
compressor_243_72 u_ca_243_72_15(.d_in(u_ca_in_15), .d_out(u_ca_out_15));
compressor_243_72 u_ca_243_72_16(.d_in(u_ca_in_16), .d_out(u_ca_out_16));
compressor_243_72 u_ca_243_72_17(.d_in(u_ca_in_17), .d_out(u_ca_out_17));
compressor_243_72 u_ca_243_72_18(.d_in(u_ca_in_18), .d_out(u_ca_out_18));
compressor_243_72 u_ca_243_72_19(.d_in(u_ca_in_19), .d_out(u_ca_out_19));
compressor_243_72 u_ca_243_72_20(.d_in(u_ca_in_20), .d_out(u_ca_out_20));
compressor_243_72 u_ca_243_72_21(.d_in(u_ca_in_21), .d_out(u_ca_out_21));
compressor_243_72 u_ca_243_72_22(.d_in(u_ca_in_22), .d_out(u_ca_out_22));
compressor_243_72 u_ca_243_72_23(.d_in(u_ca_in_23), .d_out(u_ca_out_23));
compressor_243_72 u_ca_243_72_24(.d_in(u_ca_in_24), .d_out(u_ca_out_24));
compressor_243_72 u_ca_243_72_25(.d_in(u_ca_in_25), .d_out(u_ca_out_25));
compressor_243_72 u_ca_243_72_26(.d_in(u_ca_in_26), .d_out(u_ca_out_26));
compressor_243_72 u_ca_243_72_27(.d_in(u_ca_in_27), .d_out(u_ca_out_27));
compressor_243_72 u_ca_243_72_28(.d_in(u_ca_in_28), .d_out(u_ca_out_28));
compressor_243_72 u_ca_243_72_29(.d_in(u_ca_in_29), .d_out(u_ca_out_29));
compressor_243_72 u_ca_243_72_30(.d_in(u_ca_in_30), .d_out(u_ca_out_30));
compressor_243_72 u_ca_243_72_31(.d_in(u_ca_in_31), .d_out(u_ca_out_31));
compressor_243_72 u_ca_243_72_32(.d_in(u_ca_in_32), .d_out(u_ca_out_32));
compressor_243_72 u_ca_243_72_33(.d_in(u_ca_in_33), .d_out(u_ca_out_33));
compressor_243_72 u_ca_243_72_34(.d_in(u_ca_in_34), .d_out(u_ca_out_34));
compressor_243_72 u_ca_243_72_35(.d_in(u_ca_in_35), .d_out(u_ca_out_35));
compressor_243_72 u_ca_243_72_36(.d_in(u_ca_in_36), .d_out(u_ca_out_36));
compressor_243_72 u_ca_243_72_37(.d_in(u_ca_in_37), .d_out(u_ca_out_37));
compressor_243_72 u_ca_243_72_38(.d_in(u_ca_in_38), .d_out(u_ca_out_38));
compressor_243_72 u_ca_243_72_39(.d_in(u_ca_in_39), .d_out(u_ca_out_39));
compressor_243_72 u_ca_243_72_40(.d_in(u_ca_in_40), .d_out(u_ca_out_40));
compressor_243_72 u_ca_243_72_41(.d_in(u_ca_in_41), .d_out(u_ca_out_41));
compressor_243_72 u_ca_243_72_42(.d_in(u_ca_in_42), .d_out(u_ca_out_42));
compressor_243_72 u_ca_243_72_43(.d_in(u_ca_in_43), .d_out(u_ca_out_43));
compressor_243_72 u_ca_243_72_44(.d_in(u_ca_in_44), .d_out(u_ca_out_44));
compressor_243_72 u_ca_243_72_45(.d_in(u_ca_in_45), .d_out(u_ca_out_45));
compressor_243_72 u_ca_243_72_46(.d_in(u_ca_in_46), .d_out(u_ca_out_46));
compressor_243_72 u_ca_243_72_47(.d_in(u_ca_in_47), .d_out(u_ca_out_47));
compressor_243_72 u_ca_243_72_48(.d_in(u_ca_in_48), .d_out(u_ca_out_48));
compressor_243_72 u_ca_243_72_49(.d_in(u_ca_in_49), .d_out(u_ca_out_49));
compressor_243_72 u_ca_243_72_50(.d_in(u_ca_in_50), .d_out(u_ca_out_50));
compressor_243_72 u_ca_243_72_51(.d_in(u_ca_in_51), .d_out(u_ca_out_51));
compressor_243_72 u_ca_243_72_52(.d_in(u_ca_in_52), .d_out(u_ca_out_52));
compressor_243_72 u_ca_243_72_53(.d_in(u_ca_in_53), .d_out(u_ca_out_53));
compressor_243_72 u_ca_243_72_54(.d_in(u_ca_in_54), .d_out(u_ca_out_54));
compressor_243_72 u_ca_243_72_55(.d_in(u_ca_in_55), .d_out(u_ca_out_55));
compressor_243_72 u_ca_243_72_56(.d_in(u_ca_in_56), .d_out(u_ca_out_56));
compressor_243_72 u_ca_243_72_57(.d_in(u_ca_in_57), .d_out(u_ca_out_57));
compressor_243_72 u_ca_243_72_58(.d_in(u_ca_in_58), .d_out(u_ca_out_58));
compressor_243_72 u_ca_243_72_59(.d_in(u_ca_in_59), .d_out(u_ca_out_59));
compressor_243_72 u_ca_243_72_60(.d_in(u_ca_in_60), .d_out(u_ca_out_60));
compressor_243_72 u_ca_243_72_61(.d_in(u_ca_in_61), .d_out(u_ca_out_61));
compressor_243_72 u_ca_243_72_62(.d_in(u_ca_in_62), .d_out(u_ca_out_62));
compressor_243_72 u_ca_243_72_63(.d_in(u_ca_in_63), .d_out(u_ca_out_63));
compressor_243_72 u_ca_243_72_64(.d_in(u_ca_in_64), .d_out(u_ca_out_64));
compressor_243_72 u_ca_243_72_65(.d_in(u_ca_in_65), .d_out(u_ca_out_65));
compressor_243_72 u_ca_243_72_66(.d_in(u_ca_in_66), .d_out(u_ca_out_66));
compressor_243_72 u_ca_243_72_67(.d_in(u_ca_in_67), .d_out(u_ca_out_67));
compressor_243_72 u_ca_243_72_68(.d_in(u_ca_in_68), .d_out(u_ca_out_68));
compressor_243_72 u_ca_243_72_69(.d_in(u_ca_in_69), .d_out(u_ca_out_69));
compressor_243_72 u_ca_243_72_70(.d_in(u_ca_in_70), .d_out(u_ca_out_70));
compressor_243_72 u_ca_243_72_71(.d_in(u_ca_in_71), .d_out(u_ca_out_71));
compressor_243_72 u_ca_243_72_72(.d_in(u_ca_in_72), .d_out(u_ca_out_72));
compressor_243_72 u_ca_243_72_73(.d_in(u_ca_in_73), .d_out(u_ca_out_73));
compressor_243_72 u_ca_243_72_74(.d_in(u_ca_in_74), .d_out(u_ca_out_74));
compressor_243_72 u_ca_243_72_75(.d_in(u_ca_in_75), .d_out(u_ca_out_75));
compressor_243_72 u_ca_243_72_76(.d_in(u_ca_in_76), .d_out(u_ca_out_76));
compressor_243_72 u_ca_243_72_77(.d_in(u_ca_in_77), .d_out(u_ca_out_77));
compressor_243_72 u_ca_243_72_78(.d_in(u_ca_in_78), .d_out(u_ca_out_78));
compressor_243_72 u_ca_243_72_79(.d_in(u_ca_in_79), .d_out(u_ca_out_79));
compressor_243_72 u_ca_243_72_80(.d_in(u_ca_in_80), .d_out(u_ca_out_80));
compressor_243_72 u_ca_243_72_81(.d_in(u_ca_in_81), .d_out(u_ca_out_81));
compressor_243_72 u_ca_243_72_82(.d_in(u_ca_in_82), .d_out(u_ca_out_82));
compressor_243_72 u_ca_243_72_83(.d_in(u_ca_in_83), .d_out(u_ca_out_83));
compressor_243_72 u_ca_243_72_84(.d_in(u_ca_in_84), .d_out(u_ca_out_84));
compressor_243_72 u_ca_243_72_85(.d_in(u_ca_in_85), .d_out(u_ca_out_85));
compressor_243_72 u_ca_243_72_86(.d_in(u_ca_in_86), .d_out(u_ca_out_86));
compressor_243_72 u_ca_243_72_87(.d_in(u_ca_in_87), .d_out(u_ca_out_87));
compressor_243_72 u_ca_243_72_88(.d_in(u_ca_in_88), .d_out(u_ca_out_88));
compressor_243_72 u_ca_243_72_89(.d_in(u_ca_in_89), .d_out(u_ca_out_89));
compressor_243_72 u_ca_243_72_90(.d_in(u_ca_in_90), .d_out(u_ca_out_90));
compressor_243_72 u_ca_243_72_91(.d_in(u_ca_in_91), .d_out(u_ca_out_91));
compressor_243_72 u_ca_243_72_92(.d_in(u_ca_in_92), .d_out(u_ca_out_92));
compressor_243_72 u_ca_243_72_93(.d_in(u_ca_in_93), .d_out(u_ca_out_93));
compressor_243_72 u_ca_243_72_94(.d_in(u_ca_in_94), .d_out(u_ca_out_94));
compressor_243_72 u_ca_243_72_95(.d_in(u_ca_in_95), .d_out(u_ca_out_95));
compressor_243_72 u_ca_243_72_96(.d_in(u_ca_in_96), .d_out(u_ca_out_96));
compressor_243_72 u_ca_243_72_97(.d_in(u_ca_in_97), .d_out(u_ca_out_97));
compressor_243_72 u_ca_243_72_98(.d_in(u_ca_in_98), .d_out(u_ca_out_98));
compressor_243_72 u_ca_243_72_99(.d_in(u_ca_in_99), .d_out(u_ca_out_99));
compressor_243_72 u_ca_243_72_100(.d_in(u_ca_in_100), .d_out(u_ca_out_100));
compressor_243_72 u_ca_243_72_101(.d_in(u_ca_in_101), .d_out(u_ca_out_101));
compressor_243_72 u_ca_243_72_102(.d_in(u_ca_in_102), .d_out(u_ca_out_102));
compressor_243_72 u_ca_243_72_103(.d_in(u_ca_in_103), .d_out(u_ca_out_103));
compressor_243_72 u_ca_243_72_104(.d_in(u_ca_in_104), .d_out(u_ca_out_104));
compressor_243_72 u_ca_243_72_105(.d_in(u_ca_in_105), .d_out(u_ca_out_105));
compressor_243_72 u_ca_243_72_106(.d_in(u_ca_in_106), .d_out(u_ca_out_106));
compressor_243_72 u_ca_243_72_107(.d_in(u_ca_in_107), .d_out(u_ca_out_107));
compressor_243_72 u_ca_243_72_108(.d_in(u_ca_in_108), .d_out(u_ca_out_108));
compressor_243_72 u_ca_243_72_109(.d_in(u_ca_in_109), .d_out(u_ca_out_109));
compressor_243_72 u_ca_243_72_110(.d_in(u_ca_in_110), .d_out(u_ca_out_110));
compressor_243_72 u_ca_243_72_111(.d_in(u_ca_in_111), .d_out(u_ca_out_111));
compressor_243_72 u_ca_243_72_112(.d_in(u_ca_in_112), .d_out(u_ca_out_112));
compressor_243_72 u_ca_243_72_113(.d_in(u_ca_in_113), .d_out(u_ca_out_113));
compressor_243_72 u_ca_243_72_114(.d_in(u_ca_in_114), .d_out(u_ca_out_114));
compressor_243_72 u_ca_243_72_115(.d_in(u_ca_in_115), .d_out(u_ca_out_115));
compressor_243_72 u_ca_243_72_116(.d_in(u_ca_in_116), .d_out(u_ca_out_116));
compressor_243_72 u_ca_243_72_117(.d_in(u_ca_in_117), .d_out(u_ca_out_117));
compressor_243_72 u_ca_243_72_118(.d_in(u_ca_in_118), .d_out(u_ca_out_118));
compressor_243_72 u_ca_243_72_119(.d_in(u_ca_in_119), .d_out(u_ca_out_119));
compressor_243_72 u_ca_243_72_120(.d_in(u_ca_in_120), .d_out(u_ca_out_120));
compressor_243_72 u_ca_243_72_121(.d_in(u_ca_in_121), .d_out(u_ca_out_121));
compressor_243_72 u_ca_243_72_122(.d_in(u_ca_in_122), .d_out(u_ca_out_122));
compressor_243_72 u_ca_243_72_123(.d_in(u_ca_in_123), .d_out(u_ca_out_123));
compressor_243_72 u_ca_243_72_124(.d_in(u_ca_in_124), .d_out(u_ca_out_124));
compressor_243_72 u_ca_243_72_125(.d_in(u_ca_in_125), .d_out(u_ca_out_125));
compressor_243_72 u_ca_243_72_126(.d_in(u_ca_in_126), .d_out(u_ca_out_126));
compressor_243_72 u_ca_243_72_127(.d_in(u_ca_in_127), .d_out(u_ca_out_127));
compressor_243_72 u_ca_243_72_128(.d_in(u_ca_in_128), .d_out(u_ca_out_128));
compressor_243_72 u_ca_243_72_129(.d_in(u_ca_in_129), .d_out(u_ca_out_129));
compressor_243_72 u_ca_243_72_130(.d_in(u_ca_in_130), .d_out(u_ca_out_130));
compressor_243_72 u_ca_243_72_131(.d_in(u_ca_in_131), .d_out(u_ca_out_131));
compressor_243_72 u_ca_243_72_132(.d_in(u_ca_in_132), .d_out(u_ca_out_132));
compressor_243_72 u_ca_243_72_133(.d_in(u_ca_in_133), .d_out(u_ca_out_133));
compressor_243_72 u_ca_243_72_134(.d_in(u_ca_in_134), .d_out(u_ca_out_134));
compressor_243_72 u_ca_243_72_135(.d_in(u_ca_in_135), .d_out(u_ca_out_135));
compressor_243_72 u_ca_243_72_136(.d_in(u_ca_in_136), .d_out(u_ca_out_136));
compressor_243_72 u_ca_243_72_137(.d_in(u_ca_in_137), .d_out(u_ca_out_137));
compressor_243_72 u_ca_243_72_138(.d_in(u_ca_in_138), .d_out(u_ca_out_138));
compressor_243_72 u_ca_243_72_139(.d_in(u_ca_in_139), .d_out(u_ca_out_139));
compressor_243_72 u_ca_243_72_140(.d_in(u_ca_in_140), .d_out(u_ca_out_140));
compressor_243_72 u_ca_243_72_141(.d_in(u_ca_in_141), .d_out(u_ca_out_141));
compressor_243_72 u_ca_243_72_142(.d_in(u_ca_in_142), .d_out(u_ca_out_142));
compressor_243_72 u_ca_243_72_143(.d_in(u_ca_in_143), .d_out(u_ca_out_143));
compressor_243_72 u_ca_243_72_144(.d_in(u_ca_in_144), .d_out(u_ca_out_144));
compressor_243_72 u_ca_243_72_145(.d_in(u_ca_in_145), .d_out(u_ca_out_145));
compressor_243_72 u_ca_243_72_146(.d_in(u_ca_in_146), .d_out(u_ca_out_146));
compressor_243_72 u_ca_243_72_147(.d_in(u_ca_in_147), .d_out(u_ca_out_147));
compressor_243_72 u_ca_243_72_148(.d_in(u_ca_in_148), .d_out(u_ca_out_148));
compressor_243_72 u_ca_243_72_149(.d_in(u_ca_in_149), .d_out(u_ca_out_149));
compressor_243_72 u_ca_243_72_150(.d_in(u_ca_in_150), .d_out(u_ca_out_150));
compressor_243_72 u_ca_243_72_151(.d_in(u_ca_in_151), .d_out(u_ca_out_151));
compressor_243_72 u_ca_243_72_152(.d_in(u_ca_in_152), .d_out(u_ca_out_152));
compressor_243_72 u_ca_243_72_153(.d_in(u_ca_in_153), .d_out(u_ca_out_153));
compressor_243_72 u_ca_243_72_154(.d_in(u_ca_in_154), .d_out(u_ca_out_154));
compressor_243_72 u_ca_243_72_155(.d_in(u_ca_in_155), .d_out(u_ca_out_155));
compressor_243_72 u_ca_243_72_156(.d_in(u_ca_in_156), .d_out(u_ca_out_156));
compressor_243_72 u_ca_243_72_157(.d_in(u_ca_in_157), .d_out(u_ca_out_157));
compressor_243_72 u_ca_243_72_158(.d_in(u_ca_in_158), .d_out(u_ca_out_158));
compressor_243_72 u_ca_243_72_159(.d_in(u_ca_in_159), .d_out(u_ca_out_159));
compressor_243_72 u_ca_243_72_160(.d_in(u_ca_in_160), .d_out(u_ca_out_160));
compressor_243_72 u_ca_243_72_161(.d_in(u_ca_in_161), .d_out(u_ca_out_161));
compressor_243_72 u_ca_243_72_162(.d_in(u_ca_in_162), .d_out(u_ca_out_162));
compressor_243_72 u_ca_243_72_163(.d_in(u_ca_in_163), .d_out(u_ca_out_163));
compressor_243_72 u_ca_243_72_164(.d_in(u_ca_in_164), .d_out(u_ca_out_164));
compressor_243_72 u_ca_243_72_165(.d_in(u_ca_in_165), .d_out(u_ca_out_165));
compressor_243_72 u_ca_243_72_166(.d_in(u_ca_in_166), .d_out(u_ca_out_166));
compressor_243_72 u_ca_243_72_167(.d_in(u_ca_in_167), .d_out(u_ca_out_167));
compressor_243_72 u_ca_243_72_168(.d_in(u_ca_in_168), .d_out(u_ca_out_168));
compressor_243_72 u_ca_243_72_169(.d_in(u_ca_in_169), .d_out(u_ca_out_169));
compressor_243_72 u_ca_243_72_170(.d_in(u_ca_in_170), .d_out(u_ca_out_170));
compressor_243_72 u_ca_243_72_171(.d_in(u_ca_in_171), .d_out(u_ca_out_171));
compressor_243_72 u_ca_243_72_172(.d_in(u_ca_in_172), .d_out(u_ca_out_172));
compressor_243_72 u_ca_243_72_173(.d_in(u_ca_in_173), .d_out(u_ca_out_173));
compressor_243_72 u_ca_243_72_174(.d_in(u_ca_in_174), .d_out(u_ca_out_174));
compressor_243_72 u_ca_243_72_175(.d_in(u_ca_in_175), .d_out(u_ca_out_175));
compressor_243_72 u_ca_243_72_176(.d_in(u_ca_in_176), .d_out(u_ca_out_176));
compressor_243_72 u_ca_243_72_177(.d_in(u_ca_in_177), .d_out(u_ca_out_177));
compressor_243_72 u_ca_243_72_178(.d_in(u_ca_in_178), .d_out(u_ca_out_178));
compressor_243_72 u_ca_243_72_179(.d_in(u_ca_in_179), .d_out(u_ca_out_179));
compressor_243_72 u_ca_243_72_180(.d_in(u_ca_in_180), .d_out(u_ca_out_180));
compressor_243_72 u_ca_243_72_181(.d_in(u_ca_in_181), .d_out(u_ca_out_181));
compressor_243_72 u_ca_243_72_182(.d_in(u_ca_in_182), .d_out(u_ca_out_182));
compressor_243_72 u_ca_243_72_183(.d_in(u_ca_in_183), .d_out(u_ca_out_183));
compressor_243_72 u_ca_243_72_184(.d_in(u_ca_in_184), .d_out(u_ca_out_184));
compressor_243_72 u_ca_243_72_185(.d_in(u_ca_in_185), .d_out(u_ca_out_185));
compressor_243_72 u_ca_243_72_186(.d_in(u_ca_in_186), .d_out(u_ca_out_186));
compressor_243_72 u_ca_243_72_187(.d_in(u_ca_in_187), .d_out(u_ca_out_187));
compressor_243_72 u_ca_243_72_188(.d_in(u_ca_in_188), .d_out(u_ca_out_188));
compressor_243_72 u_ca_243_72_189(.d_in(u_ca_in_189), .d_out(u_ca_out_189));
compressor_243_72 u_ca_243_72_190(.d_in(u_ca_in_190), .d_out(u_ca_out_190));
compressor_243_72 u_ca_243_72_191(.d_in(u_ca_in_191), .d_out(u_ca_out_191));
compressor_243_72 u_ca_243_72_192(.d_in(u_ca_in_192), .d_out(u_ca_out_192));
compressor_243_72 u_ca_243_72_193(.d_in(u_ca_in_193), .d_out(u_ca_out_193));
compressor_243_72 u_ca_243_72_194(.d_in(u_ca_in_194), .d_out(u_ca_out_194));
compressor_243_72 u_ca_243_72_195(.d_in(u_ca_in_195), .d_out(u_ca_out_195));
compressor_243_72 u_ca_243_72_196(.d_in(u_ca_in_196), .d_out(u_ca_out_196));
compressor_243_72 u_ca_243_72_197(.d_in(u_ca_in_197), .d_out(u_ca_out_197));
compressor_243_72 u_ca_243_72_198(.d_in(u_ca_in_198), .d_out(u_ca_out_198));
compressor_243_72 u_ca_243_72_199(.d_in(u_ca_in_199), .d_out(u_ca_out_199));
compressor_243_72 u_ca_243_72_200(.d_in(u_ca_in_200), .d_out(u_ca_out_200));
compressor_243_72 u_ca_243_72_201(.d_in(u_ca_in_201), .d_out(u_ca_out_201));
compressor_243_72 u_ca_243_72_202(.d_in(u_ca_in_202), .d_out(u_ca_out_202));
compressor_243_72 u_ca_243_72_203(.d_in(u_ca_in_203), .d_out(u_ca_out_203));
compressor_243_72 u_ca_243_72_204(.d_in(u_ca_in_204), .d_out(u_ca_out_204));
compressor_243_72 u_ca_243_72_205(.d_in(u_ca_in_205), .d_out(u_ca_out_205));
compressor_243_72 u_ca_243_72_206(.d_in(u_ca_in_206), .d_out(u_ca_out_206));
compressor_243_72 u_ca_243_72_207(.d_in(u_ca_in_207), .d_out(u_ca_out_207));
compressor_243_72 u_ca_243_72_208(.d_in(u_ca_in_208), .d_out(u_ca_out_208));
compressor_243_72 u_ca_243_72_209(.d_in(u_ca_in_209), .d_out(u_ca_out_209));
compressor_243_72 u_ca_243_72_210(.d_in(u_ca_in_210), .d_out(u_ca_out_210));
compressor_243_72 u_ca_243_72_211(.d_in(u_ca_in_211), .d_out(u_ca_out_211));
compressor_243_72 u_ca_243_72_212(.d_in(u_ca_in_212), .d_out(u_ca_out_212));
compressor_243_72 u_ca_243_72_213(.d_in(u_ca_in_213), .d_out(u_ca_out_213));
compressor_243_72 u_ca_243_72_214(.d_in(u_ca_in_214), .d_out(u_ca_out_214));
compressor_243_72 u_ca_243_72_215(.d_in(u_ca_in_215), .d_out(u_ca_out_215));
compressor_243_72 u_ca_243_72_216(.d_in(u_ca_in_216), .d_out(u_ca_out_216));
compressor_243_72 u_ca_243_72_217(.d_in(u_ca_in_217), .d_out(u_ca_out_217));
compressor_243_72 u_ca_243_72_218(.d_in(u_ca_in_218), .d_out(u_ca_out_218));
compressor_243_72 u_ca_243_72_219(.d_in(u_ca_in_219), .d_out(u_ca_out_219));
compressor_243_72 u_ca_243_72_220(.d_in(u_ca_in_220), .d_out(u_ca_out_220));
compressor_243_72 u_ca_243_72_221(.d_in(u_ca_in_221), .d_out(u_ca_out_221));
compressor_243_72 u_ca_243_72_222(.d_in(u_ca_in_222), .d_out(u_ca_out_222));
compressor_243_72 u_ca_243_72_223(.d_in(u_ca_in_223), .d_out(u_ca_out_223));
compressor_243_72 u_ca_243_72_224(.d_in(u_ca_in_224), .d_out(u_ca_out_224));
compressor_243_72 u_ca_243_72_225(.d_in(u_ca_in_225), .d_out(u_ca_out_225));
compressor_243_72 u_ca_243_72_226(.d_in(u_ca_in_226), .d_out(u_ca_out_226));
compressor_243_72 u_ca_243_72_227(.d_in(u_ca_in_227), .d_out(u_ca_out_227));
compressor_243_72 u_ca_243_72_228(.d_in(u_ca_in_228), .d_out(u_ca_out_228));
compressor_243_72 u_ca_243_72_229(.d_in(u_ca_in_229), .d_out(u_ca_out_229));
compressor_243_72 u_ca_243_72_230(.d_in(u_ca_in_230), .d_out(u_ca_out_230));
compressor_243_72 u_ca_243_72_231(.d_in(u_ca_in_231), .d_out(u_ca_out_231));
compressor_243_72 u_ca_243_72_232(.d_in(u_ca_in_232), .d_out(u_ca_out_232));
compressor_243_72 u_ca_243_72_233(.d_in(u_ca_in_233), .d_out(u_ca_out_233));
compressor_243_72 u_ca_243_72_234(.d_in(u_ca_in_234), .d_out(u_ca_out_234));
compressor_243_72 u_ca_243_72_235(.d_in(u_ca_in_235), .d_out(u_ca_out_235));
compressor_243_72 u_ca_243_72_236(.d_in(u_ca_in_236), .d_out(u_ca_out_236));
compressor_243_72 u_ca_243_72_237(.d_in(u_ca_in_237), .d_out(u_ca_out_237));
compressor_243_72 u_ca_243_72_238(.d_in(u_ca_in_238), .d_out(u_ca_out_238));
compressor_243_72 u_ca_243_72_239(.d_in(u_ca_in_239), .d_out(u_ca_out_239));
compressor_243_72 u_ca_243_72_240(.d_in(u_ca_in_240), .d_out(u_ca_out_240));
compressor_243_72 u_ca_243_72_241(.d_in(u_ca_in_241), .d_out(u_ca_out_241));
compressor_243_72 u_ca_243_72_242(.d_in(u_ca_in_242), .d_out(u_ca_out_242));
compressor_243_72 u_ca_243_72_243(.d_in(u_ca_in_243), .d_out(u_ca_out_243));
compressor_243_72 u_ca_243_72_244(.d_in(u_ca_in_244), .d_out(u_ca_out_244));
compressor_243_72 u_ca_243_72_245(.d_in(u_ca_in_245), .d_out(u_ca_out_245));
compressor_243_72 u_ca_243_72_246(.d_in(u_ca_in_246), .d_out(u_ca_out_246));
compressor_243_72 u_ca_243_72_247(.d_in(u_ca_in_247), .d_out(u_ca_out_247));
compressor_243_72 u_ca_243_72_248(.d_in(u_ca_in_248), .d_out(u_ca_out_248));
compressor_243_72 u_ca_243_72_249(.d_in(u_ca_in_249), .d_out(u_ca_out_249));
compressor_243_72 u_ca_243_72_250(.d_in(u_ca_in_250), .d_out(u_ca_out_250));
compressor_243_72 u_ca_243_72_251(.d_in(u_ca_in_251), .d_out(u_ca_out_251));
compressor_243_72 u_ca_243_72_252(.d_in(u_ca_in_252), .d_out(u_ca_out_252));
compressor_243_72 u_ca_243_72_253(.d_in(u_ca_in_253), .d_out(u_ca_out_253));
compressor_243_72 u_ca_243_72_254(.d_in(u_ca_in_254), .d_out(u_ca_out_254));
compressor_243_72 u_ca_243_72_255(.d_in(u_ca_in_255), .d_out(u_ca_out_255));
compressor_243_72 u_ca_243_72_256(.d_in(u_ca_in_256), .d_out(u_ca_out_256));
compressor_243_72 u_ca_243_72_257(.d_in(u_ca_in_257), .d_out(u_ca_out_257));
compressor_243_72 u_ca_243_72_258(.d_in(u_ca_in_258), .d_out(u_ca_out_258));
compressor_243_72 u_ca_243_72_259(.d_in(u_ca_in_259), .d_out(u_ca_out_259));
compressor_243_72 u_ca_243_72_260(.d_in(u_ca_in_260), .d_out(u_ca_out_260));
compressor_243_72 u_ca_243_72_261(.d_in(u_ca_in_261), .d_out(u_ca_out_261));
compressor_243_72 u_ca_243_72_262(.d_in(u_ca_in_262), .d_out(u_ca_out_262));
compressor_243_72 u_ca_243_72_263(.d_in(u_ca_in_263), .d_out(u_ca_out_263));
compressor_243_72 u_ca_243_72_264(.d_in(u_ca_in_264), .d_out(u_ca_out_264));
compressor_243_72 u_ca_243_72_265(.d_in(u_ca_in_265), .d_out(u_ca_out_265));
compressor_243_72 u_ca_243_72_266(.d_in(u_ca_in_266), .d_out(u_ca_out_266));
compressor_243_72 u_ca_243_72_267(.d_in(u_ca_in_267), .d_out(u_ca_out_267));
compressor_243_72 u_ca_243_72_268(.d_in(u_ca_in_268), .d_out(u_ca_out_268));
compressor_243_72 u_ca_243_72_269(.d_in(u_ca_in_269), .d_out(u_ca_out_269));
compressor_243_72 u_ca_243_72_270(.d_in(u_ca_in_270), .d_out(u_ca_out_270));
compressor_243_72 u_ca_243_72_271(.d_in(u_ca_in_271), .d_out(u_ca_out_271));
compressor_243_72 u_ca_243_72_272(.d_in(u_ca_in_272), .d_out(u_ca_out_272));
compressor_243_72 u_ca_243_72_273(.d_in(u_ca_in_273), .d_out(u_ca_out_273));
compressor_243_72 u_ca_243_72_274(.d_in(u_ca_in_274), .d_out(u_ca_out_274));
compressor_243_72 u_ca_243_72_275(.d_in(u_ca_in_275), .d_out(u_ca_out_275));
compressor_243_72 u_ca_243_72_276(.d_in(u_ca_in_276), .d_out(u_ca_out_276));
compressor_243_72 u_ca_243_72_277(.d_in(u_ca_in_277), .d_out(u_ca_out_277));
compressor_243_72 u_ca_243_72_278(.d_in(u_ca_in_278), .d_out(u_ca_out_278));
compressor_243_72 u_ca_243_72_279(.d_in(u_ca_in_279), .d_out(u_ca_out_279));
compressor_243_72 u_ca_243_72_280(.d_in(u_ca_in_280), .d_out(u_ca_out_280));
compressor_243_72 u_ca_243_72_281(.d_in(u_ca_in_281), .d_out(u_ca_out_281));
compressor_243_72 u_ca_243_72_282(.d_in(u_ca_in_282), .d_out(u_ca_out_282));
compressor_243_72 u_ca_243_72_283(.d_in(u_ca_in_283), .d_out(u_ca_out_283));
compressor_243_72 u_ca_243_72_284(.d_in(u_ca_in_284), .d_out(u_ca_out_284));
compressor_243_72 u_ca_243_72_285(.d_in(u_ca_in_285), .d_out(u_ca_out_285));
compressor_243_72 u_ca_243_72_286(.d_in(u_ca_in_286), .d_out(u_ca_out_286));
compressor_243_72 u_ca_243_72_287(.d_in(u_ca_in_287), .d_out(u_ca_out_287));
compressor_243_72 u_ca_243_72_288(.d_in(u_ca_in_288), .d_out(u_ca_out_288));
compressor_243_72 u_ca_243_72_289(.d_in(u_ca_in_289), .d_out(u_ca_out_289));
compressor_243_72 u_ca_243_72_290(.d_in(u_ca_in_290), .d_out(u_ca_out_290));
compressor_243_72 u_ca_243_72_291(.d_in(u_ca_in_291), .d_out(u_ca_out_291));
compressor_243_72 u_ca_243_72_292(.d_in(u_ca_in_292), .d_out(u_ca_out_292));
compressor_243_72 u_ca_243_72_293(.d_in(u_ca_in_293), .d_out(u_ca_out_293));
compressor_243_72 u_ca_243_72_294(.d_in(u_ca_in_294), .d_out(u_ca_out_294));
compressor_243_72 u_ca_243_72_295(.d_in(u_ca_in_295), .d_out(u_ca_out_295));
compressor_243_72 u_ca_243_72_296(.d_in(u_ca_in_296), .d_out(u_ca_out_296));
compressor_243_72 u_ca_243_72_297(.d_in(u_ca_in_297), .d_out(u_ca_out_297));
compressor_243_72 u_ca_243_72_298(.d_in(u_ca_in_298), .d_out(u_ca_out_298));
compressor_243_72 u_ca_243_72_299(.d_in(u_ca_in_299), .d_out(u_ca_out_299));
compressor_243_72 u_ca_243_72_300(.d_in(u_ca_in_300), .d_out(u_ca_out_300));
compressor_243_72 u_ca_243_72_301(.d_in(u_ca_in_301), .d_out(u_ca_out_301));
compressor_243_72 u_ca_243_72_302(.d_in(u_ca_in_302), .d_out(u_ca_out_302));
compressor_243_72 u_ca_243_72_303(.d_in(u_ca_in_303), .d_out(u_ca_out_303));
compressor_243_72 u_ca_243_72_304(.d_in(u_ca_in_304), .d_out(u_ca_out_304));
compressor_243_72 u_ca_243_72_305(.d_in(u_ca_in_305), .d_out(u_ca_out_305));
compressor_243_72 u_ca_243_72_306(.d_in(u_ca_in_306), .d_out(u_ca_out_306));
compressor_243_72 u_ca_243_72_307(.d_in(u_ca_in_307), .d_out(u_ca_out_307));
compressor_243_72 u_ca_243_72_308(.d_in(u_ca_in_308), .d_out(u_ca_out_308));
compressor_243_72 u_ca_243_72_309(.d_in(u_ca_in_309), .d_out(u_ca_out_309));
compressor_243_72 u_ca_243_72_310(.d_in(u_ca_in_310), .d_out(u_ca_out_310));
compressor_243_72 u_ca_243_72_311(.d_in(u_ca_in_311), .d_out(u_ca_out_311));
compressor_243_72 u_ca_243_72_312(.d_in(u_ca_in_312), .d_out(u_ca_out_312));
compressor_243_72 u_ca_243_72_313(.d_in(u_ca_in_313), .d_out(u_ca_out_313));
compressor_243_72 u_ca_243_72_314(.d_in(u_ca_in_314), .d_out(u_ca_out_314));
compressor_243_72 u_ca_243_72_315(.d_in(u_ca_in_315), .d_out(u_ca_out_315));
compressor_243_72 u_ca_243_72_316(.d_in(u_ca_in_316), .d_out(u_ca_out_316));
compressor_243_72 u_ca_243_72_317(.d_in(u_ca_in_317), .d_out(u_ca_out_317));
compressor_243_72 u_ca_243_72_318(.d_in(u_ca_in_318), .d_out(u_ca_out_318));
compressor_243_72 u_ca_243_72_319(.d_in(u_ca_in_319), .d_out(u_ca_out_319));
compressor_243_72 u_ca_243_72_320(.d_in(u_ca_in_320), .d_out(u_ca_out_320));
compressor_243_72 u_ca_243_72_321(.d_in(u_ca_in_321), .d_out(u_ca_out_321));
compressor_243_72 u_ca_243_72_322(.d_in(u_ca_in_322), .d_out(u_ca_out_322));
compressor_243_72 u_ca_243_72_323(.d_in(u_ca_in_323), .d_out(u_ca_out_323));
compressor_243_72 u_ca_243_72_324(.d_in(u_ca_in_324), .d_out(u_ca_out_324));
compressor_243_72 u_ca_243_72_325(.d_in(u_ca_in_325), .d_out(u_ca_out_325));
compressor_243_72 u_ca_243_72_326(.d_in(u_ca_in_326), .d_out(u_ca_out_326));
compressor_243_72 u_ca_243_72_327(.d_in(u_ca_in_327), .d_out(u_ca_out_327));
compressor_243_72 u_ca_243_72_328(.d_in(u_ca_in_328), .d_out(u_ca_out_328));
compressor_243_72 u_ca_243_72_329(.d_in(u_ca_in_329), .d_out(u_ca_out_329));
compressor_243_72 u_ca_243_72_330(.d_in(u_ca_in_330), .d_out(u_ca_out_330));
compressor_243_72 u_ca_243_72_331(.d_in(u_ca_in_331), .d_out(u_ca_out_331));
compressor_243_72 u_ca_243_72_332(.d_in(u_ca_in_332), .d_out(u_ca_out_332));
compressor_243_72 u_ca_243_72_333(.d_in(u_ca_in_333), .d_out(u_ca_out_333));
compressor_243_72 u_ca_243_72_334(.d_in(u_ca_in_334), .d_out(u_ca_out_334));
compressor_243_72 u_ca_243_72_335(.d_in(u_ca_in_335), .d_out(u_ca_out_335));
compressor_243_72 u_ca_243_72_336(.d_in(u_ca_in_336), .d_out(u_ca_out_336));
compressor_243_72 u_ca_243_72_337(.d_in(u_ca_in_337), .d_out(u_ca_out_337));
compressor_243_72 u_ca_243_72_338(.d_in(u_ca_in_338), .d_out(u_ca_out_338));
compressor_243_72 u_ca_243_72_339(.d_in(u_ca_in_339), .d_out(u_ca_out_339));
compressor_243_72 u_ca_243_72_340(.d_in(u_ca_in_340), .d_out(u_ca_out_340));
compressor_243_72 u_ca_243_72_341(.d_in(u_ca_in_341), .d_out(u_ca_out_341));
compressor_243_72 u_ca_243_72_342(.d_in(u_ca_in_342), .d_out(u_ca_out_342));
compressor_243_72 u_ca_243_72_343(.d_in(u_ca_in_343), .d_out(u_ca_out_343));
compressor_243_72 u_ca_243_72_344(.d_in(u_ca_in_344), .d_out(u_ca_out_344));
compressor_243_72 u_ca_243_72_345(.d_in(u_ca_in_345), .d_out(u_ca_out_345));
compressor_243_72 u_ca_243_72_346(.d_in(u_ca_in_346), .d_out(u_ca_out_346));
compressor_243_72 u_ca_243_72_347(.d_in(u_ca_in_347), .d_out(u_ca_out_347));
compressor_243_72 u_ca_243_72_348(.d_in(u_ca_in_348), .d_out(u_ca_out_348));
compressor_243_72 u_ca_243_72_349(.d_in(u_ca_in_349), .d_out(u_ca_out_349));
compressor_243_72 u_ca_243_72_350(.d_in(u_ca_in_350), .d_out(u_ca_out_350));
compressor_243_72 u_ca_243_72_351(.d_in(u_ca_in_351), .d_out(u_ca_out_351));
compressor_243_72 u_ca_243_72_352(.d_in(u_ca_in_352), .d_out(u_ca_out_352));
compressor_243_72 u_ca_243_72_353(.d_in(u_ca_in_353), .d_out(u_ca_out_353));
compressor_243_72 u_ca_243_72_354(.d_in(u_ca_in_354), .d_out(u_ca_out_354));
compressor_243_72 u_ca_243_72_355(.d_in(u_ca_in_355), .d_out(u_ca_out_355));
compressor_243_72 u_ca_243_72_356(.d_in(u_ca_in_356), .d_out(u_ca_out_356));
compressor_243_72 u_ca_243_72_357(.d_in(u_ca_in_357), .d_out(u_ca_out_357));
compressor_243_72 u_ca_243_72_358(.d_in(u_ca_in_358), .d_out(u_ca_out_358));
compressor_243_72 u_ca_243_72_359(.d_in(u_ca_in_359), .d_out(u_ca_out_359));
compressor_243_72 u_ca_243_72_360(.d_in(u_ca_in_360), .d_out(u_ca_out_360));
compressor_243_72 u_ca_243_72_361(.d_in(u_ca_in_361), .d_out(u_ca_out_361));
compressor_243_72 u_ca_243_72_362(.d_in(u_ca_in_362), .d_out(u_ca_out_362));
compressor_243_72 u_ca_243_72_363(.d_in(u_ca_in_363), .d_out(u_ca_out_363));
compressor_243_72 u_ca_243_72_364(.d_in(u_ca_in_364), .d_out(u_ca_out_364));
compressor_243_72 u_ca_243_72_365(.d_in(u_ca_in_365), .d_out(u_ca_out_365));
compressor_243_72 u_ca_243_72_366(.d_in(u_ca_in_366), .d_out(u_ca_out_366));
compressor_243_72 u_ca_243_72_367(.d_in(u_ca_in_367), .d_out(u_ca_out_367));
compressor_243_72 u_ca_243_72_368(.d_in(u_ca_in_368), .d_out(u_ca_out_368));
compressor_243_72 u_ca_243_72_369(.d_in(u_ca_in_369), .d_out(u_ca_out_369));
compressor_243_72 u_ca_243_72_370(.d_in(u_ca_in_370), .d_out(u_ca_out_370));
compressor_243_72 u_ca_243_72_371(.d_in(u_ca_in_371), .d_out(u_ca_out_371));
compressor_243_72 u_ca_243_72_372(.d_in(u_ca_in_372), .d_out(u_ca_out_372));
compressor_243_72 u_ca_243_72_373(.d_in(u_ca_in_373), .d_out(u_ca_out_373));
compressor_243_72 u_ca_243_72_374(.d_in(u_ca_in_374), .d_out(u_ca_out_374));
compressor_243_72 u_ca_243_72_375(.d_in(u_ca_in_375), .d_out(u_ca_out_375));
compressor_243_72 u_ca_243_72_376(.d_in(u_ca_in_376), .d_out(u_ca_out_376));
compressor_243_72 u_ca_243_72_377(.d_in(u_ca_in_377), .d_out(u_ca_out_377));
compressor_243_72 u_ca_243_72_378(.d_in(u_ca_in_378), .d_out(u_ca_out_378));
compressor_243_72 u_ca_243_72_379(.d_in(u_ca_in_379), .d_out(u_ca_out_379));
compressor_243_72 u_ca_243_72_380(.d_in(u_ca_in_380), .d_out(u_ca_out_380));
compressor_243_72 u_ca_243_72_381(.d_in(u_ca_in_381), .d_out(u_ca_out_381));
compressor_243_72 u_ca_243_72_382(.d_in(u_ca_in_382), .d_out(u_ca_out_382));
compressor_243_72 u_ca_243_72_383(.d_in(u_ca_in_383), .d_out(u_ca_out_383));
compressor_243_72 u_ca_243_72_384(.d_in(u_ca_in_384), .d_out(u_ca_out_384));
compressor_243_72 u_ca_243_72_385(.d_in(u_ca_in_385), .d_out(u_ca_out_385));
compressor_243_72 u_ca_243_72_386(.d_in(u_ca_in_386), .d_out(u_ca_out_386));
compressor_243_72 u_ca_243_72_387(.d_in(u_ca_in_387), .d_out(u_ca_out_387));
compressor_243_72 u_ca_243_72_388(.d_in(u_ca_in_388), .d_out(u_ca_out_388));
compressor_243_72 u_ca_243_72_389(.d_in(u_ca_in_389), .d_out(u_ca_out_389));
compressor_243_72 u_ca_243_72_390(.d_in(u_ca_in_390), .d_out(u_ca_out_390));
compressor_243_72 u_ca_243_72_391(.d_in(u_ca_in_391), .d_out(u_ca_out_391));
compressor_243_72 u_ca_243_72_392(.d_in(u_ca_in_392), .d_out(u_ca_out_392));
compressor_243_72 u_ca_243_72_393(.d_in(u_ca_in_393), .d_out(u_ca_out_393));
compressor_243_72 u_ca_243_72_394(.d_in(u_ca_in_394), .d_out(u_ca_out_394));
compressor_243_72 u_ca_243_72_395(.d_in(u_ca_in_395), .d_out(u_ca_out_395));
compressor_243_72 u_ca_243_72_396(.d_in(u_ca_in_396), .d_out(u_ca_out_396));
compressor_243_72 u_ca_243_72_397(.d_in(u_ca_in_397), .d_out(u_ca_out_397));
compressor_243_72 u_ca_243_72_398(.d_in(u_ca_in_398), .d_out(u_ca_out_398));
compressor_243_72 u_ca_243_72_399(.d_in(u_ca_in_399), .d_out(u_ca_out_399));
compressor_243_72 u_ca_243_72_400(.d_in(u_ca_in_400), .d_out(u_ca_out_400));
compressor_243_72 u_ca_243_72_401(.d_in(u_ca_in_401), .d_out(u_ca_out_401));
compressor_243_72 u_ca_243_72_402(.d_in(u_ca_in_402), .d_out(u_ca_out_402));
compressor_243_72 u_ca_243_72_403(.d_in(u_ca_in_403), .d_out(u_ca_out_403));
compressor_243_72 u_ca_243_72_404(.d_in(u_ca_in_404), .d_out(u_ca_out_404));
compressor_243_72 u_ca_243_72_405(.d_in(u_ca_in_405), .d_out(u_ca_out_405));
compressor_243_72 u_ca_243_72_406(.d_in(u_ca_in_406), .d_out(u_ca_out_406));
compressor_243_72 u_ca_243_72_407(.d_in(u_ca_in_407), .d_out(u_ca_out_407));
compressor_243_72 u_ca_243_72_408(.d_in(u_ca_in_408), .d_out(u_ca_out_408));
compressor_243_72 u_ca_243_72_409(.d_in(u_ca_in_409), .d_out(u_ca_out_409));
compressor_243_72 u_ca_243_72_410(.d_in(u_ca_in_410), .d_out(u_ca_out_410));
compressor_243_72 u_ca_243_72_411(.d_in(u_ca_in_411), .d_out(u_ca_out_411));
compressor_243_72 u_ca_243_72_412(.d_in(u_ca_in_412), .d_out(u_ca_out_412));
compressor_243_72 u_ca_243_72_413(.d_in(u_ca_in_413), .d_out(u_ca_out_413));
compressor_243_72 u_ca_243_72_414(.d_in(u_ca_in_414), .d_out(u_ca_out_414));
compressor_243_72 u_ca_243_72_415(.d_in(u_ca_in_415), .d_out(u_ca_out_415));
compressor_243_72 u_ca_243_72_416(.d_in(u_ca_in_416), .d_out(u_ca_out_416));
compressor_243_72 u_ca_243_72_417(.d_in(u_ca_in_417), .d_out(u_ca_out_417));
compressor_243_72 u_ca_243_72_418(.d_in(u_ca_in_418), .d_out(u_ca_out_418));
compressor_243_72 u_ca_243_72_419(.d_in(u_ca_in_419), .d_out(u_ca_out_419));
compressor_243_72 u_ca_243_72_420(.d_in(u_ca_in_420), .d_out(u_ca_out_420));
compressor_243_72 u_ca_243_72_421(.d_in(u_ca_in_421), .d_out(u_ca_out_421));
compressor_243_72 u_ca_243_72_422(.d_in(u_ca_in_422), .d_out(u_ca_out_422));
compressor_243_72 u_ca_243_72_423(.d_in(u_ca_in_423), .d_out(u_ca_out_423));
compressor_243_72 u_ca_243_72_424(.d_in(u_ca_in_424), .d_out(u_ca_out_424));
compressor_243_72 u_ca_243_72_425(.d_in(u_ca_in_425), .d_out(u_ca_out_425));
compressor_243_72 u_ca_243_72_426(.d_in(u_ca_in_426), .d_out(u_ca_out_426));
compressor_243_72 u_ca_243_72_427(.d_in(u_ca_in_427), .d_out(u_ca_out_427));
compressor_243_72 u_ca_243_72_428(.d_in(u_ca_in_428), .d_out(u_ca_out_428));
compressor_243_72 u_ca_243_72_429(.d_in(u_ca_in_429), .d_out(u_ca_out_429));
compressor_243_72 u_ca_243_72_430(.d_in(u_ca_in_430), .d_out(u_ca_out_430));
compressor_243_72 u_ca_243_72_431(.d_in(u_ca_in_431), .d_out(u_ca_out_431));
compressor_243_72 u_ca_243_72_432(.d_in(u_ca_in_432), .d_out(u_ca_out_432));
compressor_243_72 u_ca_243_72_433(.d_in(u_ca_in_433), .d_out(u_ca_out_433));
compressor_243_72 u_ca_243_72_434(.d_in(u_ca_in_434), .d_out(u_ca_out_434));
compressor_243_72 u_ca_243_72_435(.d_in(u_ca_in_435), .d_out(u_ca_out_435));
compressor_243_72 u_ca_243_72_436(.d_in(u_ca_in_436), .d_out(u_ca_out_436));
compressor_243_72 u_ca_243_72_437(.d_in(u_ca_in_437), .d_out(u_ca_out_437));
compressor_243_72 u_ca_243_72_438(.d_in(u_ca_in_438), .d_out(u_ca_out_438));
compressor_243_72 u_ca_243_72_439(.d_in(u_ca_in_439), .d_out(u_ca_out_439));
compressor_243_72 u_ca_243_72_440(.d_in(u_ca_in_440), .d_out(u_ca_out_440));
compressor_243_72 u_ca_243_72_441(.d_in(u_ca_in_441), .d_out(u_ca_out_441));
compressor_243_72 u_ca_243_72_442(.d_in(u_ca_in_442), .d_out(u_ca_out_442));
compressor_243_72 u_ca_243_72_443(.d_in(u_ca_in_443), .d_out(u_ca_out_443));
compressor_243_72 u_ca_243_72_444(.d_in(u_ca_in_444), .d_out(u_ca_out_444));
compressor_243_72 u_ca_243_72_445(.d_in(u_ca_in_445), .d_out(u_ca_out_445));
compressor_243_72 u_ca_243_72_446(.d_in(u_ca_in_446), .d_out(u_ca_out_446));
compressor_243_72 u_ca_243_72_447(.d_in(u_ca_in_447), .d_out(u_ca_out_447));
compressor_243_72 u_ca_243_72_448(.d_in(u_ca_in_448), .d_out(u_ca_out_448));
compressor_243_72 u_ca_243_72_449(.d_in(u_ca_in_449), .d_out(u_ca_out_449));
compressor_243_72 u_ca_243_72_450(.d_in(u_ca_in_450), .d_out(u_ca_out_450));
compressor_243_72 u_ca_243_72_451(.d_in(u_ca_in_451), .d_out(u_ca_out_451));
compressor_243_72 u_ca_243_72_452(.d_in(u_ca_in_452), .d_out(u_ca_out_452));
compressor_243_72 u_ca_243_72_453(.d_in(u_ca_in_453), .d_out(u_ca_out_453));
compressor_243_72 u_ca_243_72_454(.d_in(u_ca_in_454), .d_out(u_ca_out_454));
compressor_243_72 u_ca_243_72_455(.d_in(u_ca_in_455), .d_out(u_ca_out_455));
compressor_243_72 u_ca_243_72_456(.d_in(u_ca_in_456), .d_out(u_ca_out_456));
compressor_243_72 u_ca_243_72_457(.d_in(u_ca_in_457), .d_out(u_ca_out_457));
compressor_243_72 u_ca_243_72_458(.d_in(u_ca_in_458), .d_out(u_ca_out_458));
compressor_243_72 u_ca_243_72_459(.d_in(u_ca_in_459), .d_out(u_ca_out_459));
compressor_243_72 u_ca_243_72_460(.d_in(u_ca_in_460), .d_out(u_ca_out_460));
compressor_243_72 u_ca_243_72_461(.d_in(u_ca_in_461), .d_out(u_ca_out_461));
compressor_243_72 u_ca_243_72_462(.d_in(u_ca_in_462), .d_out(u_ca_out_462));
compressor_243_72 u_ca_243_72_463(.d_in(u_ca_in_463), .d_out(u_ca_out_463));
compressor_243_72 u_ca_243_72_464(.d_in(u_ca_in_464), .d_out(u_ca_out_464));
compressor_243_72 u_ca_243_72_465(.d_in(u_ca_in_465), .d_out(u_ca_out_465));
compressor_243_72 u_ca_243_72_466(.d_in(u_ca_in_466), .d_out(u_ca_out_466));
compressor_243_72 u_ca_243_72_467(.d_in(u_ca_in_467), .d_out(u_ca_out_467));
compressor_243_72 u_ca_243_72_468(.d_in(u_ca_in_468), .d_out(u_ca_out_468));
compressor_243_72 u_ca_243_72_469(.d_in(u_ca_in_469), .d_out(u_ca_out_469));
compressor_243_72 u_ca_243_72_470(.d_in(u_ca_in_470), .d_out(u_ca_out_470));
compressor_243_72 u_ca_243_72_471(.d_in(u_ca_in_471), .d_out(u_ca_out_471));
compressor_243_72 u_ca_243_72_472(.d_in(u_ca_in_472), .d_out(u_ca_out_472));
compressor_243_72 u_ca_243_72_473(.d_in(u_ca_in_473), .d_out(u_ca_out_473));
compressor_243_72 u_ca_243_72_474(.d_in(u_ca_in_474), .d_out(u_ca_out_474));
compressor_243_72 u_ca_243_72_475(.d_in(u_ca_in_475), .d_out(u_ca_out_475));
compressor_243_72 u_ca_243_72_476(.d_in(u_ca_in_476), .d_out(u_ca_out_476));
compressor_243_72 u_ca_243_72_477(.d_in(u_ca_in_477), .d_out(u_ca_out_477));
compressor_243_72 u_ca_243_72_478(.d_in(u_ca_in_478), .d_out(u_ca_out_478));
compressor_243_72 u_ca_243_72_479(.d_in(u_ca_in_479), .d_out(u_ca_out_479));
compressor_243_72 u_ca_243_72_480(.d_in(u_ca_in_480), .d_out(u_ca_out_480));
compressor_243_72 u_ca_243_72_481(.d_in(u_ca_in_481), .d_out(u_ca_out_481));
compressor_243_72 u_ca_243_72_482(.d_in(u_ca_in_482), .d_out(u_ca_out_482));
compressor_243_72 u_ca_243_72_483(.d_in(u_ca_in_483), .d_out(u_ca_out_483));
compressor_243_72 u_ca_243_72_484(.d_in(u_ca_in_484), .d_out(u_ca_out_484));
compressor_243_72 u_ca_243_72_485(.d_in(u_ca_in_485), .d_out(u_ca_out_485));
compressor_243_72 u_ca_243_72_486(.d_in(u_ca_in_486), .d_out(u_ca_out_486));
compressor_243_72 u_ca_243_72_487(.d_in(u_ca_in_487), .d_out(u_ca_out_487));
compressor_243_72 u_ca_243_72_488(.d_in(u_ca_in_488), .d_out(u_ca_out_488));
compressor_243_72 u_ca_243_72_489(.d_in(u_ca_in_489), .d_out(u_ca_out_489));
compressor_243_72 u_ca_243_72_490(.d_in(u_ca_in_490), .d_out(u_ca_out_490));
compressor_243_72 u_ca_243_72_491(.d_in(u_ca_in_491), .d_out(u_ca_out_491));
compressor_243_72 u_ca_243_72_492(.d_in(u_ca_in_492), .d_out(u_ca_out_492));
compressor_243_72 u_ca_243_72_493(.d_in(u_ca_in_493), .d_out(u_ca_out_493));
compressor_243_72 u_ca_243_72_494(.d_in(u_ca_in_494), .d_out(u_ca_out_494));
compressor_243_72 u_ca_243_72_495(.d_in(u_ca_in_495), .d_out(u_ca_out_495));
compressor_243_72 u_ca_243_72_496(.d_in(u_ca_in_496), .d_out(u_ca_out_496));
compressor_243_72 u_ca_243_72_497(.d_in(u_ca_in_497), .d_out(u_ca_out_497));
compressor_243_72 u_ca_243_72_498(.d_in(u_ca_in_498), .d_out(u_ca_out_498));
compressor_243_72 u_ca_243_72_499(.d_in(u_ca_in_499), .d_out(u_ca_out_499));
compressor_243_72 u_ca_243_72_500(.d_in(u_ca_in_500), .d_out(u_ca_out_500));
compressor_243_72 u_ca_243_72_501(.d_in(u_ca_in_501), .d_out(u_ca_out_501));
compressor_243_72 u_ca_243_72_502(.d_in(u_ca_in_502), .d_out(u_ca_out_502));
compressor_243_72 u_ca_243_72_503(.d_in(u_ca_in_503), .d_out(u_ca_out_503));
compressor_243_72 u_ca_243_72_504(.d_in(u_ca_in_504), .d_out(u_ca_out_504));
compressor_243_72 u_ca_243_72_505(.d_in(u_ca_in_505), .d_out(u_ca_out_505));
compressor_243_72 u_ca_243_72_506(.d_in(u_ca_in_506), .d_out(u_ca_out_506));
compressor_243_72 u_ca_243_72_507(.d_in(u_ca_in_507), .d_out(u_ca_out_507));
compressor_243_72 u_ca_243_72_508(.d_in(u_ca_in_508), .d_out(u_ca_out_508));
compressor_243_72 u_ca_243_72_509(.d_in(u_ca_in_509), .d_out(u_ca_out_509));
compressor_243_72 u_ca_243_72_510(.d_in(u_ca_in_510), .d_out(u_ca_out_510));
compressor_243_72 u_ca_243_72_511(.d_in(u_ca_in_511), .d_out(u_ca_out_511));
compressor_243_72 u_ca_243_72_512(.d_in(u_ca_in_512), .d_out(u_ca_out_512));
compressor_243_72 u_ca_243_72_513(.d_in(u_ca_in_513), .d_out(u_ca_out_513));
compressor_243_72 u_ca_243_72_514(.d_in(u_ca_in_514), .d_out(u_ca_out_514));
compressor_243_72 u_ca_243_72_515(.d_in(u_ca_in_515), .d_out(u_ca_out_515));
compressor_243_72 u_ca_243_72_516(.d_in(u_ca_in_516), .d_out(u_ca_out_516));
compressor_243_72 u_ca_243_72_517(.d_in(u_ca_in_517), .d_out(u_ca_out_517));
compressor_243_72 u_ca_243_72_518(.d_in(u_ca_in_518), .d_out(u_ca_out_518));
compressor_243_72 u_ca_243_72_519(.d_in(u_ca_in_519), .d_out(u_ca_out_519));
compressor_243_72 u_ca_243_72_520(.d_in(u_ca_in_520), .d_out(u_ca_out_520));
compressor_243_72 u_ca_243_72_521(.d_in(u_ca_in_521), .d_out(u_ca_out_521));
compressor_243_72 u_ca_243_72_522(.d_in(u_ca_in_522), .d_out(u_ca_out_522));
compressor_243_72 u_ca_243_72_523(.d_in(u_ca_in_523), .d_out(u_ca_out_523));
compressor_243_72 u_ca_243_72_524(.d_in(u_ca_in_524), .d_out(u_ca_out_524));
compressor_243_72 u_ca_243_72_525(.d_in(u_ca_in_525), .d_out(u_ca_out_525));
compressor_243_72 u_ca_243_72_526(.d_in(u_ca_in_526), .d_out(u_ca_out_526));
compressor_243_72 u_ca_243_72_527(.d_in(u_ca_in_527), .d_out(u_ca_out_527));
compressor_243_72 u_ca_243_72_528(.d_in(u_ca_in_528), .d_out(u_ca_out_528));
compressor_243_72 u_ca_243_72_529(.d_in(u_ca_in_529), .d_out(u_ca_out_529));
compressor_243_72 u_ca_243_72_530(.d_in(u_ca_in_530), .d_out(u_ca_out_530));
compressor_243_72 u_ca_243_72_531(.d_in(u_ca_in_531), .d_out(u_ca_out_531));
compressor_243_72 u_ca_243_72_532(.d_in(u_ca_in_532), .d_out(u_ca_out_532));
compressor_243_72 u_ca_243_72_533(.d_in(u_ca_in_533), .d_out(u_ca_out_533));
compressor_243_72 u_ca_243_72_534(.d_in(u_ca_in_534), .d_out(u_ca_out_534));
compressor_243_72 u_ca_243_72_535(.d_in(u_ca_in_535), .d_out(u_ca_out_535));
compressor_243_72 u_ca_243_72_536(.d_in(u_ca_in_536), .d_out(u_ca_out_536));
compressor_243_72 u_ca_243_72_537(.d_in(u_ca_in_537), .d_out(u_ca_out_537));
compressor_243_72 u_ca_243_72_538(.d_in(u_ca_in_538), .d_out(u_ca_out_538));
compressor_243_72 u_ca_243_72_539(.d_in(u_ca_in_539), .d_out(u_ca_out_539));
compressor_243_72 u_ca_243_72_540(.d_in(u_ca_in_540), .d_out(u_ca_out_540));
compressor_243_72 u_ca_243_72_541(.d_in(u_ca_in_541), .d_out(u_ca_out_541));
compressor_243_72 u_ca_243_72_542(.d_in(u_ca_in_542), .d_out(u_ca_out_542));
compressor_243_72 u_ca_243_72_543(.d_in(u_ca_in_543), .d_out(u_ca_out_543));
compressor_243_72 u_ca_243_72_544(.d_in(u_ca_in_544), .d_out(u_ca_out_544));
compressor_243_72 u_ca_243_72_545(.d_in(u_ca_in_545), .d_out(u_ca_out_545));
compressor_243_72 u_ca_243_72_546(.d_in(u_ca_in_546), .d_out(u_ca_out_546));
compressor_243_72 u_ca_243_72_547(.d_in(u_ca_in_547), .d_out(u_ca_out_547));
compressor_243_72 u_ca_243_72_548(.d_in(u_ca_in_548), .d_out(u_ca_out_548));
compressor_243_72 u_ca_243_72_549(.d_in(u_ca_in_549), .d_out(u_ca_out_549));
compressor_243_72 u_ca_243_72_550(.d_in(u_ca_in_550), .d_out(u_ca_out_550));
compressor_243_72 u_ca_243_72_551(.d_in(u_ca_in_551), .d_out(u_ca_out_551));
compressor_243_72 u_ca_243_72_552(.d_in(u_ca_in_552), .d_out(u_ca_out_552));
compressor_243_72 u_ca_243_72_553(.d_in(u_ca_in_553), .d_out(u_ca_out_553));
compressor_243_72 u_ca_243_72_554(.d_in(u_ca_in_554), .d_out(u_ca_out_554));
compressor_243_72 u_ca_243_72_555(.d_in(u_ca_in_555), .d_out(u_ca_out_555));
compressor_243_72 u_ca_243_72_556(.d_in(u_ca_in_556), .d_out(u_ca_out_556));
compressor_243_72 u_ca_243_72_557(.d_in(u_ca_in_557), .d_out(u_ca_out_557));
compressor_243_72 u_ca_243_72_558(.d_in(u_ca_in_558), .d_out(u_ca_out_558));
compressor_243_72 u_ca_243_72_559(.d_in(u_ca_in_559), .d_out(u_ca_out_559));
compressor_243_72 u_ca_243_72_560(.d_in(u_ca_in_560), .d_out(u_ca_out_560));
compressor_243_72 u_ca_243_72_561(.d_in(u_ca_in_561), .d_out(u_ca_out_561));
compressor_243_72 u_ca_243_72_562(.d_in(u_ca_in_562), .d_out(u_ca_out_562));
compressor_243_72 u_ca_243_72_563(.d_in(u_ca_in_563), .d_out(u_ca_out_563));
compressor_243_72 u_ca_243_72_564(.d_in(u_ca_in_564), .d_out(u_ca_out_564));
compressor_243_72 u_ca_243_72_565(.d_in(u_ca_in_565), .d_out(u_ca_out_565));
compressor_243_72 u_ca_243_72_566(.d_in(u_ca_in_566), .d_out(u_ca_out_566));
compressor_243_72 u_ca_243_72_567(.d_in(u_ca_in_567), .d_out(u_ca_out_567));
compressor_243_72 u_ca_243_72_568(.d_in(u_ca_in_568), .d_out(u_ca_out_568));
compressor_243_72 u_ca_243_72_569(.d_in(u_ca_in_569), .d_out(u_ca_out_569));
compressor_243_72 u_ca_243_72_570(.d_in(u_ca_in_570), .d_out(u_ca_out_570));
compressor_243_72 u_ca_243_72_571(.d_in(u_ca_in_571), .d_out(u_ca_out_571));
compressor_243_72 u_ca_243_72_572(.d_in(u_ca_in_572), .d_out(u_ca_out_572));
compressor_243_72 u_ca_243_72_573(.d_in(u_ca_in_573), .d_out(u_ca_out_573));
compressor_243_72 u_ca_243_72_574(.d_in(u_ca_in_574), .d_out(u_ca_out_574));
compressor_243_72 u_ca_243_72_575(.d_in(u_ca_in_575), .d_out(u_ca_out_575));
compressor_243_72 u_ca_243_72_576(.d_in(u_ca_in_576), .d_out(u_ca_out_576));
compressor_243_72 u_ca_243_72_577(.d_in(u_ca_in_577), .d_out(u_ca_out_577));
compressor_243_72 u_ca_243_72_578(.d_in(u_ca_in_578), .d_out(u_ca_out_578));
compressor_243_72 u_ca_243_72_579(.d_in(u_ca_in_579), .d_out(u_ca_out_579));
compressor_243_72 u_ca_243_72_580(.d_in(u_ca_in_580), .d_out(u_ca_out_580));
compressor_243_72 u_ca_243_72_581(.d_in(u_ca_in_581), .d_out(u_ca_out_581));
compressor_243_72 u_ca_243_72_582(.d_in(u_ca_in_582), .d_out(u_ca_out_582));
compressor_243_72 u_ca_243_72_583(.d_in(u_ca_in_583), .d_out(u_ca_out_583));
compressor_243_72 u_ca_243_72_584(.d_in(u_ca_in_584), .d_out(u_ca_out_584));
compressor_243_72 u_ca_243_72_585(.d_in(u_ca_in_585), .d_out(u_ca_out_585));
compressor_243_72 u_ca_243_72_586(.d_in(u_ca_in_586), .d_out(u_ca_out_586));
compressor_243_72 u_ca_243_72_587(.d_in(u_ca_in_587), .d_out(u_ca_out_587));
compressor_243_72 u_ca_243_72_588(.d_in(u_ca_in_588), .d_out(u_ca_out_588));
compressor_243_72 u_ca_243_72_589(.d_in(u_ca_in_589), .d_out(u_ca_out_589));
compressor_243_72 u_ca_243_72_590(.d_in(u_ca_in_590), .d_out(u_ca_out_590));
compressor_243_72 u_ca_243_72_591(.d_in(u_ca_in_591), .d_out(u_ca_out_591));
compressor_243_72 u_ca_243_72_592(.d_in(u_ca_in_592), .d_out(u_ca_out_592));
compressor_243_72 u_ca_243_72_593(.d_in(u_ca_in_593), .d_out(u_ca_out_593));
compressor_243_72 u_ca_243_72_594(.d_in(u_ca_in_594), .d_out(u_ca_out_594));
compressor_243_72 u_ca_243_72_595(.d_in(u_ca_in_595), .d_out(u_ca_out_595));
compressor_243_72 u_ca_243_72_596(.d_in(u_ca_in_596), .d_out(u_ca_out_596));
compressor_243_72 u_ca_243_72_597(.d_in(u_ca_in_597), .d_out(u_ca_out_597));
compressor_243_72 u_ca_243_72_598(.d_in(u_ca_in_598), .d_out(u_ca_out_598));
compressor_243_72 u_ca_243_72_599(.d_in(u_ca_in_599), .d_out(u_ca_out_599));
compressor_243_72 u_ca_243_72_600(.d_in(u_ca_in_600), .d_out(u_ca_out_600));
compressor_243_72 u_ca_243_72_601(.d_in(u_ca_in_601), .d_out(u_ca_out_601));
compressor_243_72 u_ca_243_72_602(.d_in(u_ca_in_602), .d_out(u_ca_out_602));
compressor_243_72 u_ca_243_72_603(.d_in(u_ca_in_603), .d_out(u_ca_out_603));
compressor_243_72 u_ca_243_72_604(.d_in(u_ca_in_604), .d_out(u_ca_out_604));
compressor_243_72 u_ca_243_72_605(.d_in(u_ca_in_605), .d_out(u_ca_out_605));
compressor_243_72 u_ca_243_72_606(.d_in(u_ca_in_606), .d_out(u_ca_out_606));
compressor_243_72 u_ca_243_72_607(.d_in(u_ca_in_607), .d_out(u_ca_out_607));
compressor_243_72 u_ca_243_72_608(.d_in(u_ca_in_608), .d_out(u_ca_out_608));
compressor_243_72 u_ca_243_72_609(.d_in(u_ca_in_609), .d_out(u_ca_out_609));
compressor_243_72 u_ca_243_72_610(.d_in(u_ca_in_610), .d_out(u_ca_out_610));
compressor_243_72 u_ca_243_72_611(.d_in(u_ca_in_611), .d_out(u_ca_out_611));
compressor_243_72 u_ca_243_72_612(.d_in(u_ca_in_612), .d_out(u_ca_out_612));
compressor_243_72 u_ca_243_72_613(.d_in(u_ca_in_613), .d_out(u_ca_out_613));
compressor_243_72 u_ca_243_72_614(.d_in(u_ca_in_614), .d_out(u_ca_out_614));
compressor_243_72 u_ca_243_72_615(.d_in(u_ca_in_615), .d_out(u_ca_out_615));
compressor_243_72 u_ca_243_72_616(.d_in(u_ca_in_616), .d_out(u_ca_out_616));
compressor_243_72 u_ca_243_72_617(.d_in(u_ca_in_617), .d_out(u_ca_out_617));
compressor_243_72 u_ca_243_72_618(.d_in(u_ca_in_618), .d_out(u_ca_out_618));
compressor_243_72 u_ca_243_72_619(.d_in(u_ca_in_619), .d_out(u_ca_out_619));
compressor_243_72 u_ca_243_72_620(.d_in(u_ca_in_620), .d_out(u_ca_out_620));
compressor_243_72 u_ca_243_72_621(.d_in(u_ca_in_621), .d_out(u_ca_out_621));
compressor_243_72 u_ca_243_72_622(.d_in(u_ca_in_622), .d_out(u_ca_out_622));
compressor_243_72 u_ca_243_72_623(.d_in(u_ca_in_623), .d_out(u_ca_out_623));
compressor_243_72 u_ca_243_72_624(.d_in(u_ca_in_624), .d_out(u_ca_out_624));
compressor_243_72 u_ca_243_72_625(.d_in(u_ca_in_625), .d_out(u_ca_out_625));
compressor_243_72 u_ca_243_72_626(.d_in(u_ca_in_626), .d_out(u_ca_out_626));
compressor_243_72 u_ca_243_72_627(.d_in(u_ca_in_627), .d_out(u_ca_out_627));
compressor_243_72 u_ca_243_72_628(.d_in(u_ca_in_628), .d_out(u_ca_out_628));
compressor_243_72 u_ca_243_72_629(.d_in(u_ca_in_629), .d_out(u_ca_out_629));
compressor_243_72 u_ca_243_72_630(.d_in(u_ca_in_630), .d_out(u_ca_out_630));
compressor_243_72 u_ca_243_72_631(.d_in(u_ca_in_631), .d_out(u_ca_out_631));
compressor_243_72 u_ca_243_72_632(.d_in(u_ca_in_632), .d_out(u_ca_out_632));
compressor_243_72 u_ca_243_72_633(.d_in(u_ca_in_633), .d_out(u_ca_out_633));
compressor_243_72 u_ca_243_72_634(.d_in(u_ca_in_634), .d_out(u_ca_out_634));
compressor_243_72 u_ca_243_72_635(.d_in(u_ca_in_635), .d_out(u_ca_out_635));
compressor_243_72 u_ca_243_72_636(.d_in(u_ca_in_636), .d_out(u_ca_out_636));
compressor_243_72 u_ca_243_72_637(.d_in(u_ca_in_637), .d_out(u_ca_out_637));
compressor_243_72 u_ca_243_72_638(.d_in(u_ca_in_638), .d_out(u_ca_out_638));
compressor_243_72 u_ca_243_72_639(.d_in(u_ca_in_639), .d_out(u_ca_out_639));
compressor_243_72 u_ca_243_72_640(.d_in(u_ca_in_640), .d_out(u_ca_out_640));
compressor_243_72 u_ca_243_72_641(.d_in(u_ca_in_641), .d_out(u_ca_out_641));
compressor_243_72 u_ca_243_72_642(.d_in(u_ca_in_642), .d_out(u_ca_out_642));
compressor_243_72 u_ca_243_72_643(.d_in(u_ca_in_643), .d_out(u_ca_out_643));
compressor_243_72 u_ca_243_72_644(.d_in(u_ca_in_644), .d_out(u_ca_out_644));
compressor_243_72 u_ca_243_72_645(.d_in(u_ca_in_645), .d_out(u_ca_out_645));
compressor_243_72 u_ca_243_72_646(.d_in(u_ca_in_646), .d_out(u_ca_out_646));
compressor_243_72 u_ca_243_72_647(.d_in(u_ca_in_647), .d_out(u_ca_out_647));
compressor_243_72 u_ca_243_72_648(.d_in(u_ca_in_648), .d_out(u_ca_out_648));
compressor_243_72 u_ca_243_72_649(.d_in(u_ca_in_649), .d_out(u_ca_out_649));
compressor_243_72 u_ca_243_72_650(.d_in(u_ca_in_650), .d_out(u_ca_out_650));
compressor_243_72 u_ca_243_72_651(.d_in(u_ca_in_651), .d_out(u_ca_out_651));
compressor_243_72 u_ca_243_72_652(.d_in(u_ca_in_652), .d_out(u_ca_out_652));
compressor_243_72 u_ca_243_72_653(.d_in(u_ca_in_653), .d_out(u_ca_out_653));
compressor_243_72 u_ca_243_72_654(.d_in(u_ca_in_654), .d_out(u_ca_out_654));
compressor_243_72 u_ca_243_72_655(.d_in(u_ca_in_655), .d_out(u_ca_out_655));
compressor_243_72 u_ca_243_72_656(.d_in(u_ca_in_656), .d_out(u_ca_out_656));
compressor_243_72 u_ca_243_72_657(.d_in(u_ca_in_657), .d_out(u_ca_out_657));
compressor_243_72 u_ca_243_72_658(.d_in(u_ca_in_658), .d_out(u_ca_out_658));
compressor_243_72 u_ca_243_72_659(.d_in(u_ca_in_659), .d_out(u_ca_out_659));
compressor_243_72 u_ca_243_72_660(.d_in(u_ca_in_660), .d_out(u_ca_out_660));
compressor_243_72 u_ca_243_72_661(.d_in(u_ca_in_661), .d_out(u_ca_out_661));
compressor_243_72 u_ca_243_72_662(.d_in(u_ca_in_662), .d_out(u_ca_out_662));
compressor_243_72 u_ca_243_72_663(.d_in(u_ca_in_663), .d_out(u_ca_out_663));
compressor_243_72 u_ca_243_72_664(.d_in(u_ca_in_664), .d_out(u_ca_out_664));
compressor_243_72 u_ca_243_72_665(.d_in(u_ca_in_665), .d_out(u_ca_out_665));
compressor_243_72 u_ca_243_72_666(.d_in(u_ca_in_666), .d_out(u_ca_out_666));
compressor_243_72 u_ca_243_72_667(.d_in(u_ca_in_667), .d_out(u_ca_out_667));
compressor_243_72 u_ca_243_72_668(.d_in(u_ca_in_668), .d_out(u_ca_out_668));
compressor_243_72 u_ca_243_72_669(.d_in(u_ca_in_669), .d_out(u_ca_out_669));
compressor_243_72 u_ca_243_72_670(.d_in(u_ca_in_670), .d_out(u_ca_out_670));
compressor_243_72 u_ca_243_72_671(.d_in(u_ca_in_671), .d_out(u_ca_out_671));
compressor_243_72 u_ca_243_72_672(.d_in(u_ca_in_672), .d_out(u_ca_out_672));
compressor_243_72 u_ca_243_72_673(.d_in(u_ca_in_673), .d_out(u_ca_out_673));
compressor_243_72 u_ca_243_72_674(.d_in(u_ca_in_674), .d_out(u_ca_out_674));
compressor_243_72 u_ca_243_72_675(.d_in(u_ca_in_675), .d_out(u_ca_out_675));
compressor_243_72 u_ca_243_72_676(.d_in(u_ca_in_676), .d_out(u_ca_out_676));
compressor_243_72 u_ca_243_72_677(.d_in(u_ca_in_677), .d_out(u_ca_out_677));
compressor_243_72 u_ca_243_72_678(.d_in(u_ca_in_678), .d_out(u_ca_out_678));
compressor_243_72 u_ca_243_72_679(.d_in(u_ca_in_679), .d_out(u_ca_out_679));
compressor_243_72 u_ca_243_72_680(.d_in(u_ca_in_680), .d_out(u_ca_out_680));
compressor_243_72 u_ca_243_72_681(.d_in(u_ca_in_681), .d_out(u_ca_out_681));
compressor_243_72 u_ca_243_72_682(.d_in(u_ca_in_682), .d_out(u_ca_out_682));
compressor_243_72 u_ca_243_72_683(.d_in(u_ca_in_683), .d_out(u_ca_out_683));
compressor_243_72 u_ca_243_72_684(.d_in(u_ca_in_684), .d_out(u_ca_out_684));
compressor_243_72 u_ca_243_72_685(.d_in(u_ca_in_685), .d_out(u_ca_out_685));
compressor_243_72 u_ca_243_72_686(.d_in(u_ca_in_686), .d_out(u_ca_out_686));
compressor_243_72 u_ca_243_72_687(.d_in(u_ca_in_687), .d_out(u_ca_out_687));
compressor_243_72 u_ca_243_72_688(.d_in(u_ca_in_688), .d_out(u_ca_out_688));
compressor_243_72 u_ca_243_72_689(.d_in(u_ca_in_689), .d_out(u_ca_out_689));
compressor_243_72 u_ca_243_72_690(.d_in(u_ca_in_690), .d_out(u_ca_out_690));
compressor_243_72 u_ca_243_72_691(.d_in(u_ca_in_691), .d_out(u_ca_out_691));
compressor_243_72 u_ca_243_72_692(.d_in(u_ca_in_692), .d_out(u_ca_out_692));
compressor_243_72 u_ca_243_72_693(.d_in(u_ca_in_693), .d_out(u_ca_out_693));
compressor_243_72 u_ca_243_72_694(.d_in(u_ca_in_694), .d_out(u_ca_out_694));
compressor_243_72 u_ca_243_72_695(.d_in(u_ca_in_695), .d_out(u_ca_out_695));
compressor_243_72 u_ca_243_72_696(.d_in(u_ca_in_696), .d_out(u_ca_out_696));
compressor_243_72 u_ca_243_72_697(.d_in(u_ca_in_697), .d_out(u_ca_out_697));
compressor_243_72 u_ca_243_72_698(.d_in(u_ca_in_698), .d_out(u_ca_out_698));
compressor_243_72 u_ca_243_72_699(.d_in(u_ca_in_699), .d_out(u_ca_out_699));
compressor_243_72 u_ca_243_72_700(.d_in(u_ca_in_700), .d_out(u_ca_out_700));
compressor_243_72 u_ca_243_72_701(.d_in(u_ca_in_701), .d_out(u_ca_out_701));
compressor_243_72 u_ca_243_72_702(.d_in(u_ca_in_702), .d_out(u_ca_out_702));
compressor_243_72 u_ca_243_72_703(.d_in(u_ca_in_703), .d_out(u_ca_out_703));
compressor_243_72 u_ca_243_72_704(.d_in(u_ca_in_704), .d_out(u_ca_out_704));
compressor_243_72 u_ca_243_72_705(.d_in(u_ca_in_705), .d_out(u_ca_out_705));
compressor_243_72 u_ca_243_72_706(.d_in(u_ca_in_706), .d_out(u_ca_out_706));
compressor_243_72 u_ca_243_72_707(.d_in(u_ca_in_707), .d_out(u_ca_out_707));
compressor_243_72 u_ca_243_72_708(.d_in(u_ca_in_708), .d_out(u_ca_out_708));
compressor_243_72 u_ca_243_72_709(.d_in(u_ca_in_709), .d_out(u_ca_out_709));
compressor_243_72 u_ca_243_72_710(.d_in(u_ca_in_710), .d_out(u_ca_out_710));
compressor_243_72 u_ca_243_72_711(.d_in(u_ca_in_711), .d_out(u_ca_out_711));
compressor_243_72 u_ca_243_72_712(.d_in(u_ca_in_712), .d_out(u_ca_out_712));
compressor_243_72 u_ca_243_72_713(.d_in(u_ca_in_713), .d_out(u_ca_out_713));
compressor_243_72 u_ca_243_72_714(.d_in(u_ca_in_714), .d_out(u_ca_out_714));
compressor_243_72 u_ca_243_72_715(.d_in(u_ca_in_715), .d_out(u_ca_out_715));
compressor_243_72 u_ca_243_72_716(.d_in(u_ca_in_716), .d_out(u_ca_out_716));
compressor_243_72 u_ca_243_72_717(.d_in(u_ca_in_717), .d_out(u_ca_out_717));
compressor_243_72 u_ca_243_72_718(.d_in(u_ca_in_718), .d_out(u_ca_out_718));
compressor_243_72 u_ca_243_72_719(.d_in(u_ca_in_719), .d_out(u_ca_out_719));
compressor_243_72 u_ca_243_72_720(.d_in(u_ca_in_720), .d_out(u_ca_out_720));
compressor_243_72 u_ca_243_72_721(.d_in(u_ca_in_721), .d_out(u_ca_out_721));
compressor_243_72 u_ca_243_72_722(.d_in(u_ca_in_722), .d_out(u_ca_out_722));
compressor_243_72 u_ca_243_72_723(.d_in(u_ca_in_723), .d_out(u_ca_out_723));
compressor_243_72 u_ca_243_72_724(.d_in(u_ca_in_724), .d_out(u_ca_out_724));
compressor_243_72 u_ca_243_72_725(.d_in(u_ca_in_725), .d_out(u_ca_out_725));
compressor_243_72 u_ca_243_72_726(.d_in(u_ca_in_726), .d_out(u_ca_out_726));
compressor_243_72 u_ca_243_72_727(.d_in(u_ca_in_727), .d_out(u_ca_out_727));
compressor_243_72 u_ca_243_72_728(.d_in(u_ca_in_728), .d_out(u_ca_out_728));
compressor_243_72 u_ca_243_72_729(.d_in(u_ca_in_729), .d_out(u_ca_out_729));
compressor_243_72 u_ca_243_72_730(.d_in(u_ca_in_730), .d_out(u_ca_out_730));
compressor_243_72 u_ca_243_72_731(.d_in(u_ca_in_731), .d_out(u_ca_out_731));
compressor_243_72 u_ca_243_72_732(.d_in(u_ca_in_732), .d_out(u_ca_out_732));
compressor_243_72 u_ca_243_72_733(.d_in(u_ca_in_733), .d_out(u_ca_out_733));
compressor_243_72 u_ca_243_72_734(.d_in(u_ca_in_734), .d_out(u_ca_out_734));
compressor_243_72 u_ca_243_72_735(.d_in(u_ca_in_735), .d_out(u_ca_out_735));
compressor_243_72 u_ca_243_72_736(.d_in(u_ca_in_736), .d_out(u_ca_out_736));
compressor_243_72 u_ca_243_72_737(.d_in(u_ca_in_737), .d_out(u_ca_out_737));
compressor_243_72 u_ca_243_72_738(.d_in(u_ca_in_738), .d_out(u_ca_out_738));
compressor_243_72 u_ca_243_72_739(.d_in(u_ca_in_739), .d_out(u_ca_out_739));
compressor_243_72 u_ca_243_72_740(.d_in(u_ca_in_740), .d_out(u_ca_out_740));
compressor_243_72 u_ca_243_72_741(.d_in(u_ca_in_741), .d_out(u_ca_out_741));
compressor_243_72 u_ca_243_72_742(.d_in(u_ca_in_742), .d_out(u_ca_out_742));
compressor_243_72 u_ca_243_72_743(.d_in(u_ca_in_743), .d_out(u_ca_out_743));
compressor_243_72 u_ca_243_72_744(.d_in(u_ca_in_744), .d_out(u_ca_out_744));
compressor_243_72 u_ca_243_72_745(.d_in(u_ca_in_745), .d_out(u_ca_out_745));
compressor_243_72 u_ca_243_72_746(.d_in(u_ca_in_746), .d_out(u_ca_out_746));
compressor_243_72 u_ca_243_72_747(.d_in(u_ca_in_747), .d_out(u_ca_out_747));
compressor_243_72 u_ca_243_72_748(.d_in(u_ca_in_748), .d_out(u_ca_out_748));
compressor_243_72 u_ca_243_72_749(.d_in(u_ca_in_749), .d_out(u_ca_out_749));
compressor_243_72 u_ca_243_72_750(.d_in(u_ca_in_750), .d_out(u_ca_out_750));
compressor_243_72 u_ca_243_72_751(.d_in(u_ca_in_751), .d_out(u_ca_out_751));
compressor_243_72 u_ca_243_72_752(.d_in(u_ca_in_752), .d_out(u_ca_out_752));
compressor_243_72 u_ca_243_72_753(.d_in(u_ca_in_753), .d_out(u_ca_out_753));
compressor_243_72 u_ca_243_72_754(.d_in(u_ca_in_754), .d_out(u_ca_out_754));
compressor_243_72 u_ca_243_72_755(.d_in(u_ca_in_755), .d_out(u_ca_out_755));
compressor_243_72 u_ca_243_72_756(.d_in(u_ca_in_756), .d_out(u_ca_out_756));
compressor_243_72 u_ca_243_72_757(.d_in(u_ca_in_757), .d_out(u_ca_out_757));
compressor_243_72 u_ca_243_72_758(.d_in(u_ca_in_758), .d_out(u_ca_out_758));
compressor_243_72 u_ca_243_72_759(.d_in(u_ca_in_759), .d_out(u_ca_out_759));
compressor_243_72 u_ca_243_72_760(.d_in(u_ca_in_760), .d_out(u_ca_out_760));
compressor_243_72 u_ca_243_72_761(.d_in(u_ca_in_761), .d_out(u_ca_out_761));
compressor_243_72 u_ca_243_72_762(.d_in(u_ca_in_762), .d_out(u_ca_out_762));
compressor_243_72 u_ca_243_72_763(.d_in(u_ca_in_763), .d_out(u_ca_out_763));
compressor_243_72 u_ca_243_72_764(.d_in(u_ca_in_764), .d_out(u_ca_out_764));
compressor_243_72 u_ca_243_72_765(.d_in(u_ca_in_765), .d_out(u_ca_out_765));
compressor_243_72 u_ca_243_72_766(.d_in(u_ca_in_766), .d_out(u_ca_out_766));
compressor_243_72 u_ca_243_72_767(.d_in(u_ca_in_767), .d_out(u_ca_out_767));
compressor_243_72 u_ca_243_72_768(.d_in(u_ca_in_768), .d_out(u_ca_out_768));
compressor_243_72 u_ca_243_72_769(.d_in(u_ca_in_769), .d_out(u_ca_out_769));
compressor_243_72 u_ca_243_72_770(.d_in(u_ca_in_770), .d_out(u_ca_out_770));
compressor_243_72 u_ca_243_72_771(.d_in(u_ca_in_771), .d_out(u_ca_out_771));
compressor_243_72 u_ca_243_72_772(.d_in(u_ca_in_772), .d_out(u_ca_out_772));
compressor_243_72 u_ca_243_72_773(.d_in(u_ca_in_773), .d_out(u_ca_out_773));
compressor_243_72 u_ca_243_72_774(.d_in(u_ca_in_774), .d_out(u_ca_out_774));
compressor_243_72 u_ca_243_72_775(.d_in(u_ca_in_775), .d_out(u_ca_out_775));
compressor_243_72 u_ca_243_72_776(.d_in(u_ca_in_776), .d_out(u_ca_out_776));
compressor_243_72 u_ca_243_72_777(.d_in(u_ca_in_777), .d_out(u_ca_out_777));
compressor_243_72 u_ca_243_72_778(.d_in(u_ca_in_778), .d_out(u_ca_out_778));
compressor_243_72 u_ca_243_72_779(.d_in(u_ca_in_779), .d_out(u_ca_out_779));
compressor_243_72 u_ca_243_72_780(.d_in(u_ca_in_780), .d_out(u_ca_out_780));
compressor_243_72 u_ca_243_72_781(.d_in(u_ca_in_781), .d_out(u_ca_out_781));
compressor_243_72 u_ca_243_72_782(.d_in(u_ca_in_782), .d_out(u_ca_out_782));
compressor_243_72 u_ca_243_72_783(.d_in(u_ca_in_783), .d_out(u_ca_out_783));
compressor_243_72 u_ca_243_72_784(.d_in(u_ca_in_784), .d_out(u_ca_out_784));
compressor_243_72 u_ca_243_72_785(.d_in(u_ca_in_785), .d_out(u_ca_out_785));
compressor_243_72 u_ca_243_72_786(.d_in(u_ca_in_786), .d_out(u_ca_out_786));
compressor_243_72 u_ca_243_72_787(.d_in(u_ca_in_787), .d_out(u_ca_out_787));
compressor_243_72 u_ca_243_72_788(.d_in(u_ca_in_788), .d_out(u_ca_out_788));
compressor_243_72 u_ca_243_72_789(.d_in(u_ca_in_789), .d_out(u_ca_out_789));
compressor_243_72 u_ca_243_72_790(.d_in(u_ca_in_790), .d_out(u_ca_out_790));
compressor_243_72 u_ca_243_72_791(.d_in(u_ca_in_791), .d_out(u_ca_out_791));
compressor_243_72 u_ca_243_72_792(.d_in(u_ca_in_792), .d_out(u_ca_out_792));
compressor_243_72 u_ca_243_72_793(.d_in(u_ca_in_793), .d_out(u_ca_out_793));
compressor_243_72 u_ca_243_72_794(.d_in(u_ca_in_794), .d_out(u_ca_out_794));
compressor_243_72 u_ca_243_72_795(.d_in(u_ca_in_795), .d_out(u_ca_out_795));
compressor_243_72 u_ca_243_72_796(.d_in(u_ca_in_796), .d_out(u_ca_out_796));
compressor_243_72 u_ca_243_72_797(.d_in(u_ca_in_797), .d_out(u_ca_out_797));
compressor_243_72 u_ca_243_72_798(.d_in(u_ca_in_798), .d_out(u_ca_out_798));
compressor_243_72 u_ca_243_72_799(.d_in(u_ca_in_799), .d_out(u_ca_out_799));
compressor_243_72 u_ca_243_72_800(.d_in(u_ca_in_800), .d_out(u_ca_out_800));
compressor_243_72 u_ca_243_72_801(.d_in(u_ca_in_801), .d_out(u_ca_out_801));
compressor_243_72 u_ca_243_72_802(.d_in(u_ca_in_802), .d_out(u_ca_out_802));
compressor_243_72 u_ca_243_72_803(.d_in(u_ca_in_803), .d_out(u_ca_out_803));
compressor_243_72 u_ca_243_72_804(.d_in(u_ca_in_804), .d_out(u_ca_out_804));
compressor_243_72 u_ca_243_72_805(.d_in(u_ca_in_805), .d_out(u_ca_out_805));
compressor_243_72 u_ca_243_72_806(.d_in(u_ca_in_806), .d_out(u_ca_out_806));
compressor_243_72 u_ca_243_72_807(.d_in(u_ca_in_807), .d_out(u_ca_out_807));
compressor_243_72 u_ca_243_72_808(.d_in(u_ca_in_808), .d_out(u_ca_out_808));
compressor_243_72 u_ca_243_72_809(.d_in(u_ca_in_809), .d_out(u_ca_out_809));
compressor_243_72 u_ca_243_72_810(.d_in(u_ca_in_810), .d_out(u_ca_out_810));
compressor_243_72 u_ca_243_72_811(.d_in(u_ca_in_811), .d_out(u_ca_out_811));
compressor_243_72 u_ca_243_72_812(.d_in(u_ca_in_812), .d_out(u_ca_out_812));
compressor_243_72 u_ca_243_72_813(.d_in(u_ca_in_813), .d_out(u_ca_out_813));
compressor_243_72 u_ca_243_72_814(.d_in(u_ca_in_814), .d_out(u_ca_out_814));
compressor_243_72 u_ca_243_72_815(.d_in(u_ca_in_815), .d_out(u_ca_out_815));
compressor_243_72 u_ca_243_72_816(.d_in(u_ca_in_816), .d_out(u_ca_out_816));
compressor_243_72 u_ca_243_72_817(.d_in(u_ca_in_817), .d_out(u_ca_out_817));
compressor_243_72 u_ca_243_72_818(.d_in(u_ca_in_818), .d_out(u_ca_out_818));
compressor_243_72 u_ca_243_72_819(.d_in(u_ca_in_819), .d_out(u_ca_out_819));
compressor_243_72 u_ca_243_72_820(.d_in(u_ca_in_820), .d_out(u_ca_out_820));
compressor_243_72 u_ca_243_72_821(.d_in(u_ca_in_821), .d_out(u_ca_out_821));
compressor_243_72 u_ca_243_72_822(.d_in(u_ca_in_822), .d_out(u_ca_out_822));
compressor_243_72 u_ca_243_72_823(.d_in(u_ca_in_823), .d_out(u_ca_out_823));
compressor_243_72 u_ca_243_72_824(.d_in(u_ca_in_824), .d_out(u_ca_out_824));
compressor_243_72 u_ca_243_72_825(.d_in(u_ca_in_825), .d_out(u_ca_out_825));
compressor_243_72 u_ca_243_72_826(.d_in(u_ca_in_826), .d_out(u_ca_out_826));
compressor_243_72 u_ca_243_72_827(.d_in(u_ca_in_827), .d_out(u_ca_out_827));
compressor_243_72 u_ca_243_72_828(.d_in(u_ca_in_828), .d_out(u_ca_out_828));
compressor_243_72 u_ca_243_72_829(.d_in(u_ca_in_829), .d_out(u_ca_out_829));
compressor_243_72 u_ca_243_72_830(.d_in(u_ca_in_830), .d_out(u_ca_out_830));
compressor_243_72 u_ca_243_72_831(.d_in(u_ca_in_831), .d_out(u_ca_out_831));
compressor_243_72 u_ca_243_72_832(.d_in(u_ca_in_832), .d_out(u_ca_out_832));
compressor_243_72 u_ca_243_72_833(.d_in(u_ca_in_833), .d_out(u_ca_out_833));
compressor_243_72 u_ca_243_72_834(.d_in(u_ca_in_834), .d_out(u_ca_out_834));
compressor_243_72 u_ca_243_72_835(.d_in(u_ca_in_835), .d_out(u_ca_out_835));
compressor_243_72 u_ca_243_72_836(.d_in(u_ca_in_836), .d_out(u_ca_out_836));
compressor_243_72 u_ca_243_72_837(.d_in(u_ca_in_837), .d_out(u_ca_out_837));
compressor_243_72 u_ca_243_72_838(.d_in(u_ca_in_838), .d_out(u_ca_out_838));
compressor_243_72 u_ca_243_72_839(.d_in(u_ca_in_839), .d_out(u_ca_out_839));
compressor_243_72 u_ca_243_72_840(.d_in(u_ca_in_840), .d_out(u_ca_out_840));
compressor_243_72 u_ca_243_72_841(.d_in(u_ca_in_841), .d_out(u_ca_out_841));
compressor_243_72 u_ca_243_72_842(.d_in(u_ca_in_842), .d_out(u_ca_out_842));
compressor_243_72 u_ca_243_72_843(.d_in(u_ca_in_843), .d_out(u_ca_out_843));
compressor_243_72 u_ca_243_72_844(.d_in(u_ca_in_844), .d_out(u_ca_out_844));
compressor_243_72 u_ca_243_72_845(.d_in(u_ca_in_845), .d_out(u_ca_out_845));
compressor_243_72 u_ca_243_72_846(.d_in(u_ca_in_846), .d_out(u_ca_out_846));
compressor_243_72 u_ca_243_72_847(.d_in(u_ca_in_847), .d_out(u_ca_out_847));
compressor_243_72 u_ca_243_72_848(.d_in(u_ca_in_848), .d_out(u_ca_out_848));
compressor_243_72 u_ca_243_72_849(.d_in(u_ca_in_849), .d_out(u_ca_out_849));
compressor_243_72 u_ca_243_72_850(.d_in(u_ca_in_850), .d_out(u_ca_out_850));
compressor_243_72 u_ca_243_72_851(.d_in(u_ca_in_851), .d_out(u_ca_out_851));
compressor_243_72 u_ca_243_72_852(.d_in(u_ca_in_852), .d_out(u_ca_out_852));
compressor_243_72 u_ca_243_72_853(.d_in(u_ca_in_853), .d_out(u_ca_out_853));
compressor_243_72 u_ca_243_72_854(.d_in(u_ca_in_854), .d_out(u_ca_out_854));
compressor_243_72 u_ca_243_72_855(.d_in(u_ca_in_855), .d_out(u_ca_out_855));
compressor_243_72 u_ca_243_72_856(.d_in(u_ca_in_856), .d_out(u_ca_out_856));
compressor_243_72 u_ca_243_72_857(.d_in(u_ca_in_857), .d_out(u_ca_out_857));
compressor_243_72 u_ca_243_72_858(.d_in(u_ca_in_858), .d_out(u_ca_out_858));
compressor_243_72 u_ca_243_72_859(.d_in(u_ca_in_859), .d_out(u_ca_out_859));
compressor_243_72 u_ca_243_72_860(.d_in(u_ca_in_860), .d_out(u_ca_out_860));
compressor_243_72 u_ca_243_72_861(.d_in(u_ca_in_861), .d_out(u_ca_out_861));
compressor_243_72 u_ca_243_72_862(.d_in(u_ca_in_862), .d_out(u_ca_out_862));
compressor_243_72 u_ca_243_72_863(.d_in(u_ca_in_863), .d_out(u_ca_out_863));
compressor_243_72 u_ca_243_72_864(.d_in(u_ca_in_864), .d_out(u_ca_out_864));
compressor_243_72 u_ca_243_72_865(.d_in(u_ca_in_865), .d_out(u_ca_out_865));
compressor_243_72 u_ca_243_72_866(.d_in(u_ca_in_866), .d_out(u_ca_out_866));
compressor_243_72 u_ca_243_72_867(.d_in(u_ca_in_867), .d_out(u_ca_out_867));
compressor_243_72 u_ca_243_72_868(.d_in(u_ca_in_868), .d_out(u_ca_out_868));
compressor_243_72 u_ca_243_72_869(.d_in(u_ca_in_869), .d_out(u_ca_out_869));
compressor_243_72 u_ca_243_72_870(.d_in(u_ca_in_870), .d_out(u_ca_out_870));
compressor_243_72 u_ca_243_72_871(.d_in(u_ca_in_871), .d_out(u_ca_out_871));
compressor_243_72 u_ca_243_72_872(.d_in(u_ca_in_872), .d_out(u_ca_out_872));
compressor_243_72 u_ca_243_72_873(.d_in(u_ca_in_873), .d_out(u_ca_out_873));
compressor_243_72 u_ca_243_72_874(.d_in(u_ca_in_874), .d_out(u_ca_out_874));
compressor_243_72 u_ca_243_72_875(.d_in(u_ca_in_875), .d_out(u_ca_out_875));
compressor_243_72 u_ca_243_72_876(.d_in(u_ca_in_876), .d_out(u_ca_out_876));
compressor_243_72 u_ca_243_72_877(.d_in(u_ca_in_877), .d_out(u_ca_out_877));
compressor_243_72 u_ca_243_72_878(.d_in(u_ca_in_878), .d_out(u_ca_out_878));
compressor_243_72 u_ca_243_72_879(.d_in(u_ca_in_879), .d_out(u_ca_out_879));
compressor_243_72 u_ca_243_72_880(.d_in(u_ca_in_880), .d_out(u_ca_out_880));
compressor_243_72 u_ca_243_72_881(.d_in(u_ca_in_881), .d_out(u_ca_out_881));
compressor_243_72 u_ca_243_72_882(.d_in(u_ca_in_882), .d_out(u_ca_out_882));
compressor_243_72 u_ca_243_72_883(.d_in(u_ca_in_883), .d_out(u_ca_out_883));
compressor_243_72 u_ca_243_72_884(.d_in(u_ca_in_884), .d_out(u_ca_out_884));
compressor_243_72 u_ca_243_72_885(.d_in(u_ca_in_885), .d_out(u_ca_out_885));
compressor_243_72 u_ca_243_72_886(.d_in(u_ca_in_886), .d_out(u_ca_out_886));
compressor_243_72 u_ca_243_72_887(.d_in(u_ca_in_887), .d_out(u_ca_out_887));
compressor_243_72 u_ca_243_72_888(.d_in(u_ca_in_888), .d_out(u_ca_out_888));
compressor_243_72 u_ca_243_72_889(.d_in(u_ca_in_889), .d_out(u_ca_out_889));
compressor_243_72 u_ca_243_72_890(.d_in(u_ca_in_890), .d_out(u_ca_out_890));
compressor_243_72 u_ca_243_72_891(.d_in(u_ca_in_891), .d_out(u_ca_out_891));
compressor_243_72 u_ca_243_72_892(.d_in(u_ca_in_892), .d_out(u_ca_out_892));
compressor_243_72 u_ca_243_72_893(.d_in(u_ca_in_893), .d_out(u_ca_out_893));
compressor_243_72 u_ca_243_72_894(.d_in(u_ca_in_894), .d_out(u_ca_out_894));
compressor_243_72 u_ca_243_72_895(.d_in(u_ca_in_895), .d_out(u_ca_out_895));
compressor_243_72 u_ca_243_72_896(.d_in(u_ca_in_896), .d_out(u_ca_out_896));
compressor_243_72 u_ca_243_72_897(.d_in(u_ca_in_897), .d_out(u_ca_out_897));
compressor_243_72 u_ca_243_72_898(.d_in(u_ca_in_898), .d_out(u_ca_out_898));
compressor_243_72 u_ca_243_72_899(.d_in(u_ca_in_899), .d_out(u_ca_out_899));
compressor_243_72 u_ca_243_72_900(.d_in(u_ca_in_900), .d_out(u_ca_out_900));
compressor_243_72 u_ca_243_72_901(.d_in(u_ca_in_901), .d_out(u_ca_out_901));
compressor_243_72 u_ca_243_72_902(.d_in(u_ca_in_902), .d_out(u_ca_out_902));
compressor_243_72 u_ca_243_72_903(.d_in(u_ca_in_903), .d_out(u_ca_out_903));
compressor_243_72 u_ca_243_72_904(.d_in(u_ca_in_904), .d_out(u_ca_out_904));
compressor_243_72 u_ca_243_72_905(.d_in(u_ca_in_905), .d_out(u_ca_out_905));
compressor_243_72 u_ca_243_72_906(.d_in(u_ca_in_906), .d_out(u_ca_out_906));
compressor_243_72 u_ca_243_72_907(.d_in(u_ca_in_907), .d_out(u_ca_out_907));
compressor_243_72 u_ca_243_72_908(.d_in(u_ca_in_908), .d_out(u_ca_out_908));
compressor_243_72 u_ca_243_72_909(.d_in(u_ca_in_909), .d_out(u_ca_out_909));
compressor_243_72 u_ca_243_72_910(.d_in(u_ca_in_910), .d_out(u_ca_out_910));
compressor_243_72 u_ca_243_72_911(.d_in(u_ca_in_911), .d_out(u_ca_out_911));
compressor_243_72 u_ca_243_72_912(.d_in(u_ca_in_912), .d_out(u_ca_out_912));
compressor_243_72 u_ca_243_72_913(.d_in(u_ca_in_913), .d_out(u_ca_out_913));
compressor_243_72 u_ca_243_72_914(.d_in(u_ca_in_914), .d_out(u_ca_out_914));
compressor_243_72 u_ca_243_72_915(.d_in(u_ca_in_915), .d_out(u_ca_out_915));
compressor_243_72 u_ca_243_72_916(.d_in(u_ca_in_916), .d_out(u_ca_out_916));
compressor_243_72 u_ca_243_72_917(.d_in(u_ca_in_917), .d_out(u_ca_out_917));
compressor_243_72 u_ca_243_72_918(.d_in(u_ca_in_918), .d_out(u_ca_out_918));
compressor_243_72 u_ca_243_72_919(.d_in(u_ca_in_919), .d_out(u_ca_out_919));
compressor_243_72 u_ca_243_72_920(.d_in(u_ca_in_920), .d_out(u_ca_out_920));
compressor_243_72 u_ca_243_72_921(.d_in(u_ca_in_921), .d_out(u_ca_out_921));
compressor_243_72 u_ca_243_72_922(.d_in(u_ca_in_922), .d_out(u_ca_out_922));
compressor_243_72 u_ca_243_72_923(.d_in(u_ca_in_923), .d_out(u_ca_out_923));
compressor_243_72 u_ca_243_72_924(.d_in(u_ca_in_924), .d_out(u_ca_out_924));
compressor_243_72 u_ca_243_72_925(.d_in(u_ca_in_925), .d_out(u_ca_out_925));
compressor_243_72 u_ca_243_72_926(.d_in(u_ca_in_926), .d_out(u_ca_out_926));
compressor_243_72 u_ca_243_72_927(.d_in(u_ca_in_927), .d_out(u_ca_out_927));
compressor_243_72 u_ca_243_72_928(.d_in(u_ca_in_928), .d_out(u_ca_out_928));
compressor_243_72 u_ca_243_72_929(.d_in(u_ca_in_929), .d_out(u_ca_out_929));
compressor_243_72 u_ca_243_72_930(.d_in(u_ca_in_930), .d_out(u_ca_out_930));
compressor_243_72 u_ca_243_72_931(.d_in(u_ca_in_931), .d_out(u_ca_out_931));
compressor_243_72 u_ca_243_72_932(.d_in(u_ca_in_932), .d_out(u_ca_out_932));
compressor_243_72 u_ca_243_72_933(.d_in(u_ca_in_933), .d_out(u_ca_out_933));
compressor_243_72 u_ca_243_72_934(.d_in(u_ca_in_934), .d_out(u_ca_out_934));
compressor_243_72 u_ca_243_72_935(.d_in(u_ca_in_935), .d_out(u_ca_out_935));
compressor_243_72 u_ca_243_72_936(.d_in(u_ca_in_936), .d_out(u_ca_out_936));
compressor_243_72 u_ca_243_72_937(.d_in(u_ca_in_937), .d_out(u_ca_out_937));
compressor_243_72 u_ca_243_72_938(.d_in(u_ca_in_938), .d_out(u_ca_out_938));
compressor_243_72 u_ca_243_72_939(.d_in(u_ca_in_939), .d_out(u_ca_out_939));
compressor_243_72 u_ca_243_72_940(.d_in(u_ca_in_940), .d_out(u_ca_out_940));
compressor_243_72 u_ca_243_72_941(.d_in(u_ca_in_941), .d_out(u_ca_out_941));
compressor_243_72 u_ca_243_72_942(.d_in(u_ca_in_942), .d_out(u_ca_out_942));
compressor_243_72 u_ca_243_72_943(.d_in(u_ca_in_943), .d_out(u_ca_out_943));
compressor_243_72 u_ca_243_72_944(.d_in(u_ca_in_944), .d_out(u_ca_out_944));
compressor_243_72 u_ca_243_72_945(.d_in(u_ca_in_945), .d_out(u_ca_out_945));
compressor_243_72 u_ca_243_72_946(.d_in(u_ca_in_946), .d_out(u_ca_out_946));
compressor_243_72 u_ca_243_72_947(.d_in(u_ca_in_947), .d_out(u_ca_out_947));
compressor_243_72 u_ca_243_72_948(.d_in(u_ca_in_948), .d_out(u_ca_out_948));
compressor_243_72 u_ca_243_72_949(.d_in(u_ca_in_949), .d_out(u_ca_out_949));
compressor_243_72 u_ca_243_72_950(.d_in(u_ca_in_950), .d_out(u_ca_out_950));
compressor_243_72 u_ca_243_72_951(.d_in(u_ca_in_951), .d_out(u_ca_out_951));
compressor_243_72 u_ca_243_72_952(.d_in(u_ca_in_952), .d_out(u_ca_out_952));
compressor_243_72 u_ca_243_72_953(.d_in(u_ca_in_953), .d_out(u_ca_out_953));
compressor_243_72 u_ca_243_72_954(.d_in(u_ca_in_954), .d_out(u_ca_out_954));
compressor_243_72 u_ca_243_72_955(.d_in(u_ca_in_955), .d_out(u_ca_out_955));
compressor_243_72 u_ca_243_72_956(.d_in(u_ca_in_956), .d_out(u_ca_out_956));
compressor_243_72 u_ca_243_72_957(.d_in(u_ca_in_957), .d_out(u_ca_out_957));
compressor_243_72 u_ca_243_72_958(.d_in(u_ca_in_958), .d_out(u_ca_out_958));
compressor_243_72 u_ca_243_72_959(.d_in(u_ca_in_959), .d_out(u_ca_out_959));
compressor_243_72 u_ca_243_72_960(.d_in(u_ca_in_960), .d_out(u_ca_out_960));
compressor_243_72 u_ca_243_72_961(.d_in(u_ca_in_961), .d_out(u_ca_out_961));
compressor_243_72 u_ca_243_72_962(.d_in(u_ca_in_962), .d_out(u_ca_out_962));
compressor_243_72 u_ca_243_72_963(.d_in(u_ca_in_963), .d_out(u_ca_out_963));
compressor_243_72 u_ca_243_72_964(.d_in(u_ca_in_964), .d_out(u_ca_out_964));
compressor_243_72 u_ca_243_72_965(.d_in(u_ca_in_965), .d_out(u_ca_out_965));
compressor_243_72 u_ca_243_72_966(.d_in(u_ca_in_966), .d_out(u_ca_out_966));
compressor_243_72 u_ca_243_72_967(.d_in(u_ca_in_967), .d_out(u_ca_out_967));
compressor_243_72 u_ca_243_72_968(.d_in(u_ca_in_968), .d_out(u_ca_out_968));
compressor_243_72 u_ca_243_72_969(.d_in(u_ca_in_969), .d_out(u_ca_out_969));
compressor_243_72 u_ca_243_72_970(.d_in(u_ca_in_970), .d_out(u_ca_out_970));
compressor_243_72 u_ca_243_72_971(.d_in(u_ca_in_971), .d_out(u_ca_out_971));
compressor_243_72 u_ca_243_72_972(.d_in(u_ca_in_972), .d_out(u_ca_out_972));
compressor_243_72 u_ca_243_72_973(.d_in(u_ca_in_973), .d_out(u_ca_out_973));
compressor_243_72 u_ca_243_72_974(.d_in(u_ca_in_974), .d_out(u_ca_out_974));
compressor_243_72 u_ca_243_72_975(.d_in(u_ca_in_975), .d_out(u_ca_out_975));
compressor_243_72 u_ca_243_72_976(.d_in(u_ca_in_976), .d_out(u_ca_out_976));
compressor_243_72 u_ca_243_72_977(.d_in(u_ca_in_977), .d_out(u_ca_out_977));
compressor_243_72 u_ca_243_72_978(.d_in(u_ca_in_978), .d_out(u_ca_out_978));
compressor_243_72 u_ca_243_72_979(.d_in(u_ca_in_979), .d_out(u_ca_out_979));
compressor_243_72 u_ca_243_72_980(.d_in(u_ca_in_980), .d_out(u_ca_out_980));
compressor_243_72 u_ca_243_72_981(.d_in(u_ca_in_981), .d_out(u_ca_out_981));
compressor_243_72 u_ca_243_72_982(.d_in(u_ca_in_982), .d_out(u_ca_out_982));
compressor_243_72 u_ca_243_72_983(.d_in(u_ca_in_983), .d_out(u_ca_out_983));
compressor_243_72 u_ca_243_72_984(.d_in(u_ca_in_984), .d_out(u_ca_out_984));
compressor_243_72 u_ca_243_72_985(.d_in(u_ca_in_985), .d_out(u_ca_out_985));
compressor_243_72 u_ca_243_72_986(.d_in(u_ca_in_986), .d_out(u_ca_out_986));
compressor_243_72 u_ca_243_72_987(.d_in(u_ca_in_987), .d_out(u_ca_out_987));
compressor_243_72 u_ca_243_72_988(.d_in(u_ca_in_988), .d_out(u_ca_out_988));
compressor_243_72 u_ca_243_72_989(.d_in(u_ca_in_989), .d_out(u_ca_out_989));
compressor_243_72 u_ca_243_72_990(.d_in(u_ca_in_990), .d_out(u_ca_out_990));
compressor_243_72 u_ca_243_72_991(.d_in(u_ca_in_991), .d_out(u_ca_out_991));
compressor_243_72 u_ca_243_72_992(.d_in(u_ca_in_992), .d_out(u_ca_out_992));
compressor_243_72 u_ca_243_72_993(.d_in(u_ca_in_993), .d_out(u_ca_out_993));
compressor_243_72 u_ca_243_72_994(.d_in(u_ca_in_994), .d_out(u_ca_out_994));
compressor_243_72 u_ca_243_72_995(.d_in(u_ca_in_995), .d_out(u_ca_out_995));
compressor_243_72 u_ca_243_72_996(.d_in(u_ca_in_996), .d_out(u_ca_out_996));
compressor_243_72 u_ca_243_72_997(.d_in(u_ca_in_997), .d_out(u_ca_out_997));
compressor_243_72 u_ca_243_72_998(.d_in(u_ca_in_998), .d_out(u_ca_out_998));
compressor_243_72 u_ca_243_72_999(.d_in(u_ca_in_999), .d_out(u_ca_out_999));
compressor_243_72 u_ca_243_72_1000(.d_in(u_ca_in_1000), .d_out(u_ca_out_1000));
compressor_243_72 u_ca_243_72_1001(.d_in(u_ca_in_1001), .d_out(u_ca_out_1001));
compressor_243_72 u_ca_243_72_1002(.d_in(u_ca_in_1002), .d_out(u_ca_out_1002));
compressor_243_72 u_ca_243_72_1003(.d_in(u_ca_in_1003), .d_out(u_ca_out_1003));
compressor_243_72 u_ca_243_72_1004(.d_in(u_ca_in_1004), .d_out(u_ca_out_1004));
compressor_243_72 u_ca_243_72_1005(.d_in(u_ca_in_1005), .d_out(u_ca_out_1005));
compressor_243_72 u_ca_243_72_1006(.d_in(u_ca_in_1006), .d_out(u_ca_out_1006));
compressor_243_72 u_ca_243_72_1007(.d_in(u_ca_in_1007), .d_out(u_ca_out_1007));
compressor_243_72 u_ca_243_72_1008(.d_in(u_ca_in_1008), .d_out(u_ca_out_1008));
compressor_243_72 u_ca_243_72_1009(.d_in(u_ca_in_1009), .d_out(u_ca_out_1009));
compressor_243_72 u_ca_243_72_1010(.d_in(u_ca_in_1010), .d_out(u_ca_out_1010));
compressor_243_72 u_ca_243_72_1011(.d_in(u_ca_in_1011), .d_out(u_ca_out_1011));
compressor_243_72 u_ca_243_72_1012(.d_in(u_ca_in_1012), .d_out(u_ca_out_1012));
compressor_243_72 u_ca_243_72_1013(.d_in(u_ca_in_1013), .d_out(u_ca_out_1013));
compressor_243_72 u_ca_243_72_1014(.d_in(u_ca_in_1014), .d_out(u_ca_out_1014));
compressor_243_72 u_ca_243_72_1015(.d_in(u_ca_in_1015), .d_out(u_ca_out_1015));
compressor_243_72 u_ca_243_72_1016(.d_in(u_ca_in_1016), .d_out(u_ca_out_1016));
compressor_243_72 u_ca_243_72_1017(.d_in(u_ca_in_1017), .d_out(u_ca_out_1017));
compressor_243_72 u_ca_243_72_1018(.d_in(u_ca_in_1018), .d_out(u_ca_out_1018));
compressor_243_72 u_ca_243_72_1019(.d_in(u_ca_in_1019), .d_out(u_ca_out_1019));
compressor_243_72 u_ca_243_72_1020(.d_in(u_ca_in_1020), .d_out(u_ca_out_1020));
compressor_243_72 u_ca_243_72_1021(.d_in(u_ca_in_1021), .d_out(u_ca_out_1021));
compressor_243_72 u_ca_243_72_1022(.d_in(u_ca_in_1022), .d_out(u_ca_out_1022));
compressor_243_72 u_ca_243_72_1023(.d_in(u_ca_in_1023), .d_out(u_ca_out_1023));
compressor_243_72 u_ca_243_72_1024(.d_in(u_ca_in_1024), .d_out(u_ca_out_1024));
compressor_243_72 u_ca_243_72_1025(.d_in(u_ca_in_1025), .d_out(u_ca_out_1025));
compressor_243_72 u_ca_243_72_1026(.d_in(u_ca_in_1026), .d_out(u_ca_out_1026));
compressor_243_72 u_ca_243_72_1027(.d_in(u_ca_in_1027), .d_out(u_ca_out_1027));
compressor_243_72 u_ca_243_72_1028(.d_in(u_ca_in_1028), .d_out(u_ca_out_1028));
compressor_243_72 u_ca_243_72_1029(.d_in(u_ca_in_1029), .d_out(u_ca_out_1029));
compressor_243_72 u_ca_243_72_1030(.d_in(u_ca_in_1030), .d_out(u_ca_out_1030));
compressor_243_72 u_ca_243_72_1031(.d_in(u_ca_in_1031), .d_out(u_ca_out_1031));
compressor_243_72 u_ca_243_72_1032(.d_in(u_ca_in_1032), .d_out(u_ca_out_1032));
compressor_243_72 u_ca_243_72_1033(.d_in(u_ca_in_1033), .d_out(u_ca_out_1033));
compressor_243_72 u_ca_243_72_1034(.d_in(u_ca_in_1034), .d_out(u_ca_out_1034));
compressor_243_72 u_ca_243_72_1035(.d_in(u_ca_in_1035), .d_out(u_ca_out_1035));
compressor_243_72 u_ca_243_72_1036(.d_in(u_ca_in_1036), .d_out(u_ca_out_1036));
compressor_243_72 u_ca_243_72_1037(.d_in(u_ca_in_1037), .d_out(u_ca_out_1037));
compressor_243_72 u_ca_243_72_1038(.d_in(u_ca_in_1038), .d_out(u_ca_out_1038));
compressor_243_72 u_ca_243_72_1039(.d_in(u_ca_in_1039), .d_out(u_ca_out_1039));
compressor_243_72 u_ca_243_72_1040(.d_in(u_ca_in_1040), .d_out(u_ca_out_1040));
compressor_243_72 u_ca_243_72_1041(.d_in(u_ca_in_1041), .d_out(u_ca_out_1041));
compressor_243_72 u_ca_243_72_1042(.d_in(u_ca_in_1042), .d_out(u_ca_out_1042));
compressor_243_72 u_ca_243_72_1043(.d_in(u_ca_in_1043), .d_out(u_ca_out_1043));
compressor_243_72 u_ca_243_72_1044(.d_in(u_ca_in_1044), .d_out(u_ca_out_1044));
compressor_243_72 u_ca_243_72_1045(.d_in(u_ca_in_1045), .d_out(u_ca_out_1045));
compressor_243_72 u_ca_243_72_1046(.d_in(u_ca_in_1046), .d_out(u_ca_out_1046));
compressor_243_72 u_ca_243_72_1047(.d_in(u_ca_in_1047), .d_out(u_ca_out_1047));
compressor_243_72 u_ca_243_72_1048(.d_in(u_ca_in_1048), .d_out(u_ca_out_1048));
compressor_243_72 u_ca_243_72_1049(.d_in(u_ca_in_1049), .d_out(u_ca_out_1049));
compressor_243_72 u_ca_243_72_1050(.d_in(u_ca_in_1050), .d_out(u_ca_out_1050));
compressor_243_72 u_ca_243_72_1051(.d_in(u_ca_in_1051), .d_out(u_ca_out_1051));
compressor_243_72 u_ca_243_72_1052(.d_in(u_ca_in_1052), .d_out(u_ca_out_1052));
compressor_243_72 u_ca_243_72_1053(.d_in(u_ca_in_1053), .d_out(u_ca_out_1053));
compressor_243_72 u_ca_243_72_1054(.d_in(u_ca_in_1054), .d_out(u_ca_out_1054));
compressor_243_72 u_ca_243_72_1055(.d_in(u_ca_in_1055), .d_out(u_ca_out_1055));
compressor_243_72 u_ca_243_72_1056(.d_in(u_ca_in_1056), .d_out(u_ca_out_1056));
compressor_243_72 u_ca_243_72_1057(.d_in(u_ca_in_1057), .d_out(u_ca_out_1057));
compressor_243_72 u_ca_243_72_1058(.d_in(u_ca_in_1058), .d_out(u_ca_out_1058));
compressor_243_72 u_ca_243_72_1059(.d_in(u_ca_in_1059), .d_out(u_ca_out_1059));
compressor_243_72 u_ca_243_72_1060(.d_in(u_ca_in_1060), .d_out(u_ca_out_1060));
compressor_243_72 u_ca_243_72_1061(.d_in(u_ca_in_1061), .d_out(u_ca_out_1061));
compressor_243_72 u_ca_243_72_1062(.d_in(u_ca_in_1062), .d_out(u_ca_out_1062));
compressor_243_72 u_ca_243_72_1063(.d_in(u_ca_in_1063), .d_out(u_ca_out_1063));
compressor_243_72 u_ca_243_72_1064(.d_in(u_ca_in_1064), .d_out(u_ca_out_1064));
compressor_243_72 u_ca_243_72_1065(.d_in(u_ca_in_1065), .d_out(u_ca_out_1065));
compressor_243_72 u_ca_243_72_1066(.d_in(u_ca_in_1066), .d_out(u_ca_out_1066));
compressor_243_72 u_ca_243_72_1067(.d_in(u_ca_in_1067), .d_out(u_ca_out_1067));
compressor_243_72 u_ca_243_72_1068(.d_in(u_ca_in_1068), .d_out(u_ca_out_1068));
compressor_243_72 u_ca_243_72_1069(.d_in(u_ca_in_1069), .d_out(u_ca_out_1069));
compressor_243_72 u_ca_243_72_1070(.d_in(u_ca_in_1070), .d_out(u_ca_out_1070));
compressor_243_72 u_ca_243_72_1071(.d_in(u_ca_in_1071), .d_out(u_ca_out_1071));
compressor_243_72 u_ca_243_72_1072(.d_in(u_ca_in_1072), .d_out(u_ca_out_1072));
compressor_243_72 u_ca_243_72_1073(.d_in(u_ca_in_1073), .d_out(u_ca_out_1073));
compressor_243_72 u_ca_243_72_1074(.d_in(u_ca_in_1074), .d_out(u_ca_out_1074));
compressor_243_72 u_ca_243_72_1075(.d_in(u_ca_in_1075), .d_out(u_ca_out_1075));
compressor_243_72 u_ca_243_72_1076(.d_in(u_ca_in_1076), .d_out(u_ca_out_1076));
compressor_243_72 u_ca_243_72_1077(.d_in(u_ca_in_1077), .d_out(u_ca_out_1077));
compressor_243_72 u_ca_243_72_1078(.d_in(u_ca_in_1078), .d_out(u_ca_out_1078));
compressor_243_72 u_ca_243_72_1079(.d_in(u_ca_in_1079), .d_out(u_ca_out_1079));
compressor_243_72 u_ca_243_72_1080(.d_in(u_ca_in_1080), .d_out(u_ca_out_1080));
compressor_243_72 u_ca_243_72_1081(.d_in(u_ca_in_1081), .d_out(u_ca_out_1081));
compressor_243_72 u_ca_243_72_1082(.d_in(u_ca_in_1082), .d_out(u_ca_out_1082));
compressor_243_72 u_ca_243_72_1083(.d_in(u_ca_in_1083), .d_out(u_ca_out_1083));
compressor_243_72 u_ca_243_72_1084(.d_in(u_ca_in_1084), .d_out(u_ca_out_1084));
compressor_243_72 u_ca_243_72_1085(.d_in(u_ca_in_1085), .d_out(u_ca_out_1085));
compressor_243_72 u_ca_243_72_1086(.d_in(u_ca_in_1086), .d_out(u_ca_out_1086));
compressor_243_72 u_ca_243_72_1087(.d_in(u_ca_in_1087), .d_out(u_ca_out_1087));
compressor_243_72 u_ca_243_72_1088(.d_in(u_ca_in_1088), .d_out(u_ca_out_1088));
compressor_243_72 u_ca_243_72_1089(.d_in(u_ca_in_1089), .d_out(u_ca_out_1089));
compressor_243_72 u_ca_243_72_1090(.d_in(u_ca_in_1090), .d_out(u_ca_out_1090));
compressor_243_72 u_ca_243_72_1091(.d_in(u_ca_in_1091), .d_out(u_ca_out_1091));
compressor_243_72 u_ca_243_72_1092(.d_in(u_ca_in_1092), .d_out(u_ca_out_1092));
compressor_243_72 u_ca_243_72_1093(.d_in(u_ca_in_1093), .d_out(u_ca_out_1093));
compressor_243_72 u_ca_243_72_1094(.d_in(u_ca_in_1094), .d_out(u_ca_out_1094));
compressor_243_72 u_ca_243_72_1095(.d_in(u_ca_in_1095), .d_out(u_ca_out_1095));
compressor_243_72 u_ca_243_72_1096(.d_in(u_ca_in_1096), .d_out(u_ca_out_1096));
compressor_243_72 u_ca_243_72_1097(.d_in(u_ca_in_1097), .d_out(u_ca_out_1097));
compressor_243_72 u_ca_243_72_1098(.d_in(u_ca_in_1098), .d_out(u_ca_out_1098));
compressor_243_72 u_ca_243_72_1099(.d_in(u_ca_in_1099), .d_out(u_ca_out_1099));
compressor_243_72 u_ca_243_72_1100(.d_in(u_ca_in_1100), .d_out(u_ca_out_1100));
compressor_243_72 u_ca_243_72_1101(.d_in(u_ca_in_1101), .d_out(u_ca_out_1101));
compressor_243_72 u_ca_243_72_1102(.d_in(u_ca_in_1102), .d_out(u_ca_out_1102));
compressor_243_72 u_ca_243_72_1103(.d_in(u_ca_in_1103), .d_out(u_ca_out_1103));
compressor_243_72 u_ca_243_72_1104(.d_in(u_ca_in_1104), .d_out(u_ca_out_1104));
compressor_243_72 u_ca_243_72_1105(.d_in(u_ca_in_1105), .d_out(u_ca_out_1105));
compressor_243_72 u_ca_243_72_1106(.d_in(u_ca_in_1106), .d_out(u_ca_out_1106));
compressor_243_72 u_ca_243_72_1107(.d_in(u_ca_in_1107), .d_out(u_ca_out_1107));
compressor_243_72 u_ca_243_72_1108(.d_in(u_ca_in_1108), .d_out(u_ca_out_1108));
compressor_243_72 u_ca_243_72_1109(.d_in(u_ca_in_1109), .d_out(u_ca_out_1109));
compressor_243_72 u_ca_243_72_1110(.d_in(u_ca_in_1110), .d_out(u_ca_out_1110));
compressor_243_72 u_ca_243_72_1111(.d_in(u_ca_in_1111), .d_out(u_ca_out_1111));
compressor_243_72 u_ca_243_72_1112(.d_in(u_ca_in_1112), .d_out(u_ca_out_1112));
compressor_243_72 u_ca_243_72_1113(.d_in(u_ca_in_1113), .d_out(u_ca_out_1113));
compressor_243_72 u_ca_243_72_1114(.d_in(u_ca_in_1114), .d_out(u_ca_out_1114));
compressor_243_72 u_ca_243_72_1115(.d_in(u_ca_in_1115), .d_out(u_ca_out_1115));
compressor_243_72 u_ca_243_72_1116(.d_in(u_ca_in_1116), .d_out(u_ca_out_1116));
compressor_243_72 u_ca_243_72_1117(.d_in(u_ca_in_1117), .d_out(u_ca_out_1117));
compressor_243_72 u_ca_243_72_1118(.d_in(u_ca_in_1118), .d_out(u_ca_out_1118));
compressor_243_72 u_ca_243_72_1119(.d_in(u_ca_in_1119), .d_out(u_ca_out_1119));
compressor_243_72 u_ca_243_72_1120(.d_in(u_ca_in_1120), .d_out(u_ca_out_1120));
compressor_243_72 u_ca_243_72_1121(.d_in(u_ca_in_1121), .d_out(u_ca_out_1121));
compressor_243_72 u_ca_243_72_1122(.d_in(u_ca_in_1122), .d_out(u_ca_out_1122));
compressor_243_72 u_ca_243_72_1123(.d_in(u_ca_in_1123), .d_out(u_ca_out_1123));
compressor_243_72 u_ca_243_72_1124(.d_in(u_ca_in_1124), .d_out(u_ca_out_1124));
compressor_243_72 u_ca_243_72_1125(.d_in(u_ca_in_1125), .d_out(u_ca_out_1125));
compressor_243_72 u_ca_243_72_1126(.d_in(u_ca_in_1126), .d_out(u_ca_out_1126));
compressor_243_72 u_ca_243_72_1127(.d_in(u_ca_in_1127), .d_out(u_ca_out_1127));
compressor_243_72 u_ca_243_72_1128(.d_in(u_ca_in_1128), .d_out(u_ca_out_1128));
compressor_243_72 u_ca_243_72_1129(.d_in(u_ca_in_1129), .d_out(u_ca_out_1129));
compressor_243_72 u_ca_243_72_1130(.d_in(u_ca_in_1130), .d_out(u_ca_out_1130));
compressor_243_72 u_ca_243_72_1131(.d_in(u_ca_in_1131), .d_out(u_ca_out_1131));
compressor_243_72 u_ca_243_72_1132(.d_in(u_ca_in_1132), .d_out(u_ca_out_1132));
compressor_243_72 u_ca_243_72_1133(.d_in(u_ca_in_1133), .d_out(u_ca_out_1133));
compressor_243_72 u_ca_243_72_1134(.d_in(u_ca_in_1134), .d_out(u_ca_out_1134));
compressor_243_72 u_ca_243_72_1135(.d_in(u_ca_in_1135), .d_out(u_ca_out_1135));
compressor_243_72 u_ca_243_72_1136(.d_in(u_ca_in_1136), .d_out(u_ca_out_1136));
compressor_243_72 u_ca_243_72_1137(.d_in(u_ca_in_1137), .d_out(u_ca_out_1137));
compressor_243_72 u_ca_243_72_1138(.d_in(u_ca_in_1138), .d_out(u_ca_out_1138));
compressor_243_72 u_ca_243_72_1139(.d_in(u_ca_in_1139), .d_out(u_ca_out_1139));
compressor_243_72 u_ca_243_72_1140(.d_in(u_ca_in_1140), .d_out(u_ca_out_1140));
compressor_243_72 u_ca_243_72_1141(.d_in(u_ca_in_1141), .d_out(u_ca_out_1141));
compressor_243_72 u_ca_243_72_1142(.d_in(u_ca_in_1142), .d_out(u_ca_out_1142));
compressor_243_72 u_ca_243_72_1143(.d_in(u_ca_in_1143), .d_out(u_ca_out_1143));
compressor_243_72 u_ca_243_72_1144(.d_in(u_ca_in_1144), .d_out(u_ca_out_1144));
compressor_243_72 u_ca_243_72_1145(.d_in(u_ca_in_1145), .d_out(u_ca_out_1145));
compressor_243_72 u_ca_243_72_1146(.d_in(u_ca_in_1146), .d_out(u_ca_out_1146));
compressor_243_72 u_ca_243_72_1147(.d_in(u_ca_in_1147), .d_out(u_ca_out_1147));
compressor_243_72 u_ca_243_72_1148(.d_in(u_ca_in_1148), .d_out(u_ca_out_1148));
compressor_243_72 u_ca_243_72_1149(.d_in(u_ca_in_1149), .d_out(u_ca_out_1149));
compressor_243_72 u_ca_243_72_1150(.d_in(u_ca_in_1150), .d_out(u_ca_out_1150));
compressor_243_72 u_ca_243_72_1151(.d_in(u_ca_in_1151), .d_out(u_ca_out_1151));
compressor_243_72 u_ca_243_72_1152(.d_in(u_ca_in_1152), .d_out(u_ca_out_1152));
compressor_243_72 u_ca_243_72_1153(.d_in(u_ca_in_1153), .d_out(u_ca_out_1153));
compressor_243_72 u_ca_243_72_1154(.d_in(u_ca_in_1154), .d_out(u_ca_out_1154));
compressor_243_72 u_ca_243_72_1155(.d_in(u_ca_in_1155), .d_out(u_ca_out_1155));
compressor_243_72 u_ca_243_72_1156(.d_in(u_ca_in_1156), .d_out(u_ca_out_1156));
compressor_243_72 u_ca_243_72_1157(.d_in(u_ca_in_1157), .d_out(u_ca_out_1157));
compressor_243_72 u_ca_243_72_1158(.d_in(u_ca_in_1158), .d_out(u_ca_out_1158));
compressor_243_72 u_ca_243_72_1159(.d_in(u_ca_in_1159), .d_out(u_ca_out_1159));
compressor_243_72 u_ca_243_72_1160(.d_in(u_ca_in_1160), .d_out(u_ca_out_1160));
compressor_243_72 u_ca_243_72_1161(.d_in(u_ca_in_1161), .d_out(u_ca_out_1161));
compressor_243_72 u_ca_243_72_1162(.d_in(u_ca_in_1162), .d_out(u_ca_out_1162));
compressor_243_72 u_ca_243_72_1163(.d_in(u_ca_in_1163), .d_out(u_ca_out_1163));
compressor_243_72 u_ca_243_72_1164(.d_in(u_ca_in_1164), .d_out(u_ca_out_1164));
compressor_243_72 u_ca_243_72_1165(.d_in(u_ca_in_1165), .d_out(u_ca_out_1165));
compressor_243_72 u_ca_243_72_1166(.d_in(u_ca_in_1166), .d_out(u_ca_out_1166));
compressor_243_72 u_ca_243_72_1167(.d_in(u_ca_in_1167), .d_out(u_ca_out_1167));
compressor_243_72 u_ca_243_72_1168(.d_in(u_ca_in_1168), .d_out(u_ca_out_1168));
compressor_243_72 u_ca_243_72_1169(.d_in(u_ca_in_1169), .d_out(u_ca_out_1169));
compressor_243_72 u_ca_243_72_1170(.d_in(u_ca_in_1170), .d_out(u_ca_out_1170));
compressor_243_72 u_ca_243_72_1171(.d_in(u_ca_in_1171), .d_out(u_ca_out_1171));
compressor_243_72 u_ca_243_72_1172(.d_in(u_ca_in_1172), .d_out(u_ca_out_1172));
compressor_243_72 u_ca_243_72_1173(.d_in(u_ca_in_1173), .d_out(u_ca_out_1173));
compressor_243_72 u_ca_243_72_1174(.d_in(u_ca_in_1174), .d_out(u_ca_out_1174));
compressor_243_72 u_ca_243_72_1175(.d_in(u_ca_in_1175), .d_out(u_ca_out_1175));
compressor_243_72 u_ca_243_72_1176(.d_in(u_ca_in_1176), .d_out(u_ca_out_1176));
compressor_243_72 u_ca_243_72_1177(.d_in(u_ca_in_1177), .d_out(u_ca_out_1177));
compressor_243_72 u_ca_243_72_1178(.d_in(u_ca_in_1178), .d_out(u_ca_out_1178));
compressor_243_72 u_ca_243_72_1179(.d_in(u_ca_in_1179), .d_out(u_ca_out_1179));
compressor_243_72 u_ca_243_72_1180(.d_in(u_ca_in_1180), .d_out(u_ca_out_1180));
compressor_243_72 u_ca_243_72_1181(.d_in(u_ca_in_1181), .d_out(u_ca_out_1181));
compressor_243_72 u_ca_243_72_1182(.d_in(u_ca_in_1182), .d_out(u_ca_out_1182));
compressor_243_72 u_ca_243_72_1183(.d_in(u_ca_in_1183), .d_out(u_ca_out_1183));
compressor_243_72 u_ca_243_72_1184(.d_in(u_ca_in_1184), .d_out(u_ca_out_1184));
compressor_243_72 u_ca_243_72_1185(.d_in(u_ca_in_1185), .d_out(u_ca_out_1185));
compressor_243_72 u_ca_243_72_1186(.d_in(u_ca_in_1186), .d_out(u_ca_out_1186));
compressor_243_72 u_ca_243_72_1187(.d_in(u_ca_in_1187), .d_out(u_ca_out_1187));
compressor_243_72 u_ca_243_72_1188(.d_in(u_ca_in_1188), .d_out(u_ca_out_1188));
compressor_243_72 u_ca_243_72_1189(.d_in(u_ca_in_1189), .d_out(u_ca_out_1189));
compressor_243_72 u_ca_243_72_1190(.d_in(u_ca_in_1190), .d_out(u_ca_out_1190));
compressor_243_72 u_ca_243_72_1191(.d_in(u_ca_in_1191), .d_out(u_ca_out_1191));
compressor_243_72 u_ca_243_72_1192(.d_in(u_ca_in_1192), .d_out(u_ca_out_1192));
compressor_243_72 u_ca_243_72_1193(.d_in(u_ca_in_1193), .d_out(u_ca_out_1193));
compressor_243_72 u_ca_243_72_1194(.d_in(u_ca_in_1194), .d_out(u_ca_out_1194));
compressor_243_72 u_ca_243_72_1195(.d_in(u_ca_in_1195), .d_out(u_ca_out_1195));
compressor_243_72 u_ca_243_72_1196(.d_in(u_ca_in_1196), .d_out(u_ca_out_1196));
compressor_243_72 u_ca_243_72_1197(.d_in(u_ca_in_1197), .d_out(u_ca_out_1197));
compressor_243_72 u_ca_243_72_1198(.d_in(u_ca_in_1198), .d_out(u_ca_out_1198));
compressor_243_72 u_ca_243_72_1199(.d_in(u_ca_in_1199), .d_out(u_ca_out_1199));
compressor_243_72 u_ca_243_72_1200(.d_in(u_ca_in_1200), .d_out(u_ca_out_1200));
compressor_243_72 u_ca_243_72_1201(.d_in(u_ca_in_1201), .d_out(u_ca_out_1201));
compressor_243_72 u_ca_243_72_1202(.d_in(u_ca_in_1202), .d_out(u_ca_out_1202));
compressor_243_72 u_ca_243_72_1203(.d_in(u_ca_in_1203), .d_out(u_ca_out_1203));
compressor_243_72 u_ca_243_72_1204(.d_in(u_ca_in_1204), .d_out(u_ca_out_1204));
compressor_243_72 u_ca_243_72_1205(.d_in(u_ca_in_1205), .d_out(u_ca_out_1205));
compressor_243_72 u_ca_243_72_1206(.d_in(u_ca_in_1206), .d_out(u_ca_out_1206));
compressor_243_72 u_ca_243_72_1207(.d_in(u_ca_in_1207), .d_out(u_ca_out_1207));
compressor_243_72 u_ca_243_72_1208(.d_in(u_ca_in_1208), .d_out(u_ca_out_1208));
compressor_243_72 u_ca_243_72_1209(.d_in(u_ca_in_1209), .d_out(u_ca_out_1209));
compressor_243_72 u_ca_243_72_1210(.d_in(u_ca_in_1210), .d_out(u_ca_out_1210));
compressor_243_72 u_ca_243_72_1211(.d_in(u_ca_in_1211), .d_out(u_ca_out_1211));
compressor_243_72 u_ca_243_72_1212(.d_in(u_ca_in_1212), .d_out(u_ca_out_1212));
compressor_243_72 u_ca_243_72_1213(.d_in(u_ca_in_1213), .d_out(u_ca_out_1213));
compressor_243_72 u_ca_243_72_1214(.d_in(u_ca_in_1214), .d_out(u_ca_out_1214));
compressor_243_72 u_ca_243_72_1215(.d_in(u_ca_in_1215), .d_out(u_ca_out_1215));
compressor_243_72 u_ca_243_72_1216(.d_in(u_ca_in_1216), .d_out(u_ca_out_1216));
compressor_243_72 u_ca_243_72_1217(.d_in(u_ca_in_1217), .d_out(u_ca_out_1217));
compressor_243_72 u_ca_243_72_1218(.d_in(u_ca_in_1218), .d_out(u_ca_out_1218));
compressor_243_72 u_ca_243_72_1219(.d_in(u_ca_in_1219), .d_out(u_ca_out_1219));
compressor_243_72 u_ca_243_72_1220(.d_in(u_ca_in_1220), .d_out(u_ca_out_1220));
compressor_243_72 u_ca_243_72_1221(.d_in(u_ca_in_1221), .d_out(u_ca_out_1221));
compressor_243_72 u_ca_243_72_1222(.d_in(u_ca_in_1222), .d_out(u_ca_out_1222));
compressor_243_72 u_ca_243_72_1223(.d_in(u_ca_in_1223), .d_out(u_ca_out_1223));
compressor_243_72 u_ca_243_72_1224(.d_in(u_ca_in_1224), .d_out(u_ca_out_1224));
compressor_243_72 u_ca_243_72_1225(.d_in(u_ca_in_1225), .d_out(u_ca_out_1225));
compressor_243_72 u_ca_243_72_1226(.d_in(u_ca_in_1226), .d_out(u_ca_out_1226));
compressor_243_72 u_ca_243_72_1227(.d_in(u_ca_in_1227), .d_out(u_ca_out_1227));
compressor_243_72 u_ca_243_72_1228(.d_in(u_ca_in_1228), .d_out(u_ca_out_1228));
compressor_243_72 u_ca_243_72_1229(.d_in(u_ca_in_1229), .d_out(u_ca_out_1229));
compressor_243_72 u_ca_243_72_1230(.d_in(u_ca_in_1230), .d_out(u_ca_out_1230));
compressor_243_72 u_ca_243_72_1231(.d_in(u_ca_in_1231), .d_out(u_ca_out_1231));
compressor_243_72 u_ca_243_72_1232(.d_in(u_ca_in_1232), .d_out(u_ca_out_1232));
compressor_243_72 u_ca_243_72_1233(.d_in(u_ca_in_1233), .d_out(u_ca_out_1233));
compressor_243_72 u_ca_243_72_1234(.d_in(u_ca_in_1234), .d_out(u_ca_out_1234));
compressor_243_72 u_ca_243_72_1235(.d_in(u_ca_in_1235), .d_out(u_ca_out_1235));
compressor_243_72 u_ca_243_72_1236(.d_in(u_ca_in_1236), .d_out(u_ca_out_1236));
compressor_243_72 u_ca_243_72_1237(.d_in(u_ca_in_1237), .d_out(u_ca_out_1237));
compressor_243_72 u_ca_243_72_1238(.d_in(u_ca_in_1238), .d_out(u_ca_out_1238));
compressor_243_72 u_ca_243_72_1239(.d_in(u_ca_in_1239), .d_out(u_ca_out_1239));
compressor_243_72 u_ca_243_72_1240(.d_in(u_ca_in_1240), .d_out(u_ca_out_1240));
compressor_243_72 u_ca_243_72_1241(.d_in(u_ca_in_1241), .d_out(u_ca_out_1241));
compressor_243_72 u_ca_243_72_1242(.d_in(u_ca_in_1242), .d_out(u_ca_out_1242));
compressor_243_72 u_ca_243_72_1243(.d_in(u_ca_in_1243), .d_out(u_ca_out_1243));
compressor_243_72 u_ca_243_72_1244(.d_in(u_ca_in_1244), .d_out(u_ca_out_1244));
compressor_243_72 u_ca_243_72_1245(.d_in(u_ca_in_1245), .d_out(u_ca_out_1245));
compressor_243_72 u_ca_243_72_1246(.d_in(u_ca_in_1246), .d_out(u_ca_out_1246));
compressor_243_72 u_ca_243_72_1247(.d_in(u_ca_in_1247), .d_out(u_ca_out_1247));
compressor_243_72 u_ca_243_72_1248(.d_in(u_ca_in_1248), .d_out(u_ca_out_1248));
compressor_243_72 u_ca_243_72_1249(.d_in(u_ca_in_1249), .d_out(u_ca_out_1249));
compressor_243_72 u_ca_243_72_1250(.d_in(u_ca_in_1250), .d_out(u_ca_out_1250));
compressor_243_72 u_ca_243_72_1251(.d_in(u_ca_in_1251), .d_out(u_ca_out_1251));
compressor_243_72 u_ca_243_72_1252(.d_in(u_ca_in_1252), .d_out(u_ca_out_1252));
compressor_243_72 u_ca_243_72_1253(.d_in(u_ca_in_1253), .d_out(u_ca_out_1253));
compressor_243_72 u_ca_243_72_1254(.d_in(u_ca_in_1254), .d_out(u_ca_out_1254));
compressor_243_72 u_ca_243_72_1255(.d_in(u_ca_in_1255), .d_out(u_ca_out_1255));
compressor_243_72 u_ca_243_72_1256(.d_in(u_ca_in_1256), .d_out(u_ca_out_1256));
compressor_243_72 u_ca_243_72_1257(.d_in(u_ca_in_1257), .d_out(u_ca_out_1257));
compressor_243_72 u_ca_243_72_1258(.d_in(u_ca_in_1258), .d_out(u_ca_out_1258));
compressor_243_72 u_ca_243_72_1259(.d_in(u_ca_in_1259), .d_out(u_ca_out_1259));
compressor_243_72 u_ca_243_72_1260(.d_in(u_ca_in_1260), .d_out(u_ca_out_1260));
compressor_243_72 u_ca_243_72_1261(.d_in(u_ca_in_1261), .d_out(u_ca_out_1261));
compressor_243_72 u_ca_243_72_1262(.d_in(u_ca_in_1262), .d_out(u_ca_out_1262));
compressor_243_72 u_ca_243_72_1263(.d_in(u_ca_in_1263), .d_out(u_ca_out_1263));
compressor_243_72 u_ca_243_72_1264(.d_in(u_ca_in_1264), .d_out(u_ca_out_1264));
compressor_243_72 u_ca_243_72_1265(.d_in(u_ca_in_1265), .d_out(u_ca_out_1265));
compressor_243_72 u_ca_243_72_1266(.d_in(u_ca_in_1266), .d_out(u_ca_out_1266));
compressor_243_72 u_ca_243_72_1267(.d_in(u_ca_in_1267), .d_out(u_ca_out_1267));
compressor_243_72 u_ca_243_72_1268(.d_in(u_ca_in_1268), .d_out(u_ca_out_1268));
compressor_243_72 u_ca_243_72_1269(.d_in(u_ca_in_1269), .d_out(u_ca_out_1269));
compressor_243_72 u_ca_243_72_1270(.d_in(u_ca_in_1270), .d_out(u_ca_out_1270));
compressor_243_72 u_ca_243_72_1271(.d_in(u_ca_in_1271), .d_out(u_ca_out_1271));
compressor_243_72 u_ca_243_72_1272(.d_in(u_ca_in_1272), .d_out(u_ca_out_1272));
compressor_243_72 u_ca_243_72_1273(.d_in(u_ca_in_1273), .d_out(u_ca_out_1273));
compressor_243_72 u_ca_243_72_1274(.d_in(u_ca_in_1274), .d_out(u_ca_out_1274));
compressor_243_72 u_ca_243_72_1275(.d_in(u_ca_in_1275), .d_out(u_ca_out_1275));
compressor_243_72 u_ca_243_72_1276(.d_in(u_ca_in_1276), .d_out(u_ca_out_1276));
compressor_243_72 u_ca_243_72_1277(.d_in(u_ca_in_1277), .d_out(u_ca_out_1277));
compressor_243_72 u_ca_243_72_1278(.d_in(u_ca_in_1278), .d_out(u_ca_out_1278));
compressor_243_72 u_ca_243_72_1279(.d_in(u_ca_in_1279), .d_out(u_ca_out_1279));

//---------------------------------------------------------



//--output-------------------------------------------------

assign col_out_0 = {{63{1'b0}}, u_ca_out_0[8:0]};
assign col_out_1 = {{36{1'b0}}, u_ca_out_1[8:0], u_ca_out_0[35:9]};
assign col_out_2 = {{9{1'b0}}, u_ca_out_2[8:0], u_ca_out_1[35:9], u_ca_out_0[62:36]};
assign col_out_3 = {u_ca_out_3[8:0],u_ca_out_2[35:9], u_ca_out_1[62:36], u_ca_out_0[71:63]};
assign col_out_4 = {u_ca_out_4[8:0],u_ca_out_3[35:9], u_ca_out_2[62:36], u_ca_out_1[71:63]};
assign col_out_5 = {u_ca_out_5[8:0],u_ca_out_4[35:9], u_ca_out_3[62:36], u_ca_out_2[71:63]};
assign col_out_6 = {u_ca_out_6[8:0],u_ca_out_5[35:9], u_ca_out_4[62:36], u_ca_out_3[71:63]};
assign col_out_7 = {u_ca_out_7[8:0],u_ca_out_6[35:9], u_ca_out_5[62:36], u_ca_out_4[71:63]};
assign col_out_8 = {u_ca_out_8[8:0],u_ca_out_7[35:9], u_ca_out_6[62:36], u_ca_out_5[71:63]};
assign col_out_9 = {u_ca_out_9[8:0],u_ca_out_8[35:9], u_ca_out_7[62:36], u_ca_out_6[71:63]};
assign col_out_10 = {u_ca_out_10[8:0],u_ca_out_9[35:9], u_ca_out_8[62:36], u_ca_out_7[71:63]};
assign col_out_11 = {u_ca_out_11[8:0],u_ca_out_10[35:9], u_ca_out_9[62:36], u_ca_out_8[71:63]};
assign col_out_12 = {u_ca_out_12[8:0],u_ca_out_11[35:9], u_ca_out_10[62:36], u_ca_out_9[71:63]};
assign col_out_13 = {u_ca_out_13[8:0],u_ca_out_12[35:9], u_ca_out_11[62:36], u_ca_out_10[71:63]};
assign col_out_14 = {u_ca_out_14[8:0],u_ca_out_13[35:9], u_ca_out_12[62:36], u_ca_out_11[71:63]};
assign col_out_15 = {u_ca_out_15[8:0],u_ca_out_14[35:9], u_ca_out_13[62:36], u_ca_out_12[71:63]};
assign col_out_16 = {u_ca_out_16[8:0],u_ca_out_15[35:9], u_ca_out_14[62:36], u_ca_out_13[71:63]};
assign col_out_17 = {u_ca_out_17[8:0],u_ca_out_16[35:9], u_ca_out_15[62:36], u_ca_out_14[71:63]};
assign col_out_18 = {u_ca_out_18[8:0],u_ca_out_17[35:9], u_ca_out_16[62:36], u_ca_out_15[71:63]};
assign col_out_19 = {u_ca_out_19[8:0],u_ca_out_18[35:9], u_ca_out_17[62:36], u_ca_out_16[71:63]};
assign col_out_20 = {u_ca_out_20[8:0],u_ca_out_19[35:9], u_ca_out_18[62:36], u_ca_out_17[71:63]};
assign col_out_21 = {u_ca_out_21[8:0],u_ca_out_20[35:9], u_ca_out_19[62:36], u_ca_out_18[71:63]};
assign col_out_22 = {u_ca_out_22[8:0],u_ca_out_21[35:9], u_ca_out_20[62:36], u_ca_out_19[71:63]};
assign col_out_23 = {u_ca_out_23[8:0],u_ca_out_22[35:9], u_ca_out_21[62:36], u_ca_out_20[71:63]};
assign col_out_24 = {u_ca_out_24[8:0],u_ca_out_23[35:9], u_ca_out_22[62:36], u_ca_out_21[71:63]};
assign col_out_25 = {u_ca_out_25[8:0],u_ca_out_24[35:9], u_ca_out_23[62:36], u_ca_out_22[71:63]};
assign col_out_26 = {u_ca_out_26[8:0],u_ca_out_25[35:9], u_ca_out_24[62:36], u_ca_out_23[71:63]};
assign col_out_27 = {u_ca_out_27[8:0],u_ca_out_26[35:9], u_ca_out_25[62:36], u_ca_out_24[71:63]};
assign col_out_28 = {u_ca_out_28[8:0],u_ca_out_27[35:9], u_ca_out_26[62:36], u_ca_out_25[71:63]};
assign col_out_29 = {u_ca_out_29[8:0],u_ca_out_28[35:9], u_ca_out_27[62:36], u_ca_out_26[71:63]};
assign col_out_30 = {u_ca_out_30[8:0],u_ca_out_29[35:9], u_ca_out_28[62:36], u_ca_out_27[71:63]};
assign col_out_31 = {u_ca_out_31[8:0],u_ca_out_30[35:9], u_ca_out_29[62:36], u_ca_out_28[71:63]};
assign col_out_32 = {u_ca_out_32[8:0],u_ca_out_31[35:9], u_ca_out_30[62:36], u_ca_out_29[71:63]};
assign col_out_33 = {u_ca_out_33[8:0],u_ca_out_32[35:9], u_ca_out_31[62:36], u_ca_out_30[71:63]};
assign col_out_34 = {u_ca_out_34[8:0],u_ca_out_33[35:9], u_ca_out_32[62:36], u_ca_out_31[71:63]};
assign col_out_35 = {u_ca_out_35[8:0],u_ca_out_34[35:9], u_ca_out_33[62:36], u_ca_out_32[71:63]};
assign col_out_36 = {u_ca_out_36[8:0],u_ca_out_35[35:9], u_ca_out_34[62:36], u_ca_out_33[71:63]};
assign col_out_37 = {u_ca_out_37[8:0],u_ca_out_36[35:9], u_ca_out_35[62:36], u_ca_out_34[71:63]};
assign col_out_38 = {u_ca_out_38[8:0],u_ca_out_37[35:9], u_ca_out_36[62:36], u_ca_out_35[71:63]};
assign col_out_39 = {u_ca_out_39[8:0],u_ca_out_38[35:9], u_ca_out_37[62:36], u_ca_out_36[71:63]};
assign col_out_40 = {u_ca_out_40[8:0],u_ca_out_39[35:9], u_ca_out_38[62:36], u_ca_out_37[71:63]};
assign col_out_41 = {u_ca_out_41[8:0],u_ca_out_40[35:9], u_ca_out_39[62:36], u_ca_out_38[71:63]};
assign col_out_42 = {u_ca_out_42[8:0],u_ca_out_41[35:9], u_ca_out_40[62:36], u_ca_out_39[71:63]};
assign col_out_43 = {u_ca_out_43[8:0],u_ca_out_42[35:9], u_ca_out_41[62:36], u_ca_out_40[71:63]};
assign col_out_44 = {u_ca_out_44[8:0],u_ca_out_43[35:9], u_ca_out_42[62:36], u_ca_out_41[71:63]};
assign col_out_45 = {u_ca_out_45[8:0],u_ca_out_44[35:9], u_ca_out_43[62:36], u_ca_out_42[71:63]};
assign col_out_46 = {u_ca_out_46[8:0],u_ca_out_45[35:9], u_ca_out_44[62:36], u_ca_out_43[71:63]};
assign col_out_47 = {u_ca_out_47[8:0],u_ca_out_46[35:9], u_ca_out_45[62:36], u_ca_out_44[71:63]};
assign col_out_48 = {u_ca_out_48[8:0],u_ca_out_47[35:9], u_ca_out_46[62:36], u_ca_out_45[71:63]};
assign col_out_49 = {u_ca_out_49[8:0],u_ca_out_48[35:9], u_ca_out_47[62:36], u_ca_out_46[71:63]};
assign col_out_50 = {u_ca_out_50[8:0],u_ca_out_49[35:9], u_ca_out_48[62:36], u_ca_out_47[71:63]};
assign col_out_51 = {u_ca_out_51[8:0],u_ca_out_50[35:9], u_ca_out_49[62:36], u_ca_out_48[71:63]};
assign col_out_52 = {u_ca_out_52[8:0],u_ca_out_51[35:9], u_ca_out_50[62:36], u_ca_out_49[71:63]};
assign col_out_53 = {u_ca_out_53[8:0],u_ca_out_52[35:9], u_ca_out_51[62:36], u_ca_out_50[71:63]};
assign col_out_54 = {u_ca_out_54[8:0],u_ca_out_53[35:9], u_ca_out_52[62:36], u_ca_out_51[71:63]};
assign col_out_55 = {u_ca_out_55[8:0],u_ca_out_54[35:9], u_ca_out_53[62:36], u_ca_out_52[71:63]};
assign col_out_56 = {u_ca_out_56[8:0],u_ca_out_55[35:9], u_ca_out_54[62:36], u_ca_out_53[71:63]};
assign col_out_57 = {u_ca_out_57[8:0],u_ca_out_56[35:9], u_ca_out_55[62:36], u_ca_out_54[71:63]};
assign col_out_58 = {u_ca_out_58[8:0],u_ca_out_57[35:9], u_ca_out_56[62:36], u_ca_out_55[71:63]};
assign col_out_59 = {u_ca_out_59[8:0],u_ca_out_58[35:9], u_ca_out_57[62:36], u_ca_out_56[71:63]};
assign col_out_60 = {u_ca_out_60[8:0],u_ca_out_59[35:9], u_ca_out_58[62:36], u_ca_out_57[71:63]};
assign col_out_61 = {u_ca_out_61[8:0],u_ca_out_60[35:9], u_ca_out_59[62:36], u_ca_out_58[71:63]};
assign col_out_62 = {u_ca_out_62[8:0],u_ca_out_61[35:9], u_ca_out_60[62:36], u_ca_out_59[71:63]};
assign col_out_63 = {u_ca_out_63[8:0],u_ca_out_62[35:9], u_ca_out_61[62:36], u_ca_out_60[71:63]};
assign col_out_64 = {u_ca_out_64[8:0],u_ca_out_63[35:9], u_ca_out_62[62:36], u_ca_out_61[71:63]};
assign col_out_65 = {u_ca_out_65[8:0],u_ca_out_64[35:9], u_ca_out_63[62:36], u_ca_out_62[71:63]};
assign col_out_66 = {u_ca_out_66[8:0],u_ca_out_65[35:9], u_ca_out_64[62:36], u_ca_out_63[71:63]};
assign col_out_67 = {u_ca_out_67[8:0],u_ca_out_66[35:9], u_ca_out_65[62:36], u_ca_out_64[71:63]};
assign col_out_68 = {u_ca_out_68[8:0],u_ca_out_67[35:9], u_ca_out_66[62:36], u_ca_out_65[71:63]};
assign col_out_69 = {u_ca_out_69[8:0],u_ca_out_68[35:9], u_ca_out_67[62:36], u_ca_out_66[71:63]};
assign col_out_70 = {u_ca_out_70[8:0],u_ca_out_69[35:9], u_ca_out_68[62:36], u_ca_out_67[71:63]};
assign col_out_71 = {u_ca_out_71[8:0],u_ca_out_70[35:9], u_ca_out_69[62:36], u_ca_out_68[71:63]};
assign col_out_72 = {u_ca_out_72[8:0],u_ca_out_71[35:9], u_ca_out_70[62:36], u_ca_out_69[71:63]};
assign col_out_73 = {u_ca_out_73[8:0],u_ca_out_72[35:9], u_ca_out_71[62:36], u_ca_out_70[71:63]};
assign col_out_74 = {u_ca_out_74[8:0],u_ca_out_73[35:9], u_ca_out_72[62:36], u_ca_out_71[71:63]};
assign col_out_75 = {u_ca_out_75[8:0],u_ca_out_74[35:9], u_ca_out_73[62:36], u_ca_out_72[71:63]};
assign col_out_76 = {u_ca_out_76[8:0],u_ca_out_75[35:9], u_ca_out_74[62:36], u_ca_out_73[71:63]};
assign col_out_77 = {u_ca_out_77[8:0],u_ca_out_76[35:9], u_ca_out_75[62:36], u_ca_out_74[71:63]};
assign col_out_78 = {u_ca_out_78[8:0],u_ca_out_77[35:9], u_ca_out_76[62:36], u_ca_out_75[71:63]};
assign col_out_79 = {u_ca_out_79[8:0],u_ca_out_78[35:9], u_ca_out_77[62:36], u_ca_out_76[71:63]};
assign col_out_80 = {u_ca_out_80[8:0],u_ca_out_79[35:9], u_ca_out_78[62:36], u_ca_out_77[71:63]};
assign col_out_81 = {u_ca_out_81[8:0],u_ca_out_80[35:9], u_ca_out_79[62:36], u_ca_out_78[71:63]};
assign col_out_82 = {u_ca_out_82[8:0],u_ca_out_81[35:9], u_ca_out_80[62:36], u_ca_out_79[71:63]};
assign col_out_83 = {u_ca_out_83[8:0],u_ca_out_82[35:9], u_ca_out_81[62:36], u_ca_out_80[71:63]};
assign col_out_84 = {u_ca_out_84[8:0],u_ca_out_83[35:9], u_ca_out_82[62:36], u_ca_out_81[71:63]};
assign col_out_85 = {u_ca_out_85[8:0],u_ca_out_84[35:9], u_ca_out_83[62:36], u_ca_out_82[71:63]};
assign col_out_86 = {u_ca_out_86[8:0],u_ca_out_85[35:9], u_ca_out_84[62:36], u_ca_out_83[71:63]};
assign col_out_87 = {u_ca_out_87[8:0],u_ca_out_86[35:9], u_ca_out_85[62:36], u_ca_out_84[71:63]};
assign col_out_88 = {u_ca_out_88[8:0],u_ca_out_87[35:9], u_ca_out_86[62:36], u_ca_out_85[71:63]};
assign col_out_89 = {u_ca_out_89[8:0],u_ca_out_88[35:9], u_ca_out_87[62:36], u_ca_out_86[71:63]};
assign col_out_90 = {u_ca_out_90[8:0],u_ca_out_89[35:9], u_ca_out_88[62:36], u_ca_out_87[71:63]};
assign col_out_91 = {u_ca_out_91[8:0],u_ca_out_90[35:9], u_ca_out_89[62:36], u_ca_out_88[71:63]};
assign col_out_92 = {u_ca_out_92[8:0],u_ca_out_91[35:9], u_ca_out_90[62:36], u_ca_out_89[71:63]};
assign col_out_93 = {u_ca_out_93[8:0],u_ca_out_92[35:9], u_ca_out_91[62:36], u_ca_out_90[71:63]};
assign col_out_94 = {u_ca_out_94[8:0],u_ca_out_93[35:9], u_ca_out_92[62:36], u_ca_out_91[71:63]};
assign col_out_95 = {u_ca_out_95[8:0],u_ca_out_94[35:9], u_ca_out_93[62:36], u_ca_out_92[71:63]};
assign col_out_96 = {u_ca_out_96[8:0],u_ca_out_95[35:9], u_ca_out_94[62:36], u_ca_out_93[71:63]};
assign col_out_97 = {u_ca_out_97[8:0],u_ca_out_96[35:9], u_ca_out_95[62:36], u_ca_out_94[71:63]};
assign col_out_98 = {u_ca_out_98[8:0],u_ca_out_97[35:9], u_ca_out_96[62:36], u_ca_out_95[71:63]};
assign col_out_99 = {u_ca_out_99[8:0],u_ca_out_98[35:9], u_ca_out_97[62:36], u_ca_out_96[71:63]};
assign col_out_100 = {u_ca_out_100[8:0],u_ca_out_99[35:9], u_ca_out_98[62:36], u_ca_out_97[71:63]};
assign col_out_101 = {u_ca_out_101[8:0],u_ca_out_100[35:9], u_ca_out_99[62:36], u_ca_out_98[71:63]};
assign col_out_102 = {u_ca_out_102[8:0],u_ca_out_101[35:9], u_ca_out_100[62:36], u_ca_out_99[71:63]};
assign col_out_103 = {u_ca_out_103[8:0],u_ca_out_102[35:9], u_ca_out_101[62:36], u_ca_out_100[71:63]};
assign col_out_104 = {u_ca_out_104[8:0],u_ca_out_103[35:9], u_ca_out_102[62:36], u_ca_out_101[71:63]};
assign col_out_105 = {u_ca_out_105[8:0],u_ca_out_104[35:9], u_ca_out_103[62:36], u_ca_out_102[71:63]};
assign col_out_106 = {u_ca_out_106[8:0],u_ca_out_105[35:9], u_ca_out_104[62:36], u_ca_out_103[71:63]};
assign col_out_107 = {u_ca_out_107[8:0],u_ca_out_106[35:9], u_ca_out_105[62:36], u_ca_out_104[71:63]};
assign col_out_108 = {u_ca_out_108[8:0],u_ca_out_107[35:9], u_ca_out_106[62:36], u_ca_out_105[71:63]};
assign col_out_109 = {u_ca_out_109[8:0],u_ca_out_108[35:9], u_ca_out_107[62:36], u_ca_out_106[71:63]};
assign col_out_110 = {u_ca_out_110[8:0],u_ca_out_109[35:9], u_ca_out_108[62:36], u_ca_out_107[71:63]};
assign col_out_111 = {u_ca_out_111[8:0],u_ca_out_110[35:9], u_ca_out_109[62:36], u_ca_out_108[71:63]};
assign col_out_112 = {u_ca_out_112[8:0],u_ca_out_111[35:9], u_ca_out_110[62:36], u_ca_out_109[71:63]};
assign col_out_113 = {u_ca_out_113[8:0],u_ca_out_112[35:9], u_ca_out_111[62:36], u_ca_out_110[71:63]};
assign col_out_114 = {u_ca_out_114[8:0],u_ca_out_113[35:9], u_ca_out_112[62:36], u_ca_out_111[71:63]};
assign col_out_115 = {u_ca_out_115[8:0],u_ca_out_114[35:9], u_ca_out_113[62:36], u_ca_out_112[71:63]};
assign col_out_116 = {u_ca_out_116[8:0],u_ca_out_115[35:9], u_ca_out_114[62:36], u_ca_out_113[71:63]};
assign col_out_117 = {u_ca_out_117[8:0],u_ca_out_116[35:9], u_ca_out_115[62:36], u_ca_out_114[71:63]};
assign col_out_118 = {u_ca_out_118[8:0],u_ca_out_117[35:9], u_ca_out_116[62:36], u_ca_out_115[71:63]};
assign col_out_119 = {u_ca_out_119[8:0],u_ca_out_118[35:9], u_ca_out_117[62:36], u_ca_out_116[71:63]};
assign col_out_120 = {u_ca_out_120[8:0],u_ca_out_119[35:9], u_ca_out_118[62:36], u_ca_out_117[71:63]};
assign col_out_121 = {u_ca_out_121[8:0],u_ca_out_120[35:9], u_ca_out_119[62:36], u_ca_out_118[71:63]};
assign col_out_122 = {u_ca_out_122[8:0],u_ca_out_121[35:9], u_ca_out_120[62:36], u_ca_out_119[71:63]};
assign col_out_123 = {u_ca_out_123[8:0],u_ca_out_122[35:9], u_ca_out_121[62:36], u_ca_out_120[71:63]};
assign col_out_124 = {u_ca_out_124[8:0],u_ca_out_123[35:9], u_ca_out_122[62:36], u_ca_out_121[71:63]};
assign col_out_125 = {u_ca_out_125[8:0],u_ca_out_124[35:9], u_ca_out_123[62:36], u_ca_out_122[71:63]};
assign col_out_126 = {u_ca_out_126[8:0],u_ca_out_125[35:9], u_ca_out_124[62:36], u_ca_out_123[71:63]};
assign col_out_127 = {u_ca_out_127[8:0],u_ca_out_126[35:9], u_ca_out_125[62:36], u_ca_out_124[71:63]};
assign col_out_128 = {u_ca_out_128[8:0],u_ca_out_127[35:9], u_ca_out_126[62:36], u_ca_out_125[71:63]};
assign col_out_129 = {u_ca_out_129[8:0],u_ca_out_128[35:9], u_ca_out_127[62:36], u_ca_out_126[71:63]};
assign col_out_130 = {u_ca_out_130[8:0],u_ca_out_129[35:9], u_ca_out_128[62:36], u_ca_out_127[71:63]};
assign col_out_131 = {u_ca_out_131[8:0],u_ca_out_130[35:9], u_ca_out_129[62:36], u_ca_out_128[71:63]};
assign col_out_132 = {u_ca_out_132[8:0],u_ca_out_131[35:9], u_ca_out_130[62:36], u_ca_out_129[71:63]};
assign col_out_133 = {u_ca_out_133[8:0],u_ca_out_132[35:9], u_ca_out_131[62:36], u_ca_out_130[71:63]};
assign col_out_134 = {u_ca_out_134[8:0],u_ca_out_133[35:9], u_ca_out_132[62:36], u_ca_out_131[71:63]};
assign col_out_135 = {u_ca_out_135[8:0],u_ca_out_134[35:9], u_ca_out_133[62:36], u_ca_out_132[71:63]};
assign col_out_136 = {u_ca_out_136[8:0],u_ca_out_135[35:9], u_ca_out_134[62:36], u_ca_out_133[71:63]};
assign col_out_137 = {u_ca_out_137[8:0],u_ca_out_136[35:9], u_ca_out_135[62:36], u_ca_out_134[71:63]};
assign col_out_138 = {u_ca_out_138[8:0],u_ca_out_137[35:9], u_ca_out_136[62:36], u_ca_out_135[71:63]};
assign col_out_139 = {u_ca_out_139[8:0],u_ca_out_138[35:9], u_ca_out_137[62:36], u_ca_out_136[71:63]};
assign col_out_140 = {u_ca_out_140[8:0],u_ca_out_139[35:9], u_ca_out_138[62:36], u_ca_out_137[71:63]};
assign col_out_141 = {u_ca_out_141[8:0],u_ca_out_140[35:9], u_ca_out_139[62:36], u_ca_out_138[71:63]};
assign col_out_142 = {u_ca_out_142[8:0],u_ca_out_141[35:9], u_ca_out_140[62:36], u_ca_out_139[71:63]};
assign col_out_143 = {u_ca_out_143[8:0],u_ca_out_142[35:9], u_ca_out_141[62:36], u_ca_out_140[71:63]};
assign col_out_144 = {u_ca_out_144[8:0],u_ca_out_143[35:9], u_ca_out_142[62:36], u_ca_out_141[71:63]};
assign col_out_145 = {u_ca_out_145[8:0],u_ca_out_144[35:9], u_ca_out_143[62:36], u_ca_out_142[71:63]};
assign col_out_146 = {u_ca_out_146[8:0],u_ca_out_145[35:9], u_ca_out_144[62:36], u_ca_out_143[71:63]};
assign col_out_147 = {u_ca_out_147[8:0],u_ca_out_146[35:9], u_ca_out_145[62:36], u_ca_out_144[71:63]};
assign col_out_148 = {u_ca_out_148[8:0],u_ca_out_147[35:9], u_ca_out_146[62:36], u_ca_out_145[71:63]};
assign col_out_149 = {u_ca_out_149[8:0],u_ca_out_148[35:9], u_ca_out_147[62:36], u_ca_out_146[71:63]};
assign col_out_150 = {u_ca_out_150[8:0],u_ca_out_149[35:9], u_ca_out_148[62:36], u_ca_out_147[71:63]};
assign col_out_151 = {u_ca_out_151[8:0],u_ca_out_150[35:9], u_ca_out_149[62:36], u_ca_out_148[71:63]};
assign col_out_152 = {u_ca_out_152[8:0],u_ca_out_151[35:9], u_ca_out_150[62:36], u_ca_out_149[71:63]};
assign col_out_153 = {u_ca_out_153[8:0],u_ca_out_152[35:9], u_ca_out_151[62:36], u_ca_out_150[71:63]};
assign col_out_154 = {u_ca_out_154[8:0],u_ca_out_153[35:9], u_ca_out_152[62:36], u_ca_out_151[71:63]};
assign col_out_155 = {u_ca_out_155[8:0],u_ca_out_154[35:9], u_ca_out_153[62:36], u_ca_out_152[71:63]};
assign col_out_156 = {u_ca_out_156[8:0],u_ca_out_155[35:9], u_ca_out_154[62:36], u_ca_out_153[71:63]};
assign col_out_157 = {u_ca_out_157[8:0],u_ca_out_156[35:9], u_ca_out_155[62:36], u_ca_out_154[71:63]};
assign col_out_158 = {u_ca_out_158[8:0],u_ca_out_157[35:9], u_ca_out_156[62:36], u_ca_out_155[71:63]};
assign col_out_159 = {u_ca_out_159[8:0],u_ca_out_158[35:9], u_ca_out_157[62:36], u_ca_out_156[71:63]};
assign col_out_160 = {u_ca_out_160[8:0],u_ca_out_159[35:9], u_ca_out_158[62:36], u_ca_out_157[71:63]};
assign col_out_161 = {u_ca_out_161[8:0],u_ca_out_160[35:9], u_ca_out_159[62:36], u_ca_out_158[71:63]};
assign col_out_162 = {u_ca_out_162[8:0],u_ca_out_161[35:9], u_ca_out_160[62:36], u_ca_out_159[71:63]};
assign col_out_163 = {u_ca_out_163[8:0],u_ca_out_162[35:9], u_ca_out_161[62:36], u_ca_out_160[71:63]};
assign col_out_164 = {u_ca_out_164[8:0],u_ca_out_163[35:9], u_ca_out_162[62:36], u_ca_out_161[71:63]};
assign col_out_165 = {u_ca_out_165[8:0],u_ca_out_164[35:9], u_ca_out_163[62:36], u_ca_out_162[71:63]};
assign col_out_166 = {u_ca_out_166[8:0],u_ca_out_165[35:9], u_ca_out_164[62:36], u_ca_out_163[71:63]};
assign col_out_167 = {u_ca_out_167[8:0],u_ca_out_166[35:9], u_ca_out_165[62:36], u_ca_out_164[71:63]};
assign col_out_168 = {u_ca_out_168[8:0],u_ca_out_167[35:9], u_ca_out_166[62:36], u_ca_out_165[71:63]};
assign col_out_169 = {u_ca_out_169[8:0],u_ca_out_168[35:9], u_ca_out_167[62:36], u_ca_out_166[71:63]};
assign col_out_170 = {u_ca_out_170[8:0],u_ca_out_169[35:9], u_ca_out_168[62:36], u_ca_out_167[71:63]};
assign col_out_171 = {u_ca_out_171[8:0],u_ca_out_170[35:9], u_ca_out_169[62:36], u_ca_out_168[71:63]};
assign col_out_172 = {u_ca_out_172[8:0],u_ca_out_171[35:9], u_ca_out_170[62:36], u_ca_out_169[71:63]};
assign col_out_173 = {u_ca_out_173[8:0],u_ca_out_172[35:9], u_ca_out_171[62:36], u_ca_out_170[71:63]};
assign col_out_174 = {u_ca_out_174[8:0],u_ca_out_173[35:9], u_ca_out_172[62:36], u_ca_out_171[71:63]};
assign col_out_175 = {u_ca_out_175[8:0],u_ca_out_174[35:9], u_ca_out_173[62:36], u_ca_out_172[71:63]};
assign col_out_176 = {u_ca_out_176[8:0],u_ca_out_175[35:9], u_ca_out_174[62:36], u_ca_out_173[71:63]};
assign col_out_177 = {u_ca_out_177[8:0],u_ca_out_176[35:9], u_ca_out_175[62:36], u_ca_out_174[71:63]};
assign col_out_178 = {u_ca_out_178[8:0],u_ca_out_177[35:9], u_ca_out_176[62:36], u_ca_out_175[71:63]};
assign col_out_179 = {u_ca_out_179[8:0],u_ca_out_178[35:9], u_ca_out_177[62:36], u_ca_out_176[71:63]};
assign col_out_180 = {u_ca_out_180[8:0],u_ca_out_179[35:9], u_ca_out_178[62:36], u_ca_out_177[71:63]};
assign col_out_181 = {u_ca_out_181[8:0],u_ca_out_180[35:9], u_ca_out_179[62:36], u_ca_out_178[71:63]};
assign col_out_182 = {u_ca_out_182[8:0],u_ca_out_181[35:9], u_ca_out_180[62:36], u_ca_out_179[71:63]};
assign col_out_183 = {u_ca_out_183[8:0],u_ca_out_182[35:9], u_ca_out_181[62:36], u_ca_out_180[71:63]};
assign col_out_184 = {u_ca_out_184[8:0],u_ca_out_183[35:9], u_ca_out_182[62:36], u_ca_out_181[71:63]};
assign col_out_185 = {u_ca_out_185[8:0],u_ca_out_184[35:9], u_ca_out_183[62:36], u_ca_out_182[71:63]};
assign col_out_186 = {u_ca_out_186[8:0],u_ca_out_185[35:9], u_ca_out_184[62:36], u_ca_out_183[71:63]};
assign col_out_187 = {u_ca_out_187[8:0],u_ca_out_186[35:9], u_ca_out_185[62:36], u_ca_out_184[71:63]};
assign col_out_188 = {u_ca_out_188[8:0],u_ca_out_187[35:9], u_ca_out_186[62:36], u_ca_out_185[71:63]};
assign col_out_189 = {u_ca_out_189[8:0],u_ca_out_188[35:9], u_ca_out_187[62:36], u_ca_out_186[71:63]};
assign col_out_190 = {u_ca_out_190[8:0],u_ca_out_189[35:9], u_ca_out_188[62:36], u_ca_out_187[71:63]};
assign col_out_191 = {u_ca_out_191[8:0],u_ca_out_190[35:9], u_ca_out_189[62:36], u_ca_out_188[71:63]};
assign col_out_192 = {u_ca_out_192[8:0],u_ca_out_191[35:9], u_ca_out_190[62:36], u_ca_out_189[71:63]};
assign col_out_193 = {u_ca_out_193[8:0],u_ca_out_192[35:9], u_ca_out_191[62:36], u_ca_out_190[71:63]};
assign col_out_194 = {u_ca_out_194[8:0],u_ca_out_193[35:9], u_ca_out_192[62:36], u_ca_out_191[71:63]};
assign col_out_195 = {u_ca_out_195[8:0],u_ca_out_194[35:9], u_ca_out_193[62:36], u_ca_out_192[71:63]};
assign col_out_196 = {u_ca_out_196[8:0],u_ca_out_195[35:9], u_ca_out_194[62:36], u_ca_out_193[71:63]};
assign col_out_197 = {u_ca_out_197[8:0],u_ca_out_196[35:9], u_ca_out_195[62:36], u_ca_out_194[71:63]};
assign col_out_198 = {u_ca_out_198[8:0],u_ca_out_197[35:9], u_ca_out_196[62:36], u_ca_out_195[71:63]};
assign col_out_199 = {u_ca_out_199[8:0],u_ca_out_198[35:9], u_ca_out_197[62:36], u_ca_out_196[71:63]};
assign col_out_200 = {u_ca_out_200[8:0],u_ca_out_199[35:9], u_ca_out_198[62:36], u_ca_out_197[71:63]};
assign col_out_201 = {u_ca_out_201[8:0],u_ca_out_200[35:9], u_ca_out_199[62:36], u_ca_out_198[71:63]};
assign col_out_202 = {u_ca_out_202[8:0],u_ca_out_201[35:9], u_ca_out_200[62:36], u_ca_out_199[71:63]};
assign col_out_203 = {u_ca_out_203[8:0],u_ca_out_202[35:9], u_ca_out_201[62:36], u_ca_out_200[71:63]};
assign col_out_204 = {u_ca_out_204[8:0],u_ca_out_203[35:9], u_ca_out_202[62:36], u_ca_out_201[71:63]};
assign col_out_205 = {u_ca_out_205[8:0],u_ca_out_204[35:9], u_ca_out_203[62:36], u_ca_out_202[71:63]};
assign col_out_206 = {u_ca_out_206[8:0],u_ca_out_205[35:9], u_ca_out_204[62:36], u_ca_out_203[71:63]};
assign col_out_207 = {u_ca_out_207[8:0],u_ca_out_206[35:9], u_ca_out_205[62:36], u_ca_out_204[71:63]};
assign col_out_208 = {u_ca_out_208[8:0],u_ca_out_207[35:9], u_ca_out_206[62:36], u_ca_out_205[71:63]};
assign col_out_209 = {u_ca_out_209[8:0],u_ca_out_208[35:9], u_ca_out_207[62:36], u_ca_out_206[71:63]};
assign col_out_210 = {u_ca_out_210[8:0],u_ca_out_209[35:9], u_ca_out_208[62:36], u_ca_out_207[71:63]};
assign col_out_211 = {u_ca_out_211[8:0],u_ca_out_210[35:9], u_ca_out_209[62:36], u_ca_out_208[71:63]};
assign col_out_212 = {u_ca_out_212[8:0],u_ca_out_211[35:9], u_ca_out_210[62:36], u_ca_out_209[71:63]};
assign col_out_213 = {u_ca_out_213[8:0],u_ca_out_212[35:9], u_ca_out_211[62:36], u_ca_out_210[71:63]};
assign col_out_214 = {u_ca_out_214[8:0],u_ca_out_213[35:9], u_ca_out_212[62:36], u_ca_out_211[71:63]};
assign col_out_215 = {u_ca_out_215[8:0],u_ca_out_214[35:9], u_ca_out_213[62:36], u_ca_out_212[71:63]};
assign col_out_216 = {u_ca_out_216[8:0],u_ca_out_215[35:9], u_ca_out_214[62:36], u_ca_out_213[71:63]};
assign col_out_217 = {u_ca_out_217[8:0],u_ca_out_216[35:9], u_ca_out_215[62:36], u_ca_out_214[71:63]};
assign col_out_218 = {u_ca_out_218[8:0],u_ca_out_217[35:9], u_ca_out_216[62:36], u_ca_out_215[71:63]};
assign col_out_219 = {u_ca_out_219[8:0],u_ca_out_218[35:9], u_ca_out_217[62:36], u_ca_out_216[71:63]};
assign col_out_220 = {u_ca_out_220[8:0],u_ca_out_219[35:9], u_ca_out_218[62:36], u_ca_out_217[71:63]};
assign col_out_221 = {u_ca_out_221[8:0],u_ca_out_220[35:9], u_ca_out_219[62:36], u_ca_out_218[71:63]};
assign col_out_222 = {u_ca_out_222[8:0],u_ca_out_221[35:9], u_ca_out_220[62:36], u_ca_out_219[71:63]};
assign col_out_223 = {u_ca_out_223[8:0],u_ca_out_222[35:9], u_ca_out_221[62:36], u_ca_out_220[71:63]};
assign col_out_224 = {u_ca_out_224[8:0],u_ca_out_223[35:9], u_ca_out_222[62:36], u_ca_out_221[71:63]};
assign col_out_225 = {u_ca_out_225[8:0],u_ca_out_224[35:9], u_ca_out_223[62:36], u_ca_out_222[71:63]};
assign col_out_226 = {u_ca_out_226[8:0],u_ca_out_225[35:9], u_ca_out_224[62:36], u_ca_out_223[71:63]};
assign col_out_227 = {u_ca_out_227[8:0],u_ca_out_226[35:9], u_ca_out_225[62:36], u_ca_out_224[71:63]};
assign col_out_228 = {u_ca_out_228[8:0],u_ca_out_227[35:9], u_ca_out_226[62:36], u_ca_out_225[71:63]};
assign col_out_229 = {u_ca_out_229[8:0],u_ca_out_228[35:9], u_ca_out_227[62:36], u_ca_out_226[71:63]};
assign col_out_230 = {u_ca_out_230[8:0],u_ca_out_229[35:9], u_ca_out_228[62:36], u_ca_out_227[71:63]};
assign col_out_231 = {u_ca_out_231[8:0],u_ca_out_230[35:9], u_ca_out_229[62:36], u_ca_out_228[71:63]};
assign col_out_232 = {u_ca_out_232[8:0],u_ca_out_231[35:9], u_ca_out_230[62:36], u_ca_out_229[71:63]};
assign col_out_233 = {u_ca_out_233[8:0],u_ca_out_232[35:9], u_ca_out_231[62:36], u_ca_out_230[71:63]};
assign col_out_234 = {u_ca_out_234[8:0],u_ca_out_233[35:9], u_ca_out_232[62:36], u_ca_out_231[71:63]};
assign col_out_235 = {u_ca_out_235[8:0],u_ca_out_234[35:9], u_ca_out_233[62:36], u_ca_out_232[71:63]};
assign col_out_236 = {u_ca_out_236[8:0],u_ca_out_235[35:9], u_ca_out_234[62:36], u_ca_out_233[71:63]};
assign col_out_237 = {u_ca_out_237[8:0],u_ca_out_236[35:9], u_ca_out_235[62:36], u_ca_out_234[71:63]};
assign col_out_238 = {u_ca_out_238[8:0],u_ca_out_237[35:9], u_ca_out_236[62:36], u_ca_out_235[71:63]};
assign col_out_239 = {u_ca_out_239[8:0],u_ca_out_238[35:9], u_ca_out_237[62:36], u_ca_out_236[71:63]};
assign col_out_240 = {u_ca_out_240[8:0],u_ca_out_239[35:9], u_ca_out_238[62:36], u_ca_out_237[71:63]};
assign col_out_241 = {u_ca_out_241[8:0],u_ca_out_240[35:9], u_ca_out_239[62:36], u_ca_out_238[71:63]};
assign col_out_242 = {u_ca_out_242[8:0],u_ca_out_241[35:9], u_ca_out_240[62:36], u_ca_out_239[71:63]};
assign col_out_243 = {u_ca_out_243[8:0],u_ca_out_242[35:9], u_ca_out_241[62:36], u_ca_out_240[71:63]};
assign col_out_244 = {u_ca_out_244[8:0],u_ca_out_243[35:9], u_ca_out_242[62:36], u_ca_out_241[71:63]};
assign col_out_245 = {u_ca_out_245[8:0],u_ca_out_244[35:9], u_ca_out_243[62:36], u_ca_out_242[71:63]};
assign col_out_246 = {u_ca_out_246[8:0],u_ca_out_245[35:9], u_ca_out_244[62:36], u_ca_out_243[71:63]};
assign col_out_247 = {u_ca_out_247[8:0],u_ca_out_246[35:9], u_ca_out_245[62:36], u_ca_out_244[71:63]};
assign col_out_248 = {u_ca_out_248[8:0],u_ca_out_247[35:9], u_ca_out_246[62:36], u_ca_out_245[71:63]};
assign col_out_249 = {u_ca_out_249[8:0],u_ca_out_248[35:9], u_ca_out_247[62:36], u_ca_out_246[71:63]};
assign col_out_250 = {u_ca_out_250[8:0],u_ca_out_249[35:9], u_ca_out_248[62:36], u_ca_out_247[71:63]};
assign col_out_251 = {u_ca_out_251[8:0],u_ca_out_250[35:9], u_ca_out_249[62:36], u_ca_out_248[71:63]};
assign col_out_252 = {u_ca_out_252[8:0],u_ca_out_251[35:9], u_ca_out_250[62:36], u_ca_out_249[71:63]};
assign col_out_253 = {u_ca_out_253[8:0],u_ca_out_252[35:9], u_ca_out_251[62:36], u_ca_out_250[71:63]};
assign col_out_254 = {u_ca_out_254[8:0],u_ca_out_253[35:9], u_ca_out_252[62:36], u_ca_out_251[71:63]};
assign col_out_255 = {u_ca_out_255[8:0],u_ca_out_254[35:9], u_ca_out_253[62:36], u_ca_out_252[71:63]};
assign col_out_256 = {u_ca_out_256[8:0],u_ca_out_255[35:9], u_ca_out_254[62:36], u_ca_out_253[71:63]};
assign col_out_257 = {u_ca_out_257[8:0],u_ca_out_256[35:9], u_ca_out_255[62:36], u_ca_out_254[71:63]};
assign col_out_258 = {u_ca_out_258[8:0],u_ca_out_257[35:9], u_ca_out_256[62:36], u_ca_out_255[71:63]};
assign col_out_259 = {u_ca_out_259[8:0],u_ca_out_258[35:9], u_ca_out_257[62:36], u_ca_out_256[71:63]};
assign col_out_260 = {u_ca_out_260[8:0],u_ca_out_259[35:9], u_ca_out_258[62:36], u_ca_out_257[71:63]};
assign col_out_261 = {u_ca_out_261[8:0],u_ca_out_260[35:9], u_ca_out_259[62:36], u_ca_out_258[71:63]};
assign col_out_262 = {u_ca_out_262[8:0],u_ca_out_261[35:9], u_ca_out_260[62:36], u_ca_out_259[71:63]};
assign col_out_263 = {u_ca_out_263[8:0],u_ca_out_262[35:9], u_ca_out_261[62:36], u_ca_out_260[71:63]};
assign col_out_264 = {u_ca_out_264[8:0],u_ca_out_263[35:9], u_ca_out_262[62:36], u_ca_out_261[71:63]};
assign col_out_265 = {u_ca_out_265[8:0],u_ca_out_264[35:9], u_ca_out_263[62:36], u_ca_out_262[71:63]};
assign col_out_266 = {u_ca_out_266[8:0],u_ca_out_265[35:9], u_ca_out_264[62:36], u_ca_out_263[71:63]};
assign col_out_267 = {u_ca_out_267[8:0],u_ca_out_266[35:9], u_ca_out_265[62:36], u_ca_out_264[71:63]};
assign col_out_268 = {u_ca_out_268[8:0],u_ca_out_267[35:9], u_ca_out_266[62:36], u_ca_out_265[71:63]};
assign col_out_269 = {u_ca_out_269[8:0],u_ca_out_268[35:9], u_ca_out_267[62:36], u_ca_out_266[71:63]};
assign col_out_270 = {u_ca_out_270[8:0],u_ca_out_269[35:9], u_ca_out_268[62:36], u_ca_out_267[71:63]};
assign col_out_271 = {u_ca_out_271[8:0],u_ca_out_270[35:9], u_ca_out_269[62:36], u_ca_out_268[71:63]};
assign col_out_272 = {u_ca_out_272[8:0],u_ca_out_271[35:9], u_ca_out_270[62:36], u_ca_out_269[71:63]};
assign col_out_273 = {u_ca_out_273[8:0],u_ca_out_272[35:9], u_ca_out_271[62:36], u_ca_out_270[71:63]};
assign col_out_274 = {u_ca_out_274[8:0],u_ca_out_273[35:9], u_ca_out_272[62:36], u_ca_out_271[71:63]};
assign col_out_275 = {u_ca_out_275[8:0],u_ca_out_274[35:9], u_ca_out_273[62:36], u_ca_out_272[71:63]};
assign col_out_276 = {u_ca_out_276[8:0],u_ca_out_275[35:9], u_ca_out_274[62:36], u_ca_out_273[71:63]};
assign col_out_277 = {u_ca_out_277[8:0],u_ca_out_276[35:9], u_ca_out_275[62:36], u_ca_out_274[71:63]};
assign col_out_278 = {u_ca_out_278[8:0],u_ca_out_277[35:9], u_ca_out_276[62:36], u_ca_out_275[71:63]};
assign col_out_279 = {u_ca_out_279[8:0],u_ca_out_278[35:9], u_ca_out_277[62:36], u_ca_out_276[71:63]};
assign col_out_280 = {u_ca_out_280[8:0],u_ca_out_279[35:9], u_ca_out_278[62:36], u_ca_out_277[71:63]};
assign col_out_281 = {u_ca_out_281[8:0],u_ca_out_280[35:9], u_ca_out_279[62:36], u_ca_out_278[71:63]};
assign col_out_282 = {u_ca_out_282[8:0],u_ca_out_281[35:9], u_ca_out_280[62:36], u_ca_out_279[71:63]};
assign col_out_283 = {u_ca_out_283[8:0],u_ca_out_282[35:9], u_ca_out_281[62:36], u_ca_out_280[71:63]};
assign col_out_284 = {u_ca_out_284[8:0],u_ca_out_283[35:9], u_ca_out_282[62:36], u_ca_out_281[71:63]};
assign col_out_285 = {u_ca_out_285[8:0],u_ca_out_284[35:9], u_ca_out_283[62:36], u_ca_out_282[71:63]};
assign col_out_286 = {u_ca_out_286[8:0],u_ca_out_285[35:9], u_ca_out_284[62:36], u_ca_out_283[71:63]};
assign col_out_287 = {u_ca_out_287[8:0],u_ca_out_286[35:9], u_ca_out_285[62:36], u_ca_out_284[71:63]};
assign col_out_288 = {u_ca_out_288[8:0],u_ca_out_287[35:9], u_ca_out_286[62:36], u_ca_out_285[71:63]};
assign col_out_289 = {u_ca_out_289[8:0],u_ca_out_288[35:9], u_ca_out_287[62:36], u_ca_out_286[71:63]};
assign col_out_290 = {u_ca_out_290[8:0],u_ca_out_289[35:9], u_ca_out_288[62:36], u_ca_out_287[71:63]};
assign col_out_291 = {u_ca_out_291[8:0],u_ca_out_290[35:9], u_ca_out_289[62:36], u_ca_out_288[71:63]};
assign col_out_292 = {u_ca_out_292[8:0],u_ca_out_291[35:9], u_ca_out_290[62:36], u_ca_out_289[71:63]};
assign col_out_293 = {u_ca_out_293[8:0],u_ca_out_292[35:9], u_ca_out_291[62:36], u_ca_out_290[71:63]};
assign col_out_294 = {u_ca_out_294[8:0],u_ca_out_293[35:9], u_ca_out_292[62:36], u_ca_out_291[71:63]};
assign col_out_295 = {u_ca_out_295[8:0],u_ca_out_294[35:9], u_ca_out_293[62:36], u_ca_out_292[71:63]};
assign col_out_296 = {u_ca_out_296[8:0],u_ca_out_295[35:9], u_ca_out_294[62:36], u_ca_out_293[71:63]};
assign col_out_297 = {u_ca_out_297[8:0],u_ca_out_296[35:9], u_ca_out_295[62:36], u_ca_out_294[71:63]};
assign col_out_298 = {u_ca_out_298[8:0],u_ca_out_297[35:9], u_ca_out_296[62:36], u_ca_out_295[71:63]};
assign col_out_299 = {u_ca_out_299[8:0],u_ca_out_298[35:9], u_ca_out_297[62:36], u_ca_out_296[71:63]};
assign col_out_300 = {u_ca_out_300[8:0],u_ca_out_299[35:9], u_ca_out_298[62:36], u_ca_out_297[71:63]};
assign col_out_301 = {u_ca_out_301[8:0],u_ca_out_300[35:9], u_ca_out_299[62:36], u_ca_out_298[71:63]};
assign col_out_302 = {u_ca_out_302[8:0],u_ca_out_301[35:9], u_ca_out_300[62:36], u_ca_out_299[71:63]};
assign col_out_303 = {u_ca_out_303[8:0],u_ca_out_302[35:9], u_ca_out_301[62:36], u_ca_out_300[71:63]};
assign col_out_304 = {u_ca_out_304[8:0],u_ca_out_303[35:9], u_ca_out_302[62:36], u_ca_out_301[71:63]};
assign col_out_305 = {u_ca_out_305[8:0],u_ca_out_304[35:9], u_ca_out_303[62:36], u_ca_out_302[71:63]};
assign col_out_306 = {u_ca_out_306[8:0],u_ca_out_305[35:9], u_ca_out_304[62:36], u_ca_out_303[71:63]};
assign col_out_307 = {u_ca_out_307[8:0],u_ca_out_306[35:9], u_ca_out_305[62:36], u_ca_out_304[71:63]};
assign col_out_308 = {u_ca_out_308[8:0],u_ca_out_307[35:9], u_ca_out_306[62:36], u_ca_out_305[71:63]};
assign col_out_309 = {u_ca_out_309[8:0],u_ca_out_308[35:9], u_ca_out_307[62:36], u_ca_out_306[71:63]};
assign col_out_310 = {u_ca_out_310[8:0],u_ca_out_309[35:9], u_ca_out_308[62:36], u_ca_out_307[71:63]};
assign col_out_311 = {u_ca_out_311[8:0],u_ca_out_310[35:9], u_ca_out_309[62:36], u_ca_out_308[71:63]};
assign col_out_312 = {u_ca_out_312[8:0],u_ca_out_311[35:9], u_ca_out_310[62:36], u_ca_out_309[71:63]};
assign col_out_313 = {u_ca_out_313[8:0],u_ca_out_312[35:9], u_ca_out_311[62:36], u_ca_out_310[71:63]};
assign col_out_314 = {u_ca_out_314[8:0],u_ca_out_313[35:9], u_ca_out_312[62:36], u_ca_out_311[71:63]};
assign col_out_315 = {u_ca_out_315[8:0],u_ca_out_314[35:9], u_ca_out_313[62:36], u_ca_out_312[71:63]};
assign col_out_316 = {u_ca_out_316[8:0],u_ca_out_315[35:9], u_ca_out_314[62:36], u_ca_out_313[71:63]};
assign col_out_317 = {u_ca_out_317[8:0],u_ca_out_316[35:9], u_ca_out_315[62:36], u_ca_out_314[71:63]};
assign col_out_318 = {u_ca_out_318[8:0],u_ca_out_317[35:9], u_ca_out_316[62:36], u_ca_out_315[71:63]};
assign col_out_319 = {u_ca_out_319[8:0],u_ca_out_318[35:9], u_ca_out_317[62:36], u_ca_out_316[71:63]};
assign col_out_320 = {u_ca_out_320[8:0],u_ca_out_319[35:9], u_ca_out_318[62:36], u_ca_out_317[71:63]};
assign col_out_321 = {u_ca_out_321[8:0],u_ca_out_320[35:9], u_ca_out_319[62:36], u_ca_out_318[71:63]};
assign col_out_322 = {u_ca_out_322[8:0],u_ca_out_321[35:9], u_ca_out_320[62:36], u_ca_out_319[71:63]};
assign col_out_323 = {u_ca_out_323[8:0],u_ca_out_322[35:9], u_ca_out_321[62:36], u_ca_out_320[71:63]};
assign col_out_324 = {u_ca_out_324[8:0],u_ca_out_323[35:9], u_ca_out_322[62:36], u_ca_out_321[71:63]};
assign col_out_325 = {u_ca_out_325[8:0],u_ca_out_324[35:9], u_ca_out_323[62:36], u_ca_out_322[71:63]};
assign col_out_326 = {u_ca_out_326[8:0],u_ca_out_325[35:9], u_ca_out_324[62:36], u_ca_out_323[71:63]};
assign col_out_327 = {u_ca_out_327[8:0],u_ca_out_326[35:9], u_ca_out_325[62:36], u_ca_out_324[71:63]};
assign col_out_328 = {u_ca_out_328[8:0],u_ca_out_327[35:9], u_ca_out_326[62:36], u_ca_out_325[71:63]};
assign col_out_329 = {u_ca_out_329[8:0],u_ca_out_328[35:9], u_ca_out_327[62:36], u_ca_out_326[71:63]};
assign col_out_330 = {u_ca_out_330[8:0],u_ca_out_329[35:9], u_ca_out_328[62:36], u_ca_out_327[71:63]};
assign col_out_331 = {u_ca_out_331[8:0],u_ca_out_330[35:9], u_ca_out_329[62:36], u_ca_out_328[71:63]};
assign col_out_332 = {u_ca_out_332[8:0],u_ca_out_331[35:9], u_ca_out_330[62:36], u_ca_out_329[71:63]};
assign col_out_333 = {u_ca_out_333[8:0],u_ca_out_332[35:9], u_ca_out_331[62:36], u_ca_out_330[71:63]};
assign col_out_334 = {u_ca_out_334[8:0],u_ca_out_333[35:9], u_ca_out_332[62:36], u_ca_out_331[71:63]};
assign col_out_335 = {u_ca_out_335[8:0],u_ca_out_334[35:9], u_ca_out_333[62:36], u_ca_out_332[71:63]};
assign col_out_336 = {u_ca_out_336[8:0],u_ca_out_335[35:9], u_ca_out_334[62:36], u_ca_out_333[71:63]};
assign col_out_337 = {u_ca_out_337[8:0],u_ca_out_336[35:9], u_ca_out_335[62:36], u_ca_out_334[71:63]};
assign col_out_338 = {u_ca_out_338[8:0],u_ca_out_337[35:9], u_ca_out_336[62:36], u_ca_out_335[71:63]};
assign col_out_339 = {u_ca_out_339[8:0],u_ca_out_338[35:9], u_ca_out_337[62:36], u_ca_out_336[71:63]};
assign col_out_340 = {u_ca_out_340[8:0],u_ca_out_339[35:9], u_ca_out_338[62:36], u_ca_out_337[71:63]};
assign col_out_341 = {u_ca_out_341[8:0],u_ca_out_340[35:9], u_ca_out_339[62:36], u_ca_out_338[71:63]};
assign col_out_342 = {u_ca_out_342[8:0],u_ca_out_341[35:9], u_ca_out_340[62:36], u_ca_out_339[71:63]};
assign col_out_343 = {u_ca_out_343[8:0],u_ca_out_342[35:9], u_ca_out_341[62:36], u_ca_out_340[71:63]};
assign col_out_344 = {u_ca_out_344[8:0],u_ca_out_343[35:9], u_ca_out_342[62:36], u_ca_out_341[71:63]};
assign col_out_345 = {u_ca_out_345[8:0],u_ca_out_344[35:9], u_ca_out_343[62:36], u_ca_out_342[71:63]};
assign col_out_346 = {u_ca_out_346[8:0],u_ca_out_345[35:9], u_ca_out_344[62:36], u_ca_out_343[71:63]};
assign col_out_347 = {u_ca_out_347[8:0],u_ca_out_346[35:9], u_ca_out_345[62:36], u_ca_out_344[71:63]};
assign col_out_348 = {u_ca_out_348[8:0],u_ca_out_347[35:9], u_ca_out_346[62:36], u_ca_out_345[71:63]};
assign col_out_349 = {u_ca_out_349[8:0],u_ca_out_348[35:9], u_ca_out_347[62:36], u_ca_out_346[71:63]};
assign col_out_350 = {u_ca_out_350[8:0],u_ca_out_349[35:9], u_ca_out_348[62:36], u_ca_out_347[71:63]};
assign col_out_351 = {u_ca_out_351[8:0],u_ca_out_350[35:9], u_ca_out_349[62:36], u_ca_out_348[71:63]};
assign col_out_352 = {u_ca_out_352[8:0],u_ca_out_351[35:9], u_ca_out_350[62:36], u_ca_out_349[71:63]};
assign col_out_353 = {u_ca_out_353[8:0],u_ca_out_352[35:9], u_ca_out_351[62:36], u_ca_out_350[71:63]};
assign col_out_354 = {u_ca_out_354[8:0],u_ca_out_353[35:9], u_ca_out_352[62:36], u_ca_out_351[71:63]};
assign col_out_355 = {u_ca_out_355[8:0],u_ca_out_354[35:9], u_ca_out_353[62:36], u_ca_out_352[71:63]};
assign col_out_356 = {u_ca_out_356[8:0],u_ca_out_355[35:9], u_ca_out_354[62:36], u_ca_out_353[71:63]};
assign col_out_357 = {u_ca_out_357[8:0],u_ca_out_356[35:9], u_ca_out_355[62:36], u_ca_out_354[71:63]};
assign col_out_358 = {u_ca_out_358[8:0],u_ca_out_357[35:9], u_ca_out_356[62:36], u_ca_out_355[71:63]};
assign col_out_359 = {u_ca_out_359[8:0],u_ca_out_358[35:9], u_ca_out_357[62:36], u_ca_out_356[71:63]};
assign col_out_360 = {u_ca_out_360[8:0],u_ca_out_359[35:9], u_ca_out_358[62:36], u_ca_out_357[71:63]};
assign col_out_361 = {u_ca_out_361[8:0],u_ca_out_360[35:9], u_ca_out_359[62:36], u_ca_out_358[71:63]};
assign col_out_362 = {u_ca_out_362[8:0],u_ca_out_361[35:9], u_ca_out_360[62:36], u_ca_out_359[71:63]};
assign col_out_363 = {u_ca_out_363[8:0],u_ca_out_362[35:9], u_ca_out_361[62:36], u_ca_out_360[71:63]};
assign col_out_364 = {u_ca_out_364[8:0],u_ca_out_363[35:9], u_ca_out_362[62:36], u_ca_out_361[71:63]};
assign col_out_365 = {u_ca_out_365[8:0],u_ca_out_364[35:9], u_ca_out_363[62:36], u_ca_out_362[71:63]};
assign col_out_366 = {u_ca_out_366[8:0],u_ca_out_365[35:9], u_ca_out_364[62:36], u_ca_out_363[71:63]};
assign col_out_367 = {u_ca_out_367[8:0],u_ca_out_366[35:9], u_ca_out_365[62:36], u_ca_out_364[71:63]};
assign col_out_368 = {u_ca_out_368[8:0],u_ca_out_367[35:9], u_ca_out_366[62:36], u_ca_out_365[71:63]};
assign col_out_369 = {u_ca_out_369[8:0],u_ca_out_368[35:9], u_ca_out_367[62:36], u_ca_out_366[71:63]};
assign col_out_370 = {u_ca_out_370[8:0],u_ca_out_369[35:9], u_ca_out_368[62:36], u_ca_out_367[71:63]};
assign col_out_371 = {u_ca_out_371[8:0],u_ca_out_370[35:9], u_ca_out_369[62:36], u_ca_out_368[71:63]};
assign col_out_372 = {u_ca_out_372[8:0],u_ca_out_371[35:9], u_ca_out_370[62:36], u_ca_out_369[71:63]};
assign col_out_373 = {u_ca_out_373[8:0],u_ca_out_372[35:9], u_ca_out_371[62:36], u_ca_out_370[71:63]};
assign col_out_374 = {u_ca_out_374[8:0],u_ca_out_373[35:9], u_ca_out_372[62:36], u_ca_out_371[71:63]};
assign col_out_375 = {u_ca_out_375[8:0],u_ca_out_374[35:9], u_ca_out_373[62:36], u_ca_out_372[71:63]};
assign col_out_376 = {u_ca_out_376[8:0],u_ca_out_375[35:9], u_ca_out_374[62:36], u_ca_out_373[71:63]};
assign col_out_377 = {u_ca_out_377[8:0],u_ca_out_376[35:9], u_ca_out_375[62:36], u_ca_out_374[71:63]};
assign col_out_378 = {u_ca_out_378[8:0],u_ca_out_377[35:9], u_ca_out_376[62:36], u_ca_out_375[71:63]};
assign col_out_379 = {u_ca_out_379[8:0],u_ca_out_378[35:9], u_ca_out_377[62:36], u_ca_out_376[71:63]};
assign col_out_380 = {u_ca_out_380[8:0],u_ca_out_379[35:9], u_ca_out_378[62:36], u_ca_out_377[71:63]};
assign col_out_381 = {u_ca_out_381[8:0],u_ca_out_380[35:9], u_ca_out_379[62:36], u_ca_out_378[71:63]};
assign col_out_382 = {u_ca_out_382[8:0],u_ca_out_381[35:9], u_ca_out_380[62:36], u_ca_out_379[71:63]};
assign col_out_383 = {u_ca_out_383[8:0],u_ca_out_382[35:9], u_ca_out_381[62:36], u_ca_out_380[71:63]};
assign col_out_384 = {u_ca_out_384[8:0],u_ca_out_383[35:9], u_ca_out_382[62:36], u_ca_out_381[71:63]};
assign col_out_385 = {u_ca_out_385[8:0],u_ca_out_384[35:9], u_ca_out_383[62:36], u_ca_out_382[71:63]};
assign col_out_386 = {u_ca_out_386[8:0],u_ca_out_385[35:9], u_ca_out_384[62:36], u_ca_out_383[71:63]};
assign col_out_387 = {u_ca_out_387[8:0],u_ca_out_386[35:9], u_ca_out_385[62:36], u_ca_out_384[71:63]};
assign col_out_388 = {u_ca_out_388[8:0],u_ca_out_387[35:9], u_ca_out_386[62:36], u_ca_out_385[71:63]};
assign col_out_389 = {u_ca_out_389[8:0],u_ca_out_388[35:9], u_ca_out_387[62:36], u_ca_out_386[71:63]};
assign col_out_390 = {u_ca_out_390[8:0],u_ca_out_389[35:9], u_ca_out_388[62:36], u_ca_out_387[71:63]};
assign col_out_391 = {u_ca_out_391[8:0],u_ca_out_390[35:9], u_ca_out_389[62:36], u_ca_out_388[71:63]};
assign col_out_392 = {u_ca_out_392[8:0],u_ca_out_391[35:9], u_ca_out_390[62:36], u_ca_out_389[71:63]};
assign col_out_393 = {u_ca_out_393[8:0],u_ca_out_392[35:9], u_ca_out_391[62:36], u_ca_out_390[71:63]};
assign col_out_394 = {u_ca_out_394[8:0],u_ca_out_393[35:9], u_ca_out_392[62:36], u_ca_out_391[71:63]};
assign col_out_395 = {u_ca_out_395[8:0],u_ca_out_394[35:9], u_ca_out_393[62:36], u_ca_out_392[71:63]};
assign col_out_396 = {u_ca_out_396[8:0],u_ca_out_395[35:9], u_ca_out_394[62:36], u_ca_out_393[71:63]};
assign col_out_397 = {u_ca_out_397[8:0],u_ca_out_396[35:9], u_ca_out_395[62:36], u_ca_out_394[71:63]};
assign col_out_398 = {u_ca_out_398[8:0],u_ca_out_397[35:9], u_ca_out_396[62:36], u_ca_out_395[71:63]};
assign col_out_399 = {u_ca_out_399[8:0],u_ca_out_398[35:9], u_ca_out_397[62:36], u_ca_out_396[71:63]};
assign col_out_400 = {u_ca_out_400[8:0],u_ca_out_399[35:9], u_ca_out_398[62:36], u_ca_out_397[71:63]};
assign col_out_401 = {u_ca_out_401[8:0],u_ca_out_400[35:9], u_ca_out_399[62:36], u_ca_out_398[71:63]};
assign col_out_402 = {u_ca_out_402[8:0],u_ca_out_401[35:9], u_ca_out_400[62:36], u_ca_out_399[71:63]};
assign col_out_403 = {u_ca_out_403[8:0],u_ca_out_402[35:9], u_ca_out_401[62:36], u_ca_out_400[71:63]};
assign col_out_404 = {u_ca_out_404[8:0],u_ca_out_403[35:9], u_ca_out_402[62:36], u_ca_out_401[71:63]};
assign col_out_405 = {u_ca_out_405[8:0],u_ca_out_404[35:9], u_ca_out_403[62:36], u_ca_out_402[71:63]};
assign col_out_406 = {u_ca_out_406[8:0],u_ca_out_405[35:9], u_ca_out_404[62:36], u_ca_out_403[71:63]};
assign col_out_407 = {u_ca_out_407[8:0],u_ca_out_406[35:9], u_ca_out_405[62:36], u_ca_out_404[71:63]};
assign col_out_408 = {u_ca_out_408[8:0],u_ca_out_407[35:9], u_ca_out_406[62:36], u_ca_out_405[71:63]};
assign col_out_409 = {u_ca_out_409[8:0],u_ca_out_408[35:9], u_ca_out_407[62:36], u_ca_out_406[71:63]};
assign col_out_410 = {u_ca_out_410[8:0],u_ca_out_409[35:9], u_ca_out_408[62:36], u_ca_out_407[71:63]};
assign col_out_411 = {u_ca_out_411[8:0],u_ca_out_410[35:9], u_ca_out_409[62:36], u_ca_out_408[71:63]};
assign col_out_412 = {u_ca_out_412[8:0],u_ca_out_411[35:9], u_ca_out_410[62:36], u_ca_out_409[71:63]};
assign col_out_413 = {u_ca_out_413[8:0],u_ca_out_412[35:9], u_ca_out_411[62:36], u_ca_out_410[71:63]};
assign col_out_414 = {u_ca_out_414[8:0],u_ca_out_413[35:9], u_ca_out_412[62:36], u_ca_out_411[71:63]};
assign col_out_415 = {u_ca_out_415[8:0],u_ca_out_414[35:9], u_ca_out_413[62:36], u_ca_out_412[71:63]};
assign col_out_416 = {u_ca_out_416[8:0],u_ca_out_415[35:9], u_ca_out_414[62:36], u_ca_out_413[71:63]};
assign col_out_417 = {u_ca_out_417[8:0],u_ca_out_416[35:9], u_ca_out_415[62:36], u_ca_out_414[71:63]};
assign col_out_418 = {u_ca_out_418[8:0],u_ca_out_417[35:9], u_ca_out_416[62:36], u_ca_out_415[71:63]};
assign col_out_419 = {u_ca_out_419[8:0],u_ca_out_418[35:9], u_ca_out_417[62:36], u_ca_out_416[71:63]};
assign col_out_420 = {u_ca_out_420[8:0],u_ca_out_419[35:9], u_ca_out_418[62:36], u_ca_out_417[71:63]};
assign col_out_421 = {u_ca_out_421[8:0],u_ca_out_420[35:9], u_ca_out_419[62:36], u_ca_out_418[71:63]};
assign col_out_422 = {u_ca_out_422[8:0],u_ca_out_421[35:9], u_ca_out_420[62:36], u_ca_out_419[71:63]};
assign col_out_423 = {u_ca_out_423[8:0],u_ca_out_422[35:9], u_ca_out_421[62:36], u_ca_out_420[71:63]};
assign col_out_424 = {u_ca_out_424[8:0],u_ca_out_423[35:9], u_ca_out_422[62:36], u_ca_out_421[71:63]};
assign col_out_425 = {u_ca_out_425[8:0],u_ca_out_424[35:9], u_ca_out_423[62:36], u_ca_out_422[71:63]};
assign col_out_426 = {u_ca_out_426[8:0],u_ca_out_425[35:9], u_ca_out_424[62:36], u_ca_out_423[71:63]};
assign col_out_427 = {u_ca_out_427[8:0],u_ca_out_426[35:9], u_ca_out_425[62:36], u_ca_out_424[71:63]};
assign col_out_428 = {u_ca_out_428[8:0],u_ca_out_427[35:9], u_ca_out_426[62:36], u_ca_out_425[71:63]};
assign col_out_429 = {u_ca_out_429[8:0],u_ca_out_428[35:9], u_ca_out_427[62:36], u_ca_out_426[71:63]};
assign col_out_430 = {u_ca_out_430[8:0],u_ca_out_429[35:9], u_ca_out_428[62:36], u_ca_out_427[71:63]};
assign col_out_431 = {u_ca_out_431[8:0],u_ca_out_430[35:9], u_ca_out_429[62:36], u_ca_out_428[71:63]};
assign col_out_432 = {u_ca_out_432[8:0],u_ca_out_431[35:9], u_ca_out_430[62:36], u_ca_out_429[71:63]};
assign col_out_433 = {u_ca_out_433[8:0],u_ca_out_432[35:9], u_ca_out_431[62:36], u_ca_out_430[71:63]};
assign col_out_434 = {u_ca_out_434[8:0],u_ca_out_433[35:9], u_ca_out_432[62:36], u_ca_out_431[71:63]};
assign col_out_435 = {u_ca_out_435[8:0],u_ca_out_434[35:9], u_ca_out_433[62:36], u_ca_out_432[71:63]};
assign col_out_436 = {u_ca_out_436[8:0],u_ca_out_435[35:9], u_ca_out_434[62:36], u_ca_out_433[71:63]};
assign col_out_437 = {u_ca_out_437[8:0],u_ca_out_436[35:9], u_ca_out_435[62:36], u_ca_out_434[71:63]};
assign col_out_438 = {u_ca_out_438[8:0],u_ca_out_437[35:9], u_ca_out_436[62:36], u_ca_out_435[71:63]};
assign col_out_439 = {u_ca_out_439[8:0],u_ca_out_438[35:9], u_ca_out_437[62:36], u_ca_out_436[71:63]};
assign col_out_440 = {u_ca_out_440[8:0],u_ca_out_439[35:9], u_ca_out_438[62:36], u_ca_out_437[71:63]};
assign col_out_441 = {u_ca_out_441[8:0],u_ca_out_440[35:9], u_ca_out_439[62:36], u_ca_out_438[71:63]};
assign col_out_442 = {u_ca_out_442[8:0],u_ca_out_441[35:9], u_ca_out_440[62:36], u_ca_out_439[71:63]};
assign col_out_443 = {u_ca_out_443[8:0],u_ca_out_442[35:9], u_ca_out_441[62:36], u_ca_out_440[71:63]};
assign col_out_444 = {u_ca_out_444[8:0],u_ca_out_443[35:9], u_ca_out_442[62:36], u_ca_out_441[71:63]};
assign col_out_445 = {u_ca_out_445[8:0],u_ca_out_444[35:9], u_ca_out_443[62:36], u_ca_out_442[71:63]};
assign col_out_446 = {u_ca_out_446[8:0],u_ca_out_445[35:9], u_ca_out_444[62:36], u_ca_out_443[71:63]};
assign col_out_447 = {u_ca_out_447[8:0],u_ca_out_446[35:9], u_ca_out_445[62:36], u_ca_out_444[71:63]};
assign col_out_448 = {u_ca_out_448[8:0],u_ca_out_447[35:9], u_ca_out_446[62:36], u_ca_out_445[71:63]};
assign col_out_449 = {u_ca_out_449[8:0],u_ca_out_448[35:9], u_ca_out_447[62:36], u_ca_out_446[71:63]};
assign col_out_450 = {u_ca_out_450[8:0],u_ca_out_449[35:9], u_ca_out_448[62:36], u_ca_out_447[71:63]};
assign col_out_451 = {u_ca_out_451[8:0],u_ca_out_450[35:9], u_ca_out_449[62:36], u_ca_out_448[71:63]};
assign col_out_452 = {u_ca_out_452[8:0],u_ca_out_451[35:9], u_ca_out_450[62:36], u_ca_out_449[71:63]};
assign col_out_453 = {u_ca_out_453[8:0],u_ca_out_452[35:9], u_ca_out_451[62:36], u_ca_out_450[71:63]};
assign col_out_454 = {u_ca_out_454[8:0],u_ca_out_453[35:9], u_ca_out_452[62:36], u_ca_out_451[71:63]};
assign col_out_455 = {u_ca_out_455[8:0],u_ca_out_454[35:9], u_ca_out_453[62:36], u_ca_out_452[71:63]};
assign col_out_456 = {u_ca_out_456[8:0],u_ca_out_455[35:9], u_ca_out_454[62:36], u_ca_out_453[71:63]};
assign col_out_457 = {u_ca_out_457[8:0],u_ca_out_456[35:9], u_ca_out_455[62:36], u_ca_out_454[71:63]};
assign col_out_458 = {u_ca_out_458[8:0],u_ca_out_457[35:9], u_ca_out_456[62:36], u_ca_out_455[71:63]};
assign col_out_459 = {u_ca_out_459[8:0],u_ca_out_458[35:9], u_ca_out_457[62:36], u_ca_out_456[71:63]};
assign col_out_460 = {u_ca_out_460[8:0],u_ca_out_459[35:9], u_ca_out_458[62:36], u_ca_out_457[71:63]};
assign col_out_461 = {u_ca_out_461[8:0],u_ca_out_460[35:9], u_ca_out_459[62:36], u_ca_out_458[71:63]};
assign col_out_462 = {u_ca_out_462[8:0],u_ca_out_461[35:9], u_ca_out_460[62:36], u_ca_out_459[71:63]};
assign col_out_463 = {u_ca_out_463[8:0],u_ca_out_462[35:9], u_ca_out_461[62:36], u_ca_out_460[71:63]};
assign col_out_464 = {u_ca_out_464[8:0],u_ca_out_463[35:9], u_ca_out_462[62:36], u_ca_out_461[71:63]};
assign col_out_465 = {u_ca_out_465[8:0],u_ca_out_464[35:9], u_ca_out_463[62:36], u_ca_out_462[71:63]};
assign col_out_466 = {u_ca_out_466[8:0],u_ca_out_465[35:9], u_ca_out_464[62:36], u_ca_out_463[71:63]};
assign col_out_467 = {u_ca_out_467[8:0],u_ca_out_466[35:9], u_ca_out_465[62:36], u_ca_out_464[71:63]};
assign col_out_468 = {u_ca_out_468[8:0],u_ca_out_467[35:9], u_ca_out_466[62:36], u_ca_out_465[71:63]};
assign col_out_469 = {u_ca_out_469[8:0],u_ca_out_468[35:9], u_ca_out_467[62:36], u_ca_out_466[71:63]};
assign col_out_470 = {u_ca_out_470[8:0],u_ca_out_469[35:9], u_ca_out_468[62:36], u_ca_out_467[71:63]};
assign col_out_471 = {u_ca_out_471[8:0],u_ca_out_470[35:9], u_ca_out_469[62:36], u_ca_out_468[71:63]};
assign col_out_472 = {u_ca_out_472[8:0],u_ca_out_471[35:9], u_ca_out_470[62:36], u_ca_out_469[71:63]};
assign col_out_473 = {u_ca_out_473[8:0],u_ca_out_472[35:9], u_ca_out_471[62:36], u_ca_out_470[71:63]};
assign col_out_474 = {u_ca_out_474[8:0],u_ca_out_473[35:9], u_ca_out_472[62:36], u_ca_out_471[71:63]};
assign col_out_475 = {u_ca_out_475[8:0],u_ca_out_474[35:9], u_ca_out_473[62:36], u_ca_out_472[71:63]};
assign col_out_476 = {u_ca_out_476[8:0],u_ca_out_475[35:9], u_ca_out_474[62:36], u_ca_out_473[71:63]};
assign col_out_477 = {u_ca_out_477[8:0],u_ca_out_476[35:9], u_ca_out_475[62:36], u_ca_out_474[71:63]};
assign col_out_478 = {u_ca_out_478[8:0],u_ca_out_477[35:9], u_ca_out_476[62:36], u_ca_out_475[71:63]};
assign col_out_479 = {u_ca_out_479[8:0],u_ca_out_478[35:9], u_ca_out_477[62:36], u_ca_out_476[71:63]};
assign col_out_480 = {u_ca_out_480[8:0],u_ca_out_479[35:9], u_ca_out_478[62:36], u_ca_out_477[71:63]};
assign col_out_481 = {u_ca_out_481[8:0],u_ca_out_480[35:9], u_ca_out_479[62:36], u_ca_out_478[71:63]};
assign col_out_482 = {u_ca_out_482[8:0],u_ca_out_481[35:9], u_ca_out_480[62:36], u_ca_out_479[71:63]};
assign col_out_483 = {u_ca_out_483[8:0],u_ca_out_482[35:9], u_ca_out_481[62:36], u_ca_out_480[71:63]};
assign col_out_484 = {u_ca_out_484[8:0],u_ca_out_483[35:9], u_ca_out_482[62:36], u_ca_out_481[71:63]};
assign col_out_485 = {u_ca_out_485[8:0],u_ca_out_484[35:9], u_ca_out_483[62:36], u_ca_out_482[71:63]};
assign col_out_486 = {u_ca_out_486[8:0],u_ca_out_485[35:9], u_ca_out_484[62:36], u_ca_out_483[71:63]};
assign col_out_487 = {u_ca_out_487[8:0],u_ca_out_486[35:9], u_ca_out_485[62:36], u_ca_out_484[71:63]};
assign col_out_488 = {u_ca_out_488[8:0],u_ca_out_487[35:9], u_ca_out_486[62:36], u_ca_out_485[71:63]};
assign col_out_489 = {u_ca_out_489[8:0],u_ca_out_488[35:9], u_ca_out_487[62:36], u_ca_out_486[71:63]};
assign col_out_490 = {u_ca_out_490[8:0],u_ca_out_489[35:9], u_ca_out_488[62:36], u_ca_out_487[71:63]};
assign col_out_491 = {u_ca_out_491[8:0],u_ca_out_490[35:9], u_ca_out_489[62:36], u_ca_out_488[71:63]};
assign col_out_492 = {u_ca_out_492[8:0],u_ca_out_491[35:9], u_ca_out_490[62:36], u_ca_out_489[71:63]};
assign col_out_493 = {u_ca_out_493[8:0],u_ca_out_492[35:9], u_ca_out_491[62:36], u_ca_out_490[71:63]};
assign col_out_494 = {u_ca_out_494[8:0],u_ca_out_493[35:9], u_ca_out_492[62:36], u_ca_out_491[71:63]};
assign col_out_495 = {u_ca_out_495[8:0],u_ca_out_494[35:9], u_ca_out_493[62:36], u_ca_out_492[71:63]};
assign col_out_496 = {u_ca_out_496[8:0],u_ca_out_495[35:9], u_ca_out_494[62:36], u_ca_out_493[71:63]};
assign col_out_497 = {u_ca_out_497[8:0],u_ca_out_496[35:9], u_ca_out_495[62:36], u_ca_out_494[71:63]};
assign col_out_498 = {u_ca_out_498[8:0],u_ca_out_497[35:9], u_ca_out_496[62:36], u_ca_out_495[71:63]};
assign col_out_499 = {u_ca_out_499[8:0],u_ca_out_498[35:9], u_ca_out_497[62:36], u_ca_out_496[71:63]};
assign col_out_500 = {u_ca_out_500[8:0],u_ca_out_499[35:9], u_ca_out_498[62:36], u_ca_out_497[71:63]};
assign col_out_501 = {u_ca_out_501[8:0],u_ca_out_500[35:9], u_ca_out_499[62:36], u_ca_out_498[71:63]};
assign col_out_502 = {u_ca_out_502[8:0],u_ca_out_501[35:9], u_ca_out_500[62:36], u_ca_out_499[71:63]};
assign col_out_503 = {u_ca_out_503[8:0],u_ca_out_502[35:9], u_ca_out_501[62:36], u_ca_out_500[71:63]};
assign col_out_504 = {u_ca_out_504[8:0],u_ca_out_503[35:9], u_ca_out_502[62:36], u_ca_out_501[71:63]};
assign col_out_505 = {u_ca_out_505[8:0],u_ca_out_504[35:9], u_ca_out_503[62:36], u_ca_out_502[71:63]};
assign col_out_506 = {u_ca_out_506[8:0],u_ca_out_505[35:9], u_ca_out_504[62:36], u_ca_out_503[71:63]};
assign col_out_507 = {u_ca_out_507[8:0],u_ca_out_506[35:9], u_ca_out_505[62:36], u_ca_out_504[71:63]};
assign col_out_508 = {u_ca_out_508[8:0],u_ca_out_507[35:9], u_ca_out_506[62:36], u_ca_out_505[71:63]};
assign col_out_509 = {u_ca_out_509[8:0],u_ca_out_508[35:9], u_ca_out_507[62:36], u_ca_out_506[71:63]};
assign col_out_510 = {u_ca_out_510[8:0],u_ca_out_509[35:9], u_ca_out_508[62:36], u_ca_out_507[71:63]};
assign col_out_511 = {u_ca_out_511[8:0],u_ca_out_510[35:9], u_ca_out_509[62:36], u_ca_out_508[71:63]};
assign col_out_512 = {u_ca_out_512[8:0],u_ca_out_511[35:9], u_ca_out_510[62:36], u_ca_out_509[71:63]};
assign col_out_513 = {u_ca_out_513[8:0],u_ca_out_512[35:9], u_ca_out_511[62:36], u_ca_out_510[71:63]};
assign col_out_514 = {u_ca_out_514[8:0],u_ca_out_513[35:9], u_ca_out_512[62:36], u_ca_out_511[71:63]};
assign col_out_515 = {u_ca_out_515[8:0],u_ca_out_514[35:9], u_ca_out_513[62:36], u_ca_out_512[71:63]};
assign col_out_516 = {u_ca_out_516[8:0],u_ca_out_515[35:9], u_ca_out_514[62:36], u_ca_out_513[71:63]};
assign col_out_517 = {u_ca_out_517[8:0],u_ca_out_516[35:9], u_ca_out_515[62:36], u_ca_out_514[71:63]};
assign col_out_518 = {u_ca_out_518[8:0],u_ca_out_517[35:9], u_ca_out_516[62:36], u_ca_out_515[71:63]};
assign col_out_519 = {u_ca_out_519[8:0],u_ca_out_518[35:9], u_ca_out_517[62:36], u_ca_out_516[71:63]};
assign col_out_520 = {u_ca_out_520[8:0],u_ca_out_519[35:9], u_ca_out_518[62:36], u_ca_out_517[71:63]};
assign col_out_521 = {u_ca_out_521[8:0],u_ca_out_520[35:9], u_ca_out_519[62:36], u_ca_out_518[71:63]};
assign col_out_522 = {u_ca_out_522[8:0],u_ca_out_521[35:9], u_ca_out_520[62:36], u_ca_out_519[71:63]};
assign col_out_523 = {u_ca_out_523[8:0],u_ca_out_522[35:9], u_ca_out_521[62:36], u_ca_out_520[71:63]};
assign col_out_524 = {u_ca_out_524[8:0],u_ca_out_523[35:9], u_ca_out_522[62:36], u_ca_out_521[71:63]};
assign col_out_525 = {u_ca_out_525[8:0],u_ca_out_524[35:9], u_ca_out_523[62:36], u_ca_out_522[71:63]};
assign col_out_526 = {u_ca_out_526[8:0],u_ca_out_525[35:9], u_ca_out_524[62:36], u_ca_out_523[71:63]};
assign col_out_527 = {u_ca_out_527[8:0],u_ca_out_526[35:9], u_ca_out_525[62:36], u_ca_out_524[71:63]};
assign col_out_528 = {u_ca_out_528[8:0],u_ca_out_527[35:9], u_ca_out_526[62:36], u_ca_out_525[71:63]};
assign col_out_529 = {u_ca_out_529[8:0],u_ca_out_528[35:9], u_ca_out_527[62:36], u_ca_out_526[71:63]};
assign col_out_530 = {u_ca_out_530[8:0],u_ca_out_529[35:9], u_ca_out_528[62:36], u_ca_out_527[71:63]};
assign col_out_531 = {u_ca_out_531[8:0],u_ca_out_530[35:9], u_ca_out_529[62:36], u_ca_out_528[71:63]};
assign col_out_532 = {u_ca_out_532[8:0],u_ca_out_531[35:9], u_ca_out_530[62:36], u_ca_out_529[71:63]};
assign col_out_533 = {u_ca_out_533[8:0],u_ca_out_532[35:9], u_ca_out_531[62:36], u_ca_out_530[71:63]};
assign col_out_534 = {u_ca_out_534[8:0],u_ca_out_533[35:9], u_ca_out_532[62:36], u_ca_out_531[71:63]};
assign col_out_535 = {u_ca_out_535[8:0],u_ca_out_534[35:9], u_ca_out_533[62:36], u_ca_out_532[71:63]};
assign col_out_536 = {u_ca_out_536[8:0],u_ca_out_535[35:9], u_ca_out_534[62:36], u_ca_out_533[71:63]};
assign col_out_537 = {u_ca_out_537[8:0],u_ca_out_536[35:9], u_ca_out_535[62:36], u_ca_out_534[71:63]};
assign col_out_538 = {u_ca_out_538[8:0],u_ca_out_537[35:9], u_ca_out_536[62:36], u_ca_out_535[71:63]};
assign col_out_539 = {u_ca_out_539[8:0],u_ca_out_538[35:9], u_ca_out_537[62:36], u_ca_out_536[71:63]};
assign col_out_540 = {u_ca_out_540[8:0],u_ca_out_539[35:9], u_ca_out_538[62:36], u_ca_out_537[71:63]};
assign col_out_541 = {u_ca_out_541[8:0],u_ca_out_540[35:9], u_ca_out_539[62:36], u_ca_out_538[71:63]};
assign col_out_542 = {u_ca_out_542[8:0],u_ca_out_541[35:9], u_ca_out_540[62:36], u_ca_out_539[71:63]};
assign col_out_543 = {u_ca_out_543[8:0],u_ca_out_542[35:9], u_ca_out_541[62:36], u_ca_out_540[71:63]};
assign col_out_544 = {u_ca_out_544[8:0],u_ca_out_543[35:9], u_ca_out_542[62:36], u_ca_out_541[71:63]};
assign col_out_545 = {u_ca_out_545[8:0],u_ca_out_544[35:9], u_ca_out_543[62:36], u_ca_out_542[71:63]};
assign col_out_546 = {u_ca_out_546[8:0],u_ca_out_545[35:9], u_ca_out_544[62:36], u_ca_out_543[71:63]};
assign col_out_547 = {u_ca_out_547[8:0],u_ca_out_546[35:9], u_ca_out_545[62:36], u_ca_out_544[71:63]};
assign col_out_548 = {u_ca_out_548[8:0],u_ca_out_547[35:9], u_ca_out_546[62:36], u_ca_out_545[71:63]};
assign col_out_549 = {u_ca_out_549[8:0],u_ca_out_548[35:9], u_ca_out_547[62:36], u_ca_out_546[71:63]};
assign col_out_550 = {u_ca_out_550[8:0],u_ca_out_549[35:9], u_ca_out_548[62:36], u_ca_out_547[71:63]};
assign col_out_551 = {u_ca_out_551[8:0],u_ca_out_550[35:9], u_ca_out_549[62:36], u_ca_out_548[71:63]};
assign col_out_552 = {u_ca_out_552[8:0],u_ca_out_551[35:9], u_ca_out_550[62:36], u_ca_out_549[71:63]};
assign col_out_553 = {u_ca_out_553[8:0],u_ca_out_552[35:9], u_ca_out_551[62:36], u_ca_out_550[71:63]};
assign col_out_554 = {u_ca_out_554[8:0],u_ca_out_553[35:9], u_ca_out_552[62:36], u_ca_out_551[71:63]};
assign col_out_555 = {u_ca_out_555[8:0],u_ca_out_554[35:9], u_ca_out_553[62:36], u_ca_out_552[71:63]};
assign col_out_556 = {u_ca_out_556[8:0],u_ca_out_555[35:9], u_ca_out_554[62:36], u_ca_out_553[71:63]};
assign col_out_557 = {u_ca_out_557[8:0],u_ca_out_556[35:9], u_ca_out_555[62:36], u_ca_out_554[71:63]};
assign col_out_558 = {u_ca_out_558[8:0],u_ca_out_557[35:9], u_ca_out_556[62:36], u_ca_out_555[71:63]};
assign col_out_559 = {u_ca_out_559[8:0],u_ca_out_558[35:9], u_ca_out_557[62:36], u_ca_out_556[71:63]};
assign col_out_560 = {u_ca_out_560[8:0],u_ca_out_559[35:9], u_ca_out_558[62:36], u_ca_out_557[71:63]};
assign col_out_561 = {u_ca_out_561[8:0],u_ca_out_560[35:9], u_ca_out_559[62:36], u_ca_out_558[71:63]};
assign col_out_562 = {u_ca_out_562[8:0],u_ca_out_561[35:9], u_ca_out_560[62:36], u_ca_out_559[71:63]};
assign col_out_563 = {u_ca_out_563[8:0],u_ca_out_562[35:9], u_ca_out_561[62:36], u_ca_out_560[71:63]};
assign col_out_564 = {u_ca_out_564[8:0],u_ca_out_563[35:9], u_ca_out_562[62:36], u_ca_out_561[71:63]};
assign col_out_565 = {u_ca_out_565[8:0],u_ca_out_564[35:9], u_ca_out_563[62:36], u_ca_out_562[71:63]};
assign col_out_566 = {u_ca_out_566[8:0],u_ca_out_565[35:9], u_ca_out_564[62:36], u_ca_out_563[71:63]};
assign col_out_567 = {u_ca_out_567[8:0],u_ca_out_566[35:9], u_ca_out_565[62:36], u_ca_out_564[71:63]};
assign col_out_568 = {u_ca_out_568[8:0],u_ca_out_567[35:9], u_ca_out_566[62:36], u_ca_out_565[71:63]};
assign col_out_569 = {u_ca_out_569[8:0],u_ca_out_568[35:9], u_ca_out_567[62:36], u_ca_out_566[71:63]};
assign col_out_570 = {u_ca_out_570[8:0],u_ca_out_569[35:9], u_ca_out_568[62:36], u_ca_out_567[71:63]};
assign col_out_571 = {u_ca_out_571[8:0],u_ca_out_570[35:9], u_ca_out_569[62:36], u_ca_out_568[71:63]};
assign col_out_572 = {u_ca_out_572[8:0],u_ca_out_571[35:9], u_ca_out_570[62:36], u_ca_out_569[71:63]};
assign col_out_573 = {u_ca_out_573[8:0],u_ca_out_572[35:9], u_ca_out_571[62:36], u_ca_out_570[71:63]};
assign col_out_574 = {u_ca_out_574[8:0],u_ca_out_573[35:9], u_ca_out_572[62:36], u_ca_out_571[71:63]};
assign col_out_575 = {u_ca_out_575[8:0],u_ca_out_574[35:9], u_ca_out_573[62:36], u_ca_out_572[71:63]};
assign col_out_576 = {u_ca_out_576[8:0],u_ca_out_575[35:9], u_ca_out_574[62:36], u_ca_out_573[71:63]};
assign col_out_577 = {u_ca_out_577[8:0],u_ca_out_576[35:9], u_ca_out_575[62:36], u_ca_out_574[71:63]};
assign col_out_578 = {u_ca_out_578[8:0],u_ca_out_577[35:9], u_ca_out_576[62:36], u_ca_out_575[71:63]};
assign col_out_579 = {u_ca_out_579[8:0],u_ca_out_578[35:9], u_ca_out_577[62:36], u_ca_out_576[71:63]};
assign col_out_580 = {u_ca_out_580[8:0],u_ca_out_579[35:9], u_ca_out_578[62:36], u_ca_out_577[71:63]};
assign col_out_581 = {u_ca_out_581[8:0],u_ca_out_580[35:9], u_ca_out_579[62:36], u_ca_out_578[71:63]};
assign col_out_582 = {u_ca_out_582[8:0],u_ca_out_581[35:9], u_ca_out_580[62:36], u_ca_out_579[71:63]};
assign col_out_583 = {u_ca_out_583[8:0],u_ca_out_582[35:9], u_ca_out_581[62:36], u_ca_out_580[71:63]};
assign col_out_584 = {u_ca_out_584[8:0],u_ca_out_583[35:9], u_ca_out_582[62:36], u_ca_out_581[71:63]};
assign col_out_585 = {u_ca_out_585[8:0],u_ca_out_584[35:9], u_ca_out_583[62:36], u_ca_out_582[71:63]};
assign col_out_586 = {u_ca_out_586[8:0],u_ca_out_585[35:9], u_ca_out_584[62:36], u_ca_out_583[71:63]};
assign col_out_587 = {u_ca_out_587[8:0],u_ca_out_586[35:9], u_ca_out_585[62:36], u_ca_out_584[71:63]};
assign col_out_588 = {u_ca_out_588[8:0],u_ca_out_587[35:9], u_ca_out_586[62:36], u_ca_out_585[71:63]};
assign col_out_589 = {u_ca_out_589[8:0],u_ca_out_588[35:9], u_ca_out_587[62:36], u_ca_out_586[71:63]};
assign col_out_590 = {u_ca_out_590[8:0],u_ca_out_589[35:9], u_ca_out_588[62:36], u_ca_out_587[71:63]};
assign col_out_591 = {u_ca_out_591[8:0],u_ca_out_590[35:9], u_ca_out_589[62:36], u_ca_out_588[71:63]};
assign col_out_592 = {u_ca_out_592[8:0],u_ca_out_591[35:9], u_ca_out_590[62:36], u_ca_out_589[71:63]};
assign col_out_593 = {u_ca_out_593[8:0],u_ca_out_592[35:9], u_ca_out_591[62:36], u_ca_out_590[71:63]};
assign col_out_594 = {u_ca_out_594[8:0],u_ca_out_593[35:9], u_ca_out_592[62:36], u_ca_out_591[71:63]};
assign col_out_595 = {u_ca_out_595[8:0],u_ca_out_594[35:9], u_ca_out_593[62:36], u_ca_out_592[71:63]};
assign col_out_596 = {u_ca_out_596[8:0],u_ca_out_595[35:9], u_ca_out_594[62:36], u_ca_out_593[71:63]};
assign col_out_597 = {u_ca_out_597[8:0],u_ca_out_596[35:9], u_ca_out_595[62:36], u_ca_out_594[71:63]};
assign col_out_598 = {u_ca_out_598[8:0],u_ca_out_597[35:9], u_ca_out_596[62:36], u_ca_out_595[71:63]};
assign col_out_599 = {u_ca_out_599[8:0],u_ca_out_598[35:9], u_ca_out_597[62:36], u_ca_out_596[71:63]};
assign col_out_600 = {u_ca_out_600[8:0],u_ca_out_599[35:9], u_ca_out_598[62:36], u_ca_out_597[71:63]};
assign col_out_601 = {u_ca_out_601[8:0],u_ca_out_600[35:9], u_ca_out_599[62:36], u_ca_out_598[71:63]};
assign col_out_602 = {u_ca_out_602[8:0],u_ca_out_601[35:9], u_ca_out_600[62:36], u_ca_out_599[71:63]};
assign col_out_603 = {u_ca_out_603[8:0],u_ca_out_602[35:9], u_ca_out_601[62:36], u_ca_out_600[71:63]};
assign col_out_604 = {u_ca_out_604[8:0],u_ca_out_603[35:9], u_ca_out_602[62:36], u_ca_out_601[71:63]};
assign col_out_605 = {u_ca_out_605[8:0],u_ca_out_604[35:9], u_ca_out_603[62:36], u_ca_out_602[71:63]};
assign col_out_606 = {u_ca_out_606[8:0],u_ca_out_605[35:9], u_ca_out_604[62:36], u_ca_out_603[71:63]};
assign col_out_607 = {u_ca_out_607[8:0],u_ca_out_606[35:9], u_ca_out_605[62:36], u_ca_out_604[71:63]};
assign col_out_608 = {u_ca_out_608[8:0],u_ca_out_607[35:9], u_ca_out_606[62:36], u_ca_out_605[71:63]};
assign col_out_609 = {u_ca_out_609[8:0],u_ca_out_608[35:9], u_ca_out_607[62:36], u_ca_out_606[71:63]};
assign col_out_610 = {u_ca_out_610[8:0],u_ca_out_609[35:9], u_ca_out_608[62:36], u_ca_out_607[71:63]};
assign col_out_611 = {u_ca_out_611[8:0],u_ca_out_610[35:9], u_ca_out_609[62:36], u_ca_out_608[71:63]};
assign col_out_612 = {u_ca_out_612[8:0],u_ca_out_611[35:9], u_ca_out_610[62:36], u_ca_out_609[71:63]};
assign col_out_613 = {u_ca_out_613[8:0],u_ca_out_612[35:9], u_ca_out_611[62:36], u_ca_out_610[71:63]};
assign col_out_614 = {u_ca_out_614[8:0],u_ca_out_613[35:9], u_ca_out_612[62:36], u_ca_out_611[71:63]};
assign col_out_615 = {u_ca_out_615[8:0],u_ca_out_614[35:9], u_ca_out_613[62:36], u_ca_out_612[71:63]};
assign col_out_616 = {u_ca_out_616[8:0],u_ca_out_615[35:9], u_ca_out_614[62:36], u_ca_out_613[71:63]};
assign col_out_617 = {u_ca_out_617[8:0],u_ca_out_616[35:9], u_ca_out_615[62:36], u_ca_out_614[71:63]};
assign col_out_618 = {u_ca_out_618[8:0],u_ca_out_617[35:9], u_ca_out_616[62:36], u_ca_out_615[71:63]};
assign col_out_619 = {u_ca_out_619[8:0],u_ca_out_618[35:9], u_ca_out_617[62:36], u_ca_out_616[71:63]};
assign col_out_620 = {u_ca_out_620[8:0],u_ca_out_619[35:9], u_ca_out_618[62:36], u_ca_out_617[71:63]};
assign col_out_621 = {u_ca_out_621[8:0],u_ca_out_620[35:9], u_ca_out_619[62:36], u_ca_out_618[71:63]};
assign col_out_622 = {u_ca_out_622[8:0],u_ca_out_621[35:9], u_ca_out_620[62:36], u_ca_out_619[71:63]};
assign col_out_623 = {u_ca_out_623[8:0],u_ca_out_622[35:9], u_ca_out_621[62:36], u_ca_out_620[71:63]};
assign col_out_624 = {u_ca_out_624[8:0],u_ca_out_623[35:9], u_ca_out_622[62:36], u_ca_out_621[71:63]};
assign col_out_625 = {u_ca_out_625[8:0],u_ca_out_624[35:9], u_ca_out_623[62:36], u_ca_out_622[71:63]};
assign col_out_626 = {u_ca_out_626[8:0],u_ca_out_625[35:9], u_ca_out_624[62:36], u_ca_out_623[71:63]};
assign col_out_627 = {u_ca_out_627[8:0],u_ca_out_626[35:9], u_ca_out_625[62:36], u_ca_out_624[71:63]};
assign col_out_628 = {u_ca_out_628[8:0],u_ca_out_627[35:9], u_ca_out_626[62:36], u_ca_out_625[71:63]};
assign col_out_629 = {u_ca_out_629[8:0],u_ca_out_628[35:9], u_ca_out_627[62:36], u_ca_out_626[71:63]};
assign col_out_630 = {u_ca_out_630[8:0],u_ca_out_629[35:9], u_ca_out_628[62:36], u_ca_out_627[71:63]};
assign col_out_631 = {u_ca_out_631[8:0],u_ca_out_630[35:9], u_ca_out_629[62:36], u_ca_out_628[71:63]};
assign col_out_632 = {u_ca_out_632[8:0],u_ca_out_631[35:9], u_ca_out_630[62:36], u_ca_out_629[71:63]};
assign col_out_633 = {u_ca_out_633[8:0],u_ca_out_632[35:9], u_ca_out_631[62:36], u_ca_out_630[71:63]};
assign col_out_634 = {u_ca_out_634[8:0],u_ca_out_633[35:9], u_ca_out_632[62:36], u_ca_out_631[71:63]};
assign col_out_635 = {u_ca_out_635[8:0],u_ca_out_634[35:9], u_ca_out_633[62:36], u_ca_out_632[71:63]};
assign col_out_636 = {u_ca_out_636[8:0],u_ca_out_635[35:9], u_ca_out_634[62:36], u_ca_out_633[71:63]};
assign col_out_637 = {u_ca_out_637[8:0],u_ca_out_636[35:9], u_ca_out_635[62:36], u_ca_out_634[71:63]};
assign col_out_638 = {u_ca_out_638[8:0],u_ca_out_637[35:9], u_ca_out_636[62:36], u_ca_out_635[71:63]};
assign col_out_639 = {u_ca_out_639[8:0],u_ca_out_638[35:9], u_ca_out_637[62:36], u_ca_out_636[71:63]};
assign col_out_640 = {u_ca_out_640[8:0],u_ca_out_639[35:9], u_ca_out_638[62:36], u_ca_out_637[71:63]};
assign col_out_641 = {u_ca_out_641[8:0],u_ca_out_640[35:9], u_ca_out_639[62:36], u_ca_out_638[71:63]};
assign col_out_642 = {u_ca_out_642[8:0],u_ca_out_641[35:9], u_ca_out_640[62:36], u_ca_out_639[71:63]};
assign col_out_643 = {u_ca_out_643[8:0],u_ca_out_642[35:9], u_ca_out_641[62:36], u_ca_out_640[71:63]};
assign col_out_644 = {u_ca_out_644[8:0],u_ca_out_643[35:9], u_ca_out_642[62:36], u_ca_out_641[71:63]};
assign col_out_645 = {u_ca_out_645[8:0],u_ca_out_644[35:9], u_ca_out_643[62:36], u_ca_out_642[71:63]};
assign col_out_646 = {u_ca_out_646[8:0],u_ca_out_645[35:9], u_ca_out_644[62:36], u_ca_out_643[71:63]};
assign col_out_647 = {u_ca_out_647[8:0],u_ca_out_646[35:9], u_ca_out_645[62:36], u_ca_out_644[71:63]};
assign col_out_648 = {u_ca_out_648[8:0],u_ca_out_647[35:9], u_ca_out_646[62:36], u_ca_out_645[71:63]};
assign col_out_649 = {u_ca_out_649[8:0],u_ca_out_648[35:9], u_ca_out_647[62:36], u_ca_out_646[71:63]};
assign col_out_650 = {u_ca_out_650[8:0],u_ca_out_649[35:9], u_ca_out_648[62:36], u_ca_out_647[71:63]};
assign col_out_651 = {u_ca_out_651[8:0],u_ca_out_650[35:9], u_ca_out_649[62:36], u_ca_out_648[71:63]};
assign col_out_652 = {u_ca_out_652[8:0],u_ca_out_651[35:9], u_ca_out_650[62:36], u_ca_out_649[71:63]};
assign col_out_653 = {u_ca_out_653[8:0],u_ca_out_652[35:9], u_ca_out_651[62:36], u_ca_out_650[71:63]};
assign col_out_654 = {u_ca_out_654[8:0],u_ca_out_653[35:9], u_ca_out_652[62:36], u_ca_out_651[71:63]};
assign col_out_655 = {u_ca_out_655[8:0],u_ca_out_654[35:9], u_ca_out_653[62:36], u_ca_out_652[71:63]};
assign col_out_656 = {u_ca_out_656[8:0],u_ca_out_655[35:9], u_ca_out_654[62:36], u_ca_out_653[71:63]};
assign col_out_657 = {u_ca_out_657[8:0],u_ca_out_656[35:9], u_ca_out_655[62:36], u_ca_out_654[71:63]};
assign col_out_658 = {u_ca_out_658[8:0],u_ca_out_657[35:9], u_ca_out_656[62:36], u_ca_out_655[71:63]};
assign col_out_659 = {u_ca_out_659[8:0],u_ca_out_658[35:9], u_ca_out_657[62:36], u_ca_out_656[71:63]};
assign col_out_660 = {u_ca_out_660[8:0],u_ca_out_659[35:9], u_ca_out_658[62:36], u_ca_out_657[71:63]};
assign col_out_661 = {u_ca_out_661[8:0],u_ca_out_660[35:9], u_ca_out_659[62:36], u_ca_out_658[71:63]};
assign col_out_662 = {u_ca_out_662[8:0],u_ca_out_661[35:9], u_ca_out_660[62:36], u_ca_out_659[71:63]};
assign col_out_663 = {u_ca_out_663[8:0],u_ca_out_662[35:9], u_ca_out_661[62:36], u_ca_out_660[71:63]};
assign col_out_664 = {u_ca_out_664[8:0],u_ca_out_663[35:9], u_ca_out_662[62:36], u_ca_out_661[71:63]};
assign col_out_665 = {u_ca_out_665[8:0],u_ca_out_664[35:9], u_ca_out_663[62:36], u_ca_out_662[71:63]};
assign col_out_666 = {u_ca_out_666[8:0],u_ca_out_665[35:9], u_ca_out_664[62:36], u_ca_out_663[71:63]};
assign col_out_667 = {u_ca_out_667[8:0],u_ca_out_666[35:9], u_ca_out_665[62:36], u_ca_out_664[71:63]};
assign col_out_668 = {u_ca_out_668[8:0],u_ca_out_667[35:9], u_ca_out_666[62:36], u_ca_out_665[71:63]};
assign col_out_669 = {u_ca_out_669[8:0],u_ca_out_668[35:9], u_ca_out_667[62:36], u_ca_out_666[71:63]};
assign col_out_670 = {u_ca_out_670[8:0],u_ca_out_669[35:9], u_ca_out_668[62:36], u_ca_out_667[71:63]};
assign col_out_671 = {u_ca_out_671[8:0],u_ca_out_670[35:9], u_ca_out_669[62:36], u_ca_out_668[71:63]};
assign col_out_672 = {u_ca_out_672[8:0],u_ca_out_671[35:9], u_ca_out_670[62:36], u_ca_out_669[71:63]};
assign col_out_673 = {u_ca_out_673[8:0],u_ca_out_672[35:9], u_ca_out_671[62:36], u_ca_out_670[71:63]};
assign col_out_674 = {u_ca_out_674[8:0],u_ca_out_673[35:9], u_ca_out_672[62:36], u_ca_out_671[71:63]};
assign col_out_675 = {u_ca_out_675[8:0],u_ca_out_674[35:9], u_ca_out_673[62:36], u_ca_out_672[71:63]};
assign col_out_676 = {u_ca_out_676[8:0],u_ca_out_675[35:9], u_ca_out_674[62:36], u_ca_out_673[71:63]};
assign col_out_677 = {u_ca_out_677[8:0],u_ca_out_676[35:9], u_ca_out_675[62:36], u_ca_out_674[71:63]};
assign col_out_678 = {u_ca_out_678[8:0],u_ca_out_677[35:9], u_ca_out_676[62:36], u_ca_out_675[71:63]};
assign col_out_679 = {u_ca_out_679[8:0],u_ca_out_678[35:9], u_ca_out_677[62:36], u_ca_out_676[71:63]};
assign col_out_680 = {u_ca_out_680[8:0],u_ca_out_679[35:9], u_ca_out_678[62:36], u_ca_out_677[71:63]};
assign col_out_681 = {u_ca_out_681[8:0],u_ca_out_680[35:9], u_ca_out_679[62:36], u_ca_out_678[71:63]};
assign col_out_682 = {u_ca_out_682[8:0],u_ca_out_681[35:9], u_ca_out_680[62:36], u_ca_out_679[71:63]};
assign col_out_683 = {u_ca_out_683[8:0],u_ca_out_682[35:9], u_ca_out_681[62:36], u_ca_out_680[71:63]};
assign col_out_684 = {u_ca_out_684[8:0],u_ca_out_683[35:9], u_ca_out_682[62:36], u_ca_out_681[71:63]};
assign col_out_685 = {u_ca_out_685[8:0],u_ca_out_684[35:9], u_ca_out_683[62:36], u_ca_out_682[71:63]};
assign col_out_686 = {u_ca_out_686[8:0],u_ca_out_685[35:9], u_ca_out_684[62:36], u_ca_out_683[71:63]};
assign col_out_687 = {u_ca_out_687[8:0],u_ca_out_686[35:9], u_ca_out_685[62:36], u_ca_out_684[71:63]};
assign col_out_688 = {u_ca_out_688[8:0],u_ca_out_687[35:9], u_ca_out_686[62:36], u_ca_out_685[71:63]};
assign col_out_689 = {u_ca_out_689[8:0],u_ca_out_688[35:9], u_ca_out_687[62:36], u_ca_out_686[71:63]};
assign col_out_690 = {u_ca_out_690[8:0],u_ca_out_689[35:9], u_ca_out_688[62:36], u_ca_out_687[71:63]};
assign col_out_691 = {u_ca_out_691[8:0],u_ca_out_690[35:9], u_ca_out_689[62:36], u_ca_out_688[71:63]};
assign col_out_692 = {u_ca_out_692[8:0],u_ca_out_691[35:9], u_ca_out_690[62:36], u_ca_out_689[71:63]};
assign col_out_693 = {u_ca_out_693[8:0],u_ca_out_692[35:9], u_ca_out_691[62:36], u_ca_out_690[71:63]};
assign col_out_694 = {u_ca_out_694[8:0],u_ca_out_693[35:9], u_ca_out_692[62:36], u_ca_out_691[71:63]};
assign col_out_695 = {u_ca_out_695[8:0],u_ca_out_694[35:9], u_ca_out_693[62:36], u_ca_out_692[71:63]};
assign col_out_696 = {u_ca_out_696[8:0],u_ca_out_695[35:9], u_ca_out_694[62:36], u_ca_out_693[71:63]};
assign col_out_697 = {u_ca_out_697[8:0],u_ca_out_696[35:9], u_ca_out_695[62:36], u_ca_out_694[71:63]};
assign col_out_698 = {u_ca_out_698[8:0],u_ca_out_697[35:9], u_ca_out_696[62:36], u_ca_out_695[71:63]};
assign col_out_699 = {u_ca_out_699[8:0],u_ca_out_698[35:9], u_ca_out_697[62:36], u_ca_out_696[71:63]};
assign col_out_700 = {u_ca_out_700[8:0],u_ca_out_699[35:9], u_ca_out_698[62:36], u_ca_out_697[71:63]};
assign col_out_701 = {u_ca_out_701[8:0],u_ca_out_700[35:9], u_ca_out_699[62:36], u_ca_out_698[71:63]};
assign col_out_702 = {u_ca_out_702[8:0],u_ca_out_701[35:9], u_ca_out_700[62:36], u_ca_out_699[71:63]};
assign col_out_703 = {u_ca_out_703[8:0],u_ca_out_702[35:9], u_ca_out_701[62:36], u_ca_out_700[71:63]};
assign col_out_704 = {u_ca_out_704[8:0],u_ca_out_703[35:9], u_ca_out_702[62:36], u_ca_out_701[71:63]};
assign col_out_705 = {u_ca_out_705[8:0],u_ca_out_704[35:9], u_ca_out_703[62:36], u_ca_out_702[71:63]};
assign col_out_706 = {u_ca_out_706[8:0],u_ca_out_705[35:9], u_ca_out_704[62:36], u_ca_out_703[71:63]};
assign col_out_707 = {u_ca_out_707[8:0],u_ca_out_706[35:9], u_ca_out_705[62:36], u_ca_out_704[71:63]};
assign col_out_708 = {u_ca_out_708[8:0],u_ca_out_707[35:9], u_ca_out_706[62:36], u_ca_out_705[71:63]};
assign col_out_709 = {u_ca_out_709[8:0],u_ca_out_708[35:9], u_ca_out_707[62:36], u_ca_out_706[71:63]};
assign col_out_710 = {u_ca_out_710[8:0],u_ca_out_709[35:9], u_ca_out_708[62:36], u_ca_out_707[71:63]};
assign col_out_711 = {u_ca_out_711[8:0],u_ca_out_710[35:9], u_ca_out_709[62:36], u_ca_out_708[71:63]};
assign col_out_712 = {u_ca_out_712[8:0],u_ca_out_711[35:9], u_ca_out_710[62:36], u_ca_out_709[71:63]};
assign col_out_713 = {u_ca_out_713[8:0],u_ca_out_712[35:9], u_ca_out_711[62:36], u_ca_out_710[71:63]};
assign col_out_714 = {u_ca_out_714[8:0],u_ca_out_713[35:9], u_ca_out_712[62:36], u_ca_out_711[71:63]};
assign col_out_715 = {u_ca_out_715[8:0],u_ca_out_714[35:9], u_ca_out_713[62:36], u_ca_out_712[71:63]};
assign col_out_716 = {u_ca_out_716[8:0],u_ca_out_715[35:9], u_ca_out_714[62:36], u_ca_out_713[71:63]};
assign col_out_717 = {u_ca_out_717[8:0],u_ca_out_716[35:9], u_ca_out_715[62:36], u_ca_out_714[71:63]};
assign col_out_718 = {u_ca_out_718[8:0],u_ca_out_717[35:9], u_ca_out_716[62:36], u_ca_out_715[71:63]};
assign col_out_719 = {u_ca_out_719[8:0],u_ca_out_718[35:9], u_ca_out_717[62:36], u_ca_out_716[71:63]};
assign col_out_720 = {u_ca_out_720[8:0],u_ca_out_719[35:9], u_ca_out_718[62:36], u_ca_out_717[71:63]};
assign col_out_721 = {u_ca_out_721[8:0],u_ca_out_720[35:9], u_ca_out_719[62:36], u_ca_out_718[71:63]};
assign col_out_722 = {u_ca_out_722[8:0],u_ca_out_721[35:9], u_ca_out_720[62:36], u_ca_out_719[71:63]};
assign col_out_723 = {u_ca_out_723[8:0],u_ca_out_722[35:9], u_ca_out_721[62:36], u_ca_out_720[71:63]};
assign col_out_724 = {u_ca_out_724[8:0],u_ca_out_723[35:9], u_ca_out_722[62:36], u_ca_out_721[71:63]};
assign col_out_725 = {u_ca_out_725[8:0],u_ca_out_724[35:9], u_ca_out_723[62:36], u_ca_out_722[71:63]};
assign col_out_726 = {u_ca_out_726[8:0],u_ca_out_725[35:9], u_ca_out_724[62:36], u_ca_out_723[71:63]};
assign col_out_727 = {u_ca_out_727[8:0],u_ca_out_726[35:9], u_ca_out_725[62:36], u_ca_out_724[71:63]};
assign col_out_728 = {u_ca_out_728[8:0],u_ca_out_727[35:9], u_ca_out_726[62:36], u_ca_out_725[71:63]};
assign col_out_729 = {u_ca_out_729[8:0],u_ca_out_728[35:9], u_ca_out_727[62:36], u_ca_out_726[71:63]};
assign col_out_730 = {u_ca_out_730[8:0],u_ca_out_729[35:9], u_ca_out_728[62:36], u_ca_out_727[71:63]};
assign col_out_731 = {u_ca_out_731[8:0],u_ca_out_730[35:9], u_ca_out_729[62:36], u_ca_out_728[71:63]};
assign col_out_732 = {u_ca_out_732[8:0],u_ca_out_731[35:9], u_ca_out_730[62:36], u_ca_out_729[71:63]};
assign col_out_733 = {u_ca_out_733[8:0],u_ca_out_732[35:9], u_ca_out_731[62:36], u_ca_out_730[71:63]};
assign col_out_734 = {u_ca_out_734[8:0],u_ca_out_733[35:9], u_ca_out_732[62:36], u_ca_out_731[71:63]};
assign col_out_735 = {u_ca_out_735[8:0],u_ca_out_734[35:9], u_ca_out_733[62:36], u_ca_out_732[71:63]};
assign col_out_736 = {u_ca_out_736[8:0],u_ca_out_735[35:9], u_ca_out_734[62:36], u_ca_out_733[71:63]};
assign col_out_737 = {u_ca_out_737[8:0],u_ca_out_736[35:9], u_ca_out_735[62:36], u_ca_out_734[71:63]};
assign col_out_738 = {u_ca_out_738[8:0],u_ca_out_737[35:9], u_ca_out_736[62:36], u_ca_out_735[71:63]};
assign col_out_739 = {u_ca_out_739[8:0],u_ca_out_738[35:9], u_ca_out_737[62:36], u_ca_out_736[71:63]};
assign col_out_740 = {u_ca_out_740[8:0],u_ca_out_739[35:9], u_ca_out_738[62:36], u_ca_out_737[71:63]};
assign col_out_741 = {u_ca_out_741[8:0],u_ca_out_740[35:9], u_ca_out_739[62:36], u_ca_out_738[71:63]};
assign col_out_742 = {u_ca_out_742[8:0],u_ca_out_741[35:9], u_ca_out_740[62:36], u_ca_out_739[71:63]};
assign col_out_743 = {u_ca_out_743[8:0],u_ca_out_742[35:9], u_ca_out_741[62:36], u_ca_out_740[71:63]};
assign col_out_744 = {u_ca_out_744[8:0],u_ca_out_743[35:9], u_ca_out_742[62:36], u_ca_out_741[71:63]};
assign col_out_745 = {u_ca_out_745[8:0],u_ca_out_744[35:9], u_ca_out_743[62:36], u_ca_out_742[71:63]};
assign col_out_746 = {u_ca_out_746[8:0],u_ca_out_745[35:9], u_ca_out_744[62:36], u_ca_out_743[71:63]};
assign col_out_747 = {u_ca_out_747[8:0],u_ca_out_746[35:9], u_ca_out_745[62:36], u_ca_out_744[71:63]};
assign col_out_748 = {u_ca_out_748[8:0],u_ca_out_747[35:9], u_ca_out_746[62:36], u_ca_out_745[71:63]};
assign col_out_749 = {u_ca_out_749[8:0],u_ca_out_748[35:9], u_ca_out_747[62:36], u_ca_out_746[71:63]};
assign col_out_750 = {u_ca_out_750[8:0],u_ca_out_749[35:9], u_ca_out_748[62:36], u_ca_out_747[71:63]};
assign col_out_751 = {u_ca_out_751[8:0],u_ca_out_750[35:9], u_ca_out_749[62:36], u_ca_out_748[71:63]};
assign col_out_752 = {u_ca_out_752[8:0],u_ca_out_751[35:9], u_ca_out_750[62:36], u_ca_out_749[71:63]};
assign col_out_753 = {u_ca_out_753[8:0],u_ca_out_752[35:9], u_ca_out_751[62:36], u_ca_out_750[71:63]};
assign col_out_754 = {u_ca_out_754[8:0],u_ca_out_753[35:9], u_ca_out_752[62:36], u_ca_out_751[71:63]};
assign col_out_755 = {u_ca_out_755[8:0],u_ca_out_754[35:9], u_ca_out_753[62:36], u_ca_out_752[71:63]};
assign col_out_756 = {u_ca_out_756[8:0],u_ca_out_755[35:9], u_ca_out_754[62:36], u_ca_out_753[71:63]};
assign col_out_757 = {u_ca_out_757[8:0],u_ca_out_756[35:9], u_ca_out_755[62:36], u_ca_out_754[71:63]};
assign col_out_758 = {u_ca_out_758[8:0],u_ca_out_757[35:9], u_ca_out_756[62:36], u_ca_out_755[71:63]};
assign col_out_759 = {u_ca_out_759[8:0],u_ca_out_758[35:9], u_ca_out_757[62:36], u_ca_out_756[71:63]};
assign col_out_760 = {u_ca_out_760[8:0],u_ca_out_759[35:9], u_ca_out_758[62:36], u_ca_out_757[71:63]};
assign col_out_761 = {u_ca_out_761[8:0],u_ca_out_760[35:9], u_ca_out_759[62:36], u_ca_out_758[71:63]};
assign col_out_762 = {u_ca_out_762[8:0],u_ca_out_761[35:9], u_ca_out_760[62:36], u_ca_out_759[71:63]};
assign col_out_763 = {u_ca_out_763[8:0],u_ca_out_762[35:9], u_ca_out_761[62:36], u_ca_out_760[71:63]};
assign col_out_764 = {u_ca_out_764[8:0],u_ca_out_763[35:9], u_ca_out_762[62:36], u_ca_out_761[71:63]};
assign col_out_765 = {u_ca_out_765[8:0],u_ca_out_764[35:9], u_ca_out_763[62:36], u_ca_out_762[71:63]};
assign col_out_766 = {u_ca_out_766[8:0],u_ca_out_765[35:9], u_ca_out_764[62:36], u_ca_out_763[71:63]};
assign col_out_767 = {u_ca_out_767[8:0],u_ca_out_766[35:9], u_ca_out_765[62:36], u_ca_out_764[71:63]};
assign col_out_768 = {u_ca_out_768[8:0],u_ca_out_767[35:9], u_ca_out_766[62:36], u_ca_out_765[71:63]};
assign col_out_769 = {u_ca_out_769[8:0],u_ca_out_768[35:9], u_ca_out_767[62:36], u_ca_out_766[71:63]};
assign col_out_770 = {u_ca_out_770[8:0],u_ca_out_769[35:9], u_ca_out_768[62:36], u_ca_out_767[71:63]};
assign col_out_771 = {u_ca_out_771[8:0],u_ca_out_770[35:9], u_ca_out_769[62:36], u_ca_out_768[71:63]};
assign col_out_772 = {u_ca_out_772[8:0],u_ca_out_771[35:9], u_ca_out_770[62:36], u_ca_out_769[71:63]};
assign col_out_773 = {u_ca_out_773[8:0],u_ca_out_772[35:9], u_ca_out_771[62:36], u_ca_out_770[71:63]};
assign col_out_774 = {u_ca_out_774[8:0],u_ca_out_773[35:9], u_ca_out_772[62:36], u_ca_out_771[71:63]};
assign col_out_775 = {u_ca_out_775[8:0],u_ca_out_774[35:9], u_ca_out_773[62:36], u_ca_out_772[71:63]};
assign col_out_776 = {u_ca_out_776[8:0],u_ca_out_775[35:9], u_ca_out_774[62:36], u_ca_out_773[71:63]};
assign col_out_777 = {u_ca_out_777[8:0],u_ca_out_776[35:9], u_ca_out_775[62:36], u_ca_out_774[71:63]};
assign col_out_778 = {u_ca_out_778[8:0],u_ca_out_777[35:9], u_ca_out_776[62:36], u_ca_out_775[71:63]};
assign col_out_779 = {u_ca_out_779[8:0],u_ca_out_778[35:9], u_ca_out_777[62:36], u_ca_out_776[71:63]};
assign col_out_780 = {u_ca_out_780[8:0],u_ca_out_779[35:9], u_ca_out_778[62:36], u_ca_out_777[71:63]};
assign col_out_781 = {u_ca_out_781[8:0],u_ca_out_780[35:9], u_ca_out_779[62:36], u_ca_out_778[71:63]};
assign col_out_782 = {u_ca_out_782[8:0],u_ca_out_781[35:9], u_ca_out_780[62:36], u_ca_out_779[71:63]};
assign col_out_783 = {u_ca_out_783[8:0],u_ca_out_782[35:9], u_ca_out_781[62:36], u_ca_out_780[71:63]};
assign col_out_784 = {u_ca_out_784[8:0],u_ca_out_783[35:9], u_ca_out_782[62:36], u_ca_out_781[71:63]};
assign col_out_785 = {u_ca_out_785[8:0],u_ca_out_784[35:9], u_ca_out_783[62:36], u_ca_out_782[71:63]};
assign col_out_786 = {u_ca_out_786[8:0],u_ca_out_785[35:9], u_ca_out_784[62:36], u_ca_out_783[71:63]};
assign col_out_787 = {u_ca_out_787[8:0],u_ca_out_786[35:9], u_ca_out_785[62:36], u_ca_out_784[71:63]};
assign col_out_788 = {u_ca_out_788[8:0],u_ca_out_787[35:9], u_ca_out_786[62:36], u_ca_out_785[71:63]};
assign col_out_789 = {u_ca_out_789[8:0],u_ca_out_788[35:9], u_ca_out_787[62:36], u_ca_out_786[71:63]};
assign col_out_790 = {u_ca_out_790[8:0],u_ca_out_789[35:9], u_ca_out_788[62:36], u_ca_out_787[71:63]};
assign col_out_791 = {u_ca_out_791[8:0],u_ca_out_790[35:9], u_ca_out_789[62:36], u_ca_out_788[71:63]};
assign col_out_792 = {u_ca_out_792[8:0],u_ca_out_791[35:9], u_ca_out_790[62:36], u_ca_out_789[71:63]};
assign col_out_793 = {u_ca_out_793[8:0],u_ca_out_792[35:9], u_ca_out_791[62:36], u_ca_out_790[71:63]};
assign col_out_794 = {u_ca_out_794[8:0],u_ca_out_793[35:9], u_ca_out_792[62:36], u_ca_out_791[71:63]};
assign col_out_795 = {u_ca_out_795[8:0],u_ca_out_794[35:9], u_ca_out_793[62:36], u_ca_out_792[71:63]};
assign col_out_796 = {u_ca_out_796[8:0],u_ca_out_795[35:9], u_ca_out_794[62:36], u_ca_out_793[71:63]};
assign col_out_797 = {u_ca_out_797[8:0],u_ca_out_796[35:9], u_ca_out_795[62:36], u_ca_out_794[71:63]};
assign col_out_798 = {u_ca_out_798[8:0],u_ca_out_797[35:9], u_ca_out_796[62:36], u_ca_out_795[71:63]};
assign col_out_799 = {u_ca_out_799[8:0],u_ca_out_798[35:9], u_ca_out_797[62:36], u_ca_out_796[71:63]};
assign col_out_800 = {u_ca_out_800[8:0],u_ca_out_799[35:9], u_ca_out_798[62:36], u_ca_out_797[71:63]};
assign col_out_801 = {u_ca_out_801[8:0],u_ca_out_800[35:9], u_ca_out_799[62:36], u_ca_out_798[71:63]};
assign col_out_802 = {u_ca_out_802[8:0],u_ca_out_801[35:9], u_ca_out_800[62:36], u_ca_out_799[71:63]};
assign col_out_803 = {u_ca_out_803[8:0],u_ca_out_802[35:9], u_ca_out_801[62:36], u_ca_out_800[71:63]};
assign col_out_804 = {u_ca_out_804[8:0],u_ca_out_803[35:9], u_ca_out_802[62:36], u_ca_out_801[71:63]};
assign col_out_805 = {u_ca_out_805[8:0],u_ca_out_804[35:9], u_ca_out_803[62:36], u_ca_out_802[71:63]};
assign col_out_806 = {u_ca_out_806[8:0],u_ca_out_805[35:9], u_ca_out_804[62:36], u_ca_out_803[71:63]};
assign col_out_807 = {u_ca_out_807[8:0],u_ca_out_806[35:9], u_ca_out_805[62:36], u_ca_out_804[71:63]};
assign col_out_808 = {u_ca_out_808[8:0],u_ca_out_807[35:9], u_ca_out_806[62:36], u_ca_out_805[71:63]};
assign col_out_809 = {u_ca_out_809[8:0],u_ca_out_808[35:9], u_ca_out_807[62:36], u_ca_out_806[71:63]};
assign col_out_810 = {u_ca_out_810[8:0],u_ca_out_809[35:9], u_ca_out_808[62:36], u_ca_out_807[71:63]};
assign col_out_811 = {u_ca_out_811[8:0],u_ca_out_810[35:9], u_ca_out_809[62:36], u_ca_out_808[71:63]};
assign col_out_812 = {u_ca_out_812[8:0],u_ca_out_811[35:9], u_ca_out_810[62:36], u_ca_out_809[71:63]};
assign col_out_813 = {u_ca_out_813[8:0],u_ca_out_812[35:9], u_ca_out_811[62:36], u_ca_out_810[71:63]};
assign col_out_814 = {u_ca_out_814[8:0],u_ca_out_813[35:9], u_ca_out_812[62:36], u_ca_out_811[71:63]};
assign col_out_815 = {u_ca_out_815[8:0],u_ca_out_814[35:9], u_ca_out_813[62:36], u_ca_out_812[71:63]};
assign col_out_816 = {u_ca_out_816[8:0],u_ca_out_815[35:9], u_ca_out_814[62:36], u_ca_out_813[71:63]};
assign col_out_817 = {u_ca_out_817[8:0],u_ca_out_816[35:9], u_ca_out_815[62:36], u_ca_out_814[71:63]};
assign col_out_818 = {u_ca_out_818[8:0],u_ca_out_817[35:9], u_ca_out_816[62:36], u_ca_out_815[71:63]};
assign col_out_819 = {u_ca_out_819[8:0],u_ca_out_818[35:9], u_ca_out_817[62:36], u_ca_out_816[71:63]};
assign col_out_820 = {u_ca_out_820[8:0],u_ca_out_819[35:9], u_ca_out_818[62:36], u_ca_out_817[71:63]};
assign col_out_821 = {u_ca_out_821[8:0],u_ca_out_820[35:9], u_ca_out_819[62:36], u_ca_out_818[71:63]};
assign col_out_822 = {u_ca_out_822[8:0],u_ca_out_821[35:9], u_ca_out_820[62:36], u_ca_out_819[71:63]};
assign col_out_823 = {u_ca_out_823[8:0],u_ca_out_822[35:9], u_ca_out_821[62:36], u_ca_out_820[71:63]};
assign col_out_824 = {u_ca_out_824[8:0],u_ca_out_823[35:9], u_ca_out_822[62:36], u_ca_out_821[71:63]};
assign col_out_825 = {u_ca_out_825[8:0],u_ca_out_824[35:9], u_ca_out_823[62:36], u_ca_out_822[71:63]};
assign col_out_826 = {u_ca_out_826[8:0],u_ca_out_825[35:9], u_ca_out_824[62:36], u_ca_out_823[71:63]};
assign col_out_827 = {u_ca_out_827[8:0],u_ca_out_826[35:9], u_ca_out_825[62:36], u_ca_out_824[71:63]};
assign col_out_828 = {u_ca_out_828[8:0],u_ca_out_827[35:9], u_ca_out_826[62:36], u_ca_out_825[71:63]};
assign col_out_829 = {u_ca_out_829[8:0],u_ca_out_828[35:9], u_ca_out_827[62:36], u_ca_out_826[71:63]};
assign col_out_830 = {u_ca_out_830[8:0],u_ca_out_829[35:9], u_ca_out_828[62:36], u_ca_out_827[71:63]};
assign col_out_831 = {u_ca_out_831[8:0],u_ca_out_830[35:9], u_ca_out_829[62:36], u_ca_out_828[71:63]};
assign col_out_832 = {u_ca_out_832[8:0],u_ca_out_831[35:9], u_ca_out_830[62:36], u_ca_out_829[71:63]};
assign col_out_833 = {u_ca_out_833[8:0],u_ca_out_832[35:9], u_ca_out_831[62:36], u_ca_out_830[71:63]};
assign col_out_834 = {u_ca_out_834[8:0],u_ca_out_833[35:9], u_ca_out_832[62:36], u_ca_out_831[71:63]};
assign col_out_835 = {u_ca_out_835[8:0],u_ca_out_834[35:9], u_ca_out_833[62:36], u_ca_out_832[71:63]};
assign col_out_836 = {u_ca_out_836[8:0],u_ca_out_835[35:9], u_ca_out_834[62:36], u_ca_out_833[71:63]};
assign col_out_837 = {u_ca_out_837[8:0],u_ca_out_836[35:9], u_ca_out_835[62:36], u_ca_out_834[71:63]};
assign col_out_838 = {u_ca_out_838[8:0],u_ca_out_837[35:9], u_ca_out_836[62:36], u_ca_out_835[71:63]};
assign col_out_839 = {u_ca_out_839[8:0],u_ca_out_838[35:9], u_ca_out_837[62:36], u_ca_out_836[71:63]};
assign col_out_840 = {u_ca_out_840[8:0],u_ca_out_839[35:9], u_ca_out_838[62:36], u_ca_out_837[71:63]};
assign col_out_841 = {u_ca_out_841[8:0],u_ca_out_840[35:9], u_ca_out_839[62:36], u_ca_out_838[71:63]};
assign col_out_842 = {u_ca_out_842[8:0],u_ca_out_841[35:9], u_ca_out_840[62:36], u_ca_out_839[71:63]};
assign col_out_843 = {u_ca_out_843[8:0],u_ca_out_842[35:9], u_ca_out_841[62:36], u_ca_out_840[71:63]};
assign col_out_844 = {u_ca_out_844[8:0],u_ca_out_843[35:9], u_ca_out_842[62:36], u_ca_out_841[71:63]};
assign col_out_845 = {u_ca_out_845[8:0],u_ca_out_844[35:9], u_ca_out_843[62:36], u_ca_out_842[71:63]};
assign col_out_846 = {u_ca_out_846[8:0],u_ca_out_845[35:9], u_ca_out_844[62:36], u_ca_out_843[71:63]};
assign col_out_847 = {u_ca_out_847[8:0],u_ca_out_846[35:9], u_ca_out_845[62:36], u_ca_out_844[71:63]};
assign col_out_848 = {u_ca_out_848[8:0],u_ca_out_847[35:9], u_ca_out_846[62:36], u_ca_out_845[71:63]};
assign col_out_849 = {u_ca_out_849[8:0],u_ca_out_848[35:9], u_ca_out_847[62:36], u_ca_out_846[71:63]};
assign col_out_850 = {u_ca_out_850[8:0],u_ca_out_849[35:9], u_ca_out_848[62:36], u_ca_out_847[71:63]};
assign col_out_851 = {u_ca_out_851[8:0],u_ca_out_850[35:9], u_ca_out_849[62:36], u_ca_out_848[71:63]};
assign col_out_852 = {u_ca_out_852[8:0],u_ca_out_851[35:9], u_ca_out_850[62:36], u_ca_out_849[71:63]};
assign col_out_853 = {u_ca_out_853[8:0],u_ca_out_852[35:9], u_ca_out_851[62:36], u_ca_out_850[71:63]};
assign col_out_854 = {u_ca_out_854[8:0],u_ca_out_853[35:9], u_ca_out_852[62:36], u_ca_out_851[71:63]};
assign col_out_855 = {u_ca_out_855[8:0],u_ca_out_854[35:9], u_ca_out_853[62:36], u_ca_out_852[71:63]};
assign col_out_856 = {u_ca_out_856[8:0],u_ca_out_855[35:9], u_ca_out_854[62:36], u_ca_out_853[71:63]};
assign col_out_857 = {u_ca_out_857[8:0],u_ca_out_856[35:9], u_ca_out_855[62:36], u_ca_out_854[71:63]};
assign col_out_858 = {u_ca_out_858[8:0],u_ca_out_857[35:9], u_ca_out_856[62:36], u_ca_out_855[71:63]};
assign col_out_859 = {u_ca_out_859[8:0],u_ca_out_858[35:9], u_ca_out_857[62:36], u_ca_out_856[71:63]};
assign col_out_860 = {u_ca_out_860[8:0],u_ca_out_859[35:9], u_ca_out_858[62:36], u_ca_out_857[71:63]};
assign col_out_861 = {u_ca_out_861[8:0],u_ca_out_860[35:9], u_ca_out_859[62:36], u_ca_out_858[71:63]};
assign col_out_862 = {u_ca_out_862[8:0],u_ca_out_861[35:9], u_ca_out_860[62:36], u_ca_out_859[71:63]};
assign col_out_863 = {u_ca_out_863[8:0],u_ca_out_862[35:9], u_ca_out_861[62:36], u_ca_out_860[71:63]};
assign col_out_864 = {u_ca_out_864[8:0],u_ca_out_863[35:9], u_ca_out_862[62:36], u_ca_out_861[71:63]};
assign col_out_865 = {u_ca_out_865[8:0],u_ca_out_864[35:9], u_ca_out_863[62:36], u_ca_out_862[71:63]};
assign col_out_866 = {u_ca_out_866[8:0],u_ca_out_865[35:9], u_ca_out_864[62:36], u_ca_out_863[71:63]};
assign col_out_867 = {u_ca_out_867[8:0],u_ca_out_866[35:9], u_ca_out_865[62:36], u_ca_out_864[71:63]};
assign col_out_868 = {u_ca_out_868[8:0],u_ca_out_867[35:9], u_ca_out_866[62:36], u_ca_out_865[71:63]};
assign col_out_869 = {u_ca_out_869[8:0],u_ca_out_868[35:9], u_ca_out_867[62:36], u_ca_out_866[71:63]};
assign col_out_870 = {u_ca_out_870[8:0],u_ca_out_869[35:9], u_ca_out_868[62:36], u_ca_out_867[71:63]};
assign col_out_871 = {u_ca_out_871[8:0],u_ca_out_870[35:9], u_ca_out_869[62:36], u_ca_out_868[71:63]};
assign col_out_872 = {u_ca_out_872[8:0],u_ca_out_871[35:9], u_ca_out_870[62:36], u_ca_out_869[71:63]};
assign col_out_873 = {u_ca_out_873[8:0],u_ca_out_872[35:9], u_ca_out_871[62:36], u_ca_out_870[71:63]};
assign col_out_874 = {u_ca_out_874[8:0],u_ca_out_873[35:9], u_ca_out_872[62:36], u_ca_out_871[71:63]};
assign col_out_875 = {u_ca_out_875[8:0],u_ca_out_874[35:9], u_ca_out_873[62:36], u_ca_out_872[71:63]};
assign col_out_876 = {u_ca_out_876[8:0],u_ca_out_875[35:9], u_ca_out_874[62:36], u_ca_out_873[71:63]};
assign col_out_877 = {u_ca_out_877[8:0],u_ca_out_876[35:9], u_ca_out_875[62:36], u_ca_out_874[71:63]};
assign col_out_878 = {u_ca_out_878[8:0],u_ca_out_877[35:9], u_ca_out_876[62:36], u_ca_out_875[71:63]};
assign col_out_879 = {u_ca_out_879[8:0],u_ca_out_878[35:9], u_ca_out_877[62:36], u_ca_out_876[71:63]};
assign col_out_880 = {u_ca_out_880[8:0],u_ca_out_879[35:9], u_ca_out_878[62:36], u_ca_out_877[71:63]};
assign col_out_881 = {u_ca_out_881[8:0],u_ca_out_880[35:9], u_ca_out_879[62:36], u_ca_out_878[71:63]};
assign col_out_882 = {u_ca_out_882[8:0],u_ca_out_881[35:9], u_ca_out_880[62:36], u_ca_out_879[71:63]};
assign col_out_883 = {u_ca_out_883[8:0],u_ca_out_882[35:9], u_ca_out_881[62:36], u_ca_out_880[71:63]};
assign col_out_884 = {u_ca_out_884[8:0],u_ca_out_883[35:9], u_ca_out_882[62:36], u_ca_out_881[71:63]};
assign col_out_885 = {u_ca_out_885[8:0],u_ca_out_884[35:9], u_ca_out_883[62:36], u_ca_out_882[71:63]};
assign col_out_886 = {u_ca_out_886[8:0],u_ca_out_885[35:9], u_ca_out_884[62:36], u_ca_out_883[71:63]};
assign col_out_887 = {u_ca_out_887[8:0],u_ca_out_886[35:9], u_ca_out_885[62:36], u_ca_out_884[71:63]};
assign col_out_888 = {u_ca_out_888[8:0],u_ca_out_887[35:9], u_ca_out_886[62:36], u_ca_out_885[71:63]};
assign col_out_889 = {u_ca_out_889[8:0],u_ca_out_888[35:9], u_ca_out_887[62:36], u_ca_out_886[71:63]};
assign col_out_890 = {u_ca_out_890[8:0],u_ca_out_889[35:9], u_ca_out_888[62:36], u_ca_out_887[71:63]};
assign col_out_891 = {u_ca_out_891[8:0],u_ca_out_890[35:9], u_ca_out_889[62:36], u_ca_out_888[71:63]};
assign col_out_892 = {u_ca_out_892[8:0],u_ca_out_891[35:9], u_ca_out_890[62:36], u_ca_out_889[71:63]};
assign col_out_893 = {u_ca_out_893[8:0],u_ca_out_892[35:9], u_ca_out_891[62:36], u_ca_out_890[71:63]};
assign col_out_894 = {u_ca_out_894[8:0],u_ca_out_893[35:9], u_ca_out_892[62:36], u_ca_out_891[71:63]};
assign col_out_895 = {u_ca_out_895[8:0],u_ca_out_894[35:9], u_ca_out_893[62:36], u_ca_out_892[71:63]};
assign col_out_896 = {u_ca_out_896[8:0],u_ca_out_895[35:9], u_ca_out_894[62:36], u_ca_out_893[71:63]};
assign col_out_897 = {u_ca_out_897[8:0],u_ca_out_896[35:9], u_ca_out_895[62:36], u_ca_out_894[71:63]};
assign col_out_898 = {u_ca_out_898[8:0],u_ca_out_897[35:9], u_ca_out_896[62:36], u_ca_out_895[71:63]};
assign col_out_899 = {u_ca_out_899[8:0],u_ca_out_898[35:9], u_ca_out_897[62:36], u_ca_out_896[71:63]};
assign col_out_900 = {u_ca_out_900[8:0],u_ca_out_899[35:9], u_ca_out_898[62:36], u_ca_out_897[71:63]};
assign col_out_901 = {u_ca_out_901[8:0],u_ca_out_900[35:9], u_ca_out_899[62:36], u_ca_out_898[71:63]};
assign col_out_902 = {u_ca_out_902[8:0],u_ca_out_901[35:9], u_ca_out_900[62:36], u_ca_out_899[71:63]};
assign col_out_903 = {u_ca_out_903[8:0],u_ca_out_902[35:9], u_ca_out_901[62:36], u_ca_out_900[71:63]};
assign col_out_904 = {u_ca_out_904[8:0],u_ca_out_903[35:9], u_ca_out_902[62:36], u_ca_out_901[71:63]};
assign col_out_905 = {u_ca_out_905[8:0],u_ca_out_904[35:9], u_ca_out_903[62:36], u_ca_out_902[71:63]};
assign col_out_906 = {u_ca_out_906[8:0],u_ca_out_905[35:9], u_ca_out_904[62:36], u_ca_out_903[71:63]};
assign col_out_907 = {u_ca_out_907[8:0],u_ca_out_906[35:9], u_ca_out_905[62:36], u_ca_out_904[71:63]};
assign col_out_908 = {u_ca_out_908[8:0],u_ca_out_907[35:9], u_ca_out_906[62:36], u_ca_out_905[71:63]};
assign col_out_909 = {u_ca_out_909[8:0],u_ca_out_908[35:9], u_ca_out_907[62:36], u_ca_out_906[71:63]};
assign col_out_910 = {u_ca_out_910[8:0],u_ca_out_909[35:9], u_ca_out_908[62:36], u_ca_out_907[71:63]};
assign col_out_911 = {u_ca_out_911[8:0],u_ca_out_910[35:9], u_ca_out_909[62:36], u_ca_out_908[71:63]};
assign col_out_912 = {u_ca_out_912[8:0],u_ca_out_911[35:9], u_ca_out_910[62:36], u_ca_out_909[71:63]};
assign col_out_913 = {u_ca_out_913[8:0],u_ca_out_912[35:9], u_ca_out_911[62:36], u_ca_out_910[71:63]};
assign col_out_914 = {u_ca_out_914[8:0],u_ca_out_913[35:9], u_ca_out_912[62:36], u_ca_out_911[71:63]};
assign col_out_915 = {u_ca_out_915[8:0],u_ca_out_914[35:9], u_ca_out_913[62:36], u_ca_out_912[71:63]};
assign col_out_916 = {u_ca_out_916[8:0],u_ca_out_915[35:9], u_ca_out_914[62:36], u_ca_out_913[71:63]};
assign col_out_917 = {u_ca_out_917[8:0],u_ca_out_916[35:9], u_ca_out_915[62:36], u_ca_out_914[71:63]};
assign col_out_918 = {u_ca_out_918[8:0],u_ca_out_917[35:9], u_ca_out_916[62:36], u_ca_out_915[71:63]};
assign col_out_919 = {u_ca_out_919[8:0],u_ca_out_918[35:9], u_ca_out_917[62:36], u_ca_out_916[71:63]};
assign col_out_920 = {u_ca_out_920[8:0],u_ca_out_919[35:9], u_ca_out_918[62:36], u_ca_out_917[71:63]};
assign col_out_921 = {u_ca_out_921[8:0],u_ca_out_920[35:9], u_ca_out_919[62:36], u_ca_out_918[71:63]};
assign col_out_922 = {u_ca_out_922[8:0],u_ca_out_921[35:9], u_ca_out_920[62:36], u_ca_out_919[71:63]};
assign col_out_923 = {u_ca_out_923[8:0],u_ca_out_922[35:9], u_ca_out_921[62:36], u_ca_out_920[71:63]};
assign col_out_924 = {u_ca_out_924[8:0],u_ca_out_923[35:9], u_ca_out_922[62:36], u_ca_out_921[71:63]};
assign col_out_925 = {u_ca_out_925[8:0],u_ca_out_924[35:9], u_ca_out_923[62:36], u_ca_out_922[71:63]};
assign col_out_926 = {u_ca_out_926[8:0],u_ca_out_925[35:9], u_ca_out_924[62:36], u_ca_out_923[71:63]};
assign col_out_927 = {u_ca_out_927[8:0],u_ca_out_926[35:9], u_ca_out_925[62:36], u_ca_out_924[71:63]};
assign col_out_928 = {u_ca_out_928[8:0],u_ca_out_927[35:9], u_ca_out_926[62:36], u_ca_out_925[71:63]};
assign col_out_929 = {u_ca_out_929[8:0],u_ca_out_928[35:9], u_ca_out_927[62:36], u_ca_out_926[71:63]};
assign col_out_930 = {u_ca_out_930[8:0],u_ca_out_929[35:9], u_ca_out_928[62:36], u_ca_out_927[71:63]};
assign col_out_931 = {u_ca_out_931[8:0],u_ca_out_930[35:9], u_ca_out_929[62:36], u_ca_out_928[71:63]};
assign col_out_932 = {u_ca_out_932[8:0],u_ca_out_931[35:9], u_ca_out_930[62:36], u_ca_out_929[71:63]};
assign col_out_933 = {u_ca_out_933[8:0],u_ca_out_932[35:9], u_ca_out_931[62:36], u_ca_out_930[71:63]};
assign col_out_934 = {u_ca_out_934[8:0],u_ca_out_933[35:9], u_ca_out_932[62:36], u_ca_out_931[71:63]};
assign col_out_935 = {u_ca_out_935[8:0],u_ca_out_934[35:9], u_ca_out_933[62:36], u_ca_out_932[71:63]};
assign col_out_936 = {u_ca_out_936[8:0],u_ca_out_935[35:9], u_ca_out_934[62:36], u_ca_out_933[71:63]};
assign col_out_937 = {u_ca_out_937[8:0],u_ca_out_936[35:9], u_ca_out_935[62:36], u_ca_out_934[71:63]};
assign col_out_938 = {u_ca_out_938[8:0],u_ca_out_937[35:9], u_ca_out_936[62:36], u_ca_out_935[71:63]};
assign col_out_939 = {u_ca_out_939[8:0],u_ca_out_938[35:9], u_ca_out_937[62:36], u_ca_out_936[71:63]};
assign col_out_940 = {u_ca_out_940[8:0],u_ca_out_939[35:9], u_ca_out_938[62:36], u_ca_out_937[71:63]};
assign col_out_941 = {u_ca_out_941[8:0],u_ca_out_940[35:9], u_ca_out_939[62:36], u_ca_out_938[71:63]};
assign col_out_942 = {u_ca_out_942[8:0],u_ca_out_941[35:9], u_ca_out_940[62:36], u_ca_out_939[71:63]};
assign col_out_943 = {u_ca_out_943[8:0],u_ca_out_942[35:9], u_ca_out_941[62:36], u_ca_out_940[71:63]};
assign col_out_944 = {u_ca_out_944[8:0],u_ca_out_943[35:9], u_ca_out_942[62:36], u_ca_out_941[71:63]};
assign col_out_945 = {u_ca_out_945[8:0],u_ca_out_944[35:9], u_ca_out_943[62:36], u_ca_out_942[71:63]};
assign col_out_946 = {u_ca_out_946[8:0],u_ca_out_945[35:9], u_ca_out_944[62:36], u_ca_out_943[71:63]};
assign col_out_947 = {u_ca_out_947[8:0],u_ca_out_946[35:9], u_ca_out_945[62:36], u_ca_out_944[71:63]};
assign col_out_948 = {u_ca_out_948[8:0],u_ca_out_947[35:9], u_ca_out_946[62:36], u_ca_out_945[71:63]};
assign col_out_949 = {u_ca_out_949[8:0],u_ca_out_948[35:9], u_ca_out_947[62:36], u_ca_out_946[71:63]};
assign col_out_950 = {u_ca_out_950[8:0],u_ca_out_949[35:9], u_ca_out_948[62:36], u_ca_out_947[71:63]};
assign col_out_951 = {u_ca_out_951[8:0],u_ca_out_950[35:9], u_ca_out_949[62:36], u_ca_out_948[71:63]};
assign col_out_952 = {u_ca_out_952[8:0],u_ca_out_951[35:9], u_ca_out_950[62:36], u_ca_out_949[71:63]};
assign col_out_953 = {u_ca_out_953[8:0],u_ca_out_952[35:9], u_ca_out_951[62:36], u_ca_out_950[71:63]};
assign col_out_954 = {u_ca_out_954[8:0],u_ca_out_953[35:9], u_ca_out_952[62:36], u_ca_out_951[71:63]};
assign col_out_955 = {u_ca_out_955[8:0],u_ca_out_954[35:9], u_ca_out_953[62:36], u_ca_out_952[71:63]};
assign col_out_956 = {u_ca_out_956[8:0],u_ca_out_955[35:9], u_ca_out_954[62:36], u_ca_out_953[71:63]};
assign col_out_957 = {u_ca_out_957[8:0],u_ca_out_956[35:9], u_ca_out_955[62:36], u_ca_out_954[71:63]};
assign col_out_958 = {u_ca_out_958[8:0],u_ca_out_957[35:9], u_ca_out_956[62:36], u_ca_out_955[71:63]};
assign col_out_959 = {u_ca_out_959[8:0],u_ca_out_958[35:9], u_ca_out_957[62:36], u_ca_out_956[71:63]};
assign col_out_960 = {u_ca_out_960[8:0],u_ca_out_959[35:9], u_ca_out_958[62:36], u_ca_out_957[71:63]};
assign col_out_961 = {u_ca_out_961[8:0],u_ca_out_960[35:9], u_ca_out_959[62:36], u_ca_out_958[71:63]};
assign col_out_962 = {u_ca_out_962[8:0],u_ca_out_961[35:9], u_ca_out_960[62:36], u_ca_out_959[71:63]};
assign col_out_963 = {u_ca_out_963[8:0],u_ca_out_962[35:9], u_ca_out_961[62:36], u_ca_out_960[71:63]};
assign col_out_964 = {u_ca_out_964[8:0],u_ca_out_963[35:9], u_ca_out_962[62:36], u_ca_out_961[71:63]};
assign col_out_965 = {u_ca_out_965[8:0],u_ca_out_964[35:9], u_ca_out_963[62:36], u_ca_out_962[71:63]};
assign col_out_966 = {u_ca_out_966[8:0],u_ca_out_965[35:9], u_ca_out_964[62:36], u_ca_out_963[71:63]};
assign col_out_967 = {u_ca_out_967[8:0],u_ca_out_966[35:9], u_ca_out_965[62:36], u_ca_out_964[71:63]};
assign col_out_968 = {u_ca_out_968[8:0],u_ca_out_967[35:9], u_ca_out_966[62:36], u_ca_out_965[71:63]};
assign col_out_969 = {u_ca_out_969[8:0],u_ca_out_968[35:9], u_ca_out_967[62:36], u_ca_out_966[71:63]};
assign col_out_970 = {u_ca_out_970[8:0],u_ca_out_969[35:9], u_ca_out_968[62:36], u_ca_out_967[71:63]};
assign col_out_971 = {u_ca_out_971[8:0],u_ca_out_970[35:9], u_ca_out_969[62:36], u_ca_out_968[71:63]};
assign col_out_972 = {u_ca_out_972[8:0],u_ca_out_971[35:9], u_ca_out_970[62:36], u_ca_out_969[71:63]};
assign col_out_973 = {u_ca_out_973[8:0],u_ca_out_972[35:9], u_ca_out_971[62:36], u_ca_out_970[71:63]};
assign col_out_974 = {u_ca_out_974[8:0],u_ca_out_973[35:9], u_ca_out_972[62:36], u_ca_out_971[71:63]};
assign col_out_975 = {u_ca_out_975[8:0],u_ca_out_974[35:9], u_ca_out_973[62:36], u_ca_out_972[71:63]};
assign col_out_976 = {u_ca_out_976[8:0],u_ca_out_975[35:9], u_ca_out_974[62:36], u_ca_out_973[71:63]};
assign col_out_977 = {u_ca_out_977[8:0],u_ca_out_976[35:9], u_ca_out_975[62:36], u_ca_out_974[71:63]};
assign col_out_978 = {u_ca_out_978[8:0],u_ca_out_977[35:9], u_ca_out_976[62:36], u_ca_out_975[71:63]};
assign col_out_979 = {u_ca_out_979[8:0],u_ca_out_978[35:9], u_ca_out_977[62:36], u_ca_out_976[71:63]};
assign col_out_980 = {u_ca_out_980[8:0],u_ca_out_979[35:9], u_ca_out_978[62:36], u_ca_out_977[71:63]};
assign col_out_981 = {u_ca_out_981[8:0],u_ca_out_980[35:9], u_ca_out_979[62:36], u_ca_out_978[71:63]};
assign col_out_982 = {u_ca_out_982[8:0],u_ca_out_981[35:9], u_ca_out_980[62:36], u_ca_out_979[71:63]};
assign col_out_983 = {u_ca_out_983[8:0],u_ca_out_982[35:9], u_ca_out_981[62:36], u_ca_out_980[71:63]};
assign col_out_984 = {u_ca_out_984[8:0],u_ca_out_983[35:9], u_ca_out_982[62:36], u_ca_out_981[71:63]};
assign col_out_985 = {u_ca_out_985[8:0],u_ca_out_984[35:9], u_ca_out_983[62:36], u_ca_out_982[71:63]};
assign col_out_986 = {u_ca_out_986[8:0],u_ca_out_985[35:9], u_ca_out_984[62:36], u_ca_out_983[71:63]};
assign col_out_987 = {u_ca_out_987[8:0],u_ca_out_986[35:9], u_ca_out_985[62:36], u_ca_out_984[71:63]};
assign col_out_988 = {u_ca_out_988[8:0],u_ca_out_987[35:9], u_ca_out_986[62:36], u_ca_out_985[71:63]};
assign col_out_989 = {u_ca_out_989[8:0],u_ca_out_988[35:9], u_ca_out_987[62:36], u_ca_out_986[71:63]};
assign col_out_990 = {u_ca_out_990[8:0],u_ca_out_989[35:9], u_ca_out_988[62:36], u_ca_out_987[71:63]};
assign col_out_991 = {u_ca_out_991[8:0],u_ca_out_990[35:9], u_ca_out_989[62:36], u_ca_out_988[71:63]};
assign col_out_992 = {u_ca_out_992[8:0],u_ca_out_991[35:9], u_ca_out_990[62:36], u_ca_out_989[71:63]};
assign col_out_993 = {u_ca_out_993[8:0],u_ca_out_992[35:9], u_ca_out_991[62:36], u_ca_out_990[71:63]};
assign col_out_994 = {u_ca_out_994[8:0],u_ca_out_993[35:9], u_ca_out_992[62:36], u_ca_out_991[71:63]};
assign col_out_995 = {u_ca_out_995[8:0],u_ca_out_994[35:9], u_ca_out_993[62:36], u_ca_out_992[71:63]};
assign col_out_996 = {u_ca_out_996[8:0],u_ca_out_995[35:9], u_ca_out_994[62:36], u_ca_out_993[71:63]};
assign col_out_997 = {u_ca_out_997[8:0],u_ca_out_996[35:9], u_ca_out_995[62:36], u_ca_out_994[71:63]};
assign col_out_998 = {u_ca_out_998[8:0],u_ca_out_997[35:9], u_ca_out_996[62:36], u_ca_out_995[71:63]};
assign col_out_999 = {u_ca_out_999[8:0],u_ca_out_998[35:9], u_ca_out_997[62:36], u_ca_out_996[71:63]};
assign col_out_1000 = {u_ca_out_1000[8:0],u_ca_out_999[35:9], u_ca_out_998[62:36], u_ca_out_997[71:63]};
assign col_out_1001 = {u_ca_out_1001[8:0],u_ca_out_1000[35:9], u_ca_out_999[62:36], u_ca_out_998[71:63]};
assign col_out_1002 = {u_ca_out_1002[8:0],u_ca_out_1001[35:9], u_ca_out_1000[62:36], u_ca_out_999[71:63]};
assign col_out_1003 = {u_ca_out_1003[8:0],u_ca_out_1002[35:9], u_ca_out_1001[62:36], u_ca_out_1000[71:63]};
assign col_out_1004 = {u_ca_out_1004[8:0],u_ca_out_1003[35:9], u_ca_out_1002[62:36], u_ca_out_1001[71:63]};
assign col_out_1005 = {u_ca_out_1005[8:0],u_ca_out_1004[35:9], u_ca_out_1003[62:36], u_ca_out_1002[71:63]};
assign col_out_1006 = {u_ca_out_1006[8:0],u_ca_out_1005[35:9], u_ca_out_1004[62:36], u_ca_out_1003[71:63]};
assign col_out_1007 = {u_ca_out_1007[8:0],u_ca_out_1006[35:9], u_ca_out_1005[62:36], u_ca_out_1004[71:63]};
assign col_out_1008 = {u_ca_out_1008[8:0],u_ca_out_1007[35:9], u_ca_out_1006[62:36], u_ca_out_1005[71:63]};
assign col_out_1009 = {u_ca_out_1009[8:0],u_ca_out_1008[35:9], u_ca_out_1007[62:36], u_ca_out_1006[71:63]};
assign col_out_1010 = {u_ca_out_1010[8:0],u_ca_out_1009[35:9], u_ca_out_1008[62:36], u_ca_out_1007[71:63]};
assign col_out_1011 = {u_ca_out_1011[8:0],u_ca_out_1010[35:9], u_ca_out_1009[62:36], u_ca_out_1008[71:63]};
assign col_out_1012 = {u_ca_out_1012[8:0],u_ca_out_1011[35:9], u_ca_out_1010[62:36], u_ca_out_1009[71:63]};
assign col_out_1013 = {u_ca_out_1013[8:0],u_ca_out_1012[35:9], u_ca_out_1011[62:36], u_ca_out_1010[71:63]};
assign col_out_1014 = {u_ca_out_1014[8:0],u_ca_out_1013[35:9], u_ca_out_1012[62:36], u_ca_out_1011[71:63]};
assign col_out_1015 = {u_ca_out_1015[8:0],u_ca_out_1014[35:9], u_ca_out_1013[62:36], u_ca_out_1012[71:63]};
assign col_out_1016 = {u_ca_out_1016[8:0],u_ca_out_1015[35:9], u_ca_out_1014[62:36], u_ca_out_1013[71:63]};
assign col_out_1017 = {u_ca_out_1017[8:0],u_ca_out_1016[35:9], u_ca_out_1015[62:36], u_ca_out_1014[71:63]};
assign col_out_1018 = {u_ca_out_1018[8:0],u_ca_out_1017[35:9], u_ca_out_1016[62:36], u_ca_out_1015[71:63]};
assign col_out_1019 = {u_ca_out_1019[8:0],u_ca_out_1018[35:9], u_ca_out_1017[62:36], u_ca_out_1016[71:63]};
assign col_out_1020 = {u_ca_out_1020[8:0],u_ca_out_1019[35:9], u_ca_out_1018[62:36], u_ca_out_1017[71:63]};
assign col_out_1021 = {u_ca_out_1021[8:0],u_ca_out_1020[35:9], u_ca_out_1019[62:36], u_ca_out_1018[71:63]};
assign col_out_1022 = {u_ca_out_1022[8:0],u_ca_out_1021[35:9], u_ca_out_1020[62:36], u_ca_out_1019[71:63]};
assign col_out_1023 = {u_ca_out_1023[8:0],u_ca_out_1022[35:9], u_ca_out_1021[62:36], u_ca_out_1020[71:63]};
assign col_out_1024 = {u_ca_out_1024[8:0],u_ca_out_1023[35:9], u_ca_out_1022[62:36], u_ca_out_1021[71:63]};
assign col_out_1025 = {u_ca_out_1025[8:0],u_ca_out_1024[35:9], u_ca_out_1023[62:36], u_ca_out_1022[71:63]};
assign col_out_1026 = {u_ca_out_1026[8:0],u_ca_out_1025[35:9], u_ca_out_1024[62:36], u_ca_out_1023[71:63]};
assign col_out_1027 = {u_ca_out_1027[8:0],u_ca_out_1026[35:9], u_ca_out_1025[62:36], u_ca_out_1024[71:63]};
assign col_out_1028 = {u_ca_out_1028[8:0],u_ca_out_1027[35:9], u_ca_out_1026[62:36], u_ca_out_1025[71:63]};
assign col_out_1029 = {u_ca_out_1029[8:0],u_ca_out_1028[35:9], u_ca_out_1027[62:36], u_ca_out_1026[71:63]};
assign col_out_1030 = {u_ca_out_1030[8:0],u_ca_out_1029[35:9], u_ca_out_1028[62:36], u_ca_out_1027[71:63]};
assign col_out_1031 = {u_ca_out_1031[8:0],u_ca_out_1030[35:9], u_ca_out_1029[62:36], u_ca_out_1028[71:63]};
assign col_out_1032 = {u_ca_out_1032[8:0],u_ca_out_1031[35:9], u_ca_out_1030[62:36], u_ca_out_1029[71:63]};
assign col_out_1033 = {u_ca_out_1033[8:0],u_ca_out_1032[35:9], u_ca_out_1031[62:36], u_ca_out_1030[71:63]};
assign col_out_1034 = {u_ca_out_1034[8:0],u_ca_out_1033[35:9], u_ca_out_1032[62:36], u_ca_out_1031[71:63]};
assign col_out_1035 = {u_ca_out_1035[8:0],u_ca_out_1034[35:9], u_ca_out_1033[62:36], u_ca_out_1032[71:63]};
assign col_out_1036 = {u_ca_out_1036[8:0],u_ca_out_1035[35:9], u_ca_out_1034[62:36], u_ca_out_1033[71:63]};
assign col_out_1037 = {u_ca_out_1037[8:0],u_ca_out_1036[35:9], u_ca_out_1035[62:36], u_ca_out_1034[71:63]};
assign col_out_1038 = {u_ca_out_1038[8:0],u_ca_out_1037[35:9], u_ca_out_1036[62:36], u_ca_out_1035[71:63]};
assign col_out_1039 = {u_ca_out_1039[8:0],u_ca_out_1038[35:9], u_ca_out_1037[62:36], u_ca_out_1036[71:63]};
assign col_out_1040 = {u_ca_out_1040[8:0],u_ca_out_1039[35:9], u_ca_out_1038[62:36], u_ca_out_1037[71:63]};
assign col_out_1041 = {u_ca_out_1041[8:0],u_ca_out_1040[35:9], u_ca_out_1039[62:36], u_ca_out_1038[71:63]};
assign col_out_1042 = {u_ca_out_1042[8:0],u_ca_out_1041[35:9], u_ca_out_1040[62:36], u_ca_out_1039[71:63]};
assign col_out_1043 = {u_ca_out_1043[8:0],u_ca_out_1042[35:9], u_ca_out_1041[62:36], u_ca_out_1040[71:63]};
assign col_out_1044 = {u_ca_out_1044[8:0],u_ca_out_1043[35:9], u_ca_out_1042[62:36], u_ca_out_1041[71:63]};
assign col_out_1045 = {u_ca_out_1045[8:0],u_ca_out_1044[35:9], u_ca_out_1043[62:36], u_ca_out_1042[71:63]};
assign col_out_1046 = {u_ca_out_1046[8:0],u_ca_out_1045[35:9], u_ca_out_1044[62:36], u_ca_out_1043[71:63]};
assign col_out_1047 = {u_ca_out_1047[8:0],u_ca_out_1046[35:9], u_ca_out_1045[62:36], u_ca_out_1044[71:63]};
assign col_out_1048 = {u_ca_out_1048[8:0],u_ca_out_1047[35:9], u_ca_out_1046[62:36], u_ca_out_1045[71:63]};
assign col_out_1049 = {u_ca_out_1049[8:0],u_ca_out_1048[35:9], u_ca_out_1047[62:36], u_ca_out_1046[71:63]};
assign col_out_1050 = {u_ca_out_1050[8:0],u_ca_out_1049[35:9], u_ca_out_1048[62:36], u_ca_out_1047[71:63]};
assign col_out_1051 = {u_ca_out_1051[8:0],u_ca_out_1050[35:9], u_ca_out_1049[62:36], u_ca_out_1048[71:63]};
assign col_out_1052 = {u_ca_out_1052[8:0],u_ca_out_1051[35:9], u_ca_out_1050[62:36], u_ca_out_1049[71:63]};
assign col_out_1053 = {u_ca_out_1053[8:0],u_ca_out_1052[35:9], u_ca_out_1051[62:36], u_ca_out_1050[71:63]};
assign col_out_1054 = {u_ca_out_1054[8:0],u_ca_out_1053[35:9], u_ca_out_1052[62:36], u_ca_out_1051[71:63]};
assign col_out_1055 = {u_ca_out_1055[8:0],u_ca_out_1054[35:9], u_ca_out_1053[62:36], u_ca_out_1052[71:63]};
assign col_out_1056 = {u_ca_out_1056[8:0],u_ca_out_1055[35:9], u_ca_out_1054[62:36], u_ca_out_1053[71:63]};
assign col_out_1057 = {u_ca_out_1057[8:0],u_ca_out_1056[35:9], u_ca_out_1055[62:36], u_ca_out_1054[71:63]};
assign col_out_1058 = {u_ca_out_1058[8:0],u_ca_out_1057[35:9], u_ca_out_1056[62:36], u_ca_out_1055[71:63]};
assign col_out_1059 = {u_ca_out_1059[8:0],u_ca_out_1058[35:9], u_ca_out_1057[62:36], u_ca_out_1056[71:63]};
assign col_out_1060 = {u_ca_out_1060[8:0],u_ca_out_1059[35:9], u_ca_out_1058[62:36], u_ca_out_1057[71:63]};
assign col_out_1061 = {u_ca_out_1061[8:0],u_ca_out_1060[35:9], u_ca_out_1059[62:36], u_ca_out_1058[71:63]};
assign col_out_1062 = {u_ca_out_1062[8:0],u_ca_out_1061[35:9], u_ca_out_1060[62:36], u_ca_out_1059[71:63]};
assign col_out_1063 = {u_ca_out_1063[8:0],u_ca_out_1062[35:9], u_ca_out_1061[62:36], u_ca_out_1060[71:63]};
assign col_out_1064 = {u_ca_out_1064[8:0],u_ca_out_1063[35:9], u_ca_out_1062[62:36], u_ca_out_1061[71:63]};
assign col_out_1065 = {u_ca_out_1065[8:0],u_ca_out_1064[35:9], u_ca_out_1063[62:36], u_ca_out_1062[71:63]};
assign col_out_1066 = {u_ca_out_1066[8:0],u_ca_out_1065[35:9], u_ca_out_1064[62:36], u_ca_out_1063[71:63]};
assign col_out_1067 = {u_ca_out_1067[8:0],u_ca_out_1066[35:9], u_ca_out_1065[62:36], u_ca_out_1064[71:63]};
assign col_out_1068 = {u_ca_out_1068[8:0],u_ca_out_1067[35:9], u_ca_out_1066[62:36], u_ca_out_1065[71:63]};
assign col_out_1069 = {u_ca_out_1069[8:0],u_ca_out_1068[35:9], u_ca_out_1067[62:36], u_ca_out_1066[71:63]};
assign col_out_1070 = {u_ca_out_1070[8:0],u_ca_out_1069[35:9], u_ca_out_1068[62:36], u_ca_out_1067[71:63]};
assign col_out_1071 = {u_ca_out_1071[8:0],u_ca_out_1070[35:9], u_ca_out_1069[62:36], u_ca_out_1068[71:63]};
assign col_out_1072 = {u_ca_out_1072[8:0],u_ca_out_1071[35:9], u_ca_out_1070[62:36], u_ca_out_1069[71:63]};
assign col_out_1073 = {u_ca_out_1073[8:0],u_ca_out_1072[35:9], u_ca_out_1071[62:36], u_ca_out_1070[71:63]};
assign col_out_1074 = {u_ca_out_1074[8:0],u_ca_out_1073[35:9], u_ca_out_1072[62:36], u_ca_out_1071[71:63]};
assign col_out_1075 = {u_ca_out_1075[8:0],u_ca_out_1074[35:9], u_ca_out_1073[62:36], u_ca_out_1072[71:63]};
assign col_out_1076 = {u_ca_out_1076[8:0],u_ca_out_1075[35:9], u_ca_out_1074[62:36], u_ca_out_1073[71:63]};
assign col_out_1077 = {u_ca_out_1077[8:0],u_ca_out_1076[35:9], u_ca_out_1075[62:36], u_ca_out_1074[71:63]};
assign col_out_1078 = {u_ca_out_1078[8:0],u_ca_out_1077[35:9], u_ca_out_1076[62:36], u_ca_out_1075[71:63]};
assign col_out_1079 = {u_ca_out_1079[8:0],u_ca_out_1078[35:9], u_ca_out_1077[62:36], u_ca_out_1076[71:63]};
assign col_out_1080 = {u_ca_out_1080[8:0],u_ca_out_1079[35:9], u_ca_out_1078[62:36], u_ca_out_1077[71:63]};
assign col_out_1081 = {u_ca_out_1081[8:0],u_ca_out_1080[35:9], u_ca_out_1079[62:36], u_ca_out_1078[71:63]};
assign col_out_1082 = {u_ca_out_1082[8:0],u_ca_out_1081[35:9], u_ca_out_1080[62:36], u_ca_out_1079[71:63]};
assign col_out_1083 = {u_ca_out_1083[8:0],u_ca_out_1082[35:9], u_ca_out_1081[62:36], u_ca_out_1080[71:63]};
assign col_out_1084 = {u_ca_out_1084[8:0],u_ca_out_1083[35:9], u_ca_out_1082[62:36], u_ca_out_1081[71:63]};
assign col_out_1085 = {u_ca_out_1085[8:0],u_ca_out_1084[35:9], u_ca_out_1083[62:36], u_ca_out_1082[71:63]};
assign col_out_1086 = {u_ca_out_1086[8:0],u_ca_out_1085[35:9], u_ca_out_1084[62:36], u_ca_out_1083[71:63]};
assign col_out_1087 = {u_ca_out_1087[8:0],u_ca_out_1086[35:9], u_ca_out_1085[62:36], u_ca_out_1084[71:63]};
assign col_out_1088 = {u_ca_out_1088[8:0],u_ca_out_1087[35:9], u_ca_out_1086[62:36], u_ca_out_1085[71:63]};
assign col_out_1089 = {u_ca_out_1089[8:0],u_ca_out_1088[35:9], u_ca_out_1087[62:36], u_ca_out_1086[71:63]};
assign col_out_1090 = {u_ca_out_1090[8:0],u_ca_out_1089[35:9], u_ca_out_1088[62:36], u_ca_out_1087[71:63]};
assign col_out_1091 = {u_ca_out_1091[8:0],u_ca_out_1090[35:9], u_ca_out_1089[62:36], u_ca_out_1088[71:63]};
assign col_out_1092 = {u_ca_out_1092[8:0],u_ca_out_1091[35:9], u_ca_out_1090[62:36], u_ca_out_1089[71:63]};
assign col_out_1093 = {u_ca_out_1093[8:0],u_ca_out_1092[35:9], u_ca_out_1091[62:36], u_ca_out_1090[71:63]};
assign col_out_1094 = {u_ca_out_1094[8:0],u_ca_out_1093[35:9], u_ca_out_1092[62:36], u_ca_out_1091[71:63]};
assign col_out_1095 = {u_ca_out_1095[8:0],u_ca_out_1094[35:9], u_ca_out_1093[62:36], u_ca_out_1092[71:63]};
assign col_out_1096 = {u_ca_out_1096[8:0],u_ca_out_1095[35:9], u_ca_out_1094[62:36], u_ca_out_1093[71:63]};
assign col_out_1097 = {u_ca_out_1097[8:0],u_ca_out_1096[35:9], u_ca_out_1095[62:36], u_ca_out_1094[71:63]};
assign col_out_1098 = {u_ca_out_1098[8:0],u_ca_out_1097[35:9], u_ca_out_1096[62:36], u_ca_out_1095[71:63]};
assign col_out_1099 = {u_ca_out_1099[8:0],u_ca_out_1098[35:9], u_ca_out_1097[62:36], u_ca_out_1096[71:63]};
assign col_out_1100 = {u_ca_out_1100[8:0],u_ca_out_1099[35:9], u_ca_out_1098[62:36], u_ca_out_1097[71:63]};
assign col_out_1101 = {u_ca_out_1101[8:0],u_ca_out_1100[35:9], u_ca_out_1099[62:36], u_ca_out_1098[71:63]};
assign col_out_1102 = {u_ca_out_1102[8:0],u_ca_out_1101[35:9], u_ca_out_1100[62:36], u_ca_out_1099[71:63]};
assign col_out_1103 = {u_ca_out_1103[8:0],u_ca_out_1102[35:9], u_ca_out_1101[62:36], u_ca_out_1100[71:63]};
assign col_out_1104 = {u_ca_out_1104[8:0],u_ca_out_1103[35:9], u_ca_out_1102[62:36], u_ca_out_1101[71:63]};
assign col_out_1105 = {u_ca_out_1105[8:0],u_ca_out_1104[35:9], u_ca_out_1103[62:36], u_ca_out_1102[71:63]};
assign col_out_1106 = {u_ca_out_1106[8:0],u_ca_out_1105[35:9], u_ca_out_1104[62:36], u_ca_out_1103[71:63]};
assign col_out_1107 = {u_ca_out_1107[8:0],u_ca_out_1106[35:9], u_ca_out_1105[62:36], u_ca_out_1104[71:63]};
assign col_out_1108 = {u_ca_out_1108[8:0],u_ca_out_1107[35:9], u_ca_out_1106[62:36], u_ca_out_1105[71:63]};
assign col_out_1109 = {u_ca_out_1109[8:0],u_ca_out_1108[35:9], u_ca_out_1107[62:36], u_ca_out_1106[71:63]};
assign col_out_1110 = {u_ca_out_1110[8:0],u_ca_out_1109[35:9], u_ca_out_1108[62:36], u_ca_out_1107[71:63]};
assign col_out_1111 = {u_ca_out_1111[8:0],u_ca_out_1110[35:9], u_ca_out_1109[62:36], u_ca_out_1108[71:63]};
assign col_out_1112 = {u_ca_out_1112[8:0],u_ca_out_1111[35:9], u_ca_out_1110[62:36], u_ca_out_1109[71:63]};
assign col_out_1113 = {u_ca_out_1113[8:0],u_ca_out_1112[35:9], u_ca_out_1111[62:36], u_ca_out_1110[71:63]};
assign col_out_1114 = {u_ca_out_1114[8:0],u_ca_out_1113[35:9], u_ca_out_1112[62:36], u_ca_out_1111[71:63]};
assign col_out_1115 = {u_ca_out_1115[8:0],u_ca_out_1114[35:9], u_ca_out_1113[62:36], u_ca_out_1112[71:63]};
assign col_out_1116 = {u_ca_out_1116[8:0],u_ca_out_1115[35:9], u_ca_out_1114[62:36], u_ca_out_1113[71:63]};
assign col_out_1117 = {u_ca_out_1117[8:0],u_ca_out_1116[35:9], u_ca_out_1115[62:36], u_ca_out_1114[71:63]};
assign col_out_1118 = {u_ca_out_1118[8:0],u_ca_out_1117[35:9], u_ca_out_1116[62:36], u_ca_out_1115[71:63]};
assign col_out_1119 = {u_ca_out_1119[8:0],u_ca_out_1118[35:9], u_ca_out_1117[62:36], u_ca_out_1116[71:63]};
assign col_out_1120 = {u_ca_out_1120[8:0],u_ca_out_1119[35:9], u_ca_out_1118[62:36], u_ca_out_1117[71:63]};
assign col_out_1121 = {u_ca_out_1121[8:0],u_ca_out_1120[35:9], u_ca_out_1119[62:36], u_ca_out_1118[71:63]};
assign col_out_1122 = {u_ca_out_1122[8:0],u_ca_out_1121[35:9], u_ca_out_1120[62:36], u_ca_out_1119[71:63]};
assign col_out_1123 = {u_ca_out_1123[8:0],u_ca_out_1122[35:9], u_ca_out_1121[62:36], u_ca_out_1120[71:63]};
assign col_out_1124 = {u_ca_out_1124[8:0],u_ca_out_1123[35:9], u_ca_out_1122[62:36], u_ca_out_1121[71:63]};
assign col_out_1125 = {u_ca_out_1125[8:0],u_ca_out_1124[35:9], u_ca_out_1123[62:36], u_ca_out_1122[71:63]};
assign col_out_1126 = {u_ca_out_1126[8:0],u_ca_out_1125[35:9], u_ca_out_1124[62:36], u_ca_out_1123[71:63]};
assign col_out_1127 = {u_ca_out_1127[8:0],u_ca_out_1126[35:9], u_ca_out_1125[62:36], u_ca_out_1124[71:63]};
assign col_out_1128 = {u_ca_out_1128[8:0],u_ca_out_1127[35:9], u_ca_out_1126[62:36], u_ca_out_1125[71:63]};
assign col_out_1129 = {u_ca_out_1129[8:0],u_ca_out_1128[35:9], u_ca_out_1127[62:36], u_ca_out_1126[71:63]};
assign col_out_1130 = {u_ca_out_1130[8:0],u_ca_out_1129[35:9], u_ca_out_1128[62:36], u_ca_out_1127[71:63]};
assign col_out_1131 = {u_ca_out_1131[8:0],u_ca_out_1130[35:9], u_ca_out_1129[62:36], u_ca_out_1128[71:63]};
assign col_out_1132 = {u_ca_out_1132[8:0],u_ca_out_1131[35:9], u_ca_out_1130[62:36], u_ca_out_1129[71:63]};
assign col_out_1133 = {u_ca_out_1133[8:0],u_ca_out_1132[35:9], u_ca_out_1131[62:36], u_ca_out_1130[71:63]};
assign col_out_1134 = {u_ca_out_1134[8:0],u_ca_out_1133[35:9], u_ca_out_1132[62:36], u_ca_out_1131[71:63]};
assign col_out_1135 = {u_ca_out_1135[8:0],u_ca_out_1134[35:9], u_ca_out_1133[62:36], u_ca_out_1132[71:63]};
assign col_out_1136 = {u_ca_out_1136[8:0],u_ca_out_1135[35:9], u_ca_out_1134[62:36], u_ca_out_1133[71:63]};
assign col_out_1137 = {u_ca_out_1137[8:0],u_ca_out_1136[35:9], u_ca_out_1135[62:36], u_ca_out_1134[71:63]};
assign col_out_1138 = {u_ca_out_1138[8:0],u_ca_out_1137[35:9], u_ca_out_1136[62:36], u_ca_out_1135[71:63]};
assign col_out_1139 = {u_ca_out_1139[8:0],u_ca_out_1138[35:9], u_ca_out_1137[62:36], u_ca_out_1136[71:63]};
assign col_out_1140 = {u_ca_out_1140[8:0],u_ca_out_1139[35:9], u_ca_out_1138[62:36], u_ca_out_1137[71:63]};
assign col_out_1141 = {u_ca_out_1141[8:0],u_ca_out_1140[35:9], u_ca_out_1139[62:36], u_ca_out_1138[71:63]};
assign col_out_1142 = {u_ca_out_1142[8:0],u_ca_out_1141[35:9], u_ca_out_1140[62:36], u_ca_out_1139[71:63]};
assign col_out_1143 = {u_ca_out_1143[8:0],u_ca_out_1142[35:9], u_ca_out_1141[62:36], u_ca_out_1140[71:63]};
assign col_out_1144 = {u_ca_out_1144[8:0],u_ca_out_1143[35:9], u_ca_out_1142[62:36], u_ca_out_1141[71:63]};
assign col_out_1145 = {u_ca_out_1145[8:0],u_ca_out_1144[35:9], u_ca_out_1143[62:36], u_ca_out_1142[71:63]};
assign col_out_1146 = {u_ca_out_1146[8:0],u_ca_out_1145[35:9], u_ca_out_1144[62:36], u_ca_out_1143[71:63]};
assign col_out_1147 = {u_ca_out_1147[8:0],u_ca_out_1146[35:9], u_ca_out_1145[62:36], u_ca_out_1144[71:63]};
assign col_out_1148 = {u_ca_out_1148[8:0],u_ca_out_1147[35:9], u_ca_out_1146[62:36], u_ca_out_1145[71:63]};
assign col_out_1149 = {u_ca_out_1149[8:0],u_ca_out_1148[35:9], u_ca_out_1147[62:36], u_ca_out_1146[71:63]};
assign col_out_1150 = {u_ca_out_1150[8:0],u_ca_out_1149[35:9], u_ca_out_1148[62:36], u_ca_out_1147[71:63]};
assign col_out_1151 = {u_ca_out_1151[8:0],u_ca_out_1150[35:9], u_ca_out_1149[62:36], u_ca_out_1148[71:63]};
assign col_out_1152 = {u_ca_out_1152[8:0],u_ca_out_1151[35:9], u_ca_out_1150[62:36], u_ca_out_1149[71:63]};
assign col_out_1153 = {u_ca_out_1153[8:0],u_ca_out_1152[35:9], u_ca_out_1151[62:36], u_ca_out_1150[71:63]};
assign col_out_1154 = {u_ca_out_1154[8:0],u_ca_out_1153[35:9], u_ca_out_1152[62:36], u_ca_out_1151[71:63]};
assign col_out_1155 = {u_ca_out_1155[8:0],u_ca_out_1154[35:9], u_ca_out_1153[62:36], u_ca_out_1152[71:63]};
assign col_out_1156 = {u_ca_out_1156[8:0],u_ca_out_1155[35:9], u_ca_out_1154[62:36], u_ca_out_1153[71:63]};
assign col_out_1157 = {u_ca_out_1157[8:0],u_ca_out_1156[35:9], u_ca_out_1155[62:36], u_ca_out_1154[71:63]};
assign col_out_1158 = {u_ca_out_1158[8:0],u_ca_out_1157[35:9], u_ca_out_1156[62:36], u_ca_out_1155[71:63]};
assign col_out_1159 = {u_ca_out_1159[8:0],u_ca_out_1158[35:9], u_ca_out_1157[62:36], u_ca_out_1156[71:63]};
assign col_out_1160 = {u_ca_out_1160[8:0],u_ca_out_1159[35:9], u_ca_out_1158[62:36], u_ca_out_1157[71:63]};
assign col_out_1161 = {u_ca_out_1161[8:0],u_ca_out_1160[35:9], u_ca_out_1159[62:36], u_ca_out_1158[71:63]};
assign col_out_1162 = {u_ca_out_1162[8:0],u_ca_out_1161[35:9], u_ca_out_1160[62:36], u_ca_out_1159[71:63]};
assign col_out_1163 = {u_ca_out_1163[8:0],u_ca_out_1162[35:9], u_ca_out_1161[62:36], u_ca_out_1160[71:63]};
assign col_out_1164 = {u_ca_out_1164[8:0],u_ca_out_1163[35:9], u_ca_out_1162[62:36], u_ca_out_1161[71:63]};
assign col_out_1165 = {u_ca_out_1165[8:0],u_ca_out_1164[35:9], u_ca_out_1163[62:36], u_ca_out_1162[71:63]};
assign col_out_1166 = {u_ca_out_1166[8:0],u_ca_out_1165[35:9], u_ca_out_1164[62:36], u_ca_out_1163[71:63]};
assign col_out_1167 = {u_ca_out_1167[8:0],u_ca_out_1166[35:9], u_ca_out_1165[62:36], u_ca_out_1164[71:63]};
assign col_out_1168 = {u_ca_out_1168[8:0],u_ca_out_1167[35:9], u_ca_out_1166[62:36], u_ca_out_1165[71:63]};
assign col_out_1169 = {u_ca_out_1169[8:0],u_ca_out_1168[35:9], u_ca_out_1167[62:36], u_ca_out_1166[71:63]};
assign col_out_1170 = {u_ca_out_1170[8:0],u_ca_out_1169[35:9], u_ca_out_1168[62:36], u_ca_out_1167[71:63]};
assign col_out_1171 = {u_ca_out_1171[8:0],u_ca_out_1170[35:9], u_ca_out_1169[62:36], u_ca_out_1168[71:63]};
assign col_out_1172 = {u_ca_out_1172[8:0],u_ca_out_1171[35:9], u_ca_out_1170[62:36], u_ca_out_1169[71:63]};
assign col_out_1173 = {u_ca_out_1173[8:0],u_ca_out_1172[35:9], u_ca_out_1171[62:36], u_ca_out_1170[71:63]};
assign col_out_1174 = {u_ca_out_1174[8:0],u_ca_out_1173[35:9], u_ca_out_1172[62:36], u_ca_out_1171[71:63]};
assign col_out_1175 = {u_ca_out_1175[8:0],u_ca_out_1174[35:9], u_ca_out_1173[62:36], u_ca_out_1172[71:63]};
assign col_out_1176 = {u_ca_out_1176[8:0],u_ca_out_1175[35:9], u_ca_out_1174[62:36], u_ca_out_1173[71:63]};
assign col_out_1177 = {u_ca_out_1177[8:0],u_ca_out_1176[35:9], u_ca_out_1175[62:36], u_ca_out_1174[71:63]};
assign col_out_1178 = {u_ca_out_1178[8:0],u_ca_out_1177[35:9], u_ca_out_1176[62:36], u_ca_out_1175[71:63]};
assign col_out_1179 = {u_ca_out_1179[8:0],u_ca_out_1178[35:9], u_ca_out_1177[62:36], u_ca_out_1176[71:63]};
assign col_out_1180 = {u_ca_out_1180[8:0],u_ca_out_1179[35:9], u_ca_out_1178[62:36], u_ca_out_1177[71:63]};
assign col_out_1181 = {u_ca_out_1181[8:0],u_ca_out_1180[35:9], u_ca_out_1179[62:36], u_ca_out_1178[71:63]};
assign col_out_1182 = {u_ca_out_1182[8:0],u_ca_out_1181[35:9], u_ca_out_1180[62:36], u_ca_out_1179[71:63]};
assign col_out_1183 = {u_ca_out_1183[8:0],u_ca_out_1182[35:9], u_ca_out_1181[62:36], u_ca_out_1180[71:63]};
assign col_out_1184 = {u_ca_out_1184[8:0],u_ca_out_1183[35:9], u_ca_out_1182[62:36], u_ca_out_1181[71:63]};
assign col_out_1185 = {u_ca_out_1185[8:0],u_ca_out_1184[35:9], u_ca_out_1183[62:36], u_ca_out_1182[71:63]};
assign col_out_1186 = {u_ca_out_1186[8:0],u_ca_out_1185[35:9], u_ca_out_1184[62:36], u_ca_out_1183[71:63]};
assign col_out_1187 = {u_ca_out_1187[8:0],u_ca_out_1186[35:9], u_ca_out_1185[62:36], u_ca_out_1184[71:63]};
assign col_out_1188 = {u_ca_out_1188[8:0],u_ca_out_1187[35:9], u_ca_out_1186[62:36], u_ca_out_1185[71:63]};
assign col_out_1189 = {u_ca_out_1189[8:0],u_ca_out_1188[35:9], u_ca_out_1187[62:36], u_ca_out_1186[71:63]};
assign col_out_1190 = {u_ca_out_1190[8:0],u_ca_out_1189[35:9], u_ca_out_1188[62:36], u_ca_out_1187[71:63]};
assign col_out_1191 = {u_ca_out_1191[8:0],u_ca_out_1190[35:9], u_ca_out_1189[62:36], u_ca_out_1188[71:63]};
assign col_out_1192 = {u_ca_out_1192[8:0],u_ca_out_1191[35:9], u_ca_out_1190[62:36], u_ca_out_1189[71:63]};
assign col_out_1193 = {u_ca_out_1193[8:0],u_ca_out_1192[35:9], u_ca_out_1191[62:36], u_ca_out_1190[71:63]};
assign col_out_1194 = {u_ca_out_1194[8:0],u_ca_out_1193[35:9], u_ca_out_1192[62:36], u_ca_out_1191[71:63]};
assign col_out_1195 = {u_ca_out_1195[8:0],u_ca_out_1194[35:9], u_ca_out_1193[62:36], u_ca_out_1192[71:63]};
assign col_out_1196 = {u_ca_out_1196[8:0],u_ca_out_1195[35:9], u_ca_out_1194[62:36], u_ca_out_1193[71:63]};
assign col_out_1197 = {u_ca_out_1197[8:0],u_ca_out_1196[35:9], u_ca_out_1195[62:36], u_ca_out_1194[71:63]};
assign col_out_1198 = {u_ca_out_1198[8:0],u_ca_out_1197[35:9], u_ca_out_1196[62:36], u_ca_out_1195[71:63]};
assign col_out_1199 = {u_ca_out_1199[8:0],u_ca_out_1198[35:9], u_ca_out_1197[62:36], u_ca_out_1196[71:63]};
assign col_out_1200 = {u_ca_out_1200[8:0],u_ca_out_1199[35:9], u_ca_out_1198[62:36], u_ca_out_1197[71:63]};
assign col_out_1201 = {u_ca_out_1201[8:0],u_ca_out_1200[35:9], u_ca_out_1199[62:36], u_ca_out_1198[71:63]};
assign col_out_1202 = {u_ca_out_1202[8:0],u_ca_out_1201[35:9], u_ca_out_1200[62:36], u_ca_out_1199[71:63]};
assign col_out_1203 = {u_ca_out_1203[8:0],u_ca_out_1202[35:9], u_ca_out_1201[62:36], u_ca_out_1200[71:63]};
assign col_out_1204 = {u_ca_out_1204[8:0],u_ca_out_1203[35:9], u_ca_out_1202[62:36], u_ca_out_1201[71:63]};
assign col_out_1205 = {u_ca_out_1205[8:0],u_ca_out_1204[35:9], u_ca_out_1203[62:36], u_ca_out_1202[71:63]};
assign col_out_1206 = {u_ca_out_1206[8:0],u_ca_out_1205[35:9], u_ca_out_1204[62:36], u_ca_out_1203[71:63]};
assign col_out_1207 = {u_ca_out_1207[8:0],u_ca_out_1206[35:9], u_ca_out_1205[62:36], u_ca_out_1204[71:63]};
assign col_out_1208 = {u_ca_out_1208[8:0],u_ca_out_1207[35:9], u_ca_out_1206[62:36], u_ca_out_1205[71:63]};
assign col_out_1209 = {u_ca_out_1209[8:0],u_ca_out_1208[35:9], u_ca_out_1207[62:36], u_ca_out_1206[71:63]};
assign col_out_1210 = {u_ca_out_1210[8:0],u_ca_out_1209[35:9], u_ca_out_1208[62:36], u_ca_out_1207[71:63]};
assign col_out_1211 = {u_ca_out_1211[8:0],u_ca_out_1210[35:9], u_ca_out_1209[62:36], u_ca_out_1208[71:63]};
assign col_out_1212 = {u_ca_out_1212[8:0],u_ca_out_1211[35:9], u_ca_out_1210[62:36], u_ca_out_1209[71:63]};
assign col_out_1213 = {u_ca_out_1213[8:0],u_ca_out_1212[35:9], u_ca_out_1211[62:36], u_ca_out_1210[71:63]};
assign col_out_1214 = {u_ca_out_1214[8:0],u_ca_out_1213[35:9], u_ca_out_1212[62:36], u_ca_out_1211[71:63]};
assign col_out_1215 = {u_ca_out_1215[8:0],u_ca_out_1214[35:9], u_ca_out_1213[62:36], u_ca_out_1212[71:63]};
assign col_out_1216 = {u_ca_out_1216[8:0],u_ca_out_1215[35:9], u_ca_out_1214[62:36], u_ca_out_1213[71:63]};
assign col_out_1217 = {u_ca_out_1217[8:0],u_ca_out_1216[35:9], u_ca_out_1215[62:36], u_ca_out_1214[71:63]};
assign col_out_1218 = {u_ca_out_1218[8:0],u_ca_out_1217[35:9], u_ca_out_1216[62:36], u_ca_out_1215[71:63]};
assign col_out_1219 = {u_ca_out_1219[8:0],u_ca_out_1218[35:9], u_ca_out_1217[62:36], u_ca_out_1216[71:63]};
assign col_out_1220 = {u_ca_out_1220[8:0],u_ca_out_1219[35:9], u_ca_out_1218[62:36], u_ca_out_1217[71:63]};
assign col_out_1221 = {u_ca_out_1221[8:0],u_ca_out_1220[35:9], u_ca_out_1219[62:36], u_ca_out_1218[71:63]};
assign col_out_1222 = {u_ca_out_1222[8:0],u_ca_out_1221[35:9], u_ca_out_1220[62:36], u_ca_out_1219[71:63]};
assign col_out_1223 = {u_ca_out_1223[8:0],u_ca_out_1222[35:9], u_ca_out_1221[62:36], u_ca_out_1220[71:63]};
assign col_out_1224 = {u_ca_out_1224[8:0],u_ca_out_1223[35:9], u_ca_out_1222[62:36], u_ca_out_1221[71:63]};
assign col_out_1225 = {u_ca_out_1225[8:0],u_ca_out_1224[35:9], u_ca_out_1223[62:36], u_ca_out_1222[71:63]};
assign col_out_1226 = {u_ca_out_1226[8:0],u_ca_out_1225[35:9], u_ca_out_1224[62:36], u_ca_out_1223[71:63]};
assign col_out_1227 = {u_ca_out_1227[8:0],u_ca_out_1226[35:9], u_ca_out_1225[62:36], u_ca_out_1224[71:63]};
assign col_out_1228 = {u_ca_out_1228[8:0],u_ca_out_1227[35:9], u_ca_out_1226[62:36], u_ca_out_1225[71:63]};
assign col_out_1229 = {u_ca_out_1229[8:0],u_ca_out_1228[35:9], u_ca_out_1227[62:36], u_ca_out_1226[71:63]};
assign col_out_1230 = {u_ca_out_1230[8:0],u_ca_out_1229[35:9], u_ca_out_1228[62:36], u_ca_out_1227[71:63]};
assign col_out_1231 = {u_ca_out_1231[8:0],u_ca_out_1230[35:9], u_ca_out_1229[62:36], u_ca_out_1228[71:63]};
assign col_out_1232 = {u_ca_out_1232[8:0],u_ca_out_1231[35:9], u_ca_out_1230[62:36], u_ca_out_1229[71:63]};
assign col_out_1233 = {u_ca_out_1233[8:0],u_ca_out_1232[35:9], u_ca_out_1231[62:36], u_ca_out_1230[71:63]};
assign col_out_1234 = {u_ca_out_1234[8:0],u_ca_out_1233[35:9], u_ca_out_1232[62:36], u_ca_out_1231[71:63]};
assign col_out_1235 = {u_ca_out_1235[8:0],u_ca_out_1234[35:9], u_ca_out_1233[62:36], u_ca_out_1232[71:63]};
assign col_out_1236 = {u_ca_out_1236[8:0],u_ca_out_1235[35:9], u_ca_out_1234[62:36], u_ca_out_1233[71:63]};
assign col_out_1237 = {u_ca_out_1237[8:0],u_ca_out_1236[35:9], u_ca_out_1235[62:36], u_ca_out_1234[71:63]};
assign col_out_1238 = {u_ca_out_1238[8:0],u_ca_out_1237[35:9], u_ca_out_1236[62:36], u_ca_out_1235[71:63]};
assign col_out_1239 = {u_ca_out_1239[8:0],u_ca_out_1238[35:9], u_ca_out_1237[62:36], u_ca_out_1236[71:63]};
assign col_out_1240 = {u_ca_out_1240[8:0],u_ca_out_1239[35:9], u_ca_out_1238[62:36], u_ca_out_1237[71:63]};
assign col_out_1241 = {u_ca_out_1241[8:0],u_ca_out_1240[35:9], u_ca_out_1239[62:36], u_ca_out_1238[71:63]};
assign col_out_1242 = {u_ca_out_1242[8:0],u_ca_out_1241[35:9], u_ca_out_1240[62:36], u_ca_out_1239[71:63]};
assign col_out_1243 = {u_ca_out_1243[8:0],u_ca_out_1242[35:9], u_ca_out_1241[62:36], u_ca_out_1240[71:63]};
assign col_out_1244 = {u_ca_out_1244[8:0],u_ca_out_1243[35:9], u_ca_out_1242[62:36], u_ca_out_1241[71:63]};
assign col_out_1245 = {u_ca_out_1245[8:0],u_ca_out_1244[35:9], u_ca_out_1243[62:36], u_ca_out_1242[71:63]};
assign col_out_1246 = {u_ca_out_1246[8:0],u_ca_out_1245[35:9], u_ca_out_1244[62:36], u_ca_out_1243[71:63]};
assign col_out_1247 = {u_ca_out_1247[8:0],u_ca_out_1246[35:9], u_ca_out_1245[62:36], u_ca_out_1244[71:63]};
assign col_out_1248 = {u_ca_out_1248[8:0],u_ca_out_1247[35:9], u_ca_out_1246[62:36], u_ca_out_1245[71:63]};
assign col_out_1249 = {u_ca_out_1249[8:0],u_ca_out_1248[35:9], u_ca_out_1247[62:36], u_ca_out_1246[71:63]};
assign col_out_1250 = {u_ca_out_1250[8:0],u_ca_out_1249[35:9], u_ca_out_1248[62:36], u_ca_out_1247[71:63]};
assign col_out_1251 = {u_ca_out_1251[8:0],u_ca_out_1250[35:9], u_ca_out_1249[62:36], u_ca_out_1248[71:63]};
assign col_out_1252 = {u_ca_out_1252[8:0],u_ca_out_1251[35:9], u_ca_out_1250[62:36], u_ca_out_1249[71:63]};
assign col_out_1253 = {u_ca_out_1253[8:0],u_ca_out_1252[35:9], u_ca_out_1251[62:36], u_ca_out_1250[71:63]};
assign col_out_1254 = {u_ca_out_1254[8:0],u_ca_out_1253[35:9], u_ca_out_1252[62:36], u_ca_out_1251[71:63]};
assign col_out_1255 = {u_ca_out_1255[8:0],u_ca_out_1254[35:9], u_ca_out_1253[62:36], u_ca_out_1252[71:63]};
assign col_out_1256 = {u_ca_out_1256[8:0],u_ca_out_1255[35:9], u_ca_out_1254[62:36], u_ca_out_1253[71:63]};
assign col_out_1257 = {u_ca_out_1257[8:0],u_ca_out_1256[35:9], u_ca_out_1255[62:36], u_ca_out_1254[71:63]};
assign col_out_1258 = {u_ca_out_1258[8:0],u_ca_out_1257[35:9], u_ca_out_1256[62:36], u_ca_out_1255[71:63]};
assign col_out_1259 = {u_ca_out_1259[8:0],u_ca_out_1258[35:9], u_ca_out_1257[62:36], u_ca_out_1256[71:63]};
assign col_out_1260 = {u_ca_out_1260[8:0],u_ca_out_1259[35:9], u_ca_out_1258[62:36], u_ca_out_1257[71:63]};
assign col_out_1261 = {u_ca_out_1261[8:0],u_ca_out_1260[35:9], u_ca_out_1259[62:36], u_ca_out_1258[71:63]};
assign col_out_1262 = {u_ca_out_1262[8:0],u_ca_out_1261[35:9], u_ca_out_1260[62:36], u_ca_out_1259[71:63]};
assign col_out_1263 = {u_ca_out_1263[8:0],u_ca_out_1262[35:9], u_ca_out_1261[62:36], u_ca_out_1260[71:63]};
assign col_out_1264 = {u_ca_out_1264[8:0],u_ca_out_1263[35:9], u_ca_out_1262[62:36], u_ca_out_1261[71:63]};
assign col_out_1265 = {u_ca_out_1265[8:0],u_ca_out_1264[35:9], u_ca_out_1263[62:36], u_ca_out_1262[71:63]};
assign col_out_1266 = {u_ca_out_1266[8:0],u_ca_out_1265[35:9], u_ca_out_1264[62:36], u_ca_out_1263[71:63]};
assign col_out_1267 = {u_ca_out_1267[8:0],u_ca_out_1266[35:9], u_ca_out_1265[62:36], u_ca_out_1264[71:63]};
assign col_out_1268 = {u_ca_out_1268[8:0],u_ca_out_1267[35:9], u_ca_out_1266[62:36], u_ca_out_1265[71:63]};
assign col_out_1269 = {u_ca_out_1269[8:0],u_ca_out_1268[35:9], u_ca_out_1267[62:36], u_ca_out_1266[71:63]};
assign col_out_1270 = {u_ca_out_1270[8:0],u_ca_out_1269[35:9], u_ca_out_1268[62:36], u_ca_out_1267[71:63]};
assign col_out_1271 = {u_ca_out_1271[8:0],u_ca_out_1270[35:9], u_ca_out_1269[62:36], u_ca_out_1268[71:63]};
assign col_out_1272 = {u_ca_out_1272[8:0],u_ca_out_1271[35:9], u_ca_out_1270[62:36], u_ca_out_1269[71:63]};
assign col_out_1273 = {u_ca_out_1273[8:0],u_ca_out_1272[35:9], u_ca_out_1271[62:36], u_ca_out_1270[71:63]};
assign col_out_1274 = {u_ca_out_1274[8:0],u_ca_out_1273[35:9], u_ca_out_1272[62:36], u_ca_out_1271[71:63]};
assign col_out_1275 = {u_ca_out_1275[8:0],u_ca_out_1274[35:9], u_ca_out_1273[62:36], u_ca_out_1272[71:63]};
assign col_out_1276 = {u_ca_out_1276[8:0],u_ca_out_1275[35:9], u_ca_out_1274[62:36], u_ca_out_1273[71:63]};
assign col_out_1277 = {u_ca_out_1277[8:0],u_ca_out_1276[35:9], u_ca_out_1275[62:36], u_ca_out_1274[71:63]};
assign col_out_1278 = {u_ca_out_1278[8:0],u_ca_out_1277[35:9], u_ca_out_1276[62:36], u_ca_out_1275[71:63]};
assign col_out_1279 = {u_ca_out_1279[8:0],u_ca_out_1278[35:9], u_ca_out_1277[62:36], u_ca_out_1276[71:63]};
assign col_out_1280 = {{9{1'b0}}, u_ca_out_1279[35:9], u_ca_out_1278[62:36], u_ca_out_1277[71:63]};
assign col_out_1281 = {{36{1'b0}}, u_ca_out_1279[62:36], u_ca_out_1278[71:63]};
assign col_out_1282 = {{63{1'b0}}, u_ca_out_1279[71:63]};

//---------------------------------------------------------


endmodule
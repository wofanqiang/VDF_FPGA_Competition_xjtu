module xpb_5_405
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h12e1db5da4496013188b918ffb856b5192d89aa69c8fa9e63c4c1ca3adcf4fab3d5a0c47586cf5cf64b33e8e9d8245545d3638b73b8e09d997373fdd3bb163e5bdd03944fc571462549b36c06c3d31375f206620c291d34ff8dc08d330c0457c6b1d36b5396f5e4c0de6122bd69351c578456a29ce8e6834cb3436617ea13ee8;
    5'b00010 : xpb = 1024'h25c3b6bb4892c0263117231ff70ad6a325b1354d391f53cc789839475b9e9f567ab4188eb0d9eb9ec9667d1d3b048aa8ba6c716e771c13b32e6e7fba7762c7cb7ba07289f8ae28c4a9366d80d87a626ebe40cc418523a69ff1b811a661808af8d63a6d6a72debc981bcc2457ad26a38af08ad4539d1cd06996686cc2fd427dd0;
    5'b00011 : xpb = 1024'h38a59218ecdc203949a2b4aff29041f4b889cff3d5aefdb2b4e455eb096def01b80e24d60946e16e2e19bbabd886cffd17a2aa25b2aa1d8cc5a5bf97b3142bb13970abcef5053d26fdd1a44144b793a61d61326247b579efea941a799240d0754157a41fac4e1ae429b2368383b9f55068d03e7d6bab389e619ca3247be3bcb8;
    5'b00100 : xpb = 1024'h4b876d769125804c622e463fee15ad464b626a9a723ea798f130728eb73d3eacf568311d61b3d73d92ccfa3a7609155174d8e2dcee3827665cdcff74eec58f96f740e513f15c5189526cdb01b0f4c4dd7c8198830a474d3fe370234cc30115f1ac74dad4e5bd7930379848af5a4d4715e115a8a73a39a0d32cd0d985fa84fba0;
    5'b00101 : xpb = 1024'h5e6948d4356ee05f7ab9d7cfe99b1897de3b05410ece517f2d7c8f32650c8e5832c23d64ba20cd0cf78038c9138b5aa5d20f1b9429c6313ff4143f522a76f37cb5111e58edb365eba70811c21d31f614dba1fea3ccd9208fdc4c2c1ff3c15b6e1792118a1f2cd77c457e5adb30e098db595b12d108c80907f8050fe779263a88;
    5'b00110 : xpb = 1024'h714b2431d9b840729345695fe52083e971139fe7ab5dfb6569c8abd612dbde03701c49ac128dc2dc5c337757b10d9ffa2f45544b65543b198b4b7f2f6628576272e1579dea0a7a4dfba34882896f274c3ac264c48f6af3dfd52834f32481a0ea82af483f589c35c853646d070773eaa0d1a07cfad756713cc3394648f7c77970;
    5'b00111 : xpb = 1024'h842cff8f7e01a085abd0faefe0a5ef3b03ec3a8e47eda54ba614c879c0ab2daead7655f36afab8abc0e6b5e64e8fe54e8c7b8d02a0e244f32282bf0ca1d9bb4830b190e2e6618eb0503e7f42f5ac588399e2cae551fcc72fce043dc65541e666edcc7ef4920b9414614a7f32de073c6649e5e724a5e4d9718e6d7caa7668b858;
    5'b01000 : xpb = 1024'h970edaed224b0098c45c8c7fdc2b5a8c96c4d534e47d4f31e260e51d6e7a7d59ead0623ac367ae7b2599f474ec122aa2e9b1c5b9dc704eccb9b9fee9dd8b1f2dee81ca27e2b8a312a4d9b60361e989baf9033106148e9a7fc6e0469986022be358e9b5a9cb7af2606f30915eb49a8e2bc22b514e747341a659a1b30bf509f740;
    5'b01001 : xpb = 1024'ha9f0b64ac69460abdce81e0fd7b0c5de299d6fdb810cf9181ead01c11c49cd05282a6e821bd4a44a8a4d330389946ff746e7fe7117fe58a650f13ec7193c8313ac52036cdf0fb774f974ecc3ce26baf258239726d7206dcfbfbc4f6cb6c2715fc406ec5f04ea50ac7d16a38a8b2ddff13a70bb784301a9db24d5e96d73ab3628;
    5'b01010 : xpb = 1024'hc254c52a8ef8bf62a6e37c8c2dbe9de4b00075148250286dd1c650f17166fa8623bfd50aa1b1b8b4fa2324b43b8a48140040f4230d9923437893f461a1b7247f5d308032bd5ce923b7620e1a18827f8c33f03af0d2c140f030bc6452d58144a001c90ea8d90b66b043cced769f10b8d63dc46bfc144b4dfa99aa4ca696a0ea5;
    5'b01011 : xpb = 1024'h1f0727b04d38ec0942f9c958be61552fddd8a1f7e4b4ac6d196881b2c4e5bf539f9609980288115ab45570d9e13ae9d59d3a47f96c679c0dcec07f2355ccd62db3a34148282ce2f4901157a20dc55930225f69cfcfbde75efbe7cf185e1859c66b39c79fc70014b71222e10340845d52dc21b0e98fd31d1474cedb2be80b4d8d;
    5'b01100 : xpb = 1024'h31e9030df1824c1c5b855ae8b9e6c08170b13c9e8144565355b49e5672b50efedcf015df5af5072a1908af687ebd2f29fa7080b0a7f5a5e765f7bf00917e3a1371737a8d2483f756e4ac8e627a028a67817fcff0924fbaaef4c3d7eb8ed89f42d656fe55006f73032008f32f1717af1854671b135e6185494003118d66ac8c75;
    5'b01101 : xpb = 1024'h44cade6b95cbac2f7410ec78b56c2bd30389d7451dd400399200bafa20845eaa1a4a2226b361fcf97dbbedf71c3f747e57a6b967e383afc0fd2efeddcd2f9df92f43b3d220db0bb93947c522e63fbb9ee0a0361154e18dfeed9fe0bebf98e4bf4174350a39ded14f2def055aedab00ddccac853d2cefed7e0b3747eee54dcb5d;
    5'b01110 : xpb = 1024'h57acb9c93a150c428c9c7e08b0f19724966271ebba63aa1fce4cd79dce53ae5557a42e6e0bcef2c8e26f2c85b9c1b9d2b4dcf21f1f11b99a94663ebb08e101deed13ed171d32201b8de2fbe3527cecd63fc09c321773614ee67be991f0592a3bac916bbf734e2f9b3bd51786c43e52a344f1ef66fb7e55b2d66b7e5063ef0a45;
    5'b01111 : xpb = 1024'h6a8e9526de5e6c55a5280f98ac770276293b0c9256f354060a98f4417c22fe0094fe3ab5643be89847226b145743ff2712132ad65a9fc3742b9d7e98449265c4aae4265c1989347de27e32a3beba1e0d9ee10252da05349edf57f26521196fb817aea274acbd8de749bb29b29ad1a468bd375990ca0cbde7a19fb4b1e290492d;
    5'b10000 : xpb = 1024'h7d70708482a7cc68bdb3a128a7fc6dc7bc13a738f382fdec46e510e529f24dabd25846fcbca8de67abd5a9a2f4c6447b6f49638d962dcd4dc2d4be758043c9aa68b45fa115e048e0371969642af74f44fe0168739c9707eed833fb3851d9b53482cbd929e62cec3357a13bde7164f62e357cc3ba989b261c6cd3eb1361318815;
    5'b10001 : xpb = 1024'h90524be226f12c7bd63f32b8a381d9194eec41df9012a7d283312d88d7c19d570fb253441515d4371088e831924889cfcc7f9c44d1bbd7275a0bfe52bbf52d90268498e612375d428bb4a0249734807c5d21ce945f28db3ed110040b8299fab0ede90fdf1f9c4a7f65874e0a47f847f3adc22de467298e5138082174dfd2c6fd;
    5'b10010 : xpb = 1024'ha334273fcb3a8c8eeecac4489f07446ae1c4dc862ca251b8bf7d4a2c8590ed024d0c5f8b6d82ca06753c26c02fcacf2429b5d4fc0d49e100f1433e2ff7a69175e454d22b0e8e71a4e04fd6e50371b1b3bc4234b521baae8ec9ec0cdeb35a402d59064694590ba8cb736d60361e8b99b92607980e35b7f686033c57d65e7405e5;
    5'b10011 : xpb = 1024'h568bd47ad95b7d93c50de018a32686b032773fbf3ba5b277decad7a805d8fa5871dee59fbc941473a912607e9ef03ae22d1e5cd26251a8ed7db3eaef88580aa2dd5d6c15b5488c222510b02d6d31eba275da13d57c654ce0d3b83b729efe317951beb1fe1b20e89fa938b82fd4ec5554f732355b3fb018a880113335432de62;
    5'b10100 : xpb = 1024'h184a98a551df17ec54dc6f9185b7d3bc96000ea2904a050dba38ca1e2e2cdf50c477faa1543637169f4464968771490280081e8461b324686f127e8c3436e48feba6100657ab9d2476ec41c343104ff1867e075e1a58281e06178c8a5ab02894003921d51b216cd608799daed3e2171ac7b88d7f828969bf53354994d2d41d4a;
    5'b10101 : xpb = 1024'h2b2c7402f62877ff6d680121813d3f0e28d8a9492cd9aef3f684e6c1dbfc2efc01d206e8aca32ce603f7a32524f38e56dd3e573b9d412e420649be696fe84875a976494b5402b186cb877883af4d8128e59e6d7edce9fb6dfef3955d8b706e106b56588a5490cb22165fafdaaa7568e03ffdf7a95117d1f41e697ff651755c32;
    5'b10110 : xpb = 1024'h3e0e4f609a71d81285f392b17cc2aa5fbbb143efc96958da32d1036589cb7ea73f2c1330051022b568aae1b3c275d3ab3a748ff2d8cf381b9d80fe46ab99ac5b674682905059c5e92022af441b8ab26044bed39f9f7bcebdf7cf9e30bc30b38cd6738f3f8e00296e2445c2068108baa5b84361d31fa63a28e99db657d0169b1a;
    5'b10111 : xpb = 1024'h50f02abe3ebb38259e7f2441784815b14e89de9665f902c06f1d2009379ace527c861f775d7d1884cd5e20425ff818ff97aac8aa145d41f534b83e23e74b10412516bbd54cb0da4b74bde60487c7e397a3df39c0620da20df0aba703ecf0f9094190c5f4c76f87ba322bd432579c0c6b3088cbfcee34a25db4d1ecb94eb7da02;
    5'b11000 : xpb = 1024'h63d2061be3049838b70ab5d173cd8102e162793d0288aca6ab693cace56a1dfdb9e02bbeb5ea0e5432115ed0fd7a5e53f4e101614feb4bcecbef7e0122fc7426e2e6f51a4907eeadc9591cc4f40514cf02ff9fe1249f755de987afd71db13e85acadfcaa00dee6064011e65e2e2f5e30a8ce3626bcc30a928006231acd5918ea;
    5'b11001 : xpb = 1024'h76b3e179874df84bcf9647616f52ec54743b13e39f18568ce7b5595093396da8f73a38060e57042396c49d5f9afca3a852173a188b7955a86326bdde5eadd80ca0b72e5f455f03101df453856042460662200601e73148ade263b8aa4e71840217cb335f3a4e44524df7f88a04c2aff62113a0508b5172c74b3a597c4bfa57d2;
    5'b11010 : xpb = 1024'h8995bcd72b97585ee821d8f16ad857a60713ae8a3ba80073240175f44108bd543494444d66c3f9f2fb77dbee387ee8fcaf4d72cfc7075f81fa5dfdbb9a5f3bf25e8767a441b61772728f8a45cc7f773dc1406c22a9c31bfddb3fc17d7f31c97e82e86a1473bda29e5bde0ab5db5601bb99590a7a59dfdafc166e8fddca9b96ba;
    5'b11011 : xpb = 1024'h9c779834cfe0b87200ad6a81665dc2f799ec4930d837aa59604d9297eed80cff71ee5094bf30efc2602b1a7cd6012e510c83ab870295695b91953d98d6109fd81c57a0e93e0d2bd4c72ac10638bca8752060d2436c54ef4dd41bca50aff20efaee05a0c9ad2d00ea69c41ce1b1e95381119e74a4286e4330e1a2c63f493cd5a2;
    5'b11100 : xpb = 1024'haf597392742a18851938fc1161e32e492cc4e3d774c7543f9c99af3b9ca75caaaf485cdc179de591c4de590b738373a569b9e43e3e23733528cc7d7611c203bdda27da2e3a6440371bc5f7c6a4f9d9ac7f8138642ee6c29dccf7d323e0b254775922d77ee69c5f3677aa2f0d887ca54689e3decdf6fcab65acd6fca0c7de148a;
    5'b11101 : xpb = 1024'h118e099a568543cf66bf15ca4d0e52494e277b4d3bdf5dae5b0912899773ff4de959ebaaa5e45cd28a3358532da7a82f62d5f50f56feacc30f647df512a0f2f223a8dec4872a57545dc72be4785b46b2ea9ca4ec64f268dd104749fc5747f76195387c0a6f42c4f4fed05a5a673fd0e2b34f6a15753fb66a319bb7fdbd9ced07;
    5'b11110 : xpb = 1024'h246fe4f7facea3e27f4aa75a4893bd9ae10015f3d86f079497552f2d45434ef926b3f7f1fe5152a1eee696e1cb29ed83c00c2dc6928cb69ca69bbdd24e5256d7e179180983816bb6b26262a4e49877ea49bd0b0d27843c2d092352cf88083cde0055b2bfa8b223410cb66c863dd322a82b94d43f43ce1e9efccfee5f3c3e2bef;
    5'b11111 : xpb = 1024'h3751c0559f1803f597d638ea441928ec73d8b09a74feb17ad3a14bd0f3129ea4640e043956be48715399d57068ac32d81d42667dce1ac0763dd2fdaf8a03babd9f49514e7fd8801906fd996550d5a921a8dd712dea160f7d01ff5ba2b8c8825a6b72e974e221818d1a9c7eb21466746da3da3e69125c86d3c80424c0badf6ad7;
    endcase
end

endmodule

module xpb_5_615
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h91795d36db13ad1787d51649859dbad552353b470ae3220cd7778279cd31483c65a2b89baf40f10ea88552b0648d39bb7b7e6dd34d97785b5f7b7291bc3f1508bc6da968aa4794db856889aa525c2ce9caa7f4075373f9f2135b55ba8213f56f9637f72e820d09cc450ab14d64daa0a3ea22d4bf7eac091a8111f3b4cb8c2512;
    5'b00010 : xpb = 1024'h72457517f439256644a4b4bbfae12e5932f4735d404ea3a231124b9de75fe370c7fcf3be945b638eb1ac6619e5bc62ac92e2b3c0787c206b0e57a5c53dabb560048c1e22a4fe2c71f83710b20bdc95a2a14aee761a61c6d3712a197a49fd484cfd685c3353511b0b03557bbbd1e51b1e856bca9cad0cb504bbb46c650e35e3b9;
    5'b00011 : xpb = 1024'h53118cf90d5e9db50174532e7024a1dd13b3ab7375ba25378aad14c2018e7ea52a572ee17975d60ebad3798366eb8b9daa46f9ada360c87abd33d8f8bf1855b74caa92dc9fb4c4086b0597b9c55cfe5b77ede8e4e14f93b4cef8dd3a11e69b2a6498c13824952c49c1a0462a3eef959920b4c079db6d60eef656e51550dfa260;
    5'b00100 : xpb = 1024'h33dda4da26841603be43f1a0e5681560f472e389ab25a6cce447dde61bbd19d98cb16a045e90488ec3fa8cece81ab48ec1ab3f9ace45708a6c100c2c4084f60e94c907969a6b5b9eddd41ec17edd67144e90e353a83d60962cc7a0f9d9cfee07cbc9263cf5d93d887feb1098abfa1013bbfdb65709ce0cd930f95dc593896107;
    5'b00101 : xpb = 1024'h14a9bcbb3fa98e527b1390135aab88e4d5321b9fe09128623de2a70a35ebb50def0ba52743aabb0ecd21a0566949dd7fd90f8587f92a189a1aec3f5fc1f19665dce77c509521f33550a2a5c9385dcfcd2533ddc26f2b2d778a9664b9a1b940e532f98b41c71d4ec73e35db0719048a8e5746ac34382eb8c36b9bd675d6331fae;
    5'b00110 : xpb = 1024'ha62319f21abd3b6a02e8a65ce04943ba276756e6eb744a6f155a2984031cfd4a54ae5dc2f2ebac1d75a6f306cdd7173b548df35b46c190f57a67b1f17e30ab6e995525b93f698810d60b2f738ab9fcb6efdbd1c9c29f27699df1ba7423cd3654c9318270492a589383408c547ddf2b32416980f3b6dac1ddecadca2aa1bf44c0;
    5'b00111 : xpb = 1024'h86ef31d333e2b3b8bfb844cf558cb73e08268efd20dfcc046ef4f2a81d4b987eb70898e5d8061e9d7ece06704f06402c6bf2394871a639052943e524ff9d4bc5e1739a733a201fa748d9b67b443a656fc67ecc38898cf44afbc07e33ebb689323061e7751a6e69d2418b56c2eae9a5acdcb276d0e53b6dc8275042dae4690367;
    5'b01000 : xpb = 1024'h67bb49b44d082c077c87e341cad02ac1e8e5c713564b4d99c88fbbcc377a33b31962d408bd20911d87f519d9d035691d83567f359c8ae114d82018588109ec1d29920f2d34d6b73dbba83d82fdbace289d21c6a7507ac12c598f41f3b39fdc0f97924c79ebb27b10ffd6213157f4202777fb6cae139c19b261f2bb8b2712c20e;
    5'b01001 : xpb = 1024'h48876195662da456395781b440139e45c9a4ff298bb6cf2f222a84f051a8cee77bbd0f2ba23b039d911c2d435164920e9abac522c76f892486fc4b8c02768c7471b083e72f8d4ed42e76c48ab73b36e173c4c11617688e0db75e05b37b892eecfec2b17ebcf68c4fbe20eb9fc4fe9aa21344628b41fcc59c9c95343b69bc80b5;
    5'b01010 : xpb = 1024'h295379767f531ca4f6272026b55711c9aa64373fc12250c47bc54e146bd76a1bde174a4e8755761d9a4340acd293baffb21f0b0ff254313435d87ebf83e32ccbb9cef8a12a43e66aa1454b9270bb9f9a4a67bb84de565aef152cc973437281ca65f316838e3a9d8e7c6bb60e3209151cae8d5868705d7186d737acebac663f5c;
    5'b01011 : xpb = 1024'ha1f9157987894f3b2f6be992a9a854d8b236f55f68dd259d560173886060550407185716c6fe89da36a541653c2e3f0c98350fd1d38d943e4b4b1f3054fcd2301ed6d5b24fa7e011413d29a2a3c0853210ab5f3a54427d072fb8d330b5bd4a7cd237b885f7eaecd3ab6807c9f138f9749d64e459ebe1d7111da259bef0ffe03;
    5'b01100 : xpb = 1024'h9b98ee8e738c420b3acbd4e2b0384022dd58aa9d0170f466acd799b253374d8ca6143e0d1bb0d9ac4befa6c6b8501dac4501bed06ad0519f44302484c18ee22bbe5b16c3cf4212dc997c5c447c98353cebb2a9faf8b821c28656e2ed8d6fca17635b72b6e18bb8997fc131ca03ee303b33f923051d6a268b92ec1950ba9c2315;
    5'b01101 : xpb = 1024'h7c65066f8cb1ba59f79b7355257bb3a6be17e2b336dc75fc067262d66d65e8c1086e793000cb4c2c5516ba30397f469d5c6604bd95b4f9aef30c57b842fb828306798b7dc9f8aa730c4ae34c36189df5c255a469bfa5eea3e425a6ad55591cf4ca8bd7bbb2cfc9d83e0bfc3870f8aab5cf4218e24bcad275cd8e9200fd45e1bc;
    5'b01110 : xpb = 1024'h5d311e50a5d732a8b46b11c79abf272a9ed71ac96c47f791600d2bfa879483f56ac8b452e5e5beac5e3dcd99baae6f8e73ca4aaac099a1bea1e88aebc46822da4e980037c4af42097f196a53ef9906ae98f89ed88693bb8541f46a6d1d426fd231bc3cc08413db16fc56c6a6de0325306a8b0ebf7a2b7e6008310ab13fefa063;
    5'b01111 : xpb = 1024'h3dfd3631befcaaf7713ab03a10029aae7f9652dfa1b37926b9a7f51ea1c31f29cd22ef75cb00312c6764e1033bdd987f8b2e9097eb7e49ce50c4be1f45d4c33196b674f1bf65d99ff1e7f15ba9196f676f9b99474d8188669fc32e2ce52bc2af98eca1c55557ec55baa191154b0d9fab05d4049ca88c2a4a42d3836182995f0a;
    5'b10000 : xpb = 1024'h1ec94e12d82223462e0a4eac85460e3260558af5d71efabc1342be42bbf1ba5e2f7d2a98b01aa3ac708bf46cbd0cc170a292d6851662f1ddffa0f152c7416388ded4e9abba1c713664b678636299d820463e93b6146f5547fd91f1ecad15158d001d06ca269bfd9478ec5b83b8181a25a11cfa79d6ecd6347d75fc11c5431db1;
    5'b10001 : xpb = 1024'hb042ab49b335d05db5df64f60ae3c907b28ac63ce2021cc8eaba40bc8923029a951fe3345f5b94bb1911471d2199fb2c1e11445863fa6a395f1c63e4838078919b42931464640611ea1f020db4f6050a10e687bd67e34f3a10ed47a72f290afc9654fdf8a8a90760bdf70cd11cf2bac98b3fcf395598df4efe87efc690cf42c3;
    5'b10010 : xpb = 1024'h910ec32acc5b48ac72af036880273c8b9349fe53176d9e5e445509e0a3519dcef77a1e574476073b22385a86a2c9241d35758a458edf12490df8971804ed18e8e36107ce5f1a9da85ced89156e766dc2e789822c2ed11c1b6ebc0b66f7125dd9fd8562fd79ed189f7c41d73f89fd35442688c51683f98b39392a6876d379016a;
    5'b10011 : xpb = 1024'h71dadb0be580c0fb2f7ea1daf56ab00f740936694cd91ff39defd304bd80390359d4597a299079bb2b5f6df023f84d0e4cd9d032b9c3ba58bcd4ca4b8659b9402b7f7c8859d1353ecfbc101d27f6d67bbe2c7c9af5bee8fccc8acf26befbb0b764b5c8024b3129de3a8ca1adf707afbec1d1baf3b25a372373cce1271622c011;
    5'b10100 : xpb = 1024'h52a6f2ecfea63949ec4e404d6aae239354c86e7f8244a188f78a9c28d7aed437bc2e949d0eaaec3b34868159a52775ff643e161fe4a862686bb0fd7f07c65997739df1425487ccd5428a9724e1773f3494cf7709bcacb5de2a5992e686e50394cbe62d071c753b1cf8d76c1c64122a395d1ab0d0e0bae30dae6f59d758cc7eb8;
    5'b10101 : xpb = 1024'h33730ace17cbb198a91ddebfdff197173587a695b7b0231e5125654cf1dd6f6c1e88cfbff3c55ebb3dad94c326569ef07ba25c0d0f8d0a781a8d30b28932f9eebbbc65fc4f3e646bb5591e2c9af7a7ed6b727178839a82bf882856a64ece56723316920bedb94c5bb722368ad11ca4b3f863a6ae0f1b8ef7e911d2879b763d5f;
    5'b10110 : xpb = 1024'h143f22af30f129e765ed7d3255350a9b1646deabed1ba4b3aac02e710c0c0aa080e30ae2d8dfd13b46d4a82ca785c7e19306a1fa3a71b287c96963e60a9f9a4603dadab649f4fc022827a534547810a642156be74a884fa0e5f71a6616b7a94f9a46f710befd5d9a756d00f93e271f2e93ac9c8b3d7c3ae223b44b37de1ffc06;
    5'b10111 : xpb = 1024'ha5b87fe60c04d6feedc2937bdad2c570687c19f2f7fec6c08237b0ead93d52dce685c37e8820c249ef59fadd0c13019d0e850fcd88092ae328e4d677c6deaf4ec048841ef43c90ddad902edea6d43d900cbd5fee9dfc4992f952702098cb9ebf307eee3f410a6766ba77b246a301bfd27dcf714abc2843fca4c63eeca9ac2118;
    5'b11000 : xpb = 1024'h868497c7252a4f4daa9231ee501638f4493b52092d6a4855dbd27a0ef36bee1148dffea16d3b34c9f8810e468d422a8e25e955bab2edd2f2d7c109ab484b4fa60866f8d8eef32874205eb5e66054a648e3605a5d64ea1674572133e060b4f19c97af5344124e78a578c27cb5100c3a4d19186727ea88efe6df68b79cec55dfbf;
    5'b11001 : xpb = 1024'h6750afa83e4fc79c6761d060c559ac7829fa8a1f62d5c9eb356d43330d9a8945ab3a39c45255a74a01a821b00e71537f3d4d9ba7ddd27b02869d3cdec9b7effd50856d92e9a9c00a932d3cee19d50f01ba0354cc2bd7e355b4eff7a0289e4479fedfb848e39289e4370d47237d16b4c7b4615d0518e99bd11a0b304d2eff9e66;
    5'b11010 : xpb = 1024'h481cc78957753feb24316ed33a9d1ffc0ab9c23598414b808f080c5727c9247a0d9474e7377019ca0acf35198fa07c7054b1e19508b72312357970124b24905498a3e24ce46057a105fbc3f5d35577ba90a64f3af2c5b03712bebb5ff087975766101d4db4d69b22f5581191ea212f424faa52e2474a47bb54ada8fd71a95d0d;
    5'b11011 : xpb = 1024'h28e8df6a709ab839e1010d45afe0937feb78fa4bcdaccd15e8a2d57b41f7bfae6feeb00a1c8a8c4a13f6488310cfa5616c162782339bcb21e455a345cc9130abe0c25706df16ef3778ca4afd8cd5e073674949a9b9b37d18708d7f1fb870ea34cd408252861aac61b3a2dc00572ba9bceaf348bf75aaf3a58f5021adb4531bb4;
    5'b11100 : xpb = 1024'h9b4f74b89c030889dd0abb825240703cc38326203184eab423d9e9f5c265ae2d248eb2d01a4feca1d1d5bec91fece52837a6d6f5e8073319331d6794dfdd10328e0cbc0d9cd86cdeb98d2054656492c3dec441880a149f9ce5c42df805a3d123470e757575ebda071eda66ec4362437863c3e9ca40b9f8fc9f29a5df6fcda5b;
    5'b11101 : xpb = 1024'h9b2e548264d3dda025a5c201aac1c1d91e6d6da90dfb70b819b521192957a31f37eba3c8b0e5efd8c5a2ae9cf68c080dfef8db42ac17eb8cf2ad490b0a3ce60be54e752984151ba971015baf98b276160894381fd41543ebe1b7989a026e3281caa8de85d96bc76cb6f857bc2910c4db705f135c22b7a8aa4b048e12c288ff6d;
    5'b11110 : xpb = 1024'h7bfa6c637df955eee27560742005355cff2ca5bf4366f24d734fea3d43863e539a45deeb96006258cec9c20677bb30ff165d212fd6fc939ca1897c3e8ba986632d6ce9e37ecbb33fe3cfe2b75232decedf37328e9b0310cd3f865c59ca57855f31d9438aaaafd8ab7543222a961b3f560ba809395118549485a706c30532be14;
    5'b11111 : xpb = 1024'h5cc68444971ece3d9f44fee69548a8e0dfebddd578d273e2cceab3615db4d987fca01a0e7b1ad4d8d7f0d56ff8ea59f02dc1671d01e13bac5065af720d1626ba758b5e9d79824ad6569e69bf0bb34787b5da2cfd61f0ddae9d5520199240d83c9909a88f7bf3e9ea338dec990325b9d0a6f0ff167f79007ec0497f7347dc7cbb;
    endcase
end

endmodule

module xpb_5_435
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h9604e039cf8ac97261c3d30faddab891c685825de2d94ca2e54f699877748c248ae16ba47a14a95e0ff9601c76f0598d100302c96ce24e4bbf9d3a17fd6ecc905ad04b3bd58b186e9e5607b5d7e077a3d530208e6df973e08a8c6341452a6ae094bdd10479724a5f2763243fe44c318c70419b7c5fda7ad0dbed25c62e560d40;
    5'b00010 : xpb = 1024'h7b5c7b1ddd275e1bf8822e484b5b29d21b95018af03af8ce4cc219db3be66b41127a59d02a02d42d809480f20a82a24fbbebddacb711cc4bce9b34d1c00b246f415161c8fb8533982a120cc916e52b16b65b47844f6cbab05f8c3487d02a332efa740fdf421b9c30c80661a0d0c83cef91a958166f699871716ad087d3c9b415;
    5'b00011 : xpb = 1024'h60b41601eac3f2c58f408980e8db9b1270a480b7fd9ca4f9b434ca1e00584a5d9a1347fbd9f0fefcf12fa1c79e14eb1267d4b89001414a4bdd992f8b82a77c4e27d27856217f4ec1b5ce11dc55e9de8997866e7a30e00180348c05ce5b29fb7d602a4eba0ac4ee0268a99f01bd444852b31114b07ef8b61206e87b49793d5aea;
    5'b00100 : xpb = 1024'h460bb0e5f860876f25fee4b9865c0c52c5b3ffe50afe51251ba77a60c4ca297a21ac362789df29cc61cac29d31a733d513bd93734b70c84bec972a454543d42d0e538ee3477969eb418a16ef94ee91fc78b1957012534850098bd714e629c3cbc5e08d94d36e3fd4094cdc62a9c053b5d478d14a8e87d3b29c66260b1eb101bf;
    5'b00101 : xpb = 1024'h2b634bca05fd1c18bcbd3ff223dc7d931ac37f12185ffd50831a2aa3893c0896a945245339cd549bd265e372c5397c97bfa66e5695a0464bfb9524ff07e02c0bf4d4a5706d738514cd461c02d3f3456f59dcbc65f3c68f1fde8ba85b71298c1a2b96cc6f9c1791a5a9f019c3963c5f18f5e08de49e16f15331e3d0ccc424a894;
    5'b00110 : xpb = 1024'h10bae6ae1399b0c2537b9b2ac15ceed36fd2fe3f25c1a97bea8cdae64dade7b330de127ee9bb7f6b4301044858cbc55a6b8f4939dfcfc44c0a931fb8ca7c83eadb55bbfd936da03e5902211612f7f8e23b07e35bd539d5efb38b79a1fc295468914d0b4a64c0e3774a93572482b86a7c17484a7eada60ef3c7617b8e69984f69;
    5'b00111 : xpb = 1024'ha6bfc6e7e3247a34b53f6e3a6f37a7653658809d089af61ecfdc447ec52273d7bbbf7e2363d028c952fa6464cfbc1ee77b924c034cb21297ca3059d0c7eb507b3626073968f8b8acf75828cbead87086103803ea433349d03e17dce34153bf49260adc4ede332dd671f67b6467049c088789e5fb0d8089c4a34ea15497ee5ca9;
    5'b01000 : xpb = 1024'h8c1761cbf0c10ede4bfdc9730cb818a58b67ffca15fca24a374ef4c1899452f443586c4f13be5398c395853a634e67aa277b26e696e19097d92e548a8a87a85a1ca71dc68ef2d3d683142ddf29dd23f8f1632ae024a690a01317ae29cc5387978bc11b29a6dc7fa81299b8c55380a76ba8f1a2951d0fa76538cc4c163d62037e;
    5'b01001 : xpb = 1024'h716efcaffe5da387e2bc24abaa3889e5e0777ef7235e4e759ec1a5044e063210caf15a7ac3ac7e683430a60ff6e0b06cd36401c9e1110e97e82c4f444d24003903283453b4ecef000ed032f268e1d76bd28e51d60619d76fe8177f7057534fe5f1775a046f85d179b33cf6263ffcb2ceca595f2f2c9ec505ce49f6d7e2d5aa53;
    5'b01010 : xpb = 1024'h56c697940bfa3831797a7fe447b8fb263586fe2430bffaa1063455471278112d528a48a6739aa937a4cbc6e58a72f92f7f4cdcad2b408c97f72a49fe0fc05817e9a94ae0dae70a299a8c3805a7e68adeb3b978cbe78d1e3fbd1750b6e2531834572d98df382f234b53e033872c78be31ebc11bc93c2de2a663c7a19988495128;
    5'b01011 : xpb = 1024'h3c1e32781996ccdb1038db1ce5396c668a967d513e21a6cc6da70589d6e9f049da2336d22388d4071566e7bb1e0541f22b35b79075700a98062844b7d25caff6d02a616e00e1255326483d18e6eb3e5194e49fc1c900650f921721fd6d52e082bce3d7ba00d8751cf48370e818f4c9950d28d8634bbd0046f9454c5b2dbcf7fd;
    5'b01100 : xpb = 1024'h2175cd5c27336184a6f7365582b9dda6dfa5fc7e4b8352f7d519b5cc9b5bcf6661bc24fdd376fed686020890b1978ab4d71e9273bf9f889815263f7194f907d5b6ab77fb26db407cb204422c25eff1c4760fc6b7aa73abdf6716f343f852a8d1229a1694c981c6ee9526ae490570d4f82e9094fd5b4c1de78ec2f71cd3309ed2;
    5'b01101 : xpb = 1024'h6cd684034cff62e3db5918e203a4ee734b57bab58e4ff233c8c660f5fcdae82e9551329836529a5f69d29664529d37783076d5709cf069824243a2b57955fb49d2c8e884cd55ba63dc0473f64f4a537573aedad8be6f2af3c16c48a8352711f8850556f922b18c035c9eba9f1ece05b4ff851976adb3b882440a1de78a445a7;
    5'b01110 : xpb = 1024'h9cd2487a045abfa09f79649dce150778fb3afe093bbe4bc621dbcfa7d7423aa774367ecdfd79d30406968982bc1a2d04930a702076b154e3e3c1744355042c44f7fcd9c422607414dc164ef53cd51cdb2c6b0e3bf9e0668fc6a327cbc87cdc001d0e26740b9d631f5d2d0fe9d63911e7c039ed13cab5b659002dc7a4a6fa52e7;
    5'b01111 : xpb = 1024'h8229e35e11f7544a3637bfd66b9578b9504a7d36491ff7f1894e7fea9bb419c3fbcf6cf9ad67fdd37731aa584fac75c73ef34b03c0e0d2e3f2bf6efd17a08423de7df051485a8f3e67d254087bd9d04e0d963531db53ad5f9ba2f912537ca44e82c4654ed446b4f0fdd04d4ac2b51d4ae1a1a9adda44d3f995ab72664c6df9bc;
    5'b10000 : xpb = 1024'h67817e421f93e8f3ccf61b0f0915e9f9a559fc635681a41cf0c1302d6025f8e083685b255d5628a2e7cccb2de33ebe89eadc25e70b1050e401bd69b6da3cdc02c4ff06de6e54aa67f38e591bbade83c0eec15c27bcc6f42f70a2ca58de7c6c9ce87aa4299cf006c29e738aabaf3128ae03096647e9d3f19a2b291d27f1e1a091;
    5'b10001 : xpb = 1024'h4cd919262d307d9d63b47647a6965b39fa697b9063e350485833e0702497d7fd0b0149510d4453725867ec0376d1074c96c500ca553fcee410bb64709cd933e1ab801d6b944ec5917f4a5e2ef9e33733cfec831d9e3a3aff45a29b9f697c34eb4e30e304659958943f16c80c9bad3411247122e1f9630f3ac0a6c7e997554766;
    5'b10010 : xpb = 1024'h3230b40a3acd1246fa72d1804416cc7a4f78fabd7144fc73bfa690b2e909b719929a377cbd327e41c9030cd90a63500f42addbad9f6f4ce41fb95f2a5f758bc0920133f8ba48e0bb0b06634238e7eaa6b117aa137fad81cf1aa26ce5f47bfd39b3e721df2e42aa65dfba056d88293f7445d8df7c08f22cdb562472ab3cc8ee3b;
    5'b10011 : xpb = 1024'h17884eee4869a6f091312cb8e1973dbaa48879ea7ea6a89f271940f5ad7b96361a3325a86d20a911399e2dae9df598d1ee96b690e99ecae42eb759e42211e39f78824a85e042fbe496c2685577ec9e199242d1096120c89eefa23e2c7f7bc588199d60b9f6ebfc37805d42ce74a54ad767409c1618814a7beba21d6ce23c9510;
    5'b10100 : xpb = 1024'had8d2f2817f47062f2f4ffc88f71f64c6b0dfc48617ff5420c68aa8e24f0225aa514914ce735526f49978dcb14e5f25efe99b95a5681192fee5493fc1f80b02fd35295c1b5ce14533518700b4fcd15bd6772f197cf1a3c7f7a2ea16dc4a63068ae5b31be705e4696a7c0670e58f17c63d7823792785bc54cc78f43331092a250;
    5'b10101 : xpb = 1024'h92e4ca0c2591050c89b35b012cf2678cc01d7b756ee1a16d73db5ad0e96201772cad7f7897237d3eba32aea0a8783b21aa82943da0b0972ffd528eb5e21d080eb9d3ac4edbc82f7cc0d4751e8ed1c930489e188db08d834f4f2e72b44fa5f8b714117099390798684863a46f456d87c6f8e9f42c87eae2ed5d0cedf4b6064925;
    5'b10110 : xpb = 1024'h783c64f0332d99b62071b639ca72d8cd152cfaa27c434d98db4e0b13add3e093b4466da44711a80e2acdcf763c0a83e4566b6f20eae015300c50896fa4b95feda054c2dc01c24aa64c907a31cdd67ca329c93f839200ca1f242e43fadaa5c10579c7af7401b0ea39e906e1d031e9932a1a51b0c6977a008df28a98b65b79effa;
    5'b10111 : xpb = 1024'h5d93ffd440ca2e5fb730117267f34a0d6a3c79cf89a4f9c442c0bb567245bfb03bdf5bcff6ffd2dd9b68f04bcf9ccca702544a04350f93301b4e84296755b7cc86d5d96927bc65cfd84c7f450cdb30160af46679737410eef92e154165a58953df7dee4eca5a3c0b89aa1f311e659e8d3bb96d60a7091e2e8808437800ed96cf;
    5'b11000 : xpb = 1024'h42eb9ab84e66c3094dee6cab0573bb4dbf4bf8fc9706a5efaa336b9936b79eccc37849fba6edfdad0c041121632f1569ae3d24e77f3f11302a4c7ee329f20fab6d56eff64db680f9640884584bdfe388ec1f8d6f54e757bece2de687f0a551a245342d2993038ddd2a4d5c920ae1a9f05d2129fab6983bcf1d85ee39a6613da4;
    5'b11001 : xpb = 1024'h2843359c5c0357b2e4acc7e3a2f42c8e145b7829a468521b11a61bdbfb297de94b11382756dc287c7c9f31f6f6c15e2c5a25ffcac96e8f30394a799cec8e678a53d8068373b09c22efc4896b8ae496fbcd4ab465365a9e8ea32db7ce7ba519f0aaea6c045bacdfaecaf099f2f75db5537e88e694c627596fb30398fb4bd4e479;
    5'b11010 : xpb = 1024'hd9ad080699fec5c7b6b231c40749dce696af756b1c9fe467918cc1ebf9b5d05d2aa265306ca534bed3a52cc8a53a6ef060edaae139e0d3048487456af2abf693a591d1099aab74c7b808e7ec9e94a6eae75db5b17cde55e782d891506a4e23f10a0aadf245631806b93d753e3d9c0b69ff0a32ed5b67710488143bcf1488b4e;
    5'b11011 : xpb = 1024'ha39fb0ba392ab5cedd2ef62bee4f56602ff079b494a34ae95e6835b7370fe92a5d8b91f780defca9fd33b2e90144007c1611dd7780805b7c07e5ae6eac998bf99529684c6f35cfbb19d69634a1c9c21283a5fbe985c7593f02b9ec564bcf4d1fa55e7be39dc87bdf92f6fb93c825f24310323eab3590f1e1246e69831f9e988e;
    5'b11100 : xpb = 1024'h88f74b9e46c74a7873ed51648bcfc7a084fff8e1a204f714c5dae5f9fb81c846e524802330cd27796dced3be94d6493ec1fab85acaafd97c16e3a9286f35e3d87baa7ed9952feae4a5929b47e0ce758564d122df673aa00ed7b9bd9cd6cf156e0b14babe6671cdb1339a38f4b4a1fda63199fb4545200f81b9ec1444c5123f63;
    5'b11101 : xpb = 1024'h6e4ee6825463df220aabac9d295038e0da0f780eaf66a3402d4d963cbff3a7636cbd6e4ee0bb5248de69f494286892016de3933e14df577c25e1a3e231d23bb7622b9566bb2a060e314ea05b1fd328f845fc49d548ade6deacb98ee361ceddbc70caf9992f1b1f82d43d7655a11e09095301b7df54af2d224f69bf066a85e638;
    5'b11110 : xpb = 1024'h53a68166620073cba16a07d5c6d0aa212f1ef73bbcc84f6b94c0467f8465867ff4565c7a90a97d184f051569bbfadac419cc6e215f0ed57c34df9e9bf46e939648acabf3e1242137bd0aa56e5ed7dc6b272770cb2a212dae81b96029eccea60ad6813873f7c4715474e0b3b68d9a146c74697479643e4ac2e4e769c80ff98d0d;
    5'b11111 : xpb = 1024'h38fe1c4a6f9d08753828630e64511b61842e7668ca29fb96fc32f6c248d7659c7bef4aa64097a7e7bfa0363f4f8d2386c5b54904a93e537c43dd9955b70aeb752f2dc281071e3c6148c6aa819ddc8fde085297c10b94747e56b9317077ce6e593c37774ec06dc3261583f1177a161fcf95d1311373cd68637a651489b56d33e2;
    endcase
end

endmodule

module xpb_5_465
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h59b47ded38a9d924fbe7472efdf68b1639704bae27faf08c5c113cd655d28ad340d075df3127f415a46f2f8584194e2dfc2f91967265e9aae0f850cd82931676bbbd4a1fe30acf0111d2cfb04209120f95b40f2bdef67046f5a9e285119bc9dd65b5f798d877e89359dc90a9e8b75c89e1f50938e129d79abb023de1e5520520;
    5'b00010 : xpb = 1024'h2bbb684af657d812cc91686eb92cedb016a942b7a7e40a13a45c056f8a2689e7e586e459829699ca9801fc424d48b919444fb46c219030a1151623cca53b83c032b5f911684a0bd110b9cbdeb365fee376324bf3166b37d35c7330f690cf1289c645d080026d8992cf93a74d99e92ea7510338f720852052f9500bf41c1a3d5;
    5'b00011 : xpb = 1024'h5c703471e80f56a628b05db5e98959f13adadfd9a279312d9656fd2d4e74f371bf28e424c9515db24def4f49a8edd9bf90748cdd347eecb4f249b30a4ce6ceb2bee8a9b0f98f6fbe22de6c6e2d3f71fdcd1733eb105d23c42b7115947aa8bb06021a54a0d89ec12c86d5cb1ec255ef7457053cc85332299fea973ea12713a8f5;
    5'b00100 : xpb = 1024'h5776d095ecafb0259922d0dd7259db602d52856f4fc8142748b80adf144d13cfcb0dc8b3052d33953003f8849a917232889f68d8432061422a2c47994a770780656bf222d09417a2217397bd66cbfdc6ec6497e62cd66fa6b8e661ed219e25138c8ba10004db13259f274e9b33d25d4ea20671ee410a40a5f2a017e838347aa;
    5'b00101 : xpb = 1024'h5f2beaf69774d4275579743cd51c28cc3c4574051cf771ced09cbd8447175c103d81526a617ac74ef76f6f0dcdc2655124b98823f697efbf039b1547173a86eec21409421014107b33ea092c1875d1ec047a58aa41c3d741613848a3e3b5ac2e9e7eb1a8d8c599c5b3cf05939bf4825ecc157057c53a7ba51a2c3f6068d54cca;
    5'b00110 : xpb = 1024'h833238e0e307883865b4394c2b86c91043fbc826f7ac1e3aed14104e9e739db7b094ad0c87c3cd5fc805f4c6e7da2b4bccef1d4464b091e33f426b65efb28b409821eb3438de2373322d639c1a31fcaa6296e3d94341a77a155992e3b26d379d52d1718007489cb86ebaf5e8cdbb8bf5f309aae5618f60f8ebf023dc544eb7f;
    5'b00111 : xpb = 1024'h61e7a17b46da51a882428ac3c0aef7a73db008309775b2700ae27ddb3fb9c4aebbd9c0aff9a430eba0ef8ed1f296f0e2b8fe836ab8b0f2c914ec7783e18e3f2ac53f68d32698b13844f5a5ea03ac31da3bdd7d69732a8abe96ff7bb34cc29d573ae30eb0d8ec725ee0c84008759315494125a3e73742cdaa49c1401faa96f09f;
    5'b01000 : xpb = 1024'haeeda12bd95f604b3245a1bae4b3b6c05aa50ade9f90284e917015be289a279f961b91660a5a672a6007f1093522e465113ed1b08640c28454588f3294ee0f00cad7e445a1282f4442e72f7acd97fb8dd8c92fcc59acdf4d71ccc3da433c4a271917420009b6264b3e4e9d3667a4ba9d440ce3dc8214814be5402fd07068f54;
    5'b01001 : xpb = 1024'h64a357fff63fcf29af0ba14aac41c6823f1a9c5c11f3f31145283e32385c2d4d3a322ef591cd9a884a6fae96176b7c744d437eb17ac9f5d3263dd9c0abe1f766c86ac8643d1d51f5560142a7eee291c87340a228a4913e3bccc6aec2b5cf8e7fd7476bb8d9134af80dc17a7d4f31a833b635d776a94b1faf795640deec589474;
    5'b01010 : xpb = 1024'hdaa90976cfb7385dfed70a299de0a470714e4d964774326235cc1b2db2c0b1877ba275bf8cf100f4f809ed4b826b9d7e558e861ca7d0f325696eb2ff3a2992c0fd8ddd5709723b1553a0fb5980fdfa714efb7bbf70181720ce3ff4d0d40b5cb0df5d12800c23afde0de24484018de94495101cd3a299a19ede903bc48c83329;
    5'b01011 : xpb = 1024'h675f0e84a5a54caadbd4b7d197d4955d408530878c7233b27f6dfe8930fe95ebb88a9d3b29f70424f3efce5a3c400805e18879f83ce2f8dd378f3bfd7635afa2cb9627f553a1f2b2670cdf65da18f1b6aaa3c6e7d5f7f1b9028de1d21edc7fa873abc8c0d93a23913abab4f228d03b1e2b460b061b5371b4a8eb419e2e1a3849;
    5'b01100 : xpb = 1024'h1066471c1c60f1070cb687298570d922087f7904def583c75da28209d3ce73b6f61295a190f879abf900be98dcfb4569799de3a88c96123c67e84d6cbdf6516813043d66871bc46e6645ac7383463f954c52dc7b286834ef42ab325c764da6f3aa5a2e3000e913970dd75ebd19b7717ebe61355cac31ec1f1d7e047b8a89d6fe;
    5'b01101 : xpb = 1024'h6a1ac509550aca2c089dce588367643841efc4b306f07453b9b3bee029a0fe8a36e30b80c2206dc19d6fee1e6114939775cd753efefbfbe748e09e3a408967decec187866a26936f78187c23c54f51a4e206eba7075ea536385514e187e970d1101025c8d960fc2a67b3ef67026ece08a0563e958d5bc3b9d880425d6fdbdc1e;
    5'b01110 : xpb = 1024'h1321fda0cbc66e88397f9db07103a7fd09ea0d305973c46897e84260cc70dc55746b03e72921e348a280de5d01cfd0fb0de2deef4eaf15467939afa9884a09a4162f9cf79da0652b775149316e7c9f8383b6013a59cee86c7872656bdf5a981c46be8b38010fec303ad09931f3560469337168ec1e3a3e244d13053acc4b7ad3;
    5'b01111 : xpb = 1024'h6cd67b8e047047ad3566e4df6efa3313435a58de816eb4f4f3f97f3722436728b53b79c65a49d75e46f00de285e91f290a127085c114fef15a3200770add201ad1ece71780ab342c892418e1b085b193196a106638c558b36e1c47f0f0f661f9ac7482d0d987d4c394ad29dbdc0d60f315667224ff6415bf0815431cb19d7ff3;
    5'b10000 : xpb = 1024'h15ddb4257b2bec096648b4375c9676d80b54a15bd3f20509d22e02b7c51344f3f2c3722cc14b4ce54c00fe2126a45c8ca227da3610c818508a8b11e6529dc1e0195afc88b42505e8885ce5ef59b2ff71bb1925f98b359be9ae39987b48678944e322e8400136c4c967c9d3a6ccf49753a8819c7b904290297ca805fa0e0d1ea8;
    5'b10001 : xpb = 1024'h6f923212b3d5c52e622ffb665a8d01ee44c4ed09fbecf5962e3f3f8e1ae5cfc73393e80bf27340faf0702da6aabdaaba9e576bcc832e01fb6b8362b3d530d856d51846a8972fd4e99a2fb59f9bbc118150cd35256a2c0c30a3e37b005a03532248d8dfd8d9aead5cc1a66450b5abf3dd8a76a5b4716c67c437aa43dbf35f23c8;
    5'b10010 : xpb = 1024'h18996aaa2a91698a9311cabe482945b30cbf35874e7045ab0c73c30ebdb5ad92711be0725974b681f5811de54b78e81e366cd57cd2e11b5a9bdc74231cf17a1c1c865c19caa9a6a5996882ad44e95f5ff27c4ab8bc9c4f66e400cb8ab1747a6d7f874548015d9d6294c30e1ba6932a3e1d91d00b024ae22eac3d06b94fcec27d;
    5'b10011 : xpb = 1024'h724de897633b42af8ef911ed461fd0c9462f8135766b36376884ffe513883865b1ec56518a9caa9799f04d6acf92364c329c6713454705057cd4c4f09f849092d843a639adb475a6ab3b525d86f2716f883059e49b92bfadd9aaae0fc310444ae53d3ce0d9d585f5ee9f9ec58f4a86c7ff86d943e374b9c9673f449b3520c79d;
    5'b10100 : xpb = 1024'h1b55212ed9f6e70bbfdae14533bc148e0e29c9b2c8ee864c46b98365b6581630ef744eb7f19e201e9f013da9704d73afcab1d0c394fa1e64ad2dd65fe74532581fb1bbaae12e4762aa741f6b301fbf4e29df6f77ee0302e419c7fe9a1a816b961beba250018475fbc1bc48908031bd2892a2039a74533433dbd2077891906652;
    5'b10101 : xpb = 1024'h75099f1c12a0c030bbc2287431b29fa4479a1560f0e976d8a2cac03c0c2aa1043044c49722c6143443706d2ef466c1ddc6e1625a0760080f8e26272d69d848cedb6f05cac4391663bc46ef1b7228d15dbf937ea3ccf9732b0f71e11f2c1d357381a199e8d9fc5e8f1b98d93a68e919b274970cd3557d0bce96d4455a76e26b72;
    5'b10110 : xpb = 1024'h1e10d7b3895c648ceca3f7cc1f4ee3690f945dde436cc6ed80ff43bcaefa7ecf6dccbcfd89c789bb48815d6d9521ff415ef6cc0a5713216ebe7f389cb198ea9422dd1b3bf7b2e81fbb7fbc291b561f3c614294371f69b6614f8f31a9838e5cbeb84fff5801ab4e94eeb5830559d0501307b23729e65b86390b670837d3520a27;
    5'b10111 : xpb = 1024'h77c555a0c2063db1e88b3efb1d456e7f4904a98c6b67b779dd10809304cd09a2ae9d32dcbaef7dd0ecf08cf3193b4d6f5b265da0c9790b199f77896a342c010ade9a655bdabdb720cd528bd95d5f314bf6f6a362fe6026a84539142e952a269c1e05f6f0da233728489213af4287ac9ce9a74062c7855dd3c6694619b8a40f47;
    5'b11000 : xpb = 1024'h20cc8e3838c1e20e196d0e530ae1b24410fef209bdeb078ebb450413a79ce76dec252b4321f0f357f2017d31b9f68ad2f33bc751192c2478cfd09ad97beca2d026087acd0e3788dccc8b58e7068c7f2a98a5b8f650d069de855664b8ec9b4de754b45c6001d2272e1baebd7a336ee2fd7cc26ab95863d83e3afc08f71513adfc;
    5'b11001 : xpb = 1024'h7a810c25716bbb331554558208d83d5a4a6f3db7e5e5f81b175640e9fd6f72412cf5a1225318e76d9670acb73e0fd900ef6b58e78b920e23b0c8eba6fe7fb946e1c5c4ecf14257ddde5e28974895913a2e59c8222fc6da257b00473dfe3717c4ba6a53f8da4a0fc1758b4e241c263f875eb773f2398dafd8f5fe46d8fa65b31c;
    5'b11010 : xpb = 1024'h238844bce8275f8f463624d9f674811f126986353869482ff58ac46aa03f500c6a7d9988ba1a5cf49b819cf5decb16648780c297db452782e121fd1646405b0c2933da5e24bc2999dd96f5a4f1c2df18d008ddb582371d5bbb1d97c855a83f0ff118b96801f8ffc748a7f7ef0d0d75e7f1d29e48ca6c2a436a9109b656d551d1;
    5'b11011 : xpb = 1024'h7d3cc2aa20d138b4421d6c08f46b0c354bd9d1e3606438bc519c0140f611dadfab4e0f67eb42510a3ff0cc7b62e4649283b0542e4dab112dc21a4de3c8d37182e4f1247e07c6f89aef69c55533cbf12865bcece1612d8da2b0c77a4d674408ed56ceb100da70e85aa2848898f5c4d271d3c7a781ab9601de259347983c2756f1;
    5'b11100 : xpb = 1024'h2643fb41978cdd1072ff3b60e2074ffa13d41a60b2e788d12fd084c198e1b8aae8d607ce5243c6914501bcba039fa1f61bc5bdde9d5e2a8cf2735f53109413482c5f39ef3b40ca56eea29262dcf93f07076c0274b39dd0d8f0e4cad7beb530388d7d1670021fd86075a13263e6ac08d266e2d1d83c747c489a260a759896f5a6;
    5'b11101 : xpb = 1024'h7ff8792ed036b6356ee6828fdffddb104d44660edae2795d8be1c197eeb4437e29a67dad836bbaa6e970ec3f87b8f02417f54f750fc41437d36bb020932729bee81c840f1e4b9958007562131f0251169d2011a09294411fe68ead5cd050fa15f3330e08da97c0f3cf7dc30dcf63655c48d7db111d9e53e3552848577de8fac6;
    5'b11110 : xpb = 1024'h28ffb1c646f25a919fc851e7cd9a1ed5153eae8c2d65c9726a16451891842149672e7613ea6d302dee81dc7e28742d87b00ab9255f772d9703c4c18fdae7cb842f8a998051c56b13ffae2f20c82f9ef53ecf2733e504845626abfde727c2216129e173780246b0f9a29a6cd8c04a9bbcdbf30567ae7cce4dc9bb0b34da58997b;
    5'b11111 : xpb = 1024'h82b42fb37f9c33b69baf9916cb90a9eb4eaefa3a5560b9fec62781eee756ac1ca7feebf31b95244392f10c03ac8d7bb5ac3a4abbd1dd1741e4bd125d5d7ae1faeb47e3a034d03a151180fed10a38b104d483365fc3faf49d1c55e06c395deb3e8f976b10dabe998cfc76fd82a901f846bde80ea08fa6a5e884bd4916bfaa9e9b;
    endcase
end

endmodule

module xpb_5_50
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h942a4a443f3f298ae03c9be8bb8f952a0f4c09a3fd9be794d67f014ddadfcf80c4df7095714ac79d9bdc7d8a1fd3c9fe1bf89e517791b1bfc9375fb8706013f3cd57d17aa519ea3017354077b4caea0645fc933307f4230b2aa937ad91c263573dd4fec9a4ef6798bcb144c0a70381e27065f15deffae7e48a45feaf1994f5b;
    5'b00010 : xpb = 1024'h1285494887e7e5315c07937d1771f2a541e981347fb37cf29acfe029bb5bf9f0189bee12ae2958f3b37b8fb143fa793fc37f13ca2ef23637f926ebf70e0c027e79aafa2f54a33d4602e6a80ef6995d40c8bf926660fe8461655526f5b2384c6ae7ba9fd9349decf31796289814e0703c4e0cbe2bbdff5cfc9148bfd5e3329eb6;
    5'b00011 : xpb = 1024'h1bc7edeccbdbd7ca0a0b5d3ba32aebf7e2de41cebf8d3b6be837d03e9909f6e824e9e51c053e056d8d395789e5f7b5dfa53e9daf466b5153f5ba61f2951203bdb6807746fef4dbe90459fc1671e60be12d1f5b99917dc69217ffba708b5472a05b97efc5ceece36ca3613ce41f50a85a75131d419cff0b7ad9ed1fc0d4cbee11;
    5'b00100 : xpb = 1024'h250a92910fcfca62b80f26fa2ee3e54a83d30268ff66f9e5359fc05376b7f3e03137dc255c52b1e766f71f6287f4f27f86fe27945de46c6ff24dd7ee1c1804fcf355f45ea9467a8c05cd501ded32ba81917f24ccc1fd08c2caaa4deb647098d5cf753fb2693bd9e62f2c513029c0e0789c197c577bfeb9f922917fabc6653d6c;
    5'b00101 : xpb = 1024'h2e4d373553c3bcfb6612f0b8ba9cde9d24c7c3033f40b85e8307b0685465f0d83d85d32eb3675e6140b4e73b29f22f1f68bdb179755d878beee14de9a31e063c302b71765398192f0740a425687f6921f5deedfff27c4af37d54e1663d8cbf0b43528f9f038ad05fbaf7657c34311896c31fdb6d5afe68776b35df96b7fe8cc7;
    5'b00110 : xpb = 1024'h378fdbd997b7af941416ba774655d7efc5bc839d7f1a76d7d06fa07d3213edd049d3ca380a7c0adb1a72af13cbef6bbf4a7d3b5e8cd6a2a7eb74c3e52a24077b6d00ee8dfde9b7d208b3f82ce3cc17c25a3eb73322fb8d242fff74e116a8e540b72fdf8b9dd9c6d946c279c83ea150b4ea263a8339fe16f5b3da3f81a997dc22;
    5'b00111 : xpb = 1024'h40d2807ddbaba22cc21a8435d20ed14266b14437bef435511dd790920fc1eac85621c1416190b754f43076ec6deca85f2c3cc543a44fbdc3e80839e0b12a08baa9d66ba5a83b56750a274c345f18c662be9e8066537acf54e2aa085befc50b762b0d2f783828bd52d28d8e14491188d3112c999918fdc573fc7e9f6c9b312b7d;
    5'b01000 : xpb = 1024'h4a1525221f9f94c5701e4df45dc7ca9507a604d1fecdf3ca6b3f80a6ed6fe7c0626fb84ab8a563cecdee3ec50fe9e4ff0dfc4f28bbc8d8dfe49bafdc383009f9e6abe8bd528cf5180b9aa03bda65750322fe499983fa118595549bd6c8e131ab9eea7f64d277b3cc5e58a2605381c0f13832f8aef7fd73f24522ff578cca7ad8;
    5'b01001 : xpb = 1024'h5357c9c66393875e1e2217b2e980c3e7a89ac56c3ea7b243b8a770bbcb1de4b86ebdaf540fba1048a7ac069db1e7219eefbbd90dd341f3fbe12f25d7bf360b39238165d4fcde93bb0d0df44355b223a3875e12ccb47953b647ff2f51a1fd57e112c7cf516cc6aa45ea23b6ac5df1f90f5f3957c4d6fd22708dc75f427e63ca33;
    5'b01010 : xpb = 1024'h5c9a6e6aa78779f6cc25e1717539bd3a498f86067e8170bd060f60d0a8cbe1b07b0ba65d66cebcc28169ce7653e45e3ed17b62f2eabb0f17ddc29bd3463c0c786056e2eca730325e0e81484ad0fed243ebbddbffe4f895e6faa9c2cc7b197e1686a51f3e0715a0bf75eecaf86862312d863fb6dab5fcd0eed66bbf2d6ffd198e;
    5'b01011 : xpb = 1024'h65dd130eeb7b6c8f7a29ab3000f2b68cea8446a0be5b2f36537750e58679dea887599d66bde3693c5b27964ef5e19adeb33aecd802342a33da5611cecd420db79d2c60045181d1010ff49c524c4b80e4501da5331577d817ad5456475435a44bfa826f2aa164973901b9df4472d2694bad4615f094fc7f6d1f101f18619668e9;
    5'b01100 : xpb = 1024'h6f1fb7b32f6f5f28282d74ee8cabafdf8b79073afe34edafa0df40fa6427dba093a7947014f815b634e55e2797ded77e94fa76bd19ad454fd6e987ca54480ef6da01dd1bfbd36fa41167f059c7982f84b47d6e6645f71a485ffee9c22d51ca816e5fbf173bb38db28d84f3907d42a169d44c750673fc2deb67b47f03532fb844;
    5'b01101 : xpb = 1024'h78625c57736351c0d6313ead1864a9322c6dc7d53e0eac28ee47310f41d5d8989ff58b796c0cc2300ea3260039dc141e76ba00a23126606bd37cfdc5db4e103616d75a33a6250e4712db446142e4de2518dd379976765c7912a97d3d066df0b6e23d0f03d602842c195007dc87b2d987fb52d41c52fbdc69b058deee44c9079f;
    5'b01110 : xpb = 1024'h81a500fbb75744598435086ba41da284cd62886f7de86aa23baf21241f83d590ac438282c3216ea9e860edd8dbd950be58798a87489f7b87d01073c16254117553acd74b5076acea144e9868be318cc57d3d00cca6f59ea9c55410b7df8a16ec561a5ef070517aa5a51b1c28922311a62259333231fb8ae7f8fd3ed9366256fa;
    5'b01111 : xpb = 1024'h8ae7a59ffb4b36f23238d22a2fd69bd76e574909bdc2291b89171138fd31d288b891798c1a361b23c21eb5b17dd68d5e3a39146c601896a3cca3e9bce95a12b490825462fac84b8d15c1ec70397e3b65e19cc9ffd774e0da77fea432b8a63d21c9f7aedd0aa0711f30e630749c9349c4495f924810fb396641a19ec427fba655;
    5'b10000 : xpb = 1024'h942a4a443f3f298ae03c9be8bb8f952a0f4c09a3fd9be794d67f014ddadfcf80c4df7095714ac79d9bdc7d8a1fd3c9fe1bf89e517791b1bfc9375fb8706013f3cd57d17aa519ea3017354077b4caea0645fc933307f4230b2aa937ad91c263573dd4fec9a4ef6798bcb144c0a70381e27065f15deffae7e48a45feaf1994f5b0;
    5'b10001 : xpb = 1024'h9d6ceee883331c238e4065a747488e7cb040ca3e3d75a60e23e6f162b88dcc78d12d679ec85f7417759a4562c1d1069dfdb828368f0accdbc5cad5b3f76615330a2d4e924f6b88d318a8947f301798a6aa5c5c663873653bdd53cb286ade898cb1b24eb63f3e5e12487c590cb173ba00976c5073cefa9662d2ea5e9a0b2e450b;
    5'b10010 : xpb = 1024'ha6af938cc7270ebc3c442f65d30187cf51358ad87d4f6487714ee177963bc970dd7b5ea81f7420914f580d3b63ce433ddf77b21ba683e7f7c25e4baf7e6c16724702cba9f9bd27761a1be886ab6447470ebc259968f2a76c8ffe5ea343faafc2258f9ea2d98d548bd4476d58bbe3f21ebe72af89adfa44e11b8ebe84fcc79466;
    5'b10011 : xpb = 1024'haff238310b1b0154ea47f9245eba8121f22a4b72bd292300beb6d18c73e9c668e9c955b17688cd0b2915d51405cb7fddc1373c00bdfd0313bef1c1ab057217b183d848c1a40ec6191b8f3c8e26b0f5e7731beecc9971e99d42a8f21e1d16d5f7996cee8f73dc4b05601281a4c6542a3ce5790e9f8cf9f35f64331e6fee60e3c1;
    5'b10100 : xpb = 1024'h887977f8d20bf24cd464b0bda19332321a908dc278b41028e42084b9e951658f2cecf420376faf663755da5c46aabb33edc9dffb2c34de40ae5f84851a5a43f4c5e912a9ecf67770a688df30921e056e376be673d6afebd3fc6f39e3c08599ade42ac525d6248f1651daf11d8f43c31bda58ed31bae44ad666803565717ccb1;
    5'b10101 : xpb = 1024'h11ca3c23d114b1bd7b4a14ca65d22c75c29dc9766764ff7bdba9f8607c431350ff1cc64b5a8ba7703d33257e6667e853209c27e4ca3c690007796e43d8aba57e89340e424921061a0bdbe1fa846e8ef747d6879a6dea40edf271871915247fd0521ffc3ef7b13f6af0e8c35de364744fe4abede8faadf32baf0c634148b11c0c;
    5'b10110 : xpb = 1024'h1b0ce0c81508a456294dde88f18b25c863928a10a73ebdf52911e87559f110490b6abd54b1a053ea16f0ed57086524f3025bb1c9e1b5841c040ce43f5fb1a6bdc6098b59f372a4bd0d4f3601ffbb3d97ac3650cd9e69831ea51c1a93ee40a605c5fd4c2b920035e47cb3d7a9edd4ac6e0bb24cfed9ada1a9f7b0c32c3a4a6b67;
    5'b10111 : xpb = 1024'h244f856c58fc96eed751a8477d441f1b04874aaae7187c6e7679d88a379f0d4117b8b45e08b50063f0aeb52faa626192e41b3baef92e9f3800a05a3ae6b7a7fd02df08719dc443600ec28a097b07ec3810961a00cee8c54f57c6ae0ec75ccc3b39da9c182c4f2c5e087eebf5f844e48c32b8ac14b8ad5028405523172be3bac2;
    5'b11000 : xpb = 1024'h2d922a109cf089878555720608fd186da57c0b4526f23ae7c3e1c89f154d0a392406ab675fc9acddca6c7d084c5f9e32c5dac59410a7ba53fd33d0366dbda93c3fb485894815e2031035de10f6549ad874f5e333ff6807800a714189a078f270adb7ec04c69e22d7944a004202b51caa59bf0b2a97acfea688f983021d7d0a1d;
    5'b11001 : xpb = 1024'h36d4ceb4e0e47c2033593bc494b611c04670cbdf66cbf9611149b8b3f2fb07313054a270b6de5957a42a44e0ee5cdad2a79a4f792820d56ff9c74631f4c3aa7b7c8a02a0f26780a611a9321871a14978d955ac672fe749b0bd1bd504799518a621953bf160ed19512015148e0d2554c880c56a4076acad24d19de2ed0f165978;
    5'b11010 : xpb = 1024'h4017735924d86eb8e15d0583206f0b12e7658c79a6a5b7da5eb1a8c8d0a904293ca2997a0df305d17de80cb9905a17728959d95e3f99f08bf65abc2d7bc9abbab95f7fb89cb91f49131c861fecedf8193db5759a60668be16fc6687f52b13edb95728bddfb3c0fcaabe028da17958ce6a7cbc95655ac5ba31a4242d800afa8d3;
    5'b11011 : xpb = 1024'h495a17fd68cc61518f60cf41ac280465885a4d13e67f7653ac1998ddae57012148f090836507b24b57a5d492325754126b19634357130ba7f2ee322902cfacf9f634fcd0470abdec148fda27683aa6b9a2153ecd90e5ce122270fbfa2bcd6511094fdbca958b064437ab3d262205c504ced2286c34ac0a2162e6a2c2f248f82e;
    5'b11100 : xpb = 1024'h529cbca1acc053ea3d64990037e0fdb8294f0dae265934ccf98188f28c04fe19553e878cbc1c5ec531639c6ad45490b24cd8ed286e8c26c3ef81a82489d5ae39330a79e7f15c5c8f16032e2ee387555a06750800c1651042d51b8f7504e98b467d2d2bb72fd9fcbdc37651722c75fd22f5d8878213abb89fab8b02ade3e24789;
    5'b11101 : xpb = 1024'h5bdf6145f0b44682eb6862bec399f70aca43ce486632f34646e9790769b2fb11618c7e9613310b3f0b2164437651cd522e98770d860541dfec151e2010dbaf786fdff6ff9badfb32177682365ed403fa6ad4d133f1e4527387c622efde05b17bf10a7ba3ca28f3374f4165be36e635411cdee697f2ab671df42f6298d57b96e4;
    5'b11110 : xpb = 1024'h652205ea34a8391b996c2c7d4f52f05d6b388ee2a60cb1bf9451691c4760f8096dda759f6a45b7b8e4df2c1c184f09f2105800f29d7e5cfbe8a8941b97e1b0b7acb5741745ff99d518e9d63dda20b29acf349a67226394a43a70b66ab721d7b164e7cb906477e9b0db0c7a0a41566d5f43e545add1ab159c3cd3c283c714e63f;
    5'b11111 : xpb = 1024'h6e64aa8e789c2bb4476ff63bdb0be9b00c2d4f7ce5e67038e1b95931250ef5017a286ca8c15a6432be9cf3f4ba4c4691f2178ad7b4f77817e53c0a171ee7b1f6e98af12ef05138781a5d2a45556d613b3394639a52e2d6d4ed1b49e5903dfde6d8c51b7cfec6e02a66d78e564bc6a57d6aeba4c3b0aac41a8578226eb8ae359a;
    endcase
end

endmodule

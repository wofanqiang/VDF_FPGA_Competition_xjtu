module xpb_5_255
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'ha72da027db07fc3f5ca2e0a03df3a43c9fab8ef13520bb204985b8e8f9efbd0dab549cc8650d4bc2c119d4650fa98e5bd2168ee67b9403c151cbfc4cd7ddc023817fb59440cc831433530dac3afd2a813cd9eccdd595710f0d00ba6acf02120acc72f6b3169c3ec9db1264957a9e8e9dd963ad14860418cedaf6a01ad712da6;
    5'b00010 : xpb = 1024'h14e5b404fb60ff87eb945c1407be748793f571de26a417640930b71d1f3df7a1b56a93990ca1a97858233a8ca1f531cb7a42d1dccf7280782a397f899afbb804702ff6b288199062866a61b5875fa550279b3d99bab2ae21e1a0174d59e04241598e5ed662d387d93b624c92af53d1d3bb2c75a290c08319db5ed4035ae25b4c;
    5'b00011 : xpb = 1024'h1f588e0779117f4be15e8a1e0b9daecb5df02acd39f623160dc912abaedcf372901fdd6592f27e348434d7d2f2efcab137643acb372bc0b43f563f4e68799406a847f20bcc265893c99f92904b0f77f83b68dc66980c0532d27022f406d0636206558e41943d4bc5d91372dc06fdbabd98c2b073d920c4a6c90e3e05085388f2;
    5'b00100 : xpb = 1024'h29cb6809f6c1ff0fd728b8280f7ce90f27eae3bc4d482ec812616e3a3e7bef436ad52732194352f0b046751943ea6396f485a3b99ee500f05472ff1335f77008e05fed65103320c50cd4c36b0ebf4aa04f367b3375655c43c3402e9ab3c08482b31cbdacc5a70fb276c499255ea7a3a77658eb4521810633b6bda806b5c4b698;
    5'b00101 : xpb = 1024'h343e420c74727ed3ccf2e632135c2352f1e59cab609a3a7a16f9c9c8ce1aeb14458a70fe9f9427acdc58125f94e4fc7cb1a70ca8069e412c698fbed803754c0b1877e8be543fe8f65009f445d26f1d4863041a0052beb354b4103a4160b0a5a35fe3ed17f710d39f1475bf6eb6518c9153ef261669e147c0a46d12086335e43e;
    5'b00110 : xpb = 1024'h3eb11c0ef222fe97c2bd143c173b5d96bbe0559a73ec462c1b9225575db9e6e5203fbacb25e4fc690869afa5e5df95626ec875966e5781687eac7e9cd0f3280d508fe417984cb127933f2520961eeff076d1b8cd30180a65a4e045e80da0c6c40cab1c83287a978bb226e5b80dfb757b318560e7b241894d921c7c0a10a711e4;
    5'b00111 : xpb = 1024'h4923f6116fd37e5bb88742461b1a97da85db0e89873e51de202a80e5ed58e2b5faf50497ac35d125347b4cec36da2e482be9de84d610c1a493c93e619e71040f88a7df70dc597958d67455fb59cec2988a9f579a0d71617695b0518eba90e7e4b9724bee59e45b784fd80c0165a55e650f1b9bb8faa1cada7fcbe60bbe183f8a;
    5'b01000 : xpb = 1024'h5396d013ed83fe1fae5170501ef9d21e4fd5c7789a905d9024c2dc747cf7de86d5aa4e643286a5e1608cea3287d4c72de90b47733dca01e0a8e5fe266beee011c0bfdaca2066418a19a986d61d7e95409e6cf666eacab88786805d356781090566397b598b4e1f64ed89324abd4f474eecb1d68a43020c676d7b500d6b896d30;
    5'b01001 : xpb = 1024'h5e09aa166b347de3a41b9e5a22d90c6219d08067ade26942295b38030c96da57b05f9830b8d77a9d8c9e8778d8cf6013a62cb061a583421cbe02bdeb396cbc13f8d7d623647309bb5cdeb7b0e12e67e8b23a9533c8240f98775068dc14712a261300aac4bcb7e3518b3a589414f93038ca48115b8b624df45b2aba0f18fa9ad6;
    5'b01010 : xpb = 1024'h687c8418e8e4fda799e5cc6426b846a5e3cb3956c13474f42df393919c35d6288b14e1fd3f284f59b8b024bf29c9f8f9634e19500d3c8258d31f7db006ea981630efd17ca87fd1eca013e88ba4de3a90c6083400a57d66a968207482c1614b46bfc7da2fee21a73e28eb7edd6ca31922a7de4c2cd3c28f8148da2410c66bc87c;
    5'b01011 : xpb = 1024'h72ef5e1b66957d6b8faffa6e2a9780e9adc5f245d48680a6328bef202bd4d1f965ca2bc9c5792415e4c1c2057ac491df206f823e74f5c294e83c3d74d46874186907ccd5ec8c9a1de3491966688e0d38d9d5d2cd82d6bdba58f080296e516c676c8f099b1f8b6b2ac69ca526c44d020c857486fe1c22d10e36898e1273dcf622;
    5'b01100 : xpb = 1024'h7d62381de445fd2f857a28782e76bb2d77c0ab34e7d88c5837244aaebb73cdca407f75964bc9f8d210d35f4bcbbf2ac4dd90eb2cdcaf02d0fd58fd39a1e6501aa11fc82f3099624f267e4a412c3ddfe0eda3719a603014cb49c08bd01b418d881956390650f52f17644dcb701bf6eaf6630ac1cf6483129b2438f814214e23c8;
    5'b01101 : xpb = 1024'h87d5122061f67cf37b4456823255f57141bb6423fb2a980a3bbca63d4b12c99b1b34bf62d21acd8e3ce4fc921cb9c3aa9ab2541b4468430d1275bcfe6f642c1cd937c38874a62a8069b37b1befedb289017110673d896bdc3a909776c831aea8c61d6871825ef30401fef1b973a0d3e040a0fca0ace3542811e86215cebf516e;
    5'b01110 : xpb = 1024'h9247ec22dfa6fcb7710e848c36352fb50bb61d130e7ca3bc405501cbdab1c56bf5ea092f586ba24a68f699d86db45c9057d3bd09ac21834927927cc33ce2081f114fbee1b8b2f2b1ace8abf6b39d8531153eaf341ae2c2ed2b60a31d7521cfc972e497dcb3c8b6f09fb01802cb4abcca1e373771f54395b4ff97cc177c307f14;
    5'b01111 : xpb = 1024'h9cbac6255d577c7b66d8b2963a1469f8d5b0d60221ceaf6e44ed5d5a6a50c13cd09f52fbdebc77069508371ebeaef57614f525f813dac3853caf3c880a5fe4214967ba3afcbfbae2f01ddcd1774d57d9290c4e00f83c19fe1c30aec42211f0ea1fabc747e5327add3d613e4c22f4a5b3fbcd72433da3d741ed47361929a1acba;
    5'b10000 : xpb = 1024'ha72da027db07fc3f5ca2e0a03df3a43c9fab8ef13520bb204985b8e8f9efbd0dab549cc8650d4bc2c119d4650fa98e5bd2168ee67b9403c151cbfc4cd7ddc023817fb59440cc831433530dac3afd2a813cd9eccdd595710f0d00ba6acf02120acc72f6b3169c3ec9db1264957a9e8e9dd963ad14860418cedaf6a01ad712da60;
    5'b10001 : xpb = 1024'hf334d496ca473a876796d33178972ef83044af72fb265ad0415b21d68c0bd682c1691c2137a1f04dcd32647d4616772b1dcfeec09a73b1b6497cb36a89277445487c3ed5484e0063ee3be465d138f85ca2920226689b0f48443416c1c790994a3293f4973d0a28f203a3ffda78515e682009037e18fd2b82368f17fba1a19b;
    5'b10010 : xpb = 1024'hb660ed7147ac6fe7d31c4dd3557d172c22afd9e864d320cd4d9b6b0662b07a75d76b2e8a78876ac79decfaace40af5ce83f38dd2853b3edcb663c78380703767d60779819551631a7236cbf29810ba0707030cf03c1f22039143fbd6eb7b1b9f6f9c35fc8a6ce158fb4ca4932223a4845b643d4c6793eb86fe5f919a912cf41;
    5'b10011 : xpb = 1024'h15d8e8d9922b46c272fbf2e739370bb68c25b68d999f3dbed972123ef5ca0378382bfcb52dd94b68a5f06cf11f3b4842a560a1cb900cf429e082fc3d0584df78b57872f15d61de62ea589d99ed30de48843dcf9be11b493129e44b641ba7d2daa3c0f2cafa1092022d65f09289cc2332234c7ea60ed980455d95631b5683fce7;
    5'b10100 : xpb = 1024'h204bc2dc0fdbc68668c620f13d1645fa56206f7cacf14970de0a6dcd8568ff4912e14681b42a2024d2020a377035e12862820ab9f7c63465f59fbc01d302bb7aed906e4aa16ea6942d8dce74b0e0b0f0980b6e68be74a0421ab4570ac897f3fb508822362b7a55eecb1716dbe1760c1c00e2b9775739c1d24b44cd1d03f52a8d;
    5'b10101 : xpb = 1024'h2abe9cde8d8c464a5e904efb40f5803e201b286bc0435522e2a2c95c1507fb19ed96904e3a7af4e0fe13a77dc1307a0e1fa373a85f7f74a20abc7bc6a080977d25a869a3e57b6ec570c2ff4f74908398abd90d359bcdf7530b8462b17588151bfd4f51a15ce419db68c83d25391ff505de78f4489f9a035f38f4371eb1665833;
    5'b10110 : xpb = 1024'h353176e10b3cc60e545a7d0544d4ba81ea15e15ad39560d4e73b24eaa4a6f6eac84bda1ac0cbc99d2a2544c4122b12f3dcc4dc96c738b4de1fd93b8b6dfe737f5dc064fd298836f6b3f8302a38405640bfa6ac0279274e63fc546e582278363caa16810c8e4dddc80679636e90c9ddefbc0f2f19e7fa44ec26a3a1205ed785d9;
    5'b10111 : xpb = 1024'h3fa450e388ed45d24a24ab0f48b3f4c5b4109a49e6e76c86ebd380793445f2bba30123e7471c9e595636e20a6325abd999e645852ef1f51a34f5fb503b7c4f8195d860566d94ff27f72d6104fbf028e8d3744acf5680a574ed2479fecf68575d56ddb077bfb7a1b4a42a89b7e873c6d999a569eb305a867914530b220c48b37f;
    5'b11000 : xpb = 1024'h4a172ae6069dc5963feed9194c932f097e0b5338fa397838f06bdc07c3e4ee8c7db66db3cd6d731582487f50b42044bf5707ae7396ab35564a12bb1508fa2b83cdf05bafb1a1c7593a6291dfbf9ffb90e741e99c33d9fc85ddf485a57c58787e03a4dfe2f12165a141dbb001401dafc3773ba4bc78bac80602027523b9b9e125;
    5'b11001 : xpb = 1024'h548a04e8844e455a35b907235072694d48060c280d8b83eaf50437965383ea5d586bb78053be47d1ae5a1c97051adda514291761fe6475925f2f7ad9d678078606085708f5ae8f8a7d97c2ba834fce38fb0f886911335396cec4914c2948999eb06c0f4e228b298ddf8cd64a97c798ad54d1df8dc11b0992efb1df25672b0ecb;
    5'b11010 : xpb = 1024'h5efcdeeb01fec51e2b83352d5451a3911200c51720dd8f9cf99c9324e322e62e3321014cda0f1c8dda6bb9dd5615768ad14a8050661db5ce744c3a9ea3f5e3883e20526239bb57bbc0ccf39546ffa0e10edd2735ee8caaa7bf949cf2d638babf5d333eb953f4ed7a7d3dfc93ef71819732681a5f097b4b1fdd614927149c3c71;
    5'b11011 : xpb = 1024'h696fb8ed7faf44e2214d63375830ddd4dbfb7e06342f9b4efe34eeb372c1e1ff0dd64b19605ff14a067d5723a7100f708e6be93ecdd6f60a8968fa637173bf8a76384dbb7dc81fed040224700aaf738922aac602cbe601b8b064a8998328dbe009fa6e24855eb1671aef22dd471b6a810ffe553051db8caccb10b328c20d6a17;
    5'b11100 : xpb = 1024'h73e292effd5fc4a6171791415c101818a5f636f54781a70102cd4a420260ddcfe88b94e5e6b0c606328ef469f80aa8564b8d522d359036469e85ba283ef19b8cae504914c1d4e81e4737554ace5f4631367864cfa93f58c9a134b4403018fd00b6c19d8fb6c87553b8a049269ec5536aed9490019a3bce39b8c01d2a6f7e97bd;
    5'b11101 : xpb = 1024'h7e556cf27b10446a0ce1bf4b5fef525c6ff0efe45ad3b2b30765a5d091ffd9a0c340deb26d019ac25ea091b04905413c08aebb1b9d497682b3a279ed0c6f778ee668446e05e1b04f8a6c8625920f18d94a46039c8698afda9204bfe6dd091e216388ccfae832394056516f6ff66f3c54cb2acad2e29c0fc6a66f872c1cefc563;
    5'b11110 : xpb = 1024'h88c846f4f8c0c42e02abed5563ce8ca039eba8d36e25be650bfe015f219ed5719df6287ef3526f7e8ab22ef699ffda21c5d0240a0502b6bec8bf39b1d9ed53911e803fc749ee7880cda1b70055beeb815e13a26963f206eb82d4cb8d89f93f42104ffc66199bfd2cf40295b94e19253ea8c105a42afc5153941ef12dca60f309;
    5'b11111 : xpb = 1024'h933b20f7767143f1f8761b5f67adc6e403e661c28177ca1710965cedb13dd14278ab724b79a3443ab6c3cc3ceafa730782f18cf86cbbf6fadddbf976a76b2f9356983b208dfb40b210d6e7db196ebe2971e14136414b5dfc73a4d73436e96062bd172bd14b05c11991b3bc02a5c30e2886574075735c92e081ce5b2f77d220af;
    endcase
end

endmodule

module xpb_5_655
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h6dc33d2a02b99bcaaf111dc7ce4cca9c297c495a95c28529917158887ba99e78489c4353ad46925b4c3a606c07475009ab6c2c805e53a22241e1a542c630d301679b0097965f0ccfba594b69342d4ac257a0e3655b752abee07cccf891b74a82e0e709059e4e106200b40068a5598af164e3bcc67f2cc0304becabd4524c5c0d;
    5'b00010 : xpb = 1024'h2ad934fe438502cc931cc3b88c3f4de6e1828f84560d69dba505f7bb44508fe88df0092e9066a627f91681912b308f48f2be311a99f473f8d3240b27518f31515ae6cc807d2d1c5a6218942fcf7ed153bb3ccd322a64286d0b6d07f66943f27392c67fe18bd328367aa819f252e2efb97aed9aaaae0e23305169dca41bb651af;
    5'b00011 : xpb = 1024'h989c7228463e9e97422de1805a8c18830afed8deebcfef0536775043bffa2e60d68c4c823dad38834550e1fd3277df529e2a5d9af848161b1505b06a17c00452c281cd18138c292a1c71df9903ac1c1612ddb09785d9532bebe9d4eefafb3cf673ad88e72a2138987b5c1a5af83c7aaadfd157712d3ae3609d5688786e02adbc;
    5'b00100 : xpb = 1024'h55b269fc870a059926398771187e9bcdc3051f08ac1ad3b74a0bef7688a11fd11be0125d20cd4c4ff22d032256611e91e57c623533e8e7f1a648164ea31e62a2b5cd9900fa5a38b4c431285f9efda2a776799a6454c850da16da0fecd287e4e7258cffc317a6506cf55033e4a5c5df72f5db35555c1c4660a2d3b948376ca35e;
    5'b00101 : xpb = 1024'h12c861d0c7d56c9b0a452d61d6711f187b0b65326c65b8695da08ea9514811416133d83803ed601c9f0924477a4a5dd12cce66cf6f89b9c8378a7c332e7cc0f2a91964e9e128483f6bf071263a4f2938da15843123b74e8841ca4aeaaa148cd7d76c769f052b68416f444d6e534f443b0be513398afda960a850ea1800d69900;
    5'b00110 : xpb = 1024'h808b9efaca8f0865b9564b29a4bde9b4a487ae8d02283d92ef11e731ccf1afb9a9d01b8bb133f277eb4384b38191addad83a934fcddd5bea796c2175f4ad93f410b465817787550f2649bc8f6e7c73fb31b667967f2c7947224717e33bcbd75ab8537fa4a37978a36ff84dd6f8a8cf2c70c8d0000a2a6990f43d95ec5322f50d;
    5'b00111 : xpb = 1024'h3da196cf0b5a6f679d61f11a62b06cff5c8df4b6c273224502a686649598a129ef23e16694540644981fa5d8a57aed1a1f8c97ea097e2dc10aae875a800bf2440400316a5e556499ce09055609cdfa8c955251634e1b76f54d3752e113587f4b6a32f68090fe9077e9ec6760a63233f486d2ade4390bcc90f9bac6bc1c8ceaaf;
    5'b01000 : xpb = 1024'hab64d3f90e140b324c730ee230fd379b860a3e115835a76e9417deed11423fa237c024ba419a989fe45a0644acc23d23caf8c46a67d1cfe34c902c9d463cc5456b9b3201f4b47169886250bf3dfb454eecf334c8a990a1b42db41fd9a50fc9ce4b19ff862f4ca0d9eaa067c94b8bbee5ebb66aaab8388cc145a772906ed946bc;
    5'b01001 : xpb = 1024'h687acbcd4edf7234307eb4d2eeefbae63e10843b18808c20a7ac7e1fd9e931127d13ea9524baac6c91362769d0ab7c63124ac904a372a1b9ddd29281d19b23955ee6fdeadb8280f430219985d94ccbe0508f1e95787f9f6258a45ad77c9c71befcf976621cd1b8ae64948152f91523ae01c0488ee719efc14b24a36038433c5e;
    5'b01010 : xpb = 1024'h2590c3a18faad936148a5ac3ace23e30f616ca64d8cb70d2bb411d52a2902282c267b07007dac0393e12488ef494bba2599ccd9edf1373906f14f8665cf981e55232c9d3c250907ed7e0e24c749e5271b42b0862476e9d10839495d5542919afaed8ed3e0a56d082de889adca69e887617ca267315fb52c150a1d43001ad3200;
    5'b01011 : xpb = 1024'h935400cb92647500c39b788b7b2f08cd1f9313bf6e8df5fc4cb275db1e39c0fb0b03f3c3b52152948a4ca8fafbdc0bac0508fa1f3d6715b2b0f69da9232a54e6b9cdca6b58af9d4e923a2db5a8cb9d340bcbebc7a2e3c7cf641162cde5e064328fbff643a8a4e0e4df3c9b454bf813677cade339952812f19c8e800453f98e0d;
    5'b01100 : xpb = 1024'h5069f89fd32fdc02a7a71e7c39218c17d79959e92ed8daae6047150de6e0b26b5057b99e984166613728ca201fc54aeb4c5afeb97907e7894239038dae88b336ad1996543f7dacd939f9767c441d23c56f67d59471d2c57d8f019dcbbd6d0c23419f6d1f9629f8b95930b4cef981782f92b7c11dc40975f1a20bb0d41d6383af;
    5'b01101 : xpb = 1024'hd7ff07413fb43048bb2c46cf7140f628f9fa012ef23bf6073dbb440af87a3db95ab7f797b617a2de404eb4543ae8a2a93ad0353b4a8b95fd37b697239e71186a065623d264bbc63e1b8bf42df6eaa56d303bf6140c1c32bb9f1d8c994f9b413f37ee3fb83af108dd324ce58a70adcf7a8c19f01f2ead8f1a788e1a3e6cd7951;
    5'b01110 : xpb = 1024'h7b432d9e16b4decf3ac3e234c560d9feb91be96d84e6448a054d0cc92b314253de47c2cd28a80c89303f4bb14af5da343f192fd412fc5b82155d0eb50017e488080062d4bcaac9339c120aac139bf5192aa4a2c69c36edea9a6ea5c226b0fe96d465ed0121fd20efd3d8cec14c6467e90da55bc872179921f3758d783919d55e;
    5'b01111 : xpb = 1024'h38592572578045d11ecf882583535d4971222f974531293c18e1abfbf3d833c4239b88a80bc82055dd1b6cd66edf1973866b346e4e9d2d58a69f74998b7642d7fb4c2ebda378d8be43d15372aeed7baa8e408c936b25eb98c55ee0bffe3da687864563dd0f8238c44dcce84af9edccb123af39aca0f8fc21f8f2be480283cb00;
    5'b10000 : xpb = 1024'ha61c629c5a39e19bcde0a5ed51a027e59a9e78f1daf3ae65aa5304846f81d23c6c37cbfbb90eb2b12955cd427626697d31d760eeacf0cf7ae88119dc51a715d962e72f5539d7e58dfe2a9edbe31ac66ce5e16ff8c69b1657a5dbadb88ff4f10a672c6ce2add049264e80e8b39f4757a28892f6732025bc5244df6a1c54d0270d;
    5'b10001 : xpb = 1024'h63325a709b05489db1ec4bde0f92ab3052a4bf1b9b3e9317bde7a3b73828c3acb18b91d69c2ec67dd631ee679a0fa8bc79296588e891a15179c37fc0dd0574295632fb3e20a5f518a5e9e7a27e6c4cfe497d59c5958a1405d0cbe8b6678198fb190be3be9b5560fac875023d4cd0bc6a9e9cd4574f071f524a5c9aec1e3a1caf;
    5'b10010 : xpb = 1024'h20485244dbd0af9f95f7f1cecd852e7b0aab05455b8977c9d17c42ea00cfb51cf6df57b17f4eda4a830e0f8cbdf8e7fbc07b6a23243273280b05e5a56863d279497ec727077404a34da9306919bdd38fad194392647911b3fbbc23b43f0e40ebcaeb5a9a88da78cf42691bc6fa5a2132b4a6b23b7de882524fd9cbbbe7a41251;
    5'b10011 : xpb = 1024'h8e0b8f6ede8a4b6a45090f969bd1f91734274e9ff14bfcf362ed9b727c7953953f7b9b052c956ca5cf486ff8c54038056be796a38286154a4ce78ae82e94a57ab119c7be9dd3117308027bd24deb1e5204ba26f7bfee3c72dc38f0acd0c58b6eabd263a027288931431d1c2f9fb3ac24198a6f01fd1542829bc6779039f06e5e;
    5'b10100 : xpb = 1024'h4b2187431f55b26c2914b58759c47c61ec2d94c9b196e1a576823aa54520450584cf60e00fb580727c24911de9297744b3399b3dbe26e720de29f0ccb9f303caa46593a784a120fdafc1c498e93ca4e3685610c48edd3a2107292baaa852335f5db1da7c14ada105bd1135b94d3d10ec2f944ce62bf6a582a143a860035a6400;
    5'b10101 : xpb = 1024'h8377f176021196e0d205b7817b6ffaca433daf371e1c6578a16d9d80dc73675ca2326baf2d5943f2900b2430d12b683fa8b9fd7f9c7b8f76f6c56b14551621a97b15f906b6f308857810d5f848e2b74cbf1fa915dcc37cf321966a87fdedb500f9151580232b8da37054f42fac675b4459e2aca5ad80882a6c0d92fccc459a2;
    5'b10110 : xpb = 1024'h75fabc4162dab538bc31793fe603ca48cdb0244e07a44b811b8832608970d4ee12bf6a0ea01c269a753b12af145a068da5f7cc58581b5b19b14dfbf40b82351bff4c602801ce3d5811da58c8b8bb76372392ddf6b941628e129633a1119625d2f0785a5da080c93c37b94faba02000a5aa81e790da04c8b2f2ad85041f10b5af;
    5'b10111 : xpb = 1024'h3310b415a3a61c3aa03d1f30a3f64d9385b66a77c7ef30332f1cd1935217c65e58132fe9833c3a67221733d4384345cced49d0f293bc2cf0429061d896e0936bf2982c10e89c4ce2b999a18f540cfcc8872ec7c38830603c3d866e9ee922cdc3a257d1398e05e110b1ad69354da9656dc08bc57508e62bb2f82ab5d3e87aab51;
    5'b11000 : xpb = 1024'ha0d3f13fa65fb8054f4e3cf87243182faf32b3d25db1b55cc08e2a1bcdc164d6a0af733d3082ccc26e5194403f8a95d698b5fd72f20fcf128472071b5d11666d5a332ca87efb59b273f2ecf8883a478adecfab28e3a58afb1e033b977ada1846833eda3f2c53f172b261699df302f05f256f823b8812ebe3441761a83ac7075e;
    5'b11001 : xpb = 1024'h5de9e913e72b1f073359e2e930359b7a6738f9fc1dfc9a0ed422c94e96685646e603391813a2e08f1b2db5656373d515e008020d2db0a0e915b46cffe86fc4bd4d7ef89165c9693d1bb235bf238bce1c426b94f5b29488a948f376955266c037351e511b19d909472c558327a08c55273b79601fb6f44ee3499492780430fd00;
    5'b11010 : xpb = 1024'h1affe0e827f68609176588d9ee281ec51f3f4025de477ec0e7b768815f0f47b72b56fef2f6c2f45bc809d68a875d1455275a06a7695172bfa6f6d2e473ce230d40cac47a4c9778c7c3717e85bedd54ada6077ec28183865773e3b19329f36827e6fdc7f7075e211ba6499cb14e15b9ef51833e03e5d5b1e34f11c347cd9af2a2;
    5'b11011 : xpb = 1024'h88c31e122ab021d3c676a6a1bc74e96148bb8980740a03ea7928c109dab8e62f73f34246a40986b7144436f68ea4645ed2c63327c7a514e1e8d8782739fef60ea865c511e2f685977dcac9eef30a9f6ffda86227dcf8b11654607e8bbbaab2aac7e4d0fca5ac317da6fd9d19f36f44e0b666faca650272139afe6f1c1fe74eaf;
    5'b11100 : xpb = 1024'h45d915e66b7b88d5aa824c927a676cac00c1cfaa3454e89c8cbd603ca35fd79fb947082187299a83c120581bb28da39e1a1837c20345e6b87a1ade0bc55d545e9bb190fac9c49522258a12b58e5c260161444bf4abe7aec47f50b98993375a9b79c447d89331495220f1b6a3a0f8a9a8cc70d8ae93e3d513a07b9febe9514451;
    5'b11101 : xpb = 1024'h2ef0dbaac46efd78e8df2833859eff6b8c815d3f49fcd4ea051ff6f6c06c90ffe9acdfc6a49ae506dfc7940d676e2dd616a3c5c3ee6b88f0b5d43f050bbb2ae8efd5ce3b092a4accd495b7c29adac92c4e035c17ad6ac72aa40f4876ac4028c2ba3beb480b661269ae5d02d4e820e70e27ab692c2c53813a5f8d0bbb2bb39f3;
    5'b11110 : xpb = 1024'h70b24ae4af008ba23d9f104b06a6ba92e2445f2e8a62527831c357f7e7b0678847371150179040abba36d9acddbe32e70cd668dc9d3a5ab14d3ee93316ec85aff6985d7b46f1b17c87a2a6e55ddaf7551c811926d64bd7318abdc17ffc7b4d0f0c8ac7ba1f0471889b99d095f3db9962475e735941f1f843f1e57c9005079600;
    5'b11111 : xpb = 1024'h2dc842b8efcbf2a421aab63bc4993ddd9a4aa5584aad372a4557f72ab05758f88c8ad72afab054786712fad201a7722654286d76d8db2c87de814f17a24ae3ffe9e429642dbfc1072f61efabf92c7de6801d02f3a53ad4dfb5adfc7dd407f4ffbe6a3e960c89895d158dea1fa164fe2a5d68513d70d35b43f762ad5fce718ba2;
    endcase
end

endmodule

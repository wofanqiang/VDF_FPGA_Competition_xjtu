module xpb_5_515
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h91fa25f12e5b6d302e920a4d54fd1154afd7ed8f779d028532f9849288ca6fe91f69ab40f55c08465e9d719bfa3ebe0ae260becd1befd9972275ea4347e33e2e16c2d397ae631dcf101c9c2845f8ad20870a74714726046ddada63653f7eb363f92f87d12e00c225c9ef72ede2c7f3ebb4a94afbbda7191d4d19c81448f6a6c;
    5'b00010 : xpb = 1024'h123f44be25cb6da605d24149aa9fa22a95fafdb1eef3a050a65f309251194dfd23ed35681eab8108cbd3ae337f47d7c15c4c17d9a37dfb32e44ebd4868fc67c5c2d85a72f5cc63b9e203938508bf15a410e14e8e28e4c08dbb5b4c6ca7efd66c7f25f0fa25c01844b93dee5dbc58fe7d7695295f77b4e323a9a33902891ed4d8;
    5'b00011 : xpb = 1024'h1b5ee71d38b1247908bb61ee7fef733fe0f87c8ae66d7078f98ec8db79a5f4fbb5e3d01c2e01418d31bd854d3eebc3a20a7223c6753cf8cc56761bec9d7a9ba8a44487ac70b29596d3055d478d1ea0761951f5d53d5720d49908f2a2fbe7c1a2beb8e97738a0246715dce58c9a857dbc31dfbe0f338f54b57e74d583cdae3f44;
    5'b00100 : xpb = 1024'h247e897c4b96db4c0ba48293553f44552bf5fb63dde740a14cbe6124a2329bfa47da6ad03d57021197a75c66fe8faf82b8982fb346fbf665c89d7a90d1f8cf8b85b0b4e5eb98c773c407270a117e2b4821c29d1c51c9811b76b698d94fdfacd8fe4be1f44b803089727bdcbb78b1fcfaed2a52beef69c64753467205123da9b0;
    5'b00101 : xpb = 1024'h2d9e2bdb5e7c921f0e8da3382a8f156a76f37a3cd56110c99fedf96dcabf42f8d9d105844cacc295fd913380be339b6366be3ba018baf3ff3ac4d9350677036e671ce21f667ef950b508f0cc95ddb61a2a334463663be16254643f0fa3d7980f3ddeda715e603cabcf1ad3ea56de7c39a874e76eab4437d928180e8656cd141c;
    5'b00110 : xpb = 1024'h36bdce3a716248f21176c3dcffdee67fc1f0f915ccdae0f1f31d91b6f34be9f76bc7a0385c02831a637b0a9a7dd7874414e4478cea79f198acec37d93af5375148890f58e1652b2da60aba8f1a3d40ec32a3ebaa7aae41a93211e545f7cf83457d71d2ee714048ce2bb9cb19350afb7863bf7c1e671ea96afce9ab079b5c7e88;
    5'b00111 : xpb = 1024'h3fdd70998447ffc5145fe481d52eb7950cee77eec454b11a464d2a001bd890f5fdbe3aec6b58439ec964e1b43d7b7324c30a5379bc38ef321f13967d6f736b3429f53c925c4b5d0a970c84519e9ccbbe3b1492f18f20a1f00fbf8b7c4bc76e7bbd04cb6b842054f08858c24813377ab71f0a10ce22f91afcd1bb4788dfebe8f4;
    5'b01000 : xpb = 1024'h48fd12f8972db69817490526aa7e88aa57ebf6c7bbce8142997cc249446537f48fb4d5a07aae04232f4eb8cdfd1f5f0571305f668df7eccb913af521a3f19f170b6169cbd7318ee7880e4e1422fc569043853a38a3930236ed6d31b29fbf59b1fc97c3e897006112e4f7b976f163f9f5da54a57dded38c8ea68ce40a247b5360;
    5'b01001 : xpb = 1024'h521cb557aa136d6b1a3225cb7fce59bfa2e975a0b348516aecac5a926cf1def321ab70548a03c4a795388fe7bcc34ae61f566b535fb6ea65036253c5d86fd2f9eccd97055217c0c4791017d6a75be1624bf5e17fb805627dcb1ad7e8f3b744e83c2abc65a9e06d354196b0a5cf907934959f3a2d9aadfe207b5e808b690abdcc;
    5'b01010 : xpb = 1024'h5b3c57b6bcf9243e1d1b4670551e2ad4ede6f479aac221933fdbf2db957e85f1b3a20b089959852bfb2267017c6736c6cd7c77403175e7fe7589b26a0cee06dcce39c43eccfdf2a16a11e1992bbb6c34546688c6cc77c2c4a8c87e1f47af301e7bbdb4e2bcc079579e35a7d4adbcf87350e9cedd56886fb250301d0cad9a2838;
    5'b01011 : xpb = 1024'h645bfa15cfdedb11200467152a6dfbea38e47352a23bf1bb930b8b24be0b2cf04598a5bca8af45b0610c3e1b3c0b22a77ba2832d0334e597e7b1110e416c3abfafa5f17847e4247e5b13ab5bb01af7065cd7300de0ea230b867624559ba71b54bb50ad5fcfa08579fad49f038be977b20c34638d1262e1442501b98df22992a4;
    5'b01100 : xpb = 1024'h6d7b9c74e2c491e422ed87b9ffbdccff83e1f22b99b5c1e3e63b236de697d3eed78f4070b8050634c6f61534fbaf0e8829c88f19d4f3e33159d86fb275ea6ea291121eb1c2ca565b4c15751e347a81d86547d754f55c83526423ca8bef9f068afae3a5dce280919c577396326a15f6f0c77ef83cce3d52d5f9d3560f36b8fd10;
    5'b01101 : xpb = 1024'h769b3ed3f5aa48b725d6a85ed50d9e14cedf7104912f920c396abbb70f247aed6985db24c75ac6b92cdfec4ebb52fa68d7ee9b06a6b2e0cacbffce56aa68a285727e4beb3db088383d173ee0b8da0caa6db87e9c09cee39941d170c24396f1c13a769e59f5609dbeb4128d614842762f82c98cec8a17c467cea4f2907b48677c;
    5'b01110 : xpb = 1024'h7fbae133088fff8a28bfc903aa5d6f2a19dcefdd88a962348c9a540037b121ebfb7c75d8d6b0873d92c9c3687af6e6498614a6f37871de643e272cfadee6d66853ea7924b896ba152e1908a33d39977c762925e31e4143e01f7f16f8978edcf77a0996d70840a9e110b18490266ef56e3e14219c45f235f9a3768f11bfd7d1e8;
    5'b01111 : xpb = 1024'h88da83921b75b65d2ba8e9a87fad403f64da6eb68023325cdfc9ec49603dc8ea8d73108ce60647c1f8b39a823a9ad22a343ab2e04a30dbfdb04e8b9f13650a4b3556a65e337cebf21f1ad265c199224e7e99cd2a32b3a426fd2cbd2eeb86c82db99c8f541b20b6036d507bbf049b74acf95eb64c01cca78b78482b9304673c54;
    5'b10000 : xpb = 1024'h91fa25f12e5b6d302e920a4d54fd1154afd7ed8f779d028532f9849288ca6fe91f69ab40f55c08465e9d719bfa3ebe0ae260becd1befd9972275ea4347e33e2e16c2d397ae631dcf101c9c2845f8ad20870a74714726046ddada63653f7eb363f92f87d12e00c225c9ef72ede2c7f3ebb4a94afbbda7191d4d19c81448f6a6c0;
    5'b10001 : xpb = 1024'h9b19c85041412403317b2af22a4ce269fad56c686f16d2ad86291cdbb15716e7b16045f504b1c8cac48748b5b9e2a9eb9086cab9edaed730949d48e77c617210f82f00d129494fac011e65eaca5837f28f7b1bb85b9864b4b888099b93769e9a38c2804e40e0ce48268e6a1cc0f4732a6ff3dfab79818aaf21eb64958d86112c;
    5'b10010 : xpb = 1024'ha4396aaf5426dad634644b96ff9cb37f45d2eb416690a2d5d958b524d9e3bde64356e0a91407894f2a711fcf798695cc3eacd6a6bf6dd4ca06c4a78bb0dfa5f3d99b2e0aa42f8188f2202fad4eb7c2c497ebc2ff700ac4fb9635afd1e76e89d0785578cb53c0da6a832d614b9f20f2692b3e745b355bfc40f6bd0116d2157b98;
    5'b10011 : xpb = 1024'had590d0e670c91a9374d6c3bd4ec849490d06a1a5e0a72fe2c884d6e027064e4d54d7b5d235d49d3905af6e9392a81acecd2e293912cd26378ec062fe55dd9d6bb075b441f15b365e321f96fd3174d96a05c6a46847d254273e356083b667506b7e8714866a0e68cdfcc587a7d4d71a7e689090af1366dd2cb8e9d9816a4e604;
    5'b10100 : xpb = 1024'h5cb6a17b80413b36f31150999e20e586a57e5c2800ca2af01db2c6177fa5edb63fb9898688c8bc956e68ebc15705cc336dec69a4038ffb13a742575df099908282453ceea6ae7fdc189c08fbe9b1437b4c817f50c6958789c046a43d533bdaac873d79bc8b7fa21b5ab68ca63a9cabd52f9bed85cc5823459f0bf14d251ea05;
    5'b10101 : xpb = 1024'heeb0c76cae9ca86721a35ae6f31df6db555649b778672d7550ac4aaa08705d9f5f2334c77e24c4dbcd065d5d51448a3e504d28711f7fd4aac9b841a1387cceb09908108655119dab28b8a5242fa9f09bd38bf3c20dbb8bf79b2107a292ba8e10806d018db980644124a5ff941d649fc0e445388189ff3c62ec25b9616e15471;
    5'b10110 : xpb = 1024'h180aaed5ddcf8159750356534481b0830052e3746f0042ffa83a5cf3c913acd887e8ce0087380cd222ba3cef94b83484932ade73e3b6fae41ec2e2be480600cdeafcae41e0374bb7a38d5414c75a29dbc5a96683354e1906575fb6b07d2394174799c895ee7812666ee957282002c93ac98ee837d47a65580393f8175b70bedd;
    5'b10111 : xpb = 1024'h212a5134f0b5382c77ec76f819d181984b50624d667a1327fb69f53cf1a053d719df68b4968dcd5688a41409545c20654150ea60b575f87d90ea41627c8434b0cc68db7b5b1d7d94948f1dd74bb9b4adce1a0dca49c0794d350d5ce6d11b7f4d872cc11301581e88cb884e56fe2f487984d97ce79054d6e9d8659498a0002949;
    5'b11000 : xpb = 1024'h2a49f394039aeeff7ad5979cef2152ad964de1265df3e3504e998d861a2cfad5abd60368a5e38ddaee8deb2314000c45ef76f64d8734f6170311a006b1026893add508b4d603af718590e799d0193f7fd68ab5115e32d99412bb031d25136a83c6bfb99014382aab28274585dc5bc7b8402411974c2f487bad373119e48f93b5;
    5'b11001 : xpb = 1024'h336995f31680a5d27dbeb841c47123c2e14b5fff556db378a1c925cf42b9a1d43dcc9e1cb5394e5f5477c23cd3a3f8269d9d023a58f3f3b07538feaae5809c768f4135ee50e9e14e7692b15c5478ca51defb5c5872a539daf068a953790b55ba0652b20d271836cd84c63cb4ba8846f6fb6ea6470809ba0d8208cd9b291efe21;
    5'b11010 : xpb = 1024'h3c89385229665ca580a7d8e699c0f4d82c48ded84ce783a0f4f8be186b4648d2cfc338d0c48f0ee3ba6199569347e4074bc30e272ab2f149e7605d4f19fed05970ad6327cbd0132b67947b1ed8d85523e76c039f87179a21ce164f89cd0340f045e5aa8a39f842efe16533e398b4c635b6b93af6c3e42b9f56da6a1c6dae688d;
    5'b11011 : xpb = 1024'h45a8dab13c4c13788390f98b6f10c5ed77465db1446153c94828566193d2efd161b9d384d3e4cf68204b707052ebcfe7f9e91a13fc71eee35987bbf34e7d043c5219906146b64508589644e15d37dff5efdcaae69b89fa68abc3f5c020fb2c268578a3074cd84f123e042b1276e145747203cfa67fbe9d312bac069db23dd2f9;
    5'b11100 : xpb = 1024'h4ec87d104f31ca4b867a1a3044609702c243dc8a3bdb23f19b57eeaabc5f96cff3b06e38e33a8fec8635478a128fbbc8a80f2600ce30ec7ccbaf1a9782fb381f3385bd9ac19c76e549980ea3e1976ac7f84d522daffc5aaf89719bf674f3175cc50b9b845fb85b349aa32241550dc4b32d4e64563b990ec3007da31ef6cd3d65;
    5'b11101 : xpb = 1024'h57e81f6f6217811e89633ad519b068180d415b633354f419ee8786f3e4ec3dce85a708ecf2905070ec1f1ea3d233a7a9563531ed9fefea163dd6793bb7796c0214f1ead43c82a8c23a99d86665f6f59a00bdf974c46ebaf6671f422cc8eb0293049e940172986756f7421970333a43f1e898f905f7738054d54f3fa03b5ca7d1;
    5'b11110 : xpb = 1024'h6107c1ce74fd37f18c4c5b79ef00392d583eda3c2acec44241b71f3d0d78e4cd179da3a101e610f55208f5bd91d7938a045b3dda71aee7afaffdd7dfebf79fe4f65e180db768da9f2b9ba228ea56806c092ea0bbd8e11b3d44cce8631ce2edc944318c7e8578737953e1109f1166c330a3e38db5b34df1e6aa20dc217fec123d;
    5'b11111 : xpb = 1024'h6a27642d87e2eec48f357c1ec4500a42a33c59152248946a94e6b78636058bcba9943e55113bd179b7f2ccd7517b7f6ab28149c7436de549222536842075d3c7d7ca4547324f0c7c1c9d6beb6eb60b3e119f4802ed537b84227a8e9970dad8ff83c484fb98587f9bb08007cdef93426f5f2e22656f2863787ef278a2c47b7ca9;
    endcase
end

endmodule

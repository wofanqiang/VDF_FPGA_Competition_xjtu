module xpb_5_30
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h890b6ca87a3180bbf82fcd040c42aeb5dca5803385fbb073b1d61a0f6815cf084322f43bd04ee2cbde071bb522186bea20610dbb3e1c29148abe9b33880461dd7aa3e8c2c09f83d0e522ab66daae0e16937eeeecfc4222265e54f8719f0de227828b10b28888223c8f5b8d12b88a1b33ddd41700ce119e451e478b4c73c81bc3;
    5'b00010 : xpb = 1024'h616993fb3274ccaf255a2231082b161a47d4fd36367fc06fe5cf7ac91d28f10882fd6afed67747091caff82360d2c709dca7f390598581dd64ddf708d5364f0980f89cd6d1ae0a5cb7ab542b1c8057fc32f8e4416bfe173c071d5ee883f121bcd60e8f3b60474beb97f733467944103e6cce4f1f4bd7df59f61f9b945eadd11b;
    5'b00011 : xpb = 1024'h39c7bb4deab818a25284775e04137d7eb3047a38e703d06c19c8db82d23c1308c2d7e1c1dc9fab465b58d4919f8d222998eed96574eedaa63efd52de22683c35874d50eae2bc90e88a33fcef5e52a1e1d272d995dbba0c51afe5c55f68d4615229920dc43806759aa092d97a39fe0548fbc8873dc99e206ecdf7abdc49938673;
    5'b00100 : xpb = 1024'h1225e2a0a2fb64957faecc8afffbe4e31e33f73b9787e0684dc23c3c874f350902b25884e2c80f839a01b0ffde477d495535bf3a9058336f191caeb36f9a29618da204fef3cb17745cbca5b3a024ebc771ecceea4b76016758ae2bd64db7a0e77d158c4d0fc59f49a92e7fadfab7fa538ac2bf5c47646183a5cfbc2434793bcb;
    5'b00101 : xpb = 1024'h9b314f491d2ce55177de998f0c3e9398fad9776f1d8390dbff98564bef65041145d54cc0b316f24f7808ccb5005fe9337596ccf5ce745c83a3db49e6f79e8b3f0845edc1b46a9b4541df511a7ad2f9de056bbdd747b8238db7032447ecc5830effa09cff984dc186388a0cc0b34215876896d65d1575ffc8c4174770a841578e;
    5'b00110 : xpb = 1024'h738f769bd5703144a508eebc0826fafd6608f471ce07a0d83391b705a478261185afc383b93f568cb6b1a9233f1a445331ddb2cae9ddb54c7dfaa5bc44d0786b0e9aa1d5c57921d11467f9debca543c3a4e5b32bb77418a35fcb8abed1a8c2a453241b88700ceb354125b2f473fc0a91f7910e7b933c40dd9bef57b893270ce6;
    5'b00111 : xpb = 1024'h4bed9dee8db37d37d23343e9040f6261d13871747e8bb0d4678b17bf598b4811c58a3a46bf67bac9f55a85917dd49f72ee2498a005470e15581a01919202659714ef55e9d687a85ce6f0a2a2fe778da9445fa88027300db90893f135b68c0239a6a79a1147cc14e449c1592834b5ff9c868b469a110281f273c768007e0cc23e;
    5'b01000 : xpb = 1024'h244bc54145f6c92aff5d9915fff7c9c63c67ee772f0fc0d09b8478790e9e6a120564b109c5901f07340361ffbc8efa92aa6b7e7520b066de32395d66df3452c31b4409fde7962ee8b9794b674049d78ee3d99dd496ec02ceb15c57ac9b6f41cefa2b189a1f8b3e93525cff5bf56ff4a715857eb88ec8c3074b9f784868f27796;
    5'b01001 : xpb = 1024'had5731e9c02849e6f78d661a0c3a787c190d6eaab50b71444d5a928876b4391a4887a54595df01d3120a7db4dea7667ccacc8c305ecc8ff2bcf7f89a6738b4a095e7f2c0a835b2b99e9bf6ce1af7e5a577588cc1932e24f50fb1501e3a7d23f67cb6294ca81360cfe1b88c6eadfa0fdaf35995b95cda614c69e70394dcba9359;
    5'b01010 : xpb = 1024'h85b5593c786b95da24b7bb470822dfe0843cebad658f81408153f3422bc75b1a88621c089c07661050b35a231d61c19c871372057a35e8bb9717546fb46aa1cc9c3ca6d4b944394571249f925cca2f8b16d2821602ea1a0ab879b6951f60638bd039a7d57fd28a7eea5432a26eb404e58253cdd7daa0a26141bf13dcc7a048b1;
    5'b01011 : xpb = 1024'h5e13808f30aee1cd51e21074040b4744ef6c68b01613913cb54d53fbe0da7d1ac83c92cba22fca4d8f5c36915c1c1cbc435a57da959f41847136b045019c8ef8a2915ae8ca52bfd143ad48569e9c7970b64c776a72a60f2061421d0c0443a32123bd265e5791b42df2efd8d62f6df9f0114e05f65866e37619972424b285fe09;
    5'b01100 : xpb = 1024'h3671a7e1e8f22dc07f0c65a0fff3aea95a9be5b2c697a138e946b4b595ed9f1b0817098ea8582e8ace0512ff9ad677dbffa13dafb1089a4d4b560c1a4ece7c24a8e60efcdb61465d1635f11ae06ec35655c66cbee26204360a0a8382e926e2b67740a4e72f50dddcfb8b7f09f027eefaa0483e14d62d248af16f346c9d6bb361;
    5'b01101 : xpb = 1024'hecfcf34a13579b3ac36bacdfbdc160dc5cb62b5771bb1351d40156f4b00c11b47f18051ae8092c80cadef6dd990d2fbbbe82384cc71f316257567ef9c006950af3ac310ec6fcce8e8be99df22410d3bf5406213521df94bb2d2e9f9ce0a224bcac423700710078c0427253db0e1e4052f42763353f3659fc94744b4885168b9;
    5'b01110 : xpb = 1024'h97db3bdd1b66fa6fa46687d2081ec4c3a270e2e8fd1761a8cf162f7eb31690238b14748d7ecf7593eab50b22fba93ee5dc4931400a8e1c2ab03403232404cb2e29deabd3ad0f50b9cde14545fcef1b5288bf51004e601b721127e26b6d1804734d4f34228f9829c89382b250696bff390d168d34220503e4e78ed000fc19847c;
    5'b01111 : xpb = 1024'h7039632fd3aa4662d190dcff04072c280da05febad9b71a5030f90386829b223caeeeb5084f7d9d1295de7913a639a059890171525f774f38a535ef87136b85a30335fe7be1dd745a069ee0a3ec1653828394654be1c1087b9f048e251fb4408a0d2b2ab675753779c1e58842a25f4439c10c5529fcb44f9bf66e048e6ff39d4;
    5'b10000 : xpb = 1024'h48978a828bed9255febb322bffef938c78cfdcee5e1f81a13708f0f21d3cd4240ac962138b203e0e6806c3ff791df52554d6fcea4160cdbc6472bacdbe68a586368813fbcf2c5dd172f296ce8093af1dc7b33ba92dd8059d62b8af5936de839df45631343f167d26a4b9feb7eadfe94e2b0afd711d91860e973ef090d1e4ef2c;
    5'b10001 : xpb = 1024'h20f5b1d54430de492be58758fbd7faf0e3ff59f10ea3919d6b0251abd24ff6244aa3d8d69148a24ba6afa06db7d85045111de2bf5cca26853e9216a30b9a92b23cdcc80fe03ae45d457b3f92c265f903672d30fd9d93fab30b8115d01bc1c33347d9afbd16d5a6d5ad55a4ebab99de58ba05358f9b57c7236f1700d8bccaa484;
    5'b10010 : xpb = 1024'haa011e7dbe625f052415545d081aa9a6c0a4da24949f42111cd86bbb3a65c52c8dc6cd126197851784b6bc22d9f0bc2f317ef07a9ae64f99c950b1d6939ef48fb780b0d2a0da682e2a9deaf99d140719faac1fea99d61cd969d60e41bacfa55aca64c06f9f5dc9123cb131fe6423f98c97d94c90696965688d5e8c253092c047;
    5'b10011 : xpb = 1024'h825f45d076a5aaf8513fa98a0403110b2bd457274523520d50d1cc74ef78e72ccda143d567bfe954c35f989118ab174eedc5d64fb64fa862a3700dabe0d0e1bbbdd564e6b1e8eeb9fd2693bddee650ff9a26153f099211ef129e74b89fb2e4f01de83ef8771cf2c1454cd83224ddee9726d384aee72fa67d65369c6d1b78759f;
    5'b10100 : xpb = 1024'h5abd6d232ee8f6eb7e69feb6ffeb786f9703d429f5a7620984cb2d2ea48c092d0d7bba986de84d92020874ff5765726eaa0cbc24d1b9012b7d8f69812e02cee7c42a18fac2f77545cfaf3c8220b89ae539a00a93794e0704bb66db2f84962485716bbd814edc1c704de87e65e597e3a1b5cdbccd64f5e7923d0eacb5065e2af7;
    5'b10101 : xpb = 1024'h331b9475e72c42deab9453e3fbd3dfd40233512ca62b7205b8c48de8599f2b2d4d56315b7410b1cf40b1516d961fcd8e6653a1f9ed2259f457aec5567b34bc13ca7ecd0ed405fbd1a237e546628ae4cad919ffe7e909fc1a642f41a66979641ac4ef3c0a269b461f56842499a651d8ac44c7f4ebe2bc28a714e6bcfcf143e04f;
    5'b10110 : xpb = 1024'hb79bbc89f6f8ed1d8bea910f7bc47386d62ce2f56af8201ecbdeea20eb24d2d8d30a81e7a39160c7f5a2ddbd4da28ae229a87cf088bb2bd31ce212bc866a93fd0d38122e514825d74c08e0aa45d2eb07893f53c58c5f1300cf7a81d4e5ca3b01872ba92fe5a6fce5f1fcacd670bcdb6d3c22d0a608269bbecbecd44dc2995a7;
    5'b10111 : xpb = 1024'h9485287119a10f8dd0ee761503fef5ee4a084e62dcab32759e9408b176c81c35d0539c5a4a87f8d85d614990f6f2949842fb958a46a7dbd1bc8cbc5f506b0b1d4b7769e5a5b4062e59e339717f0b3cc70c12e429550813566b4ca08eed6a85d79afdcb4586e2920aee7b57e01f95e8eab196440b2e9408010b0658914ff1b16a;
    5'b11000 : xpb = 1024'h6ce34fc3d1e45b80fe18cb41ffe75d52b537cb658d2f4271d28d696b2bdb3e36102e131d50b05d159c0a25ff35acefb7ff427b5f6211349a96ac18349d9cf84951cc1df9b6c28cba2c6be235c0dd86acab8cd97dc4c4086c14150705d24dc56cee8149ce5ea1bbb9f716fe13e04fddf540907c29ac5a4915e2de68d93ad766c2;
    5'b11001 : xpb = 1024'h454177168a27a7742b43206efbcfc4b7206748683db3526e0686ca24e0ee6036500889e056d8c152dab3026d74674ad7bb8961347d7a8d6370cb7409eacee5755820d20dc7d11345fef48afa02afd0924b06ced2347ffd81bcdd6d7cb73105024204c8573660e568ffb2a447a109d2ffcf8ab4482a208a2abab6792125bd1c1a;
    5'b11010 : xpb = 1024'h1d9f9e69426af367586d759bf7b82c1b8b96c56aee37626a3a802ade960182368fe300a35d012590195bdedbb321a5f777d0470998e3e62c4aeacfdf3800d2a15e758621d8df99d1d17d33be44821a77ea80c426a43bf29765a5d3f39c144497958846e00e200f18084e4a7b61c3c80a5e84ec66a7e6cb3f928e896910a2d172;
    5'b11011 : xpb = 1024'ha6ab0b11bc9c7423509d42a003fadad1683c459e743312ddec5644edfe17513ed305f4df2d50085bf762fa90d53a11e1983154c4d7000f40d5a96b12c005347ed9196ee4997f1da2b69fdf251f30288e7dffb313a07e14bdc3facc653b2226bf1813579296a8315497a9d78e1a4de33e3c59036775f86984b0d614b5846aed35;
    5'b11100 : xpb = 1024'h7f09326474dfc0167dc797ccffe34235d36bc2a124b722da204fa5a7b32a733f12e06ba233786c99360bd6ff13f46d0154783a99f2696809afc8c6e80d3721aadf6e22f8aa8da42e892887e9610272741d79a868103a09d36cc332dc200566546b96d61b6e675b03a0457dc1db07d848cb533b85f3beaa9988ae24fd6f50a28d;
    5'b11101 : xpb = 1024'h576759b72d230c09aaf1ecf9fbcba99a3e9b3fa3d53b32d654490661683d953f52bae26539a0d0d674b4b36d52aec82110bf206f0dd2c0d289e822bd5a690ed6e5c2d70cbb9c2aba5bb130ada2d4bc59bcf39dbc7ff5fee9158b995304e8a5e9bf1a54a4462684b2a8e123f59bc1cd535a4d73a47184ebae608635455a3657e5;
    5'b11110 : xpb = 1024'h2fc58109e56657fcd81c4226f7b410fea9cabca685bf42d28842671b1d50b73f929559283fc93513b35d8fdb91692340cd060644293c199b64077e92a79afc02ec178b20ccaab1462e39d971e4a7063f5c6d9310efb1f3febe53ffc9e9cbe57f129dd32d1de5ae61b17cca295c7bc25de947abc2ef4b2cc3385e458d451c0d3d;
    5'b11111 : xpb = 1024'h823a85c9da9a3f005469753f39c786314fa39a9364352cebc3bc7d4d263d93fd26fcfeb45f19950f2066c49d0237e60894cec1944a572643e26da67f4cce92ef26c3f34ddb937d200c2823626795024fbe788655f6de914671c6640ceaf2514662151b5f5a4d810ba18705d1d35b7687841e3e16d116dd8103655d53001c295;
    endcase
end

endmodule

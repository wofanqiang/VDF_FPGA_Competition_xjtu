module xpb_5_295
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h91dcc77ee5eacd0250ec5554c74517fa0f3a97acf37407f8aeb9b2d28c7700d83b6b24edd9697164320e4f3c3b4a77d05e89b054a529535ac385c3d18f1284a5a12e001b2d36b953822d685fc895f290db22be54cbf516f9b7648a491505a4ecbddf59cf13163202d62336efaf44b535af20aaa143428d4232e6889cba289bcb;
    5'b00010 : xpb = 1024'h730c49a809e7653bd6d332d27e2fe8a2acff2c2911706f79df96ac4f65eb54a8738dcc62e8ac6439c4be5f319336ded658f938c3279fd669d66c4844e3529499ce0ccb87aadc7561f1c0ce1cf85020f0c24083110b6400e2b93c82976fe0a7474cb7217475636b782586870066b944420f6776603639bd541f5d9634eb6ed12b;
    5'b00011 : xpb = 1024'h543bcbd12de3fd755cba1050351ab94b4ac3c0a52f6cd6fb1073a5cc3f5fa878abb073d7f7ef570f576e6f26eb2345dc5368c131aa165978e952ccb83792a48dfaeb96f428823170615433da280a4f50a95e47cd4ad2eacbbb147ae5cabba9a1db8ee919d7b0a4ed74e9d7111e2dd34e6fae421f2930ed660bd4a3cd1cb5068b;
    5'b00100 : xpb = 1024'h356b4dfa51e095aee2a0edcdec0589f3e88855214d693e7c41509f4918d3fc48e3d31b4d073249e4ea1e7f1c430face24dd849a02c8cdc87fc39512b8bd2b48227ca6260a627ed7ed0e7999757c47db0907c0c898a41d4b4bcec73342596abfc6a66b0bf39fdde62c44d2721d5a2625acff50dde1c281d77f84bb1654dfb3beb;
    5'b00101 : xpb = 1024'h169ad02375dd2de86887cb4ba2f05a9c864ce99d6b65a5fd722d98c5f24850191bf5c2c216753cba7cce8f119afc13e84847d20eaf035f970f1fd59ee012c47654a92dcd23cda98d407aff54877eac107799d145c9b0be9dbec46b828071ae56f93e78649c4b17d813b077328d16f167303bd99d0f1f4d89e4c2befd7f41714b;
    5'b00110 : xpb = 1024'ha87797a25bc7faeab97420a06a3572969587814a5ed9adf620e74b987ebf50f15760e7afefdeae1eaedcde4dd6468bb8a6d18263542cb2f1d2a599706f25491bf5d72de8510462e0c2a867b450149ea152bc8f9a95a5d5977628f5cb95775343b71dd233af6149dae9d3ae223c5ba69cdf5c843e5261dacc17a9479a396a0d16;
    5'b00111 : xpb = 1024'h89a719cb7fc493243f5afe1e2120433f334c15c67cd6157751c445155833a4c18f838f24ff21a0f4418cee432e32f2bea1410ad1d6a33600e58c1de3c365591022b5f954ceaa1eef323bcd717fcecd0139da5456d514bf807800ee19f052559e45f599d911ae83503936fe32f3d035a93fa34ffd45590ade042055326ab04276;
    5'b01000 : xpb = 1024'h6ad69bf4a3c12b5dc541db9bd80b13e7d110aa429ad27cf882a13e9231a7f891c7a6369a0e6493c9d43cfe38861f59c49bb093405919b90ff872a25717a569044f94c4c14c4fdafda1cf332eaf88fb6120f819131483a96979d8e6684b2d57f8d4cd617e73fbbcc5889a4e43ab44c4b59fea1bbc38503aeff09762ca9bf677d6;
    5'b01001 : xpb = 1024'h4c061e1dc7bdc3974b28b9198ef5e4906ed53ebeb8cee479b37e380f0b1c4c61ffc8de0f1da7869f66ed0e2dde0bc0ca96201baedb903c1f0b5926ca6be578f87c73902dc9f5970c116298ebdf4329c10815ddcf53f293527bb0deb6a6085a5363a52923d648f63ad7fd9e5462b953c20030e77b2b476b01dd0e7062cd3cad36;
    5'b01010 : xpb = 1024'h2d35a046ebba5bd0d10f969745e0b5390c99d33ad6cb4bfae45b318be490a03237eb85842cea7974f99d1e2335f827d0908fa41d5e06bf2e1e3fab3dc02588eca9525b9a479b531a80f5fea90efd5820ef33a28b93617d3b7d88d70500e35cadf27cf0c938962fb02760ee651a2de2ce6077b33a1e3e9b13c9857dfafe82e296;
    5'b01011 : xpb = 1024'he6522700fb6f40a56f67414fccb85e1aa5e67b6f4c7b37c15382b08be04f402700e2cf93c2d6c4a8c4d2e188de48ed68aff2c8be07d423d31262fb1146598e0d6312706c5410f28f08964663eb78680d6516747d2d067247f60cf535bbe5f088154b86e9ae3692576c43e75d1a271dac0be7ef91135cb25b5fc8b932fc917f6;
    5'b01100 : xpb = 1024'ha041e9eef5a1c10ca7e2c969c4109ddbb998ff63e83bbb74c3f1dddb4a7bf4daab7951e71596ddaebe5b7d54c92f06a6e988dce085a69597f4abf382a3781d86775f2721f277c87c72b6ccc6074d7911b174259c9ec57e1e36c5599c70c403f53f34123dadf99b284ce7756580e727106fdf299a54785867e8e3142fe9f1b3c1;
    5'b01101 : xpb = 1024'h81716c18199e59462dc9a6e77afb6e84575d93e0063822f5f4ced75823f048aae39bf95c24d9d084510b8d4a211b6dace3f8654f081d18a7079277f5f7b82d7aa43df28e701d848ae24a32833707a7719891ea58de346807389d51eacb9f064fce0bd9e31046d49d9c4ac576385bb61cd025f559476f8879d55a21c81b37e921;
    5'b01110 : xpb = 1024'h62a0ee413d9af17fb3b0846531e63f2cf522285c24348a7725abd0d4fd649c7b1bbea0d1341cc359e3bb9d3f7907d4b2de67edbd8a939bb61a78fc694bf83d6ed11cbdfaedc3409951dd984066c1d5d17fafaf151da351f03a754a39267a08aa5ce3a18872940e12ebae1586efd04529306cc1183a66b88bc1d12f604c7e1e81;
    5'b01111 : xpb = 1024'h43d0706a619789b9399761e2e8d10fd592e6bcd84230f1f85688ca51d6d8f04b53e14846435fb62f766bad34d0f43bb8d8d7762c0d0a1ec52d5f80dca0384d62fdfb89676b68fca7c170fdfd967c043166cd73d15d123bd93c4d428781550b04ebbb692dd4e147883b116597a744d43590b38cd72d5de89dae483cf87dc453e1;
    5'b10000 : xpb = 1024'h24fff293859421f2bf7e3f609fbbe07e30ab5154602d59798765c3ceb04d441b8c03efbb52a2a905091bbd2a28e0a2bed346fe9a8f80a1d44046054ff4785d572ada54d3e90eb8b6310463bac63632914deb388d9c8125c23e253ad5dc300d5f7a9330d3372e80fd8a74b5a85eb96341f0fa5896205518af9abf4a90af0a8941;
    5'b10001 : xpb = 1024'h62f74bca990ba2c45651cde56a6b126ce6fe5d07e29c0fab842bd4b89c197ebc426973061e59bda9bcbcd1f80cd09c4cdb6870911f724e3532c89c348b86d4b57b9204066b474c4a097c977f5f060f13508fd49dbf00fab3ffd3324370b0fba096af878997bba72d9d805b9162df24e51412455134c48c187365828e050bea1;
    5'b10010 : xpb = 1024'h980c3c3b8f7b872e965172331debc920ddaa7d7d719dc8f366fc701e163898c3ff91bc1e3b4f0d3ecdda1c5bbc1781952c40375db720783e16b24d94d7caf1f0f8e7205b93eb2e1822c531d7be865382102bbb9ea7e526a4f761bd6d4c10b4a6c74a5247ac91ec75affb3ca8c572a7840061cef6568ed603ba1ce0c59a795a6c;
    5'b10011 : xpb = 1024'h793bbe64b3781f681c384fb0d4d699c97b6f11f98f9a307497d9699aefacec9437b463934a920014608a2c511403e89b26afbfcc3996fb4d2998d2082c0b01e525c5ebc81190ea2692589794ee4081e1f749805ae754108df939b5bba6ebb701562219ed0edf25eaff5e8cb97ce7369060a89ab549860615a693ee5dcbbf8fcc;
    5'b10100 : xpb = 1024'h5a6b408dd774b7a1a21f2d2e8bc16a721933a675ad9697f5c8b66317c92140646fd70b0859d4f2e9f33a3c466bf04fa1211f483abc0d7e5c3c7f567b804b11d952a4b7348f36a63501ebfd521dfab041de67451726c2fa76fb11ae0a01c6b95be4f9e192712c5f604ec1dcca345bc59cc0ef66743c7d3627930afbf5fd05c52c;
    5'b10101 : xpb = 1024'h3b9ac2b6fb714fdb28060aac42ac3b1ab6f83af1cb92ff76f9935c94a2959434a7f9b27d6917e5bf85ea4c3bc3dcb6a71b8ed0a93e84016b4f65daeed48b21cd7f8382a10cdc6243717f630f4db4dea1c58509d36631e45ffce9a6585ca1bbb673d1a937d37998d59e252cdaebd054a9213632332f7466397f82098e2e4bfa8c;
    5'b10110 : xpb = 1024'h1cca44e01f6de814adece829f9970bc354bccf6de98f66f82a7056117c09e804e01c59f2785ad895189a5c311bc91dad15fe5917c0fa847a624c5f6228cb31c1ac624e0d8a821e51e112c8cc7d6f0d01aca2ce8fa5a0ce48fec19ea6b77cbe1102a970dd35c6d24aed887ceba344e3b5817cfdf2226b964b6bf917265f922fec;
    5'b10111 : xpb = 1024'haea70c5f0558b516fed93d7ec0dc23bd63f7671add036ef0d92a08e40880e8dd1b877ee051c449f94aa8ab6d5713957d7488096c6623d7d525d22333b7ddb6674d904e28b7b8d7a56340312c4604ff9287c58ce47195e542b62628efcc8262fdc088caac48dd044dc3abb3db528998eb309da89365ae238d9edf9fc319bacbb7;
    5'b11000 : xpb = 1024'h8fd68e8829554d5084c01afc77c6f46601bbfb96faffd6720a070260e1f53cad53aa265561073ccedd58bb62aefffc836ef791dae89a5ae438b8a7a70c1dc65b7a6f1995355e93b3d2d396e975bf2df26ee351a0b104cf2bb7fe213e275d65584f609251ab2a3dc3130f03ec09fe27f790e4745258a5539f8b56ad5b4b010117;
    5'b11001 : xpb = 1024'h710610b14d51e58a0aa6f87a2eb1c50e9f80901318fc3df33ae3fbddbb69907d8bcccdca704a2fa47008cb5806ec638969671a496b10ddf34b9f2c1a605dd64fa74de501b3044fc24266fca6a5795c525601165cf073b914b9d6198c823867b2de3859f70d777738627253fcc172b703f12b40114b9c83b177cdbaf37c473677;
    5'b11010 : xpb = 1024'h523592da714e7dc3908dd5f7e59c95b73d45248f36f8a5746bc0f55a94dde44dc3ef753f7f8d227a02b8db4d5ed8ca8f63d6a2b7ed8761025e85b08db49de643d42cb06e30aa0bd0b1fa6263d5338ab23d1edb192fe2a2fdbbae11dadd136a0d6d10219c6fc4b0adb1d5a40d78e7461051720bd03e93b3c36444c88bad8d6bd7;
    5'b11011 : xpb = 1024'h33651503954b15fd1674b3759c87665fdb09b90b54f50cf59c9deed76e52381dfc121cb48ed0154f9568eb42b6c531955e462b266ffde411716c350108ddf638010b7bdaae4fc7df218dc82104edb912243c9fd56f518ce6bd860a2937ee6c67fbe7e941d211ea230138f41e305bd51cb1b8d78f318ae3d550bbd623ded3a137;
    5'b11100 : xpb = 1024'h1494972cb947ae369c5b90f35372370878ce4d8772f17476cd7ae85447c68bee3434c4299e1308252818fb380eb1989b58b5b394f27467208452b9745d1e062c2dea47472bf583ed91212dde34a7e7720b5a6491aec076cfbf5e027792c96ec28abfb0e7345f2398509c442ee7d0642911ffa34e248213e73d32e3bc1019d697;
    5'b11101 : xpb = 1024'ha6715eab9f327b38ed47e6481ab74f028808e53466657c6f7c349b26d43d8cc66f9fe917777c79895a274a7449fc106bb73f63e9979dba7b47d87d45ec308ad1cf184762592c3d41134e963dfd3dda02e67d22e67ab58dc976c28cc0a7cf13af489f0ab64775559b26bf7b1e9715195ec1204def67c4a12970196c58ca427262;
    5'b11110 : xpb = 1024'h87a0e0d4c32f1372732ec3c5d1a21fab25cd79b08461e3f0ad1194a3adb1e096a7c2908c86bf6c5eecd75a69a1e87771b1aeec581a143d8a5abf01b940709ac5fbf712ced6d1f94f82e1fbfb2cf80862cd9ae7a2ba2477b2789a850f02aa1609d776d25ba9c28f107622cb2f4e89a86b216719ae5abbd13b5c9079f0fb88a7c2;
    5'b11111 : xpb = 1024'h68d062fde72bababf915a143888cf053c3920e2ca25e4b71ddee8e2087263466dfe5380196025f347f876a5ef9d4de77ac1e74c69c8ac0996da5862c94b0aaba28d5de3b5477b55df27561b85cb236c2b4b8ac5ef993619b7a727d5d5d851864664e9a010c0fc885c5861b4005fe377781ade56d4db3014d490787892ccedd22;
    endcase
end

endmodule

module xpb_5_745
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h5d0800155fc50eda9580a213491ea0bdfc3ddcfc5b0d1ab6bf8bf8f992c5814b90bdf58423b12f726377f13e843e4ad50d4c5e23954fe3dd2aa64a553a982427a87deba43f2603cd5ed14e1ee608b74e62fd405282ba364a8198dcb31d5de915b802c09015d4052116452ab82c5b6a07585a089e35334a9baa6898e53e002cd0;
    5'b00010 : xpb = 1024'h962bad4fd9be8ec5ffbcc4f81e2fa2a8705b6c7e0a294f6013b389d7288558f1e336d8f7d3be0562791a336251e84dfb67e946107ecf76ea4ad554c3a5dd39ddcaca299cebb0a55ab08999b3335aa6bd1f5870c78ee3f844da5276b80912f9940fdeef67adf11b4a5ca6e9160e6ade561da325a1a1b38070e61b6c5f31df335;
    5'b00011 : xpb = 1024'h666abaea5d60f7c6f57c6e62cb019ae8834393c43bafafacc0c73197054dd6daaef16313a0ed0fc88b099474a95ccfb4c3caf2849d3cdb4bcf539fa174f5f7c5852a8e3e0de10e2309d9e7ba193e61ba34f2c75efba875cecf3e041e9def18aef900af8690b316d5bc0f99498d4217ecba343af84f4e82a2b8ca4fab311e2005;
    5'b00100 : xpb = 1024'h12c575a9fb37d1d8bff7989f03c5f4550e0b6d8fc14529ec0276713ae510ab1e3c66db1efa77c0ac4f23466c4a3d09bf6cfd28c20fd9eedd495aaa9874bba73bb95945339d7614ab56113336666b54d7a3eb0e18f1dc7f089b4a4ed701225f3281fbddecf5be23694b94dd22c1cd5bcac3b464b43436700e1cc36d8be63be66a;
    5'b00101 : xpb = 1024'h6fcd75bf5afce0b355783ab24ce495130a494a8c1c5244a2c2026a3477d62c69cd24d0a31e28f01eb29b37aace7b54947a4986e5a529d2ba7400f4edaf53cb6361d730d7dc9c1878b4e281554c740c2606e84e6b7496b5531ce32b8a1e80484839fe9e7d0b92288a61da07daee28c5d21c0e6d526969baa9c72c0671243c133a;
    5'b00110 : xpb = 1024'h1c28307ef8d3bac51ff364ee85a8ee7f95112457a1e7bee203b1a9d8579900ad5a9a48ae77b3a10276b4e9a26f5b8e9f237bbd2317c6e64bee07ffe4af197ad99605e7cd6c311f010119ccd199a0ff4375e095256acabe8ce8ef764281b38ecbc2f9cce3709d351df15f4bb422b409b0258e970e4e51a8152b252451d959d99f;
    5'b00111 : xpb = 1024'h793030945898c99fb5740701cec78f3d914f0153fcf4d998c33da2d1ea5e81f8eb583e329b64d074da2cdae0f399d97430c81b46ad16ca2918ae4a39e9b19f013e83d371ab5722ce5feb1af07fa9b691d8ddd577ed84f4d76a8852f59f1177e17afc8d7386713a3f07a4766c4f0f73b77de89fac8384f2b0d58dbd37175a066f;
    5'b01000 : xpb = 1024'h258aeb53f66fa3b17fef313e078be8aa1c16db1f828a53d804ece275ca21563c78cdb63df4ef81589e468cd8947a137ed9fa51841fb3ddba92b55530e9774e7772b28a673aec2956ac22666cccd6a9af47d61c31e3b8fe1136949dae0244be6503f7bbd9eb7c46d29729ba45839ab7958768c968686ce01c3986db17cc77ccd4;
    5'b01001 : xpb = 1024'h8292eb695634b28c156fd35150aa89681854b81bdd976e8ec478db6f5ce6d788098babc218a0b0cb01be7e1718b85e53e746afa7b503c197bd5b9f86240f729f1b30760b7a122d240af3b48bb2df60fdaad35c846673345bb82d7a611fa2a77abbfa7c6a01504bf3ad6ee4fdaff6219cdfc2d2069da02ab7e3ef73fd0a77f9a4;
    5'b01010 : xpb = 1024'h2eeda628f40b8c9ddfeafd8d896ee2d4a31c91e7632ce8ce06281b133ca9abcb970123cd722b61aec5d8300eb998985e9078e5e527a0d5293762aa7d23d522154f5f2d0109a733ac572b0008000c541b19cba33e5ca73d958439c51982d5edfe44f5aad0665b58873cf428d6e481657ae942fbc28288182347e891ddbf95c009;
    5'b01011 : xpb = 1024'h8bf5a63e53d09b78756b9fa0d28d83929f5a6ee3be3a0384c5b4140ccf6f2d1727bf195195dc91212950214d3dd6e3339dc54408bcf0b9066208f4d25e6d463cf7dd18a548cd3779b5fc4e26e6150b697cc8e390df6173e005d2a1cca033d713fcf86b607c2f5da85339538f10dccf82419d0460b7bb62bef2512ac2fd95ecd9;
    5'b01100 : xpb = 1024'h385060fdf1a7758a3fe6c9dd0b51dcff2a2248af43cf7dc4076353b0af32015ab534915cef674204ed69d344deb71d3e46f77a462f8dcc97dc0fffc95e32f5b32c0bcf9ad8623e02023399a33341fe86ebc12a4ad5957d19d1deec8503671d9785f399c6e13a6a3be2be9768456813604b1d2e1c9ca3502a564a48a3b2b3b33e;
    5'b01101 : xpb = 1024'h95586113516c8464d5676bf054707dbd266025ab9edc987ac6ef4caa41f782a645f286e11318717750e1c48362f568135443d869c4ddb07506b64a1e98cb19dad489bb3f178841cf6104e7c2194ab5d54ebe6a9d584fb3645377c93820c506ad3df65a56f70e6f5cf903c22071c37d67a37736bad1d69ac600b2e188f0b3e00e;
    5'b01110 : xpb = 1024'h41b31bd2ef435e769fe2962c8d34d729b127ff77247212ba089e8c4e21ba56e9d367feec6ca3225b14fb767b03d5a21dfd760ea7377ac40680bd55159890c95108b87234a71d4857ad3c333e6677a8f2bdb6b1574e83bc9e1f8413f083f84d30c6f188bd5c197bf0888905f9a64ec145acf76076b6be883164abff69a5d1a673;
    5'b01111 : xpb = 1024'h9ebb1be84f086d513563383fd65377e7ad65dc737f7f2d70c82a8547b47fd8356425f470905451cd787367b98813ecf30ac26ccacccaa7e3ab639f6ad328ed78b1365dd8e6434c250c0d815d4c80604120b3f1a9d13df2e8a11cf0a3a15636467ef4494d71ed81119ece30b1d2aa2b4d05516914ebf1d2cd0f14984ee3d1d343;
    5'b10000 : xpb = 1024'h4b15d6a7ecdf4762ffde627c0f17d154382db63f0514a7b009d9c4eb9442ac78f19b6c7be9df02b13c8d19b128f426fdb3f4a3083f67bb75256aaa61d2ee9ceee56514ce75d852ad5844ccd999ad535e8fac3863c771fc226d293b5c04897cca07ef77b3d6f88da52e53748b07356f2b0ed192d0d0d9c038730db62f98ef99a8;
    5'b10001 : xpb = 1024'ha81dd6bd4ca4563d955f048f58367212346b933b6021c266c965bde527082dc4825962000d903223a0050aefad3271d2c141012bd4b79f525010f4b70d86c1168de30072b4fe567ab7161af87fb60aacf2a978b64a2c326ceec2180f21e765dfbff23843eccc92c644989f433390d932672b9b6f060d0ad41d764f14d6efc678;
    5'b10010 : xpb = 1024'h5478917cea7b304f5fda2ecb90facb7ebf336d06e5b73ca60b14fd8906cb02080fceda0b671ae307641ebce74e12abdd6a7337694754b2e3ca17ffae0d4c708cc211b76844935d03034d6674cce2fdca61a1bf7040603ba6bace62c7851aac6348ed66aa51d79f59d41de31c681c1d1070abc52aeaf4f83f816f6cf58c0d8cdd;
    5'b10011 : xpb = 1024'hd34c3c88520a612a555907c9bf24eb49fb46d26b4cb6e54cc43d2ce68dd64b9d445216c0a593eb28386edeeef2e5e813a56da6b9f1c675441f0aa50d122002f6406e5dd428638b4f84b1f11a0ff0e7d09a062a369444e086daad7fe84df2e6d1e89510b6e2abed63a326f59ca760ee7a2beee6cfdce5aae5688ad6412b5342;
    5'b10100 : xpb = 1024'h5ddb4c51e817193bbfd5fb1b12ddc5a9463923cec659d19c0c503626795357972e02479ae456c35d8bb0601d733130bd20f1cbca4f41aa526ec554fa47aa442a9ebe5a02134e6758ae5600100018a8363397467cb94e7b2b08738a3305abdbfc89eb55a0ccb6b10e79e851adc902caf5d285f785051030468fd123bb7f2b8012;
    5'b10101 : xpb = 1024'ha36071185edf34d8a5125574ba21f15d100fd9a4bef4bdb4dff75ca59162bdabb77bfa63de174414fca121514116ac7ca240207c1debde3e8cc5ff1476ff3a0d2ed10f7a2e36de0fa8d4b8c4d459b53a28f8d36af828464d47fd4eb68df228012e6840731c1bda2096d9586fd8e0ed3dc062140e9f81db1f3ca419c34494677;
    5'b10110 : xpb = 1024'h673e0726e5b302281fd1c76a94c0bfd3cd3eda96a6fc66920d8b6ec3ebdbad264c35b52a6192a3b3b3420353984fb59cd770602b572ea1c11372aa46820817c87b6afc9be20971ae595e99ab334e52a2058ccd89323cbaaf5618b19e863d0b95cae944974795c2c31fb2c03f29e978db346029df1f2b684d9e32da8172497347;
    5'b10111 : xpb = 1024'h1398c1e68389dc39ea4cf1a6cd8519405806b4622c91e0d14f3aae67cb9e8169d9ab2d35bb1d5497775bb54b392fefa780a29668c9cbb5528d79b53d81cdc73eaf99b391719e7836a595e527807b45bf748514432870c3e92224fc56e970521953e472fdaca0cf56af3804185e74bcb93de0539b041355b9022bf862276739ac;
    5'b11000 : xpb = 1024'h70a0c1fbe34eeb147fcd93ba16a3b9fe5444915e879efb880ec6a7615e6402b56a6922b9dece8409dad3a689bd6e3a7c8deef48c5f1b992fb81fff92bc65eb6658179f35b0c47c04046733466683fd0dd7825495ab2afa33a3bdd90a06ce3b2f0be7338dc274d477c57d2ed08ad026c0963a5c393946a054ac9491476567667c;
    5'b11001 : xpb = 1024'h1cfb7cbb8125c5264a48bdf64f68136adf0c6b2a0d3475c75075e7053e26d6f8f7de9ac5385934ed9eed58815e4e748737212ac9d1b8acc132270a89bc2b9adc8c46562b4059828c509e7ec2b3b0f02b467a9b4fa15f036d6fca23c26a0181b294e261f4277fe10b550272a9bf5b6a9e9fba85f51e2e8dc0108daf281a852ce1;
    5'b11010 : xpb = 1024'h7a037cd0e0ead400dfc960099886b428db4a48266841907e1001dffed0ec5844889c90495c0a6460026549bfe28cbf5c446d88ed6708909e5ccd54def6c3bf0434c441cf7f7f8659af6fcce199b9a779a977dba2241939b7f1630075875f6ac84ce522843d53e62c6b479d61ebb6d4a5f8148e935361d85bbaf6480d588559b1;
    5'b11011 : xpb = 1024'h265e37907ec1ae12aa448a45d14b0d95661221f1edd70abd51b11fa2b0af2c8816120854b5951543c67efbb7836cf966ed9fbf2ad9a5a42fd6d45fd5f6896e7a68f2f8c50f148ce1fba7185de6e69a971870225c1a4d42f1bd6f4b2dea92b14bd5e050eaa25ef2bffacce13b204218840194b84f3849c5c71eef65ee0da32016;
    5'b11100 : xpb = 1024'h836637a5de86bced3fc52c591a69ae53624ffeee48e42574113d189c4374add3a6cffdd8d94644b629f6ecf607ab443bfaec1d4e6ef5880d017aaa2b312192a21170e4694e3a90af5a78667cccef51e57b6d62ae9d07793c3f0827e107f09a618de3117ab832f7e111120bf34c9d828b59eec0ed6d7d1062c957fed34ba34ce6;
    5'b11101 : xpb = 1024'h2fc0f2657c5d96ff0a405695532e07bfed17d8b9ce799fb352ec584023378217344575e432d0f599ee109eeda88b7e46a41e538be1929b9e7b81b52230e74218459f9b5eddcf9737a6afb1f91a1c4502ea65a968933b82760b1472996b23e0e516de3fe11d3e0474a0974fcc8128c669636eeaa95264fdce2d511cb400c1134b;
    5'b11110 : xpb = 1024'h8cc8f27adc22a5d99fc0f8a89c4ca87de955b5b62986ba6a12785139b5fd0362c5036b685682250c5188902c2cc9c91bb16ab1af76e27f7ba627ff776b7f663fee1d87031cf59b05058100180024fc514d62e9bb15f5b8c08cad4f4c8881c9facee1007133120995b6dc7a84ad843070bbc8f34787984869d7b9b5993ec1401b;
    5'b11111 : xpb = 1024'h3923ad3a79f97feb6a3c22e4d51101ea741d8f81af1c34a9542790dd95bfd7a65278e373b00cd5f015a24223cdaa03265a9ce7ece97f930d202f0a6e6b4515b6224c3df8ac8aa18d51b84b944d51ef6ebc5b30750c29c1fa58b99a04ebb5107e57dc2ed7981d16294661be5de20f744ec5491d036c8035d53bb2d379f3df0680;
    endcase
end

endmodule

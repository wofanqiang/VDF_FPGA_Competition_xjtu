module xpb_5_165
(
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(*) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'hb397c9d512f82c740f84d88ffec96b27f12115d2577c729331eb028c1558ea606e1e815c9b22cdd38ac4810272f2ccd999dbfe1f4f4204a783cb372e31c442de817fabccb4dae1e07ebf5db835bbd96ae8c58dd2898a91a4fe7ee0356fc71e4b7f7d0fde4cab1d2d61a22b8ad96263143b63f363011dc91b03b322ca836c269;
    5'b00010 : xpb = 1024'h1672f93aa25f058e81f09b11ffd92d64fe2422ba4aef8e52663d605182ab1d4c0dc3d02b936459ba715890204e5e599b333b7fc3e9e84094f07966e5c638885bd02ff579969b5c3c0fd7ebb706b77b2d5d18b1ba513152349fcfdc06adf8e3c96fefa1fbc99563a5ac3445715b2c4c62876c7e6c6023b92360766459506d84d2;
    5'b00011 : xpb = 1024'h21ac75d7f38e8855c2e8e89affc5c4177d3634177067557b995c107a4400abf214a5b8415d168697aa04d830758d8668ccd93fa5dedc60df68b61a58a954cc89b847f03661e90a5a17c3e1928a1338c40ba50a9779c9fb4eefb7ca0a04f555ae27e772f9ae601578824e682a08c27293cb22bda2903595b510b19685f8a4473b;
    5'b00100 : xpb = 1024'h2ce5f27544be0b1d03e13623ffb25ac9fc48457495df1ca4cc7ac0a305563a981b87a05726c8b374e2b120409cbcb3366676ff87d3d08129e0f2cdcb8c7110b7a05feaf32d36b8781fafd76e0d6ef65aba316374a262a4693f9fb80d5bf1c792dfdf43f7932ac74b58688ae2b65898c50ed8fcd8c0477246c0ecc8b2a0db09a4;
    5'b00101 : xpb = 1024'h381f6f1295ed8de444d983acff9ef17c7b5a56d1bb56e3cdff9970cbc6abc93e2269886cf07ae0521b5d6850c3ebe0040014bf69c8c4a174592f813e6f8d54e58877e5aff8846696279bcd4990cab3f168bdbc51cafb4d838f87a610b2ee397797d714f577f5791e2e82ad9b63eebef6528f3c0ef0594ed87127fadf4911cc0d;
    5'b00110 : xpb = 1024'h4358ebafe71d10ab85d1d135ff8b882efa6c682ee0ceaaf732b820f4880157e4294b7082ba2d0d2f5409b060eb1b0cd199b27f4bbdb8c1bed16c34b152a99913708fe06cc3d214b42f87c32514267188174a152ef393f69ddf6f941409eaab5c4fcee5f35cc02af1049cd0541184e52796457b45206b2b6a21632d0bf1488e76;
    5'b00111 : xpb = 1024'h4e92684d384c9372c6ca1ebeff781ee1797e798c0646722065d6d11d4956e68a302d589883df3a0c8cb5f871124a399f33503f2db2ace20949a8e82435c5dd4158a7db298f1fc2d23773b90097822f1ec5d66e0c1c2c9fb82f57821760e71d4107c6b6f1418adcc3dab6f30cbf1b0b58d9fbba7b507d07fbd19e5f38997f50df;
    5'b01000 : xpb = 1024'h59cbe4ea897c163a07c26c47ff64b593f8908ae92bbe394998f581460aac7530370f40ae4d9166e9c56240813979666cccedff0fa7a10253c1e59b9718e2216f40bfd5e65a6d70f03f5faedc1addecb57462c6e944c548d27f3f701ab7e38f25bfbe87ef26558e96b0d115c56cb1318a1db1f9b1808ee48d81d9916541b61348;
    5'b01001 : xpb = 1024'h65056187daab990148bab9d0ff514c4677a29c4651360072cc14316ecc0203d63df128c4174393c6fe0e889160a8933a668bbef19c95229e3a224f09fbfe659d28d7d0a325bb1f0e474ba4b79e39aa4c22ef1fc66d5df1eccf275e1e0ee0010a77b658ed0b20406986eb387e1a4757bb616838e7b0a0c11f3214c391e9ecd5b1;
    5'b01010 : xpb = 1024'h703ede252bdb1bc889b30759ff3de2f8f6b4ada376adc79bff32e1978d57927c44d310d9e0f5c0a436bad0a187d7c00800297ed3918942e8b25f027cdf1aa9cb10efcb5ff108cd2c4f379a93219567e2d17b78a395f69b071f0f4c2165dc72ef2fae29eaefeaf23c5d055b36c7dd7deca51e781de0b29db0e24ff5be9223981a;
    5'b01011 : xpb = 1024'h7b785ac27d0a9e8fcaab54e2ff2a79ab75c6bf009c258ec5325191c04ead21224bb4f8efaaa7ed816f6718b1af06ecd599c73eb5867d63332a9bb5efc236edf8f907c61cbc567b4a5723906ea4f125798007d180be8f44216ef73a24bcd8e4d3e7a5fae8d4b5a40f331f7def7573a41de8d4b75410c47a42928b27eb3a5a5a83;
    5'b01100 : xpb = 1024'h86b1d75fce3a21570ba3a26bff17105df4d8d05dc19d55ee657041e91002afc85296e105745a1a5ea81360c1d63619a33364fe977b71837da2d86962a5533226e11fc0d987a429685f0f864a284ce3102e942a5de727ed3bbedf282813d556b89f9dcbe6b98055e20939a0a82309ca4f2c8af68a40d656d442c65a17e2911cec;
    5'b01101 : xpb = 1024'h91eb53fd1f69a41e4c9beff4ff03a71073eae1bae7151d17988ef211d1583e6e5978c91b3e0c473be0bfa8d1fd654670cd02be797065a3c81b151cd5886f7654c937bb9652f1d78666fb7c25aba8a0a6dd20833b0fc096560ec7162b6ad1c89d57959ce49e4b07b4df53c360d09ff080704135c070e83365f3018c448ac7df55;
    5'b01110 : xpb = 1024'h9d24d09a709926e58d943d7dfef03dc2f2fcf3180c8ce440cbada23a92adcd14605ab13107be7419196bf0e22494733e66a07e5b6559c4129351d0486b8bba82b14fb6531e3f85a46ee772012f045e3d8bacdc1838593f705eaf042ec1ce3a820f8d6de28315b987b56de6197e3616b1b3f774f6a0fa0ff7a33cbe7132fea1be;
    5'b01111 : xpb = 1024'ha85e4d37c1c8a9acce8c8b06fedcd475720f04753204ab69fecc526354035bba673c9946d170a0f6521838f24bc3a00c003e3e3d5a4de45d0b8e83bb4ea7feb09967b10fe98d33c276d367dcb2601bd43a3934f560f1e88aae96f23218caac66c7853ee067e06b5a8b8808d22bcc3ce2f7adb42cd10bec895377f09ddb356427;
    5'b10000 : xpb = 1024'h2ea847f5109f7ab447f60b8ee6f23d67fab12a18204d21bb40e493662563d586ad603e3d0fc4f44eb6641bb8f94bc0f35c1d6392c8f345bd32bf7cff6f1ce2d0d30771e0549e49b6c255b159ce01539f4c09439fd04649448f24e3ab59c7bb950757db49be2249fdae244abe1923ceaec8a1480b0d26beabd43a7c5fa89c025;
    5'b10001 : xpb = 1024'he24011ca2397a728577ae41ee5bba88febd23fea77c9944e72cf95f23abcbfe71b7ebf99aae7c22241289cbb6c3e8dccf5f961b218354a64b68ab42da0e125af54871dad09792b9741150f1203bd2d0a34ced17259d0dae98da3c3e0c98ed9e086d4eb280acd672b0fc67648f28631c304053b6e0e4487c6d7ed9f2a2c0828e;
    5'b10010 : xpb = 1024'h195d7db9f368fd39c66ffbcaee48513b7dcf355bccf4606e1a4ba987e5015aa47899d40f6460a8ff5cbed1dbddf315aa68fd55fd167774f0c3a55eb5bd2a5688dd606c979be540d77bfd46cca397906751d945f44e35b6c8e8c22a4163955f82c0651fb06577884587168a1d3cbe894d73f692ed10f6250e1dba0c1f4af744f7;
    5'b10011 : xpb = 1024'h2496fa574498800107684953ee34e7edfce146b8f26c27974d6a59b0a656e94a7f7bbc252e12d5dc956b19ec05224278029b15df0b6b953b3be21228a0469ab6c57867546732eef583e93ca826f34dfe00659ed176ce5fe338aa1844ba91d167785cf0ae4a423a185d30acd5ea54af7eb7acd2234108019fcdf53e4bf32e0760;
    5'b10100 : xpb = 1024'h2fd076f495c802c8486096dcee217ea07bf3581617e3eec0808909d967ac77f0865da43af7c502b9ce1761fc2c516f459c38d5c1005fb585b41ec59b8362dee4ad90621132809d138bd53283aa4f0b94aef1f7ae9f6708fd88920648118e434c3054c1ac2f0cebeb334acf8e97ead5affb6311597119de317e3070789b64c9c9;
    5'b10101 : xpb = 1024'h3b09f391e6f7858f8958e465ee0e1552fb0569733d5bb5e9b3a7ba02290206968d3f8c50c1772f9706c3aa0c53809c1335d695a2f553d5d02c5b790e667f231295a85ccdfdce4b3193c1285f2daac92b5d7e508bc7ffb217d879f44b688ab530e84c92aa13d79dbe0964f2474580fbe13f19508fa12bbac32e6ba2a5439b8c32;
    5'b10110 : xpb = 1024'h4643702f38270856ca5131eeedfaac057a177ad062d37d12e6c66a2aea57953c942174668b295c743f6ff21c7aafc8e0cf745584ea47f61aa4982c81499b67407dc0578ac91bf94f9bad1e3ab10686c20c0aa968f0985b322861e24ebf872715a04463a7f8a24f90df7f14fff317221282cf8fc5d13d9754dea6d4d1ebd24e9b;
    5'b10111 : xpb = 1024'h517ceccc89568b1e0b497f77ede742b7f9298c2d884b443c19e51a53abad23e29b035c7c54db8951781c3a2ca1def5ae69121566df3c16651cd4dff42cb7ab6e65d852479469a76da399141634624458ba9702461931044c7849d052168398fa583c34a5dd6d0163b59937b8a0ad4843c685cefc014f73e68ee206fe94091104;
    5'b11000 : xpb = 1024'h5cb66969da860de54c41cd00edd3d96a783b9d8aadc30b654d03ca7c6d02b288a1e544921e8db62eb0c8823cc90e227c02afd548d43036af951193670fd3ef9c4df04d045fb7558bab8509f1b7be01ef69235b2341c9ad66c831be556d800adf103405a3c237b3368bb35a714e436e750a3c0e32316150783f1d392b3c3fd36d;
    5'b11001 : xpb = 1024'h67efe6072bb590ac8d3a1a89edc0701cf74daee7d33ad28e80227aa52e58412ea8c72ca7e83fe30be974ca4cf03d4f499c4d952ac92456fa0d4e46d9f2f033ca360847c12b0503a9b370ffcd3b19bf8617afb4006a6256811819ac58c47c7cc3c82bd6a1a702650961cd7d29fbd994a64df24d6861732d09ef586b57e47695d6;
    5'b11010 : xpb = 1024'h732962a47ce51373ce326812edad06cf765fc044f8b299b7b3412acdefadcfd4afa914bdb1f20fe92221125d176c7c1735eb550cbe187744858afa4cd60c77f81e20427df652b1c7bb5cf5a8be757d1cc63c0cdd92faff9b68019a5c1b78eea88023a79f8bcd16dc37e79fe2a96fbad791a88c9e9185099b9f939d848cad583f;
    5'b11011 : xpb = 1024'h7e62df41ce14963b0f2ab59bed999d81f571d1a21e2a60e0e65fdaf6b1035e7ab68afcd37ba43cc65acd5a6d3e9ba8e4cf8914eeb30c978efdc7adbfb928bc2606383d3ac1a05fe5c348eb8441d13ab374c865babb93a8b5b7e9885f7275608d381b789d7097c8af0e01c29b5705e108d55ecbd4c196e62d4fcecfb134e41aa8;
    5'b11100 : xpb = 1024'h899c5bdf1f44190250230324ed8634347483e2ff43a2280a197e8b1f7258ed20bd6ce4e9455669a39379a27d65cad5b26926d4d0a800b7d9760461329c450053ee5037f78cee0e03cb34e15fc52cf84a2354be97e42c51d007d17662c971d271f013499b55627a81e41be554049c073a19150b0af1a8c2bf000a01dddd1add11;
    5'b11101 : xpb = 1024'h94d5d87c70739bc9911b50aded72cae6f395f45c6919ef334c9d3b4833ae7bc6c44eccff0f089680cc25ea8d8cfa028002c494b29cf4d823ee4114a57f614481d66832b4583bbc21d320d73b4888b5e0d1e117750cc4faea57b96466206e4456a80b1a993a2d2c54ba36080cb2322d6b5ccb4a4121ba9f50b045340a85519f7a;
    5'b11110 : xpb = 1024'ha00f5519c1a31e90d2139e36ed5f619972a805b98e91b65c7fbbeb70f5040a6ccb30b514d8bac35e04d2329db4292f4d9c62549491e8f86e667dc818627d88afbe802d7123896a3fdb0ccd16cbe47377806d7052355da404a7a15269776ab63b6002eb971ef7de2790502ac55fc8539ca081897751cc7be2608066372d8861e3;
    5'b11111 : xpb = 1024'hab48d1b712d2a158130bebbfed4bf84bf1ba1716b4097d85b2da9b99b6599912d2129d2aa26cf03b3d7e7aaddb585c1b3600147686dd18b8deba7b8b4599ccdda698282deed7185de2f8c2f24f40310e2ef9c92f5df64d1ef789406cce67282017fabc9503c28ffa666a4d7e0d5e79cde437c8ad81de587410bb9863d5bf244c;
    endcase
end

endmodule

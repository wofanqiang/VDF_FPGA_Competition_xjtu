module xpb_5_885
(
    input clk, 
    input [5:1] data_in, 
    output [1024:1] data_out 
); 

reg [1024:1] xpb; 

assign data_out = xpb; 

always@(posedge clk) begin
    case(data_in)
    5'b00000 : xpb = 1024'h0;
    5'b00001 : xpb = 1024'h6192805b4a097329c37827fa4203782443ab1313ffa996a7b8fb4310ad1d86ea8e04de6190a77c2e44c11dc852994fe97c95fb0648a8f6bd5aecbc2baf8ec671644cc10eb40828836876b44c15e74bffe251fd28e0e9aa9dff031115de997d6226112380cbbee251bf060fdc6bf62b5526d506ba0ae480523bd3615ab96cd198;
    5'b00010 : xpb = 1024'h1277bb60d224b18abbead81d73aca8f715e022f729db8cd7f419cccba73860cd18c13f4a572879cdea23fc49c1d48f089511ce266e9f1d2f053a38f9244b1831544a4d6eb87f53c1be5365f592f2d3ced09f00b9354d282b48799031030858321d1ab4d7e6b4cc15f74c38d9e01c3080fed02e91c57da374313747b0e9f73cc5;
    5'b00011 : xpb = 1024'h740a3bbc1c2e24b47f630017b5b0211b598b360b2985237fad150fdc5455e7b7a6c61dabe7cff5fc2ee51a12146ddef211a7c92cb74813ec6026f524d3d9dea2b8970e7d6c877c4526ca1a41a8da1fceb2f0fde21636d2c9477ca146e1a1d594432bd858b273ae67b65248b64c125bd625a5354bd06223c66d0aa90ba3640e5d;
    5'b00100 : xpb = 1024'h24ef76c1a449631577d5b03ae75951ee2bc045ee53b719afe83399974e70c19a31827e94ae50f39bd447f89383a91e112a239c4cdd3e3a5e0a7471f248963062a8949add70fea7837ca6cbeb25e5a79da13e01726a9a505690f320620610b0643a3569afcd69982bee9871b3c0386101fda05d238afb46e8626e8f61d3ee798a;
    5'b00101 : xpb = 1024'h8681f71cee52d63f3b4dd835295cca126f6b59025360b057a12edca7fb8e4884bf875cf63ef86fca1909165bd6426dfaa6b9975325e7311b65612e1df824f6d40ce15bec2506d006e51d80373bccf39d838ffe9b4b83faf48ff63177e4aa2dc660468d3099287a7dad9e81902c2e8c57247563dd95dfc73a9e41f0bc8d5b4b22;
    5'b00110 : xpb = 1024'h37673222766e14a033c088585b05fae541a068e57d92a687dc4d6662f5a922674a43bddf05796d69be6bf4dd457dad19bf356a734bdd578d0faeaaeb6ce14893fcdee84c297dfb453afa31e0b8d87b6c71dd022b9fe77881d96cb0930919089657501e87b41e6441e5e4aa8da0549182fc708bb55078ea5c93a5d712bde5b64f;
    5'b00111 : xpb = 1024'h98f9b27dc07787c9f738b0529d097309854b7bf97d3c3d2f9548a973a2c6a951d8489c409620e998032d12a59816fd033bcb657994864e4a6a9b67171c700f05612ba95add8623c8a370e62ccebfc76c542eff5480d1231fd86fc1a8e7b285f87d6142087fdd4693a4eaba6a0c4abcd82345926f5b5d6aaecf79386d775287e7;
    5'b01000 : xpb = 1024'h49deed834892c62aefab6075ceb2a3dc57808bdca76e335fd067332e9ce183346304fd295ca1e737a88ff12707523c2254473899ba7c74bc14e8e3e4912c60c5512935bae1fd4f06f94d97d64bcb4f3b427c02e4d534a0ad21e640c40c2160c8746ad35f9ad33057dd30e3678070c203fb40ba4715f68dd0c4dd1ec3a7dcf314;
    5'b01001 : xpb = 1024'hab716dde929c3954b323887010b61c009b2b9ef0a717ca078962763f49ff0a1ef109db8aed496365ed510eef59eb8c0bd0dd33a003256b796fd5a01040bb2736b575f6c99605778a61c44c2261b29b3b24ce000db61e4b4b20e951d9eabade2a9a7bf6e0669212a99c36f343ec66ed592215c10120db0e2300b0801e6149c4ac;
    5'b01010 : xpb = 1024'h5c56a8e41ab777b5ab963893425f4cd36d60aed3d149c037c480fffa4419e4017bc63c73b3ca610592b3ed70c926cb2ae95906c0291b91eb1a231cddb57778f6a57383299a7ca2c8b7a0fdcbdebe230a131b039e0a81c8d86a5fd0f50f29b8fa918588378187fc6dd47d1c41608cf284fa10e8d8db743144f614667491d42fd9;
    5'b01011 : xpb = 1024'hd3be3e9a2d2b616a408e8b674087da63f95beb6fb7bb667ff9f89b53e34bde406829d5c7a4b5ea53816cbf238620a4a01d4d9e04f11b85cc47099ab2a33cab695710f899ef3ce070d7daf755bc9aad90168072e5ee54665b3d65010339893ca888f198e9c7de6320cc3453ed4b2f7b0d20c10b0960d5466eb784ccac25e9b06;
    5'b01100 : xpb = 1024'h6ece6444ecdc2940678110b0b60bf5ca8340d1cafb254d0fb89accc5eb5244ce94877bbe0af2dad37cd7e9ba8afb5a337e6ad4e697baaf1a1f5d55d6d9c29127f9bdd09852fbf68a75f463c171b0f6d8e3ba04573fcef103b2d961261232112caea03d0f683cc883cbc9551b40a92305f8e1176aa0f1d4b9274bae257bcb6c9e;
    5'b01101 : xpb = 1024'h1fb39f4a74f767a15ff3c0d3e7b5269d5575e1ae2557433ff3b95680e56d1eb11f43dca6d173d873223ac83bfa36995296e6a806bdb0d58bc9aad2a44e7ee2e7e9bb5cf8577321c8cbd1156aeebc7ea7d20707e794326e90fc4fe04136a0ebfca5a9ce668332b248040f7e18b4cf2831d0dc3f425b8af7db1caf947bac55d7cb;
    5'b01110 : xpb = 1024'h81461fa5bf00dacb236be8ce29b89ec19920f4c22500d9e7acb49991928aa59bad48bb08621b54a166fbe6044ccfe93c137ca30d0659cc4924978ecffe0da9594e081e070b7b4a4c3447c9b704a3caa7b4590510751c192efb52f157153a695ecbbaf1e74ef19499c3158df520c55386f7b145fc666f782d5882f5d665c2a963;
    5'b01111 : xpb = 1024'h322b5aab471c192c1bde98f15b61cf946b5604a54f32d017e7d3234c8ca57f7e38051bf1289c52410c5ec485bc0b285b2bf8762d2c4ff2bacee50b9d72c9fb193e05aa670ff2758a8a247b6081af5276a2a608a0c97f96bc44c9707239a9442ec2c4833e69e77e5dfb5bb6f294eb58b2cfac6dd421089b4f4de6dc2c964d1490;
    5'b10000 : xpb = 1024'h93bddb0691258c55df56c0eb9d6547b8af0117b94edc66bfa0ce665d39c30668c609fa52b943ce6f511fe24e0ea47844a88e713374f8e97829d1c7c92258c18aa2526b75c3fa9e0df29b2fac97969e7684f805c9aa69415a43cc81881842c190e8d5a6bf35a660afba61c6cf00e18407f681748e2bed1ba189ba3d874fb9e628;
    5'b10001 : xpb = 1024'h44a3160c1940cab6d7c9710ecf0e788b8136279c790e5cefdbecf01833dde04b50c65b3b7fc4cc0ef682c0cf7ddfb763c10a44539aef0fe9d41f44969715134a924ff7d5c871c94c4877e15614a2264573450959feccbee78d4300a33cb19c60dfdf3816509c4a73f2a7efcc75078933ce7c9c65e6863ec37f1e23dd80445155;
    5'b10010 : xpb = 1024'ha6359667634a3de09b4199091111f0afc4e13ab078b7f39794e83328e0fb6735decb399d106c483d3b43de97d079074d3da03f59e39806a72f0c00c246a3d9bbf69cb8e47c79f1cfb0ee95a22a89724555970682dfb669858c4611b91b4b19c305f05b971c5b2cc5b1adffa8e0fdb488f551a31ff16abf15baf1853839b122ed;
    5'b10011 : xpb = 1024'h571ad16ceb657c4193b4492c42bb218297164a93a2e9e9c7d006bce3db16411869879a85d6ed45dce0a6bd193fb4466c561c127a098e2d18d9597d8fbb602b7be69a454480f11d0e06cb474ba794fa1443e40a133419e712d5bc90d43fb9f492fcf9ecee37511689e9f428a65523b9b4cd4ccaf7ac03e237b0556b8e6a3b8e1a;
    5'b10100 : xpb = 1024'h8000c727380baa28c26f94f74645255694b5a76cd1bdff80b25469ed5311afaf443fb6e9d6e437c86099b9aaeef858b6e97e59a2f84538a83a6fa5d301c7d3bd697d1a48568484c5ca7f8f524a081e332310da3887d64a01f330fef6428cf62f4037e455247004e223a51a3c949bee0a547f2cf669d0559a5b951e49ac5f947;
    5'b10101 : xpb = 1024'h69928ccdbd8a2dcc4f9f2149b667ca79acf66d8accc5769fc42089af824ea1e58248d9d02e15bfaacacab9630188d574eb2de0a0782d4a47de93b688dfab43ad3ae492b3397070cfc51ead413a87cde314830acc69670f3e1e36210542c24cc51a14a1c61e05e29fe1406180353fea35cc1cf989718185abe18cb33f5432cadf;
    5'b10110 : xpb = 1024'h1a77c7d345a56c2d4811d16ce810fb4c7f2b7d6df6f76ccfff3f136a7c697bc80d053ab8f496bd4a702d97e470c4149403a9b3c09e2370b988e133565467956d2ae21f133de79c0e1afb5eeab79355b202d00e5cbdca8ccb67aca02067312795111e331d38fbcc6419868a7da965ef61a41821612c1aa8cdd6f0999584bd360c;
    5'b10111 : xpb = 1024'h7c0a482e8faedf570b89f9672a147370c2d69081f6a10377b83a567b298702b29b0a191a853e3978b4eeb5acc35d647d803faec6e6cc6776e3cdef8203f65bde8f2ee021f1efc49183721336cd7aa1b1e5220b859eb4376966afb13645caa4f7372f569e04baaeb5d88c9a5a155c1ab6caed281b36ff292012c3faf03e2a07a4;
    5'b11000 : xpb = 1024'h2cef833417ca1db803fca98a5bbda443950ba06520d2f9a7f358e03623a1dc9525c67a034bbf37185a51942e3298a39c98bb81e70cc28de88e1b6c4f78b2ad9e7f2c6c81f666efcfd94ec4e04a862980d36f0f15f317b4f6b02630516a397fc72e38e7f51fb0987a10d2c35789821fe2a2e84ff2f1984c420827e1466eb472d1;
    5'b11001 : xpb = 1024'h8e82038f61d390e1c774d1849dc11c67d8b6b379207c904fac542346d0bf637fb3cb5864dc66b3469f12b1f68531f38615517ced556b84a5e908287b2841740fe3792d90aa6f185341c5792c606d7580b5c10c3ed4015f94af29416748d2fd29544a0b75eb6f7acbcfd8d333f5784b37c9bd56acfc7ccc9443fb42a128214469;
    5'b11010 : xpb = 1024'h3f673e94e9eecf42bfe781a7cf6a4d3aaaebc35c4aae867fe772ad01cada3d623e87b94da2e7b0e644759077f46d32a52dcd500d7b61ab179355a5489cfdc5cfd376b9f0aee6439197a22ad5dd78fd4fa40e0fcf2864dd21f89fc0826d41d7f94b539ccd06656490081efc31699e5063a1b87e84b715efb6395f28f758abaf96;
    5'b11011 : xpb = 1024'ha0f9bef033f8426c835fa9a2116dc55eee96d6704a581d27a06df01277f7c44ccc8c97af338f2d148936ae404706828eaa634b13c40aa1d4ee4261744c8c8c4137c37aff62ee6c150018df21f360494f86600cf8094e87bff7a2d1984bdb555b7164c04dd22446e1c7250c0dd5947bb8c88d853ec1fa700875328a521218812e;
    5'b11100 : xpb = 1024'h51def9f5bc1380cd7bd259c54316f631c0cbe653748a1357db8c79cd72129e2f5748f897fa102ab42e998cc1b641c1adc2df1e33ea00c846988fde41c148de0127c1075f6765975355f590cb706bd11e74ad10885db2054d411950b3704a302b686e51a4ed1a30a5ff6b350b49ba80e4a088ad167c93932a6a9670a842a2ec5b;
    5'b11101 : xpb = 1024'h2c434fb442ebf2e744509e874c027049300f6369ebc098816ab03886c2d7811e2055980c0912853d3fc6b43257d00ccdb5af1540ff6eeb842dd5b0f36052fc117be93bf6bdcc291abd24274ed7758ed62fa1418b21582da8a8fcfce94b90afb5f77e2fc08101a6a37b15e08bde086107883d4ee372cb64c5ffa56fe732d5788;
    5'b11110 : xpb = 1024'h6456b5568e38325837bd31e2b6c39f28d6ac094a9e65a02fcfa64699194afefc700a37e25138a48218bd890b781650b657f0ec5a589fe5759dca173ae593f6327c0b54ce1fe4eb151448f6c1035ea4ed454c114192ff2d788992e0e47352885d8589067cd3cefcbbf6b76de529d6b1659f58dba84211369e9bcdb8592c9a2920;
    5'b11111 : xpb = 1024'h153bf05c165370b9302fe205e86ccffba8e1192dc89796600ac4d0541365d8defac698cb17b9a221be20678ce7518fd5706cbf7a7e960be7481794085a5047f26c08e12e245c16536a25a86a806a2cbc339914d1e762ab05d3095fff97c1632d7c9297d3eec4e6802efd96e29dfcb6917754037ffcaa59c091319eaf5d24944d;
    endcase
end

endmodule
